module basic_3000_30000_3500_5_levels_10xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
nor U0 (N_0,In_1513,In_1550);
xor U1 (N_1,In_1510,In_560);
xor U2 (N_2,In_838,In_728);
and U3 (N_3,In_1314,In_1516);
or U4 (N_4,In_247,In_253);
or U5 (N_5,In_305,In_2218);
and U6 (N_6,In_1745,In_941);
nand U7 (N_7,In_580,In_1764);
nand U8 (N_8,In_2708,In_2827);
or U9 (N_9,In_1208,In_2257);
or U10 (N_10,In_2361,In_943);
or U11 (N_11,In_2058,In_343);
xnor U12 (N_12,In_1055,In_1290);
and U13 (N_13,In_1413,In_2598);
or U14 (N_14,In_868,In_2302);
nor U15 (N_15,In_0,In_2737);
xnor U16 (N_16,In_197,In_1593);
or U17 (N_17,In_1634,In_2146);
xnor U18 (N_18,In_1303,In_2926);
xor U19 (N_19,In_1825,In_1313);
nand U20 (N_20,In_1261,In_1424);
or U21 (N_21,In_2605,In_1352);
or U22 (N_22,In_1657,In_1796);
xor U23 (N_23,In_2213,In_427);
nand U24 (N_24,In_2687,In_1875);
nand U25 (N_25,In_2662,In_2534);
and U26 (N_26,In_3,In_526);
xor U27 (N_27,In_1073,In_1220);
nor U28 (N_28,In_1039,In_658);
nand U29 (N_29,In_830,In_2616);
and U30 (N_30,In_2289,In_726);
and U31 (N_31,In_897,In_249);
nand U32 (N_32,In_2159,In_1431);
xor U33 (N_33,In_2970,In_1536);
xnor U34 (N_34,In_1756,In_11);
xnor U35 (N_35,In_113,In_2593);
xor U36 (N_36,In_2535,In_736);
and U37 (N_37,In_956,In_255);
xnor U38 (N_38,In_1082,In_2626);
nand U39 (N_39,In_898,In_511);
or U40 (N_40,In_2176,In_2823);
or U41 (N_41,In_1471,In_2793);
or U42 (N_42,In_288,In_1125);
nand U43 (N_43,In_2814,In_317);
nor U44 (N_44,In_2460,In_1839);
or U45 (N_45,In_124,In_1722);
xor U46 (N_46,In_1395,In_1211);
nand U47 (N_47,In_91,In_592);
and U48 (N_48,In_1924,In_1305);
or U49 (N_49,In_2850,In_949);
or U50 (N_50,In_1723,In_424);
nor U51 (N_51,In_1246,In_496);
nand U52 (N_52,In_2647,In_1575);
or U53 (N_53,In_2606,In_2990);
nor U54 (N_54,In_2147,In_2009);
xnor U55 (N_55,In_2420,In_1587);
xor U56 (N_56,In_1249,In_1870);
nand U57 (N_57,In_800,In_14);
xnor U58 (N_58,In_811,In_2490);
nand U59 (N_59,In_2114,In_1886);
or U60 (N_60,In_1002,In_2689);
and U61 (N_61,In_51,In_2199);
nand U62 (N_62,In_1772,In_2017);
and U63 (N_63,In_1613,In_1411);
and U64 (N_64,In_1243,In_1770);
nand U65 (N_65,In_2193,In_1298);
nor U66 (N_66,In_660,In_2237);
nand U67 (N_67,In_613,In_1444);
nand U68 (N_68,In_222,In_1708);
or U69 (N_69,In_326,In_2056);
nand U70 (N_70,In_1336,In_1891);
nor U71 (N_71,In_1646,In_40);
or U72 (N_72,In_643,In_873);
or U73 (N_73,In_2346,In_1675);
and U74 (N_74,In_1087,In_1052);
and U75 (N_75,In_246,In_1691);
nor U76 (N_76,In_2542,In_2818);
xor U77 (N_77,In_2697,In_1136);
nand U78 (N_78,In_262,In_667);
nor U79 (N_79,In_54,In_1761);
or U80 (N_80,In_2249,In_2919);
nand U81 (N_81,In_886,In_2196);
or U82 (N_82,In_2885,In_1752);
xnor U83 (N_83,In_1194,In_703);
xnor U84 (N_84,In_1012,In_1470);
xor U85 (N_85,In_1110,In_1973);
xor U86 (N_86,In_2393,In_2841);
nand U87 (N_87,In_1578,In_21);
and U88 (N_88,In_152,In_2933);
nand U89 (N_89,In_2894,In_2281);
nor U90 (N_90,In_2629,In_77);
xnor U91 (N_91,In_2145,In_2504);
nand U92 (N_92,In_745,In_2773);
nor U93 (N_93,In_2117,In_334);
nand U94 (N_94,In_1784,In_2011);
or U95 (N_95,In_1715,In_2044);
xnor U96 (N_96,In_1416,In_976);
or U97 (N_97,In_2825,In_2955);
nor U98 (N_98,In_1589,In_1455);
nand U99 (N_99,In_1522,In_944);
nand U100 (N_100,In_1938,In_7);
xor U101 (N_101,In_2931,In_2268);
or U102 (N_102,In_1822,In_2619);
nor U103 (N_103,In_555,In_2135);
and U104 (N_104,In_1275,In_1096);
nor U105 (N_105,In_686,In_1504);
and U106 (N_106,In_286,In_2751);
nand U107 (N_107,In_1692,In_1677);
xnor U108 (N_108,In_1913,In_1626);
nor U109 (N_109,In_2803,In_2958);
nor U110 (N_110,In_1320,In_664);
xnor U111 (N_111,In_1928,In_1563);
or U112 (N_112,In_1771,In_2184);
nor U113 (N_113,In_307,In_639);
or U114 (N_114,In_623,In_2726);
and U115 (N_115,In_1454,In_1531);
nor U116 (N_116,In_965,In_423);
nand U117 (N_117,In_2764,In_236);
xor U118 (N_118,In_376,In_488);
nor U119 (N_119,In_596,In_49);
xnor U120 (N_120,In_2916,In_2585);
and U121 (N_121,In_781,In_672);
or U122 (N_122,In_599,In_1155);
nor U123 (N_123,In_707,In_2506);
xor U124 (N_124,In_1994,In_1307);
xor U125 (N_125,In_1453,In_2941);
nor U126 (N_126,In_2630,In_150);
and U127 (N_127,In_1890,In_2602);
xnor U128 (N_128,In_640,In_1193);
nand U129 (N_129,In_125,In_2376);
xor U130 (N_130,In_335,In_1366);
and U131 (N_131,In_2701,In_2334);
and U132 (N_132,In_401,In_1739);
nor U133 (N_133,In_1241,In_86);
nand U134 (N_134,In_244,In_950);
nand U135 (N_135,In_2712,In_2705);
xnor U136 (N_136,In_1250,In_922);
nor U137 (N_137,In_1067,In_1909);
nand U138 (N_138,In_2095,In_1607);
and U139 (N_139,In_2144,In_448);
xnor U140 (N_140,In_2576,In_12);
or U141 (N_141,In_2997,In_2062);
and U142 (N_142,In_2731,In_2978);
nor U143 (N_143,In_2473,In_1548);
nand U144 (N_144,In_280,In_1980);
xnor U145 (N_145,In_1623,In_2465);
nor U146 (N_146,In_2462,In_2696);
nor U147 (N_147,In_918,In_777);
or U148 (N_148,In_2076,In_1596);
nand U149 (N_149,In_1640,In_95);
xnor U150 (N_150,In_2533,In_224);
nand U151 (N_151,In_1285,In_73);
and U152 (N_152,In_2142,In_386);
nand U153 (N_153,In_827,In_768);
or U154 (N_154,In_2020,In_722);
nor U155 (N_155,In_499,In_2022);
nand U156 (N_156,In_899,In_1779);
nand U157 (N_157,In_1889,In_157);
and U158 (N_158,In_158,In_149);
xnor U159 (N_159,In_2546,In_131);
and U160 (N_160,In_2620,In_2522);
or U161 (N_161,In_1406,In_9);
xnor U162 (N_162,In_318,In_2496);
xor U163 (N_163,In_1789,In_230);
and U164 (N_164,In_85,In_2852);
and U165 (N_165,In_2792,In_558);
nor U166 (N_166,In_1074,In_2577);
and U167 (N_167,In_1355,In_215);
or U168 (N_168,In_1731,In_2758);
xnor U169 (N_169,In_702,In_2010);
xnor U170 (N_170,In_10,In_2036);
or U171 (N_171,In_544,In_2956);
nor U172 (N_172,In_1714,In_986);
nor U173 (N_173,In_1242,In_2952);
nor U174 (N_174,In_2458,In_1793);
or U175 (N_175,In_1521,In_1378);
nor U176 (N_176,In_2643,In_1166);
nor U177 (N_177,In_2007,In_2944);
nor U178 (N_178,In_104,In_1642);
or U179 (N_179,In_1868,In_48);
nor U180 (N_180,In_2560,In_931);
and U181 (N_181,In_1008,In_62);
and U182 (N_182,In_1011,In_618);
xnor U183 (N_183,In_470,In_2962);
or U184 (N_184,In_446,In_2069);
and U185 (N_185,In_2452,In_2075);
xnor U186 (N_186,In_2876,In_2536);
nand U187 (N_187,In_1168,In_795);
and U188 (N_188,In_1051,In_1629);
nor U189 (N_189,In_1617,In_2946);
and U190 (N_190,In_2703,In_2345);
nand U191 (N_191,In_1173,In_2426);
or U192 (N_192,In_1600,In_1740);
nand U193 (N_193,In_138,In_1702);
and U194 (N_194,In_274,In_539);
xnor U195 (N_195,In_1765,In_1530);
and U196 (N_196,In_507,In_1376);
and U197 (N_197,In_1143,In_2693);
nand U198 (N_198,In_1729,In_1983);
nor U199 (N_199,In_1674,In_110);
xnor U200 (N_200,In_1511,In_506);
xnor U201 (N_201,In_1207,In_1092);
nand U202 (N_202,In_1351,In_2544);
nand U203 (N_203,In_1997,In_2263);
and U204 (N_204,In_2736,In_715);
or U205 (N_205,In_1018,In_1651);
and U206 (N_206,In_2296,In_2810);
and U207 (N_207,In_2405,In_2617);
or U208 (N_208,In_2255,In_1703);
or U209 (N_209,In_1641,In_1614);
or U210 (N_210,In_142,In_2812);
and U211 (N_211,In_2379,In_2949);
and U212 (N_212,In_2867,In_2053);
and U213 (N_213,In_2206,In_2692);
or U214 (N_214,In_2203,In_1775);
xor U215 (N_215,In_2511,In_609);
xor U216 (N_216,In_2644,In_2101);
nand U217 (N_217,In_282,In_1016);
and U218 (N_218,In_1673,In_537);
or U219 (N_219,In_778,In_1618);
and U220 (N_220,In_1262,In_1192);
xor U221 (N_221,In_2648,In_835);
nand U222 (N_222,In_155,In_129);
xnor U223 (N_223,In_2864,In_1140);
nor U224 (N_224,In_240,In_354);
and U225 (N_225,In_1517,In_2344);
and U226 (N_226,In_2514,In_1068);
or U227 (N_227,In_2125,In_101);
or U228 (N_228,In_2640,In_2702);
and U229 (N_229,In_605,In_2776);
or U230 (N_230,In_1121,In_1495);
or U231 (N_231,In_2813,In_2719);
nand U232 (N_232,In_58,In_2500);
nor U233 (N_233,In_1217,In_826);
nand U234 (N_234,In_1482,In_1337);
nand U235 (N_235,In_718,In_1007);
or U236 (N_236,In_591,In_2043);
nand U237 (N_237,In_1633,In_531);
nor U238 (N_238,In_289,In_198);
xor U239 (N_239,In_2898,In_72);
nor U240 (N_240,In_571,In_2267);
nor U241 (N_241,In_1823,In_2594);
or U242 (N_242,In_2110,In_491);
and U243 (N_243,In_2408,In_996);
and U244 (N_244,In_251,In_457);
and U245 (N_245,In_1299,In_349);
or U246 (N_246,In_393,In_1499);
or U247 (N_247,In_787,In_775);
nand U248 (N_248,In_2655,In_1929);
and U249 (N_249,In_2055,In_663);
xnor U250 (N_250,In_1735,In_1390);
nand U251 (N_251,In_2632,In_1995);
nand U252 (N_252,In_375,In_2323);
nor U253 (N_253,In_476,In_202);
and U254 (N_254,In_487,In_254);
xnor U255 (N_255,In_1345,In_1106);
xor U256 (N_256,In_1577,In_1969);
nand U257 (N_257,In_720,In_1515);
and U258 (N_258,In_2651,In_1635);
or U259 (N_259,In_2637,In_2189);
or U260 (N_260,In_1377,In_2113);
or U261 (N_261,In_2437,In_2066);
and U262 (N_262,In_512,In_700);
or U263 (N_263,In_1781,In_2634);
xnor U264 (N_264,In_1152,In_2492);
nand U265 (N_265,In_422,In_1724);
nor U266 (N_266,In_2188,In_189);
nor U267 (N_267,In_352,In_1429);
xor U268 (N_268,In_813,In_1230);
nor U269 (N_269,In_2080,In_1503);
nand U270 (N_270,In_1410,In_1976);
and U271 (N_271,In_2133,In_2204);
xnor U272 (N_272,In_415,In_887);
or U273 (N_273,In_2327,In_547);
nand U274 (N_274,In_1458,In_486);
or U275 (N_275,In_2318,In_2192);
and U276 (N_276,In_1947,In_2815);
or U277 (N_277,In_801,In_834);
or U278 (N_278,In_1120,In_2603);
xor U279 (N_279,In_662,In_1292);
nor U280 (N_280,In_2720,In_2555);
or U281 (N_281,In_2895,In_540);
and U282 (N_282,In_1857,In_1310);
nor U283 (N_283,In_2012,In_2412);
or U284 (N_284,In_167,In_1170);
nand U285 (N_285,In_859,In_1196);
or U286 (N_286,In_959,In_1525);
or U287 (N_287,In_2982,In_143);
nor U288 (N_288,In_481,In_56);
or U289 (N_289,In_2586,In_2312);
or U290 (N_290,In_2609,In_2183);
or U291 (N_291,In_2964,In_1260);
nand U292 (N_292,In_2856,In_213);
nand U293 (N_293,In_862,In_2097);
and U294 (N_294,In_1697,In_709);
xor U295 (N_295,In_2911,In_1716);
nand U296 (N_296,In_2171,In_1738);
nor U297 (N_297,In_769,In_1960);
xnor U298 (N_298,In_2879,In_1043);
and U299 (N_299,In_353,In_177);
xor U300 (N_300,In_2155,In_1028);
or U301 (N_301,In_1165,In_2399);
xnor U302 (N_302,In_1887,In_372);
xnor U303 (N_303,In_206,In_1894);
nand U304 (N_304,In_1428,In_2759);
nor U305 (N_305,In_443,In_130);
xnor U306 (N_306,In_477,In_1900);
nor U307 (N_307,In_688,In_340);
xnor U308 (N_308,In_1189,In_1034);
nand U309 (N_309,In_2805,In_1943);
or U310 (N_310,In_2025,In_1149);
xor U311 (N_311,In_562,In_2513);
nand U312 (N_312,In_2178,In_2461);
and U313 (N_313,In_863,In_2571);
nand U314 (N_314,In_2407,In_2435);
or U315 (N_315,In_2633,In_2034);
nor U316 (N_316,In_2175,In_1780);
or U317 (N_317,In_882,In_1477);
nor U318 (N_318,In_1999,In_2148);
or U319 (N_319,In_2367,In_2356);
and U320 (N_320,In_2967,In_2423);
xnor U321 (N_321,In_2625,In_1726);
or U322 (N_322,In_679,In_2851);
xnor U323 (N_323,In_611,In_88);
and U324 (N_324,In_2454,In_193);
or U325 (N_325,In_1331,In_1583);
nand U326 (N_326,In_840,In_930);
xor U327 (N_327,In_2671,In_2768);
xnor U328 (N_328,In_2270,In_1302);
or U329 (N_329,In_273,In_28);
nand U330 (N_330,In_265,In_128);
and U331 (N_331,In_1683,In_2049);
xor U332 (N_332,In_758,In_502);
and U333 (N_333,In_2516,In_2953);
nor U334 (N_334,In_2992,In_2357);
and U335 (N_335,In_1667,In_1636);
xnor U336 (N_336,In_226,In_824);
nand U337 (N_337,In_955,In_1088);
and U338 (N_338,In_2313,In_2364);
or U339 (N_339,In_543,In_1599);
nand U340 (N_340,In_1218,In_1013);
nand U341 (N_341,In_103,In_704);
nand U342 (N_342,In_1371,In_348);
or U343 (N_343,In_2284,In_1743);
nor U344 (N_344,In_1417,In_2433);
or U345 (N_345,In_1758,In_964);
and U346 (N_346,In_379,In_825);
and U347 (N_347,In_2559,In_362);
nor U348 (N_348,In_1541,In_1812);
or U349 (N_349,In_430,In_2891);
and U350 (N_350,In_2241,In_84);
nor U351 (N_351,In_1508,In_1151);
or U352 (N_352,In_2439,In_1278);
xor U353 (N_353,In_1274,In_1658);
xnor U354 (N_354,In_2524,In_1233);
nor U355 (N_355,In_2561,In_593);
nor U356 (N_356,In_1546,In_313);
xnor U357 (N_357,In_214,In_2467);
or U358 (N_358,In_2607,In_856);
xnor U359 (N_359,In_2021,In_1236);
nand U360 (N_360,In_1325,In_1344);
nand U361 (N_361,In_65,In_929);
and U362 (N_362,In_920,In_875);
xor U363 (N_363,In_935,In_550);
nor U364 (N_364,In_2920,In_2304);
nor U365 (N_365,In_391,In_404);
nor U366 (N_366,In_2786,In_2324);
nand U367 (N_367,In_2610,In_139);
xor U368 (N_368,In_2569,In_1904);
nor U369 (N_369,In_2556,In_2591);
xnor U370 (N_370,In_1685,In_678);
and U371 (N_371,In_1256,In_2710);
or U372 (N_372,In_2120,In_2590);
or U373 (N_373,In_1644,In_1339);
nor U374 (N_374,In_2652,In_1954);
nor U375 (N_375,In_16,In_2972);
and U376 (N_376,In_2691,In_1671);
nand U377 (N_377,In_2169,In_432);
nand U378 (N_378,In_154,In_751);
and U379 (N_379,In_2498,In_2086);
nor U380 (N_380,In_2711,In_140);
nor U381 (N_381,In_2440,In_1252);
or U382 (N_382,In_1836,In_219);
nor U383 (N_383,In_1549,In_1277);
and U384 (N_384,In_480,In_1528);
nor U385 (N_385,In_1112,In_2830);
or U386 (N_386,In_1266,In_1681);
or U387 (N_387,In_2503,In_153);
nor U388 (N_388,In_536,In_1203);
nand U389 (N_389,In_1888,In_932);
nor U390 (N_390,In_2520,In_2352);
and U391 (N_391,In_2019,In_2874);
and U392 (N_392,In_817,In_630);
or U393 (N_393,In_1996,In_1713);
and U394 (N_394,In_1267,In_2116);
or U395 (N_395,In_2382,In_854);
or U396 (N_396,In_1844,In_1966);
and U397 (N_397,In_2293,In_1442);
xor U398 (N_398,In_2817,In_2787);
nand U399 (N_399,In_59,In_2550);
nor U400 (N_400,In_2948,In_97);
nor U401 (N_401,In_1806,In_1534);
and U402 (N_402,In_585,In_1782);
nor U403 (N_403,In_576,In_269);
xor U404 (N_404,In_1127,In_2589);
xor U405 (N_405,In_2917,In_2163);
nor U406 (N_406,In_2247,In_2713);
xor U407 (N_407,In_29,In_1209);
and U408 (N_408,In_2543,In_2799);
nand U409 (N_409,In_2238,In_564);
or U410 (N_410,In_1676,In_275);
or U411 (N_411,In_620,In_1926);
or U412 (N_412,In_44,In_1461);
or U413 (N_413,In_1955,In_2409);
and U414 (N_414,In_1554,In_1361);
nor U415 (N_415,In_2774,In_79);
and U416 (N_416,In_242,In_1711);
nand U417 (N_417,In_1319,In_2686);
or U418 (N_418,In_2051,In_896);
nor U419 (N_419,In_1650,In_463);
and U420 (N_420,In_610,In_1750);
nor U421 (N_421,In_2777,In_2548);
and U422 (N_422,In_1403,In_1059);
nor U423 (N_423,In_78,In_199);
xor U424 (N_424,In_697,In_594);
nor U425 (N_425,In_951,In_631);
nor U426 (N_426,In_773,In_2057);
nor U427 (N_427,In_1200,In_1419);
or U428 (N_428,In_1912,In_1443);
nor U429 (N_429,In_2979,In_2477);
or U430 (N_430,In_992,In_1359);
nor U431 (N_431,In_2807,In_1348);
nand U432 (N_432,In_760,In_165);
and U433 (N_433,In_985,In_1391);
and U434 (N_434,In_1690,In_1965);
or U435 (N_435,In_181,In_2210);
nand U436 (N_436,In_1672,In_1038);
and U437 (N_437,In_2838,In_2384);
nor U438 (N_438,In_126,In_441);
xor U439 (N_439,In_2960,In_2694);
nor U440 (N_440,In_2714,In_687);
or U441 (N_441,In_1452,In_708);
nand U442 (N_442,In_98,In_319);
nor U443 (N_443,In_1769,In_1434);
xor U444 (N_444,In_802,In_1078);
and U445 (N_445,In_1591,In_2578);
nand U446 (N_446,In_519,In_2123);
nand U447 (N_447,In_2672,In_64);
xnor U448 (N_448,In_2680,In_1160);
nand U449 (N_449,In_798,In_2604);
or U450 (N_450,In_1478,In_2179);
and U451 (N_451,In_122,In_363);
xor U452 (N_452,In_294,In_2674);
nor U453 (N_453,In_1879,In_1786);
nor U454 (N_454,In_18,In_1400);
xnor U455 (N_455,In_1062,In_2936);
and U456 (N_456,In_257,In_1925);
nor U457 (N_457,In_1688,In_2928);
or U458 (N_458,In_434,In_946);
or U459 (N_459,In_1834,In_654);
or U460 (N_460,In_2568,In_1485);
nor U461 (N_461,In_1540,In_622);
xor U462 (N_462,In_426,In_2305);
xor U463 (N_463,In_2715,In_350);
and U464 (N_464,In_2580,In_948);
or U465 (N_465,In_192,In_1315);
and U466 (N_466,In_1229,In_115);
nor U467 (N_467,In_32,In_2657);
nor U468 (N_468,In_998,In_2761);
and U469 (N_469,In_2762,In_1512);
nor U470 (N_470,In_1820,In_1179);
nor U471 (N_471,In_1579,In_2613);
nand U472 (N_472,In_2654,In_180);
and U473 (N_473,In_1831,In_1104);
xor U474 (N_474,In_2042,In_2753);
nand U475 (N_475,In_1340,In_1223);
or U476 (N_476,In_2747,In_1214);
nor U477 (N_477,In_1718,In_1412);
xnor U478 (N_478,In_732,In_1655);
xnor U479 (N_479,In_2728,In_680);
xnor U480 (N_480,In_1956,In_171);
or U481 (N_481,In_923,In_2325);
xor U482 (N_482,In_1805,In_2093);
xor U483 (N_483,In_883,In_2028);
xor U484 (N_484,In_1464,In_1474);
nor U485 (N_485,In_528,In_2174);
xor U486 (N_486,In_1754,In_1353);
and U487 (N_487,In_435,In_1896);
and U488 (N_488,In_1154,In_2908);
nor U489 (N_489,In_2089,In_2235);
xor U490 (N_490,In_1430,In_478);
nor U491 (N_491,In_2214,In_2314);
and U492 (N_492,In_1505,In_111);
and U493 (N_493,In_845,In_2781);
or U494 (N_494,In_1864,In_1163);
nor U495 (N_495,In_1115,In_2226);
or U496 (N_496,In_2763,In_1818);
or U497 (N_497,In_2310,In_1952);
and U498 (N_498,In_1379,In_892);
nor U499 (N_499,In_1066,In_979);
nor U500 (N_500,In_261,In_2000);
nand U501 (N_501,In_2748,In_1021);
or U502 (N_502,In_1309,In_232);
and U503 (N_503,In_617,In_2912);
and U504 (N_504,In_2868,In_1342);
xnor U505 (N_505,In_351,In_1553);
and U506 (N_506,In_1847,In_2765);
nand U507 (N_507,In_1659,In_990);
and U508 (N_508,In_548,In_2538);
and U509 (N_509,In_2315,In_727);
or U510 (N_510,In_2347,In_556);
nand U511 (N_511,In_200,In_1418);
and U512 (N_512,In_604,In_2351);
xor U513 (N_513,In_803,In_2645);
xor U514 (N_514,In_974,In_2008);
nor U515 (N_515,In_2295,In_1948);
and U516 (N_516,In_1961,In_619);
or U517 (N_517,In_2921,In_2037);
nor U518 (N_518,In_2261,In_1145);
or U519 (N_519,In_316,In_670);
or U520 (N_520,In_47,In_2635);
and U521 (N_521,In_1897,In_302);
nor U522 (N_522,In_1374,In_1524);
and U523 (N_523,In_2493,In_681);
and U524 (N_524,In_1272,In_523);
nand U525 (N_525,In_233,In_632);
xnor U526 (N_526,In_1584,In_2222);
or U527 (N_527,In_628,In_1649);
or U528 (N_528,In_1547,In_852);
or U529 (N_529,In_926,In_2137);
or U530 (N_530,In_1380,In_2592);
nand U531 (N_531,In_1821,In_2839);
and U532 (N_532,In_2335,In_1354);
and U533 (N_533,In_2115,In_1138);
or U534 (N_534,In_169,In_1562);
or U535 (N_535,In_2170,In_2515);
and U536 (N_536,In_2986,In_2269);
xor U537 (N_537,In_649,In_1005);
nor U538 (N_538,In_1235,In_2355);
or U539 (N_539,In_116,In_1231);
nand U540 (N_540,In_2227,In_2622);
or U541 (N_541,In_276,In_2965);
nor U542 (N_542,In_2678,In_1829);
xnor U543 (N_543,In_497,In_1433);
or U544 (N_544,In_2079,In_38);
or U545 (N_545,In_2366,In_541);
nand U546 (N_546,In_2182,In_1874);
xnor U547 (N_547,In_398,In_1393);
xor U548 (N_548,In_2052,In_508);
and U549 (N_549,In_2618,In_2299);
nor U550 (N_550,In_1945,In_1284);
and U551 (N_551,In_2861,In_382);
nor U552 (N_552,In_2734,In_1798);
nor U553 (N_553,In_2280,In_2158);
nand U554 (N_554,In_1114,In_1244);
nor U555 (N_555,In_1389,In_1286);
or U556 (N_556,In_1604,In_2784);
nand U557 (N_557,In_1245,In_1157);
or U558 (N_558,In_2862,In_2451);
or U559 (N_559,In_381,In_2273);
nand U560 (N_560,In_2326,In_2939);
and U561 (N_561,In_1367,In_1265);
or U562 (N_562,In_2893,In_2400);
xor U563 (N_563,In_2470,In_2285);
nor U564 (N_564,In_1071,In_1279);
nand U565 (N_565,In_1060,In_1526);
nor U566 (N_566,In_212,In_809);
or U567 (N_567,In_2664,In_993);
and U568 (N_568,In_2670,In_2478);
or U569 (N_569,In_2425,In_172);
or U570 (N_570,In_35,In_1150);
or U571 (N_571,In_2201,In_1437);
nor U572 (N_572,In_2725,In_754);
nor U573 (N_573,In_1970,In_495);
nand U574 (N_574,In_2389,In_1282);
and U575 (N_575,In_2221,In_1757);
nor U576 (N_576,In_2291,In_1533);
nor U577 (N_577,In_2195,In_2029);
or U578 (N_578,In_1122,In_1491);
nor U579 (N_579,In_960,In_2700);
xor U580 (N_580,In_962,In_2368);
nand U581 (N_581,In_1807,In_2574);
nor U582 (N_582,In_2730,In_1527);
xor U583 (N_583,In_529,In_615);
xor U584 (N_584,In_2649,In_1594);
nand U585 (N_585,In_494,In_2845);
or U586 (N_586,In_2450,In_321);
and U587 (N_587,In_1422,In_2338);
and U588 (N_588,In_119,In_743);
nand U589 (N_589,In_304,In_1105);
nor U590 (N_590,In_1932,In_2475);
nor U591 (N_591,In_2716,In_2139);
nor U592 (N_592,In_952,In_501);
xor U593 (N_593,In_1234,In_1777);
xnor U594 (N_594,In_1202,In_2416);
or U595 (N_595,In_339,In_565);
and U596 (N_596,In_2378,In_2871);
nor U597 (N_597,In_1085,In_2468);
nand U598 (N_598,In_1027,In_2834);
nand U599 (N_599,In_186,In_739);
nand U600 (N_600,In_1680,In_1656);
or U601 (N_601,In_1388,In_2775);
and U602 (N_602,In_575,In_1449);
or U603 (N_603,In_1029,In_1438);
nor U604 (N_604,In_790,In_553);
nor U605 (N_605,In_936,In_413);
nand U606 (N_606,In_1975,In_1832);
nand U607 (N_607,In_1281,In_2031);
and U608 (N_608,In_2596,In_1480);
nand U609 (N_609,In_2428,In_2039);
and U610 (N_610,In_2092,In_1564);
and U611 (N_611,In_1321,In_2077);
or U612 (N_612,In_2488,In_1025);
or U613 (N_613,In_2530,In_2112);
and U614 (N_614,In_1463,In_2791);
and U615 (N_615,In_2721,In_1301);
and U616 (N_616,In_2211,In_1210);
nand U617 (N_617,In_2394,In_1920);
and U618 (N_618,In_823,In_600);
or U619 (N_619,In_2336,In_2790);
and U620 (N_620,In_650,In_484);
nor U621 (N_621,In_939,In_2745);
xnor U622 (N_622,In_2003,In_641);
nand U623 (N_623,In_668,In_412);
and U624 (N_624,In_2185,In_42);
nor U625 (N_625,In_2527,In_2554);
nor U626 (N_626,In_730,In_1091);
xnor U627 (N_627,In_1985,In_1364);
or U628 (N_628,In_1381,In_1270);
nor U629 (N_629,In_89,In_2989);
and U630 (N_630,In_1989,In_2024);
nor U631 (N_631,In_2341,In_1332);
or U632 (N_632,In_1964,In_1863);
xor U633 (N_633,In_1686,In_2563);
nand U634 (N_634,In_1931,In_2070);
xnor U635 (N_635,In_2829,In_220);
or U636 (N_636,In_2743,In_1387);
and U637 (N_637,In_706,In_1343);
and U638 (N_638,In_1006,In_1846);
xor U639 (N_639,In_2236,In_1205);
nor U640 (N_640,In_1048,In_2976);
nand U641 (N_641,In_669,In_2482);
or U642 (N_642,In_1318,In_1664);
and U643 (N_643,In_1439,In_2331);
and U644 (N_644,In_2549,In_1316);
nor U645 (N_645,In_1719,In_2177);
xnor U646 (N_646,In_2251,In_252);
nor U647 (N_647,In_2973,In_665);
xnor U648 (N_648,In_2707,In_2250);
or U649 (N_649,In_2387,In_1603);
or U650 (N_650,In_1907,In_57);
nand U651 (N_651,In_1957,In_1312);
and U652 (N_652,In_2013,In_972);
or U653 (N_653,In_626,In_2943);
nor U654 (N_654,In_2348,In_322);
or U655 (N_655,In_637,In_136);
nand U656 (N_656,In_1061,In_400);
nor U657 (N_657,In_752,In_455);
or U658 (N_658,In_2661,In_1436);
xor U659 (N_659,In_1631,In_1009);
and U660 (N_660,In_1123,In_1481);
nor U661 (N_661,In_2359,In_2540);
xor U662 (N_662,In_1083,In_661);
or U663 (N_663,In_2252,In_869);
xor U664 (N_664,In_521,In_361);
nor U665 (N_665,In_695,In_2788);
nor U666 (N_666,In_832,In_2208);
and U667 (N_667,In_2875,In_1308);
or U668 (N_668,In_442,In_606);
nor U669 (N_669,In_2998,In_1058);
nand U670 (N_670,In_1523,In_1147);
or U671 (N_671,In_2200,In_1259);
nor U672 (N_672,In_2430,In_2666);
nor U673 (N_673,In_55,In_1432);
nor U674 (N_674,In_2811,In_52);
xor U675 (N_675,In_659,In_1802);
xnor U676 (N_676,In_1363,In_764);
nor U677 (N_677,In_2824,In_2015);
nor U678 (N_678,In_270,In_1537);
and U679 (N_679,In_2448,In_1289);
nand U680 (N_680,In_160,In_2614);
and U681 (N_681,In_2016,In_574);
xor U682 (N_682,In_829,In_1169);
nor U683 (N_683,In_2152,In_1247);
nor U684 (N_684,In_371,In_2438);
or U685 (N_685,In_90,In_1300);
nand U686 (N_686,In_2306,In_1446);
xnor U687 (N_687,In_577,In_870);
or U688 (N_688,In_1827,In_102);
and U689 (N_689,In_1111,In_201);
nor U690 (N_690,In_204,In_2349);
xor U691 (N_691,In_338,In_2947);
xor U692 (N_692,In_942,In_1561);
and U693 (N_693,In_2676,In_1188);
nand U694 (N_694,In_2782,In_595);
nand U695 (N_695,In_2853,In_1098);
or U696 (N_696,In_1551,In_766);
and U697 (N_697,In_1255,In_298);
nand U698 (N_698,In_2380,In_1253);
or U699 (N_699,In_482,In_2316);
nand U700 (N_700,In_365,In_584);
or U701 (N_701,In_166,In_2303);
or U702 (N_702,In_1862,In_176);
nor U703 (N_703,In_1056,In_2771);
and U704 (N_704,In_2131,In_2820);
nand U705 (N_705,In_2507,In_763);
or U706 (N_706,In_2499,In_2974);
or U707 (N_707,In_2870,In_291);
xnor U708 (N_708,In_1326,In_1682);
xor U709 (N_709,In_1459,In_2373);
and U710 (N_710,In_586,In_1597);
or U711 (N_711,In_2523,In_2545);
nand U712 (N_712,In_1753,In_625);
nor U713 (N_713,In_981,In_4);
nand U714 (N_714,In_1991,In_1701);
xor U715 (N_715,In_2256,In_1124);
nor U716 (N_716,In_2925,In_2588);
xnor U717 (N_717,In_910,In_310);
xnor U718 (N_718,In_156,In_1621);
nor U719 (N_719,In_355,In_812);
and U720 (N_720,In_2722,In_303);
nor U721 (N_721,In_1734,In_2981);
nor U722 (N_722,In_314,In_2048);
nand U723 (N_723,In_1198,In_2806);
xor U724 (N_724,In_738,In_1448);
or U725 (N_725,In_1500,In_1457);
xor U726 (N_726,In_2846,In_453);
nor U727 (N_727,In_357,In_671);
and U728 (N_728,In_903,In_911);
xor U729 (N_729,In_2491,In_689);
xnor U730 (N_730,In_1126,In_877);
xor U731 (N_731,In_2904,In_2292);
and U732 (N_732,In_954,In_1529);
xor U733 (N_733,In_1816,In_24);
xnor U734 (N_734,In_1707,In_2623);
xor U735 (N_735,In_2436,In_1558);
or U736 (N_736,In_2277,In_287);
nand U737 (N_737,In_2567,In_1225);
nor U738 (N_738,In_2410,In_237);
xnor U739 (N_739,In_1746,In_2509);
or U740 (N_740,In_1398,In_666);
and U741 (N_741,In_2422,In_909);
nand U742 (N_742,In_755,In_2742);
xnor U743 (N_743,In_2886,In_975);
or U744 (N_744,In_1949,In_2755);
or U745 (N_745,In_2570,In_2443);
nand U746 (N_746,In_1405,In_1978);
and U747 (N_747,In_693,In_1520);
xor U748 (N_748,In_148,In_2510);
nor U749 (N_749,In_733,In_1375);
and U750 (N_750,In_366,In_851);
and U751 (N_751,In_1630,In_184);
nor U752 (N_752,In_1611,In_1024);
nand U753 (N_753,In_2601,In_1598);
xnor U754 (N_754,In_1518,In_1615);
nand U755 (N_755,In_34,In_1662);
nand U756 (N_756,In_1176,In_905);
nor U757 (N_757,In_410,In_1737);
and U758 (N_758,In_566,In_1044);
and U759 (N_759,In_1360,In_1271);
and U760 (N_760,In_849,In_1763);
and U761 (N_761,In_677,In_308);
nor U762 (N_762,In_846,In_786);
xor U763 (N_763,In_735,In_389);
and U764 (N_764,In_2547,In_916);
or U765 (N_765,In_1800,In_2924);
and U766 (N_766,In_1040,In_578);
nand U767 (N_767,In_2882,In_1187);
and U768 (N_768,In_2733,In_2826);
nor U769 (N_769,In_945,In_2485);
and U770 (N_770,In_479,In_839);
xnor U771 (N_771,In_2519,In_1595);
xnor U772 (N_772,In_194,In_2202);
nand U773 (N_773,In_864,In_387);
or U774 (N_774,In_924,In_1565);
nand U775 (N_775,In_598,In_1687);
xor U776 (N_776,In_390,In_1030);
or U777 (N_777,In_419,In_1892);
nand U778 (N_778,In_182,In_572);
or U779 (N_779,In_1004,In_1866);
and U780 (N_780,In_1645,In_1330);
xnor U781 (N_781,In_1462,In_2108);
nor U782 (N_782,In_770,In_740);
and U783 (N_783,In_437,In_428);
nand U784 (N_784,In_306,In_2265);
and U785 (N_785,In_1288,In_753);
nand U786 (N_786,In_425,In_2424);
and U787 (N_787,In_1409,In_714);
and U788 (N_788,In_367,In_2600);
or U789 (N_789,In_2641,In_682);
xnor U790 (N_790,In_1334,In_872);
and U791 (N_791,In_705,In_983);
or U792 (N_792,In_1908,In_1819);
nor U793 (N_793,In_2558,In_1848);
or U794 (N_794,In_1415,In_170);
nand U795 (N_795,In_878,In_1460);
xnor U796 (N_796,In_2102,In_997);
nor U797 (N_797,In_1998,In_196);
or U798 (N_798,In_1498,In_961);
or U799 (N_799,In_325,In_227);
nand U800 (N_800,In_1268,In_1172);
and U801 (N_801,In_420,In_2388);
nor U802 (N_802,In_1590,In_1329);
nand U803 (N_803,In_2219,In_783);
or U804 (N_804,In_737,In_741);
nor U805 (N_805,In_2612,In_332);
and U806 (N_806,In_1899,In_2363);
nor U807 (N_807,In_590,In_762);
and U808 (N_808,In_820,In_2927);
or U809 (N_809,In_2518,In_406);
xnor U810 (N_810,In_1177,In_344);
nand U811 (N_811,In_2060,In_26);
or U812 (N_812,In_2215,In_1101);
nand U813 (N_813,In_858,In_216);
xnor U814 (N_814,In_2286,In_534);
nor U815 (N_815,In_451,In_27);
and U816 (N_816,In_524,In_1497);
xnor U817 (N_817,In_1248,In_1178);
nor U818 (N_818,In_971,In_2091);
xor U819 (N_819,In_1238,In_2072);
or U820 (N_820,In_1469,In_2001);
or U821 (N_821,In_2966,In_1134);
and U822 (N_822,In_1190,In_2350);
nor U823 (N_823,In_36,In_81);
nor U824 (N_824,In_2858,In_522);
nor U825 (N_825,In_1219,In_1346);
and U826 (N_826,In_475,In_2311);
and U827 (N_827,In_2282,In_245);
or U828 (N_828,In_2245,In_2333);
xor U829 (N_829,In_2246,In_454);
nor U830 (N_830,In_436,In_2831);
xnor U831 (N_831,In_2205,In_2887);
nand U832 (N_832,In_2038,In_1479);
or U833 (N_833,In_1185,In_2888);
or U834 (N_834,In_369,In_2040);
nand U835 (N_835,In_2995,In_1803);
nor U836 (N_836,In_2395,In_1181);
or U837 (N_837,In_836,In_853);
and U838 (N_838,In_2085,In_1776);
and U839 (N_839,In_2987,In_748);
and U840 (N_840,In_1639,In_83);
xor U841 (N_841,In_1293,In_1287);
and U842 (N_842,In_2890,In_2474);
and U843 (N_843,In_1937,In_2583);
xnor U844 (N_844,In_431,In_2332);
xnor U845 (N_845,In_934,In_1493);
nor U846 (N_846,In_1571,In_513);
xnor U847 (N_847,In_71,In_1237);
xnor U848 (N_848,In_2754,In_776);
or U849 (N_849,In_938,In_2308);
nor U850 (N_850,In_1304,In_2279);
or U851 (N_851,In_2396,In_1036);
nand U852 (N_852,In_1921,In_1624);
xnor U853 (N_853,In_2901,In_2259);
xnor U854 (N_854,In_2866,In_1506);
or U855 (N_855,In_2624,In_2685);
nor U856 (N_856,In_324,In_1100);
or U857 (N_857,In_2402,In_2584);
xnor U858 (N_858,In_1585,In_1704);
xnor U859 (N_859,In_2224,In_1660);
or U860 (N_860,In_767,In_1053);
nand U861 (N_861,In_1226,In_263);
xnor U862 (N_862,In_1322,In_1396);
or U863 (N_863,In_1368,In_2903);
and U864 (N_864,In_229,In_164);
nor U865 (N_865,In_2032,In_1171);
and U866 (N_866,In_1204,In_2107);
and U867 (N_867,In_2957,In_234);
nand U868 (N_868,In_1383,In_793);
or U869 (N_869,In_785,In_2067);
xnor U870 (N_870,In_535,In_1884);
or U871 (N_871,In_1663,In_20);
or U872 (N_872,In_300,In_2141);
or U873 (N_873,In_988,In_2228);
nand U874 (N_874,In_2230,In_107);
nand U875 (N_875,In_2118,In_603);
or U876 (N_876,In_377,In_569);
xnor U877 (N_877,In_831,In_2278);
and U878 (N_878,In_2718,In_2248);
xor U879 (N_879,In_1328,In_1971);
and U880 (N_880,In_517,In_2658);
nor U881 (N_881,In_1079,In_953);
nand U882 (N_882,In_2899,In_757);
nand U883 (N_883,In_1382,In_2431);
nand U884 (N_884,In_2971,In_1733);
xor U885 (N_885,In_2566,In_2098);
xnor U886 (N_886,In_2254,In_1679);
and U887 (N_887,In_1883,In_1972);
xnor U888 (N_888,In_657,In_673);
xnor U889 (N_889,In_1760,In_2729);
nor U890 (N_890,In_967,In_2840);
xor U891 (N_891,In_127,In_2140);
xnor U892 (N_892,In_1609,In_2172);
or U893 (N_893,In_211,In_1620);
and U894 (N_894,In_1981,In_2682);
nand U895 (N_895,In_2419,In_485);
xor U896 (N_896,In_444,In_2706);
nor U897 (N_897,In_2929,In_545);
xnor U898 (N_898,In_2968,In_2497);
nand U899 (N_899,In_2442,In_489);
and U900 (N_900,In_2595,In_2229);
or U901 (N_901,In_684,In_907);
xor U902 (N_902,In_2512,In_41);
or U903 (N_903,In_384,In_2413);
and U904 (N_904,In_1696,In_2129);
and U905 (N_905,In_1946,In_147);
nand U906 (N_906,In_311,In_2695);
nand U907 (N_907,In_208,In_2390);
xnor U908 (N_908,In_2767,In_1070);
xor U909 (N_909,In_1049,In_2415);
nor U910 (N_910,In_716,In_315);
or U911 (N_911,In_1349,In_1774);
xnor U912 (N_912,In_1035,In_515);
and U913 (N_913,In_1987,In_2126);
xor U914 (N_914,In_2054,In_624);
and U915 (N_915,In_1885,In_462);
nor U916 (N_916,In_2552,In_2531);
nand U917 (N_917,In_458,In_1762);
or U918 (N_918,In_1882,In_2071);
nand U919 (N_919,In_2599,In_272);
nor U920 (N_920,In_1851,In_1974);
nor U921 (N_921,In_80,In_217);
or U922 (N_922,In_2938,In_373);
nor U923 (N_923,In_1037,In_1982);
xor U924 (N_924,In_2587,In_1869);
and U925 (N_925,In_183,In_1759);
nand U926 (N_926,In_2529,In_937);
nor U927 (N_927,In_2913,In_1559);
xor U928 (N_928,In_1606,In_1666);
xor U929 (N_929,In_151,In_947);
and U930 (N_930,In_2087,In_1472);
nor U931 (N_931,In_467,In_921);
nand U932 (N_932,In_2103,In_2317);
or U933 (N_933,In_2795,In_1572);
and U934 (N_934,In_2963,In_2667);
nand U935 (N_935,In_205,In_588);
nand U936 (N_936,In_638,In_1254);
or U937 (N_937,In_2656,In_2863);
or U938 (N_938,In_2994,In_866);
xor U939 (N_939,In_191,In_744);
or U940 (N_940,In_1654,In_1566);
and U941 (N_941,In_2628,In_203);
and U942 (N_942,In_1146,In_1108);
or U943 (N_943,In_1918,In_120);
nand U944 (N_944,In_1435,In_2854);
nor U945 (N_945,In_1916,In_456);
or U946 (N_946,In_2168,In_1570);
nand U947 (N_947,In_330,In_2234);
nor U948 (N_948,In_902,In_2675);
nand U949 (N_949,In_2242,In_1519);
nand U950 (N_950,In_914,In_2014);
nand U951 (N_951,In_1224,In_928);
or U952 (N_952,In_1075,In_833);
nand U953 (N_953,In_2371,In_1581);
nand U954 (N_954,In_135,In_647);
nand U955 (N_955,In_2320,In_1228);
or U956 (N_956,In_2083,In_1785);
and U957 (N_957,In_1923,In_2915);
or U958 (N_958,In_2157,In_2684);
nor U959 (N_959,In_163,In_2844);
nand U960 (N_960,In_1958,In_2783);
or U961 (N_961,In_1174,In_1860);
or U962 (N_962,In_2993,In_2673);
or U963 (N_963,In_1542,In_399);
xor U964 (N_964,In_1755,In_471);
nand U965 (N_965,In_1240,In_2381);
nor U966 (N_966,In_1842,In_1576);
nor U967 (N_967,In_1856,In_2832);
nor U968 (N_968,In_1017,In_2918);
and U969 (N_969,In_1905,In_675);
or U970 (N_970,In_2074,In_1586);
nor U971 (N_971,In_2521,In_2669);
nor U972 (N_972,In_2897,In_1054);
or U973 (N_973,In_2988,In_968);
nand U974 (N_974,In_1852,In_1728);
or U975 (N_975,In_5,In_895);
nor U976 (N_976,In_1494,In_2421);
xor U977 (N_977,In_2276,In_1661);
xor U978 (N_978,In_819,In_2194);
or U979 (N_979,In_15,In_464);
nand U980 (N_980,In_516,In_2999);
or U981 (N_981,In_804,In_602);
or U982 (N_982,In_627,In_1159);
xor U983 (N_983,In_117,In_1922);
xor U984 (N_984,In_346,In_2900);
and U985 (N_985,In_195,In_1814);
nand U986 (N_986,In_2857,In_2063);
and U987 (N_987,In_1927,In_2704);
or U988 (N_988,In_433,In_2937);
xor U989 (N_989,In_1830,In_238);
nand U990 (N_990,In_2537,In_1408);
nor U991 (N_991,In_530,In_2321);
xnor U992 (N_992,In_2207,In_2934);
xnor U993 (N_993,In_1627,In_711);
nand U994 (N_994,In_561,In_418);
xnor U995 (N_995,In_121,In_50);
or U996 (N_996,In_359,In_818);
xnor U997 (N_997,In_2094,In_2068);
xor U998 (N_998,In_1849,In_1944);
or U999 (N_999,In_676,In_1601);
or U1000 (N_1000,In_231,In_1766);
nand U1001 (N_1001,In_880,In_397);
and U1002 (N_1002,In_1445,In_2106);
nor U1003 (N_1003,In_2418,In_780);
nand U1004 (N_1004,In_2096,In_168);
or U1005 (N_1005,In_2374,In_782);
and U1006 (N_1006,In_1184,In_1568);
nor U1007 (N_1007,In_1186,In_2608);
and U1008 (N_1008,In_2243,In_2878);
and U1009 (N_1009,In_2217,In_1747);
nor U1010 (N_1010,In_2239,In_1751);
nor U1011 (N_1011,In_792,In_1370);
xnor U1012 (N_1012,In_1097,In_1222);
or U1013 (N_1013,In_2244,In_893);
nor U1014 (N_1014,In_2300,In_449);
xnor U1015 (N_1015,In_538,In_1137);
or U1016 (N_1016,In_61,In_1045);
xor U1017 (N_1017,In_2253,In_1019);
xor U1018 (N_1018,In_1195,In_2262);
or U1019 (N_1019,In_1076,In_1648);
or U1020 (N_1020,In_2362,In_312);
xnor U1021 (N_1021,In_473,In_417);
nand U1022 (N_1022,In_1,In_2403);
nor U1023 (N_1023,In_2627,In_1119);
nor U1024 (N_1024,In_2945,In_500);
nand U1025 (N_1025,In_2099,In_1826);
or U1026 (N_1026,In_1148,In_2954);
nor U1027 (N_1027,In_2138,In_2836);
xnor U1028 (N_1028,In_621,In_2582);
nor U1029 (N_1029,In_2427,In_2061);
and U1030 (N_1030,In_1967,In_1795);
xor U1031 (N_1031,In_368,In_69);
or U1032 (N_1032,In_2996,In_789);
or U1033 (N_1033,In_114,In_1689);
nand U1034 (N_1034,In_2690,In_889);
or U1035 (N_1035,In_459,In_1632);
nand U1036 (N_1036,In_1914,In_784);
nand U1037 (N_1037,In_173,In_1327);
nand U1038 (N_1038,In_765,In_279);
xnor U1039 (N_1039,In_1010,In_865);
or U1040 (N_1040,In_2780,In_1560);
nor U1041 (N_1041,In_2869,In_93);
nor U1042 (N_1042,In_2328,In_966);
and U1043 (N_1043,In_358,In_2517);
nand U1044 (N_1044,In_493,In_794);
or U1045 (N_1045,In_1608,In_2059);
nor U1046 (N_1046,In_2369,In_989);
nand U1047 (N_1047,In_2688,In_1665);
xor U1048 (N_1048,In_1306,In_1295);
xor U1049 (N_1049,In_607,In_1792);
or U1050 (N_1050,In_573,In_1843);
or U1051 (N_1051,In_1099,In_1158);
xor U1052 (N_1052,In_1362,In_646);
or U1053 (N_1053,In_1787,In_2370);
nor U1054 (N_1054,In_1476,In_1475);
xor U1055 (N_1055,In_559,In_1069);
and U1056 (N_1056,In_1678,In_1557);
nor U1057 (N_1057,In_188,In_175);
nand U1058 (N_1058,In_1934,In_2023);
or U1059 (N_1059,In_2808,In_796);
or U1060 (N_1060,In_525,In_1473);
nand U1061 (N_1061,In_1538,In_2290);
nor U1062 (N_1062,In_1853,In_2445);
nand U1063 (N_1063,In_549,In_642);
nand U1064 (N_1064,In_1727,In_483);
nor U1065 (N_1065,In_1700,In_328);
nor U1066 (N_1066,In_2319,In_1131);
nor U1067 (N_1067,In_2082,In_1877);
or U1068 (N_1068,In_2472,In_1919);
or U1069 (N_1069,In_568,In_2109);
xor U1070 (N_1070,In_2848,In_1709);
xor U1071 (N_1071,In_2018,In_2398);
nand U1072 (N_1072,In_2383,In_1933);
nand U1073 (N_1073,In_2750,In_1990);
and U1074 (N_1074,In_1251,In_1492);
nand U1075 (N_1075,In_1514,In_469);
or U1076 (N_1076,In_1951,In_1065);
or U1077 (N_1077,In_656,In_2809);
or U1078 (N_1078,In_1637,In_747);
xor U1079 (N_1079,In_23,In_991);
xor U1080 (N_1080,In_2167,In_1162);
or U1081 (N_1081,In_68,In_396);
or U1082 (N_1082,In_2732,In_1768);
xor U1083 (N_1083,In_1341,In_1588);
nor U1084 (N_1084,In_133,In_2122);
or U1085 (N_1085,In_655,In_2136);
or U1086 (N_1086,In_2414,In_2124);
nand U1087 (N_1087,In_1865,In_2447);
xor U1088 (N_1088,In_1050,In_2735);
or U1089 (N_1089,In_712,In_1128);
or U1090 (N_1090,In_385,In_1720);
nand U1091 (N_1091,In_1730,In_1132);
nand U1092 (N_1092,In_583,In_2842);
or U1093 (N_1093,In_2760,In_146);
or U1094 (N_1094,In_2816,In_1414);
or U1095 (N_1095,In_1619,In_6);
nand U1096 (N_1096,In_2801,In_822);
nor U1097 (N_1097,In_725,In_958);
and U1098 (N_1098,In_1835,In_2173);
nor U1099 (N_1099,In_264,In_1732);
nand U1100 (N_1100,In_2329,In_2665);
or U1101 (N_1101,In_1042,In_2835);
and U1102 (N_1102,In_256,In_791);
nor U1103 (N_1103,In_67,In_292);
or U1104 (N_1104,In_1977,In_724);
nand U1105 (N_1105,In_651,In_933);
nand U1106 (N_1106,In_174,In_1484);
and U1107 (N_1107,In_1090,In_1717);
nor U1108 (N_1108,In_492,In_2005);
nand U1109 (N_1109,In_1706,In_395);
nor U1110 (N_1110,In_1699,In_871);
xnor U1111 (N_1111,In_1984,In_2225);
nand U1112 (N_1112,In_1323,In_1622);
nand U1113 (N_1113,In_1000,In_472);
or U1114 (N_1114,In_2065,In_2358);
nor U1115 (N_1115,In_1573,In_1963);
nor U1116 (N_1116,In_92,In_63);
nand U1117 (N_1117,In_1258,In_207);
xor U1118 (N_1118,In_2532,In_225);
and U1119 (N_1119,In_106,In_1556);
nor U1120 (N_1120,In_1291,In_2909);
and U1121 (N_1121,In_1988,In_1456);
nand U1122 (N_1122,In_2111,In_1116);
nand U1123 (N_1123,In_2727,In_1867);
xor U1124 (N_1124,In_1153,In_2837);
xor U1125 (N_1125,In_380,In_1420);
nor U1126 (N_1126,In_2397,In_842);
nor U1127 (N_1127,In_710,In_1794);
and U1128 (N_1128,In_828,In_1809);
xnor U1129 (N_1129,In_30,In_8);
xor U1130 (N_1130,In_2557,In_60);
xnor U1131 (N_1131,In_1427,In_1216);
or U1132 (N_1132,In_1509,In_99);
xnor U1133 (N_1133,In_1942,In_53);
and U1134 (N_1134,In_2770,In_1854);
or U1135 (N_1135,In_2907,In_2088);
and U1136 (N_1136,In_1426,In_579);
xor U1137 (N_1137,In_2154,In_2959);
or U1138 (N_1138,In_746,In_1451);
nand U1139 (N_1139,In_1773,In_2991);
xor U1140 (N_1140,In_374,In_70);
and U1141 (N_1141,In_414,In_1838);
xnor U1142 (N_1142,In_1135,In_1647);
or U1143 (N_1143,In_653,In_2766);
and U1144 (N_1144,In_1466,In_1273);
nor U1145 (N_1145,In_723,In_301);
nor U1146 (N_1146,In_1369,In_66);
nor U1147 (N_1147,In_2828,In_13);
nand U1148 (N_1148,In_235,In_445);
nand U1149 (N_1149,In_2466,In_1881);
xor U1150 (N_1150,In_2794,In_2581);
xnor U1151 (N_1151,In_2699,In_2914);
nand U1152 (N_1152,In_2922,In_2539);
or U1153 (N_1153,In_1670,In_141);
nand U1154 (N_1154,In_2128,In_2134);
nand U1155 (N_1155,In_2483,In_2119);
and U1156 (N_1156,In_1490,In_2307);
and U1157 (N_1157,In_39,In_2322);
nand U1158 (N_1158,In_239,In_2935);
and U1159 (N_1159,In_19,In_1941);
nand U1160 (N_1160,In_699,In_2197);
nor U1161 (N_1161,In_267,In_2984);
nand U1162 (N_1162,In_1026,In_1130);
nor U1163 (N_1163,In_1113,In_1625);
nand U1164 (N_1164,In_837,In_1778);
nand U1165 (N_1165,In_1199,In_1335);
nor U1166 (N_1166,In_2041,In_2575);
xor U1167 (N_1167,In_2471,In_2642);
xor U1168 (N_1168,In_2804,In_808);
and U1169 (N_1169,In_250,In_1047);
nor U1170 (N_1170,In_881,In_452);
nor U1171 (N_1171,In_2553,In_388);
and U1172 (N_1172,In_857,In_2160);
nor U1173 (N_1173,In_1440,In_378);
and U1174 (N_1174,In_557,In_2104);
nor U1175 (N_1175,In_498,In_2156);
xor U1176 (N_1176,In_1545,In_2342);
nor U1177 (N_1177,In_2942,In_1365);
nand U1178 (N_1178,In_190,In_2406);
and U1179 (N_1179,In_25,In_2494);
and U1180 (N_1180,In_2294,In_1197);
nor U1181 (N_1181,In_2779,In_1811);
and U1182 (N_1182,In_277,In_2789);
or U1183 (N_1183,In_1109,In_1213);
xnor U1184 (N_1184,In_2668,In_1022);
nand U1185 (N_1185,In_1935,In_1930);
nor U1186 (N_1186,In_2541,In_2266);
and U1187 (N_1187,In_977,In_2283);
nand U1188 (N_1188,In_554,In_1232);
or U1189 (N_1189,In_421,In_1693);
nand U1190 (N_1190,In_505,In_1450);
nand U1191 (N_1191,In_392,In_749);
nand U1192 (N_1192,In_1878,In_551);
nand U1193 (N_1193,In_439,In_1063);
and U1194 (N_1194,In_1567,In_1992);
nand U1195 (N_1195,In_2562,In_520);
nand U1196 (N_1196,In_503,In_2046);
nor U1197 (N_1197,In_2486,In_2484);
xor U1198 (N_1198,In_2375,In_221);
and U1199 (N_1199,In_2785,In_2045);
or U1200 (N_1200,In_694,In_567);
and U1201 (N_1201,In_1767,In_2752);
and U1202 (N_1202,In_1164,In_1496);
and U1203 (N_1203,In_2417,In_2723);
or U1204 (N_1204,In_1837,In_309);
and U1205 (N_1205,In_1129,In_1183);
and U1206 (N_1206,In_1023,In_1895);
or U1207 (N_1207,In_1483,In_1338);
and U1208 (N_1208,In_1880,In_1215);
xor U1209 (N_1209,In_2161,In_1357);
nand U1210 (N_1210,In_2528,In_2565);
xor U1211 (N_1211,In_2223,In_984);
nor U1212 (N_1212,In_1898,In_438);
and U1213 (N_1213,In_1653,In_885);
and U1214 (N_1214,In_2377,In_2526);
and U1215 (N_1215,In_1384,In_597);
xor U1216 (N_1216,In_2301,In_76);
nor U1217 (N_1217,In_636,In_1501);
nand U1218 (N_1218,In_1915,In_2231);
and U1219 (N_1219,In_2551,In_1610);
nand U1220 (N_1220,In_973,In_2724);
or U1221 (N_1221,In_904,In_1876);
or U1222 (N_1222,In_1902,In_504);
nand U1223 (N_1223,In_474,In_2969);
nand U1224 (N_1224,In_692,In_756);
or U1225 (N_1225,In_2180,In_2050);
nor U1226 (N_1226,In_218,In_1084);
xnor U1227 (N_1227,In_144,In_1296);
nor U1228 (N_1228,In_635,In_841);
nor U1229 (N_1229,In_259,In_2391);
nor U1230 (N_1230,In_1280,In_2769);
and U1231 (N_1231,In_2401,In_2459);
xnor U1232 (N_1232,In_719,In_2164);
or U1233 (N_1233,In_2386,In_1936);
nor U1234 (N_1234,In_297,In_2132);
or U1235 (N_1235,In_271,In_2501);
and U1236 (N_1236,In_2343,In_1041);
nor U1237 (N_1237,In_2220,In_2564);
nor U1238 (N_1238,In_581,In_1968);
and U1239 (N_1239,In_2035,In_2340);
or U1240 (N_1240,In_37,In_696);
or U1241 (N_1241,In_290,In_2772);
and U1242 (N_1242,In_2033,In_1239);
and U1243 (N_1243,In_1441,In_563);
or U1244 (N_1244,In_2309,In_1580);
nor U1245 (N_1245,In_2597,In_223);
nor U1246 (N_1246,In_209,In_2821);
nand U1247 (N_1247,In_2105,In_405);
and U1248 (N_1248,In_1801,In_806);
and U1249 (N_1249,In_178,In_2741);
nand U1250 (N_1250,In_2365,In_788);
xor U1251 (N_1251,In_179,In_2337);
and U1252 (N_1252,In_1817,In_587);
and U1253 (N_1253,In_2216,In_2884);
nand U1254 (N_1254,In_925,In_1081);
nor U1255 (N_1255,In_546,In_2149);
nand U1256 (N_1256,In_323,In_1616);
nand U1257 (N_1257,In_364,In_999);
nor U1258 (N_1258,In_2027,In_2573);
and U1259 (N_1259,In_821,In_2354);
nor U1260 (N_1260,In_1748,In_2487);
xor U1261 (N_1261,In_45,In_1813);
and U1262 (N_1262,In_1605,In_2985);
nor U1263 (N_1263,In_2297,In_629);
xor U1264 (N_1264,In_1133,In_1749);
nor U1265 (N_1265,In_652,In_2905);
and U1266 (N_1266,In_2681,In_1845);
or U1267 (N_1267,In_843,In_329);
xor U1268 (N_1268,In_2579,In_2631);
nor U1269 (N_1269,In_1161,In_327);
xor U1270 (N_1270,In_2881,In_860);
or U1271 (N_1271,In_1698,In_861);
or U1272 (N_1272,In_118,In_108);
nand U1273 (N_1273,In_2449,In_690);
or U1274 (N_1274,In_2385,In_2150);
and U1275 (N_1275,In_145,In_1102);
nand U1276 (N_1276,In_2638,In_1297);
nand U1277 (N_1277,In_159,In_1824);
and U1278 (N_1278,In_450,In_1543);
nand U1279 (N_1279,In_1872,In_901);
or U1280 (N_1280,In_1993,In_2877);
xor U1281 (N_1281,In_46,In_2453);
nor U1282 (N_1282,In_2639,In_1917);
xnor U1283 (N_1283,In_532,In_2392);
and U1284 (N_1284,In_2233,In_2);
xnor U1285 (N_1285,In_867,In_713);
nor U1286 (N_1286,In_2865,In_1953);
or U1287 (N_1287,In_2819,In_1791);
and U1288 (N_1288,In_683,In_408);
and U1289 (N_1289,In_1840,In_2165);
and U1290 (N_1290,In_612,In_940);
and U1291 (N_1291,In_1020,In_644);
and U1292 (N_1292,In_1077,In_582);
nand U1293 (N_1293,In_1893,In_360);
nor U1294 (N_1294,In_1392,In_2683);
nor U1295 (N_1295,In_815,In_1294);
nand U1296 (N_1296,In_342,In_1263);
nor U1297 (N_1297,In_1850,In_772);
and U1298 (N_1298,In_1103,In_1859);
nor U1299 (N_1299,In_1741,In_2444);
or U1300 (N_1300,In_691,In_1901);
and U1301 (N_1301,In_2896,In_407);
or U1302 (N_1302,In_2287,In_1276);
or U1303 (N_1303,In_1394,In_320);
nor U1304 (N_1304,In_969,In_970);
and U1305 (N_1305,In_1652,In_701);
or U1306 (N_1306,In_2339,In_1095);
or U1307 (N_1307,In_2650,In_995);
xor U1308 (N_1308,In_337,In_645);
or U1309 (N_1309,In_243,In_533);
and U1310 (N_1310,In_2653,In_761);
nand U1311 (N_1311,In_2847,In_685);
nor U1312 (N_1312,In_268,In_1080);
nand U1313 (N_1313,In_2143,In_1072);
or U1314 (N_1314,In_1489,In_2739);
and U1315 (N_1315,In_2026,In_1423);
and U1316 (N_1316,In_874,In_2798);
xnor U1317 (N_1317,In_2502,In_2889);
nor U1318 (N_1318,In_731,In_2100);
or U1319 (N_1319,In_1742,In_1093);
nand U1320 (N_1320,In_1574,In_2464);
nor U1321 (N_1321,In_1628,In_1358);
and U1322 (N_1322,In_2849,In_2081);
and U1323 (N_1323,In_1317,In_403);
nand U1324 (N_1324,In_2434,In_74);
and U1325 (N_1325,In_2121,In_2353);
and U1326 (N_1326,In_1425,In_1399);
and U1327 (N_1327,In_1532,In_2455);
nand U1328 (N_1328,In_333,In_1906);
and U1329 (N_1329,In_2621,In_2872);
nor U1330 (N_1330,In_913,In_1725);
nand U1331 (N_1331,In_345,In_2372);
xor U1332 (N_1332,In_1144,In_963);
nand U1333 (N_1333,In_132,In_2209);
or U1334 (N_1334,In_2797,In_2002);
xnor U1335 (N_1335,In_2073,In_1118);
nand U1336 (N_1336,In_2796,In_774);
nand U1337 (N_1337,In_2738,In_1873);
or U1338 (N_1338,In_1555,In_994);
and U1339 (N_1339,In_742,In_750);
nand U1340 (N_1340,In_2275,In_805);
nand U1341 (N_1341,In_601,In_1142);
xnor U1342 (N_1342,In_2084,In_518);
nor U1343 (N_1343,In_1372,In_1324);
and U1344 (N_1344,In_844,In_2778);
or U1345 (N_1345,In_2360,In_1347);
or U1346 (N_1346,In_1910,In_2910);
nand U1347 (N_1347,In_187,In_570);
nand U1348 (N_1348,In_1227,In_2940);
nor U1349 (N_1349,In_1421,In_1804);
xnor U1350 (N_1350,In_2006,In_2800);
xnor U1351 (N_1351,In_266,In_281);
or U1352 (N_1352,In_1815,In_2880);
nand U1353 (N_1353,In_2611,In_855);
or U1354 (N_1354,In_1841,In_982);
nor U1355 (N_1355,In_1283,In_17);
and U1356 (N_1356,In_2463,In_1705);
or U1357 (N_1357,In_2843,In_608);
and U1358 (N_1358,In_1788,In_2330);
and U1359 (N_1359,In_1373,In_1810);
nor U1360 (N_1360,In_1911,In_589);
nand U1361 (N_1361,In_1003,In_161);
nand U1362 (N_1362,In_2679,In_440);
xor U1363 (N_1363,In_2476,In_879);
nand U1364 (N_1364,In_1695,In_2906);
or U1365 (N_1365,In_1269,In_331);
nand U1366 (N_1366,In_552,In_616);
nand U1367 (N_1367,In_2746,In_1032);
nor U1368 (N_1368,In_894,In_2663);
xnor U1369 (N_1369,In_43,In_884);
xnor U1370 (N_1370,In_514,In_2505);
or U1371 (N_1371,In_1094,In_87);
nand U1372 (N_1372,In_1903,In_816);
nor U1373 (N_1373,In_2151,In_1940);
xor U1374 (N_1374,In_2264,In_1959);
nor U1375 (N_1375,In_105,In_370);
or U1376 (N_1376,In_1950,In_2258);
nor U1377 (N_1377,In_1721,In_1117);
nand U1378 (N_1378,In_2481,In_2615);
or U1379 (N_1379,In_185,In_2047);
xnor U1380 (N_1380,In_1939,In_927);
and U1381 (N_1381,In_2572,In_1167);
and U1382 (N_1382,In_22,In_284);
xor U1383 (N_1383,In_810,In_2030);
or U1384 (N_1384,In_2859,In_1465);
nor U1385 (N_1385,In_94,In_2411);
and U1386 (N_1386,In_1175,In_1064);
xor U1387 (N_1387,In_978,In_510);
xor U1388 (N_1388,In_1544,In_1502);
or U1389 (N_1389,In_2717,In_1712);
nor U1390 (N_1390,In_1668,In_2212);
nand U1391 (N_1391,In_2740,In_100);
or U1392 (N_1392,In_915,In_461);
and U1393 (N_1393,In_1156,In_210);
or U1394 (N_1394,In_1191,In_2757);
xor U1395 (N_1395,In_468,In_2646);
and U1396 (N_1396,In_2802,In_1141);
and U1397 (N_1397,In_1535,In_2951);
nand U1398 (N_1398,In_394,In_634);
xor U1399 (N_1399,In_2432,In_2975);
xor U1400 (N_1400,In_1833,In_416);
xor U1401 (N_1401,In_2166,In_490);
nor U1402 (N_1402,In_278,In_2078);
nand U1403 (N_1403,In_2274,In_2980);
nand U1404 (N_1404,In_1507,In_906);
nor U1405 (N_1405,In_1858,In_1986);
nor U1406 (N_1406,In_1736,In_75);
xor U1407 (N_1407,In_2064,In_1221);
xor U1408 (N_1408,In_1447,In_2677);
nor U1409 (N_1409,In_411,In_891);
xnor U1410 (N_1410,In_1402,In_2873);
xnor U1411 (N_1411,In_1356,In_1569);
and U1412 (N_1412,In_1014,In_1201);
xor U1413 (N_1413,In_162,In_2127);
nor U1414 (N_1414,In_779,In_2090);
xor U1415 (N_1415,In_2404,In_542);
xnor U1416 (N_1416,In_2186,In_2271);
xor U1417 (N_1417,In_797,In_987);
and U1418 (N_1418,In_1799,In_1783);
xnor U1419 (N_1419,In_1182,In_2855);
nor U1420 (N_1420,In_82,In_717);
xor U1421 (N_1421,In_1350,In_1257);
nor U1422 (N_1422,In_876,In_1797);
nand U1423 (N_1423,In_2181,In_1057);
xnor U1424 (N_1424,In_807,In_2525);
nand U1425 (N_1425,In_137,In_888);
nand U1426 (N_1426,In_1033,In_2636);
or U1427 (N_1427,In_734,In_1107);
or U1428 (N_1428,In_2709,In_2198);
or U1429 (N_1429,In_729,In_1487);
nor U1430 (N_1430,In_900,In_1212);
and U1431 (N_1431,In_2288,In_2749);
or U1432 (N_1432,In_2153,In_648);
or U1433 (N_1433,In_850,In_2923);
nor U1434 (N_1434,In_383,In_2822);
xor U1435 (N_1435,In_1828,In_1404);
nand U1436 (N_1436,In_1407,In_1046);
nand U1437 (N_1437,In_771,In_109);
nand U1438 (N_1438,In_721,In_2983);
nor U1439 (N_1439,In_799,In_908);
xor U1440 (N_1440,In_341,In_1468);
and U1441 (N_1441,In_2429,In_1790);
nand U1442 (N_1442,In_1684,In_96);
xor U1443 (N_1443,In_31,In_2860);
nor U1444 (N_1444,In_2479,In_1333);
nand U1445 (N_1445,In_2240,In_2191);
nor U1446 (N_1446,In_1001,In_336);
and U1447 (N_1447,In_299,In_2441);
and U1448 (N_1448,In_1397,In_2162);
nor U1449 (N_1449,In_698,In_2260);
and U1450 (N_1450,In_1385,In_912);
xor U1451 (N_1451,In_2930,In_1710);
nor U1452 (N_1452,In_1539,In_674);
xnor U1453 (N_1453,In_429,In_1602);
xnor U1454 (N_1454,In_2892,In_2950);
nor U1455 (N_1455,In_2272,In_1694);
or U1456 (N_1456,In_465,In_1855);
xnor U1457 (N_1457,In_447,In_1467);
and U1458 (N_1458,In_1669,In_2660);
nand U1459 (N_1459,In_890,In_1264);
or U1460 (N_1460,In_123,In_460);
xnor U1461 (N_1461,In_2659,In_814);
and U1462 (N_1462,In_1638,In_33);
nor U1463 (N_1463,In_296,In_409);
or U1464 (N_1464,In_1086,In_2932);
nor U1465 (N_1465,In_1962,In_1612);
or U1466 (N_1466,In_2446,In_1311);
and U1467 (N_1467,In_509,In_293);
nor U1468 (N_1468,In_2190,In_2004);
and U1469 (N_1469,In_2495,In_1488);
or U1470 (N_1470,In_980,In_2457);
nor U1471 (N_1471,In_2187,In_295);
xnor U1472 (N_1472,In_1552,In_2744);
nor U1473 (N_1473,In_2756,In_847);
nor U1474 (N_1474,In_2489,In_241);
and U1475 (N_1475,In_1386,In_1401);
xor U1476 (N_1476,In_347,In_134);
nand U1477 (N_1477,In_1582,In_1861);
nand U1478 (N_1478,In_2508,In_2130);
and U1479 (N_1479,In_283,In_1015);
and U1480 (N_1480,In_260,In_759);
xor U1481 (N_1481,In_1486,In_919);
nor U1482 (N_1482,In_2456,In_258);
and U1483 (N_1483,In_1643,In_356);
xnor U1484 (N_1484,In_957,In_248);
nor U1485 (N_1485,In_1979,In_2480);
nor U1486 (N_1486,In_1031,In_228);
and U1487 (N_1487,In_1871,In_112);
nor U1488 (N_1488,In_633,In_2883);
or U1489 (N_1489,In_1089,In_1139);
nand U1490 (N_1490,In_1808,In_466);
nand U1491 (N_1491,In_1744,In_2698);
and U1492 (N_1492,In_2298,In_2232);
and U1493 (N_1493,In_614,In_1180);
xor U1494 (N_1494,In_2469,In_2833);
nand U1495 (N_1495,In_848,In_2902);
xnor U1496 (N_1496,In_2961,In_917);
and U1497 (N_1497,In_402,In_1592);
xor U1498 (N_1498,In_2977,In_285);
or U1499 (N_1499,In_1206,In_527);
or U1500 (N_1500,In_2072,In_2628);
nor U1501 (N_1501,In_1417,In_142);
nand U1502 (N_1502,In_1998,In_2834);
nor U1503 (N_1503,In_2640,In_644);
nand U1504 (N_1504,In_466,In_1207);
xnor U1505 (N_1505,In_1180,In_863);
or U1506 (N_1506,In_1250,In_1799);
nor U1507 (N_1507,In_554,In_691);
or U1508 (N_1508,In_437,In_1592);
xor U1509 (N_1509,In_2297,In_778);
xor U1510 (N_1510,In_2322,In_1811);
or U1511 (N_1511,In_2005,In_1513);
xnor U1512 (N_1512,In_2682,In_204);
xnor U1513 (N_1513,In_2569,In_1220);
xnor U1514 (N_1514,In_1696,In_114);
nand U1515 (N_1515,In_2328,In_904);
xor U1516 (N_1516,In_1419,In_1210);
nand U1517 (N_1517,In_1027,In_844);
nor U1518 (N_1518,In_1962,In_2428);
nand U1519 (N_1519,In_2313,In_1632);
nor U1520 (N_1520,In_985,In_1332);
or U1521 (N_1521,In_2849,In_726);
nor U1522 (N_1522,In_857,In_1220);
or U1523 (N_1523,In_94,In_1109);
xor U1524 (N_1524,In_1056,In_2876);
nor U1525 (N_1525,In_799,In_1569);
xor U1526 (N_1526,In_2185,In_2093);
and U1527 (N_1527,In_395,In_2424);
nor U1528 (N_1528,In_2268,In_1545);
nand U1529 (N_1529,In_1334,In_1309);
xor U1530 (N_1530,In_1201,In_727);
nor U1531 (N_1531,In_1435,In_672);
and U1532 (N_1532,In_2229,In_2374);
xnor U1533 (N_1533,In_2370,In_1844);
and U1534 (N_1534,In_2040,In_1533);
nor U1535 (N_1535,In_2027,In_512);
and U1536 (N_1536,In_2801,In_2939);
nand U1537 (N_1537,In_319,In_950);
or U1538 (N_1538,In_1120,In_868);
xor U1539 (N_1539,In_2989,In_2791);
nand U1540 (N_1540,In_2108,In_556);
or U1541 (N_1541,In_278,In_1293);
nand U1542 (N_1542,In_833,In_905);
or U1543 (N_1543,In_2724,In_2933);
nand U1544 (N_1544,In_459,In_462);
xor U1545 (N_1545,In_1285,In_1062);
nor U1546 (N_1546,In_2170,In_2460);
nor U1547 (N_1547,In_1908,In_1138);
nor U1548 (N_1548,In_2951,In_1422);
nor U1549 (N_1549,In_2067,In_2120);
nand U1550 (N_1550,In_2649,In_1263);
xor U1551 (N_1551,In_1612,In_442);
nand U1552 (N_1552,In_2343,In_1616);
nor U1553 (N_1553,In_1238,In_2295);
and U1554 (N_1554,In_2919,In_283);
and U1555 (N_1555,In_1196,In_1633);
and U1556 (N_1556,In_997,In_1681);
nor U1557 (N_1557,In_1789,In_278);
or U1558 (N_1558,In_2903,In_2457);
and U1559 (N_1559,In_1423,In_769);
nand U1560 (N_1560,In_112,In_702);
and U1561 (N_1561,In_1293,In_88);
nor U1562 (N_1562,In_664,In_103);
nor U1563 (N_1563,In_2306,In_744);
or U1564 (N_1564,In_989,In_1743);
nand U1565 (N_1565,In_2840,In_1031);
nor U1566 (N_1566,In_919,In_918);
nand U1567 (N_1567,In_2656,In_2763);
xor U1568 (N_1568,In_2063,In_1004);
or U1569 (N_1569,In_34,In_162);
nand U1570 (N_1570,In_488,In_1791);
nand U1571 (N_1571,In_2613,In_1390);
nor U1572 (N_1572,In_2192,In_1086);
or U1573 (N_1573,In_833,In_2715);
or U1574 (N_1574,In_8,In_2574);
or U1575 (N_1575,In_1793,In_921);
and U1576 (N_1576,In_1842,In_556);
and U1577 (N_1577,In_2412,In_2506);
or U1578 (N_1578,In_381,In_1842);
xor U1579 (N_1579,In_2041,In_1681);
xor U1580 (N_1580,In_1657,In_1159);
nor U1581 (N_1581,In_2301,In_1270);
or U1582 (N_1582,In_800,In_2137);
nand U1583 (N_1583,In_191,In_148);
nor U1584 (N_1584,In_602,In_586);
or U1585 (N_1585,In_810,In_738);
nand U1586 (N_1586,In_1543,In_587);
and U1587 (N_1587,In_571,In_2229);
and U1588 (N_1588,In_587,In_2312);
xnor U1589 (N_1589,In_2040,In_1717);
nor U1590 (N_1590,In_176,In_2439);
and U1591 (N_1591,In_2695,In_2725);
xnor U1592 (N_1592,In_934,In_426);
nand U1593 (N_1593,In_2217,In_123);
xnor U1594 (N_1594,In_79,In_570);
or U1595 (N_1595,In_923,In_1969);
xnor U1596 (N_1596,In_533,In_1186);
nand U1597 (N_1597,In_2733,In_514);
or U1598 (N_1598,In_1752,In_1001);
xnor U1599 (N_1599,In_671,In_2945);
nand U1600 (N_1600,In_1900,In_1367);
nand U1601 (N_1601,In_1178,In_648);
or U1602 (N_1602,In_1814,In_1020);
nor U1603 (N_1603,In_853,In_880);
or U1604 (N_1604,In_2239,In_1006);
xnor U1605 (N_1605,In_91,In_2374);
or U1606 (N_1606,In_1154,In_473);
nor U1607 (N_1607,In_1397,In_1760);
and U1608 (N_1608,In_2203,In_1190);
nor U1609 (N_1609,In_1485,In_1170);
nor U1610 (N_1610,In_2021,In_2330);
nor U1611 (N_1611,In_2048,In_2871);
and U1612 (N_1612,In_2327,In_2838);
xnor U1613 (N_1613,In_153,In_2383);
xnor U1614 (N_1614,In_2284,In_2461);
or U1615 (N_1615,In_732,In_505);
or U1616 (N_1616,In_2281,In_2084);
nor U1617 (N_1617,In_395,In_1777);
xnor U1618 (N_1618,In_1092,In_2745);
nor U1619 (N_1619,In_486,In_568);
nor U1620 (N_1620,In_2505,In_2506);
and U1621 (N_1621,In_2235,In_115);
xnor U1622 (N_1622,In_2891,In_1222);
and U1623 (N_1623,In_2130,In_507);
nand U1624 (N_1624,In_2944,In_743);
nand U1625 (N_1625,In_835,In_225);
and U1626 (N_1626,In_1911,In_171);
or U1627 (N_1627,In_2378,In_1533);
nor U1628 (N_1628,In_2388,In_1182);
nor U1629 (N_1629,In_2872,In_654);
nor U1630 (N_1630,In_2766,In_2036);
xnor U1631 (N_1631,In_720,In_314);
or U1632 (N_1632,In_560,In_170);
or U1633 (N_1633,In_2750,In_2829);
nand U1634 (N_1634,In_544,In_2664);
nand U1635 (N_1635,In_2633,In_1943);
nor U1636 (N_1636,In_649,In_1564);
nor U1637 (N_1637,In_2000,In_2944);
xnor U1638 (N_1638,In_1113,In_1385);
nor U1639 (N_1639,In_645,In_791);
or U1640 (N_1640,In_2236,In_1586);
and U1641 (N_1641,In_1709,In_2161);
nor U1642 (N_1642,In_848,In_923);
and U1643 (N_1643,In_2821,In_840);
or U1644 (N_1644,In_856,In_2442);
nand U1645 (N_1645,In_160,In_1184);
nand U1646 (N_1646,In_2741,In_1597);
or U1647 (N_1647,In_2609,In_1600);
xor U1648 (N_1648,In_105,In_65);
and U1649 (N_1649,In_1356,In_299);
and U1650 (N_1650,In_92,In_302);
nand U1651 (N_1651,In_2202,In_627);
or U1652 (N_1652,In_2837,In_2823);
and U1653 (N_1653,In_74,In_196);
or U1654 (N_1654,In_481,In_2745);
and U1655 (N_1655,In_1874,In_2734);
and U1656 (N_1656,In_2427,In_2939);
nand U1657 (N_1657,In_2546,In_1376);
and U1658 (N_1658,In_873,In_2425);
xor U1659 (N_1659,In_845,In_525);
and U1660 (N_1660,In_299,In_848);
nor U1661 (N_1661,In_731,In_353);
nor U1662 (N_1662,In_1322,In_800);
nor U1663 (N_1663,In_963,In_2780);
xnor U1664 (N_1664,In_1655,In_1315);
nand U1665 (N_1665,In_1764,In_428);
nor U1666 (N_1666,In_2567,In_2040);
or U1667 (N_1667,In_1043,In_455);
and U1668 (N_1668,In_40,In_1613);
nor U1669 (N_1669,In_345,In_1674);
nor U1670 (N_1670,In_2309,In_1665);
xor U1671 (N_1671,In_1836,In_2638);
nor U1672 (N_1672,In_1830,In_2909);
or U1673 (N_1673,In_2017,In_2657);
and U1674 (N_1674,In_635,In_2184);
nand U1675 (N_1675,In_974,In_1742);
and U1676 (N_1676,In_485,In_2848);
and U1677 (N_1677,In_728,In_2098);
xnor U1678 (N_1678,In_479,In_2819);
or U1679 (N_1679,In_2527,In_850);
nand U1680 (N_1680,In_458,In_2609);
xor U1681 (N_1681,In_1853,In_764);
nor U1682 (N_1682,In_1082,In_328);
nand U1683 (N_1683,In_549,In_651);
nor U1684 (N_1684,In_53,In_773);
nor U1685 (N_1685,In_1292,In_310);
and U1686 (N_1686,In_230,In_1676);
nand U1687 (N_1687,In_1807,In_115);
nand U1688 (N_1688,In_796,In_2696);
xor U1689 (N_1689,In_2924,In_1363);
and U1690 (N_1690,In_2752,In_2805);
and U1691 (N_1691,In_2906,In_72);
and U1692 (N_1692,In_2256,In_2817);
nand U1693 (N_1693,In_2851,In_2702);
and U1694 (N_1694,In_2250,In_1721);
xor U1695 (N_1695,In_1629,In_1254);
and U1696 (N_1696,In_2013,In_1277);
nor U1697 (N_1697,In_2013,In_2384);
xnor U1698 (N_1698,In_921,In_1390);
xnor U1699 (N_1699,In_874,In_2630);
xnor U1700 (N_1700,In_2336,In_1674);
and U1701 (N_1701,In_2774,In_2590);
nand U1702 (N_1702,In_144,In_2979);
or U1703 (N_1703,In_2367,In_1482);
nand U1704 (N_1704,In_842,In_234);
or U1705 (N_1705,In_2477,In_2210);
nand U1706 (N_1706,In_443,In_2764);
nor U1707 (N_1707,In_721,In_968);
and U1708 (N_1708,In_1659,In_2928);
nor U1709 (N_1709,In_1269,In_1085);
and U1710 (N_1710,In_1614,In_2335);
nor U1711 (N_1711,In_2233,In_2593);
or U1712 (N_1712,In_1162,In_2494);
nand U1713 (N_1713,In_1435,In_88);
or U1714 (N_1714,In_1161,In_2183);
nand U1715 (N_1715,In_2180,In_1898);
nand U1716 (N_1716,In_1293,In_142);
or U1717 (N_1717,In_1244,In_200);
or U1718 (N_1718,In_914,In_1931);
or U1719 (N_1719,In_2687,In_1029);
or U1720 (N_1720,In_292,In_529);
and U1721 (N_1721,In_2629,In_158);
nor U1722 (N_1722,In_2816,In_843);
xnor U1723 (N_1723,In_2070,In_15);
nor U1724 (N_1724,In_885,In_60);
nor U1725 (N_1725,In_2238,In_340);
nor U1726 (N_1726,In_596,In_1845);
nor U1727 (N_1727,In_764,In_2441);
xor U1728 (N_1728,In_991,In_1470);
xor U1729 (N_1729,In_1882,In_1219);
nor U1730 (N_1730,In_2926,In_2032);
nand U1731 (N_1731,In_1199,In_2913);
or U1732 (N_1732,In_1956,In_1025);
nand U1733 (N_1733,In_2662,In_1587);
xor U1734 (N_1734,In_254,In_1517);
nor U1735 (N_1735,In_450,In_2741);
nand U1736 (N_1736,In_437,In_269);
or U1737 (N_1737,In_1541,In_2332);
and U1738 (N_1738,In_2292,In_860);
nand U1739 (N_1739,In_1486,In_2787);
and U1740 (N_1740,In_190,In_537);
xnor U1741 (N_1741,In_2335,In_230);
and U1742 (N_1742,In_1799,In_454);
and U1743 (N_1743,In_1684,In_6);
nand U1744 (N_1744,In_2718,In_480);
or U1745 (N_1745,In_2634,In_96);
xnor U1746 (N_1746,In_1984,In_767);
and U1747 (N_1747,In_2337,In_426);
nand U1748 (N_1748,In_81,In_1014);
xnor U1749 (N_1749,In_1139,In_2373);
xnor U1750 (N_1750,In_48,In_1517);
xor U1751 (N_1751,In_1022,In_370);
nor U1752 (N_1752,In_85,In_2365);
nor U1753 (N_1753,In_67,In_2195);
xor U1754 (N_1754,In_608,In_67);
nand U1755 (N_1755,In_2940,In_2925);
nand U1756 (N_1756,In_1936,In_1340);
or U1757 (N_1757,In_596,In_1860);
and U1758 (N_1758,In_1817,In_911);
nor U1759 (N_1759,In_1503,In_1806);
xnor U1760 (N_1760,In_2648,In_1059);
nand U1761 (N_1761,In_1218,In_1205);
or U1762 (N_1762,In_2136,In_642);
xnor U1763 (N_1763,In_1707,In_1054);
or U1764 (N_1764,In_2,In_2707);
nor U1765 (N_1765,In_1128,In_238);
nand U1766 (N_1766,In_2696,In_2167);
or U1767 (N_1767,In_1411,In_1077);
nand U1768 (N_1768,In_579,In_1090);
xnor U1769 (N_1769,In_931,In_793);
nor U1770 (N_1770,In_1727,In_1797);
and U1771 (N_1771,In_2308,In_2174);
xnor U1772 (N_1772,In_971,In_7);
and U1773 (N_1773,In_2162,In_2542);
and U1774 (N_1774,In_2491,In_28);
and U1775 (N_1775,In_2031,In_1380);
xnor U1776 (N_1776,In_2421,In_949);
xor U1777 (N_1777,In_2802,In_1808);
nand U1778 (N_1778,In_1874,In_1975);
xor U1779 (N_1779,In_2882,In_529);
nor U1780 (N_1780,In_44,In_2813);
or U1781 (N_1781,In_1526,In_1031);
and U1782 (N_1782,In_1339,In_2119);
or U1783 (N_1783,In_2065,In_2754);
nor U1784 (N_1784,In_1247,In_1452);
xnor U1785 (N_1785,In_2556,In_973);
or U1786 (N_1786,In_1489,In_2643);
or U1787 (N_1787,In_1838,In_2930);
and U1788 (N_1788,In_2817,In_86);
or U1789 (N_1789,In_419,In_813);
xnor U1790 (N_1790,In_1058,In_494);
and U1791 (N_1791,In_2521,In_354);
nand U1792 (N_1792,In_215,In_2016);
nand U1793 (N_1793,In_2156,In_1461);
nor U1794 (N_1794,In_2238,In_945);
or U1795 (N_1795,In_835,In_2789);
or U1796 (N_1796,In_1947,In_1905);
xor U1797 (N_1797,In_2144,In_2437);
xor U1798 (N_1798,In_1197,In_2078);
and U1799 (N_1799,In_942,In_328);
xnor U1800 (N_1800,In_1250,In_1704);
xnor U1801 (N_1801,In_2710,In_1374);
nor U1802 (N_1802,In_2659,In_1687);
and U1803 (N_1803,In_1604,In_1831);
nor U1804 (N_1804,In_1940,In_180);
xnor U1805 (N_1805,In_1218,In_1706);
xor U1806 (N_1806,In_1068,In_1514);
nand U1807 (N_1807,In_2356,In_1061);
or U1808 (N_1808,In_993,In_869);
nand U1809 (N_1809,In_1502,In_2812);
and U1810 (N_1810,In_2995,In_1274);
or U1811 (N_1811,In_2087,In_367);
and U1812 (N_1812,In_5,In_2677);
nor U1813 (N_1813,In_1577,In_1933);
xor U1814 (N_1814,In_2380,In_495);
xor U1815 (N_1815,In_1482,In_2140);
nand U1816 (N_1816,In_1340,In_2398);
and U1817 (N_1817,In_1495,In_2122);
and U1818 (N_1818,In_739,In_2554);
and U1819 (N_1819,In_1742,In_45);
nor U1820 (N_1820,In_2709,In_151);
nor U1821 (N_1821,In_1192,In_1111);
nand U1822 (N_1822,In_1215,In_136);
and U1823 (N_1823,In_315,In_2910);
nand U1824 (N_1824,In_1643,In_1070);
xor U1825 (N_1825,In_2039,In_1701);
and U1826 (N_1826,In_1334,In_1517);
nor U1827 (N_1827,In_1346,In_2095);
nand U1828 (N_1828,In_1957,In_951);
nor U1829 (N_1829,In_1363,In_719);
and U1830 (N_1830,In_2199,In_1733);
and U1831 (N_1831,In_128,In_2865);
xnor U1832 (N_1832,In_2775,In_2278);
and U1833 (N_1833,In_2490,In_350);
xor U1834 (N_1834,In_533,In_2764);
or U1835 (N_1835,In_2074,In_47);
nand U1836 (N_1836,In_1380,In_1494);
xnor U1837 (N_1837,In_2005,In_2144);
nor U1838 (N_1838,In_1411,In_1132);
xor U1839 (N_1839,In_2720,In_2122);
xor U1840 (N_1840,In_2515,In_673);
and U1841 (N_1841,In_203,In_358);
and U1842 (N_1842,In_1977,In_416);
or U1843 (N_1843,In_2738,In_1499);
nor U1844 (N_1844,In_2842,In_2817);
or U1845 (N_1845,In_1789,In_584);
and U1846 (N_1846,In_1798,In_696);
or U1847 (N_1847,In_245,In_2988);
nand U1848 (N_1848,In_467,In_1239);
or U1849 (N_1849,In_891,In_1921);
or U1850 (N_1850,In_2118,In_2871);
and U1851 (N_1851,In_1165,In_2737);
nor U1852 (N_1852,In_2003,In_618);
nand U1853 (N_1853,In_115,In_518);
nor U1854 (N_1854,In_2762,In_745);
nand U1855 (N_1855,In_1396,In_42);
xor U1856 (N_1856,In_989,In_1377);
xnor U1857 (N_1857,In_2238,In_2292);
and U1858 (N_1858,In_2598,In_2446);
nand U1859 (N_1859,In_138,In_949);
xnor U1860 (N_1860,In_2189,In_2473);
nand U1861 (N_1861,In_2955,In_214);
and U1862 (N_1862,In_2591,In_1625);
nand U1863 (N_1863,In_1638,In_177);
and U1864 (N_1864,In_1534,In_2266);
nor U1865 (N_1865,In_2203,In_290);
and U1866 (N_1866,In_2241,In_2463);
nor U1867 (N_1867,In_2669,In_2382);
and U1868 (N_1868,In_1350,In_1712);
nor U1869 (N_1869,In_310,In_1252);
nand U1870 (N_1870,In_1888,In_1717);
nor U1871 (N_1871,In_955,In_392);
and U1872 (N_1872,In_1845,In_2476);
nand U1873 (N_1873,In_1586,In_1420);
nand U1874 (N_1874,In_453,In_1985);
nand U1875 (N_1875,In_680,In_209);
xnor U1876 (N_1876,In_1678,In_1614);
or U1877 (N_1877,In_1169,In_2768);
nand U1878 (N_1878,In_2761,In_2752);
xnor U1879 (N_1879,In_922,In_2395);
and U1880 (N_1880,In_301,In_2945);
xnor U1881 (N_1881,In_1779,In_576);
and U1882 (N_1882,In_2900,In_2187);
nand U1883 (N_1883,In_1741,In_518);
or U1884 (N_1884,In_2743,In_652);
nor U1885 (N_1885,In_56,In_654);
nand U1886 (N_1886,In_2077,In_2233);
and U1887 (N_1887,In_1453,In_1070);
xor U1888 (N_1888,In_324,In_1293);
nor U1889 (N_1889,In_2483,In_2142);
or U1890 (N_1890,In_810,In_1864);
or U1891 (N_1891,In_2718,In_2751);
or U1892 (N_1892,In_801,In_140);
and U1893 (N_1893,In_1775,In_2977);
and U1894 (N_1894,In_221,In_1014);
nand U1895 (N_1895,In_1504,In_379);
nand U1896 (N_1896,In_365,In_2839);
nand U1897 (N_1897,In_217,In_739);
or U1898 (N_1898,In_539,In_2199);
or U1899 (N_1899,In_90,In_2641);
and U1900 (N_1900,In_2764,In_0);
nor U1901 (N_1901,In_2347,In_2656);
xnor U1902 (N_1902,In_1849,In_2065);
nand U1903 (N_1903,In_1476,In_2295);
nor U1904 (N_1904,In_196,In_949);
xor U1905 (N_1905,In_2622,In_2654);
nor U1906 (N_1906,In_2909,In_1938);
nand U1907 (N_1907,In_1208,In_999);
nor U1908 (N_1908,In_2633,In_1071);
xnor U1909 (N_1909,In_180,In_101);
xor U1910 (N_1910,In_1358,In_2780);
nand U1911 (N_1911,In_1980,In_1446);
nor U1912 (N_1912,In_91,In_73);
or U1913 (N_1913,In_111,In_25);
and U1914 (N_1914,In_2712,In_270);
and U1915 (N_1915,In_122,In_2083);
and U1916 (N_1916,In_2527,In_178);
nor U1917 (N_1917,In_497,In_77);
and U1918 (N_1918,In_2313,In_2219);
or U1919 (N_1919,In_797,In_1843);
and U1920 (N_1920,In_116,In_703);
nor U1921 (N_1921,In_2153,In_618);
xor U1922 (N_1922,In_1227,In_675);
and U1923 (N_1923,In_675,In_1685);
and U1924 (N_1924,In_731,In_2492);
and U1925 (N_1925,In_806,In_1769);
nor U1926 (N_1926,In_1810,In_2155);
nor U1927 (N_1927,In_354,In_1411);
xor U1928 (N_1928,In_361,In_284);
or U1929 (N_1929,In_865,In_1024);
and U1930 (N_1930,In_1678,In_1288);
or U1931 (N_1931,In_1406,In_2823);
and U1932 (N_1932,In_2970,In_370);
xor U1933 (N_1933,In_2209,In_1138);
or U1934 (N_1934,In_1167,In_2090);
xnor U1935 (N_1935,In_2530,In_2815);
and U1936 (N_1936,In_845,In_2170);
or U1937 (N_1937,In_723,In_641);
nand U1938 (N_1938,In_2874,In_2550);
or U1939 (N_1939,In_1790,In_3);
and U1940 (N_1940,In_1647,In_1242);
xnor U1941 (N_1941,In_1547,In_888);
xor U1942 (N_1942,In_790,In_1640);
nor U1943 (N_1943,In_1330,In_1355);
nand U1944 (N_1944,In_1981,In_1404);
xor U1945 (N_1945,In_121,In_2776);
xnor U1946 (N_1946,In_1782,In_1695);
and U1947 (N_1947,In_1229,In_503);
nor U1948 (N_1948,In_1782,In_1647);
or U1949 (N_1949,In_1706,In_758);
nand U1950 (N_1950,In_2600,In_992);
xnor U1951 (N_1951,In_1619,In_2652);
and U1952 (N_1952,In_84,In_2033);
xnor U1953 (N_1953,In_2073,In_2701);
or U1954 (N_1954,In_2593,In_2023);
nor U1955 (N_1955,In_2073,In_2056);
nand U1956 (N_1956,In_881,In_1066);
or U1957 (N_1957,In_688,In_2475);
and U1958 (N_1958,In_1966,In_709);
xor U1959 (N_1959,In_355,In_2152);
and U1960 (N_1960,In_114,In_677);
nor U1961 (N_1961,In_1623,In_89);
or U1962 (N_1962,In_2626,In_2701);
and U1963 (N_1963,In_245,In_1373);
nor U1964 (N_1964,In_1810,In_2453);
nor U1965 (N_1965,In_2398,In_1833);
and U1966 (N_1966,In_1628,In_677);
nand U1967 (N_1967,In_1645,In_2136);
or U1968 (N_1968,In_799,In_730);
nand U1969 (N_1969,In_742,In_2427);
and U1970 (N_1970,In_2799,In_2447);
or U1971 (N_1971,In_2336,In_1466);
nor U1972 (N_1972,In_2599,In_1080);
xnor U1973 (N_1973,In_2598,In_1903);
nor U1974 (N_1974,In_292,In_2900);
nand U1975 (N_1975,In_2028,In_1855);
nand U1976 (N_1976,In_1074,In_2068);
nor U1977 (N_1977,In_1603,In_272);
or U1978 (N_1978,In_2847,In_1323);
nor U1979 (N_1979,In_1254,In_1347);
xnor U1980 (N_1980,In_1526,In_192);
nand U1981 (N_1981,In_1306,In_2769);
or U1982 (N_1982,In_1774,In_2515);
nand U1983 (N_1983,In_1579,In_2087);
nand U1984 (N_1984,In_961,In_559);
nor U1985 (N_1985,In_1780,In_234);
nand U1986 (N_1986,In_1056,In_2585);
or U1987 (N_1987,In_1188,In_1527);
nor U1988 (N_1988,In_1473,In_70);
xnor U1989 (N_1989,In_2656,In_2082);
or U1990 (N_1990,In_2658,In_2700);
and U1991 (N_1991,In_1182,In_1313);
nor U1992 (N_1992,In_1576,In_1957);
or U1993 (N_1993,In_1509,In_72);
nand U1994 (N_1994,In_904,In_838);
or U1995 (N_1995,In_2849,In_1494);
xor U1996 (N_1996,In_449,In_933);
or U1997 (N_1997,In_2410,In_510);
or U1998 (N_1998,In_856,In_2811);
and U1999 (N_1999,In_2647,In_14);
nor U2000 (N_2000,In_557,In_1204);
nor U2001 (N_2001,In_1258,In_1130);
and U2002 (N_2002,In_735,In_1626);
or U2003 (N_2003,In_2600,In_2500);
or U2004 (N_2004,In_450,In_1593);
nand U2005 (N_2005,In_1221,In_2800);
nor U2006 (N_2006,In_613,In_2945);
or U2007 (N_2007,In_2954,In_2161);
nand U2008 (N_2008,In_2133,In_2176);
or U2009 (N_2009,In_1346,In_2618);
xnor U2010 (N_2010,In_2141,In_2100);
nor U2011 (N_2011,In_141,In_874);
xor U2012 (N_2012,In_2929,In_2380);
nor U2013 (N_2013,In_144,In_1792);
or U2014 (N_2014,In_2198,In_1701);
or U2015 (N_2015,In_2547,In_2730);
or U2016 (N_2016,In_2248,In_2296);
xnor U2017 (N_2017,In_2537,In_609);
xnor U2018 (N_2018,In_374,In_476);
and U2019 (N_2019,In_435,In_1843);
xnor U2020 (N_2020,In_2424,In_1982);
and U2021 (N_2021,In_2083,In_1544);
xor U2022 (N_2022,In_550,In_1408);
xnor U2023 (N_2023,In_1759,In_2754);
nor U2024 (N_2024,In_1743,In_1007);
and U2025 (N_2025,In_2250,In_1323);
and U2026 (N_2026,In_1196,In_1209);
nand U2027 (N_2027,In_1732,In_2093);
or U2028 (N_2028,In_2383,In_1257);
xor U2029 (N_2029,In_2661,In_2189);
and U2030 (N_2030,In_2509,In_602);
nor U2031 (N_2031,In_2763,In_859);
nor U2032 (N_2032,In_1812,In_747);
nand U2033 (N_2033,In_369,In_455);
nand U2034 (N_2034,In_2794,In_1981);
or U2035 (N_2035,In_2135,In_2524);
and U2036 (N_2036,In_1080,In_1508);
nor U2037 (N_2037,In_2769,In_770);
xnor U2038 (N_2038,In_1922,In_163);
or U2039 (N_2039,In_2799,In_255);
and U2040 (N_2040,In_1656,In_2857);
xnor U2041 (N_2041,In_1686,In_1457);
nand U2042 (N_2042,In_2928,In_13);
nor U2043 (N_2043,In_2352,In_2351);
and U2044 (N_2044,In_1285,In_313);
nand U2045 (N_2045,In_2150,In_2510);
nand U2046 (N_2046,In_2268,In_2562);
or U2047 (N_2047,In_2704,In_1351);
nand U2048 (N_2048,In_975,In_2634);
or U2049 (N_2049,In_1830,In_26);
nand U2050 (N_2050,In_546,In_1576);
or U2051 (N_2051,In_2060,In_2346);
or U2052 (N_2052,In_940,In_1612);
nor U2053 (N_2053,In_1535,In_2447);
or U2054 (N_2054,In_750,In_209);
and U2055 (N_2055,In_2474,In_1335);
or U2056 (N_2056,In_2050,In_2730);
or U2057 (N_2057,In_79,In_2731);
and U2058 (N_2058,In_1801,In_2432);
nor U2059 (N_2059,In_2017,In_474);
nor U2060 (N_2060,In_1659,In_1272);
and U2061 (N_2061,In_280,In_441);
nor U2062 (N_2062,In_681,In_58);
xnor U2063 (N_2063,In_1110,In_2647);
nand U2064 (N_2064,In_2222,In_1951);
nand U2065 (N_2065,In_1284,In_1048);
nor U2066 (N_2066,In_2580,In_892);
or U2067 (N_2067,In_1606,In_713);
or U2068 (N_2068,In_2722,In_1993);
nor U2069 (N_2069,In_572,In_1746);
or U2070 (N_2070,In_2844,In_2354);
and U2071 (N_2071,In_2130,In_1730);
nor U2072 (N_2072,In_1299,In_1140);
and U2073 (N_2073,In_836,In_2864);
nand U2074 (N_2074,In_830,In_1290);
nand U2075 (N_2075,In_2759,In_843);
nand U2076 (N_2076,In_2997,In_1800);
nand U2077 (N_2077,In_886,In_179);
or U2078 (N_2078,In_2816,In_749);
and U2079 (N_2079,In_345,In_1245);
and U2080 (N_2080,In_2655,In_566);
nand U2081 (N_2081,In_1367,In_1353);
or U2082 (N_2082,In_2193,In_2784);
or U2083 (N_2083,In_1369,In_1347);
xor U2084 (N_2084,In_861,In_1377);
xor U2085 (N_2085,In_376,In_1302);
nand U2086 (N_2086,In_563,In_1273);
and U2087 (N_2087,In_2222,In_1583);
nor U2088 (N_2088,In_2462,In_1601);
xor U2089 (N_2089,In_40,In_194);
nor U2090 (N_2090,In_1228,In_2791);
nand U2091 (N_2091,In_182,In_1867);
or U2092 (N_2092,In_2607,In_2050);
or U2093 (N_2093,In_1171,In_1735);
and U2094 (N_2094,In_2391,In_873);
xnor U2095 (N_2095,In_1184,In_1966);
or U2096 (N_2096,In_512,In_947);
nand U2097 (N_2097,In_2480,In_214);
nand U2098 (N_2098,In_1385,In_1738);
xnor U2099 (N_2099,In_345,In_778);
and U2100 (N_2100,In_1129,In_2478);
and U2101 (N_2101,In_1208,In_2417);
and U2102 (N_2102,In_602,In_328);
and U2103 (N_2103,In_592,In_2288);
xnor U2104 (N_2104,In_4,In_1397);
or U2105 (N_2105,In_1642,In_2084);
nor U2106 (N_2106,In_1993,In_1121);
nand U2107 (N_2107,In_315,In_271);
or U2108 (N_2108,In_1143,In_2527);
and U2109 (N_2109,In_2924,In_2243);
nand U2110 (N_2110,In_2747,In_2558);
xor U2111 (N_2111,In_352,In_944);
xor U2112 (N_2112,In_565,In_2789);
or U2113 (N_2113,In_399,In_1263);
nand U2114 (N_2114,In_2545,In_1024);
or U2115 (N_2115,In_1172,In_2942);
or U2116 (N_2116,In_466,In_938);
xor U2117 (N_2117,In_1479,In_1230);
and U2118 (N_2118,In_2823,In_1221);
and U2119 (N_2119,In_1495,In_2160);
xor U2120 (N_2120,In_2334,In_1042);
or U2121 (N_2121,In_356,In_732);
nand U2122 (N_2122,In_90,In_658);
xnor U2123 (N_2123,In_1034,In_2906);
xor U2124 (N_2124,In_31,In_644);
and U2125 (N_2125,In_58,In_2109);
and U2126 (N_2126,In_1418,In_2783);
nand U2127 (N_2127,In_762,In_1294);
or U2128 (N_2128,In_2843,In_1802);
nand U2129 (N_2129,In_202,In_2213);
and U2130 (N_2130,In_812,In_2668);
nor U2131 (N_2131,In_173,In_844);
nand U2132 (N_2132,In_1729,In_12);
and U2133 (N_2133,In_818,In_300);
nand U2134 (N_2134,In_2445,In_230);
nor U2135 (N_2135,In_1303,In_1026);
nand U2136 (N_2136,In_297,In_2290);
nand U2137 (N_2137,In_2817,In_827);
nand U2138 (N_2138,In_479,In_2012);
or U2139 (N_2139,In_1259,In_458);
xor U2140 (N_2140,In_233,In_1939);
nor U2141 (N_2141,In_227,In_2474);
nand U2142 (N_2142,In_881,In_2339);
xnor U2143 (N_2143,In_774,In_985);
nand U2144 (N_2144,In_2254,In_119);
and U2145 (N_2145,In_1652,In_1644);
nand U2146 (N_2146,In_2307,In_2124);
xor U2147 (N_2147,In_86,In_990);
nor U2148 (N_2148,In_538,In_5);
or U2149 (N_2149,In_126,In_2023);
or U2150 (N_2150,In_2509,In_1776);
and U2151 (N_2151,In_338,In_2129);
xor U2152 (N_2152,In_1927,In_924);
or U2153 (N_2153,In_859,In_2752);
nand U2154 (N_2154,In_279,In_184);
xor U2155 (N_2155,In_402,In_1717);
xnor U2156 (N_2156,In_801,In_2395);
and U2157 (N_2157,In_1913,In_2124);
or U2158 (N_2158,In_1719,In_982);
or U2159 (N_2159,In_2208,In_2682);
and U2160 (N_2160,In_1269,In_2218);
xnor U2161 (N_2161,In_2738,In_642);
and U2162 (N_2162,In_147,In_2841);
nand U2163 (N_2163,In_514,In_826);
xor U2164 (N_2164,In_1992,In_2887);
and U2165 (N_2165,In_2501,In_2774);
or U2166 (N_2166,In_1005,In_2619);
nand U2167 (N_2167,In_1367,In_1966);
or U2168 (N_2168,In_418,In_44);
nand U2169 (N_2169,In_2364,In_839);
nand U2170 (N_2170,In_841,In_2725);
nand U2171 (N_2171,In_1929,In_415);
nor U2172 (N_2172,In_1411,In_1061);
and U2173 (N_2173,In_741,In_1430);
nand U2174 (N_2174,In_1754,In_238);
and U2175 (N_2175,In_1453,In_1926);
or U2176 (N_2176,In_262,In_1649);
xor U2177 (N_2177,In_851,In_228);
nand U2178 (N_2178,In_349,In_569);
nand U2179 (N_2179,In_1525,In_2636);
or U2180 (N_2180,In_300,In_587);
nand U2181 (N_2181,In_1998,In_1597);
nor U2182 (N_2182,In_534,In_1759);
nand U2183 (N_2183,In_2307,In_1486);
nand U2184 (N_2184,In_291,In_165);
xor U2185 (N_2185,In_2299,In_511);
nand U2186 (N_2186,In_341,In_964);
nor U2187 (N_2187,In_1447,In_2945);
or U2188 (N_2188,In_2180,In_2283);
nand U2189 (N_2189,In_142,In_2661);
nor U2190 (N_2190,In_2012,In_2206);
nand U2191 (N_2191,In_1844,In_2817);
nor U2192 (N_2192,In_650,In_2654);
nand U2193 (N_2193,In_2710,In_1615);
nor U2194 (N_2194,In_1592,In_2430);
nor U2195 (N_2195,In_92,In_2133);
nand U2196 (N_2196,In_2053,In_795);
nor U2197 (N_2197,In_1274,In_2515);
nand U2198 (N_2198,In_1561,In_1266);
nand U2199 (N_2199,In_790,In_1565);
nor U2200 (N_2200,In_1202,In_1414);
and U2201 (N_2201,In_2346,In_765);
nand U2202 (N_2202,In_2461,In_1285);
xor U2203 (N_2203,In_321,In_324);
or U2204 (N_2204,In_795,In_2250);
and U2205 (N_2205,In_2893,In_2486);
nand U2206 (N_2206,In_269,In_761);
nor U2207 (N_2207,In_1974,In_2745);
and U2208 (N_2208,In_2889,In_840);
nand U2209 (N_2209,In_874,In_1700);
xnor U2210 (N_2210,In_1214,In_2803);
xor U2211 (N_2211,In_325,In_1625);
nor U2212 (N_2212,In_1674,In_711);
xnor U2213 (N_2213,In_2870,In_925);
nand U2214 (N_2214,In_373,In_1050);
or U2215 (N_2215,In_2365,In_1003);
or U2216 (N_2216,In_1100,In_1331);
or U2217 (N_2217,In_2726,In_832);
nor U2218 (N_2218,In_133,In_570);
nand U2219 (N_2219,In_128,In_1344);
nand U2220 (N_2220,In_2259,In_1282);
and U2221 (N_2221,In_2377,In_1302);
xor U2222 (N_2222,In_2618,In_770);
or U2223 (N_2223,In_2734,In_2462);
or U2224 (N_2224,In_1201,In_1733);
nor U2225 (N_2225,In_751,In_65);
or U2226 (N_2226,In_1674,In_1568);
or U2227 (N_2227,In_506,In_1633);
or U2228 (N_2228,In_1882,In_2815);
nor U2229 (N_2229,In_115,In_2790);
xnor U2230 (N_2230,In_2298,In_2749);
and U2231 (N_2231,In_669,In_1410);
xor U2232 (N_2232,In_1890,In_1235);
xnor U2233 (N_2233,In_2391,In_2719);
or U2234 (N_2234,In_149,In_759);
nor U2235 (N_2235,In_2539,In_2940);
nand U2236 (N_2236,In_1495,In_2381);
xor U2237 (N_2237,In_516,In_1553);
or U2238 (N_2238,In_1043,In_2048);
xor U2239 (N_2239,In_79,In_876);
or U2240 (N_2240,In_2442,In_1930);
and U2241 (N_2241,In_1602,In_552);
nor U2242 (N_2242,In_2453,In_2009);
or U2243 (N_2243,In_1424,In_1913);
or U2244 (N_2244,In_1182,In_1827);
and U2245 (N_2245,In_1175,In_2861);
nor U2246 (N_2246,In_1817,In_33);
nor U2247 (N_2247,In_1912,In_2079);
or U2248 (N_2248,In_2944,In_1370);
or U2249 (N_2249,In_2995,In_1162);
xor U2250 (N_2250,In_659,In_98);
and U2251 (N_2251,In_2991,In_57);
xnor U2252 (N_2252,In_1171,In_1039);
nor U2253 (N_2253,In_447,In_190);
nor U2254 (N_2254,In_24,In_2303);
and U2255 (N_2255,In_1181,In_80);
nor U2256 (N_2256,In_630,In_2281);
nor U2257 (N_2257,In_2670,In_2942);
nor U2258 (N_2258,In_1493,In_2476);
and U2259 (N_2259,In_1468,In_1411);
or U2260 (N_2260,In_1291,In_2408);
and U2261 (N_2261,In_898,In_1280);
xor U2262 (N_2262,In_2613,In_2457);
and U2263 (N_2263,In_1217,In_864);
nand U2264 (N_2264,In_2486,In_2153);
nor U2265 (N_2265,In_2183,In_310);
xnor U2266 (N_2266,In_123,In_1703);
nor U2267 (N_2267,In_1954,In_1993);
nor U2268 (N_2268,In_1018,In_827);
nand U2269 (N_2269,In_446,In_1984);
xor U2270 (N_2270,In_1343,In_2353);
xnor U2271 (N_2271,In_1605,In_1399);
nor U2272 (N_2272,In_1141,In_275);
or U2273 (N_2273,In_1990,In_1917);
nor U2274 (N_2274,In_1996,In_57);
or U2275 (N_2275,In_1231,In_804);
nor U2276 (N_2276,In_1568,In_1043);
or U2277 (N_2277,In_2829,In_859);
and U2278 (N_2278,In_2149,In_1335);
and U2279 (N_2279,In_295,In_358);
nor U2280 (N_2280,In_2003,In_2215);
and U2281 (N_2281,In_2773,In_2062);
xor U2282 (N_2282,In_1086,In_2700);
xor U2283 (N_2283,In_1700,In_2690);
and U2284 (N_2284,In_1580,In_1930);
nor U2285 (N_2285,In_2236,In_59);
nor U2286 (N_2286,In_2712,In_2136);
nand U2287 (N_2287,In_1966,In_317);
or U2288 (N_2288,In_1852,In_2254);
nor U2289 (N_2289,In_2058,In_2745);
xnor U2290 (N_2290,In_2241,In_569);
nor U2291 (N_2291,In_2469,In_2144);
xor U2292 (N_2292,In_1681,In_241);
and U2293 (N_2293,In_1820,In_1654);
nand U2294 (N_2294,In_2117,In_1352);
and U2295 (N_2295,In_276,In_2365);
and U2296 (N_2296,In_1196,In_2368);
nor U2297 (N_2297,In_572,In_1330);
nor U2298 (N_2298,In_619,In_2551);
xnor U2299 (N_2299,In_806,In_1891);
xor U2300 (N_2300,In_2172,In_531);
nand U2301 (N_2301,In_1531,In_2983);
nor U2302 (N_2302,In_2752,In_171);
and U2303 (N_2303,In_2975,In_2012);
and U2304 (N_2304,In_326,In_2652);
xor U2305 (N_2305,In_1733,In_412);
and U2306 (N_2306,In_2307,In_1591);
or U2307 (N_2307,In_337,In_161);
xor U2308 (N_2308,In_2678,In_2899);
xor U2309 (N_2309,In_1618,In_1748);
xnor U2310 (N_2310,In_2199,In_1498);
nand U2311 (N_2311,In_2682,In_1576);
or U2312 (N_2312,In_1930,In_649);
nor U2313 (N_2313,In_2775,In_951);
and U2314 (N_2314,In_1244,In_1545);
and U2315 (N_2315,In_2208,In_790);
nor U2316 (N_2316,In_2368,In_2629);
nand U2317 (N_2317,In_2983,In_218);
nor U2318 (N_2318,In_2115,In_1781);
or U2319 (N_2319,In_2163,In_2238);
xor U2320 (N_2320,In_2920,In_2267);
nor U2321 (N_2321,In_293,In_716);
or U2322 (N_2322,In_654,In_2986);
and U2323 (N_2323,In_617,In_2597);
or U2324 (N_2324,In_367,In_2163);
nor U2325 (N_2325,In_2450,In_404);
or U2326 (N_2326,In_1253,In_495);
nor U2327 (N_2327,In_1537,In_1433);
and U2328 (N_2328,In_93,In_2948);
or U2329 (N_2329,In_1415,In_469);
xor U2330 (N_2330,In_697,In_1504);
xnor U2331 (N_2331,In_1103,In_2694);
and U2332 (N_2332,In_1893,In_1099);
xor U2333 (N_2333,In_593,In_2859);
nor U2334 (N_2334,In_1875,In_941);
nand U2335 (N_2335,In_1209,In_2921);
nor U2336 (N_2336,In_2234,In_156);
nand U2337 (N_2337,In_2131,In_2980);
or U2338 (N_2338,In_2802,In_2097);
xnor U2339 (N_2339,In_122,In_2657);
xor U2340 (N_2340,In_444,In_1716);
and U2341 (N_2341,In_2807,In_486);
xnor U2342 (N_2342,In_923,In_315);
nor U2343 (N_2343,In_921,In_50);
nor U2344 (N_2344,In_750,In_177);
or U2345 (N_2345,In_2211,In_766);
nor U2346 (N_2346,In_1646,In_1502);
xor U2347 (N_2347,In_2844,In_1774);
nand U2348 (N_2348,In_461,In_2198);
nand U2349 (N_2349,In_2373,In_595);
xor U2350 (N_2350,In_1042,In_1349);
nor U2351 (N_2351,In_2235,In_327);
nand U2352 (N_2352,In_2902,In_826);
and U2353 (N_2353,In_275,In_566);
xnor U2354 (N_2354,In_1873,In_365);
and U2355 (N_2355,In_2975,In_2300);
and U2356 (N_2356,In_1087,In_481);
xor U2357 (N_2357,In_1996,In_2538);
or U2358 (N_2358,In_2422,In_1853);
nor U2359 (N_2359,In_364,In_2137);
or U2360 (N_2360,In_426,In_2136);
or U2361 (N_2361,In_2266,In_1099);
and U2362 (N_2362,In_2115,In_2673);
nand U2363 (N_2363,In_462,In_1116);
and U2364 (N_2364,In_1224,In_2837);
or U2365 (N_2365,In_2840,In_499);
and U2366 (N_2366,In_1734,In_1558);
xnor U2367 (N_2367,In_857,In_1747);
xor U2368 (N_2368,In_256,In_2757);
or U2369 (N_2369,In_2541,In_2702);
nand U2370 (N_2370,In_258,In_671);
and U2371 (N_2371,In_1618,In_2570);
nor U2372 (N_2372,In_2974,In_388);
nor U2373 (N_2373,In_2225,In_1242);
xor U2374 (N_2374,In_1662,In_2559);
and U2375 (N_2375,In_207,In_1733);
xnor U2376 (N_2376,In_1250,In_2547);
and U2377 (N_2377,In_1735,In_2987);
or U2378 (N_2378,In_1121,In_1275);
nand U2379 (N_2379,In_280,In_2908);
nand U2380 (N_2380,In_496,In_1565);
or U2381 (N_2381,In_618,In_2438);
nor U2382 (N_2382,In_560,In_1949);
or U2383 (N_2383,In_2259,In_629);
or U2384 (N_2384,In_2271,In_1286);
and U2385 (N_2385,In_879,In_1633);
nand U2386 (N_2386,In_1983,In_1220);
nor U2387 (N_2387,In_1659,In_1150);
xor U2388 (N_2388,In_2173,In_1417);
and U2389 (N_2389,In_2695,In_1382);
or U2390 (N_2390,In_1691,In_1763);
or U2391 (N_2391,In_955,In_680);
or U2392 (N_2392,In_2947,In_2555);
nor U2393 (N_2393,In_1142,In_1004);
and U2394 (N_2394,In_2809,In_1947);
or U2395 (N_2395,In_2383,In_1058);
nand U2396 (N_2396,In_2424,In_2294);
or U2397 (N_2397,In_448,In_216);
xnor U2398 (N_2398,In_2095,In_2331);
nand U2399 (N_2399,In_2671,In_2289);
nand U2400 (N_2400,In_2152,In_40);
nor U2401 (N_2401,In_2931,In_2131);
nor U2402 (N_2402,In_702,In_2630);
nand U2403 (N_2403,In_234,In_1140);
nor U2404 (N_2404,In_1560,In_1586);
xnor U2405 (N_2405,In_693,In_2726);
nand U2406 (N_2406,In_1942,In_527);
xor U2407 (N_2407,In_1024,In_404);
and U2408 (N_2408,In_1345,In_2743);
nor U2409 (N_2409,In_1895,In_1974);
nor U2410 (N_2410,In_1464,In_2513);
nand U2411 (N_2411,In_978,In_1619);
and U2412 (N_2412,In_1450,In_207);
xnor U2413 (N_2413,In_1174,In_669);
nand U2414 (N_2414,In_478,In_195);
nand U2415 (N_2415,In_2090,In_1891);
nand U2416 (N_2416,In_2064,In_313);
xnor U2417 (N_2417,In_1808,In_336);
xnor U2418 (N_2418,In_2321,In_2237);
xor U2419 (N_2419,In_2687,In_2212);
nor U2420 (N_2420,In_912,In_2248);
and U2421 (N_2421,In_361,In_2226);
nand U2422 (N_2422,In_1788,In_2181);
and U2423 (N_2423,In_1521,In_21);
or U2424 (N_2424,In_1899,In_2934);
nor U2425 (N_2425,In_2612,In_1652);
nand U2426 (N_2426,In_2545,In_2213);
nor U2427 (N_2427,In_645,In_158);
nor U2428 (N_2428,In_101,In_345);
and U2429 (N_2429,In_889,In_273);
and U2430 (N_2430,In_524,In_1524);
and U2431 (N_2431,In_1061,In_994);
nor U2432 (N_2432,In_1468,In_1166);
xor U2433 (N_2433,In_2065,In_41);
or U2434 (N_2434,In_259,In_2247);
and U2435 (N_2435,In_2573,In_2419);
xnor U2436 (N_2436,In_1270,In_1802);
or U2437 (N_2437,In_543,In_1738);
and U2438 (N_2438,In_1099,In_899);
and U2439 (N_2439,In_1404,In_418);
or U2440 (N_2440,In_1568,In_95);
nor U2441 (N_2441,In_1791,In_2172);
nor U2442 (N_2442,In_990,In_1639);
or U2443 (N_2443,In_354,In_483);
nand U2444 (N_2444,In_805,In_2975);
or U2445 (N_2445,In_1533,In_2097);
nand U2446 (N_2446,In_2288,In_1933);
nand U2447 (N_2447,In_1369,In_2520);
or U2448 (N_2448,In_1730,In_1477);
and U2449 (N_2449,In_1476,In_1794);
and U2450 (N_2450,In_634,In_366);
or U2451 (N_2451,In_2783,In_2859);
nand U2452 (N_2452,In_2910,In_2403);
or U2453 (N_2453,In_2569,In_2970);
xnor U2454 (N_2454,In_2190,In_2186);
xor U2455 (N_2455,In_2403,In_117);
xnor U2456 (N_2456,In_2328,In_899);
or U2457 (N_2457,In_1528,In_1932);
xnor U2458 (N_2458,In_1025,In_2858);
nand U2459 (N_2459,In_888,In_163);
xnor U2460 (N_2460,In_1031,In_2652);
or U2461 (N_2461,In_209,In_819);
nand U2462 (N_2462,In_1688,In_747);
and U2463 (N_2463,In_2940,In_148);
nand U2464 (N_2464,In_252,In_2891);
xnor U2465 (N_2465,In_1922,In_1885);
nand U2466 (N_2466,In_819,In_2510);
nand U2467 (N_2467,In_2855,In_1212);
nand U2468 (N_2468,In_2453,In_2568);
and U2469 (N_2469,In_2767,In_703);
and U2470 (N_2470,In_2219,In_1608);
and U2471 (N_2471,In_1511,In_1113);
nand U2472 (N_2472,In_291,In_820);
xnor U2473 (N_2473,In_2169,In_1483);
nand U2474 (N_2474,In_1254,In_754);
or U2475 (N_2475,In_862,In_956);
nor U2476 (N_2476,In_2427,In_1920);
nor U2477 (N_2477,In_2435,In_1667);
and U2478 (N_2478,In_2298,In_2343);
and U2479 (N_2479,In_399,In_1377);
nor U2480 (N_2480,In_1615,In_1160);
xor U2481 (N_2481,In_1691,In_524);
xnor U2482 (N_2482,In_2445,In_1584);
nor U2483 (N_2483,In_1254,In_1766);
xnor U2484 (N_2484,In_2767,In_665);
nor U2485 (N_2485,In_1762,In_2686);
nand U2486 (N_2486,In_2054,In_2513);
and U2487 (N_2487,In_1287,In_2928);
nor U2488 (N_2488,In_563,In_1197);
nor U2489 (N_2489,In_211,In_1948);
nand U2490 (N_2490,In_1582,In_1952);
nand U2491 (N_2491,In_2687,In_536);
or U2492 (N_2492,In_1357,In_583);
and U2493 (N_2493,In_1062,In_2650);
xnor U2494 (N_2494,In_1087,In_775);
or U2495 (N_2495,In_2719,In_508);
nand U2496 (N_2496,In_167,In_556);
nor U2497 (N_2497,In_2740,In_2149);
or U2498 (N_2498,In_691,In_1881);
or U2499 (N_2499,In_1823,In_1717);
or U2500 (N_2500,In_1004,In_2196);
nor U2501 (N_2501,In_741,In_516);
nor U2502 (N_2502,In_1281,In_1500);
nor U2503 (N_2503,In_2865,In_2657);
or U2504 (N_2504,In_1998,In_2261);
or U2505 (N_2505,In_2133,In_2179);
xnor U2506 (N_2506,In_1782,In_97);
nor U2507 (N_2507,In_2545,In_852);
nor U2508 (N_2508,In_2381,In_2080);
or U2509 (N_2509,In_1624,In_830);
or U2510 (N_2510,In_603,In_1306);
and U2511 (N_2511,In_1194,In_1219);
nand U2512 (N_2512,In_1556,In_1725);
nand U2513 (N_2513,In_1949,In_436);
nor U2514 (N_2514,In_2435,In_1141);
nand U2515 (N_2515,In_656,In_926);
xnor U2516 (N_2516,In_1715,In_1766);
xor U2517 (N_2517,In_2270,In_2433);
or U2518 (N_2518,In_1728,In_2893);
xor U2519 (N_2519,In_689,In_239);
xnor U2520 (N_2520,In_2599,In_2758);
and U2521 (N_2521,In_2579,In_2488);
nor U2522 (N_2522,In_667,In_2398);
nand U2523 (N_2523,In_1789,In_207);
nor U2524 (N_2524,In_1652,In_162);
xnor U2525 (N_2525,In_1726,In_409);
nor U2526 (N_2526,In_1239,In_2250);
nand U2527 (N_2527,In_2596,In_807);
nand U2528 (N_2528,In_937,In_2699);
nand U2529 (N_2529,In_2496,In_1588);
or U2530 (N_2530,In_2168,In_1530);
xnor U2531 (N_2531,In_187,In_606);
or U2532 (N_2532,In_133,In_2279);
and U2533 (N_2533,In_163,In_2169);
nor U2534 (N_2534,In_705,In_762);
or U2535 (N_2535,In_1600,In_290);
nor U2536 (N_2536,In_2621,In_1630);
or U2537 (N_2537,In_2114,In_1436);
nor U2538 (N_2538,In_305,In_1119);
nand U2539 (N_2539,In_1061,In_1852);
and U2540 (N_2540,In_2284,In_2712);
nand U2541 (N_2541,In_2935,In_1731);
and U2542 (N_2542,In_2591,In_2957);
xor U2543 (N_2543,In_1817,In_2815);
and U2544 (N_2544,In_2570,In_1728);
or U2545 (N_2545,In_1406,In_2336);
and U2546 (N_2546,In_655,In_2770);
xor U2547 (N_2547,In_436,In_606);
and U2548 (N_2548,In_275,In_37);
and U2549 (N_2549,In_846,In_2806);
or U2550 (N_2550,In_1005,In_2025);
and U2551 (N_2551,In_2928,In_346);
nor U2552 (N_2552,In_604,In_1026);
nand U2553 (N_2553,In_1539,In_533);
xor U2554 (N_2554,In_1524,In_268);
nor U2555 (N_2555,In_1394,In_2412);
nand U2556 (N_2556,In_2712,In_742);
or U2557 (N_2557,In_669,In_230);
xor U2558 (N_2558,In_398,In_2564);
nand U2559 (N_2559,In_744,In_1340);
nor U2560 (N_2560,In_1776,In_1477);
nand U2561 (N_2561,In_1639,In_191);
or U2562 (N_2562,In_125,In_2716);
nor U2563 (N_2563,In_2831,In_2428);
nand U2564 (N_2564,In_2263,In_1904);
nand U2565 (N_2565,In_1774,In_1635);
nand U2566 (N_2566,In_91,In_1243);
and U2567 (N_2567,In_1178,In_1895);
nand U2568 (N_2568,In_2182,In_1623);
nand U2569 (N_2569,In_2246,In_2213);
nand U2570 (N_2570,In_800,In_2324);
xnor U2571 (N_2571,In_679,In_1859);
and U2572 (N_2572,In_1759,In_2988);
nor U2573 (N_2573,In_1783,In_2819);
and U2574 (N_2574,In_112,In_780);
nand U2575 (N_2575,In_350,In_1426);
and U2576 (N_2576,In_1445,In_847);
nand U2577 (N_2577,In_347,In_852);
and U2578 (N_2578,In_345,In_2907);
and U2579 (N_2579,In_2643,In_676);
xnor U2580 (N_2580,In_2884,In_1651);
nor U2581 (N_2581,In_1878,In_1721);
and U2582 (N_2582,In_1677,In_2268);
or U2583 (N_2583,In_2102,In_1866);
nand U2584 (N_2584,In_949,In_2793);
nor U2585 (N_2585,In_66,In_2243);
nor U2586 (N_2586,In_2365,In_2492);
and U2587 (N_2587,In_1228,In_213);
or U2588 (N_2588,In_1300,In_2959);
nor U2589 (N_2589,In_1477,In_1509);
xnor U2590 (N_2590,In_1878,In_147);
nand U2591 (N_2591,In_288,In_1163);
nand U2592 (N_2592,In_1984,In_463);
nand U2593 (N_2593,In_302,In_2528);
nand U2594 (N_2594,In_2883,In_2924);
or U2595 (N_2595,In_1165,In_701);
xor U2596 (N_2596,In_2099,In_2052);
xnor U2597 (N_2597,In_1651,In_949);
nand U2598 (N_2598,In_42,In_1863);
and U2599 (N_2599,In_2556,In_2078);
xor U2600 (N_2600,In_489,In_267);
and U2601 (N_2601,In_989,In_2921);
nor U2602 (N_2602,In_484,In_858);
nor U2603 (N_2603,In_2017,In_183);
nor U2604 (N_2604,In_1672,In_1799);
xor U2605 (N_2605,In_1894,In_862);
xor U2606 (N_2606,In_2920,In_1003);
and U2607 (N_2607,In_2866,In_816);
nor U2608 (N_2608,In_2963,In_1254);
and U2609 (N_2609,In_433,In_2330);
nor U2610 (N_2610,In_2978,In_2062);
xor U2611 (N_2611,In_1634,In_2252);
nand U2612 (N_2612,In_410,In_2363);
xnor U2613 (N_2613,In_2011,In_2606);
nand U2614 (N_2614,In_2537,In_2902);
xor U2615 (N_2615,In_398,In_2323);
and U2616 (N_2616,In_2841,In_2550);
xnor U2617 (N_2617,In_1097,In_17);
or U2618 (N_2618,In_1546,In_1179);
xor U2619 (N_2619,In_850,In_176);
nand U2620 (N_2620,In_623,In_2607);
xnor U2621 (N_2621,In_2867,In_871);
nor U2622 (N_2622,In_1360,In_584);
nor U2623 (N_2623,In_438,In_24);
nand U2624 (N_2624,In_166,In_179);
or U2625 (N_2625,In_1149,In_1046);
xnor U2626 (N_2626,In_1009,In_326);
nor U2627 (N_2627,In_2675,In_1884);
and U2628 (N_2628,In_41,In_1540);
xor U2629 (N_2629,In_2720,In_786);
and U2630 (N_2630,In_1810,In_674);
or U2631 (N_2631,In_244,In_493);
nand U2632 (N_2632,In_1542,In_1865);
nor U2633 (N_2633,In_2590,In_300);
or U2634 (N_2634,In_1236,In_680);
or U2635 (N_2635,In_751,In_2448);
and U2636 (N_2636,In_2464,In_842);
nor U2637 (N_2637,In_2635,In_1911);
xor U2638 (N_2638,In_1916,In_879);
nor U2639 (N_2639,In_859,In_1417);
xnor U2640 (N_2640,In_811,In_1012);
nor U2641 (N_2641,In_1629,In_2355);
nand U2642 (N_2642,In_142,In_1324);
xnor U2643 (N_2643,In_711,In_2822);
and U2644 (N_2644,In_2963,In_588);
xor U2645 (N_2645,In_767,In_570);
nor U2646 (N_2646,In_2887,In_2312);
nor U2647 (N_2647,In_971,In_2521);
xor U2648 (N_2648,In_1735,In_1473);
xnor U2649 (N_2649,In_2562,In_676);
nand U2650 (N_2650,In_2028,In_2864);
or U2651 (N_2651,In_2539,In_308);
nor U2652 (N_2652,In_668,In_2902);
and U2653 (N_2653,In_2018,In_1874);
or U2654 (N_2654,In_2754,In_2372);
xnor U2655 (N_2655,In_1289,In_865);
nand U2656 (N_2656,In_930,In_1896);
or U2657 (N_2657,In_1020,In_674);
nor U2658 (N_2658,In_2298,In_2827);
and U2659 (N_2659,In_2764,In_901);
xnor U2660 (N_2660,In_1354,In_1426);
and U2661 (N_2661,In_1334,In_371);
nor U2662 (N_2662,In_566,In_2026);
xor U2663 (N_2663,In_2895,In_1511);
xor U2664 (N_2664,In_1284,In_871);
nand U2665 (N_2665,In_2034,In_2569);
nor U2666 (N_2666,In_541,In_606);
xnor U2667 (N_2667,In_2997,In_1315);
xor U2668 (N_2668,In_283,In_1194);
nor U2669 (N_2669,In_870,In_994);
nor U2670 (N_2670,In_139,In_722);
nor U2671 (N_2671,In_149,In_1195);
and U2672 (N_2672,In_1087,In_761);
nand U2673 (N_2673,In_990,In_2611);
xor U2674 (N_2674,In_2376,In_2830);
and U2675 (N_2675,In_717,In_2890);
xnor U2676 (N_2676,In_93,In_2132);
and U2677 (N_2677,In_242,In_1684);
and U2678 (N_2678,In_1512,In_803);
nor U2679 (N_2679,In_181,In_1539);
xnor U2680 (N_2680,In_386,In_2500);
and U2681 (N_2681,In_1082,In_552);
nor U2682 (N_2682,In_2911,In_317);
and U2683 (N_2683,In_1811,In_1224);
and U2684 (N_2684,In_798,In_1942);
nand U2685 (N_2685,In_826,In_1163);
and U2686 (N_2686,In_720,In_318);
and U2687 (N_2687,In_616,In_1024);
nor U2688 (N_2688,In_315,In_2694);
and U2689 (N_2689,In_1536,In_304);
or U2690 (N_2690,In_419,In_2323);
or U2691 (N_2691,In_1161,In_1771);
and U2692 (N_2692,In_2160,In_1153);
nand U2693 (N_2693,In_1957,In_248);
and U2694 (N_2694,In_372,In_583);
nor U2695 (N_2695,In_1825,In_525);
nand U2696 (N_2696,In_105,In_388);
nand U2697 (N_2697,In_574,In_2189);
nor U2698 (N_2698,In_2967,In_1503);
nand U2699 (N_2699,In_496,In_1524);
or U2700 (N_2700,In_986,In_938);
and U2701 (N_2701,In_863,In_2235);
xnor U2702 (N_2702,In_1527,In_1421);
xor U2703 (N_2703,In_1858,In_379);
nand U2704 (N_2704,In_2193,In_2862);
nor U2705 (N_2705,In_895,In_1645);
xnor U2706 (N_2706,In_49,In_477);
or U2707 (N_2707,In_1898,In_1097);
or U2708 (N_2708,In_1212,In_1997);
xnor U2709 (N_2709,In_387,In_1563);
xor U2710 (N_2710,In_1335,In_2739);
and U2711 (N_2711,In_273,In_2163);
xnor U2712 (N_2712,In_1578,In_905);
nor U2713 (N_2713,In_558,In_1093);
and U2714 (N_2714,In_2068,In_1079);
nand U2715 (N_2715,In_1985,In_1654);
xnor U2716 (N_2716,In_2329,In_1259);
nor U2717 (N_2717,In_617,In_2226);
xor U2718 (N_2718,In_2184,In_261);
or U2719 (N_2719,In_1849,In_2615);
or U2720 (N_2720,In_1755,In_487);
or U2721 (N_2721,In_1694,In_442);
or U2722 (N_2722,In_2024,In_1740);
nor U2723 (N_2723,In_173,In_1688);
or U2724 (N_2724,In_1334,In_1413);
nor U2725 (N_2725,In_1816,In_426);
nor U2726 (N_2726,In_1851,In_1782);
nor U2727 (N_2727,In_424,In_2888);
xnor U2728 (N_2728,In_53,In_899);
or U2729 (N_2729,In_55,In_2763);
xor U2730 (N_2730,In_1213,In_1052);
nor U2731 (N_2731,In_2537,In_642);
xor U2732 (N_2732,In_1597,In_2722);
nor U2733 (N_2733,In_1844,In_2101);
nor U2734 (N_2734,In_1620,In_2416);
or U2735 (N_2735,In_2017,In_1522);
and U2736 (N_2736,In_937,In_1892);
xor U2737 (N_2737,In_1581,In_969);
or U2738 (N_2738,In_688,In_467);
or U2739 (N_2739,In_1095,In_1923);
or U2740 (N_2740,In_2652,In_2589);
and U2741 (N_2741,In_1693,In_2109);
nand U2742 (N_2742,In_1216,In_944);
and U2743 (N_2743,In_1828,In_208);
nand U2744 (N_2744,In_1515,In_2513);
xnor U2745 (N_2745,In_1489,In_1732);
and U2746 (N_2746,In_1572,In_1159);
and U2747 (N_2747,In_179,In_594);
or U2748 (N_2748,In_816,In_2274);
and U2749 (N_2749,In_1665,In_1225);
or U2750 (N_2750,In_410,In_2826);
and U2751 (N_2751,In_2276,In_2513);
nor U2752 (N_2752,In_1715,In_2399);
and U2753 (N_2753,In_2068,In_1077);
and U2754 (N_2754,In_994,In_2033);
or U2755 (N_2755,In_1014,In_2826);
and U2756 (N_2756,In_2514,In_2901);
xor U2757 (N_2757,In_2373,In_803);
nand U2758 (N_2758,In_1681,In_1203);
and U2759 (N_2759,In_1145,In_826);
xor U2760 (N_2760,In_291,In_1630);
nand U2761 (N_2761,In_1329,In_1835);
or U2762 (N_2762,In_1283,In_1756);
or U2763 (N_2763,In_1362,In_81);
or U2764 (N_2764,In_1445,In_1638);
nor U2765 (N_2765,In_864,In_1486);
and U2766 (N_2766,In_1184,In_2761);
nand U2767 (N_2767,In_1854,In_2624);
xnor U2768 (N_2768,In_75,In_1851);
or U2769 (N_2769,In_1254,In_963);
and U2770 (N_2770,In_1154,In_2102);
and U2771 (N_2771,In_2022,In_1481);
nand U2772 (N_2772,In_607,In_1416);
and U2773 (N_2773,In_1669,In_2206);
nand U2774 (N_2774,In_2073,In_2425);
nor U2775 (N_2775,In_210,In_2730);
and U2776 (N_2776,In_116,In_1197);
xnor U2777 (N_2777,In_2958,In_1463);
and U2778 (N_2778,In_1586,In_2387);
xnor U2779 (N_2779,In_1203,In_1917);
xor U2780 (N_2780,In_697,In_2519);
nand U2781 (N_2781,In_2565,In_628);
or U2782 (N_2782,In_1223,In_1593);
nand U2783 (N_2783,In_2693,In_218);
nor U2784 (N_2784,In_1203,In_1639);
and U2785 (N_2785,In_1447,In_2105);
nand U2786 (N_2786,In_2133,In_1859);
and U2787 (N_2787,In_1948,In_1103);
nor U2788 (N_2788,In_2268,In_2843);
or U2789 (N_2789,In_1810,In_629);
and U2790 (N_2790,In_486,In_2276);
nor U2791 (N_2791,In_1248,In_217);
and U2792 (N_2792,In_221,In_118);
nand U2793 (N_2793,In_895,In_2782);
nor U2794 (N_2794,In_2734,In_1472);
nand U2795 (N_2795,In_2349,In_658);
nor U2796 (N_2796,In_521,In_1978);
nand U2797 (N_2797,In_1921,In_1094);
nor U2798 (N_2798,In_1863,In_1209);
nor U2799 (N_2799,In_2517,In_1241);
or U2800 (N_2800,In_2312,In_18);
xnor U2801 (N_2801,In_118,In_680);
and U2802 (N_2802,In_966,In_866);
nand U2803 (N_2803,In_1341,In_2551);
and U2804 (N_2804,In_933,In_2400);
or U2805 (N_2805,In_1512,In_227);
or U2806 (N_2806,In_2806,In_141);
nor U2807 (N_2807,In_190,In_104);
or U2808 (N_2808,In_2251,In_1641);
and U2809 (N_2809,In_1429,In_68);
or U2810 (N_2810,In_2671,In_746);
or U2811 (N_2811,In_435,In_2841);
or U2812 (N_2812,In_158,In_198);
or U2813 (N_2813,In_2121,In_1871);
xor U2814 (N_2814,In_2178,In_725);
or U2815 (N_2815,In_1055,In_117);
or U2816 (N_2816,In_1189,In_456);
nand U2817 (N_2817,In_231,In_1712);
and U2818 (N_2818,In_2967,In_2808);
nor U2819 (N_2819,In_2331,In_2430);
and U2820 (N_2820,In_2966,In_1870);
nor U2821 (N_2821,In_606,In_2288);
or U2822 (N_2822,In_1403,In_2674);
and U2823 (N_2823,In_711,In_2918);
xnor U2824 (N_2824,In_1738,In_1747);
nor U2825 (N_2825,In_1733,In_2087);
or U2826 (N_2826,In_1901,In_1600);
and U2827 (N_2827,In_1807,In_1640);
xor U2828 (N_2828,In_2558,In_2574);
nor U2829 (N_2829,In_2119,In_2840);
nand U2830 (N_2830,In_593,In_518);
nor U2831 (N_2831,In_2406,In_1728);
nor U2832 (N_2832,In_392,In_2556);
and U2833 (N_2833,In_1179,In_482);
or U2834 (N_2834,In_1486,In_1698);
xnor U2835 (N_2835,In_1879,In_286);
xor U2836 (N_2836,In_62,In_897);
or U2837 (N_2837,In_1024,In_660);
and U2838 (N_2838,In_594,In_940);
nor U2839 (N_2839,In_419,In_153);
nand U2840 (N_2840,In_926,In_2779);
and U2841 (N_2841,In_147,In_90);
and U2842 (N_2842,In_2207,In_2047);
xnor U2843 (N_2843,In_1897,In_1755);
or U2844 (N_2844,In_430,In_2668);
nor U2845 (N_2845,In_2330,In_1695);
nor U2846 (N_2846,In_44,In_94);
or U2847 (N_2847,In_1164,In_1627);
xor U2848 (N_2848,In_1408,In_562);
nand U2849 (N_2849,In_344,In_2009);
nor U2850 (N_2850,In_2802,In_1332);
nor U2851 (N_2851,In_2073,In_623);
nor U2852 (N_2852,In_54,In_885);
xor U2853 (N_2853,In_330,In_688);
xor U2854 (N_2854,In_991,In_2918);
nor U2855 (N_2855,In_1302,In_1162);
xor U2856 (N_2856,In_2746,In_1200);
nand U2857 (N_2857,In_885,In_2699);
nand U2858 (N_2858,In_2236,In_651);
xnor U2859 (N_2859,In_2256,In_1649);
and U2860 (N_2860,In_1757,In_2750);
and U2861 (N_2861,In_1653,In_748);
nand U2862 (N_2862,In_1375,In_1121);
nand U2863 (N_2863,In_892,In_1429);
nor U2864 (N_2864,In_457,In_1607);
nand U2865 (N_2865,In_2526,In_303);
or U2866 (N_2866,In_1147,In_90);
xnor U2867 (N_2867,In_726,In_1807);
and U2868 (N_2868,In_1401,In_1902);
nor U2869 (N_2869,In_1174,In_254);
nand U2870 (N_2870,In_809,In_2021);
and U2871 (N_2871,In_1600,In_1257);
nor U2872 (N_2872,In_2837,In_1980);
nor U2873 (N_2873,In_1001,In_723);
nand U2874 (N_2874,In_2273,In_1198);
and U2875 (N_2875,In_2019,In_1043);
and U2876 (N_2876,In_1673,In_989);
xnor U2877 (N_2877,In_2240,In_2065);
xnor U2878 (N_2878,In_549,In_815);
and U2879 (N_2879,In_61,In_834);
and U2880 (N_2880,In_33,In_197);
nor U2881 (N_2881,In_1804,In_2189);
or U2882 (N_2882,In_1253,In_2432);
nor U2883 (N_2883,In_2957,In_9);
nor U2884 (N_2884,In_2491,In_2742);
nand U2885 (N_2885,In_2845,In_1450);
and U2886 (N_2886,In_1313,In_929);
xnor U2887 (N_2887,In_757,In_1716);
nor U2888 (N_2888,In_1717,In_2024);
and U2889 (N_2889,In_2165,In_2605);
xor U2890 (N_2890,In_1804,In_821);
or U2891 (N_2891,In_2075,In_1775);
nor U2892 (N_2892,In_1135,In_1938);
xor U2893 (N_2893,In_1768,In_2952);
nand U2894 (N_2894,In_2042,In_2073);
xor U2895 (N_2895,In_1138,In_2813);
and U2896 (N_2896,In_2690,In_888);
or U2897 (N_2897,In_676,In_1293);
and U2898 (N_2898,In_1667,In_1378);
and U2899 (N_2899,In_1122,In_2162);
and U2900 (N_2900,In_1296,In_1788);
xor U2901 (N_2901,In_858,In_2761);
nand U2902 (N_2902,In_2721,In_1264);
or U2903 (N_2903,In_444,In_69);
nand U2904 (N_2904,In_995,In_203);
nand U2905 (N_2905,In_554,In_1097);
xnor U2906 (N_2906,In_2101,In_2703);
or U2907 (N_2907,In_614,In_2081);
xor U2908 (N_2908,In_597,In_2488);
or U2909 (N_2909,In_753,In_1476);
xnor U2910 (N_2910,In_724,In_426);
or U2911 (N_2911,In_2847,In_2897);
and U2912 (N_2912,In_2319,In_2252);
nand U2913 (N_2913,In_157,In_1060);
and U2914 (N_2914,In_1531,In_865);
and U2915 (N_2915,In_1782,In_2722);
or U2916 (N_2916,In_14,In_810);
or U2917 (N_2917,In_1422,In_1345);
and U2918 (N_2918,In_452,In_210);
nand U2919 (N_2919,In_2682,In_2495);
nor U2920 (N_2920,In_1946,In_1751);
nand U2921 (N_2921,In_1286,In_2763);
nor U2922 (N_2922,In_2562,In_510);
nor U2923 (N_2923,In_2563,In_308);
and U2924 (N_2924,In_1371,In_1336);
and U2925 (N_2925,In_587,In_2100);
nand U2926 (N_2926,In_213,In_2117);
nand U2927 (N_2927,In_2788,In_1105);
nor U2928 (N_2928,In_695,In_740);
nand U2929 (N_2929,In_2375,In_646);
or U2930 (N_2930,In_1922,In_297);
or U2931 (N_2931,In_1791,In_2555);
or U2932 (N_2932,In_427,In_552);
nand U2933 (N_2933,In_1169,In_2776);
or U2934 (N_2934,In_1350,In_1424);
or U2935 (N_2935,In_2381,In_2555);
and U2936 (N_2936,In_1187,In_2646);
nand U2937 (N_2937,In_798,In_2881);
and U2938 (N_2938,In_296,In_715);
nor U2939 (N_2939,In_668,In_2829);
or U2940 (N_2940,In_1248,In_2447);
nor U2941 (N_2941,In_1867,In_650);
xnor U2942 (N_2942,In_2307,In_2688);
nand U2943 (N_2943,In_1509,In_1457);
and U2944 (N_2944,In_2811,In_1428);
or U2945 (N_2945,In_121,In_1095);
nand U2946 (N_2946,In_1349,In_1159);
nand U2947 (N_2947,In_2603,In_1839);
or U2948 (N_2948,In_1880,In_1027);
nor U2949 (N_2949,In_1291,In_998);
or U2950 (N_2950,In_557,In_1926);
or U2951 (N_2951,In_2514,In_127);
xor U2952 (N_2952,In_2510,In_2525);
or U2953 (N_2953,In_1509,In_2204);
and U2954 (N_2954,In_1413,In_1481);
nand U2955 (N_2955,In_2552,In_2283);
xor U2956 (N_2956,In_1855,In_2611);
nand U2957 (N_2957,In_244,In_2512);
nor U2958 (N_2958,In_2223,In_229);
or U2959 (N_2959,In_2332,In_1195);
xor U2960 (N_2960,In_900,In_442);
or U2961 (N_2961,In_869,In_2002);
nor U2962 (N_2962,In_1546,In_1020);
and U2963 (N_2963,In_382,In_2610);
nor U2964 (N_2964,In_1611,In_1910);
or U2965 (N_2965,In_2981,In_1987);
nor U2966 (N_2966,In_922,In_2197);
and U2967 (N_2967,In_1345,In_122);
and U2968 (N_2968,In_489,In_288);
or U2969 (N_2969,In_826,In_254);
or U2970 (N_2970,In_1568,In_109);
or U2971 (N_2971,In_752,In_1463);
xnor U2972 (N_2972,In_1669,In_881);
nand U2973 (N_2973,In_843,In_2342);
and U2974 (N_2974,In_2361,In_1573);
and U2975 (N_2975,In_1180,In_1486);
nor U2976 (N_2976,In_595,In_631);
and U2977 (N_2977,In_2738,In_1283);
or U2978 (N_2978,In_2773,In_2298);
and U2979 (N_2979,In_1469,In_1430);
or U2980 (N_2980,In_2881,In_1946);
xnor U2981 (N_2981,In_605,In_2532);
nor U2982 (N_2982,In_915,In_1184);
nand U2983 (N_2983,In_1137,In_1686);
and U2984 (N_2984,In_701,In_1095);
nand U2985 (N_2985,In_681,In_395);
nand U2986 (N_2986,In_2697,In_1870);
nor U2987 (N_2987,In_1881,In_376);
or U2988 (N_2988,In_780,In_2103);
nand U2989 (N_2989,In_1058,In_357);
and U2990 (N_2990,In_981,In_1405);
nor U2991 (N_2991,In_1974,In_53);
or U2992 (N_2992,In_689,In_2401);
and U2993 (N_2993,In_129,In_2543);
nor U2994 (N_2994,In_1615,In_568);
nor U2995 (N_2995,In_2252,In_1481);
and U2996 (N_2996,In_2429,In_1206);
nand U2997 (N_2997,In_2297,In_235);
and U2998 (N_2998,In_1000,In_2244);
and U2999 (N_2999,In_364,In_563);
nor U3000 (N_3000,In_328,In_2708);
and U3001 (N_3001,In_362,In_481);
or U3002 (N_3002,In_2922,In_546);
nand U3003 (N_3003,In_833,In_441);
and U3004 (N_3004,In_1198,In_1222);
or U3005 (N_3005,In_2413,In_2607);
and U3006 (N_3006,In_1079,In_1760);
xor U3007 (N_3007,In_1237,In_800);
and U3008 (N_3008,In_2446,In_1738);
or U3009 (N_3009,In_622,In_46);
xnor U3010 (N_3010,In_1088,In_1117);
and U3011 (N_3011,In_1587,In_745);
or U3012 (N_3012,In_1372,In_2846);
xor U3013 (N_3013,In_2755,In_1093);
or U3014 (N_3014,In_2583,In_1524);
xor U3015 (N_3015,In_902,In_2182);
or U3016 (N_3016,In_1687,In_1806);
xnor U3017 (N_3017,In_859,In_1031);
nor U3018 (N_3018,In_552,In_1639);
and U3019 (N_3019,In_459,In_1867);
and U3020 (N_3020,In_561,In_1710);
and U3021 (N_3021,In_2229,In_1887);
nand U3022 (N_3022,In_993,In_1084);
and U3023 (N_3023,In_41,In_406);
nand U3024 (N_3024,In_1270,In_1313);
nor U3025 (N_3025,In_1482,In_477);
nor U3026 (N_3026,In_1826,In_428);
xor U3027 (N_3027,In_500,In_508);
xor U3028 (N_3028,In_1262,In_846);
xor U3029 (N_3029,In_2556,In_2270);
xor U3030 (N_3030,In_166,In_2964);
nor U3031 (N_3031,In_671,In_1218);
or U3032 (N_3032,In_1934,In_2507);
nand U3033 (N_3033,In_631,In_2986);
xnor U3034 (N_3034,In_2531,In_1837);
xnor U3035 (N_3035,In_1891,In_1317);
nand U3036 (N_3036,In_1583,In_1726);
nand U3037 (N_3037,In_1479,In_2926);
or U3038 (N_3038,In_2417,In_2901);
xnor U3039 (N_3039,In_984,In_2311);
or U3040 (N_3040,In_2783,In_2821);
nand U3041 (N_3041,In_1587,In_23);
nor U3042 (N_3042,In_1997,In_1720);
nand U3043 (N_3043,In_1490,In_608);
nor U3044 (N_3044,In_2609,In_1789);
nand U3045 (N_3045,In_1275,In_812);
and U3046 (N_3046,In_2403,In_589);
nor U3047 (N_3047,In_888,In_2039);
and U3048 (N_3048,In_710,In_2611);
and U3049 (N_3049,In_2337,In_278);
nand U3050 (N_3050,In_500,In_2944);
nor U3051 (N_3051,In_964,In_2198);
nand U3052 (N_3052,In_1329,In_177);
nor U3053 (N_3053,In_901,In_277);
and U3054 (N_3054,In_494,In_945);
and U3055 (N_3055,In_1692,In_414);
xor U3056 (N_3056,In_568,In_637);
xnor U3057 (N_3057,In_440,In_2877);
and U3058 (N_3058,In_2190,In_196);
and U3059 (N_3059,In_2944,In_1253);
nand U3060 (N_3060,In_2668,In_1382);
nand U3061 (N_3061,In_2488,In_478);
or U3062 (N_3062,In_206,In_1307);
and U3063 (N_3063,In_154,In_86);
nor U3064 (N_3064,In_2530,In_2802);
nor U3065 (N_3065,In_2854,In_2106);
nor U3066 (N_3066,In_2878,In_224);
or U3067 (N_3067,In_1210,In_721);
nand U3068 (N_3068,In_2788,In_1159);
xnor U3069 (N_3069,In_1712,In_1113);
or U3070 (N_3070,In_1407,In_1674);
or U3071 (N_3071,In_2655,In_1789);
xnor U3072 (N_3072,In_1844,In_116);
and U3073 (N_3073,In_2743,In_2322);
xnor U3074 (N_3074,In_94,In_337);
nor U3075 (N_3075,In_2300,In_2929);
or U3076 (N_3076,In_2280,In_1957);
or U3077 (N_3077,In_2209,In_1886);
and U3078 (N_3078,In_1713,In_1590);
nor U3079 (N_3079,In_2839,In_102);
xnor U3080 (N_3080,In_994,In_880);
nand U3081 (N_3081,In_2166,In_1240);
nor U3082 (N_3082,In_752,In_350);
nand U3083 (N_3083,In_398,In_1448);
or U3084 (N_3084,In_2380,In_49);
nor U3085 (N_3085,In_288,In_2195);
nor U3086 (N_3086,In_1718,In_2658);
and U3087 (N_3087,In_2972,In_802);
nor U3088 (N_3088,In_1931,In_197);
or U3089 (N_3089,In_1243,In_1437);
or U3090 (N_3090,In_2609,In_371);
nand U3091 (N_3091,In_857,In_2404);
nor U3092 (N_3092,In_1514,In_2051);
and U3093 (N_3093,In_2156,In_335);
nor U3094 (N_3094,In_1838,In_2440);
xor U3095 (N_3095,In_804,In_870);
or U3096 (N_3096,In_222,In_2912);
nor U3097 (N_3097,In_1407,In_1254);
nand U3098 (N_3098,In_1772,In_393);
nand U3099 (N_3099,In_2698,In_1892);
nand U3100 (N_3100,In_1282,In_896);
or U3101 (N_3101,In_2312,In_682);
nor U3102 (N_3102,In_724,In_392);
or U3103 (N_3103,In_1277,In_59);
and U3104 (N_3104,In_1174,In_1291);
xnor U3105 (N_3105,In_452,In_630);
xor U3106 (N_3106,In_1323,In_1758);
xnor U3107 (N_3107,In_1132,In_757);
nor U3108 (N_3108,In_62,In_2821);
and U3109 (N_3109,In_1862,In_615);
or U3110 (N_3110,In_2406,In_821);
nor U3111 (N_3111,In_2259,In_589);
and U3112 (N_3112,In_1282,In_179);
or U3113 (N_3113,In_496,In_675);
nor U3114 (N_3114,In_430,In_1966);
nand U3115 (N_3115,In_258,In_2606);
and U3116 (N_3116,In_1604,In_1262);
nor U3117 (N_3117,In_2084,In_1388);
xnor U3118 (N_3118,In_743,In_500);
nor U3119 (N_3119,In_875,In_170);
nor U3120 (N_3120,In_1530,In_1259);
xnor U3121 (N_3121,In_1701,In_599);
nor U3122 (N_3122,In_2743,In_1462);
nand U3123 (N_3123,In_1393,In_80);
nand U3124 (N_3124,In_1877,In_2092);
and U3125 (N_3125,In_1439,In_902);
and U3126 (N_3126,In_1352,In_836);
or U3127 (N_3127,In_2128,In_2545);
xnor U3128 (N_3128,In_2134,In_2885);
nand U3129 (N_3129,In_1364,In_2831);
or U3130 (N_3130,In_1373,In_2721);
or U3131 (N_3131,In_2854,In_828);
nor U3132 (N_3132,In_1379,In_2803);
nand U3133 (N_3133,In_2375,In_1115);
and U3134 (N_3134,In_1010,In_1774);
xnor U3135 (N_3135,In_2330,In_898);
or U3136 (N_3136,In_688,In_618);
nand U3137 (N_3137,In_2270,In_1826);
and U3138 (N_3138,In_1203,In_255);
nor U3139 (N_3139,In_1749,In_2637);
or U3140 (N_3140,In_2327,In_894);
or U3141 (N_3141,In_1947,In_797);
and U3142 (N_3142,In_1878,In_1615);
and U3143 (N_3143,In_710,In_2108);
nor U3144 (N_3144,In_1473,In_606);
nand U3145 (N_3145,In_829,In_1754);
nor U3146 (N_3146,In_216,In_1534);
xnor U3147 (N_3147,In_2955,In_744);
nor U3148 (N_3148,In_1479,In_2847);
and U3149 (N_3149,In_88,In_875);
nand U3150 (N_3150,In_1770,In_1217);
xor U3151 (N_3151,In_2180,In_2321);
nor U3152 (N_3152,In_2674,In_1888);
and U3153 (N_3153,In_18,In_29);
xnor U3154 (N_3154,In_2571,In_1993);
and U3155 (N_3155,In_1723,In_2885);
xor U3156 (N_3156,In_2405,In_1857);
or U3157 (N_3157,In_1883,In_834);
nand U3158 (N_3158,In_1120,In_2186);
and U3159 (N_3159,In_1621,In_220);
nor U3160 (N_3160,In_1330,In_1436);
xnor U3161 (N_3161,In_1622,In_1959);
nor U3162 (N_3162,In_2680,In_2757);
nand U3163 (N_3163,In_463,In_2943);
and U3164 (N_3164,In_2774,In_2374);
xor U3165 (N_3165,In_135,In_2877);
or U3166 (N_3166,In_527,In_1890);
or U3167 (N_3167,In_1212,In_990);
xnor U3168 (N_3168,In_2302,In_2740);
and U3169 (N_3169,In_1894,In_2171);
xor U3170 (N_3170,In_2357,In_2401);
nand U3171 (N_3171,In_616,In_240);
nor U3172 (N_3172,In_2,In_2658);
and U3173 (N_3173,In_1214,In_1152);
xnor U3174 (N_3174,In_1818,In_1026);
or U3175 (N_3175,In_985,In_435);
or U3176 (N_3176,In_308,In_2282);
xnor U3177 (N_3177,In_1364,In_1283);
xor U3178 (N_3178,In_1290,In_2070);
xor U3179 (N_3179,In_1848,In_1403);
nor U3180 (N_3180,In_1066,In_1614);
and U3181 (N_3181,In_76,In_401);
or U3182 (N_3182,In_2408,In_2660);
nand U3183 (N_3183,In_2776,In_837);
or U3184 (N_3184,In_1166,In_1008);
nor U3185 (N_3185,In_434,In_2214);
and U3186 (N_3186,In_2144,In_1106);
and U3187 (N_3187,In_2760,In_2274);
and U3188 (N_3188,In_221,In_1926);
nand U3189 (N_3189,In_368,In_106);
nor U3190 (N_3190,In_299,In_375);
nor U3191 (N_3191,In_2621,In_1884);
xor U3192 (N_3192,In_77,In_1739);
nand U3193 (N_3193,In_1106,In_1774);
nand U3194 (N_3194,In_542,In_730);
nor U3195 (N_3195,In_2940,In_2579);
nand U3196 (N_3196,In_991,In_2703);
nor U3197 (N_3197,In_1271,In_87);
and U3198 (N_3198,In_742,In_1523);
xor U3199 (N_3199,In_1102,In_2272);
nor U3200 (N_3200,In_2701,In_1533);
nand U3201 (N_3201,In_2730,In_576);
nor U3202 (N_3202,In_2904,In_801);
and U3203 (N_3203,In_2478,In_2843);
nor U3204 (N_3204,In_948,In_59);
and U3205 (N_3205,In_1328,In_1915);
nor U3206 (N_3206,In_2322,In_1243);
nor U3207 (N_3207,In_100,In_839);
nand U3208 (N_3208,In_1223,In_1059);
or U3209 (N_3209,In_2275,In_2082);
xor U3210 (N_3210,In_2616,In_730);
and U3211 (N_3211,In_161,In_2649);
or U3212 (N_3212,In_363,In_593);
and U3213 (N_3213,In_18,In_1052);
xor U3214 (N_3214,In_1060,In_2728);
and U3215 (N_3215,In_773,In_1676);
and U3216 (N_3216,In_1006,In_2036);
and U3217 (N_3217,In_641,In_484);
and U3218 (N_3218,In_1972,In_1211);
nor U3219 (N_3219,In_1493,In_784);
and U3220 (N_3220,In_2715,In_1040);
nand U3221 (N_3221,In_2459,In_1842);
nor U3222 (N_3222,In_1311,In_2187);
nor U3223 (N_3223,In_2461,In_1686);
nand U3224 (N_3224,In_2141,In_1869);
nand U3225 (N_3225,In_1624,In_1378);
nor U3226 (N_3226,In_132,In_1542);
or U3227 (N_3227,In_1937,In_38);
xnor U3228 (N_3228,In_2833,In_916);
or U3229 (N_3229,In_2326,In_817);
nor U3230 (N_3230,In_1214,In_2869);
nor U3231 (N_3231,In_1706,In_929);
nor U3232 (N_3232,In_2643,In_2087);
nand U3233 (N_3233,In_1798,In_2742);
nand U3234 (N_3234,In_1440,In_2179);
and U3235 (N_3235,In_1606,In_2544);
nor U3236 (N_3236,In_2926,In_2562);
nand U3237 (N_3237,In_106,In_2007);
nor U3238 (N_3238,In_456,In_1625);
or U3239 (N_3239,In_2622,In_1130);
and U3240 (N_3240,In_843,In_8);
xor U3241 (N_3241,In_2466,In_2790);
nand U3242 (N_3242,In_834,In_1169);
or U3243 (N_3243,In_861,In_1454);
nand U3244 (N_3244,In_2094,In_1622);
nor U3245 (N_3245,In_2632,In_2743);
xor U3246 (N_3246,In_1491,In_192);
nor U3247 (N_3247,In_1538,In_2968);
or U3248 (N_3248,In_117,In_1944);
and U3249 (N_3249,In_1037,In_1770);
xnor U3250 (N_3250,In_430,In_2486);
nor U3251 (N_3251,In_507,In_379);
nand U3252 (N_3252,In_2850,In_233);
nand U3253 (N_3253,In_2015,In_1602);
nand U3254 (N_3254,In_2626,In_1231);
nor U3255 (N_3255,In_2033,In_673);
or U3256 (N_3256,In_1277,In_1789);
or U3257 (N_3257,In_1375,In_1891);
nand U3258 (N_3258,In_702,In_2300);
nand U3259 (N_3259,In_846,In_255);
nand U3260 (N_3260,In_1987,In_2923);
or U3261 (N_3261,In_2322,In_1685);
nand U3262 (N_3262,In_1574,In_1369);
xnor U3263 (N_3263,In_2202,In_2376);
and U3264 (N_3264,In_1522,In_2064);
xnor U3265 (N_3265,In_1390,In_282);
and U3266 (N_3266,In_2227,In_2273);
and U3267 (N_3267,In_2976,In_1556);
and U3268 (N_3268,In_1350,In_2955);
xnor U3269 (N_3269,In_545,In_2074);
or U3270 (N_3270,In_90,In_80);
or U3271 (N_3271,In_847,In_552);
nor U3272 (N_3272,In_1790,In_821);
nor U3273 (N_3273,In_916,In_320);
and U3274 (N_3274,In_38,In_2960);
nor U3275 (N_3275,In_1392,In_2611);
nand U3276 (N_3276,In_2261,In_1752);
and U3277 (N_3277,In_1554,In_991);
nand U3278 (N_3278,In_96,In_2806);
or U3279 (N_3279,In_2631,In_2678);
or U3280 (N_3280,In_675,In_1115);
and U3281 (N_3281,In_2369,In_1302);
and U3282 (N_3282,In_480,In_1672);
nand U3283 (N_3283,In_62,In_2641);
and U3284 (N_3284,In_2061,In_2953);
xnor U3285 (N_3285,In_1625,In_2543);
xor U3286 (N_3286,In_2590,In_850);
xnor U3287 (N_3287,In_2052,In_1640);
xor U3288 (N_3288,In_145,In_2303);
xnor U3289 (N_3289,In_1661,In_1885);
and U3290 (N_3290,In_533,In_1101);
xnor U3291 (N_3291,In_1880,In_935);
nand U3292 (N_3292,In_604,In_2796);
nand U3293 (N_3293,In_1258,In_2463);
and U3294 (N_3294,In_1592,In_1596);
nand U3295 (N_3295,In_991,In_51);
nor U3296 (N_3296,In_1636,In_1573);
xnor U3297 (N_3297,In_2228,In_901);
nand U3298 (N_3298,In_706,In_553);
nor U3299 (N_3299,In_2718,In_53);
xnor U3300 (N_3300,In_2315,In_136);
and U3301 (N_3301,In_1958,In_1187);
or U3302 (N_3302,In_2568,In_1445);
or U3303 (N_3303,In_13,In_570);
or U3304 (N_3304,In_1247,In_887);
or U3305 (N_3305,In_1152,In_268);
nand U3306 (N_3306,In_2008,In_1212);
xor U3307 (N_3307,In_94,In_561);
and U3308 (N_3308,In_2802,In_2219);
nand U3309 (N_3309,In_2456,In_1705);
xor U3310 (N_3310,In_763,In_2947);
nor U3311 (N_3311,In_158,In_593);
or U3312 (N_3312,In_1310,In_747);
nor U3313 (N_3313,In_1440,In_1935);
and U3314 (N_3314,In_1833,In_2712);
and U3315 (N_3315,In_1717,In_2354);
and U3316 (N_3316,In_2478,In_2012);
nor U3317 (N_3317,In_2430,In_1533);
nor U3318 (N_3318,In_1488,In_463);
nor U3319 (N_3319,In_1406,In_2112);
nor U3320 (N_3320,In_1916,In_1946);
or U3321 (N_3321,In_1745,In_1848);
and U3322 (N_3322,In_2113,In_1953);
nor U3323 (N_3323,In_130,In_2836);
xor U3324 (N_3324,In_2530,In_1102);
xnor U3325 (N_3325,In_2623,In_568);
nand U3326 (N_3326,In_616,In_1236);
nor U3327 (N_3327,In_1987,In_1386);
xor U3328 (N_3328,In_2865,In_708);
or U3329 (N_3329,In_497,In_2871);
xor U3330 (N_3330,In_2024,In_656);
nand U3331 (N_3331,In_1930,In_1024);
xor U3332 (N_3332,In_474,In_313);
nand U3333 (N_3333,In_702,In_587);
nand U3334 (N_3334,In_2025,In_2637);
nand U3335 (N_3335,In_901,In_1638);
xor U3336 (N_3336,In_548,In_2348);
nor U3337 (N_3337,In_639,In_607);
and U3338 (N_3338,In_2256,In_317);
nand U3339 (N_3339,In_168,In_2793);
and U3340 (N_3340,In_2890,In_2924);
and U3341 (N_3341,In_2551,In_1240);
xnor U3342 (N_3342,In_777,In_2301);
xor U3343 (N_3343,In_713,In_815);
or U3344 (N_3344,In_1622,In_89);
nand U3345 (N_3345,In_1870,In_342);
or U3346 (N_3346,In_1399,In_1662);
and U3347 (N_3347,In_2260,In_2211);
and U3348 (N_3348,In_1622,In_2511);
or U3349 (N_3349,In_1851,In_1375);
nor U3350 (N_3350,In_1342,In_1433);
and U3351 (N_3351,In_1440,In_370);
and U3352 (N_3352,In_2360,In_609);
xor U3353 (N_3353,In_1101,In_1611);
nor U3354 (N_3354,In_1415,In_36);
or U3355 (N_3355,In_501,In_2955);
nand U3356 (N_3356,In_373,In_1795);
nor U3357 (N_3357,In_2663,In_89);
xnor U3358 (N_3358,In_2615,In_603);
or U3359 (N_3359,In_915,In_765);
xnor U3360 (N_3360,In_1798,In_38);
or U3361 (N_3361,In_953,In_942);
nand U3362 (N_3362,In_1550,In_45);
xor U3363 (N_3363,In_1135,In_74);
and U3364 (N_3364,In_1060,In_824);
or U3365 (N_3365,In_26,In_2873);
nand U3366 (N_3366,In_2064,In_668);
nor U3367 (N_3367,In_494,In_1311);
nand U3368 (N_3368,In_510,In_2125);
xor U3369 (N_3369,In_608,In_547);
xnor U3370 (N_3370,In_2901,In_1045);
and U3371 (N_3371,In_41,In_177);
nand U3372 (N_3372,In_370,In_497);
nand U3373 (N_3373,In_2837,In_1933);
and U3374 (N_3374,In_2120,In_1600);
nand U3375 (N_3375,In_2496,In_509);
xor U3376 (N_3376,In_2456,In_2100);
nand U3377 (N_3377,In_2415,In_639);
nand U3378 (N_3378,In_859,In_2123);
nand U3379 (N_3379,In_2158,In_686);
and U3380 (N_3380,In_2119,In_897);
or U3381 (N_3381,In_2446,In_24);
xor U3382 (N_3382,In_1666,In_1994);
xor U3383 (N_3383,In_2393,In_1379);
xor U3384 (N_3384,In_1217,In_860);
xnor U3385 (N_3385,In_1961,In_321);
nand U3386 (N_3386,In_203,In_2463);
xnor U3387 (N_3387,In_2477,In_2037);
and U3388 (N_3388,In_587,In_2890);
and U3389 (N_3389,In_1323,In_104);
nor U3390 (N_3390,In_1853,In_739);
or U3391 (N_3391,In_2562,In_2187);
xor U3392 (N_3392,In_128,In_923);
xor U3393 (N_3393,In_798,In_370);
nand U3394 (N_3394,In_2769,In_530);
nor U3395 (N_3395,In_41,In_582);
xor U3396 (N_3396,In_618,In_1263);
nand U3397 (N_3397,In_968,In_2231);
nor U3398 (N_3398,In_2162,In_309);
or U3399 (N_3399,In_2237,In_20);
nand U3400 (N_3400,In_2621,In_556);
nand U3401 (N_3401,In_930,In_1016);
nor U3402 (N_3402,In_1886,In_898);
xor U3403 (N_3403,In_1372,In_395);
nor U3404 (N_3404,In_506,In_1545);
nand U3405 (N_3405,In_1852,In_366);
xor U3406 (N_3406,In_387,In_1779);
nor U3407 (N_3407,In_1261,In_438);
and U3408 (N_3408,In_5,In_1965);
xor U3409 (N_3409,In_1356,In_1588);
and U3410 (N_3410,In_1437,In_835);
nand U3411 (N_3411,In_493,In_627);
or U3412 (N_3412,In_67,In_468);
and U3413 (N_3413,In_165,In_2233);
nor U3414 (N_3414,In_2545,In_1930);
nor U3415 (N_3415,In_814,In_338);
nor U3416 (N_3416,In_2835,In_1995);
xor U3417 (N_3417,In_1265,In_1813);
nand U3418 (N_3418,In_1518,In_1945);
nor U3419 (N_3419,In_2225,In_736);
nor U3420 (N_3420,In_2245,In_695);
nor U3421 (N_3421,In_2047,In_719);
nand U3422 (N_3422,In_1157,In_1286);
xnor U3423 (N_3423,In_1757,In_2078);
nand U3424 (N_3424,In_2920,In_1610);
nor U3425 (N_3425,In_1096,In_457);
nand U3426 (N_3426,In_1694,In_1284);
xnor U3427 (N_3427,In_2670,In_1331);
nand U3428 (N_3428,In_1808,In_270);
and U3429 (N_3429,In_2287,In_2574);
or U3430 (N_3430,In_389,In_947);
and U3431 (N_3431,In_1282,In_777);
nor U3432 (N_3432,In_1069,In_855);
nand U3433 (N_3433,In_1352,In_1832);
nor U3434 (N_3434,In_1513,In_1216);
nand U3435 (N_3435,In_226,In_961);
nand U3436 (N_3436,In_158,In_1640);
xnor U3437 (N_3437,In_2497,In_2397);
xor U3438 (N_3438,In_2483,In_1624);
and U3439 (N_3439,In_837,In_2506);
or U3440 (N_3440,In_2203,In_634);
and U3441 (N_3441,In_17,In_2980);
and U3442 (N_3442,In_1363,In_1956);
nand U3443 (N_3443,In_800,In_1926);
and U3444 (N_3444,In_788,In_909);
or U3445 (N_3445,In_1883,In_2648);
or U3446 (N_3446,In_1116,In_2705);
nor U3447 (N_3447,In_237,In_126);
nor U3448 (N_3448,In_1854,In_520);
xnor U3449 (N_3449,In_2173,In_2082);
nor U3450 (N_3450,In_2057,In_2805);
nand U3451 (N_3451,In_109,In_2958);
nor U3452 (N_3452,In_589,In_789);
or U3453 (N_3453,In_19,In_1993);
nand U3454 (N_3454,In_692,In_1942);
xor U3455 (N_3455,In_1286,In_693);
and U3456 (N_3456,In_326,In_2831);
xor U3457 (N_3457,In_2997,In_1683);
or U3458 (N_3458,In_374,In_739);
or U3459 (N_3459,In_1011,In_2875);
nor U3460 (N_3460,In_410,In_2581);
xor U3461 (N_3461,In_1466,In_1210);
nand U3462 (N_3462,In_1224,In_654);
or U3463 (N_3463,In_643,In_1093);
and U3464 (N_3464,In_1777,In_2850);
xnor U3465 (N_3465,In_79,In_1835);
nor U3466 (N_3466,In_2032,In_2148);
nor U3467 (N_3467,In_1248,In_1242);
nand U3468 (N_3468,In_1852,In_700);
nand U3469 (N_3469,In_1943,In_850);
nand U3470 (N_3470,In_957,In_667);
and U3471 (N_3471,In_867,In_1754);
and U3472 (N_3472,In_2278,In_2225);
and U3473 (N_3473,In_2869,In_2033);
nand U3474 (N_3474,In_379,In_2585);
and U3475 (N_3475,In_2140,In_1247);
and U3476 (N_3476,In_678,In_640);
nor U3477 (N_3477,In_1726,In_2776);
nand U3478 (N_3478,In_2461,In_2587);
nor U3479 (N_3479,In_803,In_218);
nor U3480 (N_3480,In_347,In_1863);
nor U3481 (N_3481,In_2434,In_1074);
and U3482 (N_3482,In_1207,In_572);
xnor U3483 (N_3483,In_2753,In_1882);
nand U3484 (N_3484,In_2349,In_2287);
nor U3485 (N_3485,In_2085,In_1164);
nand U3486 (N_3486,In_1866,In_195);
xnor U3487 (N_3487,In_2778,In_992);
nor U3488 (N_3488,In_1348,In_2219);
nand U3489 (N_3489,In_979,In_1933);
xor U3490 (N_3490,In_1762,In_85);
or U3491 (N_3491,In_1489,In_83);
or U3492 (N_3492,In_1130,In_1647);
or U3493 (N_3493,In_838,In_1478);
nor U3494 (N_3494,In_2225,In_1862);
nor U3495 (N_3495,In_2609,In_1865);
and U3496 (N_3496,In_1086,In_1456);
nand U3497 (N_3497,In_2802,In_1166);
xor U3498 (N_3498,In_1369,In_2547);
xor U3499 (N_3499,In_771,In_2194);
nand U3500 (N_3500,In_1853,In_1260);
and U3501 (N_3501,In_824,In_897);
and U3502 (N_3502,In_642,In_2071);
and U3503 (N_3503,In_51,In_38);
nand U3504 (N_3504,In_2840,In_909);
or U3505 (N_3505,In_2584,In_560);
xnor U3506 (N_3506,In_1689,In_1503);
nor U3507 (N_3507,In_796,In_2866);
nand U3508 (N_3508,In_1861,In_323);
or U3509 (N_3509,In_1623,In_494);
nor U3510 (N_3510,In_1270,In_1117);
or U3511 (N_3511,In_139,In_1667);
or U3512 (N_3512,In_9,In_1835);
xor U3513 (N_3513,In_338,In_557);
or U3514 (N_3514,In_2614,In_685);
xnor U3515 (N_3515,In_2441,In_255);
nor U3516 (N_3516,In_99,In_850);
and U3517 (N_3517,In_2403,In_993);
or U3518 (N_3518,In_2512,In_282);
nand U3519 (N_3519,In_2026,In_2031);
nand U3520 (N_3520,In_730,In_1298);
and U3521 (N_3521,In_2219,In_2901);
xor U3522 (N_3522,In_1752,In_1915);
and U3523 (N_3523,In_1947,In_254);
and U3524 (N_3524,In_2450,In_1561);
xnor U3525 (N_3525,In_16,In_2867);
or U3526 (N_3526,In_1460,In_572);
or U3527 (N_3527,In_1578,In_560);
or U3528 (N_3528,In_1927,In_1668);
and U3529 (N_3529,In_1270,In_1892);
or U3530 (N_3530,In_329,In_66);
nand U3531 (N_3531,In_2151,In_1884);
nor U3532 (N_3532,In_710,In_442);
or U3533 (N_3533,In_563,In_1866);
or U3534 (N_3534,In_2853,In_2194);
or U3535 (N_3535,In_2138,In_237);
nand U3536 (N_3536,In_867,In_1519);
nand U3537 (N_3537,In_1152,In_666);
and U3538 (N_3538,In_1562,In_2998);
or U3539 (N_3539,In_296,In_528);
and U3540 (N_3540,In_527,In_1565);
or U3541 (N_3541,In_2343,In_879);
nand U3542 (N_3542,In_2660,In_2644);
nor U3543 (N_3543,In_2105,In_1677);
nand U3544 (N_3544,In_351,In_1412);
or U3545 (N_3545,In_2887,In_283);
nand U3546 (N_3546,In_368,In_2061);
xor U3547 (N_3547,In_789,In_1362);
or U3548 (N_3548,In_226,In_2489);
xnor U3549 (N_3549,In_1967,In_431);
nor U3550 (N_3550,In_915,In_2996);
nand U3551 (N_3551,In_353,In_1135);
xnor U3552 (N_3552,In_2621,In_2011);
nor U3553 (N_3553,In_2701,In_2061);
nor U3554 (N_3554,In_654,In_1085);
and U3555 (N_3555,In_1123,In_2166);
or U3556 (N_3556,In_1108,In_597);
or U3557 (N_3557,In_1201,In_1763);
nor U3558 (N_3558,In_1551,In_825);
xnor U3559 (N_3559,In_1922,In_260);
nand U3560 (N_3560,In_681,In_924);
or U3561 (N_3561,In_991,In_1435);
or U3562 (N_3562,In_1360,In_1181);
and U3563 (N_3563,In_1532,In_2736);
nor U3564 (N_3564,In_2634,In_616);
nand U3565 (N_3565,In_1689,In_2273);
nor U3566 (N_3566,In_543,In_830);
nor U3567 (N_3567,In_728,In_1533);
and U3568 (N_3568,In_2435,In_2418);
nor U3569 (N_3569,In_1585,In_2211);
or U3570 (N_3570,In_2472,In_1071);
and U3571 (N_3571,In_231,In_1502);
nand U3572 (N_3572,In_657,In_2851);
nand U3573 (N_3573,In_2604,In_331);
xnor U3574 (N_3574,In_351,In_2948);
xnor U3575 (N_3575,In_1194,In_2012);
nor U3576 (N_3576,In_2419,In_2393);
nor U3577 (N_3577,In_995,In_2249);
or U3578 (N_3578,In_185,In_1058);
xor U3579 (N_3579,In_2179,In_1770);
and U3580 (N_3580,In_1447,In_1122);
xnor U3581 (N_3581,In_1499,In_1046);
xnor U3582 (N_3582,In_1590,In_2844);
nand U3583 (N_3583,In_561,In_330);
nand U3584 (N_3584,In_1281,In_1706);
xor U3585 (N_3585,In_507,In_1076);
or U3586 (N_3586,In_1135,In_1038);
nor U3587 (N_3587,In_634,In_877);
xnor U3588 (N_3588,In_1874,In_1539);
nand U3589 (N_3589,In_141,In_380);
and U3590 (N_3590,In_584,In_1008);
and U3591 (N_3591,In_1560,In_1261);
nor U3592 (N_3592,In_1726,In_939);
xnor U3593 (N_3593,In_132,In_762);
xor U3594 (N_3594,In_284,In_427);
xnor U3595 (N_3595,In_2240,In_1521);
xnor U3596 (N_3596,In_1692,In_1044);
and U3597 (N_3597,In_610,In_285);
nand U3598 (N_3598,In_19,In_1306);
or U3599 (N_3599,In_1254,In_1435);
xnor U3600 (N_3600,In_929,In_1356);
nor U3601 (N_3601,In_2743,In_2339);
xnor U3602 (N_3602,In_1148,In_2722);
nand U3603 (N_3603,In_376,In_1818);
and U3604 (N_3604,In_1012,In_2690);
nor U3605 (N_3605,In_774,In_2932);
or U3606 (N_3606,In_1400,In_1785);
nor U3607 (N_3607,In_2777,In_1944);
nand U3608 (N_3608,In_2625,In_1986);
nor U3609 (N_3609,In_1362,In_229);
or U3610 (N_3610,In_1955,In_2508);
nor U3611 (N_3611,In_729,In_495);
and U3612 (N_3612,In_190,In_592);
xor U3613 (N_3613,In_562,In_2706);
and U3614 (N_3614,In_1348,In_2586);
xor U3615 (N_3615,In_1338,In_1019);
or U3616 (N_3616,In_199,In_2402);
xnor U3617 (N_3617,In_637,In_1260);
nor U3618 (N_3618,In_1971,In_561);
and U3619 (N_3619,In_1981,In_457);
or U3620 (N_3620,In_1701,In_755);
and U3621 (N_3621,In_43,In_2986);
nor U3622 (N_3622,In_1416,In_2240);
or U3623 (N_3623,In_1056,In_2882);
and U3624 (N_3624,In_1236,In_1700);
xor U3625 (N_3625,In_1943,In_907);
or U3626 (N_3626,In_1512,In_1251);
and U3627 (N_3627,In_1361,In_1288);
and U3628 (N_3628,In_1153,In_542);
and U3629 (N_3629,In_274,In_1926);
nor U3630 (N_3630,In_792,In_1773);
and U3631 (N_3631,In_2974,In_687);
xor U3632 (N_3632,In_2215,In_2699);
or U3633 (N_3633,In_1395,In_647);
or U3634 (N_3634,In_2149,In_2315);
nand U3635 (N_3635,In_2011,In_1034);
or U3636 (N_3636,In_1816,In_640);
xor U3637 (N_3637,In_1086,In_1284);
xnor U3638 (N_3638,In_1894,In_1019);
nand U3639 (N_3639,In_176,In_2038);
xor U3640 (N_3640,In_43,In_2415);
or U3641 (N_3641,In_2544,In_514);
and U3642 (N_3642,In_482,In_2653);
nand U3643 (N_3643,In_2694,In_1161);
nand U3644 (N_3644,In_1794,In_1890);
nand U3645 (N_3645,In_2450,In_273);
or U3646 (N_3646,In_261,In_378);
nor U3647 (N_3647,In_1626,In_380);
nor U3648 (N_3648,In_427,In_939);
xor U3649 (N_3649,In_987,In_452);
nor U3650 (N_3650,In_445,In_1607);
and U3651 (N_3651,In_2720,In_1358);
nor U3652 (N_3652,In_189,In_519);
nor U3653 (N_3653,In_702,In_815);
or U3654 (N_3654,In_2635,In_2499);
and U3655 (N_3655,In_440,In_1733);
and U3656 (N_3656,In_238,In_2429);
nor U3657 (N_3657,In_510,In_1545);
or U3658 (N_3658,In_2326,In_2224);
nor U3659 (N_3659,In_871,In_2225);
nand U3660 (N_3660,In_291,In_11);
xnor U3661 (N_3661,In_1864,In_1934);
or U3662 (N_3662,In_1422,In_2083);
xnor U3663 (N_3663,In_2980,In_2740);
nor U3664 (N_3664,In_1351,In_2457);
nor U3665 (N_3665,In_218,In_2079);
and U3666 (N_3666,In_95,In_2921);
and U3667 (N_3667,In_1068,In_1274);
nand U3668 (N_3668,In_1500,In_411);
and U3669 (N_3669,In_257,In_481);
xor U3670 (N_3670,In_86,In_594);
xor U3671 (N_3671,In_574,In_1473);
xnor U3672 (N_3672,In_2711,In_2564);
nor U3673 (N_3673,In_1247,In_1142);
nand U3674 (N_3674,In_519,In_1699);
and U3675 (N_3675,In_945,In_2735);
or U3676 (N_3676,In_1647,In_2697);
and U3677 (N_3677,In_207,In_2565);
and U3678 (N_3678,In_2596,In_1261);
nand U3679 (N_3679,In_479,In_2902);
or U3680 (N_3680,In_2579,In_1768);
nand U3681 (N_3681,In_391,In_2076);
xor U3682 (N_3682,In_8,In_1017);
nor U3683 (N_3683,In_1443,In_158);
and U3684 (N_3684,In_2219,In_978);
nor U3685 (N_3685,In_653,In_2392);
nand U3686 (N_3686,In_1849,In_2088);
or U3687 (N_3687,In_2470,In_1985);
xnor U3688 (N_3688,In_1497,In_430);
nand U3689 (N_3689,In_2055,In_1156);
nand U3690 (N_3690,In_655,In_1499);
and U3691 (N_3691,In_2658,In_2230);
nor U3692 (N_3692,In_2210,In_1371);
and U3693 (N_3693,In_2782,In_970);
and U3694 (N_3694,In_1186,In_585);
xnor U3695 (N_3695,In_1423,In_2308);
nand U3696 (N_3696,In_2643,In_1782);
or U3697 (N_3697,In_597,In_1191);
or U3698 (N_3698,In_2303,In_506);
xor U3699 (N_3699,In_2777,In_632);
nor U3700 (N_3700,In_724,In_543);
xnor U3701 (N_3701,In_877,In_1271);
nand U3702 (N_3702,In_2910,In_873);
nand U3703 (N_3703,In_1616,In_2322);
xnor U3704 (N_3704,In_1815,In_2607);
or U3705 (N_3705,In_2312,In_277);
or U3706 (N_3706,In_1107,In_75);
nor U3707 (N_3707,In_1867,In_172);
xnor U3708 (N_3708,In_2848,In_1412);
or U3709 (N_3709,In_2576,In_685);
nand U3710 (N_3710,In_2321,In_2696);
and U3711 (N_3711,In_514,In_865);
nor U3712 (N_3712,In_1292,In_1071);
xnor U3713 (N_3713,In_1750,In_543);
nand U3714 (N_3714,In_1753,In_1328);
and U3715 (N_3715,In_1866,In_1205);
nor U3716 (N_3716,In_2820,In_2686);
nor U3717 (N_3717,In_203,In_1676);
and U3718 (N_3718,In_1500,In_1392);
or U3719 (N_3719,In_1983,In_1537);
and U3720 (N_3720,In_1637,In_692);
or U3721 (N_3721,In_2511,In_2796);
xor U3722 (N_3722,In_875,In_387);
and U3723 (N_3723,In_1128,In_2230);
and U3724 (N_3724,In_1154,In_2553);
nand U3725 (N_3725,In_1737,In_1915);
nor U3726 (N_3726,In_1101,In_2778);
xor U3727 (N_3727,In_744,In_435);
nand U3728 (N_3728,In_328,In_207);
or U3729 (N_3729,In_1327,In_159);
or U3730 (N_3730,In_1795,In_1931);
nor U3731 (N_3731,In_1330,In_82);
and U3732 (N_3732,In_376,In_1316);
or U3733 (N_3733,In_467,In_2929);
nand U3734 (N_3734,In_1141,In_1255);
xnor U3735 (N_3735,In_1421,In_790);
nand U3736 (N_3736,In_2595,In_1079);
or U3737 (N_3737,In_503,In_1526);
and U3738 (N_3738,In_1808,In_2970);
nor U3739 (N_3739,In_2872,In_748);
nor U3740 (N_3740,In_796,In_2023);
xnor U3741 (N_3741,In_1304,In_2614);
or U3742 (N_3742,In_325,In_1593);
nand U3743 (N_3743,In_1364,In_2024);
or U3744 (N_3744,In_1143,In_507);
xor U3745 (N_3745,In_1453,In_2844);
xor U3746 (N_3746,In_184,In_690);
xnor U3747 (N_3747,In_2872,In_1398);
and U3748 (N_3748,In_2279,In_1283);
and U3749 (N_3749,In_2557,In_755);
nor U3750 (N_3750,In_637,In_661);
or U3751 (N_3751,In_1076,In_629);
nand U3752 (N_3752,In_1646,In_514);
and U3753 (N_3753,In_1092,In_321);
nand U3754 (N_3754,In_1119,In_2658);
nand U3755 (N_3755,In_2039,In_1390);
or U3756 (N_3756,In_1710,In_1773);
nor U3757 (N_3757,In_2253,In_120);
xor U3758 (N_3758,In_198,In_123);
or U3759 (N_3759,In_2356,In_511);
nor U3760 (N_3760,In_1639,In_974);
and U3761 (N_3761,In_1992,In_1203);
nor U3762 (N_3762,In_999,In_2416);
xor U3763 (N_3763,In_2054,In_1895);
nor U3764 (N_3764,In_615,In_1973);
and U3765 (N_3765,In_2380,In_1092);
nand U3766 (N_3766,In_1956,In_1938);
nand U3767 (N_3767,In_1038,In_1033);
or U3768 (N_3768,In_2311,In_838);
nor U3769 (N_3769,In_2771,In_718);
or U3770 (N_3770,In_1837,In_2777);
xnor U3771 (N_3771,In_2202,In_49);
nand U3772 (N_3772,In_2870,In_400);
nand U3773 (N_3773,In_2042,In_567);
xnor U3774 (N_3774,In_1642,In_325);
xnor U3775 (N_3775,In_226,In_2530);
nand U3776 (N_3776,In_338,In_1746);
and U3777 (N_3777,In_2520,In_2329);
and U3778 (N_3778,In_1870,In_2420);
or U3779 (N_3779,In_2717,In_328);
or U3780 (N_3780,In_1115,In_2159);
and U3781 (N_3781,In_1124,In_2652);
nand U3782 (N_3782,In_1025,In_727);
or U3783 (N_3783,In_2531,In_1787);
nand U3784 (N_3784,In_1032,In_2621);
and U3785 (N_3785,In_101,In_1551);
xor U3786 (N_3786,In_487,In_2329);
xor U3787 (N_3787,In_1388,In_1689);
or U3788 (N_3788,In_1020,In_1890);
nor U3789 (N_3789,In_2102,In_1773);
or U3790 (N_3790,In_1235,In_732);
xor U3791 (N_3791,In_2438,In_478);
xnor U3792 (N_3792,In_117,In_1915);
nor U3793 (N_3793,In_228,In_573);
nor U3794 (N_3794,In_2769,In_2147);
nand U3795 (N_3795,In_941,In_2406);
nor U3796 (N_3796,In_2812,In_2038);
nand U3797 (N_3797,In_447,In_168);
or U3798 (N_3798,In_1444,In_963);
xor U3799 (N_3799,In_2665,In_1851);
and U3800 (N_3800,In_2509,In_764);
or U3801 (N_3801,In_489,In_1532);
and U3802 (N_3802,In_1611,In_2621);
and U3803 (N_3803,In_1458,In_2459);
or U3804 (N_3804,In_1172,In_530);
or U3805 (N_3805,In_1772,In_2067);
and U3806 (N_3806,In_2920,In_823);
nor U3807 (N_3807,In_1442,In_1510);
or U3808 (N_3808,In_2429,In_936);
and U3809 (N_3809,In_2898,In_1265);
xor U3810 (N_3810,In_2590,In_244);
or U3811 (N_3811,In_2600,In_2895);
or U3812 (N_3812,In_2685,In_2848);
nor U3813 (N_3813,In_384,In_2740);
nor U3814 (N_3814,In_2405,In_1914);
nor U3815 (N_3815,In_2430,In_1001);
or U3816 (N_3816,In_2841,In_2749);
or U3817 (N_3817,In_382,In_1353);
nor U3818 (N_3818,In_272,In_1870);
and U3819 (N_3819,In_1608,In_17);
or U3820 (N_3820,In_319,In_1004);
and U3821 (N_3821,In_2499,In_1454);
nor U3822 (N_3822,In_2029,In_682);
and U3823 (N_3823,In_169,In_651);
or U3824 (N_3824,In_1037,In_1966);
nand U3825 (N_3825,In_2579,In_1241);
or U3826 (N_3826,In_1895,In_2866);
and U3827 (N_3827,In_1345,In_54);
and U3828 (N_3828,In_1685,In_2636);
nand U3829 (N_3829,In_115,In_974);
nand U3830 (N_3830,In_2349,In_174);
xor U3831 (N_3831,In_1729,In_1978);
or U3832 (N_3832,In_2985,In_1802);
xor U3833 (N_3833,In_1565,In_2829);
nor U3834 (N_3834,In_1883,In_853);
xnor U3835 (N_3835,In_164,In_1395);
or U3836 (N_3836,In_2588,In_768);
and U3837 (N_3837,In_2006,In_63);
or U3838 (N_3838,In_1732,In_2928);
nor U3839 (N_3839,In_823,In_56);
xnor U3840 (N_3840,In_1594,In_2244);
nand U3841 (N_3841,In_383,In_2606);
nor U3842 (N_3842,In_1904,In_2723);
xnor U3843 (N_3843,In_2564,In_1364);
nand U3844 (N_3844,In_379,In_2945);
nand U3845 (N_3845,In_626,In_2114);
nand U3846 (N_3846,In_528,In_525);
or U3847 (N_3847,In_2041,In_1830);
nand U3848 (N_3848,In_1697,In_1014);
nand U3849 (N_3849,In_2742,In_231);
xor U3850 (N_3850,In_1482,In_2292);
nor U3851 (N_3851,In_685,In_265);
xnor U3852 (N_3852,In_1310,In_2611);
xor U3853 (N_3853,In_1293,In_1407);
nor U3854 (N_3854,In_31,In_2048);
or U3855 (N_3855,In_2726,In_2377);
nand U3856 (N_3856,In_1041,In_1786);
xor U3857 (N_3857,In_942,In_2334);
nand U3858 (N_3858,In_451,In_2270);
nor U3859 (N_3859,In_2429,In_1472);
and U3860 (N_3860,In_1239,In_633);
or U3861 (N_3861,In_416,In_1753);
nand U3862 (N_3862,In_746,In_2858);
or U3863 (N_3863,In_1045,In_1679);
xnor U3864 (N_3864,In_1982,In_2143);
xnor U3865 (N_3865,In_1741,In_2553);
nor U3866 (N_3866,In_149,In_260);
nand U3867 (N_3867,In_1128,In_2116);
nor U3868 (N_3868,In_2319,In_1387);
and U3869 (N_3869,In_2407,In_1442);
nor U3870 (N_3870,In_923,In_120);
xor U3871 (N_3871,In_181,In_1669);
nand U3872 (N_3872,In_1772,In_2142);
nand U3873 (N_3873,In_378,In_91);
nor U3874 (N_3874,In_1155,In_2500);
nand U3875 (N_3875,In_621,In_767);
xnor U3876 (N_3876,In_2354,In_2155);
nor U3877 (N_3877,In_378,In_2761);
and U3878 (N_3878,In_2965,In_915);
or U3879 (N_3879,In_1625,In_748);
or U3880 (N_3880,In_1330,In_2368);
or U3881 (N_3881,In_2780,In_2502);
nand U3882 (N_3882,In_976,In_1633);
or U3883 (N_3883,In_146,In_552);
and U3884 (N_3884,In_1024,In_2871);
nand U3885 (N_3885,In_742,In_2523);
nand U3886 (N_3886,In_1320,In_231);
xnor U3887 (N_3887,In_1731,In_2183);
nand U3888 (N_3888,In_994,In_2950);
or U3889 (N_3889,In_1666,In_1609);
nand U3890 (N_3890,In_1467,In_2025);
nor U3891 (N_3891,In_119,In_985);
xnor U3892 (N_3892,In_626,In_1126);
xor U3893 (N_3893,In_1060,In_2756);
nor U3894 (N_3894,In_1687,In_97);
xnor U3895 (N_3895,In_764,In_2757);
nor U3896 (N_3896,In_2788,In_2157);
nand U3897 (N_3897,In_901,In_2370);
or U3898 (N_3898,In_2493,In_23);
xnor U3899 (N_3899,In_551,In_862);
nand U3900 (N_3900,In_2744,In_2269);
nor U3901 (N_3901,In_691,In_54);
or U3902 (N_3902,In_806,In_234);
nand U3903 (N_3903,In_2006,In_2057);
nor U3904 (N_3904,In_878,In_729);
or U3905 (N_3905,In_984,In_1282);
and U3906 (N_3906,In_1721,In_1626);
nand U3907 (N_3907,In_979,In_961);
nand U3908 (N_3908,In_434,In_344);
xor U3909 (N_3909,In_1723,In_414);
nand U3910 (N_3910,In_2027,In_2718);
nor U3911 (N_3911,In_1371,In_2371);
xnor U3912 (N_3912,In_1527,In_2688);
or U3913 (N_3913,In_1120,In_1653);
or U3914 (N_3914,In_2316,In_12);
nor U3915 (N_3915,In_2569,In_2465);
and U3916 (N_3916,In_2421,In_1447);
or U3917 (N_3917,In_501,In_558);
nand U3918 (N_3918,In_2283,In_554);
xnor U3919 (N_3919,In_111,In_2340);
xor U3920 (N_3920,In_101,In_998);
nor U3921 (N_3921,In_792,In_2373);
nor U3922 (N_3922,In_2566,In_1072);
nand U3923 (N_3923,In_1724,In_2312);
and U3924 (N_3924,In_639,In_285);
xnor U3925 (N_3925,In_1672,In_1457);
nor U3926 (N_3926,In_1972,In_1337);
xnor U3927 (N_3927,In_78,In_2580);
nand U3928 (N_3928,In_21,In_1236);
xnor U3929 (N_3929,In_782,In_268);
xnor U3930 (N_3930,In_1398,In_613);
nand U3931 (N_3931,In_918,In_637);
or U3932 (N_3932,In_2907,In_2405);
or U3933 (N_3933,In_1839,In_1676);
nor U3934 (N_3934,In_954,In_1404);
or U3935 (N_3935,In_1001,In_458);
or U3936 (N_3936,In_676,In_2051);
nor U3937 (N_3937,In_2038,In_423);
and U3938 (N_3938,In_1018,In_2271);
nor U3939 (N_3939,In_2451,In_526);
or U3940 (N_3940,In_689,In_2834);
nor U3941 (N_3941,In_1488,In_473);
nand U3942 (N_3942,In_726,In_914);
nor U3943 (N_3943,In_184,In_2464);
or U3944 (N_3944,In_770,In_1600);
or U3945 (N_3945,In_1316,In_2587);
or U3946 (N_3946,In_1039,In_526);
xor U3947 (N_3947,In_230,In_159);
xor U3948 (N_3948,In_2055,In_2497);
nor U3949 (N_3949,In_2346,In_1071);
nor U3950 (N_3950,In_739,In_2120);
xnor U3951 (N_3951,In_804,In_2686);
nand U3952 (N_3952,In_118,In_376);
xnor U3953 (N_3953,In_391,In_1595);
and U3954 (N_3954,In_1317,In_1960);
nand U3955 (N_3955,In_2852,In_2744);
nand U3956 (N_3956,In_1791,In_2080);
or U3957 (N_3957,In_1607,In_1518);
and U3958 (N_3958,In_1561,In_1091);
xor U3959 (N_3959,In_2248,In_1026);
nand U3960 (N_3960,In_308,In_2280);
or U3961 (N_3961,In_1076,In_338);
nor U3962 (N_3962,In_2796,In_982);
xnor U3963 (N_3963,In_2283,In_1249);
nor U3964 (N_3964,In_2594,In_2786);
xor U3965 (N_3965,In_264,In_2711);
and U3966 (N_3966,In_555,In_1000);
or U3967 (N_3967,In_2284,In_2204);
or U3968 (N_3968,In_1491,In_548);
xnor U3969 (N_3969,In_1200,In_162);
nand U3970 (N_3970,In_1434,In_861);
xor U3971 (N_3971,In_1244,In_387);
and U3972 (N_3972,In_2075,In_1689);
nand U3973 (N_3973,In_2460,In_2743);
nor U3974 (N_3974,In_74,In_2560);
nand U3975 (N_3975,In_1230,In_55);
or U3976 (N_3976,In_2695,In_2605);
nor U3977 (N_3977,In_1686,In_362);
xor U3978 (N_3978,In_1743,In_2456);
xor U3979 (N_3979,In_2791,In_2348);
or U3980 (N_3980,In_163,In_723);
and U3981 (N_3981,In_2239,In_1483);
or U3982 (N_3982,In_2269,In_2049);
xnor U3983 (N_3983,In_2222,In_2301);
xor U3984 (N_3984,In_2630,In_1744);
and U3985 (N_3985,In_2549,In_1063);
nor U3986 (N_3986,In_505,In_1831);
xnor U3987 (N_3987,In_469,In_1238);
nand U3988 (N_3988,In_1353,In_2474);
and U3989 (N_3989,In_2096,In_107);
nand U3990 (N_3990,In_2548,In_2251);
nor U3991 (N_3991,In_181,In_1476);
nand U3992 (N_3992,In_619,In_87);
nand U3993 (N_3993,In_1423,In_1994);
nor U3994 (N_3994,In_2992,In_2158);
xnor U3995 (N_3995,In_1438,In_1081);
xnor U3996 (N_3996,In_406,In_1346);
and U3997 (N_3997,In_1028,In_1349);
nand U3998 (N_3998,In_526,In_2978);
and U3999 (N_3999,In_1133,In_641);
and U4000 (N_4000,In_1827,In_2510);
nor U4001 (N_4001,In_1946,In_323);
and U4002 (N_4002,In_691,In_1362);
or U4003 (N_4003,In_2400,In_2101);
or U4004 (N_4004,In_2722,In_183);
nor U4005 (N_4005,In_1160,In_467);
nand U4006 (N_4006,In_757,In_660);
nand U4007 (N_4007,In_892,In_1939);
and U4008 (N_4008,In_471,In_1625);
or U4009 (N_4009,In_1727,In_2503);
xor U4010 (N_4010,In_301,In_2337);
nand U4011 (N_4011,In_1227,In_337);
and U4012 (N_4012,In_1786,In_951);
nand U4013 (N_4013,In_20,In_1040);
and U4014 (N_4014,In_1517,In_2142);
xor U4015 (N_4015,In_618,In_1786);
or U4016 (N_4016,In_217,In_1062);
or U4017 (N_4017,In_1521,In_1292);
and U4018 (N_4018,In_1669,In_1230);
nand U4019 (N_4019,In_1026,In_2112);
nor U4020 (N_4020,In_1237,In_1747);
nand U4021 (N_4021,In_2793,In_1599);
xor U4022 (N_4022,In_529,In_1642);
nand U4023 (N_4023,In_2127,In_2118);
xor U4024 (N_4024,In_2313,In_2776);
xor U4025 (N_4025,In_1184,In_91);
and U4026 (N_4026,In_1089,In_1225);
xnor U4027 (N_4027,In_2166,In_2079);
and U4028 (N_4028,In_388,In_1191);
or U4029 (N_4029,In_1474,In_860);
or U4030 (N_4030,In_2530,In_31);
xor U4031 (N_4031,In_2601,In_2495);
and U4032 (N_4032,In_517,In_306);
and U4033 (N_4033,In_943,In_2145);
and U4034 (N_4034,In_959,In_625);
or U4035 (N_4035,In_36,In_862);
nor U4036 (N_4036,In_710,In_1616);
nand U4037 (N_4037,In_581,In_1855);
xor U4038 (N_4038,In_2020,In_2319);
xnor U4039 (N_4039,In_1606,In_2478);
xor U4040 (N_4040,In_2403,In_1172);
xnor U4041 (N_4041,In_2348,In_27);
nor U4042 (N_4042,In_1405,In_1543);
and U4043 (N_4043,In_1651,In_2671);
nor U4044 (N_4044,In_2226,In_1585);
nand U4045 (N_4045,In_546,In_2340);
or U4046 (N_4046,In_1259,In_37);
nor U4047 (N_4047,In_2727,In_1610);
and U4048 (N_4048,In_1193,In_817);
nor U4049 (N_4049,In_941,In_1542);
or U4050 (N_4050,In_1488,In_353);
nor U4051 (N_4051,In_1157,In_2754);
or U4052 (N_4052,In_2137,In_209);
and U4053 (N_4053,In_694,In_495);
xnor U4054 (N_4054,In_742,In_734);
and U4055 (N_4055,In_2608,In_1179);
or U4056 (N_4056,In_1423,In_369);
nor U4057 (N_4057,In_2604,In_64);
nand U4058 (N_4058,In_495,In_2387);
or U4059 (N_4059,In_2167,In_1294);
and U4060 (N_4060,In_408,In_659);
and U4061 (N_4061,In_1368,In_334);
nor U4062 (N_4062,In_1791,In_2590);
nand U4063 (N_4063,In_921,In_2610);
and U4064 (N_4064,In_400,In_1557);
and U4065 (N_4065,In_286,In_1506);
or U4066 (N_4066,In_2479,In_2912);
and U4067 (N_4067,In_1279,In_1178);
nor U4068 (N_4068,In_2268,In_2102);
or U4069 (N_4069,In_1609,In_2843);
xor U4070 (N_4070,In_469,In_2393);
nor U4071 (N_4071,In_2155,In_233);
nor U4072 (N_4072,In_2066,In_2117);
xnor U4073 (N_4073,In_1769,In_1178);
or U4074 (N_4074,In_2049,In_2672);
and U4075 (N_4075,In_2909,In_220);
or U4076 (N_4076,In_2561,In_740);
or U4077 (N_4077,In_1394,In_2812);
xnor U4078 (N_4078,In_2452,In_1497);
and U4079 (N_4079,In_967,In_189);
or U4080 (N_4080,In_2361,In_594);
nand U4081 (N_4081,In_1904,In_167);
or U4082 (N_4082,In_2286,In_426);
and U4083 (N_4083,In_1600,In_2823);
and U4084 (N_4084,In_1092,In_350);
or U4085 (N_4085,In_2034,In_2196);
xor U4086 (N_4086,In_1678,In_284);
and U4087 (N_4087,In_2126,In_1486);
nand U4088 (N_4088,In_2921,In_1483);
nand U4089 (N_4089,In_911,In_2331);
nor U4090 (N_4090,In_1929,In_2919);
xor U4091 (N_4091,In_736,In_249);
nor U4092 (N_4092,In_2321,In_2805);
nand U4093 (N_4093,In_958,In_2333);
and U4094 (N_4094,In_1081,In_673);
xor U4095 (N_4095,In_620,In_395);
and U4096 (N_4096,In_2169,In_607);
and U4097 (N_4097,In_1861,In_1068);
or U4098 (N_4098,In_1625,In_1007);
xor U4099 (N_4099,In_1079,In_433);
nand U4100 (N_4100,In_1689,In_2429);
xnor U4101 (N_4101,In_43,In_2855);
xor U4102 (N_4102,In_1341,In_2791);
nor U4103 (N_4103,In_1396,In_2331);
xor U4104 (N_4104,In_625,In_2365);
or U4105 (N_4105,In_293,In_1626);
xnor U4106 (N_4106,In_2121,In_550);
nor U4107 (N_4107,In_2121,In_1628);
xor U4108 (N_4108,In_1464,In_635);
xor U4109 (N_4109,In_1187,In_2789);
xnor U4110 (N_4110,In_593,In_484);
or U4111 (N_4111,In_1251,In_864);
nand U4112 (N_4112,In_826,In_2467);
nand U4113 (N_4113,In_2960,In_710);
nand U4114 (N_4114,In_1575,In_2821);
xor U4115 (N_4115,In_1847,In_2396);
nor U4116 (N_4116,In_2514,In_2096);
nand U4117 (N_4117,In_285,In_1298);
nor U4118 (N_4118,In_1143,In_1210);
xnor U4119 (N_4119,In_382,In_52);
and U4120 (N_4120,In_2066,In_2212);
xor U4121 (N_4121,In_1015,In_324);
nor U4122 (N_4122,In_246,In_548);
nor U4123 (N_4123,In_1400,In_1057);
and U4124 (N_4124,In_1168,In_1599);
and U4125 (N_4125,In_1077,In_1534);
nand U4126 (N_4126,In_112,In_2875);
xor U4127 (N_4127,In_2820,In_1542);
and U4128 (N_4128,In_2895,In_1501);
xnor U4129 (N_4129,In_2703,In_693);
xnor U4130 (N_4130,In_318,In_852);
xnor U4131 (N_4131,In_1505,In_256);
nor U4132 (N_4132,In_103,In_1429);
or U4133 (N_4133,In_1604,In_673);
nand U4134 (N_4134,In_1140,In_2496);
nor U4135 (N_4135,In_291,In_1162);
xor U4136 (N_4136,In_2038,In_72);
nor U4137 (N_4137,In_1477,In_224);
xnor U4138 (N_4138,In_2424,In_1362);
and U4139 (N_4139,In_494,In_789);
or U4140 (N_4140,In_2064,In_2376);
and U4141 (N_4141,In_1551,In_2140);
and U4142 (N_4142,In_531,In_1380);
xor U4143 (N_4143,In_1855,In_1613);
and U4144 (N_4144,In_250,In_1902);
nand U4145 (N_4145,In_534,In_876);
or U4146 (N_4146,In_1324,In_1216);
and U4147 (N_4147,In_1196,In_2013);
or U4148 (N_4148,In_33,In_1838);
nand U4149 (N_4149,In_1288,In_2029);
nor U4150 (N_4150,In_548,In_665);
nand U4151 (N_4151,In_1705,In_1352);
or U4152 (N_4152,In_528,In_638);
or U4153 (N_4153,In_1437,In_965);
nand U4154 (N_4154,In_577,In_579);
and U4155 (N_4155,In_1395,In_1936);
xnor U4156 (N_4156,In_1174,In_1037);
nor U4157 (N_4157,In_687,In_1444);
nor U4158 (N_4158,In_1620,In_1793);
and U4159 (N_4159,In_2021,In_214);
xnor U4160 (N_4160,In_1083,In_1414);
and U4161 (N_4161,In_2393,In_91);
nand U4162 (N_4162,In_1646,In_2880);
xnor U4163 (N_4163,In_94,In_821);
xnor U4164 (N_4164,In_1639,In_1487);
nand U4165 (N_4165,In_976,In_49);
nand U4166 (N_4166,In_705,In_160);
nand U4167 (N_4167,In_835,In_1842);
and U4168 (N_4168,In_1788,In_1565);
and U4169 (N_4169,In_2111,In_129);
nor U4170 (N_4170,In_1526,In_1512);
nand U4171 (N_4171,In_0,In_179);
nor U4172 (N_4172,In_537,In_2908);
xor U4173 (N_4173,In_361,In_2163);
or U4174 (N_4174,In_2792,In_2383);
nor U4175 (N_4175,In_411,In_867);
and U4176 (N_4176,In_2140,In_1286);
xnor U4177 (N_4177,In_2311,In_1499);
nor U4178 (N_4178,In_1976,In_2948);
or U4179 (N_4179,In_1783,In_948);
xor U4180 (N_4180,In_781,In_2570);
nor U4181 (N_4181,In_2478,In_421);
nor U4182 (N_4182,In_2276,In_702);
and U4183 (N_4183,In_2491,In_1007);
xor U4184 (N_4184,In_1508,In_1920);
and U4185 (N_4185,In_2121,In_2638);
or U4186 (N_4186,In_386,In_1986);
xnor U4187 (N_4187,In_2429,In_183);
nand U4188 (N_4188,In_126,In_782);
and U4189 (N_4189,In_1917,In_479);
xor U4190 (N_4190,In_512,In_481);
nor U4191 (N_4191,In_924,In_39);
and U4192 (N_4192,In_919,In_2851);
nor U4193 (N_4193,In_4,In_1876);
nor U4194 (N_4194,In_812,In_2633);
nor U4195 (N_4195,In_819,In_1014);
xnor U4196 (N_4196,In_728,In_1187);
and U4197 (N_4197,In_1428,In_443);
or U4198 (N_4198,In_2731,In_2819);
nor U4199 (N_4199,In_2704,In_2701);
nor U4200 (N_4200,In_2438,In_1788);
or U4201 (N_4201,In_2762,In_52);
nor U4202 (N_4202,In_56,In_1265);
nand U4203 (N_4203,In_76,In_2138);
xor U4204 (N_4204,In_1017,In_533);
nor U4205 (N_4205,In_356,In_1232);
and U4206 (N_4206,In_223,In_1535);
nor U4207 (N_4207,In_691,In_1168);
and U4208 (N_4208,In_1183,In_1143);
nand U4209 (N_4209,In_1078,In_2077);
nand U4210 (N_4210,In_1137,In_741);
and U4211 (N_4211,In_1878,In_2572);
and U4212 (N_4212,In_2377,In_1127);
nand U4213 (N_4213,In_122,In_316);
nor U4214 (N_4214,In_915,In_2666);
nor U4215 (N_4215,In_1190,In_2380);
and U4216 (N_4216,In_830,In_1281);
xor U4217 (N_4217,In_1079,In_1314);
and U4218 (N_4218,In_453,In_56);
nor U4219 (N_4219,In_1068,In_2912);
nand U4220 (N_4220,In_2282,In_314);
or U4221 (N_4221,In_2703,In_1370);
or U4222 (N_4222,In_102,In_1771);
nand U4223 (N_4223,In_1825,In_340);
nand U4224 (N_4224,In_249,In_2062);
or U4225 (N_4225,In_1509,In_274);
and U4226 (N_4226,In_2285,In_1328);
nand U4227 (N_4227,In_2338,In_305);
or U4228 (N_4228,In_886,In_1651);
xnor U4229 (N_4229,In_651,In_2678);
nor U4230 (N_4230,In_2453,In_897);
xnor U4231 (N_4231,In_130,In_2416);
xnor U4232 (N_4232,In_362,In_2741);
nand U4233 (N_4233,In_2090,In_458);
xor U4234 (N_4234,In_556,In_2457);
or U4235 (N_4235,In_1507,In_1793);
xnor U4236 (N_4236,In_1498,In_1162);
or U4237 (N_4237,In_2363,In_2809);
or U4238 (N_4238,In_2403,In_387);
or U4239 (N_4239,In_510,In_1891);
xor U4240 (N_4240,In_252,In_2494);
nor U4241 (N_4241,In_244,In_425);
nor U4242 (N_4242,In_2973,In_2722);
and U4243 (N_4243,In_2184,In_1673);
nand U4244 (N_4244,In_2599,In_1933);
and U4245 (N_4245,In_2355,In_1421);
nor U4246 (N_4246,In_1184,In_2387);
nor U4247 (N_4247,In_2897,In_1001);
xor U4248 (N_4248,In_1331,In_14);
nor U4249 (N_4249,In_794,In_1606);
nand U4250 (N_4250,In_2579,In_710);
nand U4251 (N_4251,In_1813,In_324);
nand U4252 (N_4252,In_1330,In_1291);
nand U4253 (N_4253,In_2275,In_342);
xnor U4254 (N_4254,In_279,In_227);
and U4255 (N_4255,In_2713,In_1870);
nand U4256 (N_4256,In_64,In_1922);
or U4257 (N_4257,In_302,In_440);
or U4258 (N_4258,In_2725,In_518);
or U4259 (N_4259,In_134,In_2650);
xnor U4260 (N_4260,In_1786,In_2406);
or U4261 (N_4261,In_2820,In_824);
nor U4262 (N_4262,In_2822,In_1723);
xor U4263 (N_4263,In_1791,In_2821);
nor U4264 (N_4264,In_1635,In_2335);
and U4265 (N_4265,In_2462,In_489);
nand U4266 (N_4266,In_2115,In_794);
nand U4267 (N_4267,In_1887,In_1788);
nor U4268 (N_4268,In_1635,In_97);
and U4269 (N_4269,In_870,In_1843);
nand U4270 (N_4270,In_351,In_2161);
and U4271 (N_4271,In_1276,In_55);
and U4272 (N_4272,In_1631,In_2626);
nand U4273 (N_4273,In_1087,In_1855);
nor U4274 (N_4274,In_398,In_942);
xnor U4275 (N_4275,In_2680,In_2269);
or U4276 (N_4276,In_1723,In_2921);
nand U4277 (N_4277,In_2250,In_2261);
and U4278 (N_4278,In_851,In_2091);
nor U4279 (N_4279,In_2693,In_1557);
nand U4280 (N_4280,In_2693,In_2796);
and U4281 (N_4281,In_2638,In_2482);
xnor U4282 (N_4282,In_2667,In_2570);
xnor U4283 (N_4283,In_1021,In_1854);
or U4284 (N_4284,In_2695,In_108);
or U4285 (N_4285,In_2132,In_228);
xor U4286 (N_4286,In_312,In_2244);
nand U4287 (N_4287,In_2675,In_2757);
and U4288 (N_4288,In_2759,In_1384);
or U4289 (N_4289,In_154,In_238);
nand U4290 (N_4290,In_1953,In_1075);
or U4291 (N_4291,In_1791,In_365);
nand U4292 (N_4292,In_2046,In_1219);
nor U4293 (N_4293,In_26,In_761);
xor U4294 (N_4294,In_1921,In_781);
nand U4295 (N_4295,In_918,In_2517);
nor U4296 (N_4296,In_925,In_2065);
xor U4297 (N_4297,In_2774,In_2397);
xnor U4298 (N_4298,In_449,In_1160);
nand U4299 (N_4299,In_1430,In_588);
or U4300 (N_4300,In_1528,In_1157);
xnor U4301 (N_4301,In_2651,In_89);
nor U4302 (N_4302,In_1951,In_2961);
nand U4303 (N_4303,In_1553,In_1353);
nand U4304 (N_4304,In_2421,In_1586);
xnor U4305 (N_4305,In_2987,In_210);
or U4306 (N_4306,In_2795,In_2210);
or U4307 (N_4307,In_208,In_1525);
xnor U4308 (N_4308,In_2539,In_2703);
xnor U4309 (N_4309,In_891,In_2660);
xor U4310 (N_4310,In_1248,In_2878);
or U4311 (N_4311,In_401,In_185);
nand U4312 (N_4312,In_872,In_124);
and U4313 (N_4313,In_1686,In_2324);
nor U4314 (N_4314,In_109,In_1609);
nand U4315 (N_4315,In_940,In_1749);
or U4316 (N_4316,In_1798,In_1511);
or U4317 (N_4317,In_609,In_2011);
xnor U4318 (N_4318,In_2258,In_1514);
nor U4319 (N_4319,In_2201,In_2808);
nor U4320 (N_4320,In_114,In_2224);
and U4321 (N_4321,In_1407,In_2094);
and U4322 (N_4322,In_2922,In_2076);
xor U4323 (N_4323,In_608,In_1143);
or U4324 (N_4324,In_1595,In_2970);
or U4325 (N_4325,In_985,In_711);
nor U4326 (N_4326,In_2687,In_1960);
and U4327 (N_4327,In_2362,In_1733);
nand U4328 (N_4328,In_515,In_2815);
and U4329 (N_4329,In_18,In_725);
or U4330 (N_4330,In_777,In_2586);
xor U4331 (N_4331,In_789,In_2036);
nand U4332 (N_4332,In_1302,In_51);
nor U4333 (N_4333,In_2868,In_565);
or U4334 (N_4334,In_1784,In_710);
xnor U4335 (N_4335,In_2233,In_2505);
and U4336 (N_4336,In_265,In_862);
and U4337 (N_4337,In_67,In_2215);
or U4338 (N_4338,In_2358,In_1024);
nor U4339 (N_4339,In_1051,In_1727);
and U4340 (N_4340,In_2287,In_121);
nand U4341 (N_4341,In_1355,In_1146);
xnor U4342 (N_4342,In_2231,In_2798);
nand U4343 (N_4343,In_690,In_2522);
xor U4344 (N_4344,In_763,In_1723);
and U4345 (N_4345,In_2769,In_3);
or U4346 (N_4346,In_1972,In_2118);
nor U4347 (N_4347,In_1984,In_2056);
and U4348 (N_4348,In_851,In_2581);
xor U4349 (N_4349,In_1835,In_1257);
or U4350 (N_4350,In_1020,In_1190);
nand U4351 (N_4351,In_928,In_1285);
or U4352 (N_4352,In_2670,In_1869);
nand U4353 (N_4353,In_2108,In_2479);
or U4354 (N_4354,In_2063,In_1996);
and U4355 (N_4355,In_1009,In_2475);
and U4356 (N_4356,In_773,In_1109);
and U4357 (N_4357,In_2372,In_1899);
or U4358 (N_4358,In_2588,In_1648);
and U4359 (N_4359,In_2676,In_1182);
nor U4360 (N_4360,In_2557,In_1651);
nor U4361 (N_4361,In_1850,In_1903);
xor U4362 (N_4362,In_2017,In_1413);
or U4363 (N_4363,In_1940,In_2747);
xnor U4364 (N_4364,In_124,In_1786);
xor U4365 (N_4365,In_2186,In_2781);
xnor U4366 (N_4366,In_1524,In_840);
or U4367 (N_4367,In_2199,In_2893);
and U4368 (N_4368,In_984,In_1302);
and U4369 (N_4369,In_395,In_2212);
nor U4370 (N_4370,In_584,In_318);
nor U4371 (N_4371,In_2927,In_2146);
and U4372 (N_4372,In_1066,In_2441);
xor U4373 (N_4373,In_107,In_2269);
xnor U4374 (N_4374,In_2000,In_2513);
or U4375 (N_4375,In_579,In_1098);
xnor U4376 (N_4376,In_2688,In_130);
nand U4377 (N_4377,In_1845,In_1323);
and U4378 (N_4378,In_302,In_648);
xnor U4379 (N_4379,In_572,In_696);
or U4380 (N_4380,In_2382,In_584);
nand U4381 (N_4381,In_1792,In_2497);
nand U4382 (N_4382,In_1121,In_2150);
xor U4383 (N_4383,In_967,In_346);
nand U4384 (N_4384,In_1001,In_2626);
nor U4385 (N_4385,In_516,In_2690);
nand U4386 (N_4386,In_69,In_80);
and U4387 (N_4387,In_548,In_780);
nand U4388 (N_4388,In_1940,In_2006);
or U4389 (N_4389,In_666,In_2045);
and U4390 (N_4390,In_457,In_1694);
or U4391 (N_4391,In_2552,In_1838);
and U4392 (N_4392,In_1355,In_1003);
and U4393 (N_4393,In_2638,In_1757);
xnor U4394 (N_4394,In_2234,In_1328);
xor U4395 (N_4395,In_1609,In_590);
xnor U4396 (N_4396,In_882,In_2178);
and U4397 (N_4397,In_338,In_2302);
nor U4398 (N_4398,In_2913,In_577);
nor U4399 (N_4399,In_1291,In_2013);
or U4400 (N_4400,In_258,In_2945);
or U4401 (N_4401,In_136,In_493);
nor U4402 (N_4402,In_2366,In_1818);
and U4403 (N_4403,In_493,In_1031);
xnor U4404 (N_4404,In_66,In_383);
or U4405 (N_4405,In_1996,In_541);
nor U4406 (N_4406,In_1319,In_1502);
and U4407 (N_4407,In_2146,In_2478);
or U4408 (N_4408,In_213,In_698);
and U4409 (N_4409,In_1454,In_3);
and U4410 (N_4410,In_2802,In_1773);
nor U4411 (N_4411,In_1163,In_291);
or U4412 (N_4412,In_211,In_2589);
xnor U4413 (N_4413,In_2835,In_2377);
xnor U4414 (N_4414,In_2953,In_1034);
nor U4415 (N_4415,In_1272,In_1764);
nor U4416 (N_4416,In_149,In_2223);
or U4417 (N_4417,In_2577,In_328);
xnor U4418 (N_4418,In_2616,In_2667);
xor U4419 (N_4419,In_1082,In_384);
or U4420 (N_4420,In_2724,In_2943);
nand U4421 (N_4421,In_2245,In_2758);
or U4422 (N_4422,In_888,In_370);
or U4423 (N_4423,In_352,In_2518);
or U4424 (N_4424,In_1414,In_2268);
nor U4425 (N_4425,In_2468,In_2845);
and U4426 (N_4426,In_606,In_2702);
xor U4427 (N_4427,In_1193,In_2816);
xnor U4428 (N_4428,In_487,In_2054);
or U4429 (N_4429,In_1811,In_2499);
and U4430 (N_4430,In_277,In_1941);
nor U4431 (N_4431,In_777,In_1512);
or U4432 (N_4432,In_1222,In_1330);
xnor U4433 (N_4433,In_1555,In_1881);
nand U4434 (N_4434,In_2992,In_2969);
xor U4435 (N_4435,In_2504,In_1841);
or U4436 (N_4436,In_2213,In_1685);
or U4437 (N_4437,In_1822,In_1423);
or U4438 (N_4438,In_2303,In_1843);
nand U4439 (N_4439,In_483,In_340);
xnor U4440 (N_4440,In_2620,In_1437);
nor U4441 (N_4441,In_1137,In_2612);
nor U4442 (N_4442,In_68,In_1701);
and U4443 (N_4443,In_75,In_1575);
and U4444 (N_4444,In_779,In_2812);
and U4445 (N_4445,In_184,In_719);
nor U4446 (N_4446,In_2688,In_292);
nand U4447 (N_4447,In_1838,In_603);
and U4448 (N_4448,In_416,In_1940);
nor U4449 (N_4449,In_2520,In_442);
nor U4450 (N_4450,In_2235,In_2961);
and U4451 (N_4451,In_140,In_1408);
xor U4452 (N_4452,In_1839,In_1439);
xor U4453 (N_4453,In_1598,In_2753);
nor U4454 (N_4454,In_61,In_2275);
and U4455 (N_4455,In_821,In_2199);
nor U4456 (N_4456,In_1135,In_1984);
xnor U4457 (N_4457,In_41,In_213);
and U4458 (N_4458,In_228,In_2497);
nand U4459 (N_4459,In_525,In_1593);
and U4460 (N_4460,In_887,In_2636);
or U4461 (N_4461,In_456,In_477);
nand U4462 (N_4462,In_199,In_1806);
nor U4463 (N_4463,In_1440,In_240);
xnor U4464 (N_4464,In_1576,In_1630);
nor U4465 (N_4465,In_1305,In_1956);
and U4466 (N_4466,In_1790,In_747);
or U4467 (N_4467,In_2457,In_2846);
nand U4468 (N_4468,In_2244,In_2506);
nor U4469 (N_4469,In_381,In_310);
or U4470 (N_4470,In_1094,In_1148);
xor U4471 (N_4471,In_917,In_1833);
or U4472 (N_4472,In_661,In_1247);
nand U4473 (N_4473,In_442,In_1137);
nand U4474 (N_4474,In_87,In_1353);
nor U4475 (N_4475,In_1438,In_145);
nand U4476 (N_4476,In_2750,In_1735);
and U4477 (N_4477,In_2805,In_1057);
or U4478 (N_4478,In_1452,In_587);
xor U4479 (N_4479,In_2139,In_1498);
nor U4480 (N_4480,In_2944,In_1616);
and U4481 (N_4481,In_1344,In_668);
and U4482 (N_4482,In_939,In_1247);
xnor U4483 (N_4483,In_2384,In_2687);
or U4484 (N_4484,In_1127,In_1384);
nor U4485 (N_4485,In_256,In_1638);
nand U4486 (N_4486,In_2510,In_2942);
nand U4487 (N_4487,In_1323,In_699);
nand U4488 (N_4488,In_2639,In_1543);
and U4489 (N_4489,In_1492,In_1682);
nor U4490 (N_4490,In_2296,In_1448);
xor U4491 (N_4491,In_570,In_2711);
xnor U4492 (N_4492,In_778,In_2366);
or U4493 (N_4493,In_882,In_2775);
and U4494 (N_4494,In_1776,In_2937);
xor U4495 (N_4495,In_1397,In_1747);
xnor U4496 (N_4496,In_2898,In_2764);
nor U4497 (N_4497,In_2216,In_1592);
and U4498 (N_4498,In_781,In_1364);
xnor U4499 (N_4499,In_943,In_1676);
nor U4500 (N_4500,In_1454,In_1466);
or U4501 (N_4501,In_1752,In_1507);
and U4502 (N_4502,In_198,In_425);
xor U4503 (N_4503,In_1790,In_954);
nand U4504 (N_4504,In_1559,In_2321);
nor U4505 (N_4505,In_1503,In_888);
and U4506 (N_4506,In_2791,In_2973);
nor U4507 (N_4507,In_961,In_1654);
nor U4508 (N_4508,In_2117,In_1411);
nand U4509 (N_4509,In_2697,In_1848);
and U4510 (N_4510,In_1171,In_729);
nor U4511 (N_4511,In_1721,In_1135);
nand U4512 (N_4512,In_1867,In_2590);
and U4513 (N_4513,In_712,In_386);
or U4514 (N_4514,In_2181,In_1182);
xor U4515 (N_4515,In_100,In_2968);
nor U4516 (N_4516,In_2058,In_1671);
xor U4517 (N_4517,In_2669,In_472);
nor U4518 (N_4518,In_1496,In_892);
and U4519 (N_4519,In_2255,In_2256);
xnor U4520 (N_4520,In_1113,In_493);
nand U4521 (N_4521,In_697,In_1898);
and U4522 (N_4522,In_140,In_1591);
xnor U4523 (N_4523,In_540,In_1030);
and U4524 (N_4524,In_2617,In_1919);
xor U4525 (N_4525,In_2546,In_2296);
and U4526 (N_4526,In_2375,In_2826);
xor U4527 (N_4527,In_460,In_2418);
or U4528 (N_4528,In_2944,In_1787);
and U4529 (N_4529,In_1038,In_1203);
nor U4530 (N_4530,In_757,In_1635);
or U4531 (N_4531,In_2244,In_615);
nor U4532 (N_4532,In_1463,In_233);
nand U4533 (N_4533,In_2587,In_394);
xnor U4534 (N_4534,In_2841,In_2693);
and U4535 (N_4535,In_1878,In_2509);
or U4536 (N_4536,In_182,In_1869);
and U4537 (N_4537,In_327,In_384);
xnor U4538 (N_4538,In_1036,In_2698);
and U4539 (N_4539,In_2500,In_2560);
nor U4540 (N_4540,In_859,In_750);
xnor U4541 (N_4541,In_1938,In_2403);
or U4542 (N_4542,In_330,In_2371);
and U4543 (N_4543,In_2867,In_740);
nand U4544 (N_4544,In_2684,In_2806);
nand U4545 (N_4545,In_2458,In_1284);
and U4546 (N_4546,In_1657,In_2461);
nor U4547 (N_4547,In_871,In_907);
xor U4548 (N_4548,In_1699,In_414);
nand U4549 (N_4549,In_1713,In_1855);
nand U4550 (N_4550,In_1995,In_2902);
or U4551 (N_4551,In_112,In_2622);
and U4552 (N_4552,In_803,In_2648);
or U4553 (N_4553,In_2058,In_377);
or U4554 (N_4554,In_1758,In_1619);
and U4555 (N_4555,In_448,In_625);
and U4556 (N_4556,In_2644,In_2383);
nor U4557 (N_4557,In_1735,In_2361);
and U4558 (N_4558,In_2116,In_2976);
or U4559 (N_4559,In_1389,In_1216);
nand U4560 (N_4560,In_1715,In_199);
and U4561 (N_4561,In_2153,In_406);
or U4562 (N_4562,In_1004,In_293);
nand U4563 (N_4563,In_2340,In_503);
nand U4564 (N_4564,In_1897,In_1498);
or U4565 (N_4565,In_463,In_1714);
nand U4566 (N_4566,In_2894,In_1167);
nand U4567 (N_4567,In_1336,In_219);
and U4568 (N_4568,In_1413,In_2833);
or U4569 (N_4569,In_2088,In_2569);
nand U4570 (N_4570,In_66,In_1993);
or U4571 (N_4571,In_2007,In_1937);
nor U4572 (N_4572,In_2826,In_2910);
nor U4573 (N_4573,In_298,In_1061);
nor U4574 (N_4574,In_2092,In_1963);
xor U4575 (N_4575,In_441,In_2384);
or U4576 (N_4576,In_2714,In_1361);
and U4577 (N_4577,In_2819,In_1332);
xor U4578 (N_4578,In_1515,In_1404);
and U4579 (N_4579,In_1473,In_1660);
nand U4580 (N_4580,In_2566,In_1591);
and U4581 (N_4581,In_359,In_2101);
or U4582 (N_4582,In_189,In_1781);
nand U4583 (N_4583,In_1340,In_1167);
or U4584 (N_4584,In_507,In_2841);
nor U4585 (N_4585,In_450,In_2100);
and U4586 (N_4586,In_1051,In_1801);
nor U4587 (N_4587,In_1030,In_246);
or U4588 (N_4588,In_2338,In_773);
or U4589 (N_4589,In_1575,In_956);
nand U4590 (N_4590,In_1162,In_615);
xor U4591 (N_4591,In_2250,In_1930);
xor U4592 (N_4592,In_1912,In_1019);
nor U4593 (N_4593,In_848,In_1628);
nor U4594 (N_4594,In_2079,In_2157);
xnor U4595 (N_4595,In_88,In_1810);
or U4596 (N_4596,In_1591,In_2762);
nand U4597 (N_4597,In_260,In_1086);
nand U4598 (N_4598,In_2009,In_1030);
or U4599 (N_4599,In_713,In_2524);
and U4600 (N_4600,In_587,In_2530);
and U4601 (N_4601,In_2195,In_395);
or U4602 (N_4602,In_91,In_202);
nand U4603 (N_4603,In_2489,In_2584);
or U4604 (N_4604,In_431,In_2475);
nand U4605 (N_4605,In_2769,In_1491);
nand U4606 (N_4606,In_2823,In_1910);
nor U4607 (N_4607,In_1701,In_2179);
or U4608 (N_4608,In_1934,In_2976);
or U4609 (N_4609,In_1328,In_2862);
nand U4610 (N_4610,In_1270,In_215);
xnor U4611 (N_4611,In_836,In_2382);
nor U4612 (N_4612,In_2072,In_1695);
nand U4613 (N_4613,In_1979,In_952);
nor U4614 (N_4614,In_2604,In_178);
nor U4615 (N_4615,In_662,In_743);
or U4616 (N_4616,In_1165,In_975);
xnor U4617 (N_4617,In_124,In_2782);
and U4618 (N_4618,In_758,In_122);
or U4619 (N_4619,In_1430,In_2655);
nor U4620 (N_4620,In_2026,In_543);
or U4621 (N_4621,In_2164,In_1272);
xor U4622 (N_4622,In_1085,In_232);
nand U4623 (N_4623,In_2194,In_677);
or U4624 (N_4624,In_236,In_1950);
xnor U4625 (N_4625,In_566,In_1156);
or U4626 (N_4626,In_216,In_2336);
xor U4627 (N_4627,In_2825,In_322);
nor U4628 (N_4628,In_1704,In_2053);
and U4629 (N_4629,In_2667,In_1917);
and U4630 (N_4630,In_2669,In_899);
or U4631 (N_4631,In_2638,In_664);
nand U4632 (N_4632,In_952,In_2248);
nor U4633 (N_4633,In_2822,In_1405);
and U4634 (N_4634,In_196,In_2218);
nor U4635 (N_4635,In_980,In_1813);
nand U4636 (N_4636,In_2865,In_383);
xnor U4637 (N_4637,In_2495,In_2224);
xnor U4638 (N_4638,In_1302,In_1055);
and U4639 (N_4639,In_876,In_1040);
and U4640 (N_4640,In_240,In_2160);
xnor U4641 (N_4641,In_1933,In_1918);
or U4642 (N_4642,In_778,In_2304);
xor U4643 (N_4643,In_1759,In_2739);
or U4644 (N_4644,In_488,In_2023);
xor U4645 (N_4645,In_1076,In_2456);
nand U4646 (N_4646,In_2601,In_2679);
nand U4647 (N_4647,In_121,In_2152);
and U4648 (N_4648,In_1132,In_2091);
nand U4649 (N_4649,In_1072,In_1519);
nor U4650 (N_4650,In_2614,In_1420);
or U4651 (N_4651,In_2607,In_2806);
or U4652 (N_4652,In_683,In_174);
nand U4653 (N_4653,In_569,In_485);
nand U4654 (N_4654,In_437,In_1947);
and U4655 (N_4655,In_2439,In_2474);
or U4656 (N_4656,In_2664,In_1448);
xnor U4657 (N_4657,In_2600,In_1361);
or U4658 (N_4658,In_2911,In_896);
or U4659 (N_4659,In_631,In_225);
nor U4660 (N_4660,In_656,In_1721);
or U4661 (N_4661,In_2402,In_1230);
nand U4662 (N_4662,In_253,In_82);
xnor U4663 (N_4663,In_2606,In_1771);
xor U4664 (N_4664,In_2806,In_2222);
nand U4665 (N_4665,In_2974,In_2835);
nand U4666 (N_4666,In_2551,In_877);
nor U4667 (N_4667,In_2587,In_1291);
nand U4668 (N_4668,In_38,In_421);
or U4669 (N_4669,In_1169,In_2054);
nand U4670 (N_4670,In_703,In_2861);
or U4671 (N_4671,In_1069,In_1830);
nand U4672 (N_4672,In_840,In_640);
or U4673 (N_4673,In_1717,In_1338);
xor U4674 (N_4674,In_2504,In_2597);
and U4675 (N_4675,In_298,In_2747);
and U4676 (N_4676,In_2701,In_868);
nand U4677 (N_4677,In_223,In_869);
and U4678 (N_4678,In_2983,In_2575);
nor U4679 (N_4679,In_1717,In_2371);
xnor U4680 (N_4680,In_512,In_2504);
nor U4681 (N_4681,In_2828,In_206);
and U4682 (N_4682,In_890,In_1210);
nand U4683 (N_4683,In_2175,In_236);
and U4684 (N_4684,In_2914,In_2100);
nor U4685 (N_4685,In_2628,In_681);
nor U4686 (N_4686,In_1334,In_1451);
nand U4687 (N_4687,In_2002,In_1997);
nor U4688 (N_4688,In_774,In_1064);
nor U4689 (N_4689,In_1111,In_1626);
nor U4690 (N_4690,In_1989,In_2795);
or U4691 (N_4691,In_1604,In_1846);
or U4692 (N_4692,In_256,In_479);
or U4693 (N_4693,In_200,In_2028);
or U4694 (N_4694,In_175,In_875);
nand U4695 (N_4695,In_624,In_1905);
and U4696 (N_4696,In_1669,In_43);
or U4697 (N_4697,In_1816,In_2653);
nor U4698 (N_4698,In_1837,In_1123);
xnor U4699 (N_4699,In_713,In_419);
and U4700 (N_4700,In_2150,In_2460);
nand U4701 (N_4701,In_2087,In_669);
nand U4702 (N_4702,In_2891,In_1184);
and U4703 (N_4703,In_2165,In_2944);
and U4704 (N_4704,In_1307,In_2805);
xor U4705 (N_4705,In_2055,In_1027);
nor U4706 (N_4706,In_2063,In_1236);
nand U4707 (N_4707,In_2406,In_925);
or U4708 (N_4708,In_324,In_1361);
nand U4709 (N_4709,In_2264,In_1319);
xor U4710 (N_4710,In_2097,In_823);
nor U4711 (N_4711,In_827,In_401);
and U4712 (N_4712,In_1327,In_2101);
xor U4713 (N_4713,In_1183,In_2695);
nand U4714 (N_4714,In_715,In_147);
xnor U4715 (N_4715,In_1135,In_803);
and U4716 (N_4716,In_2762,In_2633);
nand U4717 (N_4717,In_2875,In_156);
nand U4718 (N_4718,In_1268,In_573);
or U4719 (N_4719,In_1854,In_97);
xnor U4720 (N_4720,In_1756,In_2119);
and U4721 (N_4721,In_1804,In_843);
xor U4722 (N_4722,In_1845,In_461);
or U4723 (N_4723,In_1679,In_1207);
or U4724 (N_4724,In_973,In_630);
nor U4725 (N_4725,In_1057,In_487);
xor U4726 (N_4726,In_831,In_1643);
nand U4727 (N_4727,In_1938,In_2364);
xnor U4728 (N_4728,In_930,In_808);
xor U4729 (N_4729,In_2546,In_825);
and U4730 (N_4730,In_1685,In_1084);
or U4731 (N_4731,In_2392,In_1044);
xor U4732 (N_4732,In_1550,In_2504);
nand U4733 (N_4733,In_381,In_1194);
xor U4734 (N_4734,In_2665,In_1144);
nor U4735 (N_4735,In_1836,In_74);
and U4736 (N_4736,In_1052,In_2852);
and U4737 (N_4737,In_2639,In_2526);
nand U4738 (N_4738,In_139,In_735);
nand U4739 (N_4739,In_547,In_2075);
and U4740 (N_4740,In_1317,In_1159);
or U4741 (N_4741,In_18,In_2189);
nor U4742 (N_4742,In_889,In_308);
xor U4743 (N_4743,In_722,In_1648);
or U4744 (N_4744,In_1429,In_653);
xnor U4745 (N_4745,In_1374,In_2315);
or U4746 (N_4746,In_511,In_2254);
or U4747 (N_4747,In_2537,In_266);
nor U4748 (N_4748,In_1590,In_2064);
and U4749 (N_4749,In_1756,In_792);
or U4750 (N_4750,In_22,In_1210);
and U4751 (N_4751,In_2154,In_858);
nor U4752 (N_4752,In_309,In_1278);
nand U4753 (N_4753,In_2513,In_2953);
nand U4754 (N_4754,In_240,In_1244);
or U4755 (N_4755,In_1328,In_1061);
nor U4756 (N_4756,In_2424,In_2278);
nand U4757 (N_4757,In_627,In_2379);
or U4758 (N_4758,In_2925,In_2093);
nand U4759 (N_4759,In_1526,In_2610);
and U4760 (N_4760,In_588,In_2288);
xor U4761 (N_4761,In_2761,In_1889);
xnor U4762 (N_4762,In_1557,In_939);
nand U4763 (N_4763,In_752,In_272);
xnor U4764 (N_4764,In_306,In_2371);
nand U4765 (N_4765,In_142,In_1533);
or U4766 (N_4766,In_596,In_2377);
xor U4767 (N_4767,In_2179,In_1547);
or U4768 (N_4768,In_618,In_1166);
or U4769 (N_4769,In_2815,In_2241);
xnor U4770 (N_4770,In_1137,In_2433);
xnor U4771 (N_4771,In_1996,In_1598);
nand U4772 (N_4772,In_1574,In_1384);
nand U4773 (N_4773,In_2846,In_236);
or U4774 (N_4774,In_854,In_1130);
and U4775 (N_4775,In_1083,In_2737);
xnor U4776 (N_4776,In_1569,In_1576);
nand U4777 (N_4777,In_901,In_1981);
xnor U4778 (N_4778,In_1236,In_201);
and U4779 (N_4779,In_1669,In_1678);
or U4780 (N_4780,In_2120,In_121);
and U4781 (N_4781,In_2880,In_1986);
xnor U4782 (N_4782,In_2144,In_1386);
xor U4783 (N_4783,In_2666,In_1109);
and U4784 (N_4784,In_119,In_2334);
and U4785 (N_4785,In_2230,In_1858);
nor U4786 (N_4786,In_543,In_1361);
xor U4787 (N_4787,In_322,In_1987);
nand U4788 (N_4788,In_432,In_666);
or U4789 (N_4789,In_2148,In_1157);
xor U4790 (N_4790,In_400,In_1806);
nor U4791 (N_4791,In_2856,In_1571);
or U4792 (N_4792,In_2067,In_2022);
xor U4793 (N_4793,In_2177,In_841);
nor U4794 (N_4794,In_2220,In_1604);
or U4795 (N_4795,In_1671,In_705);
and U4796 (N_4796,In_2133,In_289);
nor U4797 (N_4797,In_544,In_2738);
nor U4798 (N_4798,In_2231,In_1130);
and U4799 (N_4799,In_2772,In_1153);
nand U4800 (N_4800,In_2084,In_2215);
nand U4801 (N_4801,In_2994,In_1015);
and U4802 (N_4802,In_810,In_2966);
and U4803 (N_4803,In_144,In_1712);
nor U4804 (N_4804,In_2564,In_2420);
or U4805 (N_4805,In_279,In_2164);
nand U4806 (N_4806,In_1254,In_747);
nand U4807 (N_4807,In_2696,In_1166);
and U4808 (N_4808,In_2223,In_416);
xnor U4809 (N_4809,In_1621,In_932);
nand U4810 (N_4810,In_654,In_1029);
nand U4811 (N_4811,In_1343,In_1821);
or U4812 (N_4812,In_700,In_1164);
or U4813 (N_4813,In_704,In_2432);
nor U4814 (N_4814,In_332,In_104);
xnor U4815 (N_4815,In_219,In_2846);
nand U4816 (N_4816,In_209,In_36);
xnor U4817 (N_4817,In_1907,In_2460);
or U4818 (N_4818,In_489,In_1489);
or U4819 (N_4819,In_253,In_1402);
and U4820 (N_4820,In_271,In_774);
xnor U4821 (N_4821,In_1480,In_1642);
xor U4822 (N_4822,In_1285,In_1239);
nor U4823 (N_4823,In_2918,In_1175);
xor U4824 (N_4824,In_2989,In_2079);
nor U4825 (N_4825,In_1907,In_319);
xor U4826 (N_4826,In_1354,In_661);
or U4827 (N_4827,In_1219,In_1090);
and U4828 (N_4828,In_1061,In_1192);
nor U4829 (N_4829,In_491,In_2280);
and U4830 (N_4830,In_2567,In_2239);
nand U4831 (N_4831,In_658,In_2215);
or U4832 (N_4832,In_2615,In_1241);
xor U4833 (N_4833,In_1498,In_1647);
nand U4834 (N_4834,In_2197,In_1897);
nand U4835 (N_4835,In_2538,In_2843);
and U4836 (N_4836,In_762,In_972);
and U4837 (N_4837,In_871,In_482);
xor U4838 (N_4838,In_1420,In_2529);
xnor U4839 (N_4839,In_2573,In_432);
nor U4840 (N_4840,In_142,In_2024);
or U4841 (N_4841,In_248,In_1798);
nand U4842 (N_4842,In_1339,In_2663);
xor U4843 (N_4843,In_2807,In_1254);
and U4844 (N_4844,In_729,In_2788);
nor U4845 (N_4845,In_1225,In_191);
or U4846 (N_4846,In_345,In_2582);
nand U4847 (N_4847,In_2333,In_576);
nor U4848 (N_4848,In_2766,In_1910);
nand U4849 (N_4849,In_923,In_1357);
xor U4850 (N_4850,In_1318,In_22);
nor U4851 (N_4851,In_2095,In_825);
xnor U4852 (N_4852,In_1137,In_213);
or U4853 (N_4853,In_1497,In_2591);
or U4854 (N_4854,In_2489,In_1673);
xnor U4855 (N_4855,In_616,In_1069);
or U4856 (N_4856,In_2201,In_2034);
xor U4857 (N_4857,In_1177,In_815);
nor U4858 (N_4858,In_2755,In_1657);
and U4859 (N_4859,In_1179,In_1168);
or U4860 (N_4860,In_53,In_201);
nand U4861 (N_4861,In_216,In_317);
xnor U4862 (N_4862,In_2352,In_1352);
nand U4863 (N_4863,In_498,In_930);
and U4864 (N_4864,In_1939,In_265);
or U4865 (N_4865,In_2189,In_2183);
xor U4866 (N_4866,In_1480,In_1148);
nand U4867 (N_4867,In_70,In_2675);
nor U4868 (N_4868,In_2142,In_832);
xor U4869 (N_4869,In_1608,In_1771);
nor U4870 (N_4870,In_56,In_1124);
or U4871 (N_4871,In_836,In_2286);
nor U4872 (N_4872,In_665,In_580);
nand U4873 (N_4873,In_727,In_995);
nand U4874 (N_4874,In_888,In_1353);
nor U4875 (N_4875,In_1375,In_1964);
nand U4876 (N_4876,In_581,In_2886);
nand U4877 (N_4877,In_2220,In_222);
xnor U4878 (N_4878,In_1984,In_532);
or U4879 (N_4879,In_2449,In_530);
and U4880 (N_4880,In_1981,In_730);
xnor U4881 (N_4881,In_2665,In_3);
or U4882 (N_4882,In_1550,In_2362);
xnor U4883 (N_4883,In_2220,In_2042);
xnor U4884 (N_4884,In_578,In_2);
xnor U4885 (N_4885,In_1383,In_1682);
and U4886 (N_4886,In_251,In_989);
and U4887 (N_4887,In_1406,In_765);
nand U4888 (N_4888,In_1286,In_2573);
xor U4889 (N_4889,In_1971,In_1221);
and U4890 (N_4890,In_2996,In_621);
and U4891 (N_4891,In_19,In_2887);
or U4892 (N_4892,In_2166,In_2821);
nand U4893 (N_4893,In_1173,In_2337);
xor U4894 (N_4894,In_2857,In_2910);
nand U4895 (N_4895,In_1505,In_2173);
and U4896 (N_4896,In_1808,In_788);
and U4897 (N_4897,In_2221,In_1385);
xor U4898 (N_4898,In_2402,In_607);
nand U4899 (N_4899,In_2006,In_1668);
or U4900 (N_4900,In_2525,In_970);
nand U4901 (N_4901,In_1872,In_1563);
nand U4902 (N_4902,In_1444,In_2400);
and U4903 (N_4903,In_2175,In_2690);
nand U4904 (N_4904,In_1313,In_1631);
nor U4905 (N_4905,In_1751,In_248);
xnor U4906 (N_4906,In_1436,In_2353);
nor U4907 (N_4907,In_915,In_2780);
and U4908 (N_4908,In_522,In_2087);
and U4909 (N_4909,In_390,In_187);
and U4910 (N_4910,In_2179,In_544);
nand U4911 (N_4911,In_1960,In_557);
nor U4912 (N_4912,In_1244,In_327);
or U4913 (N_4913,In_455,In_2676);
xor U4914 (N_4914,In_1970,In_288);
nand U4915 (N_4915,In_2982,In_220);
and U4916 (N_4916,In_1211,In_483);
nand U4917 (N_4917,In_1859,In_883);
nor U4918 (N_4918,In_548,In_1638);
xor U4919 (N_4919,In_240,In_2900);
nor U4920 (N_4920,In_2237,In_273);
nor U4921 (N_4921,In_1993,In_923);
nor U4922 (N_4922,In_1344,In_50);
nor U4923 (N_4923,In_460,In_1033);
xor U4924 (N_4924,In_1307,In_226);
nor U4925 (N_4925,In_257,In_2291);
nand U4926 (N_4926,In_1301,In_1835);
xnor U4927 (N_4927,In_1418,In_2892);
and U4928 (N_4928,In_2938,In_2482);
nor U4929 (N_4929,In_217,In_2500);
and U4930 (N_4930,In_2381,In_1364);
and U4931 (N_4931,In_1854,In_2040);
and U4932 (N_4932,In_2269,In_1835);
xor U4933 (N_4933,In_594,In_2590);
xor U4934 (N_4934,In_1031,In_1606);
nor U4935 (N_4935,In_50,In_1637);
xor U4936 (N_4936,In_1154,In_1419);
and U4937 (N_4937,In_1583,In_796);
xor U4938 (N_4938,In_375,In_2481);
nand U4939 (N_4939,In_2493,In_374);
or U4940 (N_4940,In_2803,In_1240);
and U4941 (N_4941,In_771,In_2178);
and U4942 (N_4942,In_1722,In_1452);
nand U4943 (N_4943,In_774,In_905);
xor U4944 (N_4944,In_34,In_1538);
nor U4945 (N_4945,In_1233,In_2675);
and U4946 (N_4946,In_2759,In_2548);
or U4947 (N_4947,In_259,In_21);
or U4948 (N_4948,In_85,In_652);
and U4949 (N_4949,In_1216,In_2248);
nor U4950 (N_4950,In_2761,In_2561);
nor U4951 (N_4951,In_398,In_1067);
or U4952 (N_4952,In_2518,In_2041);
or U4953 (N_4953,In_387,In_2795);
nand U4954 (N_4954,In_242,In_909);
and U4955 (N_4955,In_790,In_1785);
nand U4956 (N_4956,In_1665,In_2664);
xnor U4957 (N_4957,In_2753,In_85);
xor U4958 (N_4958,In_762,In_2053);
and U4959 (N_4959,In_1373,In_1425);
or U4960 (N_4960,In_1770,In_1445);
nor U4961 (N_4961,In_1161,In_555);
nor U4962 (N_4962,In_1512,In_850);
or U4963 (N_4963,In_2856,In_2973);
nor U4964 (N_4964,In_2820,In_966);
and U4965 (N_4965,In_1593,In_217);
nor U4966 (N_4966,In_210,In_1157);
or U4967 (N_4967,In_2730,In_639);
xnor U4968 (N_4968,In_219,In_1634);
and U4969 (N_4969,In_171,In_2457);
and U4970 (N_4970,In_438,In_2496);
nand U4971 (N_4971,In_2570,In_757);
and U4972 (N_4972,In_1904,In_1122);
xnor U4973 (N_4973,In_657,In_2542);
xnor U4974 (N_4974,In_2659,In_471);
and U4975 (N_4975,In_1549,In_2179);
nor U4976 (N_4976,In_858,In_970);
nor U4977 (N_4977,In_1847,In_1894);
xnor U4978 (N_4978,In_1901,In_2549);
xnor U4979 (N_4979,In_1674,In_1234);
or U4980 (N_4980,In_2638,In_2848);
xnor U4981 (N_4981,In_533,In_2086);
or U4982 (N_4982,In_2803,In_1839);
nand U4983 (N_4983,In_1999,In_2210);
xnor U4984 (N_4984,In_2797,In_878);
or U4985 (N_4985,In_742,In_80);
xnor U4986 (N_4986,In_2230,In_182);
nor U4987 (N_4987,In_2302,In_1859);
xnor U4988 (N_4988,In_531,In_2233);
nand U4989 (N_4989,In_2833,In_813);
and U4990 (N_4990,In_2345,In_2877);
nor U4991 (N_4991,In_2560,In_1962);
nor U4992 (N_4992,In_2018,In_2455);
or U4993 (N_4993,In_1148,In_608);
and U4994 (N_4994,In_1096,In_2585);
and U4995 (N_4995,In_1988,In_2494);
nor U4996 (N_4996,In_644,In_1722);
or U4997 (N_4997,In_1836,In_2411);
nor U4998 (N_4998,In_714,In_1728);
and U4999 (N_4999,In_441,In_1781);
xnor U5000 (N_5000,In_2546,In_689);
and U5001 (N_5001,In_2221,In_940);
nand U5002 (N_5002,In_2741,In_68);
or U5003 (N_5003,In_1286,In_922);
nor U5004 (N_5004,In_729,In_318);
nor U5005 (N_5005,In_413,In_1656);
or U5006 (N_5006,In_1398,In_2940);
or U5007 (N_5007,In_1705,In_1861);
or U5008 (N_5008,In_1286,In_2200);
nand U5009 (N_5009,In_2875,In_1582);
or U5010 (N_5010,In_1242,In_1208);
nand U5011 (N_5011,In_2619,In_2160);
nand U5012 (N_5012,In_2539,In_599);
and U5013 (N_5013,In_1761,In_1658);
xnor U5014 (N_5014,In_2326,In_1407);
or U5015 (N_5015,In_2846,In_850);
and U5016 (N_5016,In_1897,In_1583);
and U5017 (N_5017,In_2459,In_872);
or U5018 (N_5018,In_922,In_627);
or U5019 (N_5019,In_1720,In_601);
or U5020 (N_5020,In_2215,In_1279);
xnor U5021 (N_5021,In_1698,In_1795);
nand U5022 (N_5022,In_1231,In_1230);
or U5023 (N_5023,In_1488,In_962);
or U5024 (N_5024,In_2038,In_1251);
and U5025 (N_5025,In_394,In_1906);
xnor U5026 (N_5026,In_2920,In_223);
or U5027 (N_5027,In_2215,In_1355);
nor U5028 (N_5028,In_2326,In_2003);
nand U5029 (N_5029,In_2566,In_2479);
nor U5030 (N_5030,In_636,In_537);
xor U5031 (N_5031,In_516,In_1580);
and U5032 (N_5032,In_331,In_86);
or U5033 (N_5033,In_1630,In_2945);
or U5034 (N_5034,In_1683,In_1263);
xnor U5035 (N_5035,In_53,In_2564);
or U5036 (N_5036,In_1641,In_1825);
nand U5037 (N_5037,In_620,In_1193);
nor U5038 (N_5038,In_495,In_1968);
nor U5039 (N_5039,In_2125,In_190);
or U5040 (N_5040,In_52,In_1318);
and U5041 (N_5041,In_1161,In_309);
or U5042 (N_5042,In_979,In_1904);
xnor U5043 (N_5043,In_256,In_1735);
and U5044 (N_5044,In_484,In_1438);
nor U5045 (N_5045,In_660,In_2752);
or U5046 (N_5046,In_623,In_1920);
or U5047 (N_5047,In_2954,In_2259);
nor U5048 (N_5048,In_1188,In_997);
xor U5049 (N_5049,In_2923,In_1971);
xnor U5050 (N_5050,In_1287,In_770);
nor U5051 (N_5051,In_2753,In_1945);
and U5052 (N_5052,In_1273,In_724);
xnor U5053 (N_5053,In_567,In_2068);
nand U5054 (N_5054,In_1906,In_2474);
nand U5055 (N_5055,In_1832,In_1335);
and U5056 (N_5056,In_310,In_1708);
nor U5057 (N_5057,In_2457,In_1505);
xor U5058 (N_5058,In_1061,In_1565);
and U5059 (N_5059,In_481,In_2166);
and U5060 (N_5060,In_2022,In_2395);
and U5061 (N_5061,In_929,In_1759);
nor U5062 (N_5062,In_1655,In_1267);
nor U5063 (N_5063,In_2927,In_1136);
and U5064 (N_5064,In_2096,In_2333);
or U5065 (N_5065,In_2785,In_2188);
nor U5066 (N_5066,In_2390,In_65);
nor U5067 (N_5067,In_1992,In_572);
nand U5068 (N_5068,In_1207,In_2995);
xnor U5069 (N_5069,In_457,In_2295);
xor U5070 (N_5070,In_920,In_326);
nand U5071 (N_5071,In_799,In_628);
nand U5072 (N_5072,In_2431,In_100);
and U5073 (N_5073,In_618,In_98);
xnor U5074 (N_5074,In_679,In_2886);
and U5075 (N_5075,In_609,In_572);
nand U5076 (N_5076,In_474,In_552);
or U5077 (N_5077,In_1002,In_164);
nand U5078 (N_5078,In_285,In_2693);
xor U5079 (N_5079,In_1593,In_890);
xor U5080 (N_5080,In_1666,In_1210);
xor U5081 (N_5081,In_2287,In_1389);
and U5082 (N_5082,In_2219,In_1133);
xor U5083 (N_5083,In_2393,In_582);
or U5084 (N_5084,In_487,In_479);
xor U5085 (N_5085,In_2413,In_320);
nand U5086 (N_5086,In_1336,In_1614);
nor U5087 (N_5087,In_632,In_479);
nor U5088 (N_5088,In_2671,In_1323);
nor U5089 (N_5089,In_458,In_2286);
or U5090 (N_5090,In_2664,In_2501);
nor U5091 (N_5091,In_494,In_1804);
and U5092 (N_5092,In_70,In_1188);
xnor U5093 (N_5093,In_2948,In_2001);
nand U5094 (N_5094,In_1842,In_1362);
nor U5095 (N_5095,In_1336,In_1702);
nand U5096 (N_5096,In_2016,In_1435);
nor U5097 (N_5097,In_1413,In_1309);
nor U5098 (N_5098,In_1477,In_2047);
nor U5099 (N_5099,In_482,In_1724);
or U5100 (N_5100,In_2563,In_656);
and U5101 (N_5101,In_2974,In_2282);
or U5102 (N_5102,In_2125,In_1349);
and U5103 (N_5103,In_1042,In_1123);
nand U5104 (N_5104,In_633,In_2210);
and U5105 (N_5105,In_2600,In_1125);
or U5106 (N_5106,In_1570,In_1229);
and U5107 (N_5107,In_529,In_1345);
nor U5108 (N_5108,In_404,In_1130);
nand U5109 (N_5109,In_2034,In_518);
xor U5110 (N_5110,In_2529,In_1344);
or U5111 (N_5111,In_412,In_2543);
or U5112 (N_5112,In_1937,In_64);
and U5113 (N_5113,In_1299,In_2623);
and U5114 (N_5114,In_1982,In_1441);
or U5115 (N_5115,In_583,In_367);
or U5116 (N_5116,In_721,In_1026);
and U5117 (N_5117,In_1475,In_127);
and U5118 (N_5118,In_2185,In_55);
or U5119 (N_5119,In_1812,In_1795);
or U5120 (N_5120,In_724,In_1087);
or U5121 (N_5121,In_2828,In_455);
and U5122 (N_5122,In_605,In_342);
xnor U5123 (N_5123,In_1186,In_1085);
nand U5124 (N_5124,In_2833,In_1926);
and U5125 (N_5125,In_1529,In_853);
xnor U5126 (N_5126,In_465,In_1527);
or U5127 (N_5127,In_2164,In_1016);
or U5128 (N_5128,In_340,In_1286);
xor U5129 (N_5129,In_1155,In_1416);
nand U5130 (N_5130,In_1029,In_1247);
and U5131 (N_5131,In_2093,In_2003);
and U5132 (N_5132,In_2504,In_254);
nand U5133 (N_5133,In_2177,In_823);
nand U5134 (N_5134,In_58,In_1939);
and U5135 (N_5135,In_2643,In_2060);
nand U5136 (N_5136,In_2855,In_1874);
nor U5137 (N_5137,In_213,In_1367);
xnor U5138 (N_5138,In_958,In_2795);
nor U5139 (N_5139,In_890,In_2272);
or U5140 (N_5140,In_2654,In_508);
and U5141 (N_5141,In_891,In_1538);
or U5142 (N_5142,In_2046,In_181);
or U5143 (N_5143,In_2134,In_2939);
nor U5144 (N_5144,In_187,In_516);
nand U5145 (N_5145,In_1133,In_1199);
and U5146 (N_5146,In_254,In_1088);
and U5147 (N_5147,In_2071,In_402);
nor U5148 (N_5148,In_137,In_2979);
nand U5149 (N_5149,In_1308,In_444);
or U5150 (N_5150,In_1023,In_974);
xnor U5151 (N_5151,In_1104,In_824);
and U5152 (N_5152,In_2418,In_1342);
or U5153 (N_5153,In_2323,In_1545);
nor U5154 (N_5154,In_2545,In_2186);
and U5155 (N_5155,In_2601,In_477);
nor U5156 (N_5156,In_1909,In_1990);
nand U5157 (N_5157,In_1193,In_1211);
xor U5158 (N_5158,In_1058,In_381);
or U5159 (N_5159,In_1999,In_206);
nor U5160 (N_5160,In_448,In_882);
xnor U5161 (N_5161,In_1766,In_1600);
nor U5162 (N_5162,In_2166,In_2441);
xnor U5163 (N_5163,In_1487,In_1809);
and U5164 (N_5164,In_2513,In_1251);
and U5165 (N_5165,In_969,In_947);
and U5166 (N_5166,In_1646,In_468);
nor U5167 (N_5167,In_2238,In_365);
and U5168 (N_5168,In_87,In_349);
nand U5169 (N_5169,In_735,In_1826);
and U5170 (N_5170,In_32,In_1694);
nand U5171 (N_5171,In_2730,In_2662);
nor U5172 (N_5172,In_380,In_2584);
nor U5173 (N_5173,In_1930,In_1230);
nor U5174 (N_5174,In_741,In_72);
nand U5175 (N_5175,In_1217,In_1036);
xor U5176 (N_5176,In_1644,In_1415);
or U5177 (N_5177,In_1512,In_110);
nor U5178 (N_5178,In_2562,In_2644);
or U5179 (N_5179,In_2964,In_328);
nor U5180 (N_5180,In_1740,In_910);
nand U5181 (N_5181,In_513,In_832);
xor U5182 (N_5182,In_1585,In_913);
nor U5183 (N_5183,In_2460,In_2552);
xor U5184 (N_5184,In_181,In_577);
nand U5185 (N_5185,In_583,In_2022);
xnor U5186 (N_5186,In_2471,In_1031);
or U5187 (N_5187,In_2240,In_2415);
xor U5188 (N_5188,In_881,In_1442);
nand U5189 (N_5189,In_915,In_1356);
nor U5190 (N_5190,In_1879,In_2740);
and U5191 (N_5191,In_320,In_1853);
or U5192 (N_5192,In_636,In_1185);
xor U5193 (N_5193,In_1153,In_2823);
or U5194 (N_5194,In_1393,In_1509);
nand U5195 (N_5195,In_1187,In_1409);
and U5196 (N_5196,In_1697,In_645);
and U5197 (N_5197,In_21,In_300);
xnor U5198 (N_5198,In_1637,In_1259);
or U5199 (N_5199,In_2695,In_2740);
and U5200 (N_5200,In_50,In_2790);
nor U5201 (N_5201,In_2478,In_1761);
nor U5202 (N_5202,In_2901,In_400);
nand U5203 (N_5203,In_2187,In_190);
and U5204 (N_5204,In_1150,In_1892);
and U5205 (N_5205,In_2398,In_1024);
xor U5206 (N_5206,In_387,In_2123);
and U5207 (N_5207,In_2361,In_1408);
nor U5208 (N_5208,In_1225,In_1163);
and U5209 (N_5209,In_2255,In_1617);
nand U5210 (N_5210,In_2792,In_2434);
xnor U5211 (N_5211,In_426,In_1766);
or U5212 (N_5212,In_1438,In_1138);
xnor U5213 (N_5213,In_1517,In_2429);
xor U5214 (N_5214,In_1541,In_1190);
nor U5215 (N_5215,In_2334,In_1575);
and U5216 (N_5216,In_2935,In_989);
or U5217 (N_5217,In_1738,In_1895);
nor U5218 (N_5218,In_668,In_50);
nand U5219 (N_5219,In_363,In_1521);
and U5220 (N_5220,In_437,In_168);
xnor U5221 (N_5221,In_2934,In_549);
and U5222 (N_5222,In_2227,In_1460);
nor U5223 (N_5223,In_2240,In_37);
nand U5224 (N_5224,In_2123,In_568);
nand U5225 (N_5225,In_2683,In_2546);
xor U5226 (N_5226,In_723,In_863);
or U5227 (N_5227,In_2393,In_392);
nor U5228 (N_5228,In_2643,In_2814);
xnor U5229 (N_5229,In_2695,In_2486);
nand U5230 (N_5230,In_2504,In_957);
nand U5231 (N_5231,In_1044,In_667);
nor U5232 (N_5232,In_1523,In_663);
nor U5233 (N_5233,In_401,In_2166);
nand U5234 (N_5234,In_1734,In_985);
and U5235 (N_5235,In_1998,In_2029);
or U5236 (N_5236,In_2013,In_2051);
xor U5237 (N_5237,In_1307,In_2965);
nor U5238 (N_5238,In_696,In_567);
or U5239 (N_5239,In_704,In_750);
xnor U5240 (N_5240,In_537,In_2245);
or U5241 (N_5241,In_131,In_2036);
nor U5242 (N_5242,In_2076,In_1300);
and U5243 (N_5243,In_1368,In_1440);
or U5244 (N_5244,In_614,In_2659);
nand U5245 (N_5245,In_1607,In_546);
xnor U5246 (N_5246,In_2748,In_2926);
or U5247 (N_5247,In_1407,In_959);
nand U5248 (N_5248,In_622,In_2024);
and U5249 (N_5249,In_2802,In_1770);
nand U5250 (N_5250,In_1746,In_118);
nand U5251 (N_5251,In_25,In_2015);
nand U5252 (N_5252,In_836,In_2297);
and U5253 (N_5253,In_1640,In_74);
or U5254 (N_5254,In_1991,In_804);
nor U5255 (N_5255,In_2146,In_2740);
and U5256 (N_5256,In_966,In_860);
or U5257 (N_5257,In_1996,In_1523);
or U5258 (N_5258,In_2989,In_2718);
and U5259 (N_5259,In_2981,In_1505);
and U5260 (N_5260,In_2043,In_202);
nor U5261 (N_5261,In_1477,In_1428);
xor U5262 (N_5262,In_449,In_54);
xor U5263 (N_5263,In_2591,In_2327);
and U5264 (N_5264,In_1078,In_2241);
and U5265 (N_5265,In_797,In_1625);
xnor U5266 (N_5266,In_2733,In_627);
xnor U5267 (N_5267,In_473,In_2937);
or U5268 (N_5268,In_1844,In_2423);
xnor U5269 (N_5269,In_2634,In_211);
nor U5270 (N_5270,In_1996,In_2970);
nor U5271 (N_5271,In_542,In_1809);
nor U5272 (N_5272,In_700,In_606);
nor U5273 (N_5273,In_245,In_2184);
nor U5274 (N_5274,In_267,In_2346);
or U5275 (N_5275,In_192,In_1557);
and U5276 (N_5276,In_1144,In_1375);
nor U5277 (N_5277,In_607,In_789);
nor U5278 (N_5278,In_236,In_201);
and U5279 (N_5279,In_2707,In_1214);
nand U5280 (N_5280,In_2322,In_2921);
nand U5281 (N_5281,In_659,In_2262);
nand U5282 (N_5282,In_2537,In_1573);
or U5283 (N_5283,In_1148,In_148);
nor U5284 (N_5284,In_2359,In_1232);
xor U5285 (N_5285,In_487,In_1009);
or U5286 (N_5286,In_49,In_2396);
nand U5287 (N_5287,In_621,In_1341);
nor U5288 (N_5288,In_2310,In_2926);
or U5289 (N_5289,In_2004,In_1673);
xnor U5290 (N_5290,In_2753,In_1795);
and U5291 (N_5291,In_2624,In_928);
nand U5292 (N_5292,In_314,In_2026);
nor U5293 (N_5293,In_2752,In_53);
xnor U5294 (N_5294,In_740,In_447);
xnor U5295 (N_5295,In_1969,In_1348);
or U5296 (N_5296,In_806,In_563);
or U5297 (N_5297,In_1650,In_1521);
and U5298 (N_5298,In_2804,In_2647);
nand U5299 (N_5299,In_1662,In_2698);
nor U5300 (N_5300,In_2415,In_887);
or U5301 (N_5301,In_2424,In_2093);
xnor U5302 (N_5302,In_751,In_1656);
or U5303 (N_5303,In_1319,In_2900);
or U5304 (N_5304,In_2964,In_1094);
or U5305 (N_5305,In_1586,In_1587);
or U5306 (N_5306,In_641,In_919);
nand U5307 (N_5307,In_2742,In_1989);
nand U5308 (N_5308,In_2539,In_1177);
or U5309 (N_5309,In_966,In_2696);
nor U5310 (N_5310,In_1735,In_475);
and U5311 (N_5311,In_42,In_69);
or U5312 (N_5312,In_647,In_1087);
nand U5313 (N_5313,In_1234,In_2044);
xor U5314 (N_5314,In_1530,In_2944);
nand U5315 (N_5315,In_1539,In_2201);
xnor U5316 (N_5316,In_1565,In_178);
nor U5317 (N_5317,In_2015,In_2506);
or U5318 (N_5318,In_1063,In_822);
and U5319 (N_5319,In_2036,In_1496);
nor U5320 (N_5320,In_2268,In_517);
xnor U5321 (N_5321,In_2180,In_81);
or U5322 (N_5322,In_2156,In_2160);
nand U5323 (N_5323,In_711,In_1765);
and U5324 (N_5324,In_1047,In_1681);
xor U5325 (N_5325,In_1322,In_1927);
nor U5326 (N_5326,In_583,In_1259);
or U5327 (N_5327,In_2106,In_147);
nor U5328 (N_5328,In_1738,In_15);
or U5329 (N_5329,In_284,In_29);
nand U5330 (N_5330,In_1256,In_1340);
nand U5331 (N_5331,In_1779,In_763);
and U5332 (N_5332,In_830,In_1845);
and U5333 (N_5333,In_930,In_2385);
xnor U5334 (N_5334,In_100,In_2233);
xnor U5335 (N_5335,In_2190,In_1115);
nand U5336 (N_5336,In_1334,In_2483);
nand U5337 (N_5337,In_1111,In_1334);
nor U5338 (N_5338,In_2294,In_459);
and U5339 (N_5339,In_2786,In_1264);
nor U5340 (N_5340,In_668,In_2349);
nor U5341 (N_5341,In_1042,In_1211);
or U5342 (N_5342,In_2916,In_1375);
or U5343 (N_5343,In_2837,In_2624);
nor U5344 (N_5344,In_1169,In_1998);
or U5345 (N_5345,In_1130,In_2007);
and U5346 (N_5346,In_2405,In_1022);
and U5347 (N_5347,In_1157,In_1465);
nand U5348 (N_5348,In_655,In_2960);
nand U5349 (N_5349,In_966,In_637);
or U5350 (N_5350,In_1242,In_2712);
nand U5351 (N_5351,In_282,In_657);
xnor U5352 (N_5352,In_2971,In_2728);
nor U5353 (N_5353,In_2278,In_2175);
or U5354 (N_5354,In_1575,In_1592);
nor U5355 (N_5355,In_1546,In_1589);
and U5356 (N_5356,In_2460,In_2492);
xnor U5357 (N_5357,In_854,In_1190);
or U5358 (N_5358,In_212,In_2677);
nand U5359 (N_5359,In_1287,In_1828);
nand U5360 (N_5360,In_2045,In_1243);
nand U5361 (N_5361,In_142,In_1617);
and U5362 (N_5362,In_1585,In_2846);
xor U5363 (N_5363,In_1594,In_2141);
xor U5364 (N_5364,In_2186,In_2457);
xor U5365 (N_5365,In_1483,In_53);
nor U5366 (N_5366,In_1716,In_2138);
nand U5367 (N_5367,In_266,In_1707);
nor U5368 (N_5368,In_649,In_2272);
nand U5369 (N_5369,In_2708,In_2151);
or U5370 (N_5370,In_1933,In_1914);
or U5371 (N_5371,In_169,In_283);
nand U5372 (N_5372,In_2978,In_2868);
xor U5373 (N_5373,In_313,In_2983);
xor U5374 (N_5374,In_1860,In_1626);
xnor U5375 (N_5375,In_2840,In_2828);
or U5376 (N_5376,In_2257,In_1644);
and U5377 (N_5377,In_582,In_2104);
xor U5378 (N_5378,In_2934,In_925);
and U5379 (N_5379,In_1956,In_2197);
nor U5380 (N_5380,In_1453,In_116);
nand U5381 (N_5381,In_2842,In_2603);
or U5382 (N_5382,In_2237,In_2119);
and U5383 (N_5383,In_1163,In_1160);
xor U5384 (N_5384,In_1631,In_1637);
nand U5385 (N_5385,In_2654,In_2895);
xnor U5386 (N_5386,In_2296,In_444);
and U5387 (N_5387,In_784,In_1831);
xnor U5388 (N_5388,In_2523,In_1644);
or U5389 (N_5389,In_1227,In_2366);
and U5390 (N_5390,In_82,In_951);
and U5391 (N_5391,In_2355,In_1200);
nor U5392 (N_5392,In_2178,In_10);
xor U5393 (N_5393,In_232,In_1050);
or U5394 (N_5394,In_396,In_1061);
nand U5395 (N_5395,In_889,In_1516);
and U5396 (N_5396,In_1892,In_1834);
and U5397 (N_5397,In_12,In_1832);
xor U5398 (N_5398,In_2229,In_617);
and U5399 (N_5399,In_2557,In_83);
nand U5400 (N_5400,In_1473,In_2021);
and U5401 (N_5401,In_240,In_2003);
xnor U5402 (N_5402,In_453,In_1656);
xnor U5403 (N_5403,In_2236,In_2823);
xnor U5404 (N_5404,In_570,In_1795);
nand U5405 (N_5405,In_1819,In_124);
nand U5406 (N_5406,In_731,In_978);
nand U5407 (N_5407,In_618,In_2646);
xor U5408 (N_5408,In_2367,In_1042);
and U5409 (N_5409,In_567,In_1305);
or U5410 (N_5410,In_1350,In_2379);
and U5411 (N_5411,In_2512,In_2834);
and U5412 (N_5412,In_341,In_1562);
xnor U5413 (N_5413,In_782,In_1906);
nand U5414 (N_5414,In_2899,In_1013);
and U5415 (N_5415,In_2452,In_253);
or U5416 (N_5416,In_2245,In_346);
xor U5417 (N_5417,In_2541,In_2822);
nand U5418 (N_5418,In_1935,In_2513);
or U5419 (N_5419,In_458,In_281);
and U5420 (N_5420,In_1689,In_714);
nor U5421 (N_5421,In_2537,In_696);
nand U5422 (N_5422,In_409,In_880);
xnor U5423 (N_5423,In_286,In_2045);
or U5424 (N_5424,In_2095,In_276);
nand U5425 (N_5425,In_2191,In_2322);
and U5426 (N_5426,In_2544,In_2999);
xor U5427 (N_5427,In_96,In_253);
or U5428 (N_5428,In_1272,In_694);
and U5429 (N_5429,In_2024,In_470);
xor U5430 (N_5430,In_972,In_1114);
or U5431 (N_5431,In_2339,In_2341);
xnor U5432 (N_5432,In_34,In_1560);
and U5433 (N_5433,In_1059,In_308);
nor U5434 (N_5434,In_1529,In_470);
nor U5435 (N_5435,In_920,In_124);
nor U5436 (N_5436,In_2115,In_367);
nand U5437 (N_5437,In_2060,In_1657);
nand U5438 (N_5438,In_2493,In_655);
nor U5439 (N_5439,In_992,In_1183);
nand U5440 (N_5440,In_645,In_2602);
or U5441 (N_5441,In_2732,In_1419);
nand U5442 (N_5442,In_2282,In_349);
and U5443 (N_5443,In_784,In_2918);
xnor U5444 (N_5444,In_1573,In_1840);
nand U5445 (N_5445,In_2208,In_41);
or U5446 (N_5446,In_2857,In_915);
nand U5447 (N_5447,In_2747,In_473);
and U5448 (N_5448,In_2496,In_324);
nor U5449 (N_5449,In_2570,In_508);
xor U5450 (N_5450,In_2616,In_2069);
or U5451 (N_5451,In_2972,In_1267);
or U5452 (N_5452,In_1291,In_1661);
and U5453 (N_5453,In_2800,In_1882);
or U5454 (N_5454,In_1264,In_1745);
or U5455 (N_5455,In_2569,In_60);
and U5456 (N_5456,In_1618,In_2610);
and U5457 (N_5457,In_1389,In_2098);
nand U5458 (N_5458,In_504,In_65);
and U5459 (N_5459,In_1141,In_399);
and U5460 (N_5460,In_1658,In_1319);
or U5461 (N_5461,In_2332,In_25);
nor U5462 (N_5462,In_2749,In_2216);
or U5463 (N_5463,In_707,In_32);
xnor U5464 (N_5464,In_1532,In_2463);
and U5465 (N_5465,In_2734,In_866);
nor U5466 (N_5466,In_126,In_537);
xnor U5467 (N_5467,In_495,In_2177);
and U5468 (N_5468,In_1713,In_283);
nor U5469 (N_5469,In_604,In_1531);
and U5470 (N_5470,In_196,In_1610);
or U5471 (N_5471,In_291,In_1462);
nor U5472 (N_5472,In_843,In_2380);
and U5473 (N_5473,In_520,In_735);
nor U5474 (N_5474,In_1936,In_2210);
and U5475 (N_5475,In_1368,In_2165);
or U5476 (N_5476,In_1203,In_204);
nor U5477 (N_5477,In_2110,In_1344);
xnor U5478 (N_5478,In_1442,In_371);
nand U5479 (N_5479,In_1965,In_2956);
or U5480 (N_5480,In_1586,In_1291);
xnor U5481 (N_5481,In_124,In_1598);
nand U5482 (N_5482,In_2324,In_25);
and U5483 (N_5483,In_2403,In_2340);
nor U5484 (N_5484,In_771,In_1431);
or U5485 (N_5485,In_580,In_1214);
nand U5486 (N_5486,In_1261,In_2900);
or U5487 (N_5487,In_2953,In_2023);
nand U5488 (N_5488,In_1293,In_2630);
xnor U5489 (N_5489,In_1012,In_512);
nand U5490 (N_5490,In_1437,In_2051);
xnor U5491 (N_5491,In_107,In_2941);
nor U5492 (N_5492,In_765,In_1213);
nand U5493 (N_5493,In_2444,In_1456);
or U5494 (N_5494,In_1314,In_2578);
and U5495 (N_5495,In_2933,In_816);
nor U5496 (N_5496,In_1391,In_312);
xnor U5497 (N_5497,In_325,In_565);
or U5498 (N_5498,In_1479,In_1509);
or U5499 (N_5499,In_413,In_45);
nand U5500 (N_5500,In_2844,In_2399);
or U5501 (N_5501,In_51,In_644);
and U5502 (N_5502,In_68,In_2453);
nand U5503 (N_5503,In_2651,In_450);
and U5504 (N_5504,In_387,In_2493);
and U5505 (N_5505,In_656,In_1389);
or U5506 (N_5506,In_2338,In_231);
xor U5507 (N_5507,In_1854,In_2338);
or U5508 (N_5508,In_326,In_629);
nor U5509 (N_5509,In_1064,In_2627);
or U5510 (N_5510,In_151,In_2133);
nor U5511 (N_5511,In_760,In_350);
nor U5512 (N_5512,In_807,In_507);
nor U5513 (N_5513,In_1664,In_1308);
and U5514 (N_5514,In_2676,In_98);
or U5515 (N_5515,In_964,In_59);
or U5516 (N_5516,In_1778,In_379);
nor U5517 (N_5517,In_2368,In_1056);
and U5518 (N_5518,In_991,In_279);
nor U5519 (N_5519,In_1538,In_360);
xor U5520 (N_5520,In_1670,In_1673);
and U5521 (N_5521,In_2323,In_1417);
nor U5522 (N_5522,In_11,In_608);
nor U5523 (N_5523,In_1668,In_433);
nor U5524 (N_5524,In_2703,In_1949);
nor U5525 (N_5525,In_2294,In_828);
and U5526 (N_5526,In_2414,In_1367);
nand U5527 (N_5527,In_1434,In_174);
nand U5528 (N_5528,In_2619,In_2804);
nor U5529 (N_5529,In_1567,In_2380);
nor U5530 (N_5530,In_2807,In_109);
nor U5531 (N_5531,In_645,In_2891);
nor U5532 (N_5532,In_1699,In_1629);
xnor U5533 (N_5533,In_1012,In_149);
nand U5534 (N_5534,In_1357,In_1110);
xnor U5535 (N_5535,In_1606,In_1719);
and U5536 (N_5536,In_1288,In_2394);
nand U5537 (N_5537,In_2786,In_352);
nand U5538 (N_5538,In_2234,In_2438);
xor U5539 (N_5539,In_1895,In_1676);
nand U5540 (N_5540,In_119,In_1382);
nand U5541 (N_5541,In_2437,In_1633);
nand U5542 (N_5542,In_1716,In_2393);
and U5543 (N_5543,In_2929,In_2610);
xor U5544 (N_5544,In_2940,In_2923);
nor U5545 (N_5545,In_2567,In_1206);
xnor U5546 (N_5546,In_863,In_1060);
nor U5547 (N_5547,In_2162,In_2673);
xor U5548 (N_5548,In_1038,In_2763);
xor U5549 (N_5549,In_789,In_161);
or U5550 (N_5550,In_2468,In_1552);
xnor U5551 (N_5551,In_2664,In_2386);
nor U5552 (N_5552,In_595,In_928);
nor U5553 (N_5553,In_563,In_437);
or U5554 (N_5554,In_1860,In_1083);
nor U5555 (N_5555,In_1855,In_1552);
xor U5556 (N_5556,In_312,In_221);
nor U5557 (N_5557,In_78,In_1938);
nand U5558 (N_5558,In_2732,In_1329);
or U5559 (N_5559,In_560,In_512);
and U5560 (N_5560,In_534,In_2129);
and U5561 (N_5561,In_1479,In_1241);
xor U5562 (N_5562,In_1390,In_1918);
xnor U5563 (N_5563,In_1311,In_257);
nand U5564 (N_5564,In_711,In_2920);
and U5565 (N_5565,In_2937,In_1961);
and U5566 (N_5566,In_2241,In_1928);
xnor U5567 (N_5567,In_220,In_1692);
and U5568 (N_5568,In_2331,In_392);
xnor U5569 (N_5569,In_2551,In_1348);
nand U5570 (N_5570,In_695,In_1823);
nor U5571 (N_5571,In_137,In_2824);
xor U5572 (N_5572,In_2277,In_1313);
nor U5573 (N_5573,In_1922,In_529);
xnor U5574 (N_5574,In_462,In_497);
nor U5575 (N_5575,In_1653,In_1119);
and U5576 (N_5576,In_175,In_599);
xnor U5577 (N_5577,In_1405,In_1185);
and U5578 (N_5578,In_1742,In_1206);
nand U5579 (N_5579,In_1165,In_2987);
xor U5580 (N_5580,In_2323,In_2391);
xnor U5581 (N_5581,In_2646,In_2185);
nor U5582 (N_5582,In_1519,In_2125);
nor U5583 (N_5583,In_492,In_568);
or U5584 (N_5584,In_114,In_718);
nand U5585 (N_5585,In_1488,In_1397);
nor U5586 (N_5586,In_1425,In_2136);
nor U5587 (N_5587,In_2078,In_1303);
nor U5588 (N_5588,In_1370,In_453);
nand U5589 (N_5589,In_205,In_1350);
xnor U5590 (N_5590,In_2500,In_413);
xnor U5591 (N_5591,In_1515,In_531);
or U5592 (N_5592,In_944,In_2505);
and U5593 (N_5593,In_1382,In_2922);
nand U5594 (N_5594,In_1582,In_1718);
or U5595 (N_5595,In_1963,In_1186);
or U5596 (N_5596,In_1353,In_1716);
nor U5597 (N_5597,In_537,In_180);
nor U5598 (N_5598,In_914,In_31);
nand U5599 (N_5599,In_1325,In_2249);
nand U5600 (N_5600,In_2182,In_545);
nand U5601 (N_5601,In_1023,In_2843);
nand U5602 (N_5602,In_2913,In_975);
xnor U5603 (N_5603,In_2897,In_1221);
xor U5604 (N_5604,In_1807,In_119);
xnor U5605 (N_5605,In_62,In_1591);
nand U5606 (N_5606,In_974,In_2245);
nor U5607 (N_5607,In_474,In_1684);
nor U5608 (N_5608,In_333,In_1471);
or U5609 (N_5609,In_2900,In_2214);
nand U5610 (N_5610,In_2729,In_373);
xor U5611 (N_5611,In_2238,In_208);
and U5612 (N_5612,In_881,In_730);
and U5613 (N_5613,In_2022,In_1435);
nor U5614 (N_5614,In_421,In_1062);
or U5615 (N_5615,In_1171,In_480);
xor U5616 (N_5616,In_1438,In_705);
nor U5617 (N_5617,In_1973,In_2597);
nor U5618 (N_5618,In_2478,In_1978);
nor U5619 (N_5619,In_633,In_2936);
nand U5620 (N_5620,In_2984,In_816);
nor U5621 (N_5621,In_2526,In_1846);
and U5622 (N_5622,In_1790,In_1637);
or U5623 (N_5623,In_591,In_649);
nand U5624 (N_5624,In_1378,In_1168);
xnor U5625 (N_5625,In_2995,In_1518);
nand U5626 (N_5626,In_260,In_1513);
or U5627 (N_5627,In_65,In_2641);
xnor U5628 (N_5628,In_1006,In_1546);
or U5629 (N_5629,In_184,In_267);
and U5630 (N_5630,In_2785,In_977);
nand U5631 (N_5631,In_937,In_1423);
nor U5632 (N_5632,In_1817,In_2919);
xnor U5633 (N_5633,In_119,In_1461);
nor U5634 (N_5634,In_1339,In_2185);
xnor U5635 (N_5635,In_1009,In_2670);
and U5636 (N_5636,In_2444,In_370);
nor U5637 (N_5637,In_39,In_265);
and U5638 (N_5638,In_1027,In_1775);
or U5639 (N_5639,In_1597,In_2056);
xor U5640 (N_5640,In_356,In_1939);
nand U5641 (N_5641,In_2730,In_2115);
xor U5642 (N_5642,In_2882,In_1098);
and U5643 (N_5643,In_312,In_2768);
and U5644 (N_5644,In_1347,In_2821);
nand U5645 (N_5645,In_2694,In_1989);
and U5646 (N_5646,In_2012,In_651);
xor U5647 (N_5647,In_2003,In_523);
or U5648 (N_5648,In_1738,In_2275);
or U5649 (N_5649,In_2753,In_692);
nand U5650 (N_5650,In_2821,In_87);
nor U5651 (N_5651,In_2616,In_1035);
nand U5652 (N_5652,In_2557,In_1928);
nand U5653 (N_5653,In_1091,In_2872);
and U5654 (N_5654,In_2643,In_1960);
nand U5655 (N_5655,In_407,In_1000);
xor U5656 (N_5656,In_2169,In_2264);
xnor U5657 (N_5657,In_2050,In_2744);
nand U5658 (N_5658,In_620,In_2103);
or U5659 (N_5659,In_1666,In_1889);
and U5660 (N_5660,In_2652,In_18);
or U5661 (N_5661,In_338,In_1736);
xor U5662 (N_5662,In_328,In_2719);
xor U5663 (N_5663,In_159,In_1490);
nor U5664 (N_5664,In_2705,In_1681);
or U5665 (N_5665,In_448,In_2906);
nand U5666 (N_5666,In_1709,In_2219);
nand U5667 (N_5667,In_1019,In_390);
or U5668 (N_5668,In_114,In_1864);
and U5669 (N_5669,In_269,In_1722);
or U5670 (N_5670,In_2209,In_1031);
and U5671 (N_5671,In_824,In_1482);
nor U5672 (N_5672,In_1684,In_664);
and U5673 (N_5673,In_1686,In_681);
xnor U5674 (N_5674,In_86,In_177);
nand U5675 (N_5675,In_915,In_2868);
xor U5676 (N_5676,In_2983,In_885);
xor U5677 (N_5677,In_1059,In_1003);
or U5678 (N_5678,In_9,In_1877);
and U5679 (N_5679,In_2713,In_665);
and U5680 (N_5680,In_2958,In_1128);
or U5681 (N_5681,In_2349,In_2847);
nor U5682 (N_5682,In_542,In_1993);
and U5683 (N_5683,In_455,In_315);
xnor U5684 (N_5684,In_624,In_2001);
nor U5685 (N_5685,In_2792,In_851);
xnor U5686 (N_5686,In_1900,In_1434);
and U5687 (N_5687,In_679,In_1222);
nor U5688 (N_5688,In_885,In_1202);
and U5689 (N_5689,In_2078,In_2591);
nor U5690 (N_5690,In_710,In_1818);
or U5691 (N_5691,In_1009,In_73);
xnor U5692 (N_5692,In_1778,In_952);
and U5693 (N_5693,In_2430,In_883);
nand U5694 (N_5694,In_2586,In_89);
and U5695 (N_5695,In_31,In_1693);
and U5696 (N_5696,In_2332,In_783);
or U5697 (N_5697,In_1170,In_867);
nand U5698 (N_5698,In_2808,In_2791);
nand U5699 (N_5699,In_1406,In_1498);
xor U5700 (N_5700,In_1266,In_2435);
and U5701 (N_5701,In_327,In_1178);
xnor U5702 (N_5702,In_754,In_256);
nor U5703 (N_5703,In_2846,In_1029);
xnor U5704 (N_5704,In_1962,In_1592);
xnor U5705 (N_5705,In_1030,In_316);
or U5706 (N_5706,In_652,In_597);
or U5707 (N_5707,In_1711,In_1375);
xnor U5708 (N_5708,In_2791,In_561);
nand U5709 (N_5709,In_2974,In_213);
xnor U5710 (N_5710,In_2097,In_2609);
xor U5711 (N_5711,In_1373,In_1808);
xnor U5712 (N_5712,In_2313,In_2691);
xor U5713 (N_5713,In_1337,In_2653);
xnor U5714 (N_5714,In_1328,In_2369);
nor U5715 (N_5715,In_1288,In_2746);
xnor U5716 (N_5716,In_735,In_2006);
xnor U5717 (N_5717,In_580,In_2463);
or U5718 (N_5718,In_33,In_1843);
xor U5719 (N_5719,In_2655,In_471);
or U5720 (N_5720,In_167,In_1532);
nor U5721 (N_5721,In_1282,In_294);
nor U5722 (N_5722,In_2574,In_1051);
and U5723 (N_5723,In_1751,In_2220);
nor U5724 (N_5724,In_421,In_357);
nor U5725 (N_5725,In_253,In_1295);
nor U5726 (N_5726,In_2991,In_1510);
nor U5727 (N_5727,In_682,In_791);
nand U5728 (N_5728,In_1826,In_1527);
and U5729 (N_5729,In_833,In_2787);
and U5730 (N_5730,In_755,In_2065);
nor U5731 (N_5731,In_149,In_910);
or U5732 (N_5732,In_2596,In_999);
nor U5733 (N_5733,In_608,In_2888);
or U5734 (N_5734,In_1591,In_49);
xor U5735 (N_5735,In_1699,In_1683);
or U5736 (N_5736,In_874,In_2482);
nor U5737 (N_5737,In_1142,In_342);
and U5738 (N_5738,In_1148,In_1576);
and U5739 (N_5739,In_509,In_15);
or U5740 (N_5740,In_1328,In_2281);
nor U5741 (N_5741,In_2257,In_947);
or U5742 (N_5742,In_2253,In_877);
nor U5743 (N_5743,In_46,In_2255);
xor U5744 (N_5744,In_1604,In_1655);
nand U5745 (N_5745,In_2095,In_741);
nand U5746 (N_5746,In_672,In_429);
and U5747 (N_5747,In_1757,In_1979);
or U5748 (N_5748,In_2976,In_2516);
or U5749 (N_5749,In_666,In_2786);
nand U5750 (N_5750,In_1545,In_2878);
xnor U5751 (N_5751,In_1733,In_2289);
nor U5752 (N_5752,In_1610,In_1016);
or U5753 (N_5753,In_1295,In_2576);
xnor U5754 (N_5754,In_1177,In_938);
or U5755 (N_5755,In_843,In_867);
nor U5756 (N_5756,In_1875,In_2080);
or U5757 (N_5757,In_1797,In_2058);
and U5758 (N_5758,In_2372,In_1120);
xnor U5759 (N_5759,In_1247,In_745);
and U5760 (N_5760,In_2464,In_1664);
and U5761 (N_5761,In_1539,In_873);
nor U5762 (N_5762,In_1892,In_2466);
nor U5763 (N_5763,In_1920,In_324);
xnor U5764 (N_5764,In_290,In_589);
nor U5765 (N_5765,In_584,In_1963);
xor U5766 (N_5766,In_1964,In_966);
nand U5767 (N_5767,In_1197,In_2744);
and U5768 (N_5768,In_1411,In_868);
or U5769 (N_5769,In_1128,In_1084);
nor U5770 (N_5770,In_1236,In_148);
or U5771 (N_5771,In_2420,In_2816);
xnor U5772 (N_5772,In_266,In_1774);
xor U5773 (N_5773,In_911,In_1922);
xor U5774 (N_5774,In_1651,In_1706);
nand U5775 (N_5775,In_2197,In_772);
nor U5776 (N_5776,In_2138,In_1586);
nand U5777 (N_5777,In_2639,In_753);
nor U5778 (N_5778,In_2227,In_2560);
or U5779 (N_5779,In_2213,In_2934);
xnor U5780 (N_5780,In_2656,In_2405);
nand U5781 (N_5781,In_1241,In_2576);
nand U5782 (N_5782,In_426,In_227);
and U5783 (N_5783,In_485,In_2292);
xor U5784 (N_5784,In_2891,In_2235);
nand U5785 (N_5785,In_2073,In_1707);
nand U5786 (N_5786,In_1135,In_690);
and U5787 (N_5787,In_1670,In_1074);
nor U5788 (N_5788,In_1444,In_835);
nand U5789 (N_5789,In_2049,In_1674);
xnor U5790 (N_5790,In_314,In_737);
and U5791 (N_5791,In_1454,In_169);
nor U5792 (N_5792,In_2702,In_1639);
nor U5793 (N_5793,In_922,In_2186);
nor U5794 (N_5794,In_2032,In_2650);
nor U5795 (N_5795,In_1374,In_2322);
nor U5796 (N_5796,In_958,In_1910);
nand U5797 (N_5797,In_457,In_2795);
nor U5798 (N_5798,In_719,In_968);
nor U5799 (N_5799,In_2068,In_1152);
and U5800 (N_5800,In_1136,In_2707);
nor U5801 (N_5801,In_2652,In_234);
xor U5802 (N_5802,In_1055,In_2239);
or U5803 (N_5803,In_1811,In_2173);
and U5804 (N_5804,In_1226,In_1067);
nand U5805 (N_5805,In_2834,In_2508);
xnor U5806 (N_5806,In_2539,In_2820);
and U5807 (N_5807,In_2783,In_2885);
and U5808 (N_5808,In_2554,In_430);
nor U5809 (N_5809,In_865,In_185);
xor U5810 (N_5810,In_2689,In_2254);
or U5811 (N_5811,In_609,In_2120);
or U5812 (N_5812,In_244,In_206);
and U5813 (N_5813,In_1669,In_2389);
or U5814 (N_5814,In_585,In_202);
nand U5815 (N_5815,In_141,In_2613);
nor U5816 (N_5816,In_42,In_2084);
or U5817 (N_5817,In_1348,In_2936);
or U5818 (N_5818,In_1149,In_987);
nor U5819 (N_5819,In_1456,In_1945);
xnor U5820 (N_5820,In_2382,In_642);
xnor U5821 (N_5821,In_2856,In_2285);
xor U5822 (N_5822,In_2540,In_2521);
nand U5823 (N_5823,In_2008,In_735);
xnor U5824 (N_5824,In_2764,In_1406);
nor U5825 (N_5825,In_2321,In_1068);
or U5826 (N_5826,In_864,In_2037);
or U5827 (N_5827,In_1674,In_2059);
nand U5828 (N_5828,In_1460,In_1289);
xnor U5829 (N_5829,In_1904,In_937);
or U5830 (N_5830,In_1737,In_442);
xor U5831 (N_5831,In_1299,In_2350);
xnor U5832 (N_5832,In_467,In_2576);
nand U5833 (N_5833,In_1235,In_2129);
xnor U5834 (N_5834,In_67,In_215);
nand U5835 (N_5835,In_1196,In_2272);
and U5836 (N_5836,In_1280,In_627);
nand U5837 (N_5837,In_587,In_402);
and U5838 (N_5838,In_2650,In_835);
xnor U5839 (N_5839,In_1558,In_15);
and U5840 (N_5840,In_319,In_2603);
or U5841 (N_5841,In_1734,In_2111);
nand U5842 (N_5842,In_2530,In_425);
and U5843 (N_5843,In_2391,In_1543);
xnor U5844 (N_5844,In_2941,In_2214);
nor U5845 (N_5845,In_2113,In_2423);
xor U5846 (N_5846,In_1987,In_1444);
and U5847 (N_5847,In_33,In_1460);
nand U5848 (N_5848,In_2902,In_1485);
xnor U5849 (N_5849,In_1420,In_537);
xnor U5850 (N_5850,In_24,In_1553);
xnor U5851 (N_5851,In_521,In_1128);
nand U5852 (N_5852,In_1735,In_2359);
or U5853 (N_5853,In_2985,In_1423);
xor U5854 (N_5854,In_1146,In_301);
or U5855 (N_5855,In_28,In_464);
and U5856 (N_5856,In_252,In_595);
xnor U5857 (N_5857,In_705,In_2900);
nor U5858 (N_5858,In_2218,In_2217);
and U5859 (N_5859,In_6,In_2436);
nand U5860 (N_5860,In_2964,In_1694);
and U5861 (N_5861,In_2002,In_2331);
nand U5862 (N_5862,In_113,In_934);
and U5863 (N_5863,In_1876,In_181);
and U5864 (N_5864,In_2128,In_610);
and U5865 (N_5865,In_2428,In_2633);
and U5866 (N_5866,In_2956,In_1957);
xor U5867 (N_5867,In_2986,In_1126);
or U5868 (N_5868,In_1945,In_1401);
nand U5869 (N_5869,In_24,In_2729);
and U5870 (N_5870,In_2401,In_1559);
xnor U5871 (N_5871,In_787,In_1283);
xor U5872 (N_5872,In_2071,In_2734);
or U5873 (N_5873,In_2982,In_9);
nor U5874 (N_5874,In_1453,In_905);
xor U5875 (N_5875,In_1676,In_1478);
nand U5876 (N_5876,In_1312,In_2362);
and U5877 (N_5877,In_1338,In_2049);
nor U5878 (N_5878,In_1386,In_283);
nor U5879 (N_5879,In_2067,In_2891);
nor U5880 (N_5880,In_953,In_1919);
and U5881 (N_5881,In_934,In_1898);
and U5882 (N_5882,In_868,In_14);
xor U5883 (N_5883,In_2928,In_2987);
and U5884 (N_5884,In_2752,In_605);
nor U5885 (N_5885,In_2787,In_755);
or U5886 (N_5886,In_2201,In_38);
or U5887 (N_5887,In_460,In_140);
nor U5888 (N_5888,In_1156,In_2662);
or U5889 (N_5889,In_1424,In_683);
nand U5890 (N_5890,In_569,In_2523);
and U5891 (N_5891,In_501,In_2168);
xnor U5892 (N_5892,In_2862,In_2608);
and U5893 (N_5893,In_2166,In_2196);
or U5894 (N_5894,In_1079,In_1443);
xnor U5895 (N_5895,In_2091,In_2082);
xnor U5896 (N_5896,In_2544,In_1201);
xor U5897 (N_5897,In_1012,In_1314);
nand U5898 (N_5898,In_2299,In_2614);
nor U5899 (N_5899,In_1590,In_1947);
or U5900 (N_5900,In_852,In_2424);
xnor U5901 (N_5901,In_1096,In_1186);
nor U5902 (N_5902,In_2698,In_500);
or U5903 (N_5903,In_1365,In_1083);
and U5904 (N_5904,In_1907,In_1020);
nand U5905 (N_5905,In_1308,In_1346);
and U5906 (N_5906,In_860,In_2818);
nand U5907 (N_5907,In_928,In_2093);
nand U5908 (N_5908,In_1520,In_99);
nor U5909 (N_5909,In_667,In_2253);
and U5910 (N_5910,In_831,In_2308);
nor U5911 (N_5911,In_2239,In_1903);
xnor U5912 (N_5912,In_2872,In_1232);
nand U5913 (N_5913,In_1324,In_232);
and U5914 (N_5914,In_453,In_122);
or U5915 (N_5915,In_1397,In_750);
nand U5916 (N_5916,In_2033,In_1006);
nand U5917 (N_5917,In_693,In_121);
nor U5918 (N_5918,In_1600,In_0);
and U5919 (N_5919,In_1363,In_1895);
or U5920 (N_5920,In_1522,In_2876);
nand U5921 (N_5921,In_46,In_312);
or U5922 (N_5922,In_2513,In_826);
and U5923 (N_5923,In_2260,In_1599);
and U5924 (N_5924,In_2664,In_414);
and U5925 (N_5925,In_1470,In_2543);
xor U5926 (N_5926,In_2923,In_450);
nand U5927 (N_5927,In_1805,In_1177);
nand U5928 (N_5928,In_755,In_2340);
xor U5929 (N_5929,In_1972,In_1734);
nor U5930 (N_5930,In_1785,In_2718);
or U5931 (N_5931,In_1145,In_1015);
or U5932 (N_5932,In_864,In_1332);
xnor U5933 (N_5933,In_479,In_2401);
xor U5934 (N_5934,In_166,In_2599);
nor U5935 (N_5935,In_1429,In_1914);
and U5936 (N_5936,In_2650,In_870);
nor U5937 (N_5937,In_1631,In_1239);
nor U5938 (N_5938,In_2063,In_295);
xor U5939 (N_5939,In_1604,In_2352);
or U5940 (N_5940,In_1032,In_465);
nor U5941 (N_5941,In_2851,In_2556);
and U5942 (N_5942,In_476,In_1655);
xor U5943 (N_5943,In_566,In_179);
xnor U5944 (N_5944,In_2162,In_280);
nand U5945 (N_5945,In_626,In_522);
or U5946 (N_5946,In_1057,In_25);
and U5947 (N_5947,In_1491,In_1847);
nand U5948 (N_5948,In_2288,In_1247);
nand U5949 (N_5949,In_1715,In_2115);
or U5950 (N_5950,In_449,In_1560);
nand U5951 (N_5951,In_386,In_1299);
nor U5952 (N_5952,In_2953,In_2025);
nor U5953 (N_5953,In_103,In_2142);
nor U5954 (N_5954,In_204,In_474);
nand U5955 (N_5955,In_1272,In_1143);
and U5956 (N_5956,In_525,In_2933);
and U5957 (N_5957,In_2691,In_1306);
nand U5958 (N_5958,In_2034,In_2156);
xor U5959 (N_5959,In_2340,In_2698);
xnor U5960 (N_5960,In_102,In_389);
and U5961 (N_5961,In_2847,In_18);
nand U5962 (N_5962,In_505,In_521);
or U5963 (N_5963,In_155,In_2020);
or U5964 (N_5964,In_1042,In_2458);
nor U5965 (N_5965,In_434,In_2242);
and U5966 (N_5966,In_2768,In_2107);
or U5967 (N_5967,In_2015,In_984);
nand U5968 (N_5968,In_1157,In_906);
nor U5969 (N_5969,In_1141,In_1298);
xnor U5970 (N_5970,In_2983,In_1425);
nand U5971 (N_5971,In_2217,In_1795);
xor U5972 (N_5972,In_881,In_40);
nor U5973 (N_5973,In_1176,In_862);
nor U5974 (N_5974,In_834,In_1110);
nor U5975 (N_5975,In_1926,In_1573);
nand U5976 (N_5976,In_2301,In_1391);
nor U5977 (N_5977,In_2984,In_2956);
or U5978 (N_5978,In_1108,In_1855);
xnor U5979 (N_5979,In_2845,In_1605);
or U5980 (N_5980,In_2853,In_348);
or U5981 (N_5981,In_1480,In_244);
or U5982 (N_5982,In_727,In_1828);
or U5983 (N_5983,In_2059,In_1508);
nor U5984 (N_5984,In_1487,In_2232);
xnor U5985 (N_5985,In_2210,In_2405);
or U5986 (N_5986,In_1922,In_295);
nand U5987 (N_5987,In_2452,In_1369);
nand U5988 (N_5988,In_455,In_1857);
and U5989 (N_5989,In_2244,In_2582);
and U5990 (N_5990,In_1711,In_2278);
nand U5991 (N_5991,In_1059,In_1212);
and U5992 (N_5992,In_2644,In_772);
and U5993 (N_5993,In_20,In_625);
nor U5994 (N_5994,In_1458,In_1154);
nand U5995 (N_5995,In_1454,In_1865);
or U5996 (N_5996,In_2804,In_1670);
xor U5997 (N_5997,In_818,In_1514);
and U5998 (N_5998,In_1791,In_1482);
and U5999 (N_5999,In_443,In_1592);
or U6000 (N_6000,N_1922,N_2814);
nand U6001 (N_6001,N_4710,N_357);
nand U6002 (N_6002,N_697,N_2280);
or U6003 (N_6003,N_4215,N_3351);
nand U6004 (N_6004,N_5444,N_5646);
and U6005 (N_6005,N_3930,N_5578);
or U6006 (N_6006,N_4252,N_1881);
and U6007 (N_6007,N_3857,N_1292);
nor U6008 (N_6008,N_5759,N_3176);
nand U6009 (N_6009,N_1906,N_5615);
or U6010 (N_6010,N_1197,N_470);
nand U6011 (N_6011,N_5808,N_3321);
or U6012 (N_6012,N_5560,N_4937);
nor U6013 (N_6013,N_5075,N_4026);
xor U6014 (N_6014,N_4429,N_4806);
nand U6015 (N_6015,N_2378,N_4016);
nor U6016 (N_6016,N_1630,N_1527);
or U6017 (N_6017,N_13,N_2879);
nand U6018 (N_6018,N_1915,N_1963);
and U6019 (N_6019,N_2326,N_502);
xor U6020 (N_6020,N_2297,N_2774);
and U6021 (N_6021,N_3839,N_3311);
or U6022 (N_6022,N_4074,N_2987);
or U6023 (N_6023,N_2964,N_1543);
nor U6024 (N_6024,N_3335,N_4159);
xnor U6025 (N_6025,N_1165,N_5735);
xnor U6026 (N_6026,N_3314,N_2067);
or U6027 (N_6027,N_4824,N_4763);
and U6028 (N_6028,N_5068,N_2622);
nand U6029 (N_6029,N_1573,N_4418);
and U6030 (N_6030,N_4154,N_5472);
nor U6031 (N_6031,N_5270,N_693);
nand U6032 (N_6032,N_2702,N_909);
nor U6033 (N_6033,N_194,N_3158);
or U6034 (N_6034,N_1999,N_807);
nand U6035 (N_6035,N_1479,N_2382);
or U6036 (N_6036,N_3928,N_5458);
xnor U6037 (N_6037,N_5227,N_431);
xor U6038 (N_6038,N_3972,N_4715);
nand U6039 (N_6039,N_4441,N_3308);
nor U6040 (N_6040,N_5417,N_2670);
and U6041 (N_6041,N_3981,N_3906);
nor U6042 (N_6042,N_616,N_1582);
and U6043 (N_6043,N_5538,N_2211);
xnor U6044 (N_6044,N_4596,N_5933);
nand U6045 (N_6045,N_2085,N_3542);
or U6046 (N_6046,N_23,N_4239);
and U6047 (N_6047,N_1160,N_4156);
nor U6048 (N_6048,N_703,N_2626);
nand U6049 (N_6049,N_3221,N_4296);
nand U6050 (N_6050,N_4373,N_1576);
xnor U6051 (N_6051,N_3407,N_2205);
or U6052 (N_6052,N_340,N_113);
nand U6053 (N_6053,N_3924,N_3389);
nor U6054 (N_6054,N_1360,N_2639);
and U6055 (N_6055,N_3649,N_4845);
and U6056 (N_6056,N_769,N_56);
and U6057 (N_6057,N_4394,N_5089);
nor U6058 (N_6058,N_3433,N_463);
or U6059 (N_6059,N_3125,N_5819);
xor U6060 (N_6060,N_5035,N_973);
and U6061 (N_6061,N_52,N_5609);
nor U6062 (N_6062,N_5876,N_2552);
and U6063 (N_6063,N_1417,N_1972);
xor U6064 (N_6064,N_1955,N_135);
and U6065 (N_6065,N_5721,N_3250);
and U6066 (N_6066,N_2929,N_1715);
or U6067 (N_6067,N_2801,N_4619);
nor U6068 (N_6068,N_1718,N_3485);
and U6069 (N_6069,N_2673,N_4096);
nand U6070 (N_6070,N_3022,N_543);
nor U6071 (N_6071,N_4623,N_2535);
or U6072 (N_6072,N_551,N_5673);
nand U6073 (N_6073,N_3681,N_2782);
nor U6074 (N_6074,N_2060,N_704);
nor U6075 (N_6075,N_3801,N_4352);
nand U6076 (N_6076,N_5674,N_5670);
nor U6077 (N_6077,N_3556,N_68);
or U6078 (N_6078,N_992,N_1953);
nor U6079 (N_6079,N_455,N_2548);
nand U6080 (N_6080,N_4990,N_5138);
or U6081 (N_6081,N_4204,N_507);
or U6082 (N_6082,N_421,N_4365);
nor U6083 (N_6083,N_4166,N_3821);
nor U6084 (N_6084,N_2777,N_1453);
nand U6085 (N_6085,N_1854,N_1656);
xnor U6086 (N_6086,N_5657,N_5934);
nand U6087 (N_6087,N_145,N_2816);
or U6088 (N_6088,N_2383,N_4905);
or U6089 (N_6089,N_3148,N_2824);
and U6090 (N_6090,N_4967,N_2612);
and U6091 (N_6091,N_1609,N_2331);
xor U6092 (N_6092,N_428,N_14);
xor U6093 (N_6093,N_1956,N_4588);
xnor U6094 (N_6094,N_2808,N_1445);
xnor U6095 (N_6095,N_3716,N_4920);
or U6096 (N_6096,N_5466,N_2831);
nand U6097 (N_6097,N_5675,N_2339);
xor U6098 (N_6098,N_3073,N_1845);
and U6099 (N_6099,N_3004,N_744);
nor U6100 (N_6100,N_5800,N_3040);
nor U6101 (N_6101,N_5237,N_5151);
and U6102 (N_6102,N_822,N_4674);
or U6103 (N_6103,N_3653,N_5481);
nor U6104 (N_6104,N_696,N_2836);
or U6105 (N_6105,N_5799,N_511);
and U6106 (N_6106,N_2266,N_1572);
nand U6107 (N_6107,N_5783,N_5083);
xor U6108 (N_6108,N_3420,N_970);
xnor U6109 (N_6109,N_1986,N_4288);
and U6110 (N_6110,N_2971,N_1615);
or U6111 (N_6111,N_454,N_1105);
nand U6112 (N_6112,N_451,N_1201);
and U6113 (N_6113,N_2656,N_1739);
nor U6114 (N_6114,N_1920,N_2985);
xor U6115 (N_6115,N_1699,N_2177);
nand U6116 (N_6116,N_5985,N_1745);
and U6117 (N_6117,N_1202,N_3570);
nor U6118 (N_6118,N_3108,N_1109);
xnor U6119 (N_6119,N_3401,N_3746);
nand U6120 (N_6120,N_602,N_5376);
or U6121 (N_6121,N_1200,N_1196);
nand U6122 (N_6122,N_3275,N_2104);
xor U6123 (N_6123,N_479,N_120);
nor U6124 (N_6124,N_1566,N_2516);
or U6125 (N_6125,N_5119,N_3168);
and U6126 (N_6126,N_2410,N_5339);
nor U6127 (N_6127,N_2097,N_4549);
and U6128 (N_6128,N_1096,N_2487);
or U6129 (N_6129,N_2883,N_4102);
nor U6130 (N_6130,N_4907,N_5047);
nor U6131 (N_6131,N_2772,N_4769);
and U6132 (N_6132,N_3478,N_2446);
nand U6133 (N_6133,N_778,N_3009);
nand U6134 (N_6134,N_1541,N_1125);
and U6135 (N_6135,N_5272,N_3664);
or U6136 (N_6136,N_4283,N_1977);
xnor U6137 (N_6137,N_718,N_2329);
nand U6138 (N_6138,N_4271,N_1636);
nand U6139 (N_6139,N_781,N_5972);
nand U6140 (N_6140,N_4278,N_4950);
nand U6141 (N_6141,N_1632,N_1242);
xor U6142 (N_6142,N_5094,N_3267);
or U6143 (N_6143,N_984,N_5568);
xor U6144 (N_6144,N_1155,N_5910);
nand U6145 (N_6145,N_1450,N_1907);
or U6146 (N_6146,N_2397,N_295);
or U6147 (N_6147,N_917,N_3499);
xnor U6148 (N_6148,N_5370,N_4129);
nor U6149 (N_6149,N_4043,N_257);
xor U6150 (N_6150,N_1730,N_2235);
and U6151 (N_6151,N_2779,N_5145);
xnor U6152 (N_6152,N_4675,N_413);
and U6153 (N_6153,N_3013,N_2371);
nor U6154 (N_6154,N_228,N_2401);
nand U6155 (N_6155,N_1776,N_3956);
and U6156 (N_6156,N_1813,N_3090);
nand U6157 (N_6157,N_5400,N_3259);
nand U6158 (N_6158,N_423,N_309);
and U6159 (N_6159,N_2722,N_2030);
nand U6160 (N_6160,N_934,N_4005);
nor U6161 (N_6161,N_348,N_5719);
xnor U6162 (N_6162,N_3110,N_5822);
or U6163 (N_6163,N_1114,N_4938);
nand U6164 (N_6164,N_5590,N_4324);
xnor U6165 (N_6165,N_1713,N_5575);
and U6166 (N_6166,N_1993,N_3779);
xor U6167 (N_6167,N_4451,N_5832);
xnor U6168 (N_6168,N_4458,N_5383);
or U6169 (N_6169,N_5618,N_99);
or U6170 (N_6170,N_356,N_1128);
nor U6171 (N_6171,N_2792,N_2314);
nand U6172 (N_6172,N_1103,N_2823);
or U6173 (N_6173,N_3195,N_1001);
xor U6174 (N_6174,N_1753,N_4898);
nor U6175 (N_6175,N_1394,N_1800);
or U6176 (N_6176,N_374,N_4238);
nor U6177 (N_6177,N_5285,N_5346);
or U6178 (N_6178,N_1244,N_5108);
xnor U6179 (N_6179,N_2479,N_2684);
nor U6180 (N_6180,N_2784,N_2206);
or U6181 (N_6181,N_2385,N_473);
nor U6182 (N_6182,N_2138,N_4522);
xnor U6183 (N_6183,N_512,N_1011);
or U6184 (N_6184,N_544,N_5610);
nand U6185 (N_6185,N_2583,N_4290);
and U6186 (N_6186,N_4251,N_2467);
nand U6187 (N_6187,N_5660,N_3589);
nand U6188 (N_6188,N_3634,N_1494);
or U6189 (N_6189,N_1552,N_1760);
nand U6190 (N_6190,N_3369,N_2643);
nor U6191 (N_6191,N_219,N_1343);
xor U6192 (N_6192,N_3490,N_2947);
nand U6193 (N_6193,N_1659,N_4878);
nand U6194 (N_6194,N_854,N_5510);
nand U6195 (N_6195,N_2727,N_3309);
or U6196 (N_6196,N_1311,N_5366);
and U6197 (N_6197,N_1838,N_5511);
nor U6198 (N_6198,N_1618,N_3403);
and U6199 (N_6199,N_43,N_5261);
or U6200 (N_6200,N_5414,N_42);
nor U6201 (N_6201,N_4205,N_2995);
and U6202 (N_6202,N_5975,N_2277);
nor U6203 (N_6203,N_5943,N_5824);
or U6204 (N_6204,N_1498,N_3353);
xnor U6205 (N_6205,N_636,N_4191);
nand U6206 (N_6206,N_169,N_4038);
xor U6207 (N_6207,N_4230,N_5627);
nand U6208 (N_6208,N_1476,N_2386);
and U6209 (N_6209,N_5010,N_5267);
xnor U6210 (N_6210,N_4110,N_232);
nand U6211 (N_6211,N_5837,N_184);
xor U6212 (N_6212,N_4476,N_899);
or U6213 (N_6213,N_5203,N_1239);
and U6214 (N_6214,N_4354,N_2754);
or U6215 (N_6215,N_2146,N_5263);
nor U6216 (N_6216,N_1735,N_3937);
nor U6217 (N_6217,N_1270,N_1454);
nand U6218 (N_6218,N_3838,N_2047);
and U6219 (N_6219,N_4218,N_4537);
and U6220 (N_6220,N_119,N_5002);
or U6221 (N_6221,N_4209,N_5844);
and U6222 (N_6222,N_311,N_1828);
and U6223 (N_6223,N_3592,N_5197);
nor U6224 (N_6224,N_280,N_2550);
nor U6225 (N_6225,N_318,N_2338);
nor U6226 (N_6226,N_4217,N_504);
and U6227 (N_6227,N_4683,N_5153);
or U6228 (N_6228,N_1116,N_529);
nor U6229 (N_6229,N_3382,N_2515);
nor U6230 (N_6230,N_1875,N_3208);
nand U6231 (N_6231,N_4380,N_3487);
nor U6232 (N_6232,N_5738,N_4100);
nand U6233 (N_6233,N_3510,N_4951);
nand U6234 (N_6234,N_3896,N_692);
xnor U6235 (N_6235,N_5073,N_3751);
nor U6236 (N_6236,N_5318,N_1625);
nor U6237 (N_6237,N_5730,N_2368);
nor U6238 (N_6238,N_126,N_2086);
nor U6239 (N_6239,N_5435,N_1965);
and U6240 (N_6240,N_3772,N_203);
and U6241 (N_6241,N_418,N_121);
nand U6242 (N_6242,N_5485,N_5881);
or U6243 (N_6243,N_5654,N_399);
nand U6244 (N_6244,N_1411,N_4015);
and U6245 (N_6245,N_4449,N_2426);
and U6246 (N_6246,N_5632,N_5535);
and U6247 (N_6247,N_5186,N_1209);
and U6248 (N_6248,N_185,N_5885);
nand U6249 (N_6249,N_2288,N_4659);
and U6250 (N_6250,N_5976,N_3650);
xor U6251 (N_6251,N_1621,N_3619);
xor U6252 (N_6252,N_1617,N_953);
nand U6253 (N_6253,N_654,N_3248);
or U6254 (N_6254,N_2930,N_5322);
nor U6255 (N_6255,N_3782,N_1748);
and U6256 (N_6256,N_5701,N_5310);
xor U6257 (N_6257,N_3990,N_2263);
nor U6258 (N_6258,N_3977,N_1474);
nor U6259 (N_6259,N_133,N_4243);
xor U6260 (N_6260,N_599,N_5358);
xnor U6261 (N_6261,N_4964,N_1283);
xnor U6262 (N_6262,N_914,N_499);
nand U6263 (N_6263,N_1747,N_3819);
nor U6264 (N_6264,N_424,N_2915);
nand U6265 (N_6265,N_3234,N_74);
nand U6266 (N_6266,N_3568,N_2618);
nor U6267 (N_6267,N_4499,N_1338);
or U6268 (N_6268,N_3647,N_5781);
or U6269 (N_6269,N_1215,N_4481);
nor U6270 (N_6270,N_405,N_3093);
xor U6271 (N_6271,N_3427,N_4842);
or U6272 (N_6272,N_5296,N_3171);
and U6273 (N_6273,N_3367,N_5826);
and U6274 (N_6274,N_1939,N_2509);
nand U6275 (N_6275,N_2644,N_1810);
nor U6276 (N_6276,N_429,N_5428);
and U6277 (N_6277,N_2696,N_4104);
nand U6278 (N_6278,N_3260,N_5234);
nand U6279 (N_6279,N_3492,N_3235);
or U6280 (N_6280,N_2681,N_5054);
nor U6281 (N_6281,N_16,N_885);
nor U6282 (N_6282,N_2492,N_736);
nand U6283 (N_6283,N_5103,N_2720);
or U6284 (N_6284,N_4464,N_823);
nand U6285 (N_6285,N_324,N_2141);
nor U6286 (N_6286,N_3062,N_5231);
or U6287 (N_6287,N_5091,N_4287);
xnor U6288 (N_6288,N_918,N_4770);
nor U6289 (N_6289,N_5529,N_818);
xor U6290 (N_6290,N_3758,N_2943);
xor U6291 (N_6291,N_2178,N_5816);
and U6292 (N_6292,N_5434,N_4616);
xor U6293 (N_6293,N_2623,N_3514);
xnor U6294 (N_6294,N_4334,N_4046);
or U6295 (N_6295,N_2707,N_2563);
and U6296 (N_6296,N_5982,N_4286);
nor U6297 (N_6297,N_2376,N_1214);
or U6298 (N_6298,N_2342,N_1113);
xor U6299 (N_6299,N_4186,N_1079);
nor U6300 (N_6300,N_2901,N_3359);
xor U6301 (N_6301,N_2756,N_2723);
nand U6302 (N_6302,N_4861,N_1307);
or U6303 (N_6303,N_3464,N_1862);
or U6304 (N_6304,N_3960,N_2208);
xor U6305 (N_6305,N_4203,N_1257);
xnor U6306 (N_6306,N_3038,N_2411);
nand U6307 (N_6307,N_3631,N_5167);
xnor U6308 (N_6308,N_1396,N_5912);
or U6309 (N_6309,N_4462,N_1683);
xor U6310 (N_6310,N_4448,N_4725);
nor U6311 (N_6311,N_5744,N_88);
xnor U6312 (N_6312,N_3481,N_5028);
or U6313 (N_6313,N_2282,N_5714);
nand U6314 (N_6314,N_2462,N_3722);
and U6315 (N_6315,N_5685,N_866);
nand U6316 (N_6316,N_956,N_819);
xor U6317 (N_6317,N_3693,N_4888);
nand U6318 (N_6318,N_808,N_1110);
or U6319 (N_6319,N_978,N_5342);
nand U6320 (N_6320,N_4000,N_508);
or U6321 (N_6321,N_4862,N_1637);
nand U6322 (N_6322,N_5382,N_5565);
and U6323 (N_6323,N_1542,N_4002);
nor U6324 (N_6324,N_2120,N_830);
nand U6325 (N_6325,N_5802,N_388);
and U6326 (N_6326,N_5490,N_4656);
or U6327 (N_6327,N_2053,N_1886);
nor U6328 (N_6328,N_5359,N_38);
nor U6329 (N_6329,N_5088,N_4644);
nor U6330 (N_6330,N_2911,N_4979);
nand U6331 (N_6331,N_5789,N_41);
nand U6332 (N_6332,N_3917,N_2853);
xor U6333 (N_6333,N_4846,N_5319);
xor U6334 (N_6334,N_3200,N_753);
nor U6335 (N_6335,N_832,N_361);
xor U6336 (N_6336,N_2179,N_1412);
or U6337 (N_6337,N_2858,N_3189);
or U6338 (N_6338,N_4632,N_1727);
xnor U6339 (N_6339,N_5527,N_1503);
nand U6340 (N_6340,N_2433,N_1485);
xor U6341 (N_6341,N_1712,N_2710);
or U6342 (N_6342,N_2237,N_3261);
nand U6343 (N_6343,N_2646,N_2525);
xnor U6344 (N_6344,N_3370,N_4784);
nor U6345 (N_6345,N_5845,N_5869);
nor U6346 (N_6346,N_2762,N_5829);
or U6347 (N_6347,N_2453,N_1189);
nor U6348 (N_6348,N_3421,N_4430);
and U6349 (N_6349,N_392,N_436);
and U6350 (N_6350,N_3963,N_552);
or U6351 (N_6351,N_5354,N_3338);
nor U6352 (N_6352,N_5361,N_2088);
or U6353 (N_6353,N_5212,N_2938);
nor U6354 (N_6354,N_3974,N_3086);
and U6355 (N_6355,N_2221,N_335);
nand U6356 (N_6356,N_2501,N_3231);
and U6357 (N_6357,N_2728,N_766);
nor U6358 (N_6358,N_2864,N_671);
xnor U6359 (N_6359,N_4151,N_2340);
nor U6360 (N_6360,N_967,N_5393);
xor U6361 (N_6361,N_4311,N_2490);
xnor U6362 (N_6362,N_3518,N_5301);
xor U6363 (N_6363,N_4320,N_186);
nand U6364 (N_6364,N_2917,N_4094);
nor U6365 (N_6365,N_4345,N_4306);
nand U6366 (N_6366,N_1047,N_3915);
or U6367 (N_6367,N_3894,N_110);
or U6368 (N_6368,N_3868,N_4189);
nor U6369 (N_6369,N_5061,N_2495);
xnor U6370 (N_6370,N_2829,N_252);
nor U6371 (N_6371,N_412,N_3871);
and U6372 (N_6372,N_3745,N_5731);
or U6373 (N_6373,N_1839,N_4376);
and U6374 (N_6374,N_3786,N_994);
xnor U6375 (N_6375,N_3547,N_3177);
nor U6376 (N_6376,N_4955,N_5818);
and U6377 (N_6377,N_702,N_3340);
xor U6378 (N_6378,N_3124,N_873);
or U6379 (N_6379,N_5637,N_4941);
and U6380 (N_6380,N_974,N_5230);
nand U6381 (N_6381,N_3263,N_247);
and U6382 (N_6382,N_1143,N_1850);
nor U6383 (N_6383,N_4602,N_5462);
nand U6384 (N_6384,N_2740,N_407);
or U6385 (N_6385,N_591,N_4075);
nand U6386 (N_6386,N_2741,N_584);
or U6387 (N_6387,N_789,N_319);
nor U6388 (N_6388,N_5132,N_648);
or U6389 (N_6389,N_4400,N_4018);
xnor U6390 (N_6390,N_2513,N_4140);
xor U6391 (N_6391,N_216,N_3656);
nor U6392 (N_6392,N_5653,N_1803);
or U6393 (N_6393,N_1526,N_1385);
and U6394 (N_6394,N_2532,N_5488);
or U6395 (N_6395,N_4216,N_5865);
xor U6396 (N_6396,N_5518,N_5160);
or U6397 (N_6397,N_5664,N_1274);
nor U6398 (N_6398,N_4450,N_1166);
nand U6399 (N_6399,N_1212,N_1589);
xnor U6400 (N_6400,N_4422,N_5955);
nor U6401 (N_6401,N_5468,N_1728);
and U6402 (N_6402,N_4411,N_5540);
nand U6403 (N_6403,N_5429,N_2481);
xnor U6404 (N_6404,N_815,N_1224);
nor U6405 (N_6405,N_1276,N_5962);
and U6406 (N_6406,N_2817,N_1616);
nor U6407 (N_6407,N_3160,N_5130);
nor U6408 (N_6408,N_4673,N_5202);
nand U6409 (N_6409,N_3159,N_3114);
xor U6410 (N_6410,N_3951,N_3383);
and U6411 (N_6411,N_1408,N_4384);
or U6412 (N_6412,N_5758,N_1737);
nor U6413 (N_6413,N_5124,N_1229);
or U6414 (N_6414,N_341,N_831);
nor U6415 (N_6415,N_513,N_1271);
nand U6416 (N_6416,N_1919,N_181);
xnor U6417 (N_6417,N_5063,N_1169);
nor U6418 (N_6418,N_3783,N_293);
nor U6419 (N_6419,N_4298,N_490);
and U6420 (N_6420,N_3931,N_3301);
and U6421 (N_6421,N_224,N_2040);
xnor U6422 (N_6422,N_577,N_3670);
and U6423 (N_6423,N_5165,N_5052);
nand U6424 (N_6424,N_2409,N_4744);
nand U6425 (N_6425,N_4021,N_1104);
nand U6426 (N_6426,N_2685,N_624);
or U6427 (N_6427,N_1357,N_2028);
or U6428 (N_6428,N_459,N_660);
nand U6429 (N_6429,N_5756,N_4030);
nand U6430 (N_6430,N_737,N_4658);
and U6431 (N_6431,N_444,N_5753);
nand U6432 (N_6432,N_549,N_2770);
or U6433 (N_6433,N_667,N_1220);
nor U6434 (N_6434,N_3796,N_1668);
nor U6435 (N_6435,N_1093,N_5453);
or U6436 (N_6436,N_1159,N_2232);
nor U6437 (N_6437,N_3067,N_4488);
nand U6438 (N_6438,N_925,N_3469);
or U6439 (N_6439,N_4375,N_1978);
nor U6440 (N_6440,N_3274,N_144);
nor U6441 (N_6441,N_1921,N_2024);
nand U6442 (N_6442,N_3241,N_474);
nand U6443 (N_6443,N_1688,N_1928);
xor U6444 (N_6444,N_4319,N_638);
nand U6445 (N_6445,N_2258,N_2498);
nand U6446 (N_6446,N_2645,N_177);
and U6447 (N_6447,N_4322,N_589);
and U6448 (N_6448,N_4711,N_2704);
and U6449 (N_6449,N_1984,N_2017);
nor U6450 (N_6450,N_2281,N_3423);
nand U6451 (N_6451,N_2021,N_833);
and U6452 (N_6452,N_2921,N_1183);
nor U6453 (N_6453,N_2455,N_1329);
xnor U6454 (N_6454,N_487,N_3545);
nand U6455 (N_6455,N_5513,N_5946);
xor U6456 (N_6456,N_2175,N_3138);
xor U6457 (N_6457,N_3940,N_4913);
nor U6458 (N_6458,N_2695,N_2093);
or U6459 (N_6459,N_3289,N_1899);
nor U6460 (N_6460,N_4027,N_4275);
nor U6461 (N_6461,N_2508,N_5880);
or U6462 (N_6462,N_4007,N_2344);
nor U6463 (N_6463,N_4370,N_2002);
nand U6464 (N_6464,N_1664,N_5110);
nor U6465 (N_6465,N_570,N_3719);
or U6466 (N_6466,N_2553,N_2896);
xnor U6467 (N_6467,N_612,N_5984);
or U6468 (N_6468,N_323,N_840);
or U6469 (N_6469,N_1309,N_1514);
or U6470 (N_6470,N_3593,N_321);
xnor U6471 (N_6471,N_5288,N_5120);
or U6472 (N_6472,N_545,N_3968);
and U6473 (N_6473,N_4848,N_4641);
or U6474 (N_6474,N_1778,N_3455);
nor U6475 (N_6475,N_1891,N_5945);
nor U6476 (N_6476,N_489,N_3677);
nor U6477 (N_6477,N_2299,N_4568);
nor U6478 (N_6478,N_1871,N_1458);
nor U6479 (N_6479,N_2071,N_358);
xnor U6480 (N_6480,N_471,N_3640);
nand U6481 (N_6481,N_325,N_1949);
nor U6482 (N_6482,N_533,N_4177);
or U6483 (N_6483,N_45,N_834);
nor U6484 (N_6484,N_1258,N_1944);
nor U6485 (N_6485,N_5093,N_1994);
and U6486 (N_6486,N_859,N_1341);
nor U6487 (N_6487,N_5623,N_1491);
or U6488 (N_6488,N_614,N_8);
xnor U6489 (N_6489,N_2447,N_278);
and U6490 (N_6490,N_3803,N_4474);
xnor U6491 (N_6491,N_5062,N_814);
or U6492 (N_6492,N_3955,N_597);
or U6493 (N_6493,N_5693,N_5207);
nor U6494 (N_6494,N_1440,N_4922);
or U6495 (N_6495,N_4126,N_5209);
or U6496 (N_6496,N_4531,N_3092);
nand U6497 (N_6497,N_1792,N_2845);
or U6498 (N_6498,N_3399,N_1734);
xnor U6499 (N_6499,N_4023,N_4986);
and U6500 (N_6500,N_4771,N_576);
xor U6501 (N_6501,N_4628,N_3494);
nor U6502 (N_6502,N_5579,N_5638);
or U6503 (N_6503,N_1964,N_3907);
nor U6504 (N_6504,N_4789,N_1375);
xor U6505 (N_6505,N_2004,N_4740);
or U6506 (N_6506,N_1952,N_5862);
nor U6507 (N_6507,N_3622,N_2204);
and U6508 (N_6508,N_1492,N_5308);
nor U6509 (N_6509,N_4182,N_2610);
and U6510 (N_6510,N_2539,N_2627);
nand U6511 (N_6511,N_1876,N_249);
or U6512 (N_6512,N_2057,N_1363);
nor U6513 (N_6513,N_2881,N_2049);
nor U6514 (N_6514,N_4234,N_3759);
or U6515 (N_6515,N_5833,N_767);
and U6516 (N_6516,N_1732,N_2261);
nor U6517 (N_6517,N_3897,N_2202);
or U6518 (N_6518,N_3426,N_132);
and U6519 (N_6519,N_2254,N_4423);
nor U6520 (N_6520,N_1301,N_29);
and U6521 (N_6521,N_4621,N_3337);
and U6522 (N_6522,N_2052,N_80);
nor U6523 (N_6523,N_3098,N_5605);
or U6524 (N_6524,N_2628,N_2270);
and U6525 (N_6525,N_3018,N_1987);
nand U6526 (N_6526,N_3016,N_2542);
xnor U6527 (N_6527,N_2375,N_3295);
nor U6528 (N_6528,N_2856,N_4069);
nor U6529 (N_6529,N_4442,N_3167);
xor U6530 (N_6530,N_2228,N_5642);
xnor U6531 (N_6531,N_3290,N_3816);
or U6532 (N_6532,N_2837,N_5733);
and U6533 (N_6533,N_4523,N_5099);
nand U6534 (N_6534,N_5866,N_2918);
or U6535 (N_6535,N_2109,N_166);
and U6536 (N_6536,N_1826,N_2394);
or U6537 (N_6537,N_176,N_2868);
and U6538 (N_6538,N_5964,N_5765);
nor U6539 (N_6539,N_5619,N_4684);
xnor U6540 (N_6540,N_71,N_2732);
nor U6541 (N_6541,N_1496,N_76);
xnor U6542 (N_6542,N_5922,N_3465);
and U6543 (N_6543,N_5852,N_3162);
nand U6544 (N_6544,N_5780,N_2262);
nor U6545 (N_6545,N_5097,N_1742);
nor U6546 (N_6546,N_2337,N_1462);
or U6547 (N_6547,N_122,N_1645);
xor U6548 (N_6548,N_3654,N_4412);
xnor U6549 (N_6549,N_4586,N_5247);
nor U6550 (N_6550,N_1331,N_3802);
xor U6551 (N_6551,N_5175,N_5142);
nand U6552 (N_6552,N_5864,N_4857);
or U6553 (N_6553,N_5525,N_5014);
and U6554 (N_6554,N_608,N_5572);
and U6555 (N_6555,N_3811,N_4578);
nand U6556 (N_6556,N_2968,N_690);
nor U6557 (N_6557,N_5273,N_5078);
nand U6558 (N_6558,N_4973,N_510);
or U6559 (N_6559,N_2315,N_874);
or U6560 (N_6560,N_5051,N_3952);
nand U6561 (N_6561,N_3581,N_1150);
xnor U6562 (N_6562,N_2015,N_1690);
nand U6563 (N_6563,N_1352,N_383);
or U6564 (N_6564,N_3682,N_5636);
xor U6565 (N_6565,N_274,N_4257);
nand U6566 (N_6566,N_1406,N_4511);
nor U6567 (N_6567,N_2286,N_2888);
xnor U6568 (N_6568,N_2099,N_639);
nor U6569 (N_6569,N_5038,N_4852);
or U6570 (N_6570,N_682,N_4526);
xor U6571 (N_6571,N_2068,N_3873);
xor U6572 (N_6572,N_4087,N_3588);
nand U6573 (N_6573,N_4750,N_610);
nand U6574 (N_6574,N_4556,N_5842);
nor U6575 (N_6575,N_5678,N_4963);
or U6576 (N_6576,N_3329,N_1578);
nand U6577 (N_6577,N_4,N_4366);
and U6578 (N_6578,N_1808,N_3665);
nand U6579 (N_6579,N_5125,N_1914);
xor U6580 (N_6580,N_1433,N_1217);
nand U6581 (N_6581,N_3284,N_1590);
or U6582 (N_6582,N_4113,N_5797);
nand U6583 (N_6583,N_2859,N_2940);
and U6584 (N_6584,N_379,N_4142);
and U6585 (N_6585,N_1587,N_491);
nor U6586 (N_6586,N_2157,N_4908);
nor U6587 (N_6587,N_828,N_5431);
and U6588 (N_6588,N_1954,N_3626);
or U6589 (N_6589,N_2689,N_4535);
xnor U6590 (N_6590,N_2989,N_4220);
nand U6591 (N_6591,N_1364,N_3844);
xnor U6592 (N_6592,N_1061,N_4893);
or U6593 (N_6593,N_331,N_4592);
or U6594 (N_6594,N_4419,N_2186);
nand U6595 (N_6595,N_603,N_4503);
nor U6596 (N_6596,N_2169,N_5222);
nor U6597 (N_6597,N_2173,N_4059);
and U6598 (N_6598,N_3408,N_1393);
or U6599 (N_6599,N_5639,N_716);
nor U6600 (N_6600,N_784,N_1137);
nand U6601 (N_6601,N_4685,N_4121);
nand U6602 (N_6602,N_2894,N_4109);
nand U6603 (N_6603,N_3115,N_1610);
or U6604 (N_6604,N_67,N_415);
and U6605 (N_6605,N_862,N_1752);
and U6606 (N_6606,N_995,N_1893);
nand U6607 (N_6607,N_4525,N_3738);
nor U6608 (N_6608,N_371,N_2006);
and U6609 (N_6609,N_2967,N_4460);
nand U6610 (N_6610,N_3081,N_3632);
xor U6611 (N_6611,N_2428,N_2775);
and U6612 (N_6612,N_1455,N_109);
xnor U6613 (N_6613,N_5906,N_4970);
nand U6614 (N_6614,N_2132,N_291);
nor U6615 (N_6615,N_5096,N_3431);
nand U6616 (N_6616,N_1551,N_2677);
nand U6617 (N_6617,N_2844,N_2353);
and U6618 (N_6618,N_746,N_3151);
or U6619 (N_6619,N_2861,N_3627);
or U6620 (N_6620,N_3625,N_4805);
nor U6621 (N_6621,N_3561,N_3107);
and U6622 (N_6622,N_5709,N_4292);
xor U6623 (N_6623,N_3330,N_4524);
nor U6624 (N_6624,N_5042,N_3725);
and U6625 (N_6625,N_1868,N_1513);
nor U6626 (N_6626,N_2227,N_70);
nand U6627 (N_6627,N_897,N_336);
and U6628 (N_6628,N_2198,N_892);
or U6629 (N_6629,N_1878,N_2035);
and U6630 (N_6630,N_1709,N_3617);
nand U6631 (N_6631,N_4471,N_4082);
xnor U6632 (N_6632,N_2878,N_1228);
or U6633 (N_6633,N_2351,N_5835);
and U6634 (N_6634,N_999,N_3386);
nor U6635 (N_6635,N_1722,N_907);
or U6636 (N_6636,N_406,N_3347);
and U6637 (N_6637,N_4876,N_1108);
xnor U6638 (N_6638,N_1896,N_5191);
xnor U6639 (N_6639,N_4426,N_1426);
nor U6640 (N_6640,N_1744,N_1567);
xnor U6641 (N_6641,N_4954,N_416);
or U6642 (N_6642,N_2797,N_307);
and U6643 (N_6643,N_2847,N_1149);
or U6644 (N_6644,N_5353,N_1088);
or U6645 (N_6645,N_5734,N_1208);
nor U6646 (N_6646,N_1131,N_1380);
nor U6647 (N_6647,N_670,N_2753);
or U6648 (N_6648,N_4086,N_2230);
or U6649 (N_6649,N_2387,N_4612);
and U6650 (N_6650,N_875,N_747);
nand U6651 (N_6651,N_585,N_6);
or U6652 (N_6652,N_1980,N_5049);
and U6653 (N_6653,N_5274,N_3156);
xnor U6654 (N_6654,N_2440,N_2072);
and U6655 (N_6655,N_1288,N_1431);
nand U6656 (N_6656,N_801,N_1178);
nor U6657 (N_6657,N_3964,N_5813);
or U6658 (N_6658,N_320,N_1370);
and U6659 (N_6659,N_2591,N_3885);
and U6660 (N_6660,N_4533,N_911);
xnor U6661 (N_6661,N_432,N_3704);
or U6662 (N_6662,N_308,N_4447);
and U6663 (N_6663,N_3437,N_618);
or U6664 (N_6664,N_3520,N_3376);
nand U6665 (N_6665,N_5216,N_2962);
nor U6666 (N_6666,N_1812,N_1049);
and U6667 (N_6667,N_5890,N_1852);
nor U6668 (N_6668,N_2988,N_1872);
nand U6669 (N_6669,N_2112,N_3607);
xnor U6670 (N_6670,N_5915,N_4912);
nor U6671 (N_6671,N_3050,N_2448);
nand U6672 (N_6672,N_1389,N_2528);
xnor U6673 (N_6673,N_5131,N_5320);
xor U6674 (N_6674,N_4351,N_5725);
and U6675 (N_6675,N_1650,N_5248);
or U6676 (N_6676,N_477,N_1497);
and U6677 (N_6677,N_198,N_2485);
nor U6678 (N_6678,N_316,N_275);
or U6679 (N_6679,N_3068,N_2863);
and U6680 (N_6680,N_112,N_1859);
nand U6681 (N_6681,N_2993,N_3511);
xnor U6682 (N_6682,N_4028,N_2531);
nor U6683 (N_6683,N_1900,N_3094);
nand U6684 (N_6684,N_4572,N_2624);
and U6685 (N_6685,N_3253,N_2855);
nor U6686 (N_6686,N_5266,N_190);
xnor U6687 (N_6687,N_28,N_701);
or U6688 (N_6688,N_2886,N_5940);
xnor U6689 (N_6689,N_4395,N_2111);
nand U6690 (N_6690,N_2587,N_3019);
or U6691 (N_6691,N_2130,N_5283);
or U6692 (N_6692,N_1591,N_2506);
xor U6693 (N_6693,N_3358,N_59);
and U6694 (N_6694,N_903,N_1670);
or U6695 (N_6695,N_3483,N_3042);
nand U6696 (N_6696,N_4995,N_2018);
xnor U6697 (N_6697,N_3757,N_4477);
nand U6698 (N_6698,N_4405,N_2295);
nand U6699 (N_6699,N_3729,N_493);
or U6700 (N_6700,N_241,N_2444);
and U6701 (N_6701,N_3715,N_2977);
nand U6702 (N_6702,N_1790,N_3328);
and U6703 (N_6703,N_4008,N_600);
nor U6704 (N_6704,N_2973,N_4285);
xnor U6705 (N_6705,N_791,N_4356);
and U6706 (N_6706,N_1749,N_152);
or U6707 (N_6707,N_3135,N_4518);
xor U6708 (N_6708,N_3413,N_3770);
nor U6709 (N_6709,N_2122,N_4484);
or U6710 (N_6710,N_567,N_5406);
or U6711 (N_6711,N_5839,N_1628);
nand U6712 (N_6712,N_3336,N_1926);
nand U6713 (N_6713,N_5990,N_1510);
or U6714 (N_6714,N_3425,N_2265);
nor U6715 (N_6715,N_2380,N_1054);
or U6716 (N_6716,N_2686,N_2236);
nand U6717 (N_6717,N_1851,N_572);
xor U6718 (N_6718,N_4259,N_3447);
xor U6719 (N_6719,N_211,N_634);
nor U6720 (N_6720,N_2949,N_3995);
or U6721 (N_6721,N_384,N_2465);
nand U6722 (N_6722,N_1486,N_5174);
nor U6723 (N_6723,N_3163,N_2373);
or U6724 (N_6724,N_3166,N_3606);
xnor U6725 (N_6725,N_5304,N_5101);
and U6726 (N_6726,N_685,N_3531);
and U6727 (N_6727,N_1765,N_1773);
xor U6728 (N_6728,N_3694,N_2963);
xor U6729 (N_6729,N_1613,N_2647);
nor U6730 (N_6730,N_2229,N_4566);
nand U6731 (N_6731,N_4391,N_2882);
nor U6732 (N_6732,N_4396,N_2106);
and U6733 (N_6733,N_2815,N_642);
nand U6734 (N_6734,N_3944,N_954);
nor U6735 (N_6735,N_4826,N_5076);
and U6736 (N_6736,N_3051,N_2051);
nor U6737 (N_6737,N_304,N_3851);
xor U6738 (N_6738,N_2107,N_4355);
nand U6739 (N_6739,N_3183,N_4233);
or U6740 (N_6740,N_1674,N_178);
nand U6741 (N_6741,N_3027,N_4765);
nor U6742 (N_6742,N_2960,N_292);
and U6743 (N_6743,N_4573,N_3962);
or U6744 (N_6744,N_4108,N_1870);
and U6745 (N_6745,N_5168,N_868);
xor U6746 (N_6746,N_472,N_1091);
xnor U6747 (N_6747,N_1685,N_4392);
nand U6748 (N_6748,N_1279,N_3001);
or U6749 (N_6749,N_5604,N_1176);
nand U6750 (N_6750,N_3992,N_2916);
and U6751 (N_6751,N_1117,N_1520);
nor U6752 (N_6752,N_3814,N_786);
xor U6753 (N_6753,N_3077,N_5397);
or U6754 (N_6754,N_770,N_3555);
or U6755 (N_6755,N_3214,N_4116);
nor U6756 (N_6756,N_3430,N_4631);
nand U6757 (N_6757,N_1592,N_5450);
and U6758 (N_6758,N_4932,N_1957);
nor U6759 (N_6759,N_2209,N_192);
nand U6760 (N_6760,N_95,N_3720);
nor U6761 (N_6761,N_4083,N_3173);
nand U6762 (N_6762,N_5806,N_4809);
nand U6763 (N_6763,N_5379,N_3266);
nand U6764 (N_6764,N_1194,N_757);
xor U6765 (N_6765,N_1528,N_942);
xor U6766 (N_6766,N_5771,N_3512);
or U6767 (N_6767,N_2889,N_3462);
nand U6768 (N_6768,N_740,N_0);
nor U6769 (N_6769,N_5284,N_1318);
or U6770 (N_6770,N_4992,N_1387);
and U6771 (N_6771,N_4282,N_3572);
nor U6772 (N_6772,N_742,N_2691);
or U6773 (N_6773,N_2294,N_4314);
or U6774 (N_6774,N_1362,N_5668);
nand U6775 (N_6775,N_3840,N_5924);
or U6776 (N_6776,N_3371,N_5763);
or U6777 (N_6777,N_5104,N_3372);
nor U6778 (N_6778,N_3164,N_5969);
nor U6779 (N_6779,N_3703,N_5531);
or U6780 (N_6780,N_3812,N_5794);
nand U6781 (N_6781,N_3975,N_5298);
xor U6782 (N_6782,N_5628,N_2839);
nand U6783 (N_6783,N_5129,N_4966);
nor U6784 (N_6784,N_4745,N_1962);
or U6785 (N_6785,N_2080,N_2081);
and U6786 (N_6786,N_2945,N_4790);
xnor U6787 (N_6787,N_1879,N_4678);
or U6788 (N_6788,N_4741,N_2737);
xnor U6789 (N_6789,N_4332,N_3732);
nor U6790 (N_6790,N_4246,N_662);
or U6791 (N_6791,N_1834,N_4748);
or U6792 (N_6792,N_4385,N_5314);
and U6793 (N_6793,N_782,N_1579);
or U6794 (N_6794,N_2430,N_4112);
xnor U6795 (N_6795,N_5046,N_4837);
or U6796 (N_6796,N_4454,N_2922);
xnor U6797 (N_6797,N_2148,N_1912);
nand U6798 (N_6798,N_3564,N_4432);
and U6799 (N_6799,N_4541,N_329);
nor U6800 (N_6800,N_837,N_2890);
or U6801 (N_6801,N_2867,N_2064);
nor U6802 (N_6802,N_4328,N_4561);
or U6803 (N_6803,N_3055,N_1802);
and U6804 (N_6804,N_568,N_3030);
and U6805 (N_6805,N_2950,N_1029);
and U6806 (N_6806,N_699,N_4677);
or U6807 (N_6807,N_1627,N_4295);
and U6808 (N_6808,N_1687,N_46);
nand U6809 (N_6809,N_5961,N_1927);
xor U6810 (N_6810,N_4865,N_419);
and U6811 (N_6811,N_983,N_3463);
or U6812 (N_6812,N_3352,N_1452);
nor U6813 (N_6813,N_1807,N_4720);
xnor U6814 (N_6814,N_958,N_3959);
nand U6815 (N_6815,N_4871,N_3435);
or U6816 (N_6816,N_4461,N_1924);
nand U6817 (N_6817,N_164,N_2914);
nand U6818 (N_6818,N_3438,N_3153);
xnor U6819 (N_6819,N_447,N_5299);
and U6820 (N_6820,N_4093,N_3028);
nor U6821 (N_6821,N_151,N_4437);
or U6822 (N_6822,N_1600,N_3535);
and U6823 (N_6823,N_575,N_4703);
xnor U6824 (N_6824,N_5966,N_5577);
or U6825 (N_6825,N_422,N_3945);
or U6826 (N_6826,N_3663,N_3127);
nand U6827 (N_6827,N_5116,N_2958);
or U6828 (N_6828,N_1397,N_5606);
and U6829 (N_6829,N_4291,N_387);
xor U6830 (N_6830,N_4976,N_805);
xor U6831 (N_6831,N_2298,N_4381);
or U6832 (N_6832,N_266,N_4851);
or U6833 (N_6833,N_3755,N_2843);
nand U6834 (N_6834,N_1247,N_1941);
nor U6835 (N_6835,N_760,N_1638);
nor U6836 (N_6836,N_4987,N_1002);
or U6837 (N_6837,N_5027,N_2241);
or U6838 (N_6838,N_5498,N_5854);
xnor U6839 (N_6839,N_5105,N_3472);
xnor U6840 (N_6840,N_1420,N_678);
and U6841 (N_6841,N_2699,N_723);
nand U6842 (N_6842,N_5305,N_4253);
or U6843 (N_6843,N_4357,N_3645);
and U6844 (N_6844,N_952,N_53);
xnor U6845 (N_6845,N_5608,N_3925);
and U6846 (N_6846,N_2841,N_4732);
and U6847 (N_6847,N_3708,N_3598);
xnor U6848 (N_6848,N_611,N_1007);
and U6849 (N_6849,N_1501,N_5889);
xnor U6850 (N_6850,N_5439,N_1967);
nand U6851 (N_6851,N_2540,N_102);
or U6852 (N_6852,N_3444,N_5917);
or U6853 (N_6853,N_1602,N_1641);
nand U6854 (N_6854,N_3633,N_5043);
or U6855 (N_6855,N_1801,N_726);
or U6856 (N_6856,N_5782,N_851);
or U6857 (N_6857,N_5530,N_5546);
nand U6858 (N_6858,N_626,N_1562);
nand U6859 (N_6859,N_1711,N_3827);
nor U6860 (N_6860,N_3470,N_4309);
nor U6861 (N_6861,N_3862,N_2664);
nor U6862 (N_6862,N_37,N_4761);
xnor U6863 (N_6863,N_4456,N_1161);
xor U6864 (N_6864,N_2003,N_368);
or U6865 (N_6865,N_2210,N_1909);
nand U6866 (N_6866,N_5929,N_3505);
xnor U6867 (N_6867,N_3583,N_9);
nand U6868 (N_6868,N_521,N_3385);
nand U6869 (N_6869,N_2493,N_4486);
nor U6870 (N_6870,N_2364,N_2220);
xnor U6871 (N_6871,N_4097,N_1280);
and U6872 (N_6872,N_3024,N_1654);
or U6873 (N_6873,N_3563,N_2142);
or U6874 (N_6874,N_5790,N_5963);
xnor U6875 (N_6875,N_5190,N_1269);
and U6876 (N_6876,N_4699,N_2207);
nor U6877 (N_6877,N_1095,N_5891);
or U6878 (N_6878,N_5000,N_153);
nand U6879 (N_6879,N_515,N_5622);
nor U6880 (N_6880,N_3699,N_221);
nand U6881 (N_6881,N_951,N_5011);
nand U6882 (N_6882,N_4179,N_3205);
nand U6883 (N_6883,N_3017,N_1232);
xor U6884 (N_6884,N_643,N_2978);
xnor U6885 (N_6885,N_5313,N_1434);
nor U6886 (N_6886,N_2473,N_2798);
and U6887 (N_6887,N_4630,N_5798);
and U6888 (N_6888,N_5311,N_3061);
and U6889 (N_6889,N_2734,N_5403);
nor U6890 (N_6890,N_2321,N_3655);
nand U6891 (N_6891,N_5005,N_1521);
xor U6892 (N_6892,N_5188,N_4213);
and U6893 (N_6893,N_5686,N_3080);
nand U6894 (N_6894,N_1129,N_2766);
xor U6895 (N_6895,N_5386,N_4127);
nand U6896 (N_6896,N_30,N_2518);
nor U6897 (N_6897,N_2441,N_2807);
nand U6898 (N_6898,N_4240,N_3048);
nor U6899 (N_6899,N_1133,N_461);
xnor U6900 (N_6900,N_1548,N_2384);
or U6901 (N_6901,N_4742,N_4199);
or U6902 (N_6902,N_2305,N_582);
or U6903 (N_6903,N_2116,N_3393);
and U6904 (N_6904,N_707,N_3264);
nor U6905 (N_6905,N_5426,N_397);
nand U6906 (N_6906,N_2549,N_5474);
and U6907 (N_6907,N_1062,N_3902);
xnor U6908 (N_6908,N_197,N_2641);
and U6909 (N_6909,N_1624,N_4378);
nand U6910 (N_6910,N_2019,N_78);
and U6911 (N_6911,N_5921,N_3832);
and U6912 (N_6912,N_5874,N_2551);
xor U6913 (N_6913,N_5071,N_1213);
nand U6914 (N_6914,N_4807,N_2951);
nand U6915 (N_6915,N_3603,N_5289);
xnor U6916 (N_6916,N_5262,N_452);
xnor U6917 (N_6917,N_799,N_1706);
nor U6918 (N_6918,N_2233,N_4766);
xnor U6919 (N_6919,N_3184,N_4433);
or U6920 (N_6920,N_2022,N_2325);
nand U6921 (N_6921,N_5067,N_4443);
or U6922 (N_6922,N_4743,N_2310);
nor U6923 (N_6923,N_5219,N_3553);
nand U6924 (N_6924,N_4867,N_3339);
and U6925 (N_6925,N_896,N_4978);
xnor U6926 (N_6926,N_3479,N_3875);
xnor U6927 (N_6927,N_649,N_4414);
or U6928 (N_6928,N_4248,N_3054);
xnor U6929 (N_6929,N_3676,N_4933);
nor U6930 (N_6930,N_258,N_147);
xor U6931 (N_6931,N_2078,N_2846);
nand U6932 (N_6932,N_3618,N_1594);
nand U6933 (N_6933,N_3652,N_3842);
nor U6934 (N_6934,N_681,N_3442);
or U6935 (N_6935,N_5938,N_4900);
xor U6936 (N_6936,N_3808,N_1599);
nand U6937 (N_6937,N_5041,N_4348);
nand U6938 (N_6938,N_4054,N_4201);
xor U6939 (N_6939,N_1786,N_2423);
and U6940 (N_6940,N_5584,N_4854);
and U6941 (N_6941,N_3736,N_941);
xor U6942 (N_6942,N_4136,N_2330);
or U6943 (N_6943,N_2311,N_1052);
nand U6944 (N_6944,N_4994,N_5594);
and U6945 (N_6945,N_857,N_3238);
and U6946 (N_6946,N_83,N_4010);
nand U6947 (N_6947,N_3332,N_3377);
or U6948 (N_6948,N_2357,N_1076);
xor U6949 (N_6949,N_3948,N_4390);
nand U6950 (N_6950,N_1649,N_4668);
or U6951 (N_6951,N_3428,N_2661);
or U6952 (N_6952,N_5821,N_1959);
or U6953 (N_6953,N_142,N_5995);
nor U6954 (N_6954,N_2804,N_3630);
or U6955 (N_6955,N_4088,N_722);
xnor U6956 (N_6956,N_4799,N_4506);
nand U6957 (N_6957,N_3724,N_4084);
xnor U6958 (N_6958,N_2568,N_1971);
and U6959 (N_6959,N_5198,N_5271);
or U6960 (N_6960,N_883,N_4661);
and U6961 (N_6961,N_3918,N_2369);
and U6962 (N_6962,N_908,N_943);
xnor U6963 (N_6963,N_1238,N_3198);
or U6964 (N_6964,N_1139,N_1359);
or U6965 (N_6965,N_5587,N_1413);
nor U6966 (N_6966,N_4567,N_2098);
and U6967 (N_6967,N_5390,N_4820);
and U6968 (N_6968,N_691,N_3809);
nand U6969 (N_6969,N_1313,N_63);
nand U6970 (N_6970,N_3036,N_817);
nor U6971 (N_6971,N_3994,N_5641);
nor U6972 (N_6972,N_2176,N_5754);
nor U6973 (N_6973,N_4455,N_2302);
nand U6974 (N_6974,N_4389,N_3467);
nand U6975 (N_6975,N_1827,N_4650);
nand U6976 (N_6976,N_5030,N_4459);
and U6977 (N_6977,N_1157,N_5087);
nor U6978 (N_6978,N_2431,N_4299);
nor U6979 (N_6979,N_3005,N_4012);
xnor U6980 (N_6980,N_3222,N_3225);
nor U6981 (N_6981,N_3414,N_635);
or U6982 (N_6982,N_1067,N_4264);
xor U6983 (N_6983,N_5324,N_5045);
nand U6984 (N_6984,N_1097,N_448);
xnor U6985 (N_6985,N_4262,N_322);
xnor U6986 (N_6986,N_3180,N_1055);
and U6987 (N_6987,N_2066,N_2110);
nor U6988 (N_6988,N_4060,N_593);
or U6989 (N_6989,N_284,N_17);
nor U6990 (N_6990,N_5581,N_858);
nand U6991 (N_6991,N_1298,N_2635);
xnor U6992 (N_6992,N_2981,N_4067);
nor U6993 (N_6993,N_838,N_881);
or U6994 (N_6994,N_4493,N_1045);
nand U6995 (N_6995,N_860,N_2966);
nand U6996 (N_6996,N_732,N_2599);
nand U6997 (N_6997,N_2595,N_4928);
and U6998 (N_6998,N_2913,N_2842);
and U6999 (N_6999,N_3286,N_3227);
nand U7000 (N_7000,N_3710,N_5828);
or U7001 (N_7001,N_1135,N_890);
nand U7002 (N_7002,N_4618,N_1240);
nand U7003 (N_7003,N_5098,N_1557);
nand U7004 (N_7004,N_3075,N_460);
nor U7005 (N_7005,N_3763,N_5343);
nor U7006 (N_7006,N_4031,N_3569);
xnor U7007 (N_7007,N_712,N_2350);
or U7008 (N_7008,N_5967,N_1489);
nor U7009 (N_7009,N_5066,N_3058);
xnor U7010 (N_7010,N_5016,N_467);
or U7011 (N_7011,N_1696,N_3805);
xor U7012 (N_7012,N_1300,N_386);
or U7013 (N_7013,N_5977,N_2619);
and U7014 (N_7014,N_902,N_3877);
or U7015 (N_7015,N_5136,N_1817);
nor U7016 (N_7016,N_5785,N_5720);
nor U7017 (N_7017,N_583,N_1951);
nand U7018 (N_7018,N_5059,N_5169);
xnor U7019 (N_7019,N_5861,N_4943);
nand U7020 (N_7020,N_2794,N_3584);
and U7021 (N_7021,N_5539,N_1023);
and U7022 (N_7022,N_4709,N_5024);
nor U7023 (N_7023,N_2457,N_3065);
xor U7024 (N_7024,N_456,N_4665);
xnor U7025 (N_7025,N_1988,N_2212);
nor U7026 (N_7026,N_3744,N_5548);
xor U7027 (N_7027,N_865,N_4265);
nor U7028 (N_7028,N_4270,N_1152);
and U7029 (N_7029,N_1016,N_4363);
xnor U7030 (N_7030,N_562,N_2);
or U7031 (N_7031,N_5241,N_1697);
xnor U7032 (N_7032,N_5930,N_1584);
nor U7033 (N_7033,N_3646,N_35);
nor U7034 (N_7034,N_3590,N_1758);
and U7035 (N_7035,N_5475,N_4244);
nand U7036 (N_7036,N_1612,N_3717);
xnor U7037 (N_7037,N_5447,N_4403);
nor U7038 (N_7038,N_3973,N_4072);
and U7039 (N_7039,N_5480,N_731);
nand U7040 (N_7040,N_5662,N_5791);
and U7041 (N_7041,N_2124,N_4267);
xnor U7042 (N_7042,N_2038,N_708);
nand U7043 (N_7043,N_2745,N_4939);
xnor U7044 (N_7044,N_365,N_4694);
and U7045 (N_7045,N_1198,N_4058);
nor U7046 (N_7046,N_3552,N_5183);
or U7047 (N_7047,N_3702,N_476);
or U7048 (N_7048,N_3795,N_5614);
or U7049 (N_7049,N_1480,N_2073);
or U7050 (N_7050,N_7,N_5514);
nor U7051 (N_7051,N_1138,N_4918);
nand U7052 (N_7052,N_5309,N_173);
nor U7053 (N_7053,N_2250,N_5774);
xnor U7054 (N_7054,N_2056,N_853);
nand U7055 (N_7055,N_1058,N_5710);
xnor U7056 (N_7056,N_107,N_1295);
and U7057 (N_7057,N_779,N_1992);
nand U7058 (N_7058,N_4339,N_563);
nor U7059 (N_7059,N_1124,N_3781);
and U7060 (N_7060,N_3825,N_127);
xor U7061 (N_7061,N_2399,N_136);
xnor U7062 (N_7062,N_302,N_3243);
and U7063 (N_7063,N_1,N_2316);
and U7064 (N_7064,N_4829,N_2354);
xor U7065 (N_7065,N_5665,N_4284);
xnor U7066 (N_7066,N_3070,N_3739);
nor U7067 (N_7067,N_1069,N_5857);
or U7068 (N_7068,N_844,N_5170);
xnor U7069 (N_7069,N_2679,N_2404);
xor U7070 (N_7070,N_4662,N_2840);
nand U7071 (N_7071,N_5224,N_1070);
or U7072 (N_7072,N_4585,N_4640);
and U7073 (N_7073,N_3143,N_2393);
or U7074 (N_7074,N_5141,N_1044);
xnor U7075 (N_7075,N_5143,N_4338);
nand U7076 (N_7076,N_2511,N_271);
nor U7077 (N_7077,N_5401,N_2147);
nor U7078 (N_7078,N_3436,N_4521);
nor U7079 (N_7079,N_2370,N_5521);
xor U7080 (N_7080,N_4916,N_3281);
xnor U7081 (N_7081,N_2031,N_3121);
or U7082 (N_7082,N_84,N_3417);
or U7083 (N_7083,N_3105,N_1090);
nor U7084 (N_7084,N_115,N_4077);
xor U7085 (N_7085,N_4516,N_2536);
nand U7086 (N_7086,N_664,N_3452);
nor U7087 (N_7087,N_5566,N_5479);
nand U7088 (N_7088,N_3132,N_3341);
or U7089 (N_7089,N_4513,N_2974);
or U7090 (N_7090,N_2037,N_2872);
nand U7091 (N_7091,N_212,N_5265);
nor U7092 (N_7092,N_5074,N_5925);
nand U7093 (N_7093,N_754,N_1284);
nor U7094 (N_7094,N_3698,N_1004);
or U7095 (N_7095,N_3448,N_4409);
nand U7096 (N_7096,N_2923,N_1829);
nand U7097 (N_7097,N_2642,N_532);
and U7098 (N_7098,N_4590,N_4343);
and U7099 (N_7099,N_3031,N_5211);
or U7100 (N_7100,N_44,N_5996);
nand U7101 (N_7101,N_3379,N_516);
and U7102 (N_7102,N_1057,N_3869);
and U7103 (N_7103,N_1856,N_2090);
nand U7104 (N_7104,N_3522,N_217);
and U7105 (N_7105,N_739,N_4569);
nand U7106 (N_7106,N_4804,N_2450);
or U7107 (N_7107,N_928,N_261);
or U7108 (N_7108,N_5399,N_2043);
nand U7109 (N_7109,N_2908,N_5411);
or U7110 (N_7110,N_2392,N_4273);
xor U7111 (N_7111,N_5656,N_1432);
nor U7112 (N_7112,N_4050,N_4446);
nand U7113 (N_7113,N_3103,N_1368);
nor U7114 (N_7114,N_5250,N_4786);
and U7115 (N_7115,N_227,N_2252);
nand U7116 (N_7116,N_404,N_1100);
and U7117 (N_7117,N_3831,N_4485);
nor U7118 (N_7118,N_571,N_256);
xor U7119 (N_7119,N_1268,N_3559);
or U7120 (N_7120,N_4655,N_2810);
nand U7121 (N_7121,N_5303,N_5541);
nand U7122 (N_7122,N_2061,N_2590);
nand U7123 (N_7123,N_3562,N_4942);
or U7124 (N_7124,N_3460,N_2127);
and U7125 (N_7125,N_5980,N_2347);
nand U7126 (N_7126,N_5157,N_2920);
or U7127 (N_7127,N_2360,N_200);
xor U7128 (N_7128,N_1731,N_2062);
nand U7129 (N_7129,N_297,N_3141);
nand U7130 (N_7130,N_1754,N_5916);
nand U7131 (N_7131,N_2736,N_2887);
nor U7132 (N_7132,N_25,N_706);
or U7133 (N_7133,N_4610,N_3378);
nand U7134 (N_7134,N_5372,N_3443);
or U7135 (N_7135,N_3000,N_3539);
xor U7136 (N_7136,N_734,N_183);
and U7137 (N_7137,N_2852,N_2278);
or U7138 (N_7138,N_1424,N_10);
or U7139 (N_7139,N_5452,N_2343);
or U7140 (N_7140,N_3165,N_2748);
nor U7141 (N_7141,N_580,N_846);
and U7142 (N_7142,N_3605,N_2407);
nor U7143 (N_7143,N_5235,N_2475);
and U7144 (N_7144,N_3310,N_2032);
xnor U7145 (N_7145,N_2714,N_155);
or U7146 (N_7146,N_4539,N_3230);
nor U7147 (N_7147,N_867,N_4428);
nor U7148 (N_7148,N_2541,N_411);
or U7149 (N_7149,N_1210,N_2477);
and U7150 (N_7150,N_1018,N_2345);
nor U7151 (N_7151,N_2597,N_5717);
xnor U7152 (N_7152,N_4981,N_3283);
or U7153 (N_7153,N_5206,N_2791);
nor U7154 (N_7154,N_4639,N_5728);
or U7155 (N_7155,N_420,N_4643);
or U7156 (N_7156,N_2245,N_1451);
or U7157 (N_7157,N_3957,N_4472);
and U7158 (N_7158,N_2445,N_2301);
nor U7159 (N_7159,N_2292,N_5135);
xnor U7160 (N_7160,N_5058,N_4305);
xor U7161 (N_7161,N_4646,N_2694);
or U7162 (N_7162,N_1179,N_4057);
and U7163 (N_7163,N_4746,N_3278);
nor U7164 (N_7164,N_1372,N_4840);
nor U7165 (N_7165,N_3557,N_5173);
nand U7166 (N_7166,N_3788,N_4044);
nand U7167 (N_7167,N_4903,N_24);
nor U7168 (N_7168,N_949,N_4360);
xnor U7169 (N_7169,N_1092,N_506);
nand U7170 (N_7170,N_1897,N_4580);
or U7171 (N_7171,N_1678,N_1643);
nor U7172 (N_7172,N_2361,N_2414);
or U7173 (N_7173,N_3760,N_3987);
xnor U7174 (N_7174,N_979,N_2283);
and U7175 (N_7175,N_5743,N_4666);
or U7176 (N_7176,N_4894,N_2355);
and U7177 (N_7177,N_3881,N_1844);
nor U7178 (N_7178,N_5505,N_5457);
xor U7179 (N_7179,N_5264,N_3049);
nand U7180 (N_7180,N_2650,N_1518);
and U7181 (N_7181,N_62,N_2458);
nand U7182 (N_7182,N_3599,N_5786);
xor U7183 (N_7183,N_886,N_4025);
nor U7184 (N_7184,N_1273,N_1701);
xor U7185 (N_7185,N_1321,N_2324);
and U7186 (N_7186,N_1853,N_887);
nand U7187 (N_7187,N_1882,N_5840);
xnor U7188 (N_7188,N_5356,N_1785);
or U7189 (N_7189,N_1472,N_5804);
and U7190 (N_7190,N_1767,N_3139);
or U7191 (N_7191,N_2596,N_5700);
nand U7192 (N_7192,N_998,N_4350);
nand U7193 (N_7193,N_2724,N_5745);
nor U7194 (N_7194,N_4335,N_1467);
xor U7195 (N_7195,N_986,N_1969);
or U7196 (N_7196,N_1065,N_22);
nor U7197 (N_7197,N_3056,N_2480);
xnor U7198 (N_7198,N_1401,N_269);
nand U7199 (N_7199,N_4434,N_5533);
and U7200 (N_7200,N_4570,N_1123);
xnor U7201 (N_7201,N_1950,N_1707);
nor U7202 (N_7202,N_2016,N_1960);
and U7203 (N_7203,N_5807,N_21);
nor U7204 (N_7204,N_385,N_2983);
and U7205 (N_7205,N_5981,N_3007);
nand U7206 (N_7206,N_5122,N_1050);
and U7207 (N_7207,N_5626,N_1461);
nor U7208 (N_7208,N_751,N_5291);
nand U7209 (N_7209,N_2149,N_2948);
xnor U7210 (N_7210,N_3996,N_1439);
xor U7211 (N_7211,N_3797,N_4200);
and U7212 (N_7212,N_2434,N_4984);
nand U7213 (N_7213,N_4638,N_3916);
xor U7214 (N_7214,N_5811,N_2690);
xnor U7215 (N_7215,N_539,N_4982);
nand U7216 (N_7216,N_1344,N_1523);
nor U7217 (N_7217,N_4975,N_279);
and U7218 (N_7218,N_2869,N_5312);
or U7219 (N_7219,N_3837,N_1122);
and U7220 (N_7220,N_2367,N_627);
nor U7221 (N_7221,N_4330,N_2555);
and U7222 (N_7222,N_5204,N_5697);
or U7223 (N_7223,N_5752,N_5948);
xor U7224 (N_7224,N_4996,N_4347);
xor U7225 (N_7225,N_3186,N_3390);
or U7226 (N_7226,N_1517,N_3333);
nor U7227 (N_7227,N_5586,N_804);
xnor U7228 (N_7228,N_4819,N_4560);
nor U7229 (N_7229,N_5905,N_5179);
and U7230 (N_7230,N_4036,N_4739);
xnor U7231 (N_7231,N_3043,N_1388);
or U7232 (N_7232,N_1672,N_3471);
and U7233 (N_7233,N_4165,N_2424);
xor U7234 (N_7234,N_215,N_3315);
nand U7235 (N_7235,N_5115,N_364);
xor U7236 (N_7236,N_1484,N_891);
xor U7237 (N_7237,N_2328,N_2614);
nor U7238 (N_7238,N_69,N_3638);
and U7239 (N_7239,N_1249,N_5348);
or U7240 (N_7240,N_4232,N_2765);
xor U7241 (N_7241,N_106,N_5329);
nand U7242 (N_7242,N_1652,N_1328);
xor U7243 (N_7243,N_4509,N_1740);
or U7244 (N_7244,N_5364,N_3890);
and U7245 (N_7245,N_1219,N_4555);
and U7246 (N_7246,N_727,N_3748);
or U7247 (N_7247,N_5079,N_4346);
or U7248 (N_7248,N_4212,N_3147);
nor U7249 (N_7249,N_1795,N_3237);
xnor U7250 (N_7250,N_2582,N_4692);
nor U7251 (N_7251,N_5809,N_4052);
or U7252 (N_7252,N_5357,N_3136);
or U7253 (N_7253,N_663,N_2939);
nor U7254 (N_7254,N_5220,N_2126);
nand U7255 (N_7255,N_303,N_214);
or U7256 (N_7256,N_2668,N_1686);
nand U7257 (N_7257,N_1708,N_3223);
and U7258 (N_7258,N_1234,N_3307);
nand U7259 (N_7259,N_775,N_4051);
or U7260 (N_7260,N_3265,N_1824);
nand U7261 (N_7261,N_5275,N_3856);
or U7262 (N_7262,N_5788,N_1692);
nand U7263 (N_7263,N_5155,N_5369);
nor U7264 (N_7264,N_1887,N_2436);
or U7265 (N_7265,N_4276,N_2170);
nand U7266 (N_7266,N_5483,N_717);
xnor U7267 (N_7267,N_5095,N_1286);
and U7268 (N_7268,N_3192,N_4120);
and U7269 (N_7269,N_1101,N_1366);
nand U7270 (N_7270,N_4149,N_4767);
and U7271 (N_7271,N_4130,N_5761);
xor U7272 (N_7272,N_205,N_1846);
nand U7273 (N_7273,N_2388,N_2517);
and U7274 (N_7274,N_4085,N_2188);
xnor U7275 (N_7275,N_5292,N_5003);
nor U7276 (N_7276,N_1482,N_2255);
and U7277 (N_7277,N_2291,N_5226);
or U7278 (N_7278,N_3938,N_501);
and U7279 (N_7279,N_3639,N_4497);
nand U7280 (N_7280,N_4552,N_5630);
and U7281 (N_7281,N_5884,N_1793);
and U7282 (N_7282,N_5859,N_1761);
nor U7283 (N_7283,N_2181,N_651);
nand U7284 (N_7284,N_2503,N_2284);
and U7285 (N_7285,N_5764,N_298);
nand U7286 (N_7286,N_237,N_4985);
xor U7287 (N_7287,N_2788,N_5534);
nand U7288 (N_7288,N_2996,N_948);
or U7289 (N_7289,N_3919,N_4181);
or U7290 (N_7290,N_1425,N_4917);
xor U7291 (N_7291,N_1075,N_3524);
xnor U7292 (N_7292,N_1883,N_2421);
or U7293 (N_7293,N_2123,N_4145);
or U7294 (N_7294,N_1172,N_1074);
xnor U7295 (N_7295,N_2119,N_725);
nor U7296 (N_7296,N_4310,N_5080);
xor U7297 (N_7297,N_5199,N_3380);
nand U7298 (N_7298,N_5522,N_2497);
nand U7299 (N_7299,N_1335,N_438);
or U7300 (N_7300,N_1418,N_2726);
nand U7301 (N_7301,N_3560,N_1185);
nand U7302 (N_7302,N_3870,N_3035);
xnor U7303 (N_7303,N_1206,N_1804);
nor U7304 (N_7304,N_380,N_752);
or U7305 (N_7305,N_1865,N_5635);
xor U7306 (N_7306,N_4811,N_2813);
xor U7307 (N_7307,N_281,N_711);
xnor U7308 (N_7308,N_1512,N_4553);
nor U7309 (N_7309,N_296,N_4117);
xor U7310 (N_7310,N_270,N_541);
or U7311 (N_7311,N_5384,N_5617);
and U7312 (N_7312,N_4598,N_4173);
nor U7313 (N_7313,N_4551,N_1306);
and U7314 (N_7314,N_3045,N_1519);
nor U7315 (N_7315,N_60,N_5200);
or U7316 (N_7316,N_2290,N_4625);
nand U7317 (N_7317,N_1046,N_3411);
nor U7318 (N_7318,N_4959,N_2128);
nand U7319 (N_7319,N_4735,N_5381);
xnor U7320 (N_7320,N_2885,N_4436);
and U7321 (N_7321,N_2084,N_1008);
and U7322 (N_7322,N_3285,N_821);
nor U7323 (N_7323,N_4279,N_3224);
or U7324 (N_7324,N_3714,N_4863);
nor U7325 (N_7325,N_2984,N_3548);
xor U7326 (N_7326,N_4009,N_1634);
xnor U7327 (N_7327,N_2761,N_3971);
nor U7328 (N_7328,N_1880,N_3006);
or U7329 (N_7329,N_864,N_2529);
or U7330 (N_7330,N_3643,N_4581);
nor U7331 (N_7331,N_947,N_1588);
nand U7332 (N_7332,N_2953,N_4466);
nor U7333 (N_7333,N_780,N_3614);
or U7334 (N_7334,N_2688,N_5307);
nand U7335 (N_7335,N_441,N_4956);
nor U7336 (N_7336,N_3853,N_3747);
xnor U7337 (N_7337,N_5768,N_4404);
or U7338 (N_7338,N_352,N_1947);
or U7339 (N_7339,N_5909,N_2366);
and U7340 (N_7340,N_518,N_3629);
and U7341 (N_7341,N_187,N_5649);
nand U7342 (N_7342,N_3530,N_748);
or U7343 (N_7343,N_4821,N_2164);
or U7344 (N_7344,N_4507,N_4548);
or U7345 (N_7345,N_2001,N_1151);
xor U7346 (N_7346,N_118,N_598);
or U7347 (N_7347,N_3947,N_5001);
xor U7348 (N_7348,N_4624,N_5557);
and U7349 (N_7349,N_496,N_1031);
and U7350 (N_7350,N_2758,N_1698);
or U7351 (N_7351,N_1782,N_1843);
or U7352 (N_7352,N_1626,N_82);
xor U7353 (N_7353,N_3966,N_475);
nand U7354 (N_7354,N_5257,N_2059);
nor U7355 (N_7355,N_524,N_3251);
or U7356 (N_7356,N_3003,N_5112);
or U7357 (N_7357,N_5371,N_3388);
or U7358 (N_7358,N_1667,N_4229);
nor U7359 (N_7359,N_5696,N_334);
nand U7360 (N_7360,N_4796,N_100);
xnor U7361 (N_7361,N_2617,N_4490);
and U7362 (N_7362,N_4388,N_981);
or U7363 (N_7363,N_679,N_768);
xor U7364 (N_7364,N_2163,N_3543);
xor U7365 (N_7365,N_97,N_5607);
nor U7366 (N_7366,N_4269,N_343);
or U7367 (N_7367,N_2546,N_5860);
nand U7368 (N_7368,N_3813,N_435);
and U7369 (N_7369,N_705,N_105);
nand U7370 (N_7370,N_1361,N_5645);
xor U7371 (N_7371,N_3866,N_5044);
nand U7372 (N_7372,N_5694,N_5454);
xnor U7373 (N_7373,N_2285,N_4974);
nor U7374 (N_7374,N_2615,N_721);
nor U7375 (N_7375,N_161,N_813);
nand U7376 (N_7376,N_5723,N_117);
and U7377 (N_7377,N_5877,N_5825);
nor U7378 (N_7378,N_688,N_3256);
xnor U7379 (N_7379,N_4724,N_5302);
xor U7380 (N_7380,N_3365,N_3846);
and U7381 (N_7381,N_3775,N_2820);
and U7382 (N_7382,N_5352,N_1043);
nand U7383 (N_7383,N_5580,N_4704);
and U7384 (N_7384,N_2554,N_5544);
nor U7385 (N_7385,N_2771,N_845);
and U7386 (N_7386,N_1275,N_5515);
or U7387 (N_7387,N_2484,N_272);
nor U7388 (N_7388,N_2700,N_5459);
nand U7389 (N_7389,N_2575,N_1457);
nand U7390 (N_7390,N_4642,N_263);
nand U7391 (N_7391,N_2033,N_540);
nand U7392 (N_7392,N_4331,N_5111);
nand U7393 (N_7393,N_940,N_997);
and U7394 (N_7394,N_5404,N_835);
nand U7395 (N_7395,N_5919,N_3305);
nand U7396 (N_7396,N_2470,N_1858);
or U7397 (N_7397,N_1822,N_5236);
or U7398 (N_7398,N_4899,N_4245);
nor U7399 (N_7399,N_3785,N_191);
or U7400 (N_7400,N_3120,N_4595);
and U7401 (N_7401,N_5336,N_1500);
xor U7402 (N_7402,N_33,N_4397);
nor U7403 (N_7403,N_5181,N_2348);
xnor U7404 (N_7404,N_1068,N_5893);
xnor U7405 (N_7405,N_5321,N_2520);
or U7406 (N_7406,N_2895,N_1968);
or U7407 (N_7407,N_3229,N_2463);
and U7408 (N_7408,N_403,N_622);
nand U7409 (N_7409,N_1003,N_1884);
nand U7410 (N_7410,N_4386,N_557);
and U7411 (N_7411,N_2573,N_3268);
and U7412 (N_7412,N_2218,N_4468);
or U7413 (N_7413,N_4923,N_5959);
nor U7414 (N_7414,N_1554,N_633);
or U7415 (N_7415,N_2927,N_4369);
nor U7416 (N_7416,N_5853,N_4778);
nor U7417 (N_7417,N_4924,N_901);
nor U7418 (N_7418,N_3155,N_2925);
nand U7419 (N_7419,N_4802,N_657);
xnor U7420 (N_7420,N_5422,N_4019);
nor U7421 (N_7421,N_5006,N_3923);
and U7422 (N_7422,N_772,N_3203);
nand U7423 (N_7423,N_709,N_20);
nor U7424 (N_7424,N_3644,N_3273);
and U7425 (N_7425,N_5766,N_2415);
and U7426 (N_7426,N_3484,N_926);
and U7427 (N_7427,N_3723,N_1416);
nand U7428 (N_7428,N_5918,N_5927);
xor U7429 (N_7429,N_1441,N_305);
xnor U7430 (N_7430,N_2095,N_5036);
and U7431 (N_7431,N_620,N_2074);
xor U7432 (N_7432,N_1287,N_160);
or U7433 (N_7433,N_2400,N_5778);
nand U7434 (N_7434,N_464,N_5690);
or U7435 (N_7435,N_4382,N_3792);
nor U7436 (N_7436,N_3933,N_3491);
xnor U7437 (N_7437,N_4702,N_1720);
or U7438 (N_7438,N_1820,N_1290);
xor U7439 (N_7439,N_3255,N_741);
xor U7440 (N_7440,N_4731,N_5643);
xor U7441 (N_7441,N_5601,N_975);
xor U7442 (N_7442,N_1187,N_2703);
nor U7443 (N_7443,N_3984,N_3025);
nor U7444 (N_7444,N_268,N_724);
xor U7445 (N_7445,N_3601,N_5896);
nor U7446 (N_7446,N_764,N_5563);
xnor U7447 (N_7447,N_2083,N_669);
nand U7448 (N_7448,N_653,N_5050);
or U7449 (N_7449,N_5009,N_1020);
or U7450 (N_7450,N_3735,N_4055);
nand U7451 (N_7451,N_2743,N_637);
and U7452 (N_7452,N_2713,N_2488);
nand U7453 (N_7453,N_4841,N_4372);
or U7454 (N_7454,N_1989,N_4307);
and U7455 (N_7455,N_2137,N_2621);
nand U7456 (N_7456,N_4801,N_4368);
or U7457 (N_7457,N_2491,N_2267);
nor U7458 (N_7458,N_430,N_3958);
or U7459 (N_7459,N_1053,N_2069);
nor U7460 (N_7460,N_480,N_2937);
nand U7461 (N_7461,N_5576,N_3236);
or U7462 (N_7462,N_4591,N_1225);
or U7463 (N_7463,N_1471,N_3326);
and U7464 (N_7464,N_2629,N_4241);
and U7465 (N_7465,N_3097,N_1757);
nor U7466 (N_7466,N_5715,N_3039);
and U7467 (N_7467,N_802,N_4480);
and U7468 (N_7468,N_4947,N_3817);
xor U7469 (N_7469,N_519,N_1772);
and U7470 (N_7470,N_893,N_3773);
or U7471 (N_7471,N_3686,N_1180);
nor U7472 (N_7472,N_209,N_5741);
xor U7473 (N_7473,N_2159,N_3997);
or U7474 (N_7474,N_5997,N_1901);
nor U7475 (N_7475,N_2739,N_4708);
xnor U7476 (N_7476,N_3623,N_1633);
nor U7477 (N_7477,N_2416,N_3976);
nand U7478 (N_7478,N_3701,N_3910);
nor U7479 (N_7479,N_333,N_5118);
nand U7480 (N_7480,N_3591,N_2372);
nor U7481 (N_7481,N_2821,N_1233);
nor U7482 (N_7482,N_3573,N_3980);
nand U7483 (N_7483,N_1938,N_2318);
nor U7484 (N_7484,N_2658,N_2190);
nor U7485 (N_7485,N_1205,N_5213);
xor U7486 (N_7486,N_1918,N_4636);
xor U7487 (N_7487,N_1877,N_5391);
or U7488 (N_7488,N_5424,N_579);
or U7489 (N_7489,N_4049,N_2133);
nand U7490 (N_7490,N_3434,N_4961);
or U7491 (N_7491,N_149,N_442);
nand U7492 (N_7492,N_3178,N_40);
xor U7493 (N_7493,N_1449,N_1182);
and U7494 (N_7494,N_2192,N_4487);
nand U7495 (N_7495,N_3602,N_3179);
nand U7496 (N_7496,N_1156,N_1866);
or U7497 (N_7497,N_3597,N_494);
nand U7498 (N_7498,N_2406,N_2044);
or U7499 (N_7499,N_5692,N_4020);
xnor U7500 (N_7500,N_3033,N_5394);
nor U7501 (N_7501,N_193,N_3220);
xnor U7502 (N_7502,N_5315,N_5218);
xor U7503 (N_7503,N_776,N_1118);
nor U7504 (N_7504,N_1538,N_372);
xor U7505 (N_7505,N_2139,N_4536);
xnor U7506 (N_7506,N_4413,N_4705);
nor U7507 (N_7507,N_5750,N_2332);
or U7508 (N_7508,N_2654,N_4814);
nor U7509 (N_7509,N_3182,N_1746);
nand U7510 (N_7510,N_3922,N_2663);
or U7511 (N_7511,N_730,N_3368);
nand U7512 (N_7512,N_1028,N_1014);
nand U7513 (N_7513,N_4712,N_3324);
nor U7514 (N_7514,N_4224,N_3441);
nor U7515 (N_7515,N_285,N_5585);
nand U7516 (N_7516,N_5355,N_1535);
or U7517 (N_7517,N_1504,N_1534);
and U7518 (N_7518,N_5297,N_1723);
and U7519 (N_7519,N_5532,N_1981);
nand U7520 (N_7520,N_3468,N_3778);
and U7521 (N_7521,N_5873,N_2959);
nor U7522 (N_7522,N_1577,N_1032);
nand U7523 (N_7523,N_49,N_3667);
or U7524 (N_7524,N_2955,N_154);
and U7525 (N_7525,N_900,N_2891);
and U7526 (N_7526,N_3496,N_2070);
nor U7527 (N_7527,N_1371,N_668);
nor U7528 (N_7528,N_1305,N_5620);
xor U7529 (N_7529,N_2594,N_96);
and U7530 (N_7530,N_5360,N_1775);
nand U7531 (N_7531,N_4326,N_5140);
nor U7532 (N_7532,N_3683,N_3546);
or U7533 (N_7533,N_1755,N_4207);
nand U7534 (N_7534,N_328,N_2519);
nand U7535 (N_7535,N_4834,N_1173);
xnor U7536 (N_7536,N_2780,N_3541);
nand U7537 (N_7537,N_4637,N_5669);
nand U7538 (N_7538,N_3806,N_3600);
xor U7539 (N_7539,N_2747,N_5847);
nor U7540 (N_7540,N_3516,N_2751);
and U7541 (N_7541,N_3841,N_3293);
and U7542 (N_7542,N_4105,N_4651);
or U7543 (N_7543,N_4697,N_5625);
or U7544 (N_7544,N_5691,N_4608);
nor U7545 (N_7545,N_3053,N_1842);
and U7546 (N_7546,N_3807,N_773);
xnor U7547 (N_7547,N_282,N_4914);
nor U7548 (N_7548,N_1714,N_4169);
nand U7549 (N_7549,N_2787,N_1098);
xor U7550 (N_7550,N_1071,N_2274);
or U7551 (N_7551,N_4124,N_408);
nand U7552 (N_7552,N_2408,N_1864);
and U7553 (N_7553,N_5992,N_2957);
nand U7554 (N_7554,N_5547,N_5260);
nand U7555 (N_7555,N_4185,N_4696);
nand U7556 (N_7556,N_4723,N_5971);
nand U7557 (N_7557,N_1237,N_2349);
xor U7558 (N_7558,N_3199,N_5726);
or U7559 (N_7559,N_3410,N_4542);
nand U7560 (N_7560,N_3836,N_4800);
or U7561 (N_7561,N_936,N_1917);
or U7562 (N_7562,N_4664,N_4686);
nand U7563 (N_7563,N_3845,N_3527);
xor U7564 (N_7564,N_5810,N_2648);
and U7565 (N_7565,N_171,N_528);
nand U7566 (N_7566,N_1019,N_4853);
nand U7567 (N_7567,N_5255,N_2854);
or U7568 (N_7568,N_3325,N_1561);
nor U7569 (N_7569,N_2377,N_3689);
nor U7570 (N_7570,N_458,N_2039);
or U7571 (N_7571,N_3519,N_3381);
xor U7572 (N_7572,N_116,N_2502);
and U7573 (N_7573,N_4958,N_1398);
xnor U7574 (N_7574,N_985,N_2838);
or U7575 (N_7575,N_5449,N_3888);
nand U7576 (N_7576,N_5256,N_3612);
nand U7577 (N_7577,N_4594,N_3887);
or U7578 (N_7578,N_5253,N_1743);
nand U7579 (N_7579,N_4565,N_3100);
or U7580 (N_7580,N_2749,N_2640);
nor U7581 (N_7581,N_4634,N_4883);
nand U7582 (N_7582,N_5747,N_3217);
or U7583 (N_7583,N_1005,N_1657);
xor U7584 (N_7584,N_4465,N_945);
and U7585 (N_7585,N_1040,N_3304);
nor U7586 (N_7586,N_5501,N_5571);
nor U7587 (N_7587,N_172,N_1848);
xor U7588 (N_7588,N_2041,N_2975);
nand U7589 (N_7589,N_15,N_1483);
and U7590 (N_7590,N_3718,N_4629);
or U7591 (N_7591,N_2580,N_4263);
or U7592 (N_7592,N_3753,N_2692);
nand U7593 (N_7593,N_4808,N_3257);
nand U7594 (N_7594,N_2909,N_1903);
or U7595 (N_7595,N_3532,N_2674);
or U7596 (N_7596,N_1874,N_5491);
nand U7597 (N_7597,N_91,N_5504);
and U7598 (N_7598,N_5834,N_3047);
or U7599 (N_7599,N_5564,N_3727);
nand U7600 (N_7600,N_1203,N_5317);
nand U7601 (N_7601,N_4064,N_1606);
nor U7602 (N_7602,N_2672,N_4184);
nor U7603 (N_7603,N_3202,N_5294);
or U7604 (N_7604,N_4538,N_2055);
xnor U7605 (N_7605,N_4901,N_3794);
xnor U7606 (N_7606,N_5440,N_3889);
nor U7607 (N_7607,N_294,N_929);
xor U7608 (N_7608,N_2767,N_2600);
xor U7609 (N_7609,N_565,N_4803);
nand U7610 (N_7610,N_3685,N_4255);
or U7611 (N_7611,N_1855,N_1985);
nand U7612 (N_7612,N_4874,N_2970);
nor U7613 (N_7613,N_3059,N_1631);
nand U7614 (N_7614,N_3395,N_4776);
nor U7615 (N_7615,N_4371,N_4663);
nand U7616 (N_7616,N_3446,N_2276);
or U7617 (N_7617,N_3021,N_550);
nand U7618 (N_7618,N_5351,N_4070);
nand U7619 (N_7619,N_888,N_3815);
and U7620 (N_7620,N_5520,N_980);
nor U7621 (N_7621,N_4304,N_2427);
and U7622 (N_7622,N_2335,N_5894);
xor U7623 (N_7623,N_3577,N_239);
xnor U7624 (N_7624,N_163,N_1264);
nor U7625 (N_7625,N_3943,N_3843);
and U7626 (N_7626,N_2514,N_5037);
or U7627 (N_7627,N_1419,N_522);
or U7628 (N_7628,N_5899,N_5603);
xnor U7629 (N_7629,N_1119,N_483);
xnor U7630 (N_7630,N_3458,N_2476);
xor U7631 (N_7631,N_3525,N_207);
or U7632 (N_7632,N_1459,N_2296);
nor U7633 (N_7633,N_2910,N_792);
or U7634 (N_7634,N_1022,N_3415);
or U7635 (N_7635,N_2818,N_2011);
nor U7636 (N_7636,N_3254,N_749);
and U7637 (N_7637,N_3998,N_5228);
and U7638 (N_7638,N_2460,N_1571);
xor U7639 (N_7639,N_4470,N_5090);
xnor U7640 (N_7640,N_1895,N_1036);
or U7641 (N_7641,N_4689,N_553);
or U7642 (N_7642,N_1030,N_631);
and U7643 (N_7643,N_2752,N_4615);
xor U7644 (N_7644,N_5987,N_312);
or U7645 (N_7645,N_51,N_2478);
nand U7646 (N_7646,N_2317,N_1996);
and U7647 (N_7647,N_5554,N_1444);
nor U7648 (N_7648,N_3211,N_4755);
or U7649 (N_7649,N_2870,N_5192);
nand U7650 (N_7650,N_3142,N_5092);
or U7651 (N_7651,N_1682,N_1231);
and U7652 (N_7652,N_946,N_5026);
nand U7653 (N_7653,N_5109,N_1167);
xor U7654 (N_7654,N_5259,N_4927);
nand U7655 (N_7655,N_714,N_806);
nor U7656 (N_7656,N_588,N_3824);
or U7657 (N_7657,N_2830,N_3488);
xor U7658 (N_7658,N_3258,N_4558);
and U7659 (N_7659,N_871,N_836);
nand U7660 (N_7660,N_1310,N_90);
xor U7661 (N_7661,N_4730,N_5177);
or U7662 (N_7662,N_581,N_2174);
or U7663 (N_7663,N_4672,N_4300);
or U7664 (N_7664,N_5,N_1565);
nand U7665 (N_7665,N_4520,N_564);
nand U7666 (N_7666,N_4308,N_5937);
xnor U7667 (N_7667,N_4071,N_81);
and U7668 (N_7668,N_3099,N_5022);
xor U7669 (N_7669,N_3345,N_5650);
nand U7670 (N_7670,N_3409,N_5613);
and U7671 (N_7671,N_5201,N_1195);
or U7672 (N_7672,N_3800,N_2980);
nor U7673 (N_7673,N_1716,N_4877);
nor U7674 (N_7674,N_3071,N_4543);
nor U7675 (N_7675,N_560,N_125);
or U7676 (N_7676,N_347,N_795);
and U7677 (N_7677,N_2537,N_5276);
nand U7678 (N_7678,N_310,N_1511);
and U7679 (N_7679,N_2253,N_3620);
and U7680 (N_7680,N_5868,N_5388);
or U7681 (N_7681,N_990,N_2182);
nor U7682 (N_7682,N_849,N_1598);
and U7683 (N_7683,N_1788,N_5438);
nand U7684 (N_7684,N_2680,N_1353);
and U7685 (N_7685,N_839,N_4550);
xnor U7686 (N_7686,N_3082,N_797);
and U7687 (N_7687,N_19,N_3074);
and U7688 (N_7688,N_2313,N_574);
nand U7689 (N_7689,N_3322,N_3762);
nand U7690 (N_7690,N_1857,N_3580);
and U7691 (N_7691,N_175,N_2249);
or U7692 (N_7692,N_3538,N_1556);
or U7693 (N_7693,N_3312,N_1000);
and U7694 (N_7694,N_5755,N_4421);
and U7695 (N_7695,N_85,N_5897);
or U7696 (N_7696,N_1367,N_1932);
nor U7697 (N_7697,N_3244,N_2952);
nor U7698 (N_7698,N_2545,N_538);
and U7699 (N_7699,N_5015,N_5817);
nor U7700 (N_7700,N_4333,N_1508);
nor U7701 (N_7701,N_1488,N_4514);
nor U7702 (N_7702,N_3787,N_1819);
nor U7703 (N_7703,N_3109,N_5347);
and U7704 (N_7704,N_5699,N_2924);
or U7705 (N_7705,N_1327,N_4855);
nand U7706 (N_7706,N_3790,N_523);
xor U7707 (N_7707,N_4601,N_2560);
nand U7708 (N_7708,N_114,N_2020);
nand U7709 (N_7709,N_2363,N_4527);
nor U7710 (N_7710,N_2135,N_3969);
nor U7711 (N_7711,N_4473,N_351);
nor U7712 (N_7712,N_1493,N_3635);
and U7713 (N_7713,N_3424,N_4435);
nand U7714 (N_7714,N_2799,N_3628);
and U7715 (N_7715,N_3354,N_5423);
nand U7716 (N_7716,N_2390,N_5497);
nand U7717 (N_7717,N_655,N_962);
or U7718 (N_7718,N_1369,N_5221);
nor U7719 (N_7719,N_790,N_1377);
nand U7720 (N_7720,N_1254,N_2213);
and U7721 (N_7721,N_4237,N_2605);
or U7722 (N_7722,N_3863,N_3422);
nor U7723 (N_7723,N_4815,N_5281);
or U7724 (N_7724,N_1648,N_1863);
nor U7725 (N_7725,N_369,N_1979);
nor U7726 (N_7726,N_1033,N_5176);
or U7727 (N_7727,N_4501,N_689);
or U7728 (N_7728,N_661,N_4983);
nor U7729 (N_7729,N_3903,N_4141);
or U7730 (N_7730,N_4670,N_5461);
nand U7731 (N_7731,N_1889,N_11);
and U7732 (N_7732,N_2438,N_3721);
or U7733 (N_7733,N_2224,N_1929);
nor U7734 (N_7734,N_2606,N_4138);
or U7735 (N_7735,N_332,N_5965);
xnor U7736 (N_7736,N_2652,N_4393);
or U7737 (N_7737,N_5850,N_3765);
nand U7738 (N_7738,N_1970,N_5932);
or U7739 (N_7739,N_5127,N_796);
nor U7740 (N_7740,N_1355,N_1407);
and U7741 (N_7741,N_349,N_287);
nor U7742 (N_7742,N_4143,N_4144);
xnor U7743 (N_7743,N_2500,N_3641);
or U7744 (N_7744,N_1304,N_3766);
and U7745 (N_7745,N_1410,N_1259);
and U7746 (N_7746,N_4367,N_4424);
or U7747 (N_7747,N_5331,N_1931);
xor U7748 (N_7748,N_5689,N_3213);
and U7749 (N_7749,N_695,N_2578);
and U7750 (N_7750,N_1935,N_338);
and U7751 (N_7751,N_5947,N_950);
xor U7752 (N_7752,N_641,N_913);
nor U7753 (N_7753,N_1809,N_1115);
xnor U7754 (N_7754,N_1861,N_4174);
or U7755 (N_7755,N_5239,N_872);
and U7756 (N_7756,N_3012,N_2833);
or U7757 (N_7757,N_2876,N_3874);
and U7758 (N_7758,N_1302,N_3014);
nor U7759 (N_7759,N_2403,N_2632);
nand U7760 (N_7760,N_1256,N_26);
and U7761 (N_7761,N_5032,N_2136);
nand U7762 (N_7762,N_254,N_1779);
xor U7763 (N_7763,N_5558,N_5823);
nand U7764 (N_7764,N_488,N_2800);
nor U7765 (N_7765,N_1188,N_4325);
xor U7766 (N_7766,N_2898,N_2682);
nand U7767 (N_7767,N_1680,N_4496);
and U7768 (N_7768,N_3129,N_3551);
nand U7769 (N_7769,N_3104,N_2333);
xor U7770 (N_7770,N_4737,N_2089);
nor U7771 (N_7771,N_5345,N_5815);
nand U7772 (N_7772,N_1569,N_4024);
nor U7773 (N_7773,N_3544,N_1888);
nand U7774 (N_7774,N_4752,N_5240);
or U7775 (N_7775,N_3170,N_4564);
and U7776 (N_7776,N_478,N_2425);
nor U7777 (N_7777,N_1316,N_2092);
xor U7778 (N_7778,N_5350,N_2358);
xnor U7779 (N_7779,N_4787,N_5335);
or U7780 (N_7780,N_3920,N_1230);
or U7781 (N_7781,N_378,N_2613);
or U7782 (N_7782,N_1263,N_4440);
xor U7783 (N_7783,N_3743,N_5385);
nand U7784 (N_7784,N_4823,N_536);
or U7785 (N_7785,N_687,N_4860);
and U7786 (N_7786,N_3497,N_4301);
and U7787 (N_7787,N_1559,N_596);
and U7788 (N_7788,N_2396,N_3939);
or U7789 (N_7789,N_5193,N_5573);
nand U7790 (N_7790,N_2100,N_5114);
nand U7791 (N_7791,N_4417,N_4045);
and U7792 (N_7792,N_5467,N_665);
nor U7793 (N_7793,N_5746,N_484);
and U7794 (N_7794,N_4362,N_1382);
nor U7795 (N_7795,N_3076,N_4047);
xor U7796 (N_7796,N_586,N_4881);
xor U7797 (N_7797,N_2456,N_4280);
nand U7798 (N_7798,N_898,N_971);
nor U7799 (N_7799,N_2320,N_924);
and U7800 (N_7800,N_3088,N_3913);
and U7801 (N_7801,N_2151,N_5306);
or U7802 (N_7802,N_4210,N_3204);
and U7803 (N_7803,N_4453,N_4534);
nor U7804 (N_7804,N_3754,N_2731);
or U7805 (N_7805,N_842,N_3932);
or U7806 (N_7806,N_3549,N_4929);
xor U7807 (N_7807,N_4175,N_382);
xor U7808 (N_7808,N_556,N_1502);
and U7809 (N_7809,N_5367,N_3865);
xnor U7810 (N_7810,N_2101,N_3355);
nand U7811 (N_7811,N_3884,N_1145);
and U7812 (N_7812,N_2598,N_2494);
or U7813 (N_7813,N_1342,N_5100);
or U7814 (N_7814,N_1134,N_2795);
xor U7815 (N_7815,N_47,N_1580);
or U7816 (N_7816,N_2936,N_4196);
and U7817 (N_7817,N_912,N_1035);
nor U7818 (N_7818,N_1478,N_2932);
xor U7819 (N_7819,N_1395,N_4042);
and U7820 (N_7820,N_546,N_1112);
nand U7821 (N_7821,N_3587,N_4873);
nand U7822 (N_7822,N_4626,N_4161);
nand U7823 (N_7823,N_3449,N_3849);
or U7824 (N_7824,N_3228,N_2307);
xnor U7825 (N_7825,N_204,N_756);
and U7826 (N_7826,N_4797,N_3594);
nor U7827 (N_7827,N_1266,N_646);
or U7828 (N_7828,N_50,N_4921);
or U7829 (N_7829,N_960,N_5707);
nand U7830 (N_7830,N_213,N_5500);
and U7831 (N_7831,N_2023,N_4997);
xor U7832 (N_7832,N_3688,N_3023);
xor U7833 (N_7833,N_1308,N_381);
nand U7834 (N_7834,N_1892,N_2300);
and U7835 (N_7835,N_989,N_927);
nand U7836 (N_7836,N_3502,N_5827);
or U7837 (N_7837,N_1171,N_2571);
nor U7838 (N_7838,N_1973,N_623);
or U7839 (N_7839,N_27,N_3130);
nand U7840 (N_7840,N_1835,N_5737);
xnor U7841 (N_7841,N_1660,N_1751);
nor U7842 (N_7842,N_1806,N_3060);
or U7843 (N_7843,N_658,N_486);
nor U7844 (N_7844,N_2272,N_5172);
nand U7845 (N_7845,N_273,N_1607);
xor U7846 (N_7846,N_5072,N_1351);
nand U7847 (N_7847,N_4063,N_4344);
xnor U7848 (N_7848,N_5463,N_4223);
nand U7849 (N_7849,N_3123,N_2102);
nand U7850 (N_7850,N_5008,N_2589);
xnor U7851 (N_7851,N_2114,N_5180);
or U7852 (N_7852,N_1184,N_1771);
xnor U7853 (N_7853,N_92,N_5280);
xnor U7854 (N_7854,N_4600,N_537);
nor U7855 (N_7855,N_4945,N_4915);
and U7856 (N_7856,N_79,N_3691);
nor U7857 (N_7857,N_2630,N_1620);
nor U7858 (N_7858,N_5327,N_4260);
or U7859 (N_7859,N_1789,N_525);
and U7860 (N_7860,N_5246,N_2785);
nor U7861 (N_7861,N_930,N_465);
nand U7862 (N_7862,N_5410,N_1428);
or U7863 (N_7863,N_4882,N_3342);
or U7864 (N_7864,N_4838,N_2633);
xnor U7865 (N_7865,N_5018,N_1409);
nand U7866 (N_7866,N_3361,N_1226);
nand U7867 (N_7867,N_2166,N_672);
nand U7868 (N_7868,N_3102,N_2557);
or U7869 (N_7869,N_2226,N_1825);
or U7870 (N_7870,N_2565,N_4146);
xor U7871 (N_7871,N_3828,N_3500);
xnor U7872 (N_7872,N_1106,N_4781);
and U7873 (N_7873,N_4700,N_3306);
nor U7874 (N_7874,N_5460,N_882);
and U7875 (N_7875,N_5487,N_2809);
and U7876 (N_7876,N_809,N_4839);
or U7877 (N_7877,N_5879,N_225);
nor U7878 (N_7878,N_5895,N_5911);
nor U7879 (N_7879,N_2435,N_2625);
or U7880 (N_7880,N_3911,N_894);
xnor U7881 (N_7881,N_4092,N_1756);
or U7882 (N_7882,N_1322,N_5855);
and U7883 (N_7883,N_2155,N_5599);
and U7884 (N_7884,N_5365,N_3936);
nand U7885 (N_7885,N_5333,N_3218);
nor U7886 (N_7886,N_5214,N_5555);
nand U7887 (N_7887,N_174,N_1423);
nor U7888 (N_7888,N_2905,N_2676);
and U7889 (N_7889,N_1085,N_1324);
xor U7890 (N_7890,N_4864,N_3515);
nor U7891 (N_7891,N_4660,N_2334);
xor U7892 (N_7892,N_1346,N_3892);
xnor U7893 (N_7893,N_4037,N_111);
nor U7894 (N_7894,N_3002,N_5667);
or U7895 (N_7895,N_288,N_856);
nand U7896 (N_7896,N_4131,N_3010);
or U7897 (N_7897,N_3495,N_3506);
and U7898 (N_7898,N_3829,N_1831);
nor U7899 (N_7899,N_4359,N_2219);
nand U7900 (N_7900,N_167,N_1354);
nand U7901 (N_7901,N_4828,N_3317);
nand U7902 (N_7902,N_3387,N_3615);
or U7903 (N_7903,N_5166,N_3015);
or U7904 (N_7904,N_4870,N_884);
or U7905 (N_7905,N_2365,N_3684);
nor U7906 (N_7906,N_5415,N_276);
or U7907 (N_7907,N_617,N_2902);
nor U7908 (N_7908,N_394,N_4098);
or U7909 (N_7909,N_3503,N_3190);
and U7910 (N_7910,N_3905,N_3219);
or U7911 (N_7911,N_376,N_2769);
xnor U7912 (N_7912,N_1340,N_5225);
nor U7913 (N_7913,N_5598,N_5178);
xor U7914 (N_7914,N_4090,N_1038);
nand U7915 (N_7915,N_1507,N_450);
nor U7916 (N_7916,N_965,N_4302);
nor U7917 (N_7917,N_229,N_2871);
and U7918 (N_7918,N_4653,N_3859);
nand U7919 (N_7919,N_3970,N_5021);
xnor U7920 (N_7920,N_1336,N_2999);
xnor U7921 (N_7921,N_3596,N_5107);
xor U7922 (N_7922,N_3675,N_841);
and U7923 (N_7923,N_4313,N_5567);
or U7924 (N_7924,N_1175,N_3690);
and U7925 (N_7925,N_462,N_2036);
xnor U7926 (N_7926,N_2042,N_3651);
and U7927 (N_7927,N_3879,N_5793);
nand U7928 (N_7928,N_4342,N_2156);
xor U7929 (N_7929,N_3929,N_4850);
or U7930 (N_7930,N_5029,N_2108);
and U7931 (N_7931,N_3820,N_2158);
or U7932 (N_7932,N_3319,N_4107);
xnor U7933 (N_7933,N_5941,N_188);
nand U7934 (N_7934,N_4297,N_4249);
xor U7935 (N_7935,N_4847,N_592);
and U7936 (N_7936,N_4733,N_1285);
and U7937 (N_7937,N_2593,N_1702);
nor U7938 (N_7938,N_2096,N_3331);
nor U7939 (N_7939,N_5421,N_5395);
nand U7940 (N_7940,N_1515,N_698);
nor U7941 (N_7941,N_4825,N_5551);
nand U7942 (N_7942,N_2706,N_2755);
or U7943 (N_7943,N_4029,N_5740);
nand U7944 (N_7944,N_2860,N_2584);
nand U7945 (N_7945,N_2660,N_3118);
and U7946 (N_7946,N_2903,N_1726);
and U7947 (N_7947,N_1422,N_4944);
nand U7948 (N_7948,N_3406,N_4544);
nor U7949 (N_7949,N_1199,N_1153);
xnor U7950 (N_7950,N_2140,N_4152);
nor U7951 (N_7951,N_3191,N_2926);
nand U7952 (N_7952,N_5711,N_4896);
and U7953 (N_7953,N_4101,N_554);
xnor U7954 (N_7954,N_1463,N_2547);
xnor U7955 (N_7955,N_5341,N_5477);
nand U7956 (N_7956,N_3172,N_5703);
xor U7957 (N_7957,N_5293,N_3793);
xnor U7958 (N_7958,N_1442,N_5902);
xor U7959 (N_7959,N_1658,N_630);
nor U7960 (N_7960,N_4972,N_1506);
nand U7961 (N_7961,N_1770,N_2783);
xor U7962 (N_7962,N_2125,N_2187);
xnor U7963 (N_7963,N_3818,N_1585);
xnor U7964 (N_7964,N_1663,N_3473);
or U7965 (N_7965,N_2046,N_2711);
xor U7966 (N_7966,N_5019,N_4952);
or U7967 (N_7967,N_3193,N_3461);
and U7968 (N_7968,N_761,N_5378);
and U7969 (N_7969,N_5597,N_5238);
and U7970 (N_7970,N_3700,N_569);
nand U7971 (N_7971,N_1783,N_1516);
nor U7972 (N_7972,N_3210,N_4340);
nor U7973 (N_7973,N_5841,N_5158);
nor U7974 (N_7974,N_2322,N_5883);
nor U7975 (N_7975,N_5727,N_264);
nor U7976 (N_7976,N_3072,N_4792);
or U7977 (N_7977,N_1374,N_1564);
nor U7978 (N_7978,N_5184,N_4597);
or U7979 (N_7979,N_4574,N_5760);
and U7980 (N_7980,N_389,N_4722);
or U7981 (N_7981,N_5957,N_3298);
nor U7982 (N_7982,N_3297,N_5020);
or U7983 (N_7983,N_4777,N_3864);
nand U7984 (N_7984,N_159,N_4957);
or U7985 (N_7985,N_1015,N_4247);
nand U7986 (N_7986,N_5998,N_5040);
or U7987 (N_7987,N_2251,N_2201);
nand U7988 (N_7988,N_5682,N_1465);
xnor U7989 (N_7989,N_3872,N_1265);
and U7990 (N_7990,N_4756,N_5496);
xnor U7991 (N_7991,N_4936,N_2786);
nand U7992 (N_7992,N_2461,N_5413);
nand U7993 (N_7993,N_4869,N_4774);
or U7994 (N_7994,N_2586,N_2572);
or U7995 (N_7995,N_1908,N_1710);
and U7996 (N_7996,N_1111,N_5507);
or U7997 (N_7997,N_2185,N_5334);
nor U7998 (N_7998,N_2742,N_2260);
nor U7999 (N_7999,N_5086,N_3921);
xnor U8000 (N_8000,N_4148,N_2576);
nor U8001 (N_8001,N_5517,N_4969);
and U8002 (N_8002,N_5923,N_5776);
and U8003 (N_8003,N_1060,N_566);
or U8004 (N_8004,N_1933,N_4341);
nor U8005 (N_8005,N_3078,N_1823);
nor U8006 (N_8006,N_3276,N_2912);
xnor U8007 (N_8007,N_3826,N_2907);
xnor U8008 (N_8008,N_2168,N_3299);
nor U8009 (N_8009,N_5330,N_87);
or U8010 (N_8010,N_4118,N_5373);
or U8011 (N_8011,N_5681,N_4053);
xnor U8012 (N_8012,N_2577,N_4633);
nor U8013 (N_8013,N_2152,N_5113);
nor U8014 (N_8014,N_4782,N_850);
or U8015 (N_8015,N_2144,N_4791);
or U8016 (N_8016,N_878,N_5053);
and U8017 (N_8017,N_2087,N_4576);
or U8018 (N_8018,N_2161,N_4971);
or U8019 (N_8019,N_4849,N_931);
nand U8020 (N_8020,N_3280,N_2725);
xor U8021 (N_8021,N_573,N_1017);
or U8022 (N_8022,N_3185,N_1414);
and U8023 (N_8023,N_5553,N_1390);
and U8024 (N_8024,N_3934,N_4605);
xor U8025 (N_8025,N_439,N_2063);
nor U8026 (N_8026,N_1539,N_5624);
nor U8027 (N_8027,N_5416,N_1403);
or U8028 (N_8028,N_745,N_3901);
or U8029 (N_8029,N_675,N_1386);
xor U8030 (N_8030,N_5150,N_5363);
xnor U8031 (N_8031,N_1642,N_5677);
nor U8032 (N_8032,N_1154,N_4892);
xor U8033 (N_8033,N_4977,N_3188);
nand U8034 (N_8034,N_3052,N_4926);
nand U8035 (N_8035,N_921,N_735);
nor U8036 (N_8036,N_3020,N_4897);
or U8037 (N_8037,N_977,N_3648);
nor U8038 (N_8038,N_4254,N_2248);
nand U8039 (N_8039,N_2562,N_2405);
nand U8040 (N_8040,N_4272,N_5007);
nand U8041 (N_8041,N_935,N_2990);
and U8042 (N_8042,N_2880,N_561);
nand U8043 (N_8043,N_1916,N_1622);
or U8044 (N_8044,N_4377,N_5666);
and U8045 (N_8045,N_201,N_3011);
nor U8046 (N_8046,N_4099,N_2866);
nor U8047 (N_8047,N_4827,N_2271);
xnor U8048 (N_8048,N_4374,N_137);
nor U8049 (N_8049,N_2275,N_4895);
xor U8050 (N_8050,N_5757,N_1222);
xor U8051 (N_8051,N_2773,N_5446);
or U8052 (N_8052,N_1646,N_1724);
and U8053 (N_8053,N_1383,N_5762);
nor U8054 (N_8054,N_4599,N_2678);
and U8055 (N_8055,N_1818,N_4691);
xor U8056 (N_8056,N_1653,N_3637);
and U8057 (N_8057,N_401,N_5742);
xnor U8058 (N_8058,N_3880,N_812);
xor U8059 (N_8059,N_440,N_2103);
or U8060 (N_8060,N_2543,N_2524);
xor U8061 (N_8061,N_4652,N_2165);
or U8062 (N_8062,N_3318,N_1597);
nor U8063 (N_8063,N_4647,N_2851);
or U8064 (N_8064,N_3741,N_150);
xor U8065 (N_8065,N_3882,N_1750);
nand U8066 (N_8066,N_4753,N_3373);
and U8067 (N_8067,N_5831,N_3761);
nand U8068 (N_8068,N_2523,N_1126);
or U8069 (N_8069,N_253,N_5278);
xor U8070 (N_8070,N_1904,N_277);
and U8071 (N_8071,N_4530,N_3950);
xnor U8072 (N_8072,N_1261,N_2507);
nor U8073 (N_8073,N_1080,N_2559);
xor U8074 (N_8074,N_4123,N_3398);
nor U8075 (N_8075,N_803,N_1107);
nand U8076 (N_8076,N_4081,N_1384);
or U8077 (N_8077,N_5773,N_3709);
nand U8078 (N_8078,N_5412,N_2634);
nor U8079 (N_8079,N_4001,N_3586);
nand U8080 (N_8080,N_3201,N_5684);
nor U8081 (N_8081,N_3154,N_4195);
or U8082 (N_8082,N_5277,N_3249);
nand U8083 (N_8083,N_4816,N_1937);
nand U8084 (N_8084,N_4162,N_3774);
xor U8085 (N_8085,N_4439,N_5471);
or U8086 (N_8086,N_3137,N_4793);
xnor U8087 (N_8087,N_5126,N_826);
nor U8088 (N_8088,N_255,N_1830);
nand U8089 (N_8089,N_2418,N_5974);
and U8090 (N_8090,N_1840,N_3616);
nor U8091 (N_8091,N_5589,N_3303);
nand U8092 (N_8092,N_3823,N_453);
nand U8093 (N_8093,N_5914,N_3291);
and U8094 (N_8094,N_4690,N_1349);
and U8095 (N_8095,N_156,N_5482);
nor U8096 (N_8096,N_5493,N_5337);
and U8097 (N_8097,N_5559,N_2374);
nor U8098 (N_8098,N_5196,N_1675);
nand U8099 (N_8099,N_5409,N_5128);
or U8100 (N_8100,N_3397,N_1766);
and U8101 (N_8101,N_2933,N_2793);
nand U8102 (N_8102,N_2715,N_4158);
and U8103 (N_8103,N_4810,N_4337);
nand U8104 (N_8104,N_5875,N_1337);
and U8105 (N_8105,N_4452,N_4431);
or U8106 (N_8106,N_1191,N_5903);
nand U8107 (N_8107,N_531,N_4728);
or U8108 (N_8108,N_345,N_4727);
xnor U8109 (N_8109,N_3269,N_5233);
and U8110 (N_8110,N_1193,N_3245);
and U8111 (N_8111,N_2665,N_923);
nor U8112 (N_8112,N_2439,N_2356);
nand U8113 (N_8113,N_5803,N_1781);
or U8114 (N_8114,N_1048,N_1669);
and U8115 (N_8115,N_1661,N_89);
and U8116 (N_8116,N_4281,N_4294);
or U8117 (N_8117,N_5907,N_2671);
xor U8118 (N_8118,N_1034,N_906);
or U8119 (N_8119,N_2834,N_2802);
or U8120 (N_8120,N_1087,N_1144);
nand U8121 (N_8121,N_3466,N_359);
nor U8122 (N_8122,N_1312,N_1391);
and U8123 (N_8123,N_3671,N_1358);
nand U8124 (N_8124,N_5147,N_1121);
nor U8125 (N_8125,N_2825,N_5736);
and U8126 (N_8126,N_2712,N_3063);
or U8127 (N_8127,N_5508,N_5716);
and U8128 (N_8128,N_1532,N_5251);
or U8129 (N_8129,N_3320,N_1608);
and U8130 (N_8130,N_3713,N_243);
or U8131 (N_8131,N_2203,N_3692);
nand U8132 (N_8132,N_5134,N_5978);
and U8133 (N_8133,N_755,N_2145);
or U8134 (N_8134,N_3860,N_218);
and U8135 (N_8135,N_3965,N_5739);
or U8136 (N_8136,N_3611,N_1429);
or U8137 (N_8137,N_3032,N_2976);
or U8138 (N_8138,N_3364,N_1252);
xor U8139 (N_8139,N_2259,N_5920);
nor U8140 (N_8140,N_647,N_4998);
or U8141 (N_8141,N_2214,N_2234);
xnor U8142 (N_8142,N_3157,N_1297);
nand U8143 (N_8143,N_2972,N_5189);
nor U8144 (N_8144,N_2759,N_5878);
and U8145 (N_8145,N_123,N_2429);
nor U8146 (N_8146,N_4949,N_4718);
or U8147 (N_8147,N_659,N_3705);
and U8148 (N_8148,N_3789,N_250);
nand U8149 (N_8149,N_4125,N_1041);
or U8150 (N_8150,N_1446,N_5194);
or U8151 (N_8151,N_2698,N_4930);
nand U8152 (N_8152,N_4772,N_1997);
nand U8153 (N_8153,N_2131,N_4387);
and U8154 (N_8154,N_3898,N_65);
xnor U8155 (N_8155,N_75,N_223);
nor U8156 (N_8156,N_3979,N_1595);
xnor U8157 (N_8157,N_5332,N_5611);
and U8158 (N_8158,N_4833,N_4039);
nor U8159 (N_8159,N_4822,N_5084);
nand U8160 (N_8160,N_3375,N_5159);
or U8161 (N_8161,N_5065,N_2693);
nand U8162 (N_8162,N_5901,N_5616);
and U8163 (N_8163,N_5070,N_4813);
nor U8164 (N_8164,N_4764,N_595);
and U8165 (N_8165,N_1186,N_3323);
nand U8166 (N_8166,N_2527,N_3400);
or U8167 (N_8167,N_1549,N_1794);
nand U8168 (N_8168,N_3540,N_2304);
or U8169 (N_8169,N_4463,N_3212);
xnor U8170 (N_8170,N_5908,N_3697);
nand U8171 (N_8171,N_410,N_3226);
and U8172 (N_8172,N_2544,N_1241);
nand U8173 (N_8173,N_5064,N_4318);
nand U8174 (N_8174,N_5252,N_1245);
nor U8175 (N_8175,N_1470,N_785);
nand U8176 (N_8176,N_1815,N_1555);
xor U8177 (N_8177,N_3734,N_2873);
nand U8178 (N_8178,N_1560,N_1639);
and U8179 (N_8179,N_2215,N_4989);
or U8180 (N_8180,N_2279,N_996);
and U8181 (N_8181,N_1677,N_829);
or U8182 (N_8182,N_1456,N_1025);
nand U8183 (N_8183,N_4830,N_2803);
and U8184 (N_8184,N_5887,N_4980);
or U8185 (N_8185,N_1094,N_4235);
xnor U8186 (N_8186,N_3983,N_5545);
and U8187 (N_8187,N_1787,N_5602);
or U8188 (N_8188,N_1665,N_4228);
nor U8189 (N_8189,N_5537,N_2402);
nand U8190 (N_8190,N_1317,N_94);
xor U8191 (N_8191,N_3440,N_3041);
xor U8192 (N_8192,N_2223,N_4695);
and U8193 (N_8193,N_5820,N_220);
xor U8194 (N_8194,N_1330,N_5316);
xnor U8195 (N_8195,N_3537,N_5983);
and U8196 (N_8196,N_5732,N_4226);
nand U8197 (N_8197,N_3926,N_3777);
and U8198 (N_8198,N_1181,N_3595);
or U8199 (N_8199,N_3207,N_2482);
and U8200 (N_8200,N_3954,N_4589);
nor U8201 (N_8201,N_2117,N_4080);
xnor U8202 (N_8202,N_4504,N_492);
nor U8203 (N_8203,N_559,N_5300);
xor U8204 (N_8204,N_2391,N_2709);
or U8205 (N_8205,N_259,N_2183);
nand U8206 (N_8206,N_4062,N_1207);
or U8207 (N_8207,N_5362,N_4563);
or U8208 (N_8208,N_680,N_939);
xnor U8209 (N_8209,N_104,N_615);
and U8210 (N_8210,N_640,N_1436);
nand U8211 (N_8211,N_547,N_1759);
nor U8212 (N_8212,N_4353,N_3509);
and U8213 (N_8213,N_2675,N_141);
nor U8214 (N_8214,N_2651,N_5991);
xor U8215 (N_8215,N_1603,N_2289);
xnor U8216 (N_8216,N_3985,N_222);
nand U8217 (N_8217,N_1260,N_3585);
nor U8218 (N_8218,N_905,N_1596);
and U8219 (N_8219,N_246,N_4225);
or U8220 (N_8220,N_373,N_1246);
or U8221 (N_8221,N_3696,N_5082);
or U8222 (N_8222,N_4261,N_4794);
or U8223 (N_8223,N_34,N_3900);
xnor U8224 (N_8224,N_3111,N_1990);
xnor U8225 (N_8225,N_4135,N_61);
nor U8226 (N_8226,N_2483,N_5688);
and U8227 (N_8227,N_5455,N_39);
nor U8228 (N_8228,N_2352,N_5805);
xor U8229 (N_8229,N_3391,N_5672);
and U8230 (N_8230,N_2076,N_18);
xnor U8231 (N_8231,N_1430,N_5775);
or U8232 (N_8232,N_3891,N_4953);
xnor U8233 (N_8233,N_4119,N_4236);
or U8234 (N_8234,N_3737,N_5402);
xor U8235 (N_8235,N_1763,N_395);
and U8236 (N_8236,N_1402,N_4277);
and U8237 (N_8237,N_3416,N_2442);
nor U8238 (N_8238,N_1120,N_3662);
and U8239 (N_8239,N_3008,N_3095);
nand U8240 (N_8240,N_449,N_3636);
xor U8241 (N_8241,N_2050,N_5863);
nand U8242 (N_8242,N_2998,N_235);
nor U8243 (N_8243,N_3252,N_759);
and U8244 (N_8244,N_3742,N_4843);
or U8245 (N_8245,N_5970,N_4736);
or U8246 (N_8246,N_2216,N_2196);
or U8247 (N_8247,N_4163,N_5232);
nor U8248 (N_8248,N_2293,N_3350);
xor U8249 (N_8249,N_601,N_2760);
and U8250 (N_8250,N_1147,N_4268);
xor U8251 (N_8251,N_5593,N_4844);
and U8252 (N_8252,N_4785,N_503);
nor U8253 (N_8253,N_4935,N_4222);
nor U8254 (N_8254,N_1326,N_4698);
xor U8255 (N_8255,N_2094,N_3144);
or U8256 (N_8256,N_5287,N_5375);
xor U8257 (N_8257,N_139,N_798);
nand U8258 (N_8258,N_2243,N_4408);
nand U8259 (N_8259,N_4559,N_4754);
and U8260 (N_8260,N_3804,N_526);
or U8261 (N_8261,N_879,N_904);
or U8262 (N_8262,N_1073,N_2750);
and U8263 (N_8263,N_621,N_5465);
nor U8264 (N_8264,N_1614,N_3993);
and U8265 (N_8265,N_4714,N_3432);
nand U8266 (N_8266,N_578,N_1545);
xor U8267 (N_8267,N_425,N_3658);
nand U8268 (N_8268,N_4190,N_976);
nand U8269 (N_8269,N_2979,N_3418);
or U8270 (N_8270,N_2805,N_2075);
nor U8271 (N_8271,N_1255,N_4547);
xor U8272 (N_8272,N_4170,N_77);
nand U8273 (N_8273,N_848,N_138);
and U8274 (N_8274,N_4545,N_1320);
nor U8275 (N_8275,N_4303,N_2359);
xor U8276 (N_8276,N_4734,N_827);
nor U8277 (N_8277,N_2395,N_2581);
xnor U8278 (N_8278,N_2464,N_4258);
nand U8279 (N_8279,N_1676,N_2091);
or U8280 (N_8280,N_3292,N_3346);
nor U8281 (N_8281,N_3949,N_982);
or U8282 (N_8282,N_3174,N_656);
nor U8283 (N_8283,N_2417,N_2954);
nand U8284 (N_8284,N_5033,N_4579);
or U8285 (N_8285,N_3504,N_3574);
nor U8286 (N_8286,N_1691,N_3833);
xnor U8287 (N_8287,N_2768,N_1797);
nor U8288 (N_8288,N_4546,N_587);
nor U8289 (N_8289,N_1894,N_482);
or U8290 (N_8290,N_535,N_73);
and U8291 (N_8291,N_4584,N_4168);
xor U8292 (N_8292,N_2077,N_938);
xnor U8293 (N_8293,N_5574,N_339);
and U8294 (N_8294,N_1934,N_377);
nand U8295 (N_8295,N_2835,N_86);
nand U8296 (N_8296,N_1798,N_3731);
or U8297 (N_8297,N_3852,N_2601);
xor U8298 (N_8298,N_2113,N_3679);
and U8299 (N_8299,N_4192,N_5926);
nand U8300 (N_8300,N_5679,N_1768);
and U8301 (N_8301,N_5057,N_824);
and U8302 (N_8302,N_3621,N_5561);
xnor U8303 (N_8303,N_4940,N_4515);
or U8304 (N_8304,N_206,N_4407);
nor U8305 (N_8305,N_1158,N_3579);
xor U8306 (N_8306,N_1350,N_3362);
or U8307 (N_8307,N_5056,N_1629);
or U8308 (N_8308,N_4469,N_957);
xnor U8309 (N_8309,N_4482,N_4103);
xnor U8310 (N_8310,N_3571,N_1833);
nand U8311 (N_8311,N_2007,N_4132);
or U8312 (N_8312,N_1905,N_4738);
nor U8313 (N_8313,N_4835,N_4583);
nor U8314 (N_8314,N_3294,N_1533);
nand U8315 (N_8315,N_5655,N_820);
xor U8316 (N_8316,N_4401,N_4575);
nand U8317 (N_8317,N_5249,N_2567);
nand U8318 (N_8318,N_306,N_2362);
and U8319 (N_8319,N_3343,N_2257);
nand U8320 (N_8320,N_262,N_3867);
nand U8321 (N_8321,N_1550,N_390);
and U8322 (N_8322,N_2934,N_2244);
or U8323 (N_8323,N_3953,N_5596);
nand U8324 (N_8324,N_4562,N_765);
nand U8325 (N_8325,N_3396,N_1860);
nand U8326 (N_8326,N_4779,N_3978);
xnor U8327 (N_8327,N_146,N_4747);
and U8328 (N_8328,N_3886,N_4398);
or U8329 (N_8329,N_1325,N_1296);
or U8330 (N_8330,N_1063,N_4399);
xor U8331 (N_8331,N_5888,N_4410);
nor U8332 (N_8332,N_2323,N_4991);
nand U8333 (N_8333,N_2217,N_2496);
nand U8334 (N_8334,N_3419,N_793);
nand U8335 (N_8335,N_3287,N_548);
nand U8336 (N_8336,N_2717,N_3069);
nand U8337 (N_8337,N_1415,N_1404);
and U8338 (N_8338,N_2579,N_3904);
and U8339 (N_8339,N_4003,N_1221);
nand U8340 (N_8340,N_2991,N_1435);
nand U8341 (N_8341,N_2790,N_2045);
and U8342 (N_8342,N_2222,N_4751);
nor U8343 (N_8343,N_2184,N_1799);
nand U8344 (N_8344,N_1381,N_5139);
or U8345 (N_8345,N_5244,N_5268);
or U8346 (N_8346,N_2716,N_4517);
and U8347 (N_8347,N_2757,N_4919);
or U8348 (N_8348,N_1948,N_520);
or U8349 (N_8349,N_2570,N_810);
nor U8350 (N_8350,N_337,N_2398);
xor U8351 (N_8351,N_783,N_605);
xor U8352 (N_8352,N_5398,N_2687);
or U8353 (N_8353,N_2729,N_4438);
xor U8354 (N_8354,N_1477,N_355);
or U8355 (N_8355,N_409,N_3277);
nor U8356 (N_8356,N_3550,N_157);
xnor U8357 (N_8357,N_5913,N_2469);
or U8358 (N_8358,N_1024,N_3991);
nor U8359 (N_8359,N_2472,N_5060);
nand U8360 (N_8360,N_4773,N_4312);
nand U8361 (N_8361,N_2997,N_3521);
xor U8362 (N_8362,N_4164,N_4788);
and U8363 (N_8363,N_1177,N_2079);
xor U8364 (N_8364,N_5344,N_4999);
and U8365 (N_8365,N_3672,N_1583);
xor U8366 (N_8366,N_3089,N_5205);
and U8367 (N_8367,N_2556,N_843);
or U8368 (N_8368,N_4032,N_919);
nor U8369 (N_8369,N_4577,N_5215);
nor U8370 (N_8370,N_677,N_433);
and U8371 (N_8371,N_481,N_1400);
xor U8372 (N_8372,N_683,N_825);
and U8373 (N_8373,N_3313,N_4817);
and U8374 (N_8374,N_3927,N_5013);
nand U8375 (N_8375,N_1281,N_4934);
and U8376 (N_8376,N_3327,N_5148);
and U8377 (N_8377,N_3768,N_4617);
and U8378 (N_8378,N_2857,N_684);
nand U8379 (N_8379,N_5456,N_2510);
xor U8380 (N_8380,N_4040,N_2904);
nor U8381 (N_8381,N_987,N_5340);
xnor U8382 (N_8382,N_1021,N_3711);
and U8383 (N_8383,N_1529,N_3475);
or U8384 (N_8384,N_2826,N_5950);
xnor U8385 (N_8385,N_3752,N_3822);
nor U8386 (N_8386,N_162,N_5569);
xor U8387 (N_8387,N_3534,N_5156);
and U8388 (N_8388,N_240,N_3196);
and U8389 (N_8389,N_1443,N_1647);
and U8390 (N_8390,N_5772,N_2609);
xor U8391 (N_8391,N_1898,N_4242);
nand U8392 (N_8392,N_4188,N_5217);
xnor U8393 (N_8393,N_788,N_5836);
and U8394 (N_8394,N_5582,N_632);
or U8395 (N_8395,N_3084,N_3554);
nand U8396 (N_8396,N_4721,N_5121);
nor U8397 (N_8397,N_1345,N_66);
and U8398 (N_8398,N_2566,N_2048);
or U8399 (N_8399,N_4176,N_5698);
or U8400 (N_8400,N_517,N_2167);
or U8401 (N_8401,N_5374,N_5146);
xnor U8402 (N_8402,N_5085,N_5936);
nand U8403 (N_8403,N_231,N_4033);
nand U8404 (N_8404,N_1162,N_1530);
xor U8405 (N_8405,N_2919,N_1902);
xor U8406 (N_8406,N_1243,N_4622);
nor U8407 (N_8407,N_1913,N_1392);
and U8408 (N_8408,N_1943,N_3982);
and U8409 (N_8409,N_1673,N_3131);
or U8410 (N_8410,N_3661,N_2708);
nand U8411 (N_8411,N_5149,N_3296);
or U8412 (N_8412,N_558,N_2308);
and U8413 (N_8413,N_5687,N_245);
nor U8414 (N_8414,N_3728,N_4048);
or U8415 (N_8415,N_4885,N_350);
or U8416 (N_8416,N_1272,N_4293);
and U8417 (N_8417,N_4557,N_728);
xor U8418 (N_8418,N_4289,N_3316);
nand U8419 (N_8419,N_5543,N_4649);
or U8420 (N_8420,N_2986,N_666);
nand U8421 (N_8421,N_5017,N_1251);
nor U8422 (N_8422,N_5552,N_497);
or U8423 (N_8423,N_2806,N_2602);
nand U8424 (N_8424,N_645,N_437);
nand U8425 (N_8425,N_5368,N_5856);
nor U8426 (N_8426,N_1303,N_1689);
or U8427 (N_8427,N_1575,N_2451);
xnor U8428 (N_8428,N_326,N_5956);
nor U8429 (N_8429,N_743,N_5671);
xor U8430 (N_8430,N_1662,N_199);
or U8431 (N_8431,N_4609,N_1784);
xnor U8432 (N_8432,N_4150,N_1605);
nand U8433 (N_8433,N_5279,N_4178);
nand U8434 (N_8434,N_750,N_4968);
and U8435 (N_8435,N_72,N_5979);
xnor U8436 (N_8436,N_1378,N_5069);
and U8437 (N_8437,N_2034,N_916);
nand U8438 (N_8438,N_4505,N_534);
nand U8439 (N_8439,N_2604,N_5338);
xnor U8440 (N_8440,N_4886,N_5443);
xnor U8441 (N_8441,N_3513,N_4317);
and U8442 (N_8442,N_542,N_3909);
nor U8443 (N_8443,N_5704,N_3999);
xnor U8444 (N_8444,N_629,N_4512);
or U8445 (N_8445,N_4606,N_3899);
nor U8446 (N_8446,N_3942,N_417);
xor U8447 (N_8447,N_1651,N_1741);
nand U8448 (N_8448,N_1086,N_4783);
xor U8449 (N_8449,N_2180,N_1294);
or U8450 (N_8450,N_4798,N_317);
nor U8451 (N_8451,N_5396,N_4716);
xor U8452 (N_8452,N_3096,N_1236);
or U8453 (N_8453,N_2657,N_3197);
nand U8454 (N_8454,N_4611,N_861);
nand U8455 (N_8455,N_260,N_1841);
nand U8456 (N_8456,N_5652,N_4073);
nor U8457 (N_8457,N_1365,N_2499);
and U8458 (N_8458,N_179,N_5749);
xnor U8459 (N_8459,N_4155,N_1873);
or U8460 (N_8460,N_5648,N_5161);
nand U8461 (N_8461,N_5787,N_3181);
xor U8462 (N_8462,N_1348,N_2134);
and U8463 (N_8463,N_1890,N_283);
xnor U8464 (N_8464,N_1936,N_3668);
nand U8465 (N_8465,N_5600,N_2812);
nand U8466 (N_8466,N_5898,N_5519);
xnor U8467 (N_8467,N_5651,N_2631);
or U8468 (N_8468,N_4491,N_2561);
and U8469 (N_8469,N_498,N_5871);
and U8470 (N_8470,N_2242,N_3079);
or U8471 (N_8471,N_1051,N_5986);
xor U8472 (N_8472,N_5958,N_2701);
or U8473 (N_8473,N_1289,N_5048);
xor U8474 (N_8474,N_2819,N_3272);
nor U8475 (N_8475,N_3847,N_5795);
nor U8476 (N_8476,N_2319,N_774);
or U8477 (N_8477,N_3576,N_3526);
or U8478 (N_8478,N_4256,N_3057);
or U8479 (N_8479,N_3405,N_889);
xor U8480 (N_8480,N_5892,N_3112);
and U8481 (N_8481,N_1146,N_4427);
nand U8482 (N_8482,N_3674,N_3064);
nor U8483 (N_8483,N_1081,N_763);
and U8484 (N_8484,N_3659,N_2118);
xnor U8485 (N_8485,N_1089,N_353);
nor U8486 (N_8486,N_2009,N_555);
and U8487 (N_8487,N_4227,N_5451);
or U8488 (N_8488,N_2225,N_54);
nand U8489 (N_8489,N_1524,N_876);
nand U8490 (N_8490,N_1885,N_1481);
nor U8491 (N_8491,N_4946,N_1769);
xor U8492 (N_8492,N_713,N_2327);
xor U8493 (N_8493,N_4079,N_3946);
xor U8494 (N_8494,N_4627,N_5993);
nor U8495 (N_8495,N_4925,N_3044);
nand U8496 (N_8496,N_2486,N_3799);
or U8497 (N_8497,N_1460,N_1553);
nand U8498 (N_8498,N_4603,N_5484);
nor U8499 (N_8499,N_3482,N_500);
nor U8500 (N_8500,N_5470,N_5973);
xnor U8501 (N_8501,N_4880,N_3582);
nand U8502 (N_8502,N_140,N_1522);
xor U8503 (N_8503,N_4111,N_4115);
nor U8504 (N_8504,N_3604,N_1982);
xor U8505 (N_8505,N_3145,N_3784);
nand U8506 (N_8506,N_402,N_3429);
nor U8507 (N_8507,N_2730,N_1923);
and U8508 (N_8508,N_5152,N_4193);
or U8509 (N_8509,N_314,N_3523);
and U8510 (N_8510,N_330,N_2341);
nand U8511 (N_8511,N_5994,N_3457);
xor U8512 (N_8512,N_3680,N_226);
and U8513 (N_8513,N_4445,N_1427);
nor U8514 (N_8514,N_2892,N_180);
nor U8515 (N_8515,N_2776,N_2303);
nor U8516 (N_8516,N_4206,N_4965);
nand U8517 (N_8517,N_4406,N_4868);
nor U8518 (N_8518,N_1704,N_445);
and U8519 (N_8519,N_2893,N_3456);
nand U8520 (N_8520,N_2522,N_1163);
xnor U8521 (N_8521,N_2154,N_2014);
and U8522 (N_8522,N_2941,N_2420);
nand U8523 (N_8523,N_3232,N_5846);
xor U8524 (N_8524,N_4122,N_4818);
xnor U8525 (N_8525,N_5988,N_2437);
and U8526 (N_8526,N_3769,N_2468);
xor U8527 (N_8527,N_3480,N_148);
and U8528 (N_8528,N_3876,N_1640);
and U8529 (N_8529,N_3666,N_3858);
or U8530 (N_8530,N_3810,N_2306);
and U8531 (N_8531,N_3302,N_426);
xnor U8532 (N_8532,N_2010,N_4532);
nand U8533 (N_8533,N_5729,N_1544);
nand U8534 (N_8534,N_3578,N_189);
nor U8535 (N_8535,N_4582,N_4540);
xor U8536 (N_8536,N_590,N_4134);
or U8537 (N_8537,N_5185,N_1725);
nor U8538 (N_8538,N_3780,N_5591);
and U8539 (N_8539,N_1505,N_771);
and U8540 (N_8540,N_988,N_1250);
xor U8541 (N_8541,N_5801,N_5621);
xor U8542 (N_8542,N_4383,N_5506);
or U8543 (N_8543,N_196,N_3161);
xnor U8544 (N_8544,N_915,N_2162);
xnor U8545 (N_8545,N_5420,N_468);
or U8546 (N_8546,N_4180,N_5478);
xnor U8547 (N_8547,N_2849,N_4004);
nand U8548 (N_8548,N_2667,N_3187);
nor U8549 (N_8549,N_4065,N_3344);
and U8550 (N_8550,N_5812,N_2449);
or U8551 (N_8551,N_5509,N_5182);
or U8552 (N_8552,N_375,N_4701);
nand U8553 (N_8553,N_2200,N_5469);
nand U8554 (N_8554,N_5295,N_2683);
nand U8555 (N_8555,N_485,N_877);
or U8556 (N_8556,N_1437,N_4494);
nor U8557 (N_8557,N_3445,N_1211);
or U8558 (N_8558,N_4681,N_5387);
or U8559 (N_8559,N_289,N_158);
and U8560 (N_8560,N_961,N_2603);
xor U8561 (N_8561,N_4078,N_5770);
xor U8562 (N_8562,N_5830,N_251);
and U8563 (N_8563,N_5427,N_1009);
or U8564 (N_8564,N_5702,N_1700);
xor U8565 (N_8565,N_3239,N_5473);
xnor U8566 (N_8566,N_5705,N_1333);
nand U8567 (N_8567,N_2412,N_3101);
nand U8568 (N_8568,N_3149,N_5870);
and U8569 (N_8569,N_2828,N_4478);
and U8570 (N_8570,N_5724,N_3206);
nand U8571 (N_8571,N_606,N_2381);
xor U8572 (N_8572,N_3117,N_3240);
xnor U8573 (N_8573,N_1278,N_2865);
and U8574 (N_8574,N_4645,N_530);
and U8575 (N_8575,N_4856,N_5210);
and U8576 (N_8576,N_5243,N_2195);
nor U8577 (N_8577,N_5323,N_4654);
and U8578 (N_8578,N_3489,N_2848);
or U8579 (N_8579,N_5433,N_5695);
xor U8580 (N_8580,N_5779,N_5872);
nand U8581 (N_8581,N_370,N_1946);
nor U8582 (N_8582,N_3169,N_4492);
and U8583 (N_8583,N_2026,N_1339);
nor U8584 (N_8584,N_393,N_5867);
xnor U8585 (N_8585,N_1130,N_210);
or U8586 (N_8586,N_1013,N_2264);
and U8587 (N_8587,N_686,N_1469);
xnor U8588 (N_8588,N_1466,N_1282);
and U8589 (N_8589,N_5448,N_5767);
or U8590 (N_8590,N_800,N_5254);
xor U8591 (N_8591,N_344,N_1299);
and U8592 (N_8592,N_1684,N_3366);
nor U8593 (N_8593,N_870,N_1223);
nand U8594 (N_8594,N_2065,N_4508);
nor U8595 (N_8595,N_3,N_4167);
or U8596 (N_8596,N_5282,N_1644);
and U8597 (N_8597,N_3029,N_3356);
and U8598 (N_8598,N_4667,N_3300);
nor U8599 (N_8599,N_4183,N_1619);
nor U8600 (N_8600,N_1066,N_4266);
or U8601 (N_8601,N_5164,N_609);
xor U8602 (N_8602,N_4911,N_1568);
or U8603 (N_8603,N_1525,N_4960);
and U8604 (N_8604,N_208,N_4171);
or U8605 (N_8605,N_4056,N_4208);
xor U8606 (N_8606,N_4415,N_327);
and U8607 (N_8607,N_5290,N_787);
nor U8608 (N_8608,N_5258,N_4219);
nor U8609 (N_8609,N_5542,N_4425);
nor U8610 (N_8610,N_1253,N_1991);
nand U8611 (N_8611,N_5432,N_5502);
xnor U8612 (N_8612,N_1867,N_5495);
xnor U8613 (N_8613,N_1910,N_5634);
xnor U8614 (N_8614,N_959,N_182);
nor U8615 (N_8615,N_1601,N_128);
and U8616 (N_8616,N_2025,N_12);
nand U8617 (N_8617,N_5077,N_1099);
nand U8618 (N_8618,N_93,N_2189);
xor U8619 (N_8619,N_4889,N_4013);
or U8620 (N_8620,N_1399,N_2160);
nor U8621 (N_8621,N_2705,N_847);
nor U8622 (N_8622,N_143,N_4106);
and U8623 (N_8623,N_3536,N_5858);
xnor U8624 (N_8624,N_3279,N_2256);
or U8625 (N_8625,N_3533,N_1940);
xnor U8626 (N_8626,N_1695,N_3756);
and U8627 (N_8627,N_1170,N_4160);
xnor U8628 (N_8628,N_895,N_5436);
nor U8629 (N_8629,N_2636,N_5489);
nand U8630 (N_8630,N_3477,N_3726);
nor U8631 (N_8631,N_4858,N_4128);
and U8632 (N_8632,N_4859,N_720);
nor U8633 (N_8633,N_2121,N_2153);
and U8634 (N_8634,N_4076,N_267);
xor U8635 (N_8635,N_2992,N_5269);
or U8636 (N_8636,N_3215,N_1438);
and U8637 (N_8637,N_5968,N_5407);
and U8638 (N_8638,N_3175,N_972);
and U8639 (N_8639,N_1037,N_3608);
and U8640 (N_8640,N_2029,N_4231);
xnor U8641 (N_8641,N_4887,N_4034);
and U8642 (N_8642,N_2005,N_4133);
or U8643 (N_8643,N_2982,N_1764);
xor U8644 (N_8644,N_3216,N_2874);
or U8645 (N_8645,N_4688,N_4211);
xnor U8646 (N_8646,N_134,N_2900);
xor U8647 (N_8647,N_4719,N_5562);
nor U8648 (N_8648,N_5171,N_5494);
or U8649 (N_8649,N_2419,N_5025);
or U8650 (N_8650,N_1010,N_3392);
nand U8651 (N_8651,N_5242,N_4904);
and U8652 (N_8652,N_5229,N_4250);
nand U8653 (N_8653,N_3669,N_55);
nand U8654 (N_8654,N_2862,N_2827);
nand U8655 (N_8655,N_5644,N_5588);
or U8656 (N_8656,N_4676,N_1148);
and U8657 (N_8657,N_993,N_5486);
nor U8658 (N_8658,N_57,N_1679);
nor U8659 (N_8659,N_2666,N_1468);
xnor U8660 (N_8660,N_1102,N_4274);
and U8661 (N_8661,N_1623,N_5595);
xnor U8662 (N_8662,N_5939,N_3989);
nor U8663 (N_8663,N_2649,N_1586);
or U8664 (N_8664,N_4483,N_2906);
xnor U8665 (N_8665,N_1976,N_5748);
nor U8666 (N_8666,N_3348,N_3855);
or U8667 (N_8667,N_1666,N_5706);
nor U8668 (N_8668,N_4593,N_2764);
and U8669 (N_8669,N_1447,N_3360);
or U8670 (N_8670,N_5012,N_4035);
xor U8671 (N_8671,N_131,N_1717);
nand U8672 (N_8672,N_3660,N_2027);
xnor U8673 (N_8673,N_4759,N_5245);
xor U8674 (N_8674,N_3152,N_2505);
nand U8675 (N_8675,N_2620,N_1039);
nand U8676 (N_8676,N_443,N_2240);
xnor U8677 (N_8677,N_5549,N_1376);
nor U8678 (N_8678,N_2942,N_1056);
or U8679 (N_8679,N_1218,N_3026);
nor U8680 (N_8680,N_2454,N_230);
or U8681 (N_8681,N_2512,N_1027);
and U8682 (N_8682,N_5640,N_2735);
and U8683 (N_8683,N_3374,N_955);
nor U8684 (N_8684,N_3941,N_2608);
nand U8685 (N_8685,N_2000,N_2336);
nor U8686 (N_8686,N_3673,N_4669);
and U8687 (N_8687,N_2811,N_5208);
nor U8688 (N_8688,N_4671,N_4017);
xor U8689 (N_8689,N_2659,N_2054);
or U8690 (N_8690,N_4336,N_363);
or U8691 (N_8691,N_2346,N_5659);
or U8692 (N_8692,N_1574,N_1635);
nor U8693 (N_8693,N_2899,N_505);
and U8694 (N_8694,N_2521,N_1604);
or U8695 (N_8695,N_4760,N_594);
and U8696 (N_8696,N_3609,N_1811);
or U8697 (N_8697,N_5325,N_108);
xor U8698 (N_8698,N_3412,N_4137);
xor U8699 (N_8699,N_1581,N_2850);
or U8700 (N_8700,N_2875,N_2172);
xor U8701 (N_8701,N_5683,N_58);
and U8702 (N_8702,N_5661,N_3349);
and U8703 (N_8703,N_2721,N_5405);
xnor U8704 (N_8704,N_2533,N_676);
xnor U8705 (N_8705,N_4172,N_48);
nand U8706 (N_8706,N_5117,N_103);
nor U8707 (N_8707,N_5425,N_1509);
xnor U8708 (N_8708,N_5528,N_5163);
or U8709 (N_8709,N_362,N_3678);
nor U8710 (N_8710,N_1082,N_4706);
and U8711 (N_8711,N_3567,N_674);
nand U8712 (N_8712,N_5769,N_4948);
nor U8713 (N_8713,N_1537,N_3791);
and U8714 (N_8714,N_4758,N_1869);
xnor U8715 (N_8715,N_3091,N_2607);
or U8716 (N_8716,N_2082,N_1315);
nor U8717 (N_8717,N_3508,N_1777);
or U8718 (N_8718,N_4402,N_4988);
and U8719 (N_8719,N_3116,N_1127);
nor U8720 (N_8720,N_1762,N_342);
nor U8721 (N_8721,N_607,N_3613);
nor U8722 (N_8722,N_2763,N_466);
nor U8723 (N_8723,N_5954,N_1821);
nor U8724 (N_8724,N_1475,N_2413);
or U8725 (N_8725,N_1805,N_2389);
and U8726 (N_8726,N_969,N_1942);
and U8727 (N_8727,N_3233,N_5777);
and U8728 (N_8728,N_4147,N_2662);
xnor U8729 (N_8729,N_3749,N_4729);
nand U8730 (N_8730,N_2961,N_963);
nor U8731 (N_8731,N_1334,N_5708);
and U8732 (N_8732,N_968,N_4780);
nand U8733 (N_8733,N_3986,N_5843);
nand U8734 (N_8734,N_2638,N_2312);
and U8735 (N_8735,N_2193,N_4349);
nand U8736 (N_8736,N_3610,N_758);
or U8737 (N_8737,N_1780,N_5838);
nand U8738 (N_8738,N_3835,N_4139);
nor U8739 (N_8739,N_1983,N_1059);
and U8740 (N_8740,N_398,N_5900);
nand U8741 (N_8741,N_4832,N_2199);
nand U8742 (N_8742,N_3507,N_4198);
xor U8743 (N_8743,N_5389,N_3776);
xnor U8744 (N_8744,N_3517,N_1072);
or U8745 (N_8745,N_1227,N_4416);
nand U8746 (N_8746,N_1174,N_4519);
xnor U8747 (N_8747,N_1487,N_3566);
and U8748 (N_8748,N_1558,N_5712);
nand U8749 (N_8749,N_3733,N_4479);
xnor U8750 (N_8750,N_4890,N_944);
nand U8751 (N_8751,N_863,N_3486);
or U8752 (N_8752,N_1736,N_937);
xnor U8753 (N_8753,N_1721,N_1655);
nand U8754 (N_8754,N_4221,N_5408);
or U8755 (N_8755,N_4726,N_5952);
xor U8756 (N_8756,N_4607,N_2239);
nand U8757 (N_8757,N_1966,N_5154);
xnor U8758 (N_8758,N_1719,N_1084);
xnor U8759 (N_8759,N_4089,N_3133);
xnor U8760 (N_8760,N_5144,N_3439);
or U8761 (N_8761,N_613,N_933);
nor U8762 (N_8762,N_4604,N_4444);
nor U8763 (N_8763,N_5102,N_2269);
or U8764 (N_8764,N_5583,N_5851);
or U8765 (N_8765,N_1356,N_2115);
nor U8766 (N_8766,N_738,N_346);
or U8767 (N_8767,N_354,N_2558);
nand U8768 (N_8768,N_852,N_4529);
or U8769 (N_8769,N_1998,N_5951);
or U8770 (N_8770,N_855,N_694);
nor U8771 (N_8771,N_391,N_4475);
nand U8772 (N_8772,N_1849,N_3453);
xor U8773 (N_8773,N_2781,N_3830);
nor U8774 (N_8774,N_966,N_1083);
nand U8775 (N_8775,N_3113,N_202);
or U8776 (N_8776,N_628,N_4657);
and U8777 (N_8777,N_495,N_619);
xnor U8778 (N_8778,N_2247,N_3961);
nand U8779 (N_8779,N_4909,N_165);
and U8780 (N_8780,N_1796,N_3854);
nor U8781 (N_8781,N_5476,N_400);
and U8782 (N_8782,N_4812,N_3529);
xor U8783 (N_8783,N_1141,N_5442);
nor U8784 (N_8784,N_811,N_5195);
or U8785 (N_8785,N_129,N_170);
and U8786 (N_8786,N_2719,N_2969);
xnor U8787 (N_8787,N_5550,N_2944);
and U8788 (N_8788,N_4528,N_5133);
xnor U8789 (N_8789,N_4872,N_719);
xor U8790 (N_8790,N_1323,N_932);
nor U8791 (N_8791,N_1192,N_4420);
xor U8792 (N_8792,N_4006,N_2574);
or U8793 (N_8793,N_1836,N_3565);
and U8794 (N_8794,N_5647,N_1064);
nand U8795 (N_8795,N_1681,N_242);
nand U8796 (N_8796,N_2669,N_1593);
xor U8797 (N_8797,N_4902,N_5106);
or U8798 (N_8798,N_4095,N_3034);
and U8799 (N_8799,N_1405,N_5081);
or U8800 (N_8800,N_2489,N_3087);
nand U8801 (N_8801,N_5137,N_4358);
nand U8802 (N_8802,N_1570,N_4648);
or U8803 (N_8803,N_64,N_3270);
xnor U8804 (N_8804,N_710,N_3122);
nand U8805 (N_8805,N_4713,N_168);
and U8806 (N_8806,N_3194,N_869);
or U8807 (N_8807,N_3908,N_396);
nand U8808 (N_8808,N_1291,N_4762);
and U8809 (N_8809,N_5418,N_1332);
xnor U8810 (N_8810,N_2946,N_3066);
nor U8811 (N_8811,N_2569,N_5039);
nand U8812 (N_8812,N_4775,N_3706);
nor U8813 (N_8813,N_3912,N_3764);
nand U8814 (N_8814,N_1347,N_5612);
and U8815 (N_8815,N_3363,N_5523);
nor U8816 (N_8816,N_5445,N_3767);
xor U8817 (N_8817,N_5516,N_1293);
nor U8818 (N_8818,N_2452,N_1705);
nor U8819 (N_8819,N_3883,N_290);
and U8820 (N_8820,N_233,N_2789);
nor U8821 (N_8821,N_3037,N_2238);
and U8822 (N_8822,N_733,N_4457);
nor U8823 (N_8823,N_4795,N_991);
and U8824 (N_8824,N_1495,N_457);
xnor U8825 (N_8825,N_4910,N_644);
xnor U8826 (N_8826,N_5492,N_4836);
and U8827 (N_8827,N_5123,N_3083);
nand U8828 (N_8828,N_1546,N_2526);
and U8829 (N_8829,N_3140,N_3128);
xnor U8830 (N_8830,N_2150,N_5055);
and U8831 (N_8831,N_5034,N_4329);
or U8832 (N_8832,N_4993,N_3575);
nor U8833 (N_8833,N_1738,N_5792);
nand U8834 (N_8834,N_1490,N_5886);
nand U8835 (N_8835,N_4620,N_2268);
and U8836 (N_8836,N_4757,N_1235);
xnor U8837 (N_8837,N_4011,N_1136);
or U8838 (N_8838,N_3334,N_366);
and U8839 (N_8839,N_964,N_5526);
xor U8840 (N_8840,N_244,N_3282);
and U8841 (N_8841,N_5499,N_5848);
nand U8842 (N_8842,N_5223,N_1132);
nand U8843 (N_8843,N_5784,N_2443);
and U8844 (N_8844,N_2309,N_5722);
xnor U8845 (N_8845,N_2637,N_5392);
nor U8846 (N_8846,N_2718,N_2273);
or U8847 (N_8847,N_4327,N_3493);
and U8848 (N_8848,N_1563,N_3134);
or U8849 (N_8849,N_124,N_2956);
xnor U8850 (N_8850,N_286,N_4197);
and U8851 (N_8851,N_3451,N_673);
or U8852 (N_8852,N_5751,N_1248);
and U8853 (N_8853,N_5380,N_5849);
xnor U8854 (N_8854,N_1671,N_920);
xor U8855 (N_8855,N_5592,N_1930);
nand U8856 (N_8856,N_604,N_1694);
nand U8857 (N_8857,N_4153,N_1319);
nand U8858 (N_8858,N_1961,N_4157);
or U8859 (N_8859,N_4498,N_4068);
and U8860 (N_8860,N_5953,N_1190);
and U8861 (N_8861,N_3474,N_1540);
nand U8862 (N_8862,N_238,N_313);
xor U8863 (N_8863,N_5556,N_3242);
nor U8864 (N_8864,N_414,N_4500);
xor U8865 (N_8865,N_4489,N_4879);
and U8866 (N_8866,N_1816,N_1499);
or U8867 (N_8867,N_5377,N_300);
xnor U8868 (N_8868,N_4768,N_794);
and U8869 (N_8869,N_2459,N_2965);
xnor U8870 (N_8870,N_469,N_650);
nor U8871 (N_8871,N_5814,N_5419);
nor U8872 (N_8872,N_1531,N_2538);
and U8873 (N_8873,N_5989,N_2197);
or U8874 (N_8874,N_4962,N_2616);
xnor U8875 (N_8875,N_1204,N_360);
or U8876 (N_8876,N_3914,N_301);
or U8877 (N_8877,N_32,N_5658);
xor U8878 (N_8878,N_5935,N_427);
or U8879 (N_8879,N_1729,N_880);
and U8880 (N_8880,N_31,N_434);
xnor U8881 (N_8881,N_3798,N_1547);
or U8882 (N_8882,N_652,N_2738);
and U8883 (N_8883,N_1448,N_1267);
or U8884 (N_8884,N_3384,N_3848);
nor U8885 (N_8885,N_5286,N_5629);
or U8886 (N_8886,N_1216,N_3895);
nor U8887 (N_8887,N_729,N_2585);
nor U8888 (N_8888,N_2655,N_1611);
and U8889 (N_8889,N_2171,N_4891);
nor U8890 (N_8890,N_2935,N_1536);
xnor U8891 (N_8891,N_4467,N_5944);
nand U8892 (N_8892,N_1421,N_2588);
and U8893 (N_8893,N_130,N_3528);
nand U8894 (N_8894,N_2432,N_5536);
and U8895 (N_8895,N_5680,N_3707);
and U8896 (N_8896,N_3450,N_2129);
xnor U8897 (N_8897,N_3642,N_4510);
nor U8898 (N_8898,N_625,N_4379);
xnor U8899 (N_8899,N_4361,N_2287);
and U8900 (N_8900,N_2466,N_2653);
nand U8901 (N_8901,N_4635,N_3246);
xor U8902 (N_8902,N_1012,N_5713);
and U8903 (N_8903,N_2592,N_5904);
or U8904 (N_8904,N_4687,N_3454);
nor U8905 (N_8905,N_3750,N_3935);
nor U8906 (N_8906,N_4682,N_265);
nor U8907 (N_8907,N_2931,N_1945);
and U8908 (N_8908,N_5503,N_1164);
or U8909 (N_8909,N_4194,N_1925);
nand U8910 (N_8910,N_3146,N_4707);
nor U8911 (N_8911,N_1847,N_2105);
nor U8912 (N_8912,N_2832,N_5931);
xnor U8913 (N_8913,N_367,N_2191);
or U8914 (N_8914,N_2733,N_5942);
and U8915 (N_8915,N_1464,N_5187);
and U8916 (N_8916,N_4680,N_101);
or U8917 (N_8917,N_1473,N_2928);
xor U8918 (N_8918,N_4831,N_3657);
and U8919 (N_8919,N_4679,N_4091);
nor U8920 (N_8920,N_5326,N_3558);
nor U8921 (N_8921,N_4931,N_4014);
nand U8922 (N_8922,N_2778,N_2471);
and U8923 (N_8923,N_4554,N_4495);
and U8924 (N_8924,N_1006,N_1042);
and U8925 (N_8925,N_2504,N_4717);
nand U8926 (N_8926,N_3850,N_1693);
and U8927 (N_8927,N_2058,N_4316);
and U8928 (N_8928,N_2994,N_3740);
xnor U8929 (N_8929,N_4693,N_777);
xor U8930 (N_8930,N_910,N_2379);
xor U8931 (N_8931,N_5023,N_3498);
xor U8932 (N_8932,N_2877,N_1814);
or U8933 (N_8933,N_816,N_2744);
nor U8934 (N_8934,N_248,N_4041);
and U8935 (N_8935,N_4613,N_3861);
xnor U8936 (N_8936,N_2564,N_5676);
or U8937 (N_8937,N_2012,N_3730);
nor U8938 (N_8938,N_5349,N_3085);
nand U8939 (N_8939,N_514,N_3687);
and U8940 (N_8940,N_3402,N_1791);
xnor U8941 (N_8941,N_5663,N_195);
xor U8942 (N_8942,N_4587,N_3046);
or U8943 (N_8943,N_5441,N_3624);
and U8944 (N_8944,N_236,N_2422);
nor U8945 (N_8945,N_3459,N_3262);
nor U8946 (N_8946,N_1026,N_2822);
nand U8947 (N_8947,N_5928,N_2530);
or U8948 (N_8948,N_2013,N_3126);
and U8949 (N_8949,N_700,N_5631);
xor U8950 (N_8950,N_1262,N_1277);
nand U8951 (N_8951,N_2697,N_4614);
nand U8952 (N_8952,N_299,N_2796);
nor U8953 (N_8953,N_36,N_4061);
or U8954 (N_8954,N_4364,N_5796);
and U8955 (N_8955,N_3247,N_446);
and U8956 (N_8956,N_1703,N_527);
xor U8957 (N_8957,N_1140,N_3893);
nand U8958 (N_8958,N_3834,N_2746);
and U8959 (N_8959,N_3394,N_5949);
nand U8960 (N_8960,N_5430,N_1142);
nand U8961 (N_8961,N_4321,N_4066);
nand U8962 (N_8962,N_2884,N_4323);
nor U8963 (N_8963,N_1995,N_1958);
xnor U8964 (N_8964,N_4114,N_509);
nand U8965 (N_8965,N_4866,N_1975);
xor U8966 (N_8966,N_2474,N_3404);
nor U8967 (N_8967,N_2143,N_1379);
nand U8968 (N_8968,N_4502,N_5718);
xor U8969 (N_8969,N_715,N_3288);
nand U8970 (N_8970,N_5882,N_4906);
and U8971 (N_8971,N_1373,N_2194);
or U8972 (N_8972,N_3271,N_5031);
nand U8973 (N_8973,N_3695,N_1832);
nor U8974 (N_8974,N_2897,N_234);
xnor U8975 (N_8975,N_5328,N_3878);
and U8976 (N_8976,N_3476,N_315);
nor U8977 (N_8977,N_1733,N_5570);
and U8978 (N_8978,N_1911,N_3501);
or U8979 (N_8979,N_3771,N_98);
or U8980 (N_8980,N_4875,N_5004);
and U8981 (N_8981,N_1314,N_5999);
or U8982 (N_8982,N_4571,N_1974);
nand U8983 (N_8983,N_3357,N_4214);
xor U8984 (N_8984,N_5437,N_3119);
or U8985 (N_8985,N_2611,N_922);
xor U8986 (N_8986,N_2534,N_3106);
nand U8987 (N_8987,N_2231,N_1837);
nor U8988 (N_8988,N_1168,N_4749);
or U8989 (N_8989,N_5464,N_1774);
xnor U8990 (N_8990,N_5162,N_2246);
nor U8991 (N_8991,N_3988,N_3967);
xor U8992 (N_8992,N_1078,N_5960);
and U8993 (N_8993,N_1077,N_4022);
nand U8994 (N_8994,N_3712,N_5512);
or U8995 (N_8995,N_4884,N_3209);
nand U8996 (N_8996,N_5524,N_3150);
nand U8997 (N_8997,N_762,N_4202);
and U8998 (N_8998,N_5633,N_4315);
nor U8999 (N_8999,N_2008,N_4187);
xor U9000 (N_9000,N_2603,N_4977);
nand U9001 (N_9001,N_560,N_249);
xor U9002 (N_9002,N_2253,N_2133);
or U9003 (N_9003,N_231,N_3118);
nand U9004 (N_9004,N_5574,N_5537);
nand U9005 (N_9005,N_3608,N_5669);
or U9006 (N_9006,N_5443,N_1775);
xnor U9007 (N_9007,N_1111,N_4381);
nor U9008 (N_9008,N_5395,N_3510);
or U9009 (N_9009,N_786,N_3483);
xor U9010 (N_9010,N_2191,N_5906);
or U9011 (N_9011,N_4004,N_4969);
nand U9012 (N_9012,N_4595,N_4686);
xnor U9013 (N_9013,N_5674,N_771);
nor U9014 (N_9014,N_2743,N_1533);
xnor U9015 (N_9015,N_237,N_1229);
nor U9016 (N_9016,N_5558,N_1303);
or U9017 (N_9017,N_4825,N_5589);
and U9018 (N_9018,N_2844,N_3698);
xor U9019 (N_9019,N_212,N_3347);
or U9020 (N_9020,N_5638,N_2124);
and U9021 (N_9021,N_5258,N_964);
nor U9022 (N_9022,N_3702,N_4458);
and U9023 (N_9023,N_3993,N_2917);
and U9024 (N_9024,N_1874,N_2932);
xnor U9025 (N_9025,N_4191,N_2827);
or U9026 (N_9026,N_1815,N_2447);
nand U9027 (N_9027,N_2075,N_362);
nor U9028 (N_9028,N_2831,N_5406);
nor U9029 (N_9029,N_1216,N_2860);
nand U9030 (N_9030,N_3972,N_5821);
nand U9031 (N_9031,N_2451,N_2679);
and U9032 (N_9032,N_4158,N_3726);
xor U9033 (N_9033,N_981,N_4018);
nand U9034 (N_9034,N_3881,N_3531);
xor U9035 (N_9035,N_965,N_4471);
xnor U9036 (N_9036,N_3085,N_1229);
or U9037 (N_9037,N_3637,N_5967);
xnor U9038 (N_9038,N_1649,N_3027);
xnor U9039 (N_9039,N_3414,N_970);
nand U9040 (N_9040,N_232,N_4949);
or U9041 (N_9041,N_3603,N_1888);
or U9042 (N_9042,N_4541,N_2655);
nor U9043 (N_9043,N_1974,N_5414);
nor U9044 (N_9044,N_3903,N_4917);
xor U9045 (N_9045,N_2416,N_1719);
xnor U9046 (N_9046,N_2820,N_2277);
or U9047 (N_9047,N_346,N_891);
nand U9048 (N_9048,N_5122,N_2008);
or U9049 (N_9049,N_2666,N_1465);
nor U9050 (N_9050,N_5660,N_5796);
or U9051 (N_9051,N_2592,N_4832);
nand U9052 (N_9052,N_4925,N_5591);
xnor U9053 (N_9053,N_5312,N_1457);
nand U9054 (N_9054,N_1414,N_3880);
and U9055 (N_9055,N_613,N_3862);
or U9056 (N_9056,N_4991,N_3908);
or U9057 (N_9057,N_3484,N_2026);
xor U9058 (N_9058,N_4631,N_745);
nand U9059 (N_9059,N_2148,N_1189);
nor U9060 (N_9060,N_2046,N_4644);
xnor U9061 (N_9061,N_3196,N_5336);
or U9062 (N_9062,N_4973,N_792);
nand U9063 (N_9063,N_5874,N_3550);
xnor U9064 (N_9064,N_4483,N_583);
nor U9065 (N_9065,N_1328,N_3902);
nand U9066 (N_9066,N_237,N_3427);
nor U9067 (N_9067,N_5072,N_3151);
nand U9068 (N_9068,N_4254,N_5421);
and U9069 (N_9069,N_4998,N_2192);
or U9070 (N_9070,N_4770,N_1164);
nor U9071 (N_9071,N_1593,N_958);
or U9072 (N_9072,N_3045,N_2279);
and U9073 (N_9073,N_2237,N_5678);
and U9074 (N_9074,N_5818,N_3983);
and U9075 (N_9075,N_5049,N_3800);
and U9076 (N_9076,N_2726,N_289);
nor U9077 (N_9077,N_2633,N_2183);
xor U9078 (N_9078,N_2569,N_439);
xor U9079 (N_9079,N_1142,N_5633);
and U9080 (N_9080,N_5772,N_5113);
xor U9081 (N_9081,N_3599,N_140);
nand U9082 (N_9082,N_4061,N_2175);
nand U9083 (N_9083,N_2371,N_4252);
nand U9084 (N_9084,N_1289,N_2020);
and U9085 (N_9085,N_3294,N_129);
xnor U9086 (N_9086,N_5699,N_3431);
and U9087 (N_9087,N_4446,N_4787);
nor U9088 (N_9088,N_1380,N_4967);
nand U9089 (N_9089,N_346,N_5762);
nor U9090 (N_9090,N_2068,N_4918);
nand U9091 (N_9091,N_5323,N_2182);
nand U9092 (N_9092,N_3083,N_853);
nor U9093 (N_9093,N_1245,N_1568);
xor U9094 (N_9094,N_5310,N_3961);
nor U9095 (N_9095,N_22,N_1862);
nor U9096 (N_9096,N_921,N_1118);
nand U9097 (N_9097,N_4735,N_3831);
xor U9098 (N_9098,N_5114,N_3769);
and U9099 (N_9099,N_3613,N_565);
or U9100 (N_9100,N_4316,N_3040);
nand U9101 (N_9101,N_4661,N_2189);
nand U9102 (N_9102,N_5469,N_3202);
xor U9103 (N_9103,N_1203,N_341);
nor U9104 (N_9104,N_1295,N_1806);
nor U9105 (N_9105,N_3292,N_1759);
nor U9106 (N_9106,N_3723,N_880);
xor U9107 (N_9107,N_1136,N_3420);
nor U9108 (N_9108,N_2883,N_4696);
and U9109 (N_9109,N_649,N_1242);
xnor U9110 (N_9110,N_1659,N_5621);
or U9111 (N_9111,N_5453,N_3073);
and U9112 (N_9112,N_3839,N_1663);
nor U9113 (N_9113,N_5734,N_5352);
or U9114 (N_9114,N_1669,N_1407);
or U9115 (N_9115,N_4720,N_4128);
and U9116 (N_9116,N_34,N_2300);
nand U9117 (N_9117,N_4720,N_1003);
nor U9118 (N_9118,N_1222,N_5360);
nand U9119 (N_9119,N_2719,N_4525);
xor U9120 (N_9120,N_4443,N_4041);
nor U9121 (N_9121,N_1923,N_2899);
and U9122 (N_9122,N_80,N_3084);
and U9123 (N_9123,N_1054,N_2069);
nor U9124 (N_9124,N_1895,N_3797);
xnor U9125 (N_9125,N_2182,N_4217);
nand U9126 (N_9126,N_4580,N_3116);
nand U9127 (N_9127,N_5053,N_528);
or U9128 (N_9128,N_2852,N_926);
nand U9129 (N_9129,N_2000,N_3860);
nor U9130 (N_9130,N_2809,N_5511);
or U9131 (N_9131,N_2907,N_2555);
or U9132 (N_9132,N_1257,N_1815);
nand U9133 (N_9133,N_1330,N_3761);
and U9134 (N_9134,N_3250,N_4775);
xor U9135 (N_9135,N_1540,N_3884);
or U9136 (N_9136,N_4634,N_528);
xnor U9137 (N_9137,N_2722,N_5693);
xor U9138 (N_9138,N_1904,N_124);
and U9139 (N_9139,N_2841,N_2724);
nor U9140 (N_9140,N_3674,N_3613);
nor U9141 (N_9141,N_3278,N_5359);
xnor U9142 (N_9142,N_1517,N_1338);
or U9143 (N_9143,N_4361,N_2909);
nor U9144 (N_9144,N_4467,N_5829);
nor U9145 (N_9145,N_5251,N_1840);
nor U9146 (N_9146,N_3799,N_368);
and U9147 (N_9147,N_2436,N_467);
nor U9148 (N_9148,N_3281,N_1081);
or U9149 (N_9149,N_5691,N_2889);
nor U9150 (N_9150,N_2388,N_805);
nor U9151 (N_9151,N_3748,N_1731);
xor U9152 (N_9152,N_3570,N_4772);
or U9153 (N_9153,N_1001,N_4313);
or U9154 (N_9154,N_4798,N_3453);
nand U9155 (N_9155,N_28,N_1984);
and U9156 (N_9156,N_4134,N_3264);
or U9157 (N_9157,N_536,N_2330);
and U9158 (N_9158,N_1493,N_5288);
or U9159 (N_9159,N_3748,N_3462);
or U9160 (N_9160,N_3488,N_2282);
nand U9161 (N_9161,N_3084,N_2650);
xor U9162 (N_9162,N_730,N_4576);
nor U9163 (N_9163,N_88,N_71);
nor U9164 (N_9164,N_3110,N_4707);
nor U9165 (N_9165,N_5626,N_4353);
and U9166 (N_9166,N_953,N_4094);
nor U9167 (N_9167,N_1879,N_2622);
xor U9168 (N_9168,N_2833,N_2298);
nand U9169 (N_9169,N_4267,N_2155);
xnor U9170 (N_9170,N_5975,N_4386);
nand U9171 (N_9171,N_5190,N_3630);
nor U9172 (N_9172,N_5189,N_4354);
xor U9173 (N_9173,N_5406,N_5363);
or U9174 (N_9174,N_3107,N_5612);
and U9175 (N_9175,N_5215,N_2752);
and U9176 (N_9176,N_4730,N_3574);
nor U9177 (N_9177,N_1532,N_3646);
and U9178 (N_9178,N_4377,N_5049);
and U9179 (N_9179,N_4698,N_5869);
nand U9180 (N_9180,N_2168,N_4696);
and U9181 (N_9181,N_1950,N_3119);
or U9182 (N_9182,N_472,N_5281);
nand U9183 (N_9183,N_2488,N_418);
xnor U9184 (N_9184,N_5932,N_2427);
nor U9185 (N_9185,N_5311,N_611);
nor U9186 (N_9186,N_4957,N_4502);
and U9187 (N_9187,N_4938,N_2557);
nand U9188 (N_9188,N_165,N_133);
and U9189 (N_9189,N_5217,N_1556);
or U9190 (N_9190,N_1590,N_1076);
or U9191 (N_9191,N_5974,N_3312);
xnor U9192 (N_9192,N_4994,N_2697);
xnor U9193 (N_9193,N_579,N_1531);
nor U9194 (N_9194,N_737,N_1063);
nand U9195 (N_9195,N_3657,N_2248);
and U9196 (N_9196,N_1276,N_594);
and U9197 (N_9197,N_2773,N_2568);
nor U9198 (N_9198,N_5010,N_5799);
xor U9199 (N_9199,N_4981,N_4821);
xnor U9200 (N_9200,N_2481,N_4727);
xor U9201 (N_9201,N_2889,N_1262);
nor U9202 (N_9202,N_2040,N_2563);
nand U9203 (N_9203,N_3238,N_180);
nand U9204 (N_9204,N_2081,N_3018);
xnor U9205 (N_9205,N_5854,N_868);
nor U9206 (N_9206,N_2994,N_1106);
nand U9207 (N_9207,N_5536,N_2578);
and U9208 (N_9208,N_1774,N_4909);
xnor U9209 (N_9209,N_2639,N_3316);
or U9210 (N_9210,N_62,N_4759);
or U9211 (N_9211,N_878,N_2154);
and U9212 (N_9212,N_1554,N_3706);
nand U9213 (N_9213,N_5523,N_4379);
and U9214 (N_9214,N_2670,N_5926);
nor U9215 (N_9215,N_3968,N_5491);
and U9216 (N_9216,N_4350,N_4802);
xnor U9217 (N_9217,N_1978,N_2074);
nor U9218 (N_9218,N_373,N_5378);
or U9219 (N_9219,N_730,N_2866);
and U9220 (N_9220,N_4939,N_2346);
nor U9221 (N_9221,N_1481,N_4326);
nor U9222 (N_9222,N_254,N_4552);
and U9223 (N_9223,N_1209,N_1200);
and U9224 (N_9224,N_2998,N_2109);
xor U9225 (N_9225,N_112,N_4393);
and U9226 (N_9226,N_4008,N_5920);
xnor U9227 (N_9227,N_3038,N_3583);
nand U9228 (N_9228,N_3766,N_2149);
xor U9229 (N_9229,N_223,N_5098);
and U9230 (N_9230,N_1196,N_4275);
xor U9231 (N_9231,N_4429,N_2136);
or U9232 (N_9232,N_1183,N_3153);
nor U9233 (N_9233,N_1246,N_361);
xnor U9234 (N_9234,N_2514,N_3165);
xor U9235 (N_9235,N_2655,N_1874);
xor U9236 (N_9236,N_5033,N_4578);
xnor U9237 (N_9237,N_5673,N_1295);
or U9238 (N_9238,N_2036,N_2849);
xor U9239 (N_9239,N_4553,N_2699);
and U9240 (N_9240,N_2386,N_3428);
nor U9241 (N_9241,N_1140,N_820);
or U9242 (N_9242,N_1503,N_5473);
nand U9243 (N_9243,N_837,N_2068);
nand U9244 (N_9244,N_5092,N_4239);
nand U9245 (N_9245,N_1567,N_2178);
and U9246 (N_9246,N_1162,N_3314);
xor U9247 (N_9247,N_2248,N_1754);
and U9248 (N_9248,N_5387,N_42);
and U9249 (N_9249,N_1061,N_4527);
xnor U9250 (N_9250,N_2132,N_2570);
nor U9251 (N_9251,N_1183,N_3928);
nand U9252 (N_9252,N_3957,N_3466);
xnor U9253 (N_9253,N_4840,N_5830);
or U9254 (N_9254,N_5485,N_3542);
or U9255 (N_9255,N_2578,N_27);
nor U9256 (N_9256,N_426,N_3527);
xnor U9257 (N_9257,N_3580,N_2687);
or U9258 (N_9258,N_2307,N_1525);
or U9259 (N_9259,N_1204,N_309);
nand U9260 (N_9260,N_1147,N_1711);
nor U9261 (N_9261,N_7,N_2532);
nor U9262 (N_9262,N_1147,N_5418);
xor U9263 (N_9263,N_3296,N_2771);
xnor U9264 (N_9264,N_921,N_541);
or U9265 (N_9265,N_5348,N_4429);
and U9266 (N_9266,N_671,N_1106);
nand U9267 (N_9267,N_4824,N_3654);
or U9268 (N_9268,N_714,N_2151);
xor U9269 (N_9269,N_3547,N_4702);
nand U9270 (N_9270,N_3889,N_2142);
xnor U9271 (N_9271,N_368,N_1357);
nor U9272 (N_9272,N_1081,N_3406);
and U9273 (N_9273,N_3122,N_2741);
xnor U9274 (N_9274,N_5805,N_4219);
xnor U9275 (N_9275,N_1410,N_3258);
xnor U9276 (N_9276,N_5410,N_5948);
xnor U9277 (N_9277,N_2837,N_834);
nor U9278 (N_9278,N_1122,N_576);
or U9279 (N_9279,N_1,N_3823);
nand U9280 (N_9280,N_1136,N_3718);
and U9281 (N_9281,N_1596,N_1006);
or U9282 (N_9282,N_4969,N_2455);
xnor U9283 (N_9283,N_2799,N_3397);
nor U9284 (N_9284,N_2912,N_2949);
and U9285 (N_9285,N_4015,N_1306);
and U9286 (N_9286,N_3684,N_1565);
nor U9287 (N_9287,N_3731,N_2574);
or U9288 (N_9288,N_4404,N_3302);
or U9289 (N_9289,N_4213,N_2956);
nor U9290 (N_9290,N_5440,N_2908);
and U9291 (N_9291,N_4786,N_1301);
or U9292 (N_9292,N_315,N_2192);
and U9293 (N_9293,N_4687,N_3896);
nor U9294 (N_9294,N_4712,N_3933);
nand U9295 (N_9295,N_5917,N_5615);
or U9296 (N_9296,N_5911,N_4745);
or U9297 (N_9297,N_2233,N_1522);
or U9298 (N_9298,N_2351,N_3918);
nor U9299 (N_9299,N_4139,N_532);
xor U9300 (N_9300,N_666,N_2984);
nand U9301 (N_9301,N_3046,N_509);
xor U9302 (N_9302,N_1435,N_302);
nor U9303 (N_9303,N_3394,N_5495);
or U9304 (N_9304,N_5133,N_2813);
and U9305 (N_9305,N_4072,N_3786);
and U9306 (N_9306,N_1568,N_59);
and U9307 (N_9307,N_1900,N_3896);
and U9308 (N_9308,N_4742,N_484);
and U9309 (N_9309,N_1090,N_5554);
xor U9310 (N_9310,N_1503,N_2592);
xor U9311 (N_9311,N_2902,N_1079);
and U9312 (N_9312,N_5949,N_492);
nand U9313 (N_9313,N_3525,N_52);
nor U9314 (N_9314,N_1036,N_1637);
nand U9315 (N_9315,N_3096,N_2715);
xor U9316 (N_9316,N_4767,N_754);
xor U9317 (N_9317,N_1430,N_3483);
and U9318 (N_9318,N_3425,N_3720);
nor U9319 (N_9319,N_159,N_5262);
nor U9320 (N_9320,N_4286,N_1776);
xnor U9321 (N_9321,N_4572,N_5106);
or U9322 (N_9322,N_3530,N_2579);
xor U9323 (N_9323,N_3098,N_4164);
and U9324 (N_9324,N_1939,N_1299);
nand U9325 (N_9325,N_5264,N_5379);
xnor U9326 (N_9326,N_4906,N_3572);
nor U9327 (N_9327,N_2803,N_5196);
nor U9328 (N_9328,N_4959,N_2018);
nor U9329 (N_9329,N_3853,N_1036);
or U9330 (N_9330,N_4090,N_5518);
nor U9331 (N_9331,N_5795,N_3413);
nand U9332 (N_9332,N_1876,N_1012);
nand U9333 (N_9333,N_283,N_1112);
and U9334 (N_9334,N_2312,N_1401);
or U9335 (N_9335,N_4325,N_2802);
xnor U9336 (N_9336,N_3574,N_4987);
or U9337 (N_9337,N_4095,N_2547);
and U9338 (N_9338,N_840,N_1263);
and U9339 (N_9339,N_251,N_5784);
or U9340 (N_9340,N_3148,N_1651);
nor U9341 (N_9341,N_4068,N_3964);
xor U9342 (N_9342,N_5226,N_5583);
nor U9343 (N_9343,N_3675,N_3822);
or U9344 (N_9344,N_3109,N_2168);
and U9345 (N_9345,N_4780,N_813);
or U9346 (N_9346,N_4097,N_4282);
or U9347 (N_9347,N_1709,N_2608);
and U9348 (N_9348,N_2593,N_345);
nand U9349 (N_9349,N_4924,N_5502);
or U9350 (N_9350,N_5994,N_2221);
nor U9351 (N_9351,N_4613,N_1989);
and U9352 (N_9352,N_3696,N_5925);
xor U9353 (N_9353,N_4989,N_4170);
nand U9354 (N_9354,N_3535,N_4428);
nor U9355 (N_9355,N_5440,N_4465);
xor U9356 (N_9356,N_4775,N_2957);
nor U9357 (N_9357,N_1247,N_4317);
nand U9358 (N_9358,N_4042,N_1055);
and U9359 (N_9359,N_1607,N_4902);
and U9360 (N_9360,N_1279,N_1529);
or U9361 (N_9361,N_5026,N_4565);
nand U9362 (N_9362,N_1500,N_3327);
nor U9363 (N_9363,N_1607,N_5588);
xor U9364 (N_9364,N_644,N_2434);
or U9365 (N_9365,N_1069,N_3506);
nand U9366 (N_9366,N_5819,N_4185);
nand U9367 (N_9367,N_2248,N_4293);
nor U9368 (N_9368,N_5636,N_1313);
or U9369 (N_9369,N_3498,N_2707);
nor U9370 (N_9370,N_5670,N_2115);
xor U9371 (N_9371,N_4674,N_3936);
nor U9372 (N_9372,N_5702,N_5115);
or U9373 (N_9373,N_1976,N_1462);
nand U9374 (N_9374,N_4352,N_4284);
and U9375 (N_9375,N_5387,N_791);
nand U9376 (N_9376,N_1818,N_4335);
xnor U9377 (N_9377,N_1249,N_54);
and U9378 (N_9378,N_5342,N_3642);
nand U9379 (N_9379,N_207,N_47);
nor U9380 (N_9380,N_5847,N_505);
xnor U9381 (N_9381,N_4989,N_4123);
xor U9382 (N_9382,N_4667,N_1634);
nor U9383 (N_9383,N_4635,N_1800);
or U9384 (N_9384,N_5829,N_5084);
or U9385 (N_9385,N_86,N_965);
xnor U9386 (N_9386,N_5190,N_3355);
xor U9387 (N_9387,N_1136,N_4704);
xor U9388 (N_9388,N_3443,N_2855);
or U9389 (N_9389,N_4976,N_1695);
nand U9390 (N_9390,N_5839,N_5037);
nor U9391 (N_9391,N_3387,N_626);
nand U9392 (N_9392,N_3599,N_5485);
xnor U9393 (N_9393,N_838,N_4202);
and U9394 (N_9394,N_2340,N_5689);
nand U9395 (N_9395,N_2315,N_3482);
and U9396 (N_9396,N_2703,N_1223);
nand U9397 (N_9397,N_3273,N_353);
and U9398 (N_9398,N_2792,N_5112);
nand U9399 (N_9399,N_1893,N_3553);
xor U9400 (N_9400,N_634,N_5051);
nor U9401 (N_9401,N_4032,N_3622);
xnor U9402 (N_9402,N_2531,N_3421);
and U9403 (N_9403,N_4618,N_4906);
and U9404 (N_9404,N_544,N_5207);
nor U9405 (N_9405,N_1928,N_4664);
xor U9406 (N_9406,N_1753,N_2220);
nor U9407 (N_9407,N_487,N_5824);
nor U9408 (N_9408,N_2286,N_647);
nand U9409 (N_9409,N_1583,N_2373);
and U9410 (N_9410,N_4028,N_155);
nor U9411 (N_9411,N_3943,N_4271);
xnor U9412 (N_9412,N_3360,N_4145);
and U9413 (N_9413,N_3712,N_4765);
nor U9414 (N_9414,N_1612,N_5214);
xnor U9415 (N_9415,N_5978,N_1915);
nor U9416 (N_9416,N_1247,N_3217);
or U9417 (N_9417,N_3158,N_2180);
and U9418 (N_9418,N_3155,N_625);
or U9419 (N_9419,N_858,N_2192);
nor U9420 (N_9420,N_2737,N_4356);
and U9421 (N_9421,N_5089,N_2007);
nor U9422 (N_9422,N_1031,N_4713);
and U9423 (N_9423,N_1729,N_3223);
nand U9424 (N_9424,N_574,N_2830);
and U9425 (N_9425,N_2028,N_4112);
and U9426 (N_9426,N_2566,N_2873);
nor U9427 (N_9427,N_192,N_2855);
and U9428 (N_9428,N_2070,N_197);
xnor U9429 (N_9429,N_5208,N_3542);
nand U9430 (N_9430,N_3042,N_451);
and U9431 (N_9431,N_614,N_3636);
and U9432 (N_9432,N_3565,N_2584);
nand U9433 (N_9433,N_5485,N_663);
xnor U9434 (N_9434,N_2945,N_3348);
xnor U9435 (N_9435,N_5466,N_5978);
xor U9436 (N_9436,N_4332,N_3648);
nor U9437 (N_9437,N_1702,N_5972);
xor U9438 (N_9438,N_362,N_5403);
xnor U9439 (N_9439,N_791,N_413);
or U9440 (N_9440,N_522,N_3703);
and U9441 (N_9441,N_3322,N_4364);
xor U9442 (N_9442,N_42,N_4663);
and U9443 (N_9443,N_3216,N_2391);
nor U9444 (N_9444,N_3876,N_3804);
xnor U9445 (N_9445,N_4519,N_5219);
or U9446 (N_9446,N_1538,N_318);
nor U9447 (N_9447,N_1454,N_5829);
and U9448 (N_9448,N_1738,N_3536);
xor U9449 (N_9449,N_2268,N_2972);
or U9450 (N_9450,N_5491,N_140);
nand U9451 (N_9451,N_3287,N_154);
nand U9452 (N_9452,N_1118,N_983);
xor U9453 (N_9453,N_5677,N_2892);
or U9454 (N_9454,N_4854,N_302);
or U9455 (N_9455,N_3292,N_2204);
nand U9456 (N_9456,N_2363,N_2380);
xor U9457 (N_9457,N_3110,N_1686);
nand U9458 (N_9458,N_2207,N_2726);
nor U9459 (N_9459,N_1494,N_5817);
xor U9460 (N_9460,N_1692,N_5011);
or U9461 (N_9461,N_3812,N_1541);
and U9462 (N_9462,N_5760,N_436);
or U9463 (N_9463,N_4327,N_5041);
xnor U9464 (N_9464,N_5428,N_3212);
xor U9465 (N_9465,N_639,N_3969);
or U9466 (N_9466,N_1071,N_3675);
or U9467 (N_9467,N_255,N_5923);
nor U9468 (N_9468,N_847,N_300);
xor U9469 (N_9469,N_4961,N_637);
or U9470 (N_9470,N_1453,N_4581);
or U9471 (N_9471,N_213,N_190);
nor U9472 (N_9472,N_4021,N_1119);
and U9473 (N_9473,N_3123,N_2667);
and U9474 (N_9474,N_918,N_962);
or U9475 (N_9475,N_3522,N_2952);
xor U9476 (N_9476,N_1213,N_4208);
or U9477 (N_9477,N_563,N_2042);
nand U9478 (N_9478,N_321,N_1221);
nand U9479 (N_9479,N_5153,N_2225);
nor U9480 (N_9480,N_3547,N_3615);
nand U9481 (N_9481,N_5543,N_4100);
nand U9482 (N_9482,N_2342,N_2396);
nand U9483 (N_9483,N_327,N_4029);
xor U9484 (N_9484,N_3940,N_3920);
nand U9485 (N_9485,N_4567,N_5252);
xor U9486 (N_9486,N_4260,N_3172);
or U9487 (N_9487,N_5109,N_2887);
nand U9488 (N_9488,N_1977,N_3849);
and U9489 (N_9489,N_5815,N_5700);
or U9490 (N_9490,N_428,N_4147);
nor U9491 (N_9491,N_5426,N_1357);
or U9492 (N_9492,N_3067,N_4358);
or U9493 (N_9493,N_957,N_5038);
nor U9494 (N_9494,N_2500,N_5513);
xor U9495 (N_9495,N_4486,N_4589);
xor U9496 (N_9496,N_4914,N_2797);
nand U9497 (N_9497,N_1508,N_500);
xor U9498 (N_9498,N_4214,N_1461);
and U9499 (N_9499,N_3305,N_3945);
nor U9500 (N_9500,N_3130,N_2843);
nand U9501 (N_9501,N_5531,N_4297);
nor U9502 (N_9502,N_767,N_1592);
or U9503 (N_9503,N_2082,N_2617);
nand U9504 (N_9504,N_525,N_5349);
and U9505 (N_9505,N_5775,N_5081);
and U9506 (N_9506,N_4349,N_1393);
xnor U9507 (N_9507,N_716,N_5775);
and U9508 (N_9508,N_4919,N_3403);
nand U9509 (N_9509,N_3207,N_2848);
nor U9510 (N_9510,N_3080,N_5017);
or U9511 (N_9511,N_167,N_287);
and U9512 (N_9512,N_3546,N_4985);
and U9513 (N_9513,N_4251,N_5831);
nand U9514 (N_9514,N_54,N_4628);
nand U9515 (N_9515,N_3329,N_814);
xor U9516 (N_9516,N_2395,N_4102);
or U9517 (N_9517,N_5105,N_800);
and U9518 (N_9518,N_5798,N_4144);
nand U9519 (N_9519,N_5079,N_2457);
nor U9520 (N_9520,N_1892,N_4977);
xnor U9521 (N_9521,N_4070,N_2718);
or U9522 (N_9522,N_3762,N_1682);
xor U9523 (N_9523,N_1341,N_3231);
xor U9524 (N_9524,N_5962,N_5722);
nor U9525 (N_9525,N_5047,N_4941);
nor U9526 (N_9526,N_1992,N_3704);
and U9527 (N_9527,N_1652,N_2254);
or U9528 (N_9528,N_4614,N_5715);
nand U9529 (N_9529,N_3397,N_964);
or U9530 (N_9530,N_1629,N_1496);
or U9531 (N_9531,N_1478,N_5418);
and U9532 (N_9532,N_1319,N_1493);
and U9533 (N_9533,N_2286,N_4195);
or U9534 (N_9534,N_5854,N_4361);
and U9535 (N_9535,N_4180,N_5807);
nor U9536 (N_9536,N_4085,N_188);
nand U9537 (N_9537,N_1310,N_135);
or U9538 (N_9538,N_2429,N_2043);
and U9539 (N_9539,N_1580,N_3254);
and U9540 (N_9540,N_141,N_3777);
nand U9541 (N_9541,N_1278,N_418);
and U9542 (N_9542,N_3118,N_5871);
or U9543 (N_9543,N_773,N_3515);
nor U9544 (N_9544,N_4875,N_839);
nand U9545 (N_9545,N_2238,N_2178);
nor U9546 (N_9546,N_1433,N_472);
xnor U9547 (N_9547,N_1437,N_4842);
and U9548 (N_9548,N_1653,N_2244);
nand U9549 (N_9549,N_594,N_4172);
and U9550 (N_9550,N_5743,N_5887);
nand U9551 (N_9551,N_5034,N_1522);
nand U9552 (N_9552,N_3268,N_2055);
nand U9553 (N_9553,N_3496,N_5279);
nor U9554 (N_9554,N_1960,N_3085);
and U9555 (N_9555,N_521,N_1918);
or U9556 (N_9556,N_3295,N_592);
xor U9557 (N_9557,N_3289,N_5645);
or U9558 (N_9558,N_3526,N_1008);
and U9559 (N_9559,N_5989,N_2661);
xor U9560 (N_9560,N_1196,N_4155);
nand U9561 (N_9561,N_3847,N_2325);
nor U9562 (N_9562,N_3049,N_5744);
nand U9563 (N_9563,N_363,N_927);
xnor U9564 (N_9564,N_1785,N_4322);
or U9565 (N_9565,N_4515,N_2510);
and U9566 (N_9566,N_3614,N_4888);
and U9567 (N_9567,N_1277,N_3327);
or U9568 (N_9568,N_4072,N_5937);
xnor U9569 (N_9569,N_5968,N_1213);
nor U9570 (N_9570,N_2602,N_4151);
or U9571 (N_9571,N_3131,N_1195);
xor U9572 (N_9572,N_562,N_3769);
or U9573 (N_9573,N_3938,N_1788);
xor U9574 (N_9574,N_3239,N_606);
nand U9575 (N_9575,N_1076,N_836);
or U9576 (N_9576,N_1663,N_847);
and U9577 (N_9577,N_289,N_4245);
xor U9578 (N_9578,N_275,N_5552);
nand U9579 (N_9579,N_4364,N_4372);
nor U9580 (N_9580,N_2987,N_2395);
xor U9581 (N_9581,N_655,N_3421);
nor U9582 (N_9582,N_306,N_850);
xor U9583 (N_9583,N_4220,N_4266);
and U9584 (N_9584,N_790,N_3862);
nor U9585 (N_9585,N_5549,N_2862);
nand U9586 (N_9586,N_2263,N_2209);
xor U9587 (N_9587,N_944,N_1376);
xnor U9588 (N_9588,N_2835,N_5756);
nand U9589 (N_9589,N_1643,N_514);
nor U9590 (N_9590,N_4603,N_2972);
or U9591 (N_9591,N_178,N_506);
xor U9592 (N_9592,N_4900,N_815);
or U9593 (N_9593,N_1450,N_5132);
and U9594 (N_9594,N_3225,N_5405);
xnor U9595 (N_9595,N_923,N_2816);
xor U9596 (N_9596,N_4753,N_2842);
nand U9597 (N_9597,N_628,N_603);
or U9598 (N_9598,N_1732,N_2491);
xor U9599 (N_9599,N_959,N_134);
or U9600 (N_9600,N_657,N_5473);
and U9601 (N_9601,N_4720,N_3761);
xor U9602 (N_9602,N_2449,N_2643);
nor U9603 (N_9603,N_5793,N_3146);
nand U9604 (N_9604,N_4451,N_1266);
nor U9605 (N_9605,N_23,N_5540);
xnor U9606 (N_9606,N_1516,N_329);
xnor U9607 (N_9607,N_5821,N_1257);
nor U9608 (N_9608,N_2166,N_1226);
nand U9609 (N_9609,N_1150,N_5127);
nand U9610 (N_9610,N_306,N_437);
nor U9611 (N_9611,N_5804,N_3935);
nand U9612 (N_9612,N_4017,N_5718);
or U9613 (N_9613,N_251,N_3783);
and U9614 (N_9614,N_5949,N_5427);
nor U9615 (N_9615,N_4927,N_1418);
nor U9616 (N_9616,N_4539,N_1120);
nand U9617 (N_9617,N_534,N_2397);
xnor U9618 (N_9618,N_5574,N_2034);
or U9619 (N_9619,N_4119,N_5361);
xor U9620 (N_9620,N_1213,N_5778);
nand U9621 (N_9621,N_3505,N_5152);
nor U9622 (N_9622,N_4579,N_4356);
nor U9623 (N_9623,N_1554,N_3267);
or U9624 (N_9624,N_4070,N_2681);
xor U9625 (N_9625,N_1185,N_5522);
and U9626 (N_9626,N_851,N_4137);
and U9627 (N_9627,N_947,N_3193);
nand U9628 (N_9628,N_2024,N_2516);
nor U9629 (N_9629,N_3772,N_5189);
nand U9630 (N_9630,N_840,N_2618);
nor U9631 (N_9631,N_14,N_1538);
and U9632 (N_9632,N_3697,N_4260);
xnor U9633 (N_9633,N_2973,N_3851);
nor U9634 (N_9634,N_1251,N_4750);
and U9635 (N_9635,N_2872,N_2460);
nor U9636 (N_9636,N_1578,N_586);
xor U9637 (N_9637,N_2550,N_4756);
xnor U9638 (N_9638,N_5440,N_5530);
or U9639 (N_9639,N_4116,N_3346);
xor U9640 (N_9640,N_5219,N_2544);
or U9641 (N_9641,N_3100,N_5404);
or U9642 (N_9642,N_3354,N_992);
or U9643 (N_9643,N_5907,N_3551);
or U9644 (N_9644,N_107,N_2158);
nand U9645 (N_9645,N_2189,N_1896);
nor U9646 (N_9646,N_904,N_1378);
xnor U9647 (N_9647,N_2502,N_199);
nand U9648 (N_9648,N_5734,N_4704);
and U9649 (N_9649,N_249,N_2721);
nand U9650 (N_9650,N_759,N_2923);
nand U9651 (N_9651,N_1994,N_4246);
nor U9652 (N_9652,N_4801,N_1497);
and U9653 (N_9653,N_1823,N_5022);
nand U9654 (N_9654,N_3151,N_870);
or U9655 (N_9655,N_554,N_4689);
nand U9656 (N_9656,N_3377,N_396);
and U9657 (N_9657,N_283,N_5750);
xor U9658 (N_9658,N_3176,N_4211);
nor U9659 (N_9659,N_2947,N_5826);
nand U9660 (N_9660,N_3824,N_361);
and U9661 (N_9661,N_4021,N_4566);
nor U9662 (N_9662,N_3137,N_5092);
or U9663 (N_9663,N_1890,N_3585);
or U9664 (N_9664,N_2423,N_2570);
or U9665 (N_9665,N_301,N_1402);
nand U9666 (N_9666,N_2013,N_1881);
or U9667 (N_9667,N_1950,N_1916);
xor U9668 (N_9668,N_2284,N_325);
nand U9669 (N_9669,N_1281,N_541);
nor U9670 (N_9670,N_3725,N_1499);
or U9671 (N_9671,N_364,N_5760);
or U9672 (N_9672,N_733,N_4717);
nand U9673 (N_9673,N_4784,N_4940);
nor U9674 (N_9674,N_2335,N_4422);
nor U9675 (N_9675,N_321,N_4776);
nand U9676 (N_9676,N_2460,N_7);
nand U9677 (N_9677,N_3798,N_4685);
nor U9678 (N_9678,N_2643,N_2193);
and U9679 (N_9679,N_4053,N_2512);
and U9680 (N_9680,N_1176,N_3949);
and U9681 (N_9681,N_700,N_5126);
nand U9682 (N_9682,N_3797,N_972);
xnor U9683 (N_9683,N_5239,N_2321);
or U9684 (N_9684,N_4478,N_4485);
nor U9685 (N_9685,N_5785,N_422);
and U9686 (N_9686,N_4875,N_2807);
and U9687 (N_9687,N_2810,N_2323);
nand U9688 (N_9688,N_4371,N_1180);
nor U9689 (N_9689,N_4905,N_5551);
xor U9690 (N_9690,N_5928,N_3954);
nor U9691 (N_9691,N_955,N_628);
xnor U9692 (N_9692,N_4546,N_5931);
nor U9693 (N_9693,N_2139,N_3429);
and U9694 (N_9694,N_4598,N_3644);
nor U9695 (N_9695,N_284,N_3700);
and U9696 (N_9696,N_4301,N_5185);
nor U9697 (N_9697,N_3975,N_3633);
and U9698 (N_9698,N_2210,N_247);
nor U9699 (N_9699,N_5072,N_5310);
nor U9700 (N_9700,N_2068,N_1694);
or U9701 (N_9701,N_1397,N_2361);
nand U9702 (N_9702,N_69,N_447);
and U9703 (N_9703,N_3410,N_2852);
xnor U9704 (N_9704,N_5076,N_5074);
nor U9705 (N_9705,N_4679,N_2670);
nand U9706 (N_9706,N_3232,N_3440);
or U9707 (N_9707,N_2367,N_1116);
xnor U9708 (N_9708,N_4457,N_1804);
or U9709 (N_9709,N_3604,N_123);
or U9710 (N_9710,N_3216,N_3524);
xor U9711 (N_9711,N_1105,N_3466);
nand U9712 (N_9712,N_3,N_2942);
nand U9713 (N_9713,N_4595,N_942);
xnor U9714 (N_9714,N_401,N_1046);
nand U9715 (N_9715,N_4825,N_4506);
and U9716 (N_9716,N_5253,N_4169);
or U9717 (N_9717,N_5504,N_4894);
or U9718 (N_9718,N_5548,N_5039);
and U9719 (N_9719,N_1118,N_3265);
nand U9720 (N_9720,N_2304,N_3917);
xnor U9721 (N_9721,N_2927,N_4508);
xnor U9722 (N_9722,N_1551,N_3574);
nand U9723 (N_9723,N_4036,N_414);
and U9724 (N_9724,N_606,N_318);
or U9725 (N_9725,N_4559,N_1151);
and U9726 (N_9726,N_671,N_3348);
xor U9727 (N_9727,N_2713,N_4026);
xnor U9728 (N_9728,N_5385,N_922);
nor U9729 (N_9729,N_3953,N_2627);
and U9730 (N_9730,N_5299,N_2036);
xnor U9731 (N_9731,N_2693,N_4258);
nand U9732 (N_9732,N_2296,N_5520);
and U9733 (N_9733,N_1754,N_5572);
or U9734 (N_9734,N_3434,N_2774);
and U9735 (N_9735,N_4928,N_108);
nor U9736 (N_9736,N_579,N_1286);
and U9737 (N_9737,N_5466,N_2616);
or U9738 (N_9738,N_3169,N_5006);
nor U9739 (N_9739,N_3766,N_237);
nor U9740 (N_9740,N_4515,N_1814);
or U9741 (N_9741,N_99,N_4570);
or U9742 (N_9742,N_2295,N_5853);
and U9743 (N_9743,N_4657,N_4605);
xor U9744 (N_9744,N_5494,N_2949);
and U9745 (N_9745,N_1656,N_1577);
nor U9746 (N_9746,N_3852,N_2026);
nand U9747 (N_9747,N_2471,N_1825);
nor U9748 (N_9748,N_255,N_3999);
nand U9749 (N_9749,N_5396,N_1058);
nor U9750 (N_9750,N_2338,N_5383);
nor U9751 (N_9751,N_1528,N_268);
or U9752 (N_9752,N_4262,N_512);
and U9753 (N_9753,N_2371,N_1508);
and U9754 (N_9754,N_774,N_3342);
nor U9755 (N_9755,N_3195,N_273);
xnor U9756 (N_9756,N_5447,N_5641);
nor U9757 (N_9757,N_4724,N_4577);
nand U9758 (N_9758,N_1693,N_2300);
nand U9759 (N_9759,N_2933,N_134);
nor U9760 (N_9760,N_39,N_5150);
and U9761 (N_9761,N_5870,N_2313);
and U9762 (N_9762,N_5722,N_5683);
nor U9763 (N_9763,N_3267,N_385);
nor U9764 (N_9764,N_3563,N_1434);
or U9765 (N_9765,N_5998,N_1659);
xnor U9766 (N_9766,N_3810,N_1492);
nand U9767 (N_9767,N_2126,N_2111);
or U9768 (N_9768,N_5708,N_2450);
or U9769 (N_9769,N_4030,N_3886);
nor U9770 (N_9770,N_1799,N_5695);
or U9771 (N_9771,N_3213,N_3977);
nor U9772 (N_9772,N_4353,N_4894);
nor U9773 (N_9773,N_402,N_3772);
and U9774 (N_9774,N_1710,N_442);
and U9775 (N_9775,N_3999,N_3616);
nand U9776 (N_9776,N_1843,N_4961);
nand U9777 (N_9777,N_2150,N_4456);
xnor U9778 (N_9778,N_4854,N_230);
xor U9779 (N_9779,N_5747,N_2523);
or U9780 (N_9780,N_3894,N_1226);
and U9781 (N_9781,N_5707,N_3030);
and U9782 (N_9782,N_4079,N_5873);
xnor U9783 (N_9783,N_2871,N_2038);
and U9784 (N_9784,N_3849,N_3561);
nor U9785 (N_9785,N_166,N_3484);
nand U9786 (N_9786,N_1110,N_3361);
nand U9787 (N_9787,N_2623,N_1044);
nor U9788 (N_9788,N_2366,N_2239);
xor U9789 (N_9789,N_5462,N_4050);
or U9790 (N_9790,N_3662,N_3255);
nand U9791 (N_9791,N_1754,N_5075);
xor U9792 (N_9792,N_3516,N_2711);
or U9793 (N_9793,N_1352,N_2646);
and U9794 (N_9794,N_3161,N_3843);
or U9795 (N_9795,N_1002,N_3685);
and U9796 (N_9796,N_501,N_4380);
nand U9797 (N_9797,N_5967,N_2496);
nor U9798 (N_9798,N_3004,N_1208);
xnor U9799 (N_9799,N_1188,N_5424);
or U9800 (N_9800,N_1214,N_3470);
xnor U9801 (N_9801,N_465,N_1819);
or U9802 (N_9802,N_1904,N_2079);
nand U9803 (N_9803,N_4765,N_1082);
xor U9804 (N_9804,N_4847,N_4065);
and U9805 (N_9805,N_1487,N_353);
nor U9806 (N_9806,N_5050,N_2675);
or U9807 (N_9807,N_1444,N_4291);
and U9808 (N_9808,N_4116,N_5410);
xor U9809 (N_9809,N_3854,N_2433);
nor U9810 (N_9810,N_3312,N_2874);
nand U9811 (N_9811,N_765,N_1387);
nor U9812 (N_9812,N_1863,N_3443);
and U9813 (N_9813,N_3511,N_5647);
nand U9814 (N_9814,N_5739,N_3356);
nand U9815 (N_9815,N_1258,N_5363);
or U9816 (N_9816,N_4668,N_1734);
xor U9817 (N_9817,N_3123,N_5859);
and U9818 (N_9818,N_2100,N_759);
xor U9819 (N_9819,N_116,N_1714);
nor U9820 (N_9820,N_4438,N_4437);
and U9821 (N_9821,N_1668,N_1413);
and U9822 (N_9822,N_4948,N_4684);
nor U9823 (N_9823,N_655,N_4832);
or U9824 (N_9824,N_4683,N_2880);
and U9825 (N_9825,N_4561,N_2260);
or U9826 (N_9826,N_5554,N_2345);
and U9827 (N_9827,N_2756,N_3098);
nor U9828 (N_9828,N_200,N_3559);
or U9829 (N_9829,N_619,N_1034);
or U9830 (N_9830,N_5692,N_974);
nand U9831 (N_9831,N_1611,N_5624);
or U9832 (N_9832,N_4928,N_5308);
and U9833 (N_9833,N_4377,N_902);
xnor U9834 (N_9834,N_3195,N_5228);
xor U9835 (N_9835,N_1091,N_2864);
or U9836 (N_9836,N_3755,N_4142);
or U9837 (N_9837,N_5144,N_3474);
or U9838 (N_9838,N_2699,N_2713);
nand U9839 (N_9839,N_5503,N_2403);
or U9840 (N_9840,N_3945,N_4934);
or U9841 (N_9841,N_2899,N_1800);
xor U9842 (N_9842,N_458,N_4240);
nor U9843 (N_9843,N_5606,N_4490);
xor U9844 (N_9844,N_643,N_5753);
nor U9845 (N_9845,N_4272,N_5753);
nor U9846 (N_9846,N_1809,N_5944);
nor U9847 (N_9847,N_1440,N_5683);
nor U9848 (N_9848,N_1022,N_4170);
and U9849 (N_9849,N_582,N_5644);
nand U9850 (N_9850,N_5350,N_1568);
xor U9851 (N_9851,N_2600,N_1536);
nand U9852 (N_9852,N_4635,N_5079);
and U9853 (N_9853,N_3022,N_3203);
nor U9854 (N_9854,N_5666,N_773);
xnor U9855 (N_9855,N_4990,N_174);
nor U9856 (N_9856,N_2454,N_1610);
and U9857 (N_9857,N_2532,N_5176);
or U9858 (N_9858,N_4856,N_1806);
nor U9859 (N_9859,N_4580,N_2431);
nor U9860 (N_9860,N_3388,N_3576);
xor U9861 (N_9861,N_245,N_2588);
and U9862 (N_9862,N_2664,N_747);
or U9863 (N_9863,N_177,N_52);
and U9864 (N_9864,N_4613,N_2516);
nor U9865 (N_9865,N_2380,N_3728);
or U9866 (N_9866,N_4483,N_5091);
nand U9867 (N_9867,N_1964,N_5972);
nand U9868 (N_9868,N_814,N_284);
nand U9869 (N_9869,N_847,N_2671);
nand U9870 (N_9870,N_945,N_4425);
or U9871 (N_9871,N_1307,N_408);
and U9872 (N_9872,N_328,N_3291);
nor U9873 (N_9873,N_1527,N_2566);
or U9874 (N_9874,N_165,N_112);
and U9875 (N_9875,N_5643,N_689);
and U9876 (N_9876,N_3393,N_4348);
nand U9877 (N_9877,N_2390,N_591);
or U9878 (N_9878,N_2923,N_4822);
xor U9879 (N_9879,N_3236,N_2938);
or U9880 (N_9880,N_2471,N_3456);
nand U9881 (N_9881,N_1935,N_3926);
and U9882 (N_9882,N_2107,N_5637);
nand U9883 (N_9883,N_4059,N_1941);
nand U9884 (N_9884,N_5849,N_364);
and U9885 (N_9885,N_3732,N_61);
nor U9886 (N_9886,N_4245,N_3659);
or U9887 (N_9887,N_1301,N_1744);
nor U9888 (N_9888,N_3676,N_5118);
nand U9889 (N_9889,N_386,N_1035);
nand U9890 (N_9890,N_575,N_5265);
or U9891 (N_9891,N_4451,N_5423);
or U9892 (N_9892,N_3304,N_4973);
nand U9893 (N_9893,N_787,N_978);
nor U9894 (N_9894,N_2160,N_5372);
nor U9895 (N_9895,N_2793,N_4059);
xnor U9896 (N_9896,N_4366,N_3932);
or U9897 (N_9897,N_2563,N_3763);
nor U9898 (N_9898,N_4654,N_4813);
and U9899 (N_9899,N_616,N_2529);
or U9900 (N_9900,N_2400,N_3354);
and U9901 (N_9901,N_2470,N_1055);
and U9902 (N_9902,N_5049,N_5613);
nand U9903 (N_9903,N_5202,N_2003);
and U9904 (N_9904,N_2746,N_3156);
or U9905 (N_9905,N_4916,N_5377);
xnor U9906 (N_9906,N_4905,N_1808);
or U9907 (N_9907,N_695,N_1277);
xor U9908 (N_9908,N_4748,N_4142);
nor U9909 (N_9909,N_4894,N_4048);
nand U9910 (N_9910,N_1027,N_3413);
or U9911 (N_9911,N_3543,N_1947);
xnor U9912 (N_9912,N_280,N_2139);
or U9913 (N_9913,N_3707,N_711);
or U9914 (N_9914,N_628,N_5634);
and U9915 (N_9915,N_2000,N_4213);
xor U9916 (N_9916,N_5584,N_4953);
nand U9917 (N_9917,N_1683,N_2950);
nor U9918 (N_9918,N_5777,N_842);
and U9919 (N_9919,N_1404,N_5461);
nand U9920 (N_9920,N_971,N_3412);
xnor U9921 (N_9921,N_3485,N_3700);
xnor U9922 (N_9922,N_1151,N_3603);
nand U9923 (N_9923,N_3029,N_5688);
and U9924 (N_9924,N_4731,N_1562);
nor U9925 (N_9925,N_2072,N_754);
xor U9926 (N_9926,N_5425,N_1654);
and U9927 (N_9927,N_2504,N_125);
and U9928 (N_9928,N_2874,N_3687);
nand U9929 (N_9929,N_5900,N_2410);
nand U9930 (N_9930,N_1939,N_2582);
nor U9931 (N_9931,N_4943,N_4652);
or U9932 (N_9932,N_2336,N_4528);
xnor U9933 (N_9933,N_5953,N_2126);
or U9934 (N_9934,N_3775,N_2329);
xnor U9935 (N_9935,N_1321,N_1078);
xnor U9936 (N_9936,N_2271,N_2071);
or U9937 (N_9937,N_5612,N_4438);
or U9938 (N_9938,N_4053,N_3315);
nand U9939 (N_9939,N_1169,N_3586);
nor U9940 (N_9940,N_1269,N_1600);
nand U9941 (N_9941,N_4428,N_2436);
or U9942 (N_9942,N_5411,N_1485);
xnor U9943 (N_9943,N_160,N_701);
xor U9944 (N_9944,N_3928,N_2252);
nor U9945 (N_9945,N_5482,N_2183);
nand U9946 (N_9946,N_4013,N_2373);
xnor U9947 (N_9947,N_5233,N_3725);
xnor U9948 (N_9948,N_5236,N_679);
or U9949 (N_9949,N_3180,N_716);
xor U9950 (N_9950,N_227,N_2854);
xnor U9951 (N_9951,N_3763,N_4088);
and U9952 (N_9952,N_3770,N_1181);
nand U9953 (N_9953,N_4954,N_4038);
and U9954 (N_9954,N_2302,N_4671);
and U9955 (N_9955,N_4889,N_4530);
xnor U9956 (N_9956,N_1730,N_3257);
or U9957 (N_9957,N_2853,N_3172);
nand U9958 (N_9958,N_5237,N_4045);
nand U9959 (N_9959,N_1271,N_2874);
and U9960 (N_9960,N_299,N_4937);
and U9961 (N_9961,N_5835,N_399);
xor U9962 (N_9962,N_4585,N_3474);
and U9963 (N_9963,N_986,N_1872);
xnor U9964 (N_9964,N_4628,N_5506);
nor U9965 (N_9965,N_55,N_5634);
nor U9966 (N_9966,N_3494,N_1918);
nor U9967 (N_9967,N_2660,N_5260);
nand U9968 (N_9968,N_3868,N_5292);
and U9969 (N_9969,N_4390,N_5382);
nor U9970 (N_9970,N_5234,N_4286);
nand U9971 (N_9971,N_4081,N_5330);
nand U9972 (N_9972,N_687,N_234);
xor U9973 (N_9973,N_5175,N_3898);
nor U9974 (N_9974,N_694,N_4375);
xor U9975 (N_9975,N_3132,N_3704);
or U9976 (N_9976,N_77,N_3377);
or U9977 (N_9977,N_1154,N_503);
xnor U9978 (N_9978,N_2499,N_2635);
and U9979 (N_9979,N_4803,N_152);
xor U9980 (N_9980,N_243,N_603);
nor U9981 (N_9981,N_2922,N_1886);
and U9982 (N_9982,N_4221,N_2888);
nor U9983 (N_9983,N_2376,N_118);
nor U9984 (N_9984,N_484,N_2016);
and U9985 (N_9985,N_1671,N_3827);
xnor U9986 (N_9986,N_3739,N_2780);
and U9987 (N_9987,N_1864,N_3106);
and U9988 (N_9988,N_1757,N_701);
and U9989 (N_9989,N_411,N_3470);
and U9990 (N_9990,N_1072,N_423);
or U9991 (N_9991,N_4998,N_3549);
nand U9992 (N_9992,N_325,N_5809);
xnor U9993 (N_9993,N_664,N_4070);
nand U9994 (N_9994,N_3114,N_668);
nor U9995 (N_9995,N_1747,N_5432);
and U9996 (N_9996,N_4312,N_415);
xor U9997 (N_9997,N_1061,N_818);
or U9998 (N_9998,N_5530,N_4764);
or U9999 (N_9999,N_5207,N_874);
or U10000 (N_10000,N_2408,N_3829);
and U10001 (N_10001,N_96,N_2107);
xor U10002 (N_10002,N_4178,N_3152);
and U10003 (N_10003,N_1276,N_1429);
or U10004 (N_10004,N_1793,N_413);
xor U10005 (N_10005,N_3408,N_4933);
and U10006 (N_10006,N_4985,N_3540);
or U10007 (N_10007,N_1137,N_1944);
and U10008 (N_10008,N_4926,N_751);
nand U10009 (N_10009,N_4376,N_3488);
xnor U10010 (N_10010,N_1411,N_4677);
xnor U10011 (N_10011,N_5021,N_1342);
nand U10012 (N_10012,N_1036,N_3297);
xor U10013 (N_10013,N_318,N_1224);
xor U10014 (N_10014,N_4755,N_1980);
and U10015 (N_10015,N_5739,N_813);
or U10016 (N_10016,N_5189,N_298);
nand U10017 (N_10017,N_257,N_1608);
or U10018 (N_10018,N_3334,N_4516);
and U10019 (N_10019,N_388,N_1151);
xor U10020 (N_10020,N_2218,N_4090);
nor U10021 (N_10021,N_3502,N_5040);
or U10022 (N_10022,N_5895,N_5079);
or U10023 (N_10023,N_1216,N_519);
or U10024 (N_10024,N_5948,N_890);
xnor U10025 (N_10025,N_5727,N_5615);
or U10026 (N_10026,N_748,N_865);
xor U10027 (N_10027,N_1057,N_4766);
xnor U10028 (N_10028,N_628,N_3425);
and U10029 (N_10029,N_3948,N_3801);
xnor U10030 (N_10030,N_229,N_1579);
xor U10031 (N_10031,N_3578,N_3700);
nand U10032 (N_10032,N_1698,N_963);
nor U10033 (N_10033,N_1642,N_2532);
or U10034 (N_10034,N_3084,N_3765);
xor U10035 (N_10035,N_4502,N_1057);
or U10036 (N_10036,N_4463,N_3152);
nand U10037 (N_10037,N_1804,N_678);
and U10038 (N_10038,N_4738,N_3210);
nand U10039 (N_10039,N_5850,N_2128);
and U10040 (N_10040,N_3364,N_3558);
nor U10041 (N_10041,N_1184,N_4149);
and U10042 (N_10042,N_280,N_3296);
xnor U10043 (N_10043,N_3399,N_5148);
and U10044 (N_10044,N_2504,N_1068);
xor U10045 (N_10045,N_3770,N_3107);
and U10046 (N_10046,N_4739,N_2825);
nand U10047 (N_10047,N_3537,N_4982);
nor U10048 (N_10048,N_3739,N_838);
and U10049 (N_10049,N_897,N_5409);
xor U10050 (N_10050,N_4451,N_1171);
and U10051 (N_10051,N_2218,N_5668);
xor U10052 (N_10052,N_2719,N_3876);
xnor U10053 (N_10053,N_490,N_5456);
nand U10054 (N_10054,N_1327,N_4306);
xor U10055 (N_10055,N_4331,N_4144);
nor U10056 (N_10056,N_5076,N_3724);
or U10057 (N_10057,N_252,N_1193);
nand U10058 (N_10058,N_4923,N_2609);
and U10059 (N_10059,N_2790,N_5523);
or U10060 (N_10060,N_4244,N_1047);
nor U10061 (N_10061,N_1683,N_3512);
or U10062 (N_10062,N_2765,N_4469);
and U10063 (N_10063,N_1857,N_4742);
or U10064 (N_10064,N_3831,N_4075);
or U10065 (N_10065,N_4402,N_585);
nor U10066 (N_10066,N_1564,N_2907);
or U10067 (N_10067,N_1972,N_3971);
xnor U10068 (N_10068,N_5454,N_5274);
nor U10069 (N_10069,N_5730,N_1667);
nor U10070 (N_10070,N_2404,N_2049);
and U10071 (N_10071,N_3314,N_2946);
or U10072 (N_10072,N_973,N_3946);
xor U10073 (N_10073,N_4210,N_3959);
and U10074 (N_10074,N_5883,N_5277);
nor U10075 (N_10075,N_1006,N_826);
and U10076 (N_10076,N_1395,N_1837);
nand U10077 (N_10077,N_5891,N_3361);
or U10078 (N_10078,N_3990,N_1061);
or U10079 (N_10079,N_1603,N_3301);
nand U10080 (N_10080,N_4815,N_5499);
nor U10081 (N_10081,N_2599,N_3564);
or U10082 (N_10082,N_5008,N_1665);
or U10083 (N_10083,N_1525,N_2215);
xor U10084 (N_10084,N_1541,N_165);
and U10085 (N_10085,N_2840,N_3301);
xor U10086 (N_10086,N_4241,N_1291);
nor U10087 (N_10087,N_2252,N_1414);
and U10088 (N_10088,N_2728,N_2614);
xor U10089 (N_10089,N_5516,N_743);
or U10090 (N_10090,N_128,N_873);
nand U10091 (N_10091,N_1838,N_3903);
or U10092 (N_10092,N_3711,N_724);
nand U10093 (N_10093,N_2460,N_186);
nand U10094 (N_10094,N_1272,N_2154);
xor U10095 (N_10095,N_173,N_493);
and U10096 (N_10096,N_710,N_1493);
xor U10097 (N_10097,N_3695,N_1617);
and U10098 (N_10098,N_5614,N_4039);
xor U10099 (N_10099,N_2922,N_3065);
or U10100 (N_10100,N_3808,N_5521);
xnor U10101 (N_10101,N_2522,N_2704);
nor U10102 (N_10102,N_1909,N_5943);
or U10103 (N_10103,N_1675,N_520);
or U10104 (N_10104,N_1109,N_2767);
nand U10105 (N_10105,N_404,N_5446);
nor U10106 (N_10106,N_4870,N_3385);
or U10107 (N_10107,N_1197,N_4455);
and U10108 (N_10108,N_1728,N_2990);
xor U10109 (N_10109,N_2545,N_1005);
nor U10110 (N_10110,N_411,N_3713);
or U10111 (N_10111,N_2697,N_208);
nor U10112 (N_10112,N_3060,N_1945);
or U10113 (N_10113,N_1744,N_4504);
nor U10114 (N_10114,N_2672,N_4508);
and U10115 (N_10115,N_1283,N_2385);
and U10116 (N_10116,N_3401,N_2051);
nand U10117 (N_10117,N_5647,N_1331);
nand U10118 (N_10118,N_343,N_5220);
nand U10119 (N_10119,N_5969,N_1381);
nor U10120 (N_10120,N_3015,N_1161);
or U10121 (N_10121,N_3472,N_5428);
nor U10122 (N_10122,N_4337,N_3383);
and U10123 (N_10123,N_1680,N_2693);
xor U10124 (N_10124,N_4187,N_5948);
nand U10125 (N_10125,N_387,N_5932);
or U10126 (N_10126,N_1676,N_5452);
and U10127 (N_10127,N_1403,N_4546);
xor U10128 (N_10128,N_4051,N_4744);
or U10129 (N_10129,N_5675,N_5930);
nor U10130 (N_10130,N_5791,N_1103);
xnor U10131 (N_10131,N_4472,N_990);
nor U10132 (N_10132,N_2134,N_2148);
nand U10133 (N_10133,N_3631,N_2323);
and U10134 (N_10134,N_1132,N_2734);
and U10135 (N_10135,N_2449,N_2378);
nor U10136 (N_10136,N_3752,N_2030);
nand U10137 (N_10137,N_5177,N_3690);
or U10138 (N_10138,N_5994,N_485);
nand U10139 (N_10139,N_3931,N_5073);
xnor U10140 (N_10140,N_3145,N_1045);
nand U10141 (N_10141,N_708,N_5631);
nand U10142 (N_10142,N_827,N_2065);
or U10143 (N_10143,N_4161,N_4102);
and U10144 (N_10144,N_4754,N_2784);
or U10145 (N_10145,N_1024,N_504);
and U10146 (N_10146,N_5864,N_629);
xnor U10147 (N_10147,N_5556,N_2170);
or U10148 (N_10148,N_854,N_4046);
nor U10149 (N_10149,N_3160,N_3625);
xnor U10150 (N_10150,N_5812,N_3736);
xnor U10151 (N_10151,N_3054,N_2840);
or U10152 (N_10152,N_289,N_5179);
nor U10153 (N_10153,N_4641,N_4108);
and U10154 (N_10154,N_490,N_4404);
nand U10155 (N_10155,N_3778,N_3219);
and U10156 (N_10156,N_242,N_1450);
and U10157 (N_10157,N_1157,N_4990);
xor U10158 (N_10158,N_586,N_4724);
nor U10159 (N_10159,N_1984,N_3105);
nand U10160 (N_10160,N_4367,N_940);
nand U10161 (N_10161,N_4871,N_1137);
and U10162 (N_10162,N_2867,N_5951);
or U10163 (N_10163,N_4192,N_4407);
and U10164 (N_10164,N_2018,N_1185);
nor U10165 (N_10165,N_2527,N_134);
nand U10166 (N_10166,N_4333,N_949);
nand U10167 (N_10167,N_2267,N_4382);
or U10168 (N_10168,N_2122,N_3312);
nand U10169 (N_10169,N_1714,N_820);
nand U10170 (N_10170,N_1882,N_4162);
and U10171 (N_10171,N_1129,N_3547);
and U10172 (N_10172,N_3900,N_4580);
or U10173 (N_10173,N_5217,N_3617);
xnor U10174 (N_10174,N_1679,N_177);
nand U10175 (N_10175,N_1008,N_2404);
nand U10176 (N_10176,N_683,N_5452);
and U10177 (N_10177,N_4495,N_259);
nor U10178 (N_10178,N_3165,N_5323);
or U10179 (N_10179,N_2594,N_2107);
xor U10180 (N_10180,N_3327,N_3713);
nor U10181 (N_10181,N_928,N_3769);
or U10182 (N_10182,N_2239,N_514);
and U10183 (N_10183,N_4844,N_5449);
or U10184 (N_10184,N_2770,N_5526);
and U10185 (N_10185,N_5782,N_4915);
and U10186 (N_10186,N_3441,N_4920);
xnor U10187 (N_10187,N_980,N_1120);
or U10188 (N_10188,N_5009,N_799);
and U10189 (N_10189,N_1103,N_3475);
nand U10190 (N_10190,N_108,N_5243);
xnor U10191 (N_10191,N_3833,N_4095);
xor U10192 (N_10192,N_4442,N_1712);
nor U10193 (N_10193,N_4891,N_146);
nand U10194 (N_10194,N_3347,N_5978);
nor U10195 (N_10195,N_5128,N_222);
nor U10196 (N_10196,N_530,N_5488);
nor U10197 (N_10197,N_214,N_2986);
or U10198 (N_10198,N_2511,N_1273);
or U10199 (N_10199,N_4248,N_2836);
nand U10200 (N_10200,N_5918,N_2789);
nor U10201 (N_10201,N_4752,N_5093);
or U10202 (N_10202,N_4433,N_4294);
nor U10203 (N_10203,N_3057,N_494);
nor U10204 (N_10204,N_2463,N_1185);
nor U10205 (N_10205,N_4466,N_2271);
nor U10206 (N_10206,N_312,N_2375);
nand U10207 (N_10207,N_361,N_4983);
xor U10208 (N_10208,N_3489,N_5241);
and U10209 (N_10209,N_5209,N_1080);
and U10210 (N_10210,N_4289,N_957);
xnor U10211 (N_10211,N_2613,N_2352);
nor U10212 (N_10212,N_2934,N_5628);
and U10213 (N_10213,N_2419,N_4839);
nor U10214 (N_10214,N_1238,N_95);
or U10215 (N_10215,N_3033,N_3594);
xor U10216 (N_10216,N_1692,N_3987);
nor U10217 (N_10217,N_5873,N_3281);
and U10218 (N_10218,N_2961,N_210);
and U10219 (N_10219,N_3556,N_3054);
nor U10220 (N_10220,N_3404,N_3793);
nand U10221 (N_10221,N_1534,N_3145);
nor U10222 (N_10222,N_3452,N_1081);
or U10223 (N_10223,N_1811,N_5362);
nor U10224 (N_10224,N_1527,N_4351);
nand U10225 (N_10225,N_4778,N_3657);
xnor U10226 (N_10226,N_1932,N_1687);
nor U10227 (N_10227,N_3733,N_5218);
or U10228 (N_10228,N_4123,N_5184);
and U10229 (N_10229,N_3979,N_5588);
nor U10230 (N_10230,N_1342,N_2187);
xnor U10231 (N_10231,N_531,N_2332);
xnor U10232 (N_10232,N_320,N_3345);
nand U10233 (N_10233,N_5890,N_2399);
nor U10234 (N_10234,N_4572,N_5067);
nand U10235 (N_10235,N_5807,N_4462);
or U10236 (N_10236,N_4064,N_1946);
nand U10237 (N_10237,N_61,N_978);
xnor U10238 (N_10238,N_1141,N_1578);
xor U10239 (N_10239,N_3724,N_2295);
and U10240 (N_10240,N_1281,N_5267);
xnor U10241 (N_10241,N_2178,N_5130);
and U10242 (N_10242,N_5497,N_2087);
nor U10243 (N_10243,N_2370,N_393);
xnor U10244 (N_10244,N_3047,N_4430);
or U10245 (N_10245,N_4992,N_1457);
and U10246 (N_10246,N_5332,N_3887);
and U10247 (N_10247,N_1716,N_2909);
or U10248 (N_10248,N_4325,N_4778);
and U10249 (N_10249,N_3974,N_5820);
and U10250 (N_10250,N_4359,N_5393);
nand U10251 (N_10251,N_2917,N_2310);
xnor U10252 (N_10252,N_2038,N_1309);
and U10253 (N_10253,N_4241,N_3699);
nor U10254 (N_10254,N_4849,N_2780);
nand U10255 (N_10255,N_5147,N_4618);
xnor U10256 (N_10256,N_1336,N_496);
nor U10257 (N_10257,N_5065,N_3155);
nor U10258 (N_10258,N_866,N_1704);
nor U10259 (N_10259,N_4559,N_543);
xor U10260 (N_10260,N_3635,N_2753);
and U10261 (N_10261,N_5125,N_2735);
nor U10262 (N_10262,N_377,N_486);
nor U10263 (N_10263,N_1289,N_4878);
or U10264 (N_10264,N_5027,N_807);
nand U10265 (N_10265,N_1204,N_4790);
nor U10266 (N_10266,N_1469,N_439);
xor U10267 (N_10267,N_4896,N_4779);
nand U10268 (N_10268,N_4182,N_4410);
xnor U10269 (N_10269,N_1184,N_1355);
nand U10270 (N_10270,N_1329,N_4182);
nor U10271 (N_10271,N_2380,N_533);
or U10272 (N_10272,N_1804,N_1037);
xnor U10273 (N_10273,N_5808,N_4121);
nand U10274 (N_10274,N_4689,N_5372);
xnor U10275 (N_10275,N_2910,N_4901);
or U10276 (N_10276,N_490,N_4854);
and U10277 (N_10277,N_4310,N_1442);
nor U10278 (N_10278,N_5715,N_1744);
or U10279 (N_10279,N_1580,N_5091);
nand U10280 (N_10280,N_2677,N_4128);
or U10281 (N_10281,N_5398,N_5929);
or U10282 (N_10282,N_3034,N_4809);
or U10283 (N_10283,N_5482,N_4063);
or U10284 (N_10284,N_4901,N_3875);
nand U10285 (N_10285,N_268,N_1192);
and U10286 (N_10286,N_5952,N_4824);
and U10287 (N_10287,N_717,N_3195);
and U10288 (N_10288,N_3462,N_1432);
nor U10289 (N_10289,N_4374,N_1347);
nor U10290 (N_10290,N_2625,N_1995);
or U10291 (N_10291,N_806,N_3814);
or U10292 (N_10292,N_2583,N_354);
and U10293 (N_10293,N_714,N_742);
nand U10294 (N_10294,N_3021,N_2468);
xnor U10295 (N_10295,N_4386,N_5812);
nand U10296 (N_10296,N_1241,N_4063);
xnor U10297 (N_10297,N_1472,N_5148);
nand U10298 (N_10298,N_5760,N_1657);
nand U10299 (N_10299,N_5639,N_967);
xnor U10300 (N_10300,N_3703,N_4109);
nor U10301 (N_10301,N_1872,N_1077);
and U10302 (N_10302,N_4702,N_4301);
xnor U10303 (N_10303,N_5096,N_2142);
nor U10304 (N_10304,N_1150,N_4921);
and U10305 (N_10305,N_2755,N_5443);
nor U10306 (N_10306,N_3960,N_5171);
nor U10307 (N_10307,N_1072,N_2209);
or U10308 (N_10308,N_378,N_3624);
and U10309 (N_10309,N_3660,N_2918);
or U10310 (N_10310,N_287,N_1962);
xor U10311 (N_10311,N_5320,N_5858);
xnor U10312 (N_10312,N_2838,N_3826);
and U10313 (N_10313,N_4029,N_1199);
and U10314 (N_10314,N_5526,N_2403);
and U10315 (N_10315,N_4578,N_2732);
nand U10316 (N_10316,N_28,N_5860);
nand U10317 (N_10317,N_1348,N_5695);
and U10318 (N_10318,N_3755,N_1739);
nor U10319 (N_10319,N_4907,N_3545);
and U10320 (N_10320,N_1106,N_377);
and U10321 (N_10321,N_2502,N_4375);
nand U10322 (N_10322,N_42,N_2145);
nand U10323 (N_10323,N_5520,N_4319);
nor U10324 (N_10324,N_1652,N_4075);
or U10325 (N_10325,N_5533,N_3876);
xnor U10326 (N_10326,N_3021,N_2999);
nand U10327 (N_10327,N_128,N_1991);
nand U10328 (N_10328,N_223,N_4457);
nand U10329 (N_10329,N_5382,N_1664);
nor U10330 (N_10330,N_4982,N_2433);
nand U10331 (N_10331,N_412,N_4523);
xor U10332 (N_10332,N_4456,N_2568);
nor U10333 (N_10333,N_3703,N_1340);
nand U10334 (N_10334,N_3261,N_2049);
and U10335 (N_10335,N_3825,N_3256);
xor U10336 (N_10336,N_4223,N_2778);
and U10337 (N_10337,N_459,N_1125);
and U10338 (N_10338,N_2075,N_5746);
and U10339 (N_10339,N_240,N_3686);
nor U10340 (N_10340,N_4495,N_138);
nand U10341 (N_10341,N_5837,N_1337);
nand U10342 (N_10342,N_1698,N_4148);
and U10343 (N_10343,N_309,N_2523);
nor U10344 (N_10344,N_5579,N_1396);
or U10345 (N_10345,N_636,N_401);
nor U10346 (N_10346,N_2089,N_1456);
or U10347 (N_10347,N_5075,N_603);
xnor U10348 (N_10348,N_4222,N_717);
xnor U10349 (N_10349,N_712,N_2965);
nor U10350 (N_10350,N_182,N_1142);
or U10351 (N_10351,N_1860,N_3441);
or U10352 (N_10352,N_3215,N_659);
and U10353 (N_10353,N_893,N_760);
xor U10354 (N_10354,N_4201,N_295);
nor U10355 (N_10355,N_5837,N_2606);
nor U10356 (N_10356,N_1174,N_4115);
or U10357 (N_10357,N_1254,N_82);
xnor U10358 (N_10358,N_5521,N_3773);
xnor U10359 (N_10359,N_389,N_1851);
nor U10360 (N_10360,N_5667,N_5487);
and U10361 (N_10361,N_2418,N_1433);
and U10362 (N_10362,N_3832,N_2678);
nor U10363 (N_10363,N_2386,N_4651);
xnor U10364 (N_10364,N_1105,N_5677);
xor U10365 (N_10365,N_2510,N_3224);
nand U10366 (N_10366,N_3425,N_2663);
nor U10367 (N_10367,N_3148,N_653);
nor U10368 (N_10368,N_1107,N_1249);
xor U10369 (N_10369,N_196,N_3261);
xnor U10370 (N_10370,N_5206,N_3216);
or U10371 (N_10371,N_3979,N_2261);
and U10372 (N_10372,N_1492,N_5158);
nand U10373 (N_10373,N_161,N_4625);
nand U10374 (N_10374,N_3971,N_173);
xor U10375 (N_10375,N_506,N_3165);
xnor U10376 (N_10376,N_4947,N_5740);
nor U10377 (N_10377,N_5541,N_2509);
nand U10378 (N_10378,N_882,N_1255);
nor U10379 (N_10379,N_5155,N_436);
xnor U10380 (N_10380,N_5735,N_3255);
nand U10381 (N_10381,N_1300,N_1866);
nor U10382 (N_10382,N_147,N_5147);
xor U10383 (N_10383,N_5664,N_3843);
or U10384 (N_10384,N_1190,N_2285);
and U10385 (N_10385,N_4125,N_4014);
xnor U10386 (N_10386,N_687,N_865);
and U10387 (N_10387,N_5790,N_4939);
xor U10388 (N_10388,N_2558,N_1737);
xnor U10389 (N_10389,N_3089,N_3529);
or U10390 (N_10390,N_4105,N_2381);
nor U10391 (N_10391,N_3461,N_3453);
and U10392 (N_10392,N_2705,N_4798);
xor U10393 (N_10393,N_4539,N_2913);
nor U10394 (N_10394,N_4981,N_3175);
nand U10395 (N_10395,N_1231,N_3069);
or U10396 (N_10396,N_5998,N_207);
and U10397 (N_10397,N_1488,N_263);
nand U10398 (N_10398,N_3903,N_1681);
or U10399 (N_10399,N_3860,N_5912);
nor U10400 (N_10400,N_169,N_810);
xnor U10401 (N_10401,N_129,N_1802);
or U10402 (N_10402,N_1593,N_2998);
or U10403 (N_10403,N_5770,N_5542);
nand U10404 (N_10404,N_3909,N_4179);
nor U10405 (N_10405,N_2914,N_128);
xnor U10406 (N_10406,N_1512,N_5811);
xor U10407 (N_10407,N_3093,N_4361);
nor U10408 (N_10408,N_4253,N_5044);
and U10409 (N_10409,N_967,N_2501);
and U10410 (N_10410,N_4772,N_4049);
and U10411 (N_10411,N_5670,N_1340);
nor U10412 (N_10412,N_2787,N_2675);
nand U10413 (N_10413,N_556,N_1569);
nor U10414 (N_10414,N_3937,N_4495);
or U10415 (N_10415,N_1399,N_1196);
or U10416 (N_10416,N_3046,N_1892);
or U10417 (N_10417,N_3120,N_3971);
nor U10418 (N_10418,N_575,N_1910);
and U10419 (N_10419,N_3361,N_2757);
and U10420 (N_10420,N_5972,N_1590);
and U10421 (N_10421,N_1801,N_4129);
and U10422 (N_10422,N_1648,N_5097);
nor U10423 (N_10423,N_2034,N_1717);
nand U10424 (N_10424,N_709,N_3552);
nand U10425 (N_10425,N_5507,N_5537);
nand U10426 (N_10426,N_2559,N_3097);
nor U10427 (N_10427,N_5857,N_3532);
or U10428 (N_10428,N_2478,N_434);
xnor U10429 (N_10429,N_2285,N_2910);
or U10430 (N_10430,N_1102,N_365);
xor U10431 (N_10431,N_3264,N_5425);
nand U10432 (N_10432,N_2883,N_3036);
xnor U10433 (N_10433,N_5558,N_1043);
or U10434 (N_10434,N_1663,N_5148);
xnor U10435 (N_10435,N_5551,N_4504);
xnor U10436 (N_10436,N_3603,N_3571);
and U10437 (N_10437,N_1958,N_173);
or U10438 (N_10438,N_4523,N_4866);
or U10439 (N_10439,N_2766,N_5034);
xor U10440 (N_10440,N_5518,N_4765);
and U10441 (N_10441,N_5111,N_178);
xor U10442 (N_10442,N_2685,N_5447);
xnor U10443 (N_10443,N_4087,N_5965);
nor U10444 (N_10444,N_5778,N_1445);
or U10445 (N_10445,N_2919,N_434);
nand U10446 (N_10446,N_2207,N_1512);
and U10447 (N_10447,N_2058,N_5681);
nor U10448 (N_10448,N_2358,N_2659);
and U10449 (N_10449,N_4697,N_3962);
nand U10450 (N_10450,N_3425,N_3509);
xnor U10451 (N_10451,N_2793,N_5554);
or U10452 (N_10452,N_3418,N_3397);
xnor U10453 (N_10453,N_5810,N_5460);
nor U10454 (N_10454,N_1063,N_520);
nor U10455 (N_10455,N_5786,N_3809);
xor U10456 (N_10456,N_990,N_4551);
nor U10457 (N_10457,N_1956,N_1539);
nand U10458 (N_10458,N_2955,N_632);
nand U10459 (N_10459,N_14,N_2155);
or U10460 (N_10460,N_2422,N_4484);
nand U10461 (N_10461,N_4411,N_5295);
or U10462 (N_10462,N_2318,N_5567);
and U10463 (N_10463,N_2667,N_375);
nand U10464 (N_10464,N_1685,N_3459);
nor U10465 (N_10465,N_1851,N_4377);
or U10466 (N_10466,N_813,N_5269);
nor U10467 (N_10467,N_57,N_4778);
and U10468 (N_10468,N_944,N_5887);
nor U10469 (N_10469,N_628,N_3936);
nor U10470 (N_10470,N_1027,N_2673);
nand U10471 (N_10471,N_1496,N_2602);
nand U10472 (N_10472,N_1232,N_2226);
xor U10473 (N_10473,N_4889,N_1162);
or U10474 (N_10474,N_1533,N_3416);
nor U10475 (N_10475,N_1390,N_1372);
nand U10476 (N_10476,N_2944,N_5067);
nor U10477 (N_10477,N_4962,N_2456);
and U10478 (N_10478,N_5522,N_2854);
and U10479 (N_10479,N_3877,N_4659);
or U10480 (N_10480,N_2742,N_4837);
nor U10481 (N_10481,N_3835,N_3504);
xor U10482 (N_10482,N_636,N_4190);
nor U10483 (N_10483,N_2473,N_618);
or U10484 (N_10484,N_2185,N_816);
xor U10485 (N_10485,N_5213,N_2741);
nand U10486 (N_10486,N_174,N_3113);
or U10487 (N_10487,N_5268,N_2142);
and U10488 (N_10488,N_2112,N_1574);
and U10489 (N_10489,N_4179,N_5889);
or U10490 (N_10490,N_3548,N_1924);
nor U10491 (N_10491,N_4304,N_1890);
xnor U10492 (N_10492,N_5993,N_2290);
nor U10493 (N_10493,N_5391,N_2860);
and U10494 (N_10494,N_1494,N_3798);
xnor U10495 (N_10495,N_3043,N_966);
xor U10496 (N_10496,N_3502,N_404);
nor U10497 (N_10497,N_1516,N_2070);
nor U10498 (N_10498,N_4044,N_1522);
nand U10499 (N_10499,N_1355,N_3531);
nor U10500 (N_10500,N_1628,N_2379);
nand U10501 (N_10501,N_227,N_3822);
and U10502 (N_10502,N_302,N_3523);
or U10503 (N_10503,N_2190,N_4298);
xor U10504 (N_10504,N_100,N_3037);
and U10505 (N_10505,N_3058,N_2643);
nand U10506 (N_10506,N_4954,N_3490);
xnor U10507 (N_10507,N_3699,N_989);
nor U10508 (N_10508,N_1727,N_2934);
and U10509 (N_10509,N_4874,N_3095);
nor U10510 (N_10510,N_4915,N_894);
and U10511 (N_10511,N_4994,N_2545);
or U10512 (N_10512,N_3882,N_619);
xnor U10513 (N_10513,N_1687,N_5829);
nor U10514 (N_10514,N_4213,N_4254);
nor U10515 (N_10515,N_1659,N_3210);
and U10516 (N_10516,N_1763,N_467);
nor U10517 (N_10517,N_1652,N_4690);
or U10518 (N_10518,N_5214,N_5099);
or U10519 (N_10519,N_1614,N_3725);
nand U10520 (N_10520,N_5840,N_5381);
or U10521 (N_10521,N_4525,N_1202);
and U10522 (N_10522,N_5318,N_1928);
or U10523 (N_10523,N_574,N_3650);
and U10524 (N_10524,N_2071,N_245);
or U10525 (N_10525,N_5842,N_2284);
or U10526 (N_10526,N_3096,N_1638);
and U10527 (N_10527,N_1738,N_5967);
nor U10528 (N_10528,N_3719,N_3008);
and U10529 (N_10529,N_1748,N_844);
and U10530 (N_10530,N_1857,N_5809);
or U10531 (N_10531,N_523,N_5828);
and U10532 (N_10532,N_1876,N_4183);
and U10533 (N_10533,N_2629,N_1003);
and U10534 (N_10534,N_1032,N_5131);
nand U10535 (N_10535,N_4802,N_4336);
nand U10536 (N_10536,N_3921,N_3211);
nand U10537 (N_10537,N_2015,N_4663);
xor U10538 (N_10538,N_536,N_3055);
xnor U10539 (N_10539,N_732,N_1723);
nor U10540 (N_10540,N_3152,N_4854);
xor U10541 (N_10541,N_584,N_5833);
nand U10542 (N_10542,N_3876,N_5760);
and U10543 (N_10543,N_407,N_2080);
and U10544 (N_10544,N_2710,N_5997);
or U10545 (N_10545,N_1689,N_1365);
and U10546 (N_10546,N_2666,N_4878);
or U10547 (N_10547,N_61,N_2902);
or U10548 (N_10548,N_4179,N_5007);
nand U10549 (N_10549,N_4082,N_4539);
nor U10550 (N_10550,N_3349,N_3897);
or U10551 (N_10551,N_1752,N_5558);
and U10552 (N_10552,N_1895,N_254);
or U10553 (N_10553,N_5930,N_3392);
nand U10554 (N_10554,N_5428,N_3904);
and U10555 (N_10555,N_1391,N_61);
nand U10556 (N_10556,N_1304,N_2956);
and U10557 (N_10557,N_3324,N_2812);
nand U10558 (N_10558,N_3929,N_4220);
xnor U10559 (N_10559,N_5756,N_3443);
nor U10560 (N_10560,N_436,N_5452);
nand U10561 (N_10561,N_4338,N_14);
nand U10562 (N_10562,N_5431,N_4408);
nor U10563 (N_10563,N_5777,N_5600);
or U10564 (N_10564,N_2375,N_3298);
nand U10565 (N_10565,N_5335,N_4444);
xnor U10566 (N_10566,N_2088,N_2362);
or U10567 (N_10567,N_1166,N_4432);
or U10568 (N_10568,N_3438,N_3150);
or U10569 (N_10569,N_5919,N_5651);
and U10570 (N_10570,N_5723,N_4346);
and U10571 (N_10571,N_185,N_2817);
xnor U10572 (N_10572,N_5197,N_1238);
nor U10573 (N_10573,N_2378,N_3523);
nor U10574 (N_10574,N_33,N_1680);
xnor U10575 (N_10575,N_3566,N_5774);
or U10576 (N_10576,N_2999,N_382);
nand U10577 (N_10577,N_4401,N_1342);
xnor U10578 (N_10578,N_1394,N_431);
or U10579 (N_10579,N_5343,N_4832);
xor U10580 (N_10580,N_5551,N_4907);
xor U10581 (N_10581,N_3520,N_527);
nor U10582 (N_10582,N_3735,N_558);
nor U10583 (N_10583,N_1953,N_2167);
nor U10584 (N_10584,N_3993,N_81);
xor U10585 (N_10585,N_1338,N_2590);
or U10586 (N_10586,N_3649,N_4503);
nand U10587 (N_10587,N_2081,N_1925);
or U10588 (N_10588,N_2882,N_3130);
nand U10589 (N_10589,N_3494,N_1868);
or U10590 (N_10590,N_986,N_1944);
xnor U10591 (N_10591,N_1807,N_3224);
or U10592 (N_10592,N_1933,N_5237);
nor U10593 (N_10593,N_1729,N_594);
and U10594 (N_10594,N_205,N_3822);
nand U10595 (N_10595,N_2415,N_3931);
xnor U10596 (N_10596,N_4019,N_1400);
or U10597 (N_10597,N_3747,N_137);
nor U10598 (N_10598,N_4959,N_2862);
and U10599 (N_10599,N_4880,N_4411);
xnor U10600 (N_10600,N_1251,N_739);
and U10601 (N_10601,N_4193,N_4626);
and U10602 (N_10602,N_5411,N_3004);
and U10603 (N_10603,N_2715,N_1259);
xor U10604 (N_10604,N_2553,N_740);
nor U10605 (N_10605,N_5353,N_5073);
nor U10606 (N_10606,N_1216,N_1253);
nor U10607 (N_10607,N_759,N_1774);
xnor U10608 (N_10608,N_2671,N_1515);
and U10609 (N_10609,N_1885,N_0);
nor U10610 (N_10610,N_1009,N_830);
and U10611 (N_10611,N_2427,N_4341);
nand U10612 (N_10612,N_312,N_3483);
xor U10613 (N_10613,N_398,N_3029);
nand U10614 (N_10614,N_2075,N_5925);
nor U10615 (N_10615,N_5470,N_874);
and U10616 (N_10616,N_556,N_1345);
nor U10617 (N_10617,N_81,N_264);
nor U10618 (N_10618,N_4834,N_2946);
and U10619 (N_10619,N_266,N_1458);
or U10620 (N_10620,N_120,N_5755);
and U10621 (N_10621,N_5578,N_5576);
nand U10622 (N_10622,N_2093,N_156);
nor U10623 (N_10623,N_817,N_5423);
nand U10624 (N_10624,N_2619,N_167);
or U10625 (N_10625,N_2202,N_4630);
nor U10626 (N_10626,N_5634,N_1976);
and U10627 (N_10627,N_2017,N_2814);
xor U10628 (N_10628,N_2641,N_2823);
xor U10629 (N_10629,N_866,N_3747);
nand U10630 (N_10630,N_4475,N_3839);
and U10631 (N_10631,N_3307,N_1114);
and U10632 (N_10632,N_1798,N_384);
nor U10633 (N_10633,N_5287,N_214);
or U10634 (N_10634,N_1282,N_259);
xnor U10635 (N_10635,N_1288,N_4911);
nand U10636 (N_10636,N_1513,N_3953);
nand U10637 (N_10637,N_1726,N_354);
or U10638 (N_10638,N_3310,N_1491);
xor U10639 (N_10639,N_2959,N_4003);
or U10640 (N_10640,N_4491,N_4538);
or U10641 (N_10641,N_5459,N_5170);
nand U10642 (N_10642,N_2981,N_5640);
or U10643 (N_10643,N_2064,N_747);
nor U10644 (N_10644,N_1608,N_727);
and U10645 (N_10645,N_3914,N_3341);
xor U10646 (N_10646,N_1053,N_642);
xor U10647 (N_10647,N_2652,N_3253);
nor U10648 (N_10648,N_5971,N_3889);
nand U10649 (N_10649,N_2894,N_39);
xor U10650 (N_10650,N_105,N_1182);
nand U10651 (N_10651,N_4510,N_5516);
xnor U10652 (N_10652,N_3338,N_3082);
xor U10653 (N_10653,N_502,N_4922);
and U10654 (N_10654,N_5694,N_3445);
or U10655 (N_10655,N_2392,N_3864);
nor U10656 (N_10656,N_5674,N_1402);
and U10657 (N_10657,N_1569,N_295);
xnor U10658 (N_10658,N_4675,N_2840);
nor U10659 (N_10659,N_4728,N_2018);
nand U10660 (N_10660,N_1060,N_1101);
nor U10661 (N_10661,N_3480,N_2337);
or U10662 (N_10662,N_5673,N_479);
nand U10663 (N_10663,N_2740,N_772);
and U10664 (N_10664,N_1797,N_3882);
nor U10665 (N_10665,N_5814,N_4290);
and U10666 (N_10666,N_4186,N_1922);
nor U10667 (N_10667,N_1573,N_3026);
nand U10668 (N_10668,N_1783,N_5871);
nor U10669 (N_10669,N_3503,N_3104);
nand U10670 (N_10670,N_3082,N_4670);
nor U10671 (N_10671,N_3528,N_4690);
nor U10672 (N_10672,N_5130,N_5305);
xnor U10673 (N_10673,N_5491,N_2267);
nand U10674 (N_10674,N_3705,N_492);
and U10675 (N_10675,N_241,N_1095);
nand U10676 (N_10676,N_5650,N_3299);
nor U10677 (N_10677,N_2871,N_4421);
nand U10678 (N_10678,N_1515,N_2439);
xnor U10679 (N_10679,N_3134,N_610);
nand U10680 (N_10680,N_3553,N_3631);
nand U10681 (N_10681,N_5652,N_1802);
nand U10682 (N_10682,N_326,N_4528);
and U10683 (N_10683,N_4573,N_5144);
nor U10684 (N_10684,N_5278,N_611);
nor U10685 (N_10685,N_3780,N_1931);
and U10686 (N_10686,N_1726,N_3657);
and U10687 (N_10687,N_2782,N_548);
and U10688 (N_10688,N_3417,N_5342);
nor U10689 (N_10689,N_2575,N_5195);
nor U10690 (N_10690,N_389,N_4709);
nand U10691 (N_10691,N_3028,N_3295);
and U10692 (N_10692,N_2036,N_3413);
and U10693 (N_10693,N_4689,N_5252);
xor U10694 (N_10694,N_4198,N_5834);
nor U10695 (N_10695,N_5188,N_1829);
xnor U10696 (N_10696,N_5229,N_4106);
xnor U10697 (N_10697,N_3426,N_5387);
nand U10698 (N_10698,N_3324,N_4153);
xnor U10699 (N_10699,N_5484,N_4892);
xor U10700 (N_10700,N_2181,N_4439);
nand U10701 (N_10701,N_257,N_2671);
and U10702 (N_10702,N_2925,N_3848);
or U10703 (N_10703,N_3791,N_2449);
xnor U10704 (N_10704,N_5455,N_2831);
nor U10705 (N_10705,N_2953,N_165);
and U10706 (N_10706,N_1341,N_4387);
xor U10707 (N_10707,N_1260,N_5731);
nand U10708 (N_10708,N_1406,N_2928);
and U10709 (N_10709,N_2662,N_1098);
xor U10710 (N_10710,N_1378,N_3981);
or U10711 (N_10711,N_1703,N_2718);
xnor U10712 (N_10712,N_1250,N_2880);
xor U10713 (N_10713,N_3215,N_5638);
nand U10714 (N_10714,N_1801,N_1735);
xor U10715 (N_10715,N_2383,N_2133);
or U10716 (N_10716,N_3718,N_4895);
and U10717 (N_10717,N_3385,N_2909);
or U10718 (N_10718,N_3724,N_2258);
xor U10719 (N_10719,N_1607,N_4758);
nor U10720 (N_10720,N_2005,N_3648);
and U10721 (N_10721,N_16,N_2522);
nor U10722 (N_10722,N_3363,N_162);
nor U10723 (N_10723,N_1891,N_3766);
nand U10724 (N_10724,N_1055,N_3895);
and U10725 (N_10725,N_5597,N_3546);
or U10726 (N_10726,N_357,N_3638);
nand U10727 (N_10727,N_1123,N_3575);
or U10728 (N_10728,N_3619,N_1345);
nor U10729 (N_10729,N_3941,N_520);
nor U10730 (N_10730,N_5357,N_1545);
xor U10731 (N_10731,N_3065,N_4710);
nand U10732 (N_10732,N_5801,N_3940);
xor U10733 (N_10733,N_5997,N_1216);
nand U10734 (N_10734,N_2256,N_4888);
and U10735 (N_10735,N_2211,N_5179);
nor U10736 (N_10736,N_4049,N_1955);
or U10737 (N_10737,N_2233,N_1514);
xor U10738 (N_10738,N_965,N_3220);
and U10739 (N_10739,N_339,N_717);
and U10740 (N_10740,N_2139,N_3667);
nand U10741 (N_10741,N_2281,N_3445);
nor U10742 (N_10742,N_5359,N_520);
nand U10743 (N_10743,N_5693,N_707);
nor U10744 (N_10744,N_5668,N_2797);
nand U10745 (N_10745,N_5551,N_4977);
and U10746 (N_10746,N_5730,N_4177);
and U10747 (N_10747,N_1127,N_3243);
xnor U10748 (N_10748,N_3864,N_5717);
nor U10749 (N_10749,N_1172,N_2816);
nand U10750 (N_10750,N_2295,N_427);
nor U10751 (N_10751,N_1555,N_1774);
or U10752 (N_10752,N_4870,N_4479);
nand U10753 (N_10753,N_2065,N_2426);
and U10754 (N_10754,N_4273,N_3963);
nor U10755 (N_10755,N_3621,N_1573);
nor U10756 (N_10756,N_801,N_2941);
or U10757 (N_10757,N_506,N_432);
and U10758 (N_10758,N_2959,N_1559);
nor U10759 (N_10759,N_2719,N_1801);
or U10760 (N_10760,N_2153,N_2388);
xor U10761 (N_10761,N_4522,N_3727);
and U10762 (N_10762,N_5418,N_3827);
nand U10763 (N_10763,N_5367,N_5394);
nand U10764 (N_10764,N_4894,N_2882);
or U10765 (N_10765,N_2932,N_2145);
nor U10766 (N_10766,N_5740,N_4528);
xor U10767 (N_10767,N_561,N_5005);
or U10768 (N_10768,N_2481,N_753);
nand U10769 (N_10769,N_4773,N_233);
nand U10770 (N_10770,N_4097,N_712);
or U10771 (N_10771,N_3059,N_5637);
xnor U10772 (N_10772,N_4680,N_5205);
nand U10773 (N_10773,N_4452,N_1156);
xor U10774 (N_10774,N_1026,N_5648);
xor U10775 (N_10775,N_302,N_3860);
and U10776 (N_10776,N_2528,N_4477);
nand U10777 (N_10777,N_4222,N_3087);
xor U10778 (N_10778,N_2176,N_4713);
or U10779 (N_10779,N_4413,N_1418);
xnor U10780 (N_10780,N_2842,N_853);
and U10781 (N_10781,N_783,N_1350);
nor U10782 (N_10782,N_5548,N_5589);
nor U10783 (N_10783,N_5394,N_4962);
or U10784 (N_10784,N_5164,N_275);
nor U10785 (N_10785,N_2232,N_1252);
or U10786 (N_10786,N_2076,N_5106);
or U10787 (N_10787,N_3422,N_3364);
xor U10788 (N_10788,N_2902,N_2756);
and U10789 (N_10789,N_4880,N_4824);
nor U10790 (N_10790,N_2513,N_4468);
and U10791 (N_10791,N_323,N_143);
nand U10792 (N_10792,N_1833,N_2094);
nand U10793 (N_10793,N_3494,N_3724);
nand U10794 (N_10794,N_470,N_3065);
and U10795 (N_10795,N_2959,N_905);
xor U10796 (N_10796,N_5807,N_1399);
nand U10797 (N_10797,N_4093,N_5392);
nand U10798 (N_10798,N_1115,N_2189);
and U10799 (N_10799,N_2961,N_3610);
nand U10800 (N_10800,N_1357,N_2329);
xor U10801 (N_10801,N_2523,N_4733);
and U10802 (N_10802,N_4667,N_275);
nor U10803 (N_10803,N_1422,N_4156);
and U10804 (N_10804,N_2566,N_2780);
or U10805 (N_10805,N_4357,N_1732);
or U10806 (N_10806,N_752,N_4343);
nand U10807 (N_10807,N_5378,N_2108);
xnor U10808 (N_10808,N_2483,N_1273);
nor U10809 (N_10809,N_3458,N_1886);
nand U10810 (N_10810,N_4986,N_5111);
nor U10811 (N_10811,N_1534,N_5928);
or U10812 (N_10812,N_3256,N_2773);
and U10813 (N_10813,N_1051,N_2004);
nand U10814 (N_10814,N_2208,N_608);
nor U10815 (N_10815,N_1018,N_4862);
nand U10816 (N_10816,N_4601,N_12);
or U10817 (N_10817,N_1617,N_3887);
nand U10818 (N_10818,N_4239,N_1784);
nor U10819 (N_10819,N_394,N_3637);
nor U10820 (N_10820,N_4508,N_3681);
or U10821 (N_10821,N_5568,N_1433);
and U10822 (N_10822,N_4525,N_421);
nor U10823 (N_10823,N_1577,N_5958);
and U10824 (N_10824,N_4128,N_4143);
xor U10825 (N_10825,N_5841,N_3605);
nand U10826 (N_10826,N_2228,N_5618);
or U10827 (N_10827,N_1178,N_4727);
nor U10828 (N_10828,N_1431,N_1019);
nand U10829 (N_10829,N_2679,N_1132);
xor U10830 (N_10830,N_2685,N_2860);
xor U10831 (N_10831,N_1122,N_4443);
nand U10832 (N_10832,N_2897,N_2560);
nor U10833 (N_10833,N_1443,N_5495);
nor U10834 (N_10834,N_1813,N_3307);
and U10835 (N_10835,N_4560,N_4035);
xnor U10836 (N_10836,N_4173,N_560);
nor U10837 (N_10837,N_4530,N_1578);
and U10838 (N_10838,N_877,N_2329);
xor U10839 (N_10839,N_4561,N_2204);
xnor U10840 (N_10840,N_3864,N_4460);
or U10841 (N_10841,N_1149,N_4453);
or U10842 (N_10842,N_3762,N_3715);
and U10843 (N_10843,N_5518,N_2535);
or U10844 (N_10844,N_5594,N_2519);
or U10845 (N_10845,N_2419,N_1560);
xor U10846 (N_10846,N_3737,N_4058);
nor U10847 (N_10847,N_4758,N_5195);
nor U10848 (N_10848,N_1921,N_5618);
or U10849 (N_10849,N_2881,N_922);
or U10850 (N_10850,N_1604,N_1717);
or U10851 (N_10851,N_4730,N_2382);
xnor U10852 (N_10852,N_5661,N_3075);
nand U10853 (N_10853,N_5102,N_1429);
and U10854 (N_10854,N_1665,N_517);
nor U10855 (N_10855,N_5507,N_4299);
and U10856 (N_10856,N_565,N_4083);
or U10857 (N_10857,N_929,N_3826);
nor U10858 (N_10858,N_5138,N_3045);
and U10859 (N_10859,N_2851,N_2604);
nor U10860 (N_10860,N_3035,N_1174);
and U10861 (N_10861,N_3030,N_3073);
nor U10862 (N_10862,N_4248,N_1396);
or U10863 (N_10863,N_4239,N_2463);
or U10864 (N_10864,N_1541,N_4607);
nor U10865 (N_10865,N_5234,N_132);
and U10866 (N_10866,N_2099,N_5921);
xnor U10867 (N_10867,N_5995,N_3437);
nor U10868 (N_10868,N_4433,N_2972);
or U10869 (N_10869,N_2704,N_2628);
or U10870 (N_10870,N_3009,N_1394);
nand U10871 (N_10871,N_2275,N_1607);
nor U10872 (N_10872,N_4227,N_4796);
xor U10873 (N_10873,N_5747,N_5619);
xnor U10874 (N_10874,N_549,N_1010);
nor U10875 (N_10875,N_254,N_1777);
nor U10876 (N_10876,N_4554,N_3373);
xnor U10877 (N_10877,N_2951,N_3955);
and U10878 (N_10878,N_5496,N_5744);
and U10879 (N_10879,N_5096,N_5028);
or U10880 (N_10880,N_2278,N_4077);
xnor U10881 (N_10881,N_5484,N_899);
nand U10882 (N_10882,N_2517,N_78);
and U10883 (N_10883,N_827,N_1219);
and U10884 (N_10884,N_3821,N_5491);
or U10885 (N_10885,N_3318,N_1997);
nand U10886 (N_10886,N_4461,N_2100);
nor U10887 (N_10887,N_239,N_392);
and U10888 (N_10888,N_5254,N_2768);
nor U10889 (N_10889,N_5695,N_4712);
and U10890 (N_10890,N_4046,N_5218);
or U10891 (N_10891,N_98,N_2249);
or U10892 (N_10892,N_3259,N_1897);
nor U10893 (N_10893,N_4291,N_3875);
and U10894 (N_10894,N_5155,N_390);
xnor U10895 (N_10895,N_1595,N_1043);
or U10896 (N_10896,N_4154,N_3805);
nor U10897 (N_10897,N_1617,N_2687);
or U10898 (N_10898,N_2230,N_3906);
or U10899 (N_10899,N_3447,N_4770);
or U10900 (N_10900,N_374,N_4470);
or U10901 (N_10901,N_4360,N_4015);
nand U10902 (N_10902,N_3225,N_1190);
xnor U10903 (N_10903,N_2042,N_100);
xnor U10904 (N_10904,N_2482,N_656);
xnor U10905 (N_10905,N_2834,N_3983);
xnor U10906 (N_10906,N_351,N_3178);
nor U10907 (N_10907,N_5757,N_2175);
or U10908 (N_10908,N_3153,N_1061);
and U10909 (N_10909,N_390,N_5957);
nor U10910 (N_10910,N_1342,N_2354);
nor U10911 (N_10911,N_856,N_2080);
nand U10912 (N_10912,N_2467,N_151);
xnor U10913 (N_10913,N_424,N_480);
nand U10914 (N_10914,N_1963,N_4871);
nand U10915 (N_10915,N_2107,N_3953);
nor U10916 (N_10916,N_3791,N_5315);
nor U10917 (N_10917,N_474,N_2535);
and U10918 (N_10918,N_2622,N_1118);
nand U10919 (N_10919,N_1078,N_4795);
or U10920 (N_10920,N_4931,N_964);
xor U10921 (N_10921,N_4515,N_1855);
and U10922 (N_10922,N_1955,N_5785);
xor U10923 (N_10923,N_3818,N_2634);
nand U10924 (N_10924,N_5099,N_1040);
and U10925 (N_10925,N_4948,N_5786);
and U10926 (N_10926,N_1148,N_1218);
and U10927 (N_10927,N_3586,N_5930);
and U10928 (N_10928,N_3284,N_5027);
or U10929 (N_10929,N_596,N_4288);
nor U10930 (N_10930,N_3157,N_2976);
nor U10931 (N_10931,N_5160,N_2234);
xor U10932 (N_10932,N_5766,N_4463);
xnor U10933 (N_10933,N_1790,N_5977);
xnor U10934 (N_10934,N_94,N_398);
xor U10935 (N_10935,N_5934,N_3530);
xnor U10936 (N_10936,N_3398,N_2012);
nor U10937 (N_10937,N_1210,N_922);
nor U10938 (N_10938,N_1300,N_3903);
and U10939 (N_10939,N_240,N_1218);
and U10940 (N_10940,N_1475,N_4848);
or U10941 (N_10941,N_1434,N_4746);
nand U10942 (N_10942,N_5305,N_5360);
or U10943 (N_10943,N_3190,N_5617);
or U10944 (N_10944,N_4745,N_3);
or U10945 (N_10945,N_145,N_2780);
or U10946 (N_10946,N_5544,N_3338);
and U10947 (N_10947,N_4056,N_4694);
nand U10948 (N_10948,N_4141,N_5516);
or U10949 (N_10949,N_968,N_5694);
nand U10950 (N_10950,N_2972,N_1925);
or U10951 (N_10951,N_739,N_1185);
or U10952 (N_10952,N_2357,N_2286);
and U10953 (N_10953,N_3846,N_5760);
and U10954 (N_10954,N_5874,N_5262);
or U10955 (N_10955,N_3822,N_4616);
and U10956 (N_10956,N_1552,N_3673);
xor U10957 (N_10957,N_69,N_4969);
nor U10958 (N_10958,N_2537,N_4577);
nand U10959 (N_10959,N_5954,N_474);
and U10960 (N_10960,N_688,N_4989);
or U10961 (N_10961,N_724,N_558);
and U10962 (N_10962,N_2159,N_1513);
nor U10963 (N_10963,N_5956,N_1701);
nand U10964 (N_10964,N_4565,N_3206);
nand U10965 (N_10965,N_3941,N_5584);
xor U10966 (N_10966,N_5951,N_5663);
nor U10967 (N_10967,N_4718,N_5170);
or U10968 (N_10968,N_1165,N_891);
nand U10969 (N_10969,N_3786,N_5240);
nor U10970 (N_10970,N_4499,N_4960);
or U10971 (N_10971,N_5511,N_3718);
nand U10972 (N_10972,N_782,N_5511);
nor U10973 (N_10973,N_3975,N_3593);
nand U10974 (N_10974,N_1773,N_2843);
xor U10975 (N_10975,N_4150,N_3154);
or U10976 (N_10976,N_2854,N_191);
nor U10977 (N_10977,N_1563,N_2518);
nor U10978 (N_10978,N_4233,N_2966);
xnor U10979 (N_10979,N_3227,N_2624);
xor U10980 (N_10980,N_4890,N_4299);
or U10981 (N_10981,N_2058,N_3667);
nand U10982 (N_10982,N_928,N_570);
nor U10983 (N_10983,N_288,N_2661);
or U10984 (N_10984,N_673,N_3246);
and U10985 (N_10985,N_4674,N_1593);
nor U10986 (N_10986,N_5626,N_3862);
nand U10987 (N_10987,N_2577,N_369);
nor U10988 (N_10988,N_5484,N_5828);
or U10989 (N_10989,N_4452,N_5351);
or U10990 (N_10990,N_4726,N_3786);
or U10991 (N_10991,N_1828,N_3358);
xor U10992 (N_10992,N_4163,N_477);
nor U10993 (N_10993,N_2028,N_4737);
nand U10994 (N_10994,N_2815,N_3974);
or U10995 (N_10995,N_5177,N_32);
xor U10996 (N_10996,N_5146,N_1825);
or U10997 (N_10997,N_5525,N_1020);
and U10998 (N_10998,N_689,N_1881);
nor U10999 (N_10999,N_1276,N_3485);
nand U11000 (N_11000,N_3466,N_44);
xor U11001 (N_11001,N_1307,N_1355);
xnor U11002 (N_11002,N_2120,N_1525);
nand U11003 (N_11003,N_4246,N_4223);
nor U11004 (N_11004,N_958,N_4120);
nor U11005 (N_11005,N_3505,N_5159);
xnor U11006 (N_11006,N_3414,N_3207);
xor U11007 (N_11007,N_2570,N_5827);
nor U11008 (N_11008,N_1536,N_5327);
and U11009 (N_11009,N_4295,N_444);
and U11010 (N_11010,N_5309,N_3208);
nor U11011 (N_11011,N_442,N_3124);
and U11012 (N_11012,N_3954,N_5552);
nand U11013 (N_11013,N_3744,N_1125);
xnor U11014 (N_11014,N_2182,N_5597);
xnor U11015 (N_11015,N_700,N_5773);
and U11016 (N_11016,N_4562,N_1854);
nor U11017 (N_11017,N_4881,N_3647);
or U11018 (N_11018,N_707,N_2037);
nand U11019 (N_11019,N_1686,N_4915);
xor U11020 (N_11020,N_5942,N_1875);
nand U11021 (N_11021,N_5119,N_4547);
xnor U11022 (N_11022,N_3069,N_2655);
and U11023 (N_11023,N_1621,N_634);
nor U11024 (N_11024,N_4638,N_263);
or U11025 (N_11025,N_5600,N_300);
nand U11026 (N_11026,N_1960,N_379);
xor U11027 (N_11027,N_1783,N_1436);
xor U11028 (N_11028,N_4092,N_1612);
and U11029 (N_11029,N_3446,N_4197);
nand U11030 (N_11030,N_3005,N_4511);
or U11031 (N_11031,N_3798,N_4640);
or U11032 (N_11032,N_5401,N_4618);
nand U11033 (N_11033,N_5786,N_2612);
nand U11034 (N_11034,N_5414,N_255);
nor U11035 (N_11035,N_2705,N_2307);
xor U11036 (N_11036,N_4454,N_2408);
or U11037 (N_11037,N_4069,N_1008);
nor U11038 (N_11038,N_3631,N_5289);
nand U11039 (N_11039,N_5359,N_5123);
nand U11040 (N_11040,N_266,N_367);
nor U11041 (N_11041,N_1166,N_3906);
nor U11042 (N_11042,N_4533,N_2702);
or U11043 (N_11043,N_497,N_5086);
or U11044 (N_11044,N_3134,N_54);
nor U11045 (N_11045,N_5381,N_479);
nand U11046 (N_11046,N_5576,N_5239);
nand U11047 (N_11047,N_1226,N_550);
or U11048 (N_11048,N_1271,N_908);
and U11049 (N_11049,N_5389,N_321);
nand U11050 (N_11050,N_4602,N_873);
or U11051 (N_11051,N_1166,N_2533);
nand U11052 (N_11052,N_4312,N_5341);
nor U11053 (N_11053,N_1233,N_764);
and U11054 (N_11054,N_676,N_5239);
xnor U11055 (N_11055,N_722,N_1138);
or U11056 (N_11056,N_5774,N_1407);
xor U11057 (N_11057,N_202,N_5975);
or U11058 (N_11058,N_2125,N_2475);
nand U11059 (N_11059,N_2108,N_2390);
or U11060 (N_11060,N_5852,N_5098);
or U11061 (N_11061,N_1104,N_3680);
xnor U11062 (N_11062,N_516,N_1174);
nand U11063 (N_11063,N_2056,N_576);
nor U11064 (N_11064,N_2982,N_3238);
nor U11065 (N_11065,N_3182,N_3148);
and U11066 (N_11066,N_3022,N_4303);
or U11067 (N_11067,N_5482,N_5813);
or U11068 (N_11068,N_4329,N_5990);
nand U11069 (N_11069,N_2811,N_4961);
nor U11070 (N_11070,N_5310,N_2136);
or U11071 (N_11071,N_3715,N_3367);
nor U11072 (N_11072,N_3257,N_2645);
or U11073 (N_11073,N_5782,N_4054);
nor U11074 (N_11074,N_362,N_703);
xor U11075 (N_11075,N_1468,N_3412);
or U11076 (N_11076,N_566,N_3838);
nand U11077 (N_11077,N_4417,N_4367);
xor U11078 (N_11078,N_490,N_2675);
nor U11079 (N_11079,N_4556,N_4779);
and U11080 (N_11080,N_1868,N_5874);
or U11081 (N_11081,N_2731,N_2210);
and U11082 (N_11082,N_739,N_1950);
or U11083 (N_11083,N_1178,N_2602);
and U11084 (N_11084,N_2339,N_2551);
nand U11085 (N_11085,N_3356,N_3171);
nand U11086 (N_11086,N_4467,N_5458);
nor U11087 (N_11087,N_5523,N_700);
nand U11088 (N_11088,N_5934,N_45);
or U11089 (N_11089,N_5183,N_3539);
nor U11090 (N_11090,N_1301,N_2687);
nor U11091 (N_11091,N_4459,N_802);
nand U11092 (N_11092,N_380,N_4752);
and U11093 (N_11093,N_1543,N_4880);
and U11094 (N_11094,N_1843,N_5083);
and U11095 (N_11095,N_513,N_1364);
or U11096 (N_11096,N_3650,N_2121);
or U11097 (N_11097,N_2123,N_431);
or U11098 (N_11098,N_4604,N_4434);
nor U11099 (N_11099,N_1768,N_1747);
or U11100 (N_11100,N_2222,N_1486);
and U11101 (N_11101,N_292,N_5658);
nor U11102 (N_11102,N_241,N_2309);
nor U11103 (N_11103,N_3913,N_1250);
nand U11104 (N_11104,N_24,N_3031);
nor U11105 (N_11105,N_4546,N_890);
nor U11106 (N_11106,N_4125,N_3427);
and U11107 (N_11107,N_2027,N_3044);
nand U11108 (N_11108,N_5868,N_4128);
or U11109 (N_11109,N_5262,N_698);
xor U11110 (N_11110,N_3731,N_5675);
xnor U11111 (N_11111,N_4833,N_4329);
or U11112 (N_11112,N_3664,N_5316);
and U11113 (N_11113,N_5280,N_5676);
and U11114 (N_11114,N_3313,N_1723);
or U11115 (N_11115,N_5047,N_4785);
xnor U11116 (N_11116,N_2753,N_4878);
xor U11117 (N_11117,N_3167,N_4400);
or U11118 (N_11118,N_3471,N_3305);
xor U11119 (N_11119,N_2161,N_1060);
nand U11120 (N_11120,N_2804,N_3526);
nor U11121 (N_11121,N_2348,N_2711);
or U11122 (N_11122,N_2741,N_731);
and U11123 (N_11123,N_678,N_4342);
or U11124 (N_11124,N_3958,N_2305);
and U11125 (N_11125,N_276,N_4406);
xor U11126 (N_11126,N_966,N_4270);
xor U11127 (N_11127,N_2789,N_1715);
xnor U11128 (N_11128,N_1637,N_5483);
and U11129 (N_11129,N_5096,N_3620);
nor U11130 (N_11130,N_3849,N_749);
nand U11131 (N_11131,N_428,N_4751);
xnor U11132 (N_11132,N_5063,N_515);
and U11133 (N_11133,N_5302,N_49);
nor U11134 (N_11134,N_1595,N_130);
nor U11135 (N_11135,N_4522,N_4635);
xnor U11136 (N_11136,N_1242,N_2646);
and U11137 (N_11137,N_325,N_1987);
nand U11138 (N_11138,N_5003,N_2125);
nor U11139 (N_11139,N_3122,N_1445);
nand U11140 (N_11140,N_4575,N_5584);
xnor U11141 (N_11141,N_158,N_5845);
nor U11142 (N_11142,N_5578,N_2182);
or U11143 (N_11143,N_1863,N_1457);
nand U11144 (N_11144,N_1733,N_5382);
or U11145 (N_11145,N_3174,N_5130);
nor U11146 (N_11146,N_5700,N_2297);
and U11147 (N_11147,N_405,N_666);
nor U11148 (N_11148,N_796,N_4067);
nor U11149 (N_11149,N_2559,N_1517);
nor U11150 (N_11150,N_1879,N_4821);
nand U11151 (N_11151,N_3995,N_3380);
or U11152 (N_11152,N_2296,N_1243);
and U11153 (N_11153,N_4661,N_5219);
xor U11154 (N_11154,N_1422,N_3273);
xnor U11155 (N_11155,N_3972,N_1036);
and U11156 (N_11156,N_1124,N_949);
nand U11157 (N_11157,N_885,N_1353);
or U11158 (N_11158,N_5130,N_661);
nor U11159 (N_11159,N_3262,N_2948);
xnor U11160 (N_11160,N_4413,N_417);
nor U11161 (N_11161,N_2946,N_2303);
nor U11162 (N_11162,N_1038,N_335);
xnor U11163 (N_11163,N_5840,N_406);
nand U11164 (N_11164,N_5998,N_1307);
xor U11165 (N_11165,N_4568,N_4541);
nand U11166 (N_11166,N_4599,N_4587);
nand U11167 (N_11167,N_3679,N_3819);
or U11168 (N_11168,N_5445,N_222);
xnor U11169 (N_11169,N_4488,N_3448);
and U11170 (N_11170,N_1778,N_3609);
or U11171 (N_11171,N_4079,N_76);
nand U11172 (N_11172,N_3023,N_3298);
or U11173 (N_11173,N_1181,N_574);
or U11174 (N_11174,N_2495,N_3386);
nor U11175 (N_11175,N_5407,N_2309);
xnor U11176 (N_11176,N_3049,N_591);
nand U11177 (N_11177,N_2629,N_2757);
nand U11178 (N_11178,N_1625,N_1418);
xor U11179 (N_11179,N_106,N_174);
nand U11180 (N_11180,N_1389,N_3880);
and U11181 (N_11181,N_4697,N_4505);
and U11182 (N_11182,N_5867,N_4115);
nand U11183 (N_11183,N_1298,N_2093);
and U11184 (N_11184,N_3283,N_5203);
or U11185 (N_11185,N_1437,N_3630);
xnor U11186 (N_11186,N_3178,N_3735);
xnor U11187 (N_11187,N_4490,N_119);
xnor U11188 (N_11188,N_5486,N_4019);
xor U11189 (N_11189,N_1564,N_1947);
or U11190 (N_11190,N_3823,N_1135);
and U11191 (N_11191,N_3662,N_5653);
nor U11192 (N_11192,N_3226,N_5921);
nand U11193 (N_11193,N_4811,N_421);
nand U11194 (N_11194,N_4245,N_2021);
nand U11195 (N_11195,N_3740,N_4397);
xnor U11196 (N_11196,N_5476,N_3987);
and U11197 (N_11197,N_2777,N_2933);
and U11198 (N_11198,N_5575,N_3397);
xnor U11199 (N_11199,N_4212,N_910);
xor U11200 (N_11200,N_4165,N_5492);
xnor U11201 (N_11201,N_2748,N_4048);
and U11202 (N_11202,N_4607,N_2868);
and U11203 (N_11203,N_3310,N_4312);
nand U11204 (N_11204,N_2348,N_1654);
and U11205 (N_11205,N_5263,N_5206);
or U11206 (N_11206,N_1612,N_2923);
or U11207 (N_11207,N_5669,N_5706);
and U11208 (N_11208,N_3350,N_5149);
xnor U11209 (N_11209,N_686,N_752);
or U11210 (N_11210,N_5485,N_2817);
xor U11211 (N_11211,N_3589,N_3997);
xnor U11212 (N_11212,N_3319,N_5748);
or U11213 (N_11213,N_5006,N_1039);
nand U11214 (N_11214,N_3354,N_3718);
or U11215 (N_11215,N_2956,N_3073);
and U11216 (N_11216,N_5238,N_801);
xor U11217 (N_11217,N_1627,N_2586);
and U11218 (N_11218,N_5977,N_452);
xor U11219 (N_11219,N_5984,N_981);
xor U11220 (N_11220,N_2507,N_4107);
or U11221 (N_11221,N_2145,N_4875);
nand U11222 (N_11222,N_2400,N_4693);
and U11223 (N_11223,N_2284,N_1485);
or U11224 (N_11224,N_4304,N_458);
or U11225 (N_11225,N_454,N_4111);
nor U11226 (N_11226,N_1690,N_5169);
nor U11227 (N_11227,N_2219,N_149);
nor U11228 (N_11228,N_5267,N_5876);
nor U11229 (N_11229,N_1634,N_3073);
or U11230 (N_11230,N_1481,N_3179);
nand U11231 (N_11231,N_4233,N_3341);
nand U11232 (N_11232,N_3281,N_798);
nor U11233 (N_11233,N_5509,N_5854);
nand U11234 (N_11234,N_3551,N_1156);
nor U11235 (N_11235,N_465,N_3328);
nor U11236 (N_11236,N_1273,N_982);
xnor U11237 (N_11237,N_2390,N_5227);
nor U11238 (N_11238,N_4685,N_4528);
or U11239 (N_11239,N_3933,N_2115);
nand U11240 (N_11240,N_5544,N_3685);
and U11241 (N_11241,N_3054,N_3512);
and U11242 (N_11242,N_4565,N_3056);
or U11243 (N_11243,N_1179,N_3649);
nand U11244 (N_11244,N_223,N_505);
nor U11245 (N_11245,N_4001,N_1937);
xor U11246 (N_11246,N_2304,N_1566);
xor U11247 (N_11247,N_2413,N_2439);
nand U11248 (N_11248,N_5943,N_4632);
nor U11249 (N_11249,N_2977,N_4412);
or U11250 (N_11250,N_2131,N_1688);
xor U11251 (N_11251,N_966,N_94);
and U11252 (N_11252,N_998,N_1600);
and U11253 (N_11253,N_3061,N_1310);
nand U11254 (N_11254,N_3251,N_5923);
or U11255 (N_11255,N_1196,N_3930);
nor U11256 (N_11256,N_4031,N_5996);
xor U11257 (N_11257,N_3463,N_4684);
nor U11258 (N_11258,N_2929,N_2350);
and U11259 (N_11259,N_4633,N_2772);
nor U11260 (N_11260,N_22,N_3656);
xnor U11261 (N_11261,N_1617,N_987);
and U11262 (N_11262,N_2623,N_2265);
nand U11263 (N_11263,N_3849,N_37);
nor U11264 (N_11264,N_906,N_4964);
and U11265 (N_11265,N_5545,N_871);
and U11266 (N_11266,N_915,N_4628);
or U11267 (N_11267,N_1989,N_2746);
xnor U11268 (N_11268,N_3523,N_450);
or U11269 (N_11269,N_2837,N_5983);
xnor U11270 (N_11270,N_2599,N_700);
nand U11271 (N_11271,N_1953,N_1675);
nand U11272 (N_11272,N_5280,N_4268);
nor U11273 (N_11273,N_2970,N_5326);
and U11274 (N_11274,N_3278,N_3350);
or U11275 (N_11275,N_2704,N_2418);
or U11276 (N_11276,N_5262,N_5898);
or U11277 (N_11277,N_2025,N_5420);
and U11278 (N_11278,N_3346,N_4857);
or U11279 (N_11279,N_4914,N_3501);
nand U11280 (N_11280,N_300,N_4579);
or U11281 (N_11281,N_1256,N_1477);
xnor U11282 (N_11282,N_3773,N_1184);
xor U11283 (N_11283,N_5099,N_2399);
xor U11284 (N_11284,N_528,N_4141);
and U11285 (N_11285,N_2556,N_5655);
xor U11286 (N_11286,N_5990,N_4429);
or U11287 (N_11287,N_5697,N_2392);
nor U11288 (N_11288,N_3500,N_2227);
nor U11289 (N_11289,N_1471,N_5099);
or U11290 (N_11290,N_1534,N_1557);
nor U11291 (N_11291,N_1232,N_3352);
nand U11292 (N_11292,N_3740,N_359);
xnor U11293 (N_11293,N_4393,N_3422);
nor U11294 (N_11294,N_5907,N_3909);
nand U11295 (N_11295,N_929,N_1677);
and U11296 (N_11296,N_4707,N_1429);
nor U11297 (N_11297,N_4031,N_5830);
xnor U11298 (N_11298,N_3942,N_2648);
nand U11299 (N_11299,N_3417,N_3054);
and U11300 (N_11300,N_5548,N_2717);
and U11301 (N_11301,N_2155,N_2082);
or U11302 (N_11302,N_1081,N_521);
xor U11303 (N_11303,N_31,N_5232);
nor U11304 (N_11304,N_5695,N_2159);
nor U11305 (N_11305,N_1302,N_3176);
or U11306 (N_11306,N_1812,N_1156);
nor U11307 (N_11307,N_1616,N_5807);
nand U11308 (N_11308,N_5415,N_2130);
xor U11309 (N_11309,N_2064,N_5659);
xnor U11310 (N_11310,N_3211,N_4609);
nor U11311 (N_11311,N_3675,N_3287);
or U11312 (N_11312,N_1764,N_1934);
xnor U11313 (N_11313,N_5448,N_1619);
and U11314 (N_11314,N_5646,N_2041);
nand U11315 (N_11315,N_604,N_2115);
and U11316 (N_11316,N_339,N_1570);
nor U11317 (N_11317,N_4331,N_3065);
or U11318 (N_11318,N_5756,N_2286);
nand U11319 (N_11319,N_5961,N_3236);
or U11320 (N_11320,N_846,N_634);
xnor U11321 (N_11321,N_5794,N_4406);
nand U11322 (N_11322,N_1216,N_5440);
or U11323 (N_11323,N_2112,N_1518);
or U11324 (N_11324,N_5476,N_2912);
nor U11325 (N_11325,N_4980,N_5773);
or U11326 (N_11326,N_2741,N_2627);
and U11327 (N_11327,N_5032,N_1480);
xor U11328 (N_11328,N_3883,N_657);
nand U11329 (N_11329,N_4850,N_2009);
nand U11330 (N_11330,N_3781,N_3142);
nand U11331 (N_11331,N_3123,N_4493);
or U11332 (N_11332,N_4776,N_32);
and U11333 (N_11333,N_5175,N_2250);
xor U11334 (N_11334,N_4629,N_2378);
nor U11335 (N_11335,N_1844,N_1851);
nand U11336 (N_11336,N_5266,N_762);
or U11337 (N_11337,N_5172,N_76);
nand U11338 (N_11338,N_47,N_5675);
or U11339 (N_11339,N_3744,N_3395);
nand U11340 (N_11340,N_319,N_3117);
nor U11341 (N_11341,N_4698,N_1443);
or U11342 (N_11342,N_2451,N_3896);
or U11343 (N_11343,N_1803,N_3244);
and U11344 (N_11344,N_4576,N_1911);
and U11345 (N_11345,N_1446,N_2832);
nand U11346 (N_11346,N_2123,N_890);
or U11347 (N_11347,N_2087,N_2591);
nand U11348 (N_11348,N_2695,N_5053);
nand U11349 (N_11349,N_3356,N_461);
nor U11350 (N_11350,N_4500,N_3543);
or U11351 (N_11351,N_3973,N_2250);
nor U11352 (N_11352,N_1026,N_2355);
nand U11353 (N_11353,N_1065,N_1975);
xor U11354 (N_11354,N_5437,N_22);
xor U11355 (N_11355,N_5567,N_5478);
or U11356 (N_11356,N_3185,N_3268);
or U11357 (N_11357,N_5391,N_347);
xor U11358 (N_11358,N_5396,N_4473);
and U11359 (N_11359,N_3536,N_4927);
and U11360 (N_11360,N_2021,N_155);
nand U11361 (N_11361,N_614,N_554);
nand U11362 (N_11362,N_2945,N_984);
and U11363 (N_11363,N_4626,N_4751);
or U11364 (N_11364,N_5500,N_2546);
xnor U11365 (N_11365,N_73,N_2568);
or U11366 (N_11366,N_682,N_4363);
nand U11367 (N_11367,N_1623,N_5898);
nor U11368 (N_11368,N_5848,N_3316);
and U11369 (N_11369,N_5451,N_1163);
or U11370 (N_11370,N_1845,N_5993);
nor U11371 (N_11371,N_4656,N_99);
and U11372 (N_11372,N_3988,N_3650);
xor U11373 (N_11373,N_3932,N_1778);
nor U11374 (N_11374,N_5583,N_3668);
nand U11375 (N_11375,N_3442,N_4010);
nand U11376 (N_11376,N_3244,N_5499);
nand U11377 (N_11377,N_4136,N_5732);
and U11378 (N_11378,N_1724,N_1910);
and U11379 (N_11379,N_1855,N_4486);
xnor U11380 (N_11380,N_994,N_2072);
and U11381 (N_11381,N_255,N_3117);
or U11382 (N_11382,N_4383,N_224);
nor U11383 (N_11383,N_4628,N_1122);
xnor U11384 (N_11384,N_2173,N_4332);
and U11385 (N_11385,N_1175,N_88);
nor U11386 (N_11386,N_894,N_5493);
xnor U11387 (N_11387,N_2774,N_4900);
nand U11388 (N_11388,N_2159,N_1799);
nand U11389 (N_11389,N_4704,N_5984);
nand U11390 (N_11390,N_1940,N_1353);
xnor U11391 (N_11391,N_1242,N_4158);
and U11392 (N_11392,N_3752,N_5177);
or U11393 (N_11393,N_2539,N_5840);
or U11394 (N_11394,N_5806,N_1448);
xor U11395 (N_11395,N_1876,N_158);
xor U11396 (N_11396,N_4308,N_1535);
nand U11397 (N_11397,N_4907,N_5630);
nand U11398 (N_11398,N_3888,N_5767);
xor U11399 (N_11399,N_702,N_4230);
xnor U11400 (N_11400,N_4447,N_1129);
xnor U11401 (N_11401,N_1278,N_2111);
or U11402 (N_11402,N_2396,N_5134);
or U11403 (N_11403,N_2762,N_506);
and U11404 (N_11404,N_3077,N_1551);
xnor U11405 (N_11405,N_2683,N_89);
or U11406 (N_11406,N_5518,N_3123);
nand U11407 (N_11407,N_1433,N_3098);
xnor U11408 (N_11408,N_1033,N_942);
nor U11409 (N_11409,N_3215,N_2246);
nor U11410 (N_11410,N_968,N_3917);
or U11411 (N_11411,N_747,N_841);
or U11412 (N_11412,N_3136,N_4799);
nor U11413 (N_11413,N_1273,N_4768);
and U11414 (N_11414,N_36,N_5812);
nand U11415 (N_11415,N_4262,N_4354);
nand U11416 (N_11416,N_5100,N_2938);
or U11417 (N_11417,N_2760,N_3327);
or U11418 (N_11418,N_5345,N_43);
or U11419 (N_11419,N_4379,N_341);
and U11420 (N_11420,N_542,N_791);
nor U11421 (N_11421,N_4396,N_4999);
or U11422 (N_11422,N_3802,N_1204);
and U11423 (N_11423,N_5754,N_1732);
xor U11424 (N_11424,N_1802,N_3370);
xor U11425 (N_11425,N_2730,N_5177);
or U11426 (N_11426,N_3225,N_1039);
or U11427 (N_11427,N_3944,N_4497);
nor U11428 (N_11428,N_2549,N_3361);
nand U11429 (N_11429,N_3895,N_533);
nor U11430 (N_11430,N_2104,N_2097);
or U11431 (N_11431,N_5569,N_908);
nor U11432 (N_11432,N_4359,N_825);
and U11433 (N_11433,N_595,N_5715);
nand U11434 (N_11434,N_3937,N_4683);
xnor U11435 (N_11435,N_3396,N_2484);
nor U11436 (N_11436,N_5542,N_5995);
nand U11437 (N_11437,N_3985,N_762);
nand U11438 (N_11438,N_2784,N_3353);
xor U11439 (N_11439,N_1101,N_1788);
or U11440 (N_11440,N_5220,N_727);
nand U11441 (N_11441,N_2741,N_1771);
xor U11442 (N_11442,N_3208,N_1039);
xor U11443 (N_11443,N_1699,N_5587);
and U11444 (N_11444,N_1073,N_2714);
nand U11445 (N_11445,N_2654,N_2598);
nor U11446 (N_11446,N_975,N_4618);
and U11447 (N_11447,N_1212,N_240);
xnor U11448 (N_11448,N_4884,N_3336);
nor U11449 (N_11449,N_765,N_4410);
xor U11450 (N_11450,N_4131,N_1027);
xnor U11451 (N_11451,N_3659,N_222);
nor U11452 (N_11452,N_2,N_281);
or U11453 (N_11453,N_1452,N_4610);
nor U11454 (N_11454,N_1086,N_5075);
nor U11455 (N_11455,N_5816,N_1692);
or U11456 (N_11456,N_5906,N_114);
and U11457 (N_11457,N_3904,N_3259);
nand U11458 (N_11458,N_4459,N_4600);
xor U11459 (N_11459,N_5686,N_4471);
and U11460 (N_11460,N_4228,N_2674);
xor U11461 (N_11461,N_4732,N_3600);
and U11462 (N_11462,N_4580,N_944);
or U11463 (N_11463,N_4888,N_2838);
xor U11464 (N_11464,N_2326,N_639);
and U11465 (N_11465,N_1614,N_5625);
or U11466 (N_11466,N_5760,N_5508);
and U11467 (N_11467,N_3718,N_4679);
nand U11468 (N_11468,N_240,N_4509);
and U11469 (N_11469,N_677,N_1440);
or U11470 (N_11470,N_3147,N_3251);
or U11471 (N_11471,N_755,N_5641);
xnor U11472 (N_11472,N_4538,N_5252);
and U11473 (N_11473,N_187,N_4365);
or U11474 (N_11474,N_1629,N_3978);
and U11475 (N_11475,N_3469,N_3614);
and U11476 (N_11476,N_2244,N_286);
nand U11477 (N_11477,N_1493,N_4115);
or U11478 (N_11478,N_4569,N_1826);
nand U11479 (N_11479,N_4817,N_3342);
or U11480 (N_11480,N_4729,N_4512);
and U11481 (N_11481,N_3358,N_5455);
xnor U11482 (N_11482,N_4007,N_4967);
xnor U11483 (N_11483,N_4701,N_5915);
and U11484 (N_11484,N_3398,N_680);
xor U11485 (N_11485,N_2407,N_383);
and U11486 (N_11486,N_4326,N_3520);
xor U11487 (N_11487,N_1635,N_5158);
or U11488 (N_11488,N_793,N_2520);
nand U11489 (N_11489,N_4389,N_4230);
nand U11490 (N_11490,N_4489,N_1284);
nor U11491 (N_11491,N_1394,N_3136);
nor U11492 (N_11492,N_3174,N_5053);
or U11493 (N_11493,N_2095,N_386);
or U11494 (N_11494,N_2478,N_5704);
and U11495 (N_11495,N_646,N_760);
or U11496 (N_11496,N_3905,N_5279);
nand U11497 (N_11497,N_5172,N_1434);
or U11498 (N_11498,N_1240,N_3004);
or U11499 (N_11499,N_3300,N_789);
xnor U11500 (N_11500,N_5763,N_1367);
or U11501 (N_11501,N_2066,N_4409);
xnor U11502 (N_11502,N_4967,N_3298);
and U11503 (N_11503,N_508,N_1083);
xor U11504 (N_11504,N_5509,N_2557);
nor U11505 (N_11505,N_84,N_1535);
nor U11506 (N_11506,N_1130,N_4128);
nand U11507 (N_11507,N_4811,N_3977);
nand U11508 (N_11508,N_5209,N_2587);
or U11509 (N_11509,N_4065,N_4689);
and U11510 (N_11510,N_2498,N_2367);
nor U11511 (N_11511,N_1318,N_2281);
nand U11512 (N_11512,N_4609,N_2865);
xnor U11513 (N_11513,N_1408,N_1465);
xnor U11514 (N_11514,N_1349,N_2982);
nand U11515 (N_11515,N_3314,N_2520);
or U11516 (N_11516,N_5094,N_3800);
and U11517 (N_11517,N_2075,N_5668);
or U11518 (N_11518,N_1142,N_838);
or U11519 (N_11519,N_4114,N_4054);
nor U11520 (N_11520,N_4281,N_5830);
nor U11521 (N_11521,N_3221,N_4967);
nand U11522 (N_11522,N_3922,N_2771);
xnor U11523 (N_11523,N_1159,N_703);
xor U11524 (N_11524,N_5613,N_3735);
xnor U11525 (N_11525,N_1339,N_1506);
xnor U11526 (N_11526,N_5395,N_1128);
and U11527 (N_11527,N_2250,N_3997);
and U11528 (N_11528,N_3316,N_4297);
nor U11529 (N_11529,N_4417,N_2128);
xor U11530 (N_11530,N_3804,N_5573);
xor U11531 (N_11531,N_3037,N_4695);
and U11532 (N_11532,N_1012,N_379);
nor U11533 (N_11533,N_3069,N_904);
nand U11534 (N_11534,N_4652,N_3761);
nand U11535 (N_11535,N_3508,N_3964);
xnor U11536 (N_11536,N_2210,N_1410);
or U11537 (N_11537,N_3288,N_1617);
nand U11538 (N_11538,N_5199,N_5892);
and U11539 (N_11539,N_3311,N_400);
or U11540 (N_11540,N_4631,N_430);
xor U11541 (N_11541,N_4214,N_169);
and U11542 (N_11542,N_5523,N_2297);
xnor U11543 (N_11543,N_374,N_1739);
nand U11544 (N_11544,N_4842,N_2325);
nand U11545 (N_11545,N_3744,N_4045);
nor U11546 (N_11546,N_4393,N_527);
nor U11547 (N_11547,N_5205,N_216);
or U11548 (N_11548,N_4237,N_4838);
nand U11549 (N_11549,N_5416,N_4025);
nor U11550 (N_11550,N_3096,N_1169);
xor U11551 (N_11551,N_2405,N_3175);
or U11552 (N_11552,N_1693,N_3025);
nand U11553 (N_11553,N_5468,N_5126);
xor U11554 (N_11554,N_3323,N_4706);
or U11555 (N_11555,N_2686,N_4857);
nand U11556 (N_11556,N_2548,N_1290);
or U11557 (N_11557,N_2066,N_2655);
and U11558 (N_11558,N_3235,N_3383);
nor U11559 (N_11559,N_4280,N_1514);
and U11560 (N_11560,N_3623,N_910);
xnor U11561 (N_11561,N_1617,N_4977);
nand U11562 (N_11562,N_939,N_4773);
nand U11563 (N_11563,N_5773,N_4513);
or U11564 (N_11564,N_4199,N_5334);
nor U11565 (N_11565,N_816,N_2811);
nand U11566 (N_11566,N_4080,N_4990);
or U11567 (N_11567,N_567,N_5929);
nor U11568 (N_11568,N_288,N_1985);
or U11569 (N_11569,N_1181,N_3217);
or U11570 (N_11570,N_1864,N_1708);
or U11571 (N_11571,N_4414,N_2578);
or U11572 (N_11572,N_3886,N_1003);
and U11573 (N_11573,N_859,N_5);
nor U11574 (N_11574,N_788,N_4760);
and U11575 (N_11575,N_4854,N_4297);
or U11576 (N_11576,N_480,N_4824);
xor U11577 (N_11577,N_3365,N_4672);
or U11578 (N_11578,N_180,N_2752);
and U11579 (N_11579,N_825,N_2268);
or U11580 (N_11580,N_1657,N_3176);
nor U11581 (N_11581,N_5869,N_329);
nor U11582 (N_11582,N_1549,N_1220);
and U11583 (N_11583,N_3455,N_3491);
nor U11584 (N_11584,N_3087,N_3672);
and U11585 (N_11585,N_1185,N_191);
xor U11586 (N_11586,N_3857,N_1277);
and U11587 (N_11587,N_4739,N_1055);
nor U11588 (N_11588,N_5076,N_4738);
nor U11589 (N_11589,N_1837,N_3190);
or U11590 (N_11590,N_2318,N_2274);
nand U11591 (N_11591,N_1388,N_1595);
and U11592 (N_11592,N_5074,N_3914);
xnor U11593 (N_11593,N_5844,N_3271);
and U11594 (N_11594,N_2711,N_4398);
nor U11595 (N_11595,N_3635,N_3162);
and U11596 (N_11596,N_3445,N_872);
nor U11597 (N_11597,N_5926,N_2058);
xor U11598 (N_11598,N_2674,N_3);
nand U11599 (N_11599,N_1526,N_560);
xnor U11600 (N_11600,N_252,N_2434);
xor U11601 (N_11601,N_2804,N_456);
nand U11602 (N_11602,N_4994,N_2377);
nor U11603 (N_11603,N_1798,N_2060);
nand U11604 (N_11604,N_1750,N_550);
xor U11605 (N_11605,N_5107,N_1912);
and U11606 (N_11606,N_178,N_4038);
or U11607 (N_11607,N_2251,N_5908);
nor U11608 (N_11608,N_208,N_4616);
xnor U11609 (N_11609,N_1033,N_4395);
nor U11610 (N_11610,N_2236,N_4885);
xnor U11611 (N_11611,N_3371,N_4592);
and U11612 (N_11612,N_4464,N_4326);
nand U11613 (N_11613,N_2881,N_4235);
nor U11614 (N_11614,N_424,N_4299);
and U11615 (N_11615,N_4855,N_1168);
or U11616 (N_11616,N_1664,N_2553);
xor U11617 (N_11617,N_5235,N_1652);
xnor U11618 (N_11618,N_3427,N_1262);
xor U11619 (N_11619,N_4057,N_5843);
nand U11620 (N_11620,N_2801,N_2362);
nor U11621 (N_11621,N_1249,N_4909);
nor U11622 (N_11622,N_819,N_3761);
and U11623 (N_11623,N_1588,N_2155);
xor U11624 (N_11624,N_5310,N_5738);
nand U11625 (N_11625,N_3831,N_2822);
xnor U11626 (N_11626,N_5932,N_1466);
and U11627 (N_11627,N_4224,N_1538);
or U11628 (N_11628,N_4693,N_4899);
and U11629 (N_11629,N_39,N_1264);
or U11630 (N_11630,N_287,N_3428);
and U11631 (N_11631,N_1444,N_4052);
xnor U11632 (N_11632,N_4774,N_436);
nor U11633 (N_11633,N_5436,N_3054);
nor U11634 (N_11634,N_1446,N_2575);
nand U11635 (N_11635,N_5874,N_4051);
xnor U11636 (N_11636,N_4749,N_1057);
nor U11637 (N_11637,N_3103,N_4245);
nand U11638 (N_11638,N_3912,N_3659);
xor U11639 (N_11639,N_1191,N_4207);
or U11640 (N_11640,N_646,N_4632);
nand U11641 (N_11641,N_3189,N_314);
and U11642 (N_11642,N_959,N_2507);
or U11643 (N_11643,N_3692,N_2433);
nand U11644 (N_11644,N_1410,N_3695);
nand U11645 (N_11645,N_1665,N_3274);
xor U11646 (N_11646,N_1894,N_5467);
or U11647 (N_11647,N_3910,N_2087);
xor U11648 (N_11648,N_5807,N_3732);
or U11649 (N_11649,N_4462,N_5205);
or U11650 (N_11650,N_4519,N_5993);
nor U11651 (N_11651,N_5136,N_1487);
and U11652 (N_11652,N_5186,N_2558);
xor U11653 (N_11653,N_1302,N_1546);
and U11654 (N_11654,N_1722,N_2668);
nor U11655 (N_11655,N_1437,N_2283);
nand U11656 (N_11656,N_1092,N_5416);
and U11657 (N_11657,N_3781,N_1532);
and U11658 (N_11658,N_2421,N_4398);
or U11659 (N_11659,N_5360,N_3632);
nor U11660 (N_11660,N_1247,N_5318);
nand U11661 (N_11661,N_2387,N_2352);
nand U11662 (N_11662,N_1167,N_3643);
and U11663 (N_11663,N_3240,N_2498);
nand U11664 (N_11664,N_5494,N_2098);
or U11665 (N_11665,N_1365,N_5877);
xor U11666 (N_11666,N_2584,N_324);
xor U11667 (N_11667,N_680,N_5434);
nand U11668 (N_11668,N_353,N_2986);
nand U11669 (N_11669,N_2562,N_5404);
nor U11670 (N_11670,N_4391,N_5930);
and U11671 (N_11671,N_3573,N_4979);
nand U11672 (N_11672,N_3752,N_2577);
xnor U11673 (N_11673,N_4334,N_4218);
nor U11674 (N_11674,N_4730,N_3926);
or U11675 (N_11675,N_5995,N_5251);
or U11676 (N_11676,N_1992,N_976);
or U11677 (N_11677,N_1361,N_5059);
or U11678 (N_11678,N_1800,N_3798);
xor U11679 (N_11679,N_1939,N_5260);
or U11680 (N_11680,N_4064,N_4678);
and U11681 (N_11681,N_3141,N_442);
and U11682 (N_11682,N_152,N_3585);
nand U11683 (N_11683,N_2831,N_5034);
nor U11684 (N_11684,N_4961,N_5449);
and U11685 (N_11685,N_2069,N_913);
xnor U11686 (N_11686,N_5271,N_3389);
nand U11687 (N_11687,N_5944,N_3932);
or U11688 (N_11688,N_4791,N_3200);
or U11689 (N_11689,N_3344,N_231);
or U11690 (N_11690,N_4716,N_664);
and U11691 (N_11691,N_4958,N_1408);
nor U11692 (N_11692,N_2028,N_2761);
and U11693 (N_11693,N_2969,N_1730);
nand U11694 (N_11694,N_2990,N_5617);
and U11695 (N_11695,N_1797,N_3330);
and U11696 (N_11696,N_948,N_2455);
nor U11697 (N_11697,N_3598,N_106);
nor U11698 (N_11698,N_2260,N_828);
nand U11699 (N_11699,N_3205,N_5821);
or U11700 (N_11700,N_4349,N_5649);
or U11701 (N_11701,N_2671,N_199);
xnor U11702 (N_11702,N_2808,N_138);
xor U11703 (N_11703,N_687,N_3124);
and U11704 (N_11704,N_112,N_5481);
and U11705 (N_11705,N_230,N_4078);
xor U11706 (N_11706,N_5682,N_4789);
and U11707 (N_11707,N_2271,N_1640);
nand U11708 (N_11708,N_858,N_189);
and U11709 (N_11709,N_1020,N_2023);
nand U11710 (N_11710,N_437,N_2646);
nor U11711 (N_11711,N_569,N_2622);
xnor U11712 (N_11712,N_1342,N_512);
and U11713 (N_11713,N_2527,N_2240);
or U11714 (N_11714,N_1755,N_2431);
nand U11715 (N_11715,N_112,N_4917);
or U11716 (N_11716,N_5248,N_5866);
or U11717 (N_11717,N_2869,N_4275);
nand U11718 (N_11718,N_5727,N_1075);
nor U11719 (N_11719,N_1403,N_5058);
nor U11720 (N_11720,N_866,N_5077);
xor U11721 (N_11721,N_82,N_1742);
or U11722 (N_11722,N_2002,N_2663);
nor U11723 (N_11723,N_196,N_5244);
and U11724 (N_11724,N_4911,N_1876);
and U11725 (N_11725,N_4003,N_1774);
and U11726 (N_11726,N_2491,N_578);
xnor U11727 (N_11727,N_4317,N_2772);
and U11728 (N_11728,N_6,N_809);
or U11729 (N_11729,N_4117,N_5139);
nand U11730 (N_11730,N_3829,N_2317);
and U11731 (N_11731,N_984,N_5281);
nor U11732 (N_11732,N_1583,N_5346);
and U11733 (N_11733,N_1146,N_1534);
and U11734 (N_11734,N_3998,N_4565);
and U11735 (N_11735,N_3707,N_1422);
nor U11736 (N_11736,N_3943,N_3119);
nand U11737 (N_11737,N_2718,N_5711);
xnor U11738 (N_11738,N_4422,N_2896);
and U11739 (N_11739,N_984,N_5937);
xor U11740 (N_11740,N_3983,N_4248);
and U11741 (N_11741,N_185,N_5005);
nand U11742 (N_11742,N_2945,N_283);
xor U11743 (N_11743,N_522,N_5014);
xnor U11744 (N_11744,N_5311,N_1663);
nand U11745 (N_11745,N_5714,N_568);
nand U11746 (N_11746,N_3528,N_3261);
xor U11747 (N_11747,N_844,N_4401);
nor U11748 (N_11748,N_2664,N_2214);
nand U11749 (N_11749,N_5833,N_3672);
nand U11750 (N_11750,N_1055,N_3584);
nand U11751 (N_11751,N_2814,N_5512);
nand U11752 (N_11752,N_549,N_4863);
xnor U11753 (N_11753,N_2909,N_2147);
or U11754 (N_11754,N_1265,N_1409);
nand U11755 (N_11755,N_4792,N_4088);
nor U11756 (N_11756,N_1863,N_5251);
nand U11757 (N_11757,N_2057,N_3954);
and U11758 (N_11758,N_2275,N_3634);
nand U11759 (N_11759,N_2155,N_5459);
nand U11760 (N_11760,N_104,N_1136);
or U11761 (N_11761,N_3814,N_5363);
and U11762 (N_11762,N_555,N_116);
xor U11763 (N_11763,N_1538,N_1696);
xnor U11764 (N_11764,N_980,N_3867);
or U11765 (N_11765,N_4550,N_2157);
and U11766 (N_11766,N_4575,N_604);
nand U11767 (N_11767,N_4384,N_5482);
nand U11768 (N_11768,N_130,N_4127);
or U11769 (N_11769,N_4505,N_1782);
xor U11770 (N_11770,N_2502,N_2457);
and U11771 (N_11771,N_5860,N_1592);
nor U11772 (N_11772,N_5356,N_4006);
or U11773 (N_11773,N_5080,N_927);
and U11774 (N_11774,N_5366,N_1001);
nand U11775 (N_11775,N_3738,N_5129);
nor U11776 (N_11776,N_1780,N_2552);
xnor U11777 (N_11777,N_5962,N_2140);
nor U11778 (N_11778,N_1452,N_1866);
xnor U11779 (N_11779,N_4415,N_5436);
nand U11780 (N_11780,N_801,N_5770);
or U11781 (N_11781,N_410,N_4558);
nor U11782 (N_11782,N_4274,N_62);
xnor U11783 (N_11783,N_2353,N_251);
or U11784 (N_11784,N_1781,N_396);
nand U11785 (N_11785,N_1124,N_4926);
or U11786 (N_11786,N_5151,N_1119);
xor U11787 (N_11787,N_890,N_4013);
nand U11788 (N_11788,N_3911,N_4450);
nand U11789 (N_11789,N_5731,N_4603);
nor U11790 (N_11790,N_1930,N_4536);
or U11791 (N_11791,N_392,N_3657);
xnor U11792 (N_11792,N_776,N_3353);
nand U11793 (N_11793,N_2948,N_5365);
and U11794 (N_11794,N_3102,N_4987);
and U11795 (N_11795,N_3150,N_2452);
nor U11796 (N_11796,N_2428,N_5943);
or U11797 (N_11797,N_4094,N_1366);
or U11798 (N_11798,N_2089,N_3523);
and U11799 (N_11799,N_3401,N_764);
and U11800 (N_11800,N_1403,N_369);
nand U11801 (N_11801,N_4382,N_4568);
or U11802 (N_11802,N_3368,N_4014);
or U11803 (N_11803,N_4840,N_4536);
nand U11804 (N_11804,N_2509,N_1458);
xnor U11805 (N_11805,N_3597,N_647);
or U11806 (N_11806,N_602,N_4653);
or U11807 (N_11807,N_5633,N_4677);
xor U11808 (N_11808,N_1163,N_5864);
xor U11809 (N_11809,N_4221,N_3857);
nand U11810 (N_11810,N_476,N_2974);
xnor U11811 (N_11811,N_912,N_3536);
or U11812 (N_11812,N_1140,N_4060);
and U11813 (N_11813,N_23,N_1393);
or U11814 (N_11814,N_5430,N_3560);
and U11815 (N_11815,N_4872,N_5640);
or U11816 (N_11816,N_5493,N_4260);
and U11817 (N_11817,N_5295,N_3452);
xnor U11818 (N_11818,N_3239,N_5423);
and U11819 (N_11819,N_730,N_4825);
or U11820 (N_11820,N_4610,N_1123);
xnor U11821 (N_11821,N_4748,N_3608);
and U11822 (N_11822,N_4575,N_4370);
nand U11823 (N_11823,N_3806,N_780);
nor U11824 (N_11824,N_2967,N_5783);
nor U11825 (N_11825,N_2778,N_251);
or U11826 (N_11826,N_5005,N_5931);
xnor U11827 (N_11827,N_5930,N_1255);
nand U11828 (N_11828,N_2308,N_4485);
and U11829 (N_11829,N_870,N_1116);
and U11830 (N_11830,N_2852,N_156);
nand U11831 (N_11831,N_3518,N_4480);
or U11832 (N_11832,N_4929,N_4261);
nand U11833 (N_11833,N_3814,N_5268);
xor U11834 (N_11834,N_1792,N_3763);
nand U11835 (N_11835,N_4068,N_2607);
nor U11836 (N_11836,N_4945,N_1151);
xor U11837 (N_11837,N_3060,N_5453);
and U11838 (N_11838,N_158,N_5597);
or U11839 (N_11839,N_2317,N_1474);
nor U11840 (N_11840,N_13,N_701);
and U11841 (N_11841,N_3942,N_5764);
nor U11842 (N_11842,N_2871,N_505);
nor U11843 (N_11843,N_2596,N_4810);
and U11844 (N_11844,N_4939,N_857);
or U11845 (N_11845,N_3696,N_291);
nor U11846 (N_11846,N_267,N_750);
and U11847 (N_11847,N_3599,N_4490);
nor U11848 (N_11848,N_1508,N_4894);
and U11849 (N_11849,N_1956,N_3929);
nand U11850 (N_11850,N_171,N_5840);
nor U11851 (N_11851,N_4079,N_649);
xnor U11852 (N_11852,N_4089,N_4529);
and U11853 (N_11853,N_755,N_2053);
nor U11854 (N_11854,N_3113,N_542);
nand U11855 (N_11855,N_4087,N_1665);
nor U11856 (N_11856,N_2044,N_2140);
nor U11857 (N_11857,N_3849,N_182);
nor U11858 (N_11858,N_5424,N_2914);
nand U11859 (N_11859,N_5125,N_4921);
nand U11860 (N_11860,N_2567,N_4595);
and U11861 (N_11861,N_2189,N_1392);
or U11862 (N_11862,N_1064,N_3697);
or U11863 (N_11863,N_2250,N_686);
xnor U11864 (N_11864,N_900,N_5531);
nor U11865 (N_11865,N_466,N_4459);
nand U11866 (N_11866,N_3626,N_4628);
xor U11867 (N_11867,N_3519,N_5687);
xor U11868 (N_11868,N_5821,N_1701);
or U11869 (N_11869,N_1932,N_2523);
nor U11870 (N_11870,N_1794,N_4778);
nand U11871 (N_11871,N_2651,N_190);
or U11872 (N_11872,N_5736,N_564);
and U11873 (N_11873,N_1700,N_4824);
nor U11874 (N_11874,N_5057,N_822);
nand U11875 (N_11875,N_3320,N_5337);
nand U11876 (N_11876,N_3312,N_3095);
nor U11877 (N_11877,N_603,N_890);
xor U11878 (N_11878,N_3746,N_911);
or U11879 (N_11879,N_4965,N_5865);
nor U11880 (N_11880,N_5813,N_1444);
or U11881 (N_11881,N_3899,N_5425);
nand U11882 (N_11882,N_2337,N_4001);
and U11883 (N_11883,N_708,N_4487);
nor U11884 (N_11884,N_4971,N_1210);
nor U11885 (N_11885,N_42,N_2272);
nor U11886 (N_11886,N_3572,N_5784);
or U11887 (N_11887,N_1402,N_1595);
or U11888 (N_11888,N_4419,N_1601);
and U11889 (N_11889,N_4001,N_4930);
nand U11890 (N_11890,N_4157,N_5967);
nor U11891 (N_11891,N_4366,N_4557);
or U11892 (N_11892,N_2221,N_3525);
and U11893 (N_11893,N_997,N_4007);
or U11894 (N_11894,N_3207,N_1228);
nor U11895 (N_11895,N_1591,N_3689);
xor U11896 (N_11896,N_292,N_2049);
and U11897 (N_11897,N_238,N_4788);
and U11898 (N_11898,N_4073,N_5591);
xnor U11899 (N_11899,N_4431,N_3075);
and U11900 (N_11900,N_2822,N_2002);
or U11901 (N_11901,N_239,N_2659);
and U11902 (N_11902,N_2789,N_2818);
or U11903 (N_11903,N_5005,N_1523);
nand U11904 (N_11904,N_58,N_5173);
nand U11905 (N_11905,N_5002,N_4123);
nor U11906 (N_11906,N_999,N_5585);
xnor U11907 (N_11907,N_1826,N_4007);
or U11908 (N_11908,N_4854,N_3654);
nand U11909 (N_11909,N_5786,N_970);
nor U11910 (N_11910,N_2485,N_4461);
or U11911 (N_11911,N_3841,N_223);
nand U11912 (N_11912,N_4484,N_2984);
nand U11913 (N_11913,N_4726,N_3732);
and U11914 (N_11914,N_3651,N_4110);
or U11915 (N_11915,N_5477,N_4506);
or U11916 (N_11916,N_4915,N_1817);
xor U11917 (N_11917,N_1704,N_5347);
xnor U11918 (N_11918,N_3109,N_1546);
xnor U11919 (N_11919,N_1171,N_962);
xnor U11920 (N_11920,N_1854,N_2288);
nor U11921 (N_11921,N_4189,N_2893);
xor U11922 (N_11922,N_5374,N_355);
xor U11923 (N_11923,N_3372,N_89);
xor U11924 (N_11924,N_2643,N_2731);
nor U11925 (N_11925,N_3857,N_1364);
xor U11926 (N_11926,N_472,N_4562);
or U11927 (N_11927,N_411,N_2701);
or U11928 (N_11928,N_1129,N_1677);
xor U11929 (N_11929,N_5841,N_3845);
and U11930 (N_11930,N_4353,N_1251);
nor U11931 (N_11931,N_4137,N_3284);
and U11932 (N_11932,N_5422,N_3995);
nand U11933 (N_11933,N_31,N_3742);
xor U11934 (N_11934,N_1731,N_3656);
xnor U11935 (N_11935,N_4751,N_4995);
nor U11936 (N_11936,N_5401,N_3686);
and U11937 (N_11937,N_3142,N_310);
or U11938 (N_11938,N_1126,N_4992);
and U11939 (N_11939,N_2411,N_1349);
xor U11940 (N_11940,N_2454,N_104);
nand U11941 (N_11941,N_1627,N_1524);
or U11942 (N_11942,N_5968,N_4270);
and U11943 (N_11943,N_1089,N_5379);
nor U11944 (N_11944,N_5031,N_73);
and U11945 (N_11945,N_139,N_1605);
xnor U11946 (N_11946,N_777,N_5973);
nor U11947 (N_11947,N_1903,N_3469);
nor U11948 (N_11948,N_4181,N_3762);
nor U11949 (N_11949,N_4631,N_5098);
nor U11950 (N_11950,N_139,N_797);
or U11951 (N_11951,N_5157,N_3883);
or U11952 (N_11952,N_1387,N_3887);
xnor U11953 (N_11953,N_4683,N_5548);
or U11954 (N_11954,N_190,N_5686);
or U11955 (N_11955,N_365,N_3983);
and U11956 (N_11956,N_1328,N_1999);
or U11957 (N_11957,N_701,N_919);
and U11958 (N_11958,N_1481,N_2092);
or U11959 (N_11959,N_466,N_2327);
nor U11960 (N_11960,N_4600,N_784);
nor U11961 (N_11961,N_207,N_5983);
nand U11962 (N_11962,N_700,N_5401);
nor U11963 (N_11963,N_3744,N_5696);
or U11964 (N_11964,N_4153,N_5126);
nor U11965 (N_11965,N_1388,N_3883);
and U11966 (N_11966,N_3313,N_2733);
and U11967 (N_11967,N_1904,N_1809);
nand U11968 (N_11968,N_3014,N_165);
nand U11969 (N_11969,N_3167,N_289);
and U11970 (N_11970,N_3689,N_1041);
nand U11971 (N_11971,N_4661,N_2731);
and U11972 (N_11972,N_5541,N_4016);
nor U11973 (N_11973,N_4021,N_5359);
and U11974 (N_11974,N_5337,N_5024);
nor U11975 (N_11975,N_2417,N_3199);
and U11976 (N_11976,N_820,N_4843);
or U11977 (N_11977,N_3728,N_5699);
or U11978 (N_11978,N_3424,N_2737);
xnor U11979 (N_11979,N_3582,N_4190);
or U11980 (N_11980,N_540,N_5677);
nor U11981 (N_11981,N_2862,N_1600);
and U11982 (N_11982,N_5988,N_5676);
and U11983 (N_11983,N_775,N_5987);
xnor U11984 (N_11984,N_4550,N_3447);
nor U11985 (N_11985,N_3864,N_633);
nand U11986 (N_11986,N_1979,N_4082);
xor U11987 (N_11987,N_367,N_375);
xor U11988 (N_11988,N_2920,N_5981);
and U11989 (N_11989,N_2379,N_1157);
or U11990 (N_11990,N_5793,N_1782);
nor U11991 (N_11991,N_2452,N_5393);
nor U11992 (N_11992,N_5004,N_1735);
and U11993 (N_11993,N_5491,N_1336);
or U11994 (N_11994,N_4657,N_2175);
and U11995 (N_11995,N_4081,N_5979);
and U11996 (N_11996,N_5372,N_5297);
xnor U11997 (N_11997,N_940,N_3832);
and U11998 (N_11998,N_4928,N_2557);
nor U11999 (N_11999,N_1292,N_1334);
nand U12000 (N_12000,N_7919,N_8425);
nand U12001 (N_12001,N_9490,N_8306);
or U12002 (N_12002,N_7322,N_9093);
and U12003 (N_12003,N_7856,N_6477);
and U12004 (N_12004,N_8043,N_7518);
and U12005 (N_12005,N_7472,N_6496);
or U12006 (N_12006,N_8569,N_9341);
or U12007 (N_12007,N_11534,N_8935);
xnor U12008 (N_12008,N_6253,N_8252);
xor U12009 (N_12009,N_7481,N_9729);
nand U12010 (N_12010,N_7475,N_8205);
nand U12011 (N_12011,N_6019,N_9267);
nor U12012 (N_12012,N_6135,N_6879);
xnor U12013 (N_12013,N_11997,N_8866);
nand U12014 (N_12014,N_7609,N_8154);
or U12015 (N_12015,N_9582,N_11348);
and U12016 (N_12016,N_8641,N_9057);
or U12017 (N_12017,N_8948,N_11741);
nor U12018 (N_12018,N_8611,N_11602);
or U12019 (N_12019,N_7950,N_10019);
nor U12020 (N_12020,N_7975,N_6747);
and U12021 (N_12021,N_7151,N_10628);
or U12022 (N_12022,N_10625,N_10945);
and U12023 (N_12023,N_11736,N_7574);
and U12024 (N_12024,N_6616,N_11347);
nor U12025 (N_12025,N_10252,N_11965);
nor U12026 (N_12026,N_11287,N_8086);
nor U12027 (N_12027,N_9215,N_11100);
or U12028 (N_12028,N_9122,N_7109);
xor U12029 (N_12029,N_10388,N_9842);
and U12030 (N_12030,N_7144,N_10537);
and U12031 (N_12031,N_9749,N_11119);
or U12032 (N_12032,N_7153,N_7276);
or U12033 (N_12033,N_8942,N_6041);
or U12034 (N_12034,N_6183,N_10694);
nor U12035 (N_12035,N_6150,N_9029);
or U12036 (N_12036,N_11669,N_8818);
nor U12037 (N_12037,N_9562,N_11476);
or U12038 (N_12038,N_7218,N_11343);
xnor U12039 (N_12039,N_6736,N_7514);
nand U12040 (N_12040,N_11002,N_10636);
nor U12041 (N_12041,N_11521,N_11744);
or U12042 (N_12042,N_8858,N_9873);
xor U12043 (N_12043,N_11978,N_6503);
nand U12044 (N_12044,N_7311,N_9959);
and U12045 (N_12045,N_8962,N_11837);
nor U12046 (N_12046,N_9513,N_10235);
or U12047 (N_12047,N_10843,N_7460);
nand U12048 (N_12048,N_9089,N_10820);
nor U12049 (N_12049,N_9328,N_6394);
nand U12050 (N_12050,N_6449,N_6053);
nand U12051 (N_12051,N_9604,N_6087);
or U12052 (N_12052,N_6969,N_11330);
nor U12053 (N_12053,N_6110,N_8113);
or U12054 (N_12054,N_7331,N_10509);
nand U12055 (N_12055,N_8864,N_7516);
and U12056 (N_12056,N_6141,N_7171);
or U12057 (N_12057,N_8173,N_9630);
nor U12058 (N_12058,N_6954,N_10260);
nor U12059 (N_12059,N_7849,N_11331);
nor U12060 (N_12060,N_7913,N_11230);
and U12061 (N_12061,N_11597,N_11887);
or U12062 (N_12062,N_10651,N_7567);
nor U12063 (N_12063,N_10976,N_11758);
and U12064 (N_12064,N_9982,N_9367);
nor U12065 (N_12065,N_10370,N_7454);
xor U12066 (N_12066,N_9943,N_10285);
or U12067 (N_12067,N_10085,N_11326);
or U12068 (N_12068,N_10750,N_7360);
xnor U12069 (N_12069,N_6124,N_11339);
or U12070 (N_12070,N_8199,N_7077);
and U12071 (N_12071,N_7683,N_6781);
nor U12072 (N_12072,N_8365,N_11353);
nor U12073 (N_12073,N_7699,N_8591);
or U12074 (N_12074,N_8091,N_10481);
nand U12075 (N_12075,N_6923,N_10873);
nand U12076 (N_12076,N_11131,N_11462);
and U12077 (N_12077,N_6127,N_6578);
nand U12078 (N_12078,N_9395,N_6085);
and U12079 (N_12079,N_7924,N_6684);
xor U12080 (N_12080,N_10339,N_7253);
nor U12081 (N_12081,N_9740,N_8082);
and U12082 (N_12082,N_8501,N_11715);
nor U12083 (N_12083,N_9546,N_9659);
xor U12084 (N_12084,N_9411,N_11647);
nor U12085 (N_12085,N_10814,N_10077);
nor U12086 (N_12086,N_9866,N_10435);
or U12087 (N_12087,N_9793,N_10834);
or U12088 (N_12088,N_7983,N_7860);
nand U12089 (N_12089,N_8129,N_10101);
or U12090 (N_12090,N_7263,N_8369);
nand U12091 (N_12091,N_6900,N_8331);
or U12092 (N_12092,N_9098,N_9882);
and U12093 (N_12093,N_7623,N_9786);
and U12094 (N_12094,N_7798,N_6515);
nand U12095 (N_12095,N_11310,N_9741);
and U12096 (N_12096,N_11572,N_11478);
nand U12097 (N_12097,N_7309,N_7048);
and U12098 (N_12098,N_11248,N_10833);
nand U12099 (N_12099,N_9008,N_11018);
nand U12100 (N_12100,N_7018,N_8795);
or U12101 (N_12101,N_7359,N_9876);
nor U12102 (N_12102,N_10254,N_10661);
nor U12103 (N_12103,N_10718,N_10624);
and U12104 (N_12104,N_7176,N_6604);
xnor U12105 (N_12105,N_7193,N_11692);
xor U12106 (N_12106,N_9508,N_10355);
nor U12107 (N_12107,N_10057,N_8906);
nand U12108 (N_12108,N_6476,N_6484);
and U12109 (N_12109,N_9832,N_11070);
nand U12110 (N_12110,N_9248,N_11408);
or U12111 (N_12111,N_8761,N_8116);
nor U12112 (N_12112,N_8430,N_9885);
and U12113 (N_12113,N_7887,N_10804);
or U12114 (N_12114,N_10487,N_6162);
nor U12115 (N_12115,N_9902,N_7202);
xor U12116 (N_12116,N_7626,N_11678);
xnor U12117 (N_12117,N_10511,N_7869);
nand U12118 (N_12118,N_9129,N_10732);
nand U12119 (N_12119,N_9572,N_7282);
nor U12120 (N_12120,N_7380,N_11227);
xor U12121 (N_12121,N_7762,N_8808);
nand U12122 (N_12122,N_9196,N_10476);
nor U12123 (N_12123,N_11481,N_11432);
xnor U12124 (N_12124,N_8322,N_7734);
nor U12125 (N_12125,N_10070,N_10360);
and U12126 (N_12126,N_8260,N_8603);
and U12127 (N_12127,N_6103,N_7008);
nand U12128 (N_12128,N_10679,N_10379);
nand U12129 (N_12129,N_11969,N_8269);
xor U12130 (N_12130,N_8422,N_11667);
xnor U12131 (N_12131,N_8355,N_7458);
nand U12132 (N_12132,N_8427,N_9884);
and U12133 (N_12133,N_10570,N_11025);
nor U12134 (N_12134,N_7836,N_8338);
nor U12135 (N_12135,N_11846,N_10910);
xor U12136 (N_12136,N_9552,N_8056);
or U12137 (N_12137,N_6857,N_10192);
nor U12138 (N_12138,N_9431,N_10114);
and U12139 (N_12139,N_10176,N_8980);
nor U12140 (N_12140,N_7469,N_7003);
and U12141 (N_12141,N_7985,N_11603);
nand U12142 (N_12142,N_10632,N_10432);
nor U12143 (N_12143,N_9983,N_11288);
or U12144 (N_12144,N_9190,N_9219);
and U12145 (N_12145,N_6094,N_6935);
or U12146 (N_12146,N_10730,N_10686);
nor U12147 (N_12147,N_9990,N_11295);
nor U12148 (N_12148,N_7854,N_11553);
or U12149 (N_12149,N_8834,N_6222);
and U12150 (N_12150,N_8662,N_6952);
or U12151 (N_12151,N_6936,N_11249);
nor U12152 (N_12152,N_8149,N_10564);
and U12153 (N_12153,N_9357,N_8142);
nand U12154 (N_12154,N_10734,N_7411);
nor U12155 (N_12155,N_11033,N_6594);
nand U12156 (N_12156,N_7838,N_11868);
nor U12157 (N_12157,N_9951,N_11982);
xor U12158 (N_12158,N_9401,N_6082);
or U12159 (N_12159,N_10967,N_10451);
nand U12160 (N_12160,N_6215,N_8739);
or U12161 (N_12161,N_8747,N_8323);
nand U12162 (N_12162,N_8098,N_9266);
nor U12163 (N_12163,N_7535,N_8133);
nand U12164 (N_12164,N_11421,N_9626);
nor U12165 (N_12165,N_6149,N_6458);
xor U12166 (N_12166,N_6855,N_6509);
or U12167 (N_12167,N_8936,N_7900);
or U12168 (N_12168,N_10830,N_8595);
and U12169 (N_12169,N_6607,N_10773);
and U12170 (N_12170,N_9007,N_6847);
or U12171 (N_12171,N_8372,N_11694);
or U12172 (N_12172,N_11776,N_11086);
and U12173 (N_12173,N_10995,N_6014);
nor U12174 (N_12174,N_9948,N_11134);
nor U12175 (N_12175,N_7873,N_9409);
xnor U12176 (N_12176,N_8716,N_9949);
and U12177 (N_12177,N_7706,N_7367);
or U12178 (N_12178,N_7168,N_11121);
or U12179 (N_12179,N_7586,N_8623);
nand U12180 (N_12180,N_11925,N_9693);
xnor U12181 (N_12181,N_7560,N_7818);
and U12182 (N_12182,N_9090,N_7281);
nor U12183 (N_12183,N_8674,N_9026);
xor U12184 (N_12184,N_9775,N_6884);
nand U12185 (N_12185,N_8754,N_10117);
nand U12186 (N_12186,N_8105,N_6440);
xor U12187 (N_12187,N_11773,N_6171);
nand U12188 (N_12188,N_8725,N_10222);
nand U12189 (N_12189,N_6332,N_10095);
or U12190 (N_12190,N_11900,N_6310);
or U12191 (N_12191,N_10038,N_11458);
and U12192 (N_12192,N_9118,N_10884);
nor U12193 (N_12193,N_6567,N_7437);
nor U12194 (N_12194,N_11608,N_6520);
or U12195 (N_12195,N_7994,N_7657);
nand U12196 (N_12196,N_7233,N_7254);
and U12197 (N_12197,N_7786,N_6734);
and U12198 (N_12198,N_11621,N_7273);
xor U12199 (N_12199,N_8497,N_6888);
nand U12200 (N_12200,N_8757,N_7912);
or U12201 (N_12201,N_9897,N_9911);
xnor U12202 (N_12202,N_8245,N_9589);
nor U12203 (N_12203,N_7045,N_9049);
and U12204 (N_12204,N_7952,N_9108);
or U12205 (N_12205,N_7748,N_8524);
nor U12206 (N_12206,N_7494,N_7929);
nand U12207 (N_12207,N_7806,N_7346);
xor U12208 (N_12208,N_9414,N_7769);
nand U12209 (N_12209,N_6582,N_9590);
or U12210 (N_12210,N_9020,N_11931);
and U12211 (N_12211,N_7713,N_6179);
nand U12212 (N_12212,N_9788,N_10985);
nor U12213 (N_12213,N_11219,N_11162);
and U12214 (N_12214,N_8162,N_6910);
and U12215 (N_12215,N_9001,N_6480);
and U12216 (N_12216,N_6345,N_9473);
or U12217 (N_12217,N_8351,N_7513);
and U12218 (N_12218,N_7252,N_9650);
or U12219 (N_12219,N_10558,N_10157);
and U12220 (N_12220,N_11390,N_7552);
nor U12221 (N_12221,N_8687,N_9514);
nor U12222 (N_12222,N_11668,N_8261);
nor U12223 (N_12223,N_8981,N_8698);
and U12224 (N_12224,N_7100,N_6730);
and U12225 (N_12225,N_11581,N_8462);
and U12226 (N_12226,N_8258,N_11051);
and U12227 (N_12227,N_6610,N_6761);
xnor U12228 (N_12228,N_11161,N_11963);
and U12229 (N_12229,N_10179,N_10365);
xnor U12230 (N_12230,N_8114,N_8538);
nand U12231 (N_12231,N_7006,N_6333);
and U12232 (N_12232,N_8530,N_9170);
nand U12233 (N_12233,N_11163,N_10139);
nand U12234 (N_12234,N_11907,N_11964);
or U12235 (N_12235,N_6994,N_9868);
or U12236 (N_12236,N_11810,N_11735);
and U12237 (N_12237,N_10406,N_9726);
and U12238 (N_12238,N_7307,N_7194);
nand U12239 (N_12239,N_7878,N_9308);
and U12240 (N_12240,N_6280,N_8577);
nor U12241 (N_12241,N_11237,N_9442);
nor U12242 (N_12242,N_6868,N_7379);
and U12243 (N_12243,N_10714,N_8843);
nand U12244 (N_12244,N_7811,N_11065);
nand U12245 (N_12245,N_6628,N_10229);
and U12246 (N_12246,N_8943,N_10507);
and U12247 (N_12247,N_7079,N_8064);
nor U12248 (N_12248,N_6837,N_7789);
or U12249 (N_12249,N_7409,N_7728);
and U12250 (N_12250,N_11210,N_6360);
xor U12251 (N_12251,N_7729,N_10171);
xnor U12252 (N_12252,N_11664,N_6733);
xnor U12253 (N_12253,N_8104,N_11723);
or U12254 (N_12254,N_10323,N_6627);
and U12255 (N_12255,N_10950,N_7258);
nor U12256 (N_12256,N_8361,N_10215);
or U12257 (N_12257,N_6185,N_6010);
or U12258 (N_12258,N_9703,N_10554);
xor U12259 (N_12259,N_8379,N_6187);
xor U12260 (N_12260,N_8387,N_10751);
nor U12261 (N_12261,N_7092,N_6738);
and U12262 (N_12262,N_9912,N_11819);
nor U12263 (N_12263,N_7526,N_8450);
xor U12264 (N_12264,N_6791,N_8574);
or U12265 (N_12265,N_11165,N_6782);
or U12266 (N_12266,N_7232,N_6443);
and U12267 (N_12267,N_11616,N_11798);
nor U12268 (N_12268,N_10735,N_8014);
and U12269 (N_12269,N_10003,N_6676);
xnor U12270 (N_12270,N_11142,N_9751);
and U12271 (N_12271,N_9327,N_10190);
xor U12272 (N_12272,N_6334,N_9255);
nand U12273 (N_12273,N_10934,N_8771);
nor U12274 (N_12274,N_7754,N_10227);
nand U12275 (N_12275,N_10011,N_10327);
nor U12276 (N_12276,N_7700,N_11243);
nor U12277 (N_12277,N_6982,N_10069);
xnor U12278 (N_12278,N_6040,N_6959);
nand U12279 (N_12279,N_11254,N_7538);
or U12280 (N_12280,N_9715,N_8030);
nand U12281 (N_12281,N_8610,N_10068);
nand U12282 (N_12282,N_10450,N_11088);
nor U12283 (N_12283,N_10658,N_11683);
or U12284 (N_12284,N_8287,N_8176);
xnor U12285 (N_12285,N_10931,N_11081);
xnor U12286 (N_12286,N_11190,N_11494);
or U12287 (N_12287,N_7721,N_8328);
xnor U12288 (N_12288,N_11180,N_7392);
nor U12289 (N_12289,N_6309,N_11027);
nand U12290 (N_12290,N_8811,N_9692);
xor U12291 (N_12291,N_10051,N_10753);
nor U12292 (N_12292,N_6406,N_6227);
xor U12293 (N_12293,N_6177,N_9452);
nand U12294 (N_12294,N_9984,N_9771);
and U12295 (N_12295,N_7744,N_6897);
nor U12296 (N_12296,N_9437,N_7782);
and U12297 (N_12297,N_11628,N_10706);
or U12298 (N_12298,N_11674,N_8308);
xor U12299 (N_12299,N_6438,N_7047);
and U12300 (N_12300,N_9717,N_7189);
and U12301 (N_12301,N_8336,N_9689);
nor U12302 (N_12302,N_7801,N_8903);
or U12303 (N_12303,N_9286,N_11836);
nor U12304 (N_12304,N_11460,N_8778);
xnor U12305 (N_12305,N_10471,N_9469);
nor U12306 (N_12306,N_9000,N_8015);
or U12307 (N_12307,N_6835,N_8673);
and U12308 (N_12308,N_7260,N_8676);
xnor U12309 (N_12309,N_9879,N_11291);
nand U12310 (N_12310,N_8366,N_7658);
xor U12311 (N_12311,N_10698,N_9838);
xor U12312 (N_12312,N_10186,N_9321);
xor U12313 (N_12313,N_6107,N_11909);
nand U12314 (N_12314,N_11858,N_8349);
nor U12315 (N_12315,N_10899,N_6322);
or U12316 (N_12316,N_10258,N_8998);
and U12317 (N_12317,N_9175,N_9702);
nand U12318 (N_12318,N_11215,N_10486);
or U12319 (N_12319,N_6213,N_11457);
and U12320 (N_12320,N_8152,N_9737);
and U12321 (N_12321,N_6919,N_8931);
nor U12322 (N_12322,N_7397,N_7834);
nor U12323 (N_12323,N_9526,N_11748);
xor U12324 (N_12324,N_11133,N_7456);
or U12325 (N_12325,N_8634,N_8780);
nand U12326 (N_12326,N_11952,N_9045);
xor U12327 (N_12327,N_6037,N_8773);
nand U12328 (N_12328,N_10547,N_7280);
nand U12329 (N_12329,N_10249,N_9687);
nor U12330 (N_12330,N_11084,N_9533);
xnor U12331 (N_12331,N_10189,N_10639);
or U12332 (N_12332,N_7415,N_8491);
and U12333 (N_12333,N_7587,N_11985);
xor U12334 (N_12334,N_11654,N_6865);
and U12335 (N_12335,N_6690,N_11045);
nor U12336 (N_12336,N_9654,N_6170);
nand U12337 (N_12337,N_10840,N_8505);
nand U12338 (N_12338,N_8679,N_7137);
nor U12339 (N_12339,N_8658,N_6963);
nand U12340 (N_12340,N_11280,N_6203);
or U12341 (N_12341,N_11447,N_11713);
nor U12342 (N_12342,N_10489,N_7382);
xnor U12343 (N_12343,N_10480,N_9128);
and U12344 (N_12344,N_8590,N_11046);
or U12345 (N_12345,N_10294,N_9148);
or U12346 (N_12346,N_6875,N_6192);
nor U12347 (N_12347,N_6346,N_6816);
and U12348 (N_12348,N_9426,N_7921);
and U12349 (N_12349,N_9850,N_10932);
nor U12350 (N_12350,N_6387,N_8150);
xor U12351 (N_12351,N_8703,N_11399);
nor U12352 (N_12352,N_7443,N_11058);
xor U12353 (N_12353,N_10572,N_7743);
xnor U12354 (N_12354,N_8292,N_7669);
nand U12355 (N_12355,N_7827,N_6510);
nand U12356 (N_12356,N_8122,N_10377);
nand U12357 (N_12357,N_10277,N_7234);
nor U12358 (N_12358,N_10352,N_9714);
nor U12359 (N_12359,N_10597,N_10047);
nor U12360 (N_12360,N_8418,N_11261);
xor U12361 (N_12361,N_11580,N_10711);
nor U12362 (N_12362,N_8939,N_7134);
or U12363 (N_12363,N_9597,N_11918);
nand U12364 (N_12364,N_7491,N_7319);
and U12365 (N_12365,N_8976,N_8549);
or U12366 (N_12366,N_10453,N_10783);
nor U12367 (N_12367,N_6472,N_7991);
and U12368 (N_12368,N_8999,N_11951);
xor U12369 (N_12369,N_7654,N_11930);
nor U12370 (N_12370,N_10505,N_6099);
nand U12371 (N_12371,N_10600,N_8143);
xnor U12372 (N_12372,N_8347,N_9713);
nor U12373 (N_12373,N_8156,N_10150);
and U12374 (N_12374,N_11530,N_9011);
xor U12375 (N_12375,N_7088,N_8821);
or U12376 (N_12376,N_7547,N_11896);
nand U12377 (N_12377,N_6169,N_9887);
nor U12378 (N_12378,N_6494,N_9636);
or U12379 (N_12379,N_11558,N_7423);
nor U12380 (N_12380,N_7817,N_7131);
or U12381 (N_12381,N_9960,N_8183);
nor U12382 (N_12382,N_6519,N_11496);
xnor U12383 (N_12383,N_7870,N_7770);
nor U12384 (N_12384,N_6341,N_11844);
or U12385 (N_12385,N_6652,N_11706);
xor U12386 (N_12386,N_9928,N_9223);
or U12387 (N_12387,N_11720,N_6967);
and U12388 (N_12388,N_8300,N_9547);
and U12389 (N_12389,N_7156,N_11318);
or U12390 (N_12390,N_7237,N_11059);
or U12391 (N_12391,N_8360,N_11841);
or U12392 (N_12392,N_10064,N_7501);
nor U12393 (N_12393,N_6680,N_8236);
nand U12394 (N_12394,N_8469,N_9795);
nand U12395 (N_12395,N_6822,N_9602);
or U12396 (N_12396,N_7235,N_6722);
or U12397 (N_12397,N_8263,N_7376);
nor U12398 (N_12398,N_11625,N_10579);
nor U12399 (N_12399,N_8562,N_7196);
or U12400 (N_12400,N_6725,N_6365);
nand U12401 (N_12401,N_8402,N_11737);
xor U12402 (N_12402,N_9283,N_8022);
xnor U12403 (N_12403,N_10279,N_9998);
nand U12404 (N_12404,N_6799,N_6410);
nor U12405 (N_12405,N_11413,N_10082);
nand U12406 (N_12406,N_11954,N_7776);
or U12407 (N_12407,N_6525,N_7433);
xor U12408 (N_12408,N_11252,N_6927);
nand U12409 (N_12409,N_10845,N_10670);
and U12410 (N_12410,N_8225,N_11937);
nand U12411 (N_12411,N_11173,N_11426);
xor U12412 (N_12412,N_7705,N_11157);
nand U12413 (N_12413,N_6375,N_8836);
xnor U12414 (N_12414,N_9688,N_6491);
nor U12415 (N_12415,N_10387,N_11835);
nor U12416 (N_12416,N_11302,N_9801);
nor U12417 (N_12417,N_9432,N_9829);
xor U12418 (N_12418,N_10994,N_7594);
or U12419 (N_12419,N_9083,N_7444);
nor U12420 (N_12420,N_11415,N_9553);
and U12421 (N_12421,N_11140,N_6386);
and U12422 (N_12422,N_10862,N_10116);
nor U12423 (N_12423,N_6599,N_8324);
nand U12424 (N_12424,N_6444,N_9097);
and U12425 (N_12425,N_6841,N_8649);
and U12426 (N_12426,N_11443,N_8612);
or U12427 (N_12427,N_7546,N_7681);
or U12428 (N_12428,N_10074,N_10292);
nand U12429 (N_12429,N_6549,N_9593);
xor U12430 (N_12430,N_6818,N_8576);
or U12431 (N_12431,N_7822,N_10589);
and U12432 (N_12432,N_11223,N_10635);
nand U12433 (N_12433,N_9558,N_8659);
and U12434 (N_12434,N_6361,N_9407);
xnor U12435 (N_12435,N_6313,N_10781);
xor U12436 (N_12436,N_10402,N_8353);
nor U12437 (N_12437,N_7796,N_7661);
or U12438 (N_12438,N_10497,N_10087);
nand U12439 (N_12439,N_6682,N_7531);
nand U12440 (N_12440,N_6479,N_6949);
xor U12441 (N_12441,N_6415,N_9149);
nand U12442 (N_12442,N_10519,N_11681);
or U12443 (N_12443,N_8776,N_10244);
and U12444 (N_12444,N_11203,N_11587);
or U12445 (N_12445,N_11196,N_8290);
xor U12446 (N_12446,N_6259,N_11916);
or U12447 (N_12447,N_9560,N_10996);
or U12448 (N_12448,N_9588,N_7327);
and U12449 (N_12449,N_7373,N_8449);
or U12450 (N_12450,N_7441,N_11751);
nor U12451 (N_12451,N_10680,N_9133);
and U12452 (N_12452,N_8782,N_8415);
nor U12453 (N_12453,N_7422,N_8218);
and U12454 (N_12454,N_7357,N_10330);
or U12455 (N_12455,N_7909,N_7390);
or U12456 (N_12456,N_11239,N_7752);
and U12457 (N_12457,N_9101,N_8699);
or U12458 (N_12458,N_7603,N_7606);
xor U12459 (N_12459,N_11260,N_9835);
and U12460 (N_12460,N_6843,N_6231);
nor U12461 (N_12461,N_11361,N_7333);
and U12462 (N_12462,N_8012,N_11220);
and U12463 (N_12463,N_10307,N_9387);
nand U12464 (N_12464,N_10728,N_8629);
nand U12465 (N_12465,N_11834,N_11630);
nand U12466 (N_12466,N_8672,N_10304);
nand U12467 (N_12467,N_10447,N_10322);
xor U12468 (N_12468,N_10801,N_9712);
and U12469 (N_12469,N_7001,N_7148);
and U12470 (N_12470,N_11060,N_9581);
or U12471 (N_12471,N_6252,N_6401);
nor U12472 (N_12472,N_6060,N_8410);
or U12473 (N_12473,N_7034,N_10765);
nor U12474 (N_12474,N_8046,N_6506);
and U12475 (N_12475,N_6299,N_9371);
and U12476 (N_12476,N_9260,N_11623);
and U12477 (N_12477,N_9601,N_7691);
or U12478 (N_12478,N_8206,N_11975);
or U12479 (N_12479,N_11933,N_7453);
nor U12480 (N_12480,N_11434,N_9673);
xnor U12481 (N_12481,N_10147,N_6077);
xor U12482 (N_12482,N_8504,N_6005);
nand U12483 (N_12483,N_8651,N_11812);
nand U12484 (N_12484,N_9814,N_6021);
or U12485 (N_12485,N_6988,N_8915);
nor U12486 (N_12486,N_10948,N_8058);
and U12487 (N_12487,N_11908,N_11075);
nor U12488 (N_12488,N_11409,N_9018);
nand U12489 (N_12489,N_9694,N_8277);
xnor U12490 (N_12490,N_10065,N_6079);
or U12491 (N_12491,N_8832,N_7846);
and U12492 (N_12492,N_11842,N_7462);
xnor U12493 (N_12493,N_11449,N_11860);
nand U12494 (N_12494,N_11831,N_6554);
or U12495 (N_12495,N_11657,N_11961);
or U12496 (N_12496,N_9381,N_10230);
and U12497 (N_12497,N_7356,N_11405);
xnor U12498 (N_12498,N_11772,N_6300);
xnor U12499 (N_12499,N_10060,N_10002);
or U12500 (N_12500,N_11263,N_7350);
and U12501 (N_12501,N_6330,N_7255);
nor U12502 (N_12502,N_9439,N_7667);
and U12503 (N_12503,N_6814,N_10593);
or U12504 (N_12504,N_11800,N_6538);
or U12505 (N_12505,N_9246,N_6100);
nor U12506 (N_12506,N_11346,N_8837);
nor U12507 (N_12507,N_9807,N_11801);
xnor U12508 (N_12508,N_8485,N_8002);
and U12509 (N_12509,N_11639,N_7668);
nand U12510 (N_12510,N_8933,N_6880);
or U12511 (N_12511,N_7876,N_9950);
and U12512 (N_12512,N_7338,N_8131);
or U12513 (N_12513,N_9969,N_8025);
xnor U12514 (N_12514,N_8424,N_9259);
nand U12515 (N_12515,N_10477,N_7108);
or U12516 (N_12516,N_10484,N_7297);
or U12517 (N_12517,N_8991,N_9355);
or U12518 (N_12518,N_7779,N_11889);
nand U12519 (N_12519,N_8033,N_6180);
nand U12520 (N_12520,N_7624,N_9235);
xnor U12521 (N_12521,N_7763,N_8708);
xor U12522 (N_12522,N_11850,N_11696);
nand U12523 (N_12523,N_8667,N_9450);
nand U12524 (N_12524,N_9753,N_9221);
and U12525 (N_12525,N_6468,N_11710);
xnor U12526 (N_12526,N_6109,N_10668);
and U12527 (N_12527,N_6901,N_11679);
nand U12528 (N_12528,N_7716,N_8481);
and U12529 (N_12529,N_6144,N_10076);
or U12530 (N_12530,N_6980,N_6251);
and U12531 (N_12531,N_8758,N_11769);
nand U12532 (N_12532,N_8625,N_11999);
and U12533 (N_12533,N_10241,N_9198);
or U12534 (N_12534,N_9464,N_8850);
or U12535 (N_12535,N_8346,N_6874);
and U12536 (N_12536,N_6987,N_8638);
xnor U12537 (N_12537,N_10425,N_10006);
or U12538 (N_12538,N_11382,N_8974);
or U12539 (N_12539,N_6036,N_9537);
nor U12540 (N_12540,N_9394,N_11726);
xor U12541 (N_12541,N_10348,N_8010);
and U12542 (N_12542,N_8271,N_9857);
xnor U12543 (N_12543,N_11212,N_10867);
and U12544 (N_12544,N_6753,N_8249);
nand U12545 (N_12545,N_9927,N_8342);
nand U12546 (N_12546,N_11077,N_6618);
xnor U12547 (N_12547,N_10905,N_11672);
xor U12548 (N_12548,N_10568,N_10269);
xnor U12549 (N_12549,N_11301,N_7484);
and U12550 (N_12550,N_9979,N_10708);
nor U12551 (N_12551,N_7662,N_11096);
and U12552 (N_12552,N_7505,N_10384);
nor U12553 (N_12553,N_7485,N_7941);
nand U12554 (N_12554,N_8362,N_9292);
and U12555 (N_12555,N_7352,N_6829);
xor U12556 (N_12556,N_8140,N_8877);
nand U12557 (N_12557,N_11360,N_8777);
and U12558 (N_12558,N_11821,N_6199);
or U12559 (N_12559,N_7911,N_10913);
nor U12560 (N_12560,N_7726,N_11765);
or U12561 (N_12561,N_7625,N_7601);
nor U12562 (N_12562,N_9145,N_9318);
nand U12563 (N_12563,N_9178,N_8040);
nand U12564 (N_12564,N_10705,N_10059);
xnor U12565 (N_12565,N_9172,N_7496);
and U12566 (N_12566,N_9095,N_8912);
or U12567 (N_12567,N_6216,N_8146);
nor U12568 (N_12568,N_9757,N_8557);
or U12569 (N_12569,N_10791,N_6145);
xnor U12570 (N_12570,N_6016,N_7886);
and U12571 (N_12571,N_8700,N_10007);
nor U12572 (N_12572,N_10397,N_9368);
xnor U12573 (N_12573,N_7335,N_6075);
or U12574 (N_12574,N_6964,N_10697);
xor U12575 (N_12575,N_10922,N_9577);
nand U12576 (N_12576,N_8161,N_11281);
or U12577 (N_12577,N_10858,N_8069);
and U12578 (N_12578,N_11130,N_10214);
xnor U12579 (N_12579,N_7427,N_6342);
nor U12580 (N_12580,N_8134,N_6836);
xor U12581 (N_12581,N_6941,N_9212);
or U12582 (N_12582,N_9287,N_6518);
nor U12583 (N_12583,N_8070,N_9611);
and U12584 (N_12584,N_6122,N_10496);
or U12585 (N_12585,N_8350,N_9282);
or U12586 (N_12586,N_6088,N_7998);
xnor U12587 (N_12587,N_7759,N_7577);
or U12588 (N_12588,N_10464,N_8412);
xor U12589 (N_12589,N_11004,N_11319);
nor U12590 (N_12590,N_7094,N_10829);
nand U12591 (N_12591,N_6777,N_9400);
and U12592 (N_12592,N_10374,N_10461);
or U12593 (N_12593,N_7965,N_8594);
or U12594 (N_12594,N_8726,N_6929);
xnor U12595 (N_12595,N_8856,N_7421);
nand U12596 (N_12596,N_7162,N_9510);
nand U12597 (N_12597,N_8175,N_8447);
nand U12598 (N_12598,N_10523,N_7621);
nor U12599 (N_12599,N_10436,N_10309);
nand U12600 (N_12600,N_8184,N_8454);
nor U12601 (N_12601,N_6225,N_6686);
xnor U12602 (N_12602,N_7095,N_8859);
or U12603 (N_12603,N_7561,N_6920);
nor U12604 (N_12604,N_10018,N_10604);
xor U12605 (N_12605,N_10120,N_8413);
or U12606 (N_12606,N_8309,N_6431);
nand U12607 (N_12607,N_6242,N_6452);
nor U12608 (N_12608,N_6625,N_11093);
and U12609 (N_12609,N_6381,N_6832);
xor U12610 (N_12610,N_10278,N_8313);
nor U12611 (N_12611,N_6962,N_11642);
and U12612 (N_12612,N_11606,N_9970);
or U12613 (N_12613,N_6266,N_6751);
xnor U12614 (N_12614,N_10337,N_10417);
nand U12615 (N_12615,N_9686,N_8171);
and U12616 (N_12616,N_10467,N_10818);
nor U12617 (N_12617,N_7940,N_8814);
and U12618 (N_12618,N_6072,N_6678);
or U12619 (N_12619,N_9862,N_11467);
or U12620 (N_12620,N_6808,N_8390);
xor U12621 (N_12621,N_7733,N_9030);
and U12622 (N_12622,N_9307,N_6850);
or U12623 (N_12623,N_7875,N_6647);
nand U12624 (N_12624,N_9051,N_6514);
nor U12625 (N_12625,N_6527,N_11818);
nor U12626 (N_12626,N_6671,N_10495);
or U12627 (N_12627,N_7591,N_11924);
and U12628 (N_12628,N_11151,N_10124);
and U12629 (N_12629,N_9529,N_7987);
or U12630 (N_12630,N_11238,N_6609);
or U12631 (N_12631,N_9515,N_8124);
nor U12632 (N_12632,N_7839,N_7330);
and U12633 (N_12633,N_8262,N_9704);
nor U12634 (N_12634,N_7989,N_11505);
or U12635 (N_12635,N_7678,N_6111);
nor U12636 (N_12636,N_11973,N_7031);
or U12637 (N_12637,N_7042,N_11218);
xnor U12638 (N_12638,N_7302,N_7523);
xor U12639 (N_12639,N_11517,N_9613);
or U12640 (N_12640,N_10565,N_7946);
or U12641 (N_12641,N_6172,N_8861);
and U12642 (N_12642,N_9099,N_10674);
nor U12643 (N_12643,N_11791,N_10357);
or U12644 (N_12644,N_11804,N_8740);
nor U12645 (N_12645,N_8367,N_11636);
and U12646 (N_12646,N_7612,N_11338);
xor U12647 (N_12647,N_8074,N_6297);
and U12648 (N_12648,N_11032,N_9016);
or U12649 (N_12649,N_8096,N_9670);
and U12650 (N_12650,N_8755,N_11928);
or U12651 (N_12651,N_7931,N_9388);
nor U12652 (N_12652,N_10975,N_11541);
nor U12653 (N_12653,N_6441,N_11807);
xor U12654 (N_12654,N_9985,N_10264);
or U12655 (N_12655,N_11983,N_7555);
and U12656 (N_12656,N_7541,N_9378);
and U12657 (N_12657,N_8655,N_11564);
or U12658 (N_12658,N_8585,N_7928);
nor U12659 (N_12659,N_10618,N_10122);
nand U12660 (N_12660,N_6117,N_10917);
and U12661 (N_12661,N_11479,N_8047);
xor U12662 (N_12662,N_7347,N_10266);
xnor U12663 (N_12663,N_7139,N_9893);
or U12664 (N_12664,N_6557,N_10305);
and U12665 (N_12665,N_8916,N_6459);
nand U12666 (N_12666,N_7324,N_11365);
and U12667 (N_12667,N_6785,N_11507);
or U12668 (N_12668,N_6696,N_7755);
or U12669 (N_12669,N_10382,N_11910);
and U12670 (N_12670,N_6221,N_7326);
nand U12671 (N_12671,N_7372,N_10557);
or U12672 (N_12672,N_8774,N_11991);
and U12673 (N_12673,N_9706,N_6337);
nand U12674 (N_12674,N_6767,N_6624);
and U12675 (N_12675,N_10131,N_6323);
nand U12676 (N_12676,N_9666,N_7121);
nor U12677 (N_12677,N_10919,N_10393);
xor U12678 (N_12678,N_8075,N_11095);
nor U12679 (N_12679,N_6655,N_8436);
nor U12680 (N_12680,N_10351,N_7771);
nand U12681 (N_12681,N_8445,N_8207);
xor U12682 (N_12682,N_7011,N_11158);
nand U12683 (N_12683,N_7054,N_6500);
or U12684 (N_12684,N_11650,N_7066);
or U12685 (N_12685,N_8586,N_6456);
and U12686 (N_12686,N_11396,N_11491);
nand U12687 (N_12687,N_9792,N_10616);
or U12688 (N_12688,N_6766,N_9312);
and U12689 (N_12689,N_9725,N_11446);
nand U12690 (N_12690,N_10739,N_6461);
and U12691 (N_12691,N_8849,N_6140);
and U12692 (N_12692,N_7502,N_11069);
and U12693 (N_12693,N_7685,N_10142);
or U12694 (N_12694,N_6121,N_10908);
nor U12695 (N_12695,N_6974,N_10363);
nand U12696 (N_12696,N_7483,N_6247);
and U12697 (N_12697,N_6973,N_8038);
nand U12698 (N_12698,N_9858,N_7476);
xor U12699 (N_12699,N_8049,N_11728);
or U12700 (N_12700,N_6432,N_11006);
and U12701 (N_12701,N_8835,N_7701);
xor U12702 (N_12702,N_10871,N_11946);
and U12703 (N_12703,N_6068,N_6511);
and U12704 (N_12704,N_6469,N_8296);
nor U12705 (N_12705,N_7385,N_11438);
nor U12706 (N_12706,N_10946,N_6388);
xor U12707 (N_12707,N_6434,N_6721);
nand U12708 (N_12708,N_7467,N_10944);
xor U12709 (N_12709,N_6702,N_7163);
xor U12710 (N_12710,N_9563,N_7648);
nand U12711 (N_12711,N_10361,N_10665);
nand U12712 (N_12712,N_6255,N_8657);
nand U12713 (N_12713,N_11972,N_8752);
and U12714 (N_12714,N_6552,N_6125);
nand U12715 (N_12715,N_11745,N_6258);
nor U12716 (N_12716,N_6304,N_11440);
and U12717 (N_12717,N_10979,N_6977);
nor U12718 (N_12718,N_10198,N_7203);
xnor U12719 (N_12719,N_6023,N_7060);
xor U12720 (N_12720,N_10457,N_8354);
nand U12721 (N_12721,N_11739,N_9534);
xnor U12722 (N_12722,N_11501,N_9931);
nand U12723 (N_12723,N_7303,N_6052);
nand U12724 (N_12724,N_7656,N_9036);
and U12725 (N_12725,N_9697,N_6915);
nand U12726 (N_12726,N_11487,N_6559);
nor U12727 (N_12727,N_10331,N_11247);
nand U12728 (N_12728,N_9640,N_11743);
nand U12729 (N_12729,N_6528,N_10503);
nor U12730 (N_12730,N_11510,N_8368);
and U12731 (N_12731,N_11734,N_6889);
or U12732 (N_12732,N_11293,N_10770);
nor U12733 (N_12733,N_9279,N_7226);
or U12734 (N_12734,N_6163,N_10924);
nand U12735 (N_12735,N_6285,N_11463);
nor U12736 (N_12736,N_11559,N_6435);
xnor U12737 (N_12737,N_7542,N_6523);
xor U12738 (N_12738,N_6279,N_6984);
nand U12739 (N_12739,N_11950,N_10306);
xor U12740 (N_12740,N_11883,N_8580);
nor U12741 (N_12741,N_7071,N_10468);
xnor U12742 (N_12742,N_10872,N_9232);
nor U12743 (N_12743,N_11369,N_9836);
nand U12744 (N_12744,N_7199,N_6807);
nor U12745 (N_12745,N_11523,N_8370);
and U12746 (N_12746,N_9682,N_9789);
nor U12747 (N_12747,N_11367,N_10418);
xnor U12748 (N_12748,N_6854,N_9494);
nand U12749 (N_12749,N_8601,N_7893);
nand U12750 (N_12750,N_10896,N_10390);
and U12751 (N_12751,N_6256,N_6467);
and U12752 (N_12752,N_11662,N_8515);
nand U12753 (N_12753,N_10338,N_9889);
xnor U12754 (N_12754,N_9299,N_8949);
and U12755 (N_12755,N_11483,N_10515);
xor U12756 (N_12756,N_10276,N_7917);
nor U12757 (N_12757,N_8552,N_7395);
and U12758 (N_12758,N_8461,N_6786);
nand U12759 (N_12759,N_6998,N_9362);
nand U12760 (N_12760,N_10280,N_9921);
or U12761 (N_12761,N_10000,N_9280);
xor U12762 (N_12762,N_11214,N_10110);
or U12763 (N_12763,N_9894,N_9073);
or U12764 (N_12764,N_10103,N_6278);
nor U12765 (N_12765,N_8111,N_7783);
or U12766 (N_12766,N_7463,N_7970);
xnor U12767 (N_12767,N_11213,N_10098);
and U12768 (N_12768,N_11160,N_11866);
xor U12769 (N_12769,N_7036,N_9453);
xor U12770 (N_12770,N_8181,N_11849);
and U12771 (N_12771,N_11884,N_8613);
nor U12772 (N_12772,N_6471,N_8317);
and U12773 (N_12773,N_7639,N_10385);
nor U12774 (N_12774,N_7178,N_10875);
xor U12775 (N_12775,N_11193,N_11940);
nor U12776 (N_12776,N_9973,N_9482);
or U12777 (N_12777,N_9479,N_10283);
or U12778 (N_12778,N_6735,N_6670);
xor U12779 (N_12779,N_9890,N_11493);
or U12780 (N_12780,N_9549,N_6315);
or U12781 (N_12781,N_11941,N_7445);
xor U12782 (N_12782,N_8624,N_7207);
xor U12783 (N_12783,N_10611,N_10137);
xnor U12784 (N_12784,N_8378,N_10815);
and U12785 (N_12785,N_9591,N_10013);
and U12786 (N_12786,N_9963,N_11698);
xnor U12787 (N_12787,N_10842,N_9609);
or U12788 (N_12788,N_11150,N_9035);
or U12789 (N_12789,N_9980,N_9785);
and U12790 (N_12790,N_7600,N_7879);
or U12791 (N_12791,N_10971,N_7703);
nand U12792 (N_12792,N_9071,N_11809);
and U12793 (N_12793,N_8297,N_7127);
xor U12794 (N_12794,N_7328,N_11036);
and U12795 (N_12795,N_10929,N_9824);
and U12796 (N_12796,N_11155,N_6641);
xnor U12797 (N_12797,N_9752,N_11389);
xor U12798 (N_12798,N_7439,N_6732);
and U12799 (N_12799,N_10719,N_11617);
nor U12800 (N_12800,N_10373,N_11110);
and U12801 (N_12801,N_9352,N_11400);
and U12802 (N_12802,N_7118,N_7106);
xor U12803 (N_12803,N_11228,N_10965);
nor U12804 (N_12804,N_9337,N_7405);
xnor U12805 (N_12805,N_7291,N_10359);
xnor U12806 (N_12806,N_8844,N_7190);
nor U12807 (N_12807,N_10737,N_8628);
and U12808 (N_12808,N_10423,N_8490);
nand U12809 (N_12809,N_8197,N_8177);
nand U12810 (N_12810,N_11276,N_6961);
nand U12811 (N_12811,N_10617,N_11750);
or U12812 (N_12812,N_6402,N_10392);
nor U12813 (N_12813,N_10607,N_8724);
nand U12814 (N_12814,N_8132,N_10391);
xnor U12815 (N_12815,N_7334,N_10093);
or U12816 (N_12816,N_10610,N_6921);
nor U12817 (N_12817,N_9153,N_10383);
or U12818 (N_12818,N_6188,N_10500);
and U12819 (N_12819,N_8960,N_11143);
nor U12820 (N_12820,N_8303,N_6396);
xor U12821 (N_12821,N_9297,N_11082);
xor U12822 (N_12822,N_9194,N_6759);
and U12823 (N_12823,N_8988,N_6813);
xor U12824 (N_12824,N_8224,N_6542);
nor U12825 (N_12825,N_6896,N_11787);
xnor U12826 (N_12826,N_10485,N_11565);
nor U12827 (N_12827,N_10806,N_6746);
xnor U12828 (N_12828,N_10588,N_8914);
nor U12829 (N_12829,N_6495,N_8204);
or U12830 (N_12830,N_9127,N_6243);
xnor U12831 (N_12831,N_10056,N_9406);
or U12832 (N_12832,N_11671,N_10776);
or U12833 (N_12833,N_7843,N_11094);
or U12834 (N_12834,N_8399,N_8275);
or U12835 (N_12835,N_8816,N_7794);
nand U12836 (N_12836,N_8357,N_7161);
or U12837 (N_12837,N_7165,N_7671);
and U12838 (N_12838,N_9878,N_8229);
xnor U12839 (N_12839,N_6996,N_8539);
nand U12840 (N_12840,N_9819,N_8558);
or U12841 (N_12841,N_9773,N_9933);
and U12842 (N_12842,N_11644,N_10936);
and U12843 (N_12843,N_7859,N_9966);
and U12844 (N_12844,N_7942,N_7201);
nor U12845 (N_12845,N_10785,N_7960);
xnor U12846 (N_12846,N_7023,N_9142);
nand U12847 (N_12847,N_9860,N_11136);
and U12848 (N_12848,N_6234,N_8910);
or U12849 (N_12849,N_7580,N_11345);
nor U12850 (N_12850,N_11990,N_9180);
or U12851 (N_12851,N_11645,N_11670);
nand U12852 (N_12852,N_9975,N_6886);
xor U12853 (N_12853,N_11358,N_11848);
nor U12854 (N_12854,N_7775,N_6138);
nand U12855 (N_12855,N_10656,N_10581);
nor U12856 (N_12856,N_11308,N_9491);
or U12857 (N_12857,N_7717,N_9113);
or U12858 (N_12858,N_8745,N_7293);
and U12859 (N_12859,N_6917,N_6774);
xor U12860 (N_12860,N_6442,N_10183);
xnor U12861 (N_12861,N_9478,N_6958);
nand U12862 (N_12862,N_6537,N_11863);
or U12863 (N_12863,N_9353,N_6794);
nor U12864 (N_12864,N_8337,N_8940);
or U12865 (N_12865,N_9441,N_10812);
or U12866 (N_12866,N_10463,N_10797);
or U12867 (N_12867,N_10130,N_6139);
xnor U12868 (N_12868,N_6933,N_11864);
nor U12869 (N_12869,N_6133,N_10626);
and U12870 (N_12870,N_9833,N_8018);
and U12871 (N_12871,N_9230,N_7115);
nor U12872 (N_12872,N_9067,N_8769);
or U12873 (N_12873,N_11688,N_7736);
and U12874 (N_12874,N_7317,N_6955);
nand U12875 (N_12875,N_9520,N_7358);
and U12876 (N_12876,N_6908,N_11721);
nor U12877 (N_12877,N_7831,N_7428);
or U12878 (N_12878,N_10398,N_8918);
nand U12879 (N_12879,N_11468,N_10302);
xor U12880 (N_12880,N_7186,N_6451);
nand U12881 (N_12881,N_11181,N_10823);
xor U12882 (N_12882,N_8163,N_9661);
or U12883 (N_12883,N_6535,N_10102);
and U12884 (N_12884,N_6558,N_6211);
nand U12885 (N_12885,N_7461,N_8982);
nor U12886 (N_12886,N_9800,N_8520);
nor U12887 (N_12887,N_7059,N_9895);
and U12888 (N_12888,N_8715,N_10445);
nor U12889 (N_12889,N_6486,N_6326);
or U12890 (N_12890,N_6499,N_7388);
or U12891 (N_12891,N_10218,N_10291);
and U12892 (N_12892,N_8953,N_9557);
nor U12893 (N_12893,N_11441,N_9920);
nor U12894 (N_12894,N_11053,N_11585);
or U12895 (N_12895,N_8201,N_10050);
nand U12896 (N_12896,N_8001,N_9903);
nand U12897 (N_12897,N_11829,N_6487);
and U12898 (N_12898,N_11711,N_8804);
or U12899 (N_12899,N_7533,N_8006);
xor U12900 (N_12900,N_10535,N_11418);
nand U12901 (N_12901,N_9214,N_10257);
or U12902 (N_12902,N_9538,N_11544);
and U12903 (N_12903,N_11092,N_8989);
or U12904 (N_12904,N_6013,N_9138);
xor U12905 (N_12905,N_6045,N_11364);
nand U12906 (N_12906,N_8868,N_9664);
or U12907 (N_12907,N_11911,N_7820);
and U12908 (N_12908,N_8384,N_8714);
and U12909 (N_12909,N_9363,N_10895);
or U12910 (N_12910,N_8071,N_11177);
xnor U12911 (N_12911,N_8564,N_6153);
nand U12912 (N_12912,N_7809,N_6693);
nand U12913 (N_12913,N_8489,N_9732);
and U12914 (N_12914,N_10313,N_7198);
xnor U12915 (N_12915,N_7519,N_10440);
and U12916 (N_12916,N_8059,N_8790);
nand U12917 (N_12917,N_10527,N_7916);
xor U12918 (N_12918,N_11349,N_9440);
nor U12919 (N_12919,N_6595,N_10548);
and U12920 (N_12920,N_8508,N_9164);
nand U12921 (N_12921,N_8519,N_8970);
and U12922 (N_12922,N_6631,N_11888);
or U12923 (N_12923,N_11998,N_10855);
xnor U12924 (N_12924,N_9599,N_6945);
xnor U12925 (N_12925,N_6934,N_10689);
xor U12926 (N_12926,N_6776,N_10533);
and U12927 (N_12927,N_11590,N_11275);
nor U12928 (N_12928,N_8896,N_7697);
xnor U12929 (N_12929,N_6032,N_7053);
and U12930 (N_12930,N_11023,N_10008);
nor U12931 (N_12931,N_9516,N_6572);
and U12932 (N_12932,N_7693,N_6290);
and U12933 (N_12933,N_11066,N_11939);
xor U12934 (N_12934,N_9764,N_6723);
and U12935 (N_12935,N_8395,N_6119);
or U12936 (N_12936,N_6811,N_8975);
nand U12937 (N_12937,N_6350,N_9781);
nor U12938 (N_12938,N_7720,N_10638);
and U12939 (N_12939,N_8499,N_8830);
and U12940 (N_12940,N_10517,N_9476);
nor U12941 (N_12941,N_8645,N_6516);
or U12942 (N_12942,N_7102,N_7393);
or U12943 (N_12943,N_10715,N_8044);
xnor U12944 (N_12944,N_8627,N_6056);
xor U12945 (N_12945,N_11499,N_9454);
and U12946 (N_12946,N_9004,N_8879);
nor U12947 (N_12947,N_6409,N_6073);
xnor U12948 (N_12948,N_9218,N_6801);
xnor U12949 (N_12949,N_10154,N_9730);
or U12950 (N_12950,N_9856,N_11768);
and U12951 (N_12951,N_10621,N_9863);
xor U12952 (N_12952,N_11871,N_6293);
xor U12953 (N_12953,N_6521,N_11936);
xnor U12954 (N_12954,N_10427,N_11270);
and U12955 (N_12955,N_9606,N_11988);
nand U12956 (N_12956,N_9329,N_9968);
nand U12957 (N_12957,N_6371,N_7517);
and U12958 (N_12958,N_6105,N_8315);
nand U12959 (N_12959,N_7459,N_7660);
xor U12960 (N_12960,N_11375,N_10324);
xnor U12961 (N_12961,N_7366,N_11600);
and U12962 (N_12962,N_10408,N_8345);
or U12963 (N_12963,N_6683,N_10727);
nor U12964 (N_12964,N_11586,N_6630);
and U12965 (N_12965,N_7948,N_8241);
or U12966 (N_12966,N_11112,N_8578);
nor U12967 (N_12967,N_10634,N_9236);
xnor U12968 (N_12968,N_8102,N_10930);
nor U12969 (N_12969,N_6336,N_7564);
nor U12970 (N_12970,N_7084,N_8081);
and U12971 (N_12971,N_7592,N_9988);
and U12972 (N_12972,N_9258,N_9252);
or U12973 (N_12973,N_11898,N_10207);
nand U12974 (N_12974,N_7068,N_9031);
nand U12975 (N_12975,N_7709,N_6704);
xor U12976 (N_12976,N_11452,N_10746);
or U12977 (N_12977,N_9995,N_9567);
or U12978 (N_12978,N_7318,N_11200);
or U12979 (N_12979,N_6240,N_6206);
nor U12980 (N_12980,N_10521,N_6860);
xor U12981 (N_12981,N_9116,N_9124);
xor U12982 (N_12982,N_6883,N_6596);
or U12983 (N_12983,N_10516,N_8810);
xor U12984 (N_12984,N_6076,N_7294);
xor U12985 (N_12985,N_11015,N_8571);
and U12986 (N_12986,N_11044,N_11761);
nor U12987 (N_12987,N_8455,N_6639);
and U12988 (N_12988,N_10119,N_8696);
nand U12989 (N_12989,N_10455,N_6780);
nand U12990 (N_12990,N_10483,N_6898);
or U12991 (N_12991,N_6750,N_9405);
xnor U12992 (N_12992,N_11225,N_7019);
or U12993 (N_12993,N_7889,N_8189);
or U12994 (N_12994,N_11611,N_7767);
or U12995 (N_12995,N_9499,N_10395);
nor U12996 (N_12996,N_10576,N_7119);
xnor U12997 (N_12997,N_8575,N_10821);
or U12998 (N_12998,N_9137,N_7634);
nor U12999 (N_12999,N_8421,N_7548);
and U13000 (N_13000,N_7244,N_6895);
and U13001 (N_13001,N_11354,N_10696);
or U13002 (N_13002,N_11039,N_11823);
xnor U13003 (N_13003,N_6593,N_11786);
nor U13004 (N_13004,N_9271,N_9675);
and U13005 (N_13005,N_9396,N_11851);
xnor U13006 (N_13006,N_7845,N_6556);
nand U13007 (N_13007,N_7787,N_9720);
or U13008 (N_13008,N_10852,N_7455);
nand U13009 (N_13009,N_8474,N_10165);
or U13010 (N_13010,N_7978,N_9074);
nor U13011 (N_13011,N_9945,N_11204);
xnor U13012 (N_13012,N_11469,N_7598);
or U13013 (N_13013,N_11108,N_8215);
or U13014 (N_13014,N_7936,N_9237);
and U13015 (N_13015,N_8460,N_10811);
nor U13016 (N_13016,N_9656,N_7016);
and U13017 (N_13017,N_7884,N_8432);
xor U13018 (N_13018,N_10605,N_6217);
nand U13019 (N_13019,N_6580,N_8274);
nor U13020 (N_13020,N_6061,N_11803);
and U13021 (N_13021,N_11147,N_6570);
xnor U13022 (N_13022,N_6224,N_9272);
nor U13023 (N_13023,N_9722,N_9334);
nand U13024 (N_13024,N_8514,N_8846);
nand U13025 (N_13025,N_8471,N_7425);
and U13026 (N_13026,N_11509,N_7375);
or U13027 (N_13027,N_8281,N_10630);
nand U13028 (N_13028,N_7543,N_8797);
xnor U13029 (N_13029,N_8053,N_7049);
nor U13030 (N_13030,N_10541,N_8257);
nor U13031 (N_13031,N_6067,N_9241);
and U13032 (N_13032,N_8165,N_6353);
nand U13033 (N_13033,N_9992,N_11172);
and U13034 (N_13034,N_7631,N_8103);
xnor U13035 (N_13035,N_7486,N_6308);
and U13036 (N_13036,N_6840,N_9662);
xnor U13037 (N_13037,N_8541,N_10799);
nor U13038 (N_13038,N_7438,N_7185);
nand U13039 (N_13039,N_10380,N_7675);
xnor U13040 (N_13040,N_7374,N_9937);
nand U13041 (N_13041,N_11475,N_9851);
and U13042 (N_13042,N_8466,N_8213);
xnor U13043 (N_13043,N_10980,N_7808);
nor U13044 (N_13044,N_11682,N_9962);
or U13045 (N_13045,N_6118,N_10566);
nand U13046 (N_13046,N_9112,N_9410);
xor U13047 (N_13047,N_9285,N_10514);
nor U13048 (N_13048,N_8770,N_9700);
xnor U13049 (N_13049,N_7730,N_10025);
xor U13050 (N_13050,N_11913,N_11746);
or U13051 (N_13051,N_8005,N_7332);
nor U13052 (N_13052,N_8796,N_8533);
or U13053 (N_13053,N_6960,N_9542);
and U13054 (N_13054,N_11185,N_7096);
or U13055 (N_13055,N_6529,N_9055);
nand U13056 (N_13056,N_10353,N_8458);
and U13057 (N_13057,N_8905,N_7768);
nand U13058 (N_13058,N_11030,N_6427);
or U13059 (N_13059,N_10831,N_6286);
xnor U13060 (N_13060,N_7236,N_6658);
nor U13061 (N_13061,N_10401,N_11854);
xnor U13062 (N_13062,N_9250,N_8339);
nand U13063 (N_13063,N_9222,N_9971);
nand U13064 (N_13064,N_9104,N_10311);
nand U13065 (N_13065,N_11929,N_10040);
and U13066 (N_13066,N_9234,N_6062);
nor U13067 (N_13067,N_8791,N_9339);
nor U13068 (N_13068,N_10699,N_6517);
nand U13069 (N_13069,N_10777,N_6178);
nor U13070 (N_13070,N_6878,N_10424);
nor U13071 (N_13071,N_10973,N_7166);
nand U13072 (N_13072,N_9669,N_6729);
xnor U13073 (N_13073,N_7908,N_11782);
and U13074 (N_13074,N_10430,N_8494);
nor U13075 (N_13075,N_7339,N_7741);
and U13076 (N_13076,N_8551,N_9620);
xnor U13077 (N_13077,N_8196,N_10083);
xor U13078 (N_13078,N_6849,N_6882);
nor U13079 (N_13079,N_10567,N_11729);
xnor U13080 (N_13080,N_7647,N_9754);
xor U13081 (N_13081,N_10286,N_8492);
xor U13082 (N_13082,N_10506,N_11980);
xnor U13083 (N_13083,N_7349,N_6493);
and U13084 (N_13084,N_9657,N_10690);
and U13085 (N_13085,N_7964,N_6665);
nor U13086 (N_13086,N_9981,N_8887);
nor U13087 (N_13087,N_9110,N_8397);
xor U13088 (N_13088,N_11470,N_6389);
xnor U13089 (N_13089,N_7225,N_8050);
nand U13090 (N_13090,N_7204,N_7573);
or U13091 (N_13091,N_8476,N_11285);
xnor U13092 (N_13092,N_7136,N_6629);
nand U13093 (N_13093,N_7773,N_8453);
nor U13094 (N_13094,N_7278,N_8968);
nand U13095 (N_13095,N_9150,N_7493);
nor U13096 (N_13096,N_6359,N_7457);
nand U13097 (N_13097,N_6789,N_11777);
and U13098 (N_13098,N_8243,N_6287);
xnor U13099 (N_13099,N_9628,N_11690);
xnor U13100 (N_13100,N_7672,N_9445);
and U13101 (N_13101,N_6420,N_11317);
nand U13102 (N_13102,N_7885,N_11838);
or U13103 (N_13103,N_7781,N_10544);
nor U13104 (N_13104,N_11167,N_10498);
nor U13105 (N_13105,N_8920,N_9467);
nand U13106 (N_13106,N_9151,N_11057);
nor U13107 (N_13107,N_8884,N_7938);
and U13108 (N_13108,N_7643,N_6489);
or U13109 (N_13109,N_9923,N_6239);
nor U13110 (N_13110,N_6748,N_6951);
xnor U13111 (N_13111,N_7664,N_11719);
nand U13112 (N_13112,N_8750,N_10020);
and U13113 (N_13113,N_8635,N_10882);
nand U13114 (N_13114,N_8969,N_6956);
xnor U13115 (N_13115,N_11226,N_11064);
nor U13116 (N_13116,N_10620,N_8148);
nand U13117 (N_13117,N_6237,N_10167);
and U13118 (N_13118,N_9867,N_6914);
nand U13119 (N_13119,N_8602,N_11047);
xor U13120 (N_13120,N_7979,N_9707);
or U13121 (N_13121,N_9721,N_11344);
or U13122 (N_13122,N_10528,N_11649);
nor U13123 (N_13123,N_9191,N_11865);
nand U13124 (N_13124,N_11102,N_7097);
or U13125 (N_13125,N_9346,N_10162);
nand U13126 (N_13126,N_7784,N_6276);
nor U13127 (N_13127,N_9228,N_8004);
or U13128 (N_13128,N_8169,N_7894);
nor U13129 (N_13129,N_6355,N_7259);
xor U13130 (N_13130,N_9817,N_8442);
nor U13131 (N_13131,N_7673,N_11904);
nor U13132 (N_13132,N_10595,N_11342);
nand U13133 (N_13133,N_10303,N_11949);
xnor U13134 (N_13134,N_8669,N_11927);
or U13135 (N_13135,N_6049,N_8815);
nand U13136 (N_13136,N_9791,N_7249);
and U13137 (N_13137,N_10526,N_11279);
or U13138 (N_13138,N_9326,N_9443);
or U13139 (N_13139,N_8957,N_8130);
nor U13140 (N_13140,N_11637,N_8853);
or U13141 (N_13141,N_9161,N_9002);
or U13142 (N_13142,N_7183,N_8011);
nand U13143 (N_13143,N_10344,N_9616);
and U13144 (N_13144,N_7829,N_7028);
and U13145 (N_13145,N_6797,N_9277);
xnor U13146 (N_13146,N_9861,N_7104);
xnor U13147 (N_13147,N_6416,N_11704);
xnor U13148 (N_13148,N_8477,N_8037);
or U13149 (N_13149,N_6740,N_7841);
or U13150 (N_13150,N_7684,N_6195);
nor U13151 (N_13151,N_10046,N_7637);
or U13152 (N_13152,N_6241,N_10926);
nand U13153 (N_13153,N_9471,N_8531);
or U13154 (N_13154,N_10121,N_11503);
or U13155 (N_13155,N_10809,N_7143);
xnor U13156 (N_13156,N_9974,N_10067);
and U13157 (N_13157,N_8404,N_7329);
xnor U13158 (N_13158,N_10420,N_10492);
xor U13159 (N_13159,N_11591,N_7642);
nor U13160 (N_13160,N_9569,N_10608);
xnor U13161 (N_13161,N_11497,N_7521);
and U13162 (N_13162,N_11500,N_9154);
xnor U13163 (N_13163,N_8954,N_6566);
xor U13164 (N_13164,N_9179,N_10284);
and U13165 (N_13165,N_6055,N_10903);
nor U13166 (N_13166,N_9313,N_11545);
or U13167 (N_13167,N_11599,N_9874);
and U13168 (N_13168,N_8604,N_10267);
xor U13169 (N_13169,N_11118,N_6160);
and U13170 (N_13170,N_11531,N_9417);
nand U13171 (N_13171,N_10577,N_6146);
nand U13172 (N_13172,N_6042,N_6708);
and U13173 (N_13173,N_6701,N_10700);
or U13174 (N_13174,N_8863,N_6749);
xor U13175 (N_13175,N_10429,N_10640);
nor U13176 (N_13176,N_6798,N_11101);
and U13177 (N_13177,N_9088,N_7864);
nand U13178 (N_13178,N_11984,N_10835);
xor U13179 (N_13179,N_10010,N_8054);
or U13180 (N_13180,N_8950,N_6674);
nand U13181 (N_13181,N_11169,N_8209);
nor U13182 (N_13182,N_8068,N_8316);
or U13183 (N_13183,N_10584,N_9309);
xnor U13184 (N_13184,N_6710,N_10774);
nor U13185 (N_13185,N_11539,N_6632);
nor U13186 (N_13186,N_9204,N_11699);
or U13187 (N_13187,N_8097,N_10216);
or U13188 (N_13188,N_9976,N_11570);
xnor U13189 (N_13189,N_7903,N_7400);
or U13190 (N_13190,N_10736,N_6619);
xnor U13191 (N_13191,N_9681,N_7930);
nand U13192 (N_13192,N_9961,N_10891);
or U13193 (N_13193,N_9135,N_11474);
and U13194 (N_13194,N_11320,N_11012);
or U13195 (N_13195,N_8518,N_6091);
and U13196 (N_13196,N_9069,N_7765);
xor U13197 (N_13197,N_10779,N_10062);
nor U13198 (N_13198,N_11419,N_7805);
or U13199 (N_13199,N_9361,N_9987);
nor U13200 (N_13200,N_8079,N_7285);
xor U13201 (N_13201,N_6779,N_9523);
xor U13202 (N_13202,N_7628,N_10629);
or U13203 (N_13203,N_8987,N_6190);
and U13204 (N_13204,N_8468,N_7804);
nand U13205 (N_13205,N_8788,N_8396);
nand U13206 (N_13206,N_8496,N_6979);
or U13207 (N_13207,N_7154,N_10970);
nor U13208 (N_13208,N_10376,N_8605);
nor U13209 (N_13209,N_7570,N_7509);
nor U13210 (N_13210,N_8444,N_8728);
xor U13211 (N_13211,N_9209,N_6248);
and U13212 (N_13212,N_8528,N_7434);
xor U13213 (N_13213,N_8352,N_7746);
and U13214 (N_13214,N_6391,N_11528);
and U13215 (N_13215,N_9195,N_8772);
xnor U13216 (N_13216,N_9084,N_8823);
or U13217 (N_13217,N_7583,N_6903);
and U13218 (N_13218,N_9126,N_11569);
nand U13219 (N_13219,N_8389,N_8854);
nor U13220 (N_13220,N_11199,N_7435);
nand U13221 (N_13221,N_10692,N_6718);
xnor U13222 (N_13222,N_11489,N_10034);
or U13223 (N_13223,N_8693,N_9924);
or U13224 (N_13224,N_8329,N_7696);
or U13225 (N_13225,N_11139,N_6048);
xnor U13226 (N_13226,N_8310,N_8984);
nand U13227 (N_13227,N_11944,N_11914);
and U13228 (N_13228,N_10029,N_11368);
nor U13229 (N_13229,N_7069,N_7022);
and U13230 (N_13230,N_8304,N_9763);
xnor U13231 (N_13231,N_6548,N_8619);
nor U13232 (N_13232,N_11753,N_10522);
nand U13233 (N_13233,N_11206,N_8710);
or U13234 (N_13234,N_8871,N_8452);
and U13235 (N_13235,N_9365,N_9528);
and U13236 (N_13236,N_6233,N_6803);
nand U13237 (N_13237,N_10297,N_9211);
nor U13238 (N_13238,N_8995,N_7112);
nand U13239 (N_13239,N_9123,N_11899);
or U13240 (N_13240,N_8802,N_6788);
xnor U13241 (N_13241,N_10188,N_9938);
or U13242 (N_13242,N_11689,N_9415);
xnor U13243 (N_13243,N_6362,N_6373);
nand U13244 (N_13244,N_7680,N_8785);
and U13245 (N_13245,N_9047,N_7219);
xnor U13246 (N_13246,N_6651,N_8220);
nor U13247 (N_13247,N_10857,N_11971);
or U13248 (N_13248,N_6876,N_10778);
nand U13249 (N_13249,N_9502,N_7365);
xor U13250 (N_13250,N_6478,N_10296);
or U13251 (N_13251,N_9156,N_8087);
or U13252 (N_13252,N_11009,N_9598);
nand U13253 (N_13253,N_7712,N_7057);
nand U13254 (N_13254,N_8568,N_8233);
nor U13255 (N_13255,N_8803,N_7412);
xor U13256 (N_13256,N_11471,N_10529);
nand U13257 (N_13257,N_7267,N_11437);
xor U13258 (N_13258,N_6283,N_10601);
nor U13259 (N_13259,N_10854,N_6621);
xor U13260 (N_13260,N_8534,N_10738);
and U13261 (N_13261,N_6688,N_9028);
xor U13262 (N_13262,N_7424,N_7027);
xnor U13263 (N_13263,N_10771,N_9244);
xnor U13264 (N_13264,N_11054,N_10657);
xor U13265 (N_13265,N_6302,N_7065);
nor U13266 (N_13266,N_7021,N_7772);
or U13267 (N_13267,N_8222,N_6561);
nand U13268 (N_13268,N_9883,N_10880);
nor U13269 (N_13269,N_10048,N_7961);
nand U13270 (N_13270,N_10341,N_10441);
or U13271 (N_13271,N_7962,N_9481);
or U13272 (N_13272,N_8020,N_6204);
xnor U13273 (N_13273,N_8198,N_8617);
or U13274 (N_13274,N_10969,N_8221);
xnor U13275 (N_13275,N_9459,N_11874);
xnor U13276 (N_13276,N_7800,N_7420);
nor U13277 (N_13277,N_6575,N_6426);
or U13278 (N_13278,N_8717,N_11996);
xnor U13279 (N_13279,N_6856,N_11732);
nand U13280 (N_13280,N_7528,N_7450);
nor U13281 (N_13281,N_11268,N_8654);
nand U13282 (N_13282,N_11283,N_7742);
or U13283 (N_13283,N_11763,N_7299);
xnor U13284 (N_13284,N_10717,N_10448);
nand U13285 (N_13285,N_11380,N_8718);
nand U13286 (N_13286,N_6483,N_6372);
nor U13287 (N_13287,N_8013,N_9392);
xnor U13288 (N_13288,N_6966,N_10407);
and U13289 (N_13289,N_10143,N_7749);
nor U13290 (N_13290,N_9559,N_6752);
nand U13291 (N_13291,N_6397,N_11879);
nor U13292 (N_13292,N_10687,N_7690);
or U13293 (N_13293,N_6210,N_7963);
or U13294 (N_13294,N_7314,N_9638);
xnor U13295 (N_13295,N_6050,N_8827);
nand U13296 (N_13296,N_11378,N_11775);
nand U13297 (N_13297,N_10682,N_6830);
xnor U13298 (N_13298,N_10729,N_11673);
or U13299 (N_13299,N_11700,N_9294);
or U13300 (N_13300,N_11407,N_6114);
nand U13301 (N_13301,N_8587,N_10443);
or U13302 (N_13302,N_9859,N_10135);
nand U13303 (N_13303,N_9125,N_7320);
and U13304 (N_13304,N_8500,N_8650);
xnor U13305 (N_13305,N_9169,N_11880);
and U13306 (N_13306,N_8695,N_8779);
and U13307 (N_13307,N_11010,N_10921);
nand U13308 (N_13308,N_7832,N_11783);
nor U13309 (N_13309,N_10681,N_8298);
and U13310 (N_13310,N_10104,N_7751);
and U13311 (N_13311,N_7342,N_10475);
nor U13312 (N_13312,N_6264,N_8809);
nand U13313 (N_13313,N_10901,N_6464);
or U13314 (N_13314,N_8112,N_7855);
nor U13315 (N_13315,N_8273,N_7933);
and U13316 (N_13316,N_7217,N_10223);
or U13317 (N_13317,N_11146,N_6327);
nand U13318 (N_13318,N_11905,N_9853);
and U13319 (N_13319,N_10090,N_11762);
nor U13320 (N_13320,N_9316,N_6136);
nor U13321 (N_13321,N_10712,N_10232);
and U13322 (N_13322,N_6993,N_10328);
xor U13323 (N_13323,N_9457,N_8800);
nor U13324 (N_13324,N_7122,N_6282);
and U13325 (N_13325,N_6261,N_7925);
or U13326 (N_13326,N_11620,N_6600);
nor U13327 (N_13327,N_6202,N_9210);
xnor U13328 (N_13328,N_7937,N_9488);
nor U13329 (N_13329,N_9658,N_6944);
nor U13330 (N_13330,N_8266,N_9265);
xnor U13331 (N_13331,N_10164,N_10832);
nor U13332 (N_13332,N_10755,N_9419);
nand U13333 (N_13333,N_8376,N_11087);
xnor U13334 (N_13334,N_10757,N_8270);
or U13335 (N_13335,N_10403,N_8536);
or U13336 (N_13336,N_9637,N_6905);
or U13337 (N_13337,N_7325,N_11444);
xnor U13338 (N_13338,N_9336,N_6744);
xor U13339 (N_13339,N_8553,N_8254);
nand U13340 (N_13340,N_6975,N_7527);
or U13341 (N_13341,N_8480,N_9061);
and U13342 (N_13342,N_6574,N_11197);
or U13343 (N_13343,N_8382,N_6018);
or U13344 (N_13344,N_11182,N_9910);
nor U13345 (N_13345,N_10984,N_10371);
xnor U13346 (N_13346,N_6384,N_10968);
xnor U13347 (N_13347,N_6398,N_6112);
nand U13348 (N_13348,N_8250,N_7803);
or U13349 (N_13349,N_10329,N_11659);
nor U13350 (N_13350,N_8109,N_11363);
nor U13351 (N_13351,N_11072,N_10318);
and U13352 (N_13352,N_8117,N_8872);
or U13353 (N_13353,N_11020,N_8609);
nor U13354 (N_13354,N_9076,N_6218);
xnor U13355 (N_13355,N_7085,N_7549);
nor U13356 (N_13356,N_11445,N_9276);
and U13357 (N_13357,N_9615,N_8760);
xor U13358 (N_13358,N_7419,N_10713);
xnor U13359 (N_13359,N_7402,N_11784);
or U13360 (N_13360,N_8735,N_6184);
or U13361 (N_13361,N_7015,N_9544);
and U13362 (N_13362,N_9310,N_8817);
xor U13363 (N_13363,N_9782,N_7901);
and U13364 (N_13364,N_11749,N_10627);
nor U13365 (N_13365,N_9325,N_10844);
nor U13366 (N_13366,N_6006,N_9594);
xnor U13367 (N_13367,N_9778,N_10394);
nor U13368 (N_13368,N_10909,N_11430);
and U13369 (N_13369,N_8567,N_11314);
nand U13370 (N_13370,N_11351,N_10602);
and U13371 (N_13371,N_9967,N_10071);
nor U13372 (N_13372,N_10562,N_7559);
nand U13373 (N_13373,N_9550,N_11780);
xnor U13374 (N_13374,N_11640,N_7790);
nand U13375 (N_13375,N_6408,N_10502);
xnor U13376 (N_13376,N_11062,N_10707);
and U13377 (N_13377,N_10637,N_6672);
nand U13378 (N_13378,N_10479,N_10105);
xor U13379 (N_13379,N_8212,N_8517);
nand U13380 (N_13380,N_6965,N_7440);
nor U13381 (N_13381,N_7130,N_11245);
and U13382 (N_13382,N_8388,N_7061);
and U13383 (N_13383,N_9333,N_9932);
or U13384 (N_13384,N_6564,N_7431);
or U13385 (N_13385,N_8238,N_7515);
nand U13386 (N_13386,N_10281,N_6470);
or U13387 (N_13387,N_6577,N_10058);
or U13388 (N_13388,N_10592,N_9382);
nor U13389 (N_13389,N_11945,N_6292);
nor U13390 (N_13390,N_9019,N_7969);
and U13391 (N_13391,N_8048,N_8253);
and U13392 (N_13392,N_8472,N_6063);
nor U13393 (N_13393,N_6668,N_9922);
and U13394 (N_13394,N_10676,N_8341);
xor U13395 (N_13395,N_8036,N_8632);
nand U13396 (N_13396,N_11148,N_11439);
or U13397 (N_13397,N_10358,N_8441);
xnor U13398 (N_13398,N_6679,N_7630);
nor U13399 (N_13399,N_9808,N_9220);
and U13400 (N_13400,N_8234,N_9070);
nor U13401 (N_13401,N_8913,N_10504);
nor U13402 (N_13402,N_9919,N_11410);
nor U13403 (N_13403,N_6863,N_7213);
nand U13404 (N_13404,N_11495,N_11691);
nor U13405 (N_13405,N_8633,N_6501);
or U13406 (N_13406,N_9100,N_7968);
xor U13407 (N_13407,N_8255,N_11272);
nand U13408 (N_13408,N_8705,N_10466);
nor U13409 (N_13409,N_11257,N_9356);
nor U13410 (N_13410,N_11901,N_6544);
xnor U13411 (N_13411,N_9519,N_10396);
and U13412 (N_13412,N_11309,N_7608);
nand U13413 (N_13413,N_8684,N_10226);
nand U13414 (N_13414,N_6403,N_8675);
or U13415 (N_13415,N_7050,N_7417);
or U13416 (N_13416,N_8190,N_8139);
nand U13417 (N_13417,N_8685,N_8042);
nand U13418 (N_13418,N_8256,N_6870);
xnor U13419 (N_13419,N_6737,N_9163);
xor U13420 (N_13420,N_11537,N_11658);
nor U13421 (N_13421,N_7295,N_7208);
or U13422 (N_13422,N_11166,N_8168);
or U13423 (N_13423,N_9632,N_10653);
or U13424 (N_13424,N_11103,N_6007);
xor U13425 (N_13425,N_7735,N_10963);
nor U13426 (N_13426,N_10128,N_8596);
nand U13427 (N_13427,N_7012,N_8406);
xnor U13428 (N_13428,N_6726,N_7602);
nand U13429 (N_13429,N_7169,N_7738);
and U13430 (N_13430,N_7310,N_6465);
xor U13431 (N_13431,N_6284,N_6597);
nand U13432 (N_13432,N_9102,N_8701);
nor U13433 (N_13433,N_6638,N_6821);
or U13434 (N_13434,N_11265,N_10655);
and U13435 (N_13435,N_9521,N_11395);
nand U13436 (N_13436,N_6182,N_7002);
nor U13437 (N_13437,N_11423,N_8125);
xnor U13438 (N_13438,N_8847,N_7896);
or U13439 (N_13439,N_10709,N_6490);
and U13440 (N_13440,N_7566,N_9430);
nor U13441 (N_13441,N_7802,N_9496);
xnor U13442 (N_13442,N_8686,N_6165);
or U13443 (N_13443,N_9139,N_7534);
or U13444 (N_13444,N_8880,N_9977);
nand U13445 (N_13445,N_6871,N_7035);
or U13446 (N_13446,N_11648,N_8979);
or U13447 (N_13447,N_8806,N_9390);
or U13448 (N_13448,N_7140,N_10148);
and U13449 (N_13449,N_10259,N_9724);
and U13450 (N_13450,N_7340,N_9570);
and U13451 (N_13451,N_9424,N_11549);
and U13452 (N_13452,N_7492,N_8833);
xnor U13453 (N_13453,N_11808,N_9568);
nor U13454 (N_13454,N_7221,N_11414);
and U13455 (N_13455,N_6894,N_6852);
or U13456 (N_13456,N_9427,N_10349);
or U13457 (N_13457,N_9332,N_10367);
xor U13458 (N_13458,N_6024,N_8682);
nand U13459 (N_13459,N_11333,N_10274);
nor U13460 (N_13460,N_9812,N_11557);
and U13461 (N_13461,N_11722,N_6046);
or U13462 (N_13462,N_9952,N_11370);
nor U13463 (N_13463,N_10839,N_8664);
nor U13464 (N_13464,N_7212,N_9736);
nand U13465 (N_13465,N_8291,N_6004);
xor U13466 (N_13466,N_9622,N_8375);
nand U13467 (N_13467,N_9077,N_7128);
xor U13468 (N_13468,N_9115,N_7835);
and U13469 (N_13469,N_7792,N_9571);
xnor U13470 (N_13470,N_8227,N_10856);
or U13471 (N_13471,N_9227,N_6364);
nor U13472 (N_13472,N_7337,N_9811);
and U13473 (N_13473,N_6953,N_8801);
or U13474 (N_13474,N_11912,N_10561);
and U13475 (N_13475,N_11472,N_7575);
nor U13476 (N_13476,N_7589,N_9174);
xor U13477 (N_13477,N_6986,N_11307);
and U13478 (N_13478,N_10666,N_8340);
or U13479 (N_13479,N_10036,N_10248);
nor U13480 (N_13480,N_7966,N_9900);
nand U13481 (N_13481,N_10591,N_9465);
xnor U13482 (N_13482,N_9079,N_7270);
xnor U13483 (N_13483,N_8993,N_6976);
and U13484 (N_13484,N_10454,N_11563);
and U13485 (N_13485,N_9864,N_8446);
and U13486 (N_13486,N_6229,N_11962);
and U13487 (N_13487,N_10691,N_7877);
nor U13488 (N_13488,N_10208,N_11618);
and U13489 (N_13489,N_8392,N_9784);
or U13490 (N_13490,N_7607,N_11847);
and U13491 (N_13491,N_6219,N_6724);
or U13492 (N_13492,N_7904,N_7394);
and U13493 (N_13493,N_8765,N_7089);
or U13494 (N_13494,N_11893,N_7120);
nor U13495 (N_13495,N_8938,N_10586);
nor U13496 (N_13496,N_8733,N_7209);
nor U13497 (N_13497,N_7308,N_11526);
or U13498 (N_13498,N_10573,N_6411);
nand U13499 (N_13499,N_10041,N_9224);
nand U13500 (N_13500,N_11816,N_10174);
xor U13501 (N_13501,N_8876,N_8573);
and U13502 (N_13502,N_9841,N_9370);
and U13503 (N_13503,N_9477,N_7914);
nand U13504 (N_13504,N_10030,N_6379);
and U13505 (N_13505,N_6102,N_8923);
xor U13506 (N_13506,N_6598,N_8743);
xnor U13507 (N_13507,N_11294,N_10955);
and U13508 (N_13508,N_11014,N_7125);
and U13509 (N_13509,N_6661,N_9871);
xnor U13510 (N_13510,N_9843,N_6288);
nand U13511 (N_13511,N_7954,N_6773);
and U13512 (N_13512,N_8267,N_9865);
nor U13513 (N_13513,N_8875,N_10428);
nor U13514 (N_13514,N_8526,N_6555);
nor U13515 (N_13515,N_8966,N_10701);
xnor U13516 (N_13516,N_7223,N_8670);
and U13517 (N_13517,N_6839,N_10320);
and U13518 (N_13518,N_10026,N_9892);
nand U13519 (N_13519,N_11216,N_8947);
xnor U13520 (N_13520,N_7981,N_8475);
and U13521 (N_13521,N_10987,N_9458);
xor U13522 (N_13522,N_9399,N_9042);
nand U13523 (N_13523,N_6430,N_8762);
and U13524 (N_13524,N_11341,N_6931);
xor U13525 (N_13525,N_6606,N_11981);
nor U13526 (N_13526,N_11222,N_6637);
and U13527 (N_13527,N_7210,N_8120);
xor U13528 (N_13528,N_8631,N_8194);
or U13529 (N_13529,N_10578,N_6475);
nor U13530 (N_13530,N_6223,N_8326);
xnor U13531 (N_13531,N_11607,N_7272);
nor U13532 (N_13532,N_10206,N_6833);
or U13533 (N_13533,N_10859,N_10237);
nor U13534 (N_13534,N_10758,N_7973);
nor U13535 (N_13535,N_6612,N_6712);
nand U13536 (N_13536,N_8838,N_9830);
nor U13537 (N_13537,N_7920,N_11629);
xor U13538 (N_13538,N_8997,N_9790);
nand U13539 (N_13539,N_9311,N_8023);
nand U13540 (N_13540,N_8400,N_6214);
or U13541 (N_13541,N_11651,N_11697);
nor U13542 (N_13542,N_10928,N_10841);
xnor U13543 (N_13543,N_7442,N_9060);
or U13544 (N_13544,N_10938,N_8272);
xor U13545 (N_13545,N_8798,N_8231);
nand U13546 (N_13546,N_11655,N_6453);
nand U13547 (N_13547,N_6756,N_7191);
and U13548 (N_13548,N_7384,N_6504);
nor U13549 (N_13549,N_7449,N_9319);
nand U13550 (N_13550,N_8007,N_7757);
and U13551 (N_13551,N_8239,N_6358);
xnor U13552 (N_13552,N_10004,N_7584);
or U13553 (N_13553,N_9397,N_6584);
and U13554 (N_13554,N_8487,N_11817);
and U13555 (N_13555,N_7944,N_6070);
or U13556 (N_13556,N_9187,N_8897);
nand U13557 (N_13557,N_8668,N_6348);
nor U13558 (N_13558,N_7487,N_8293);
and U13559 (N_13559,N_9173,N_6134);
xor U13560 (N_13560,N_7214,N_11540);
and U13561 (N_13561,N_7164,N_8956);
or U13562 (N_13562,N_8886,N_10805);
and U13563 (N_13563,N_11547,N_8666);
or U13564 (N_13564,N_11325,N_11156);
and U13565 (N_13565,N_8930,N_7116);
nand U13566 (N_13566,N_11402,N_8080);
xnor U13567 (N_13567,N_10808,N_8597);
nor U13568 (N_13568,N_7396,N_8683);
nand U13569 (N_13569,N_8032,N_9733);
nand U13570 (N_13570,N_6482,N_10299);
nand U13571 (N_13571,N_9408,N_6298);
nor U13572 (N_13572,N_11373,N_7044);
nand U13573 (N_13573,N_8746,N_6097);
nor U13574 (N_13574,N_6071,N_6349);
or U13575 (N_13575,N_7857,N_10731);
xor U13576 (N_13576,N_11085,N_9420);
or U13577 (N_13577,N_7823,N_9595);
xor U13578 (N_13578,N_7520,N_6601);
xor U13579 (N_13579,N_8543,N_7740);
nand U13580 (N_13580,N_9779,N_8108);
nor U13581 (N_13581,N_10828,N_9708);
and U13582 (N_13582,N_9556,N_6912);
xnor U13583 (N_13583,N_9685,N_6885);
nand U13584 (N_13584,N_7853,N_11524);
nor U13585 (N_13585,N_8653,N_7996);
xnor U13586 (N_13586,N_9242,N_8784);
nand U13587 (N_13587,N_10136,N_9460);
or U13588 (N_13588,N_8008,N_7718);
and U13589 (N_13589,N_10293,N_6143);
nand U13590 (N_13590,N_8459,N_7480);
nor U13591 (N_13591,N_9840,N_8155);
or U13592 (N_13592,N_6547,N_6235);
or U13593 (N_13593,N_9936,N_10219);
or U13594 (N_13594,N_9758,N_9273);
xnor U13595 (N_13595,N_9727,N_6950);
nand U13596 (N_13596,N_10883,N_9942);
nand U13597 (N_13597,N_9750,N_7569);
and U13598 (N_13598,N_7710,N_6711);
and U13599 (N_13599,N_7175,N_7283);
xnor U13600 (N_13600,N_11856,N_10140);
and U13601 (N_13601,N_11175,N_11381);
or U13602 (N_13602,N_9456,N_7711);
nor U13603 (N_13603,N_11561,N_11311);
xor U13604 (N_13604,N_6694,N_6142);
xor U13605 (N_13605,N_7403,N_8235);
xor U13606 (N_13606,N_11511,N_11289);
nor U13607 (N_13607,N_9852,N_11527);
xnor U13608 (N_13608,N_6645,N_10543);
xor U13609 (N_13609,N_9709,N_9503);
and U13610 (N_13610,N_7387,N_6126);
and U13611 (N_13611,N_7949,N_6220);
nand U13612 (N_13612,N_8027,N_9540);
nor U13613 (N_13613,N_10220,N_9705);
nor U13614 (N_13614,N_11259,N_7257);
or U13615 (N_13615,N_10066,N_7404);
nor U13616 (N_13616,N_9810,N_6667);
and U13617 (N_13617,N_8090,N_9649);
and U13618 (N_13618,N_6152,N_10246);
or U13619 (N_13619,N_6603,N_11194);
nand U13620 (N_13620,N_10460,N_9909);
nand U13621 (N_13621,N_8138,N_11646);
xor U13622 (N_13622,N_11461,N_10197);
xor U13623 (N_13623,N_9783,N_8503);
xnor U13624 (N_13624,N_10091,N_7655);
or U13625 (N_13625,N_8467,N_9281);
and U13626 (N_13626,N_7000,N_9338);
or U13627 (N_13627,N_9794,N_10180);
nor U13628 (N_13628,N_11052,N_11703);
and U13629 (N_13629,N_10782,N_11393);
xnor U13630 (N_13630,N_6644,N_9999);
nor U13631 (N_13631,N_9583,N_11922);
nand U13632 (N_13632,N_7640,N_7348);
nand U13633 (N_13633,N_10693,N_6131);
nor U13634 (N_13634,N_10242,N_11377);
nor U13635 (N_13635,N_6972,N_10314);
xor U13636 (N_13636,N_6132,N_6636);
and U13637 (N_13637,N_11208,N_7692);
nor U13638 (N_13638,N_11089,N_10957);
or U13639 (N_13639,N_11666,N_9064);
and U13640 (N_13640,N_9451,N_11705);
xor U13641 (N_13641,N_10958,N_8420);
xnor U13642 (N_13642,N_6760,N_10228);
xnor U13643 (N_13643,N_9554,N_11442);
nand U13644 (N_13644,N_9263,N_11178);
nand U13645 (N_13645,N_8793,N_9298);
xnor U13646 (N_13646,N_6928,N_11324);
nor U13647 (N_13647,N_7336,N_9295);
xor U13648 (N_13648,N_6343,N_11653);
nand U13649 (N_13649,N_11562,N_9918);
nand U13650 (N_13650,N_6108,N_6828);
nor U13651 (N_13651,N_11435,N_11123);
nor U13652 (N_13652,N_7825,N_11388);
xor U13653 (N_13653,N_10053,N_10860);
xor U13654 (N_13654,N_10452,N_7636);
xnor U13655 (N_13655,N_11250,N_10288);
or U13656 (N_13656,N_8720,N_6197);
nor U13657 (N_13657,N_10807,N_11870);
nor U13658 (N_13658,N_11665,N_9522);
xor U13659 (N_13659,N_7899,N_7653);
and U13660 (N_13660,N_9374,N_8593);
and U13661 (N_13661,N_9192,N_6877);
xnor U13662 (N_13662,N_11114,N_8394);
or U13663 (N_13663,N_7264,N_6065);
nor U13664 (N_13664,N_11048,N_6445);
nand U13665 (N_13665,N_9404,N_8971);
and U13666 (N_13666,N_9475,N_9772);
or U13667 (N_13667,N_7275,N_6034);
nand U13668 (N_13668,N_10052,N_8437);
xnor U13669 (N_13669,N_9511,N_9022);
or U13670 (N_13670,N_9188,N_6926);
xor U13671 (N_13671,N_6755,N_8640);
xor U13672 (N_13672,N_10112,N_9755);
nor U13673 (N_13673,N_9130,N_10211);
or U13674 (N_13674,N_7997,N_6271);
nand U13675 (N_13675,N_10470,N_8121);
nand U13676 (N_13676,N_10894,N_9044);
or U13677 (N_13677,N_11754,N_7999);
or U13678 (N_13678,N_10720,N_6784);
xnor U13679 (N_13679,N_7101,N_8885);
nor U13680 (N_13680,N_6787,N_10433);
nand U13681 (N_13681,N_10474,N_10916);
and U13682 (N_13682,N_10342,N_7017);
nor U13683 (N_13683,N_11195,N_6719);
xnor U13684 (N_13684,N_7861,N_10160);
nand U13685 (N_13685,N_8812,N_7797);
nor U13686 (N_13686,N_6648,N_6588);
nor U13687 (N_13687,N_9618,N_7391);
nand U13688 (N_13688,N_11477,N_9147);
xnor U13689 (N_13689,N_11074,N_8622);
nand U13690 (N_13690,N_9888,N_9804);
or U13691 (N_13691,N_7890,N_8211);
xnor U13692 (N_13692,N_6568,N_6709);
xnor U13693 (N_13693,N_8302,N_6815);
xor U13694 (N_13694,N_9377,N_10039);
or U13695 (N_13695,N_10663,N_6834);
or U13696 (N_13696,N_9317,N_11398);
or U13697 (N_13697,N_9393,N_10664);
and U13698 (N_13698,N_10422,N_10166);
and U13699 (N_13699,N_11264,N_6844);
and U13700 (N_13700,N_9787,N_10788);
xor U13701 (N_13701,N_7025,N_10710);
nor U13702 (N_13702,N_10962,N_7599);
or U13703 (N_13703,N_11428,N_11878);
and U13704 (N_13704,N_9607,N_10414);
xor U13705 (N_13705,N_10107,N_6990);
and U13706 (N_13706,N_11149,N_6296);
nand U13707 (N_13707,N_6546,N_10999);
nor U13708 (N_13708,N_11567,N_11026);
and U13709 (N_13709,N_7172,N_11832);
or U13710 (N_13710,N_9438,N_11417);
nor U13711 (N_13711,N_7620,N_10108);
and U13712 (N_13712,N_9291,N_7489);
xnor U13713 (N_13713,N_9182,N_8416);
nand U13714 (N_13714,N_10989,N_11138);
xor U13715 (N_13715,N_8451,N_11335);
and U13716 (N_13716,N_9119,N_6316);
or U13717 (N_13717,N_9527,N_8144);
and U13718 (N_13718,N_6758,N_7362);
and U13719 (N_13719,N_7892,N_6576);
or U13720 (N_13720,N_11656,N_6089);
nand U13721 (N_13721,N_6399,N_8902);
nor U13722 (N_13722,N_7113,N_8652);
and U13723 (N_13723,N_9461,N_6249);
nand U13724 (N_13724,N_11356,N_11482);
xor U13725 (N_13725,N_9012,N_6455);
nor U13726 (N_13726,N_7083,N_10410);
xnor U13727 (N_13727,N_8911,N_11306);
and U13728 (N_13728,N_11757,N_11286);
xnor U13729 (N_13729,N_9498,N_10027);
and U13730 (N_13730,N_11845,N_11582);
nor U13731 (N_13731,N_10181,N_8391);
nand U13732 (N_13732,N_7635,N_9831);
xnor U13733 (N_13733,N_11894,N_6826);
nand U13734 (N_13734,N_11080,N_7479);
or U13735 (N_13735,N_7616,N_6862);
and U13736 (N_13736,N_7043,N_10942);
nor U13737 (N_13737,N_11120,N_11813);
nor U13738 (N_13738,N_10144,N_11366);
nand U13739 (N_13739,N_11770,N_8223);
nand U13740 (N_13740,N_11725,N_11099);
nand U13741 (N_13741,N_8282,N_7262);
xor U13742 (N_13742,N_6433,N_9208);
and U13743 (N_13743,N_9845,N_8417);
or U13744 (N_13744,N_10822,N_6831);
nor U13745 (N_13745,N_10031,N_6728);
or U13746 (N_13746,N_8484,N_6273);
nor U13747 (N_13747,N_6858,N_11755);
and U13748 (N_13748,N_9117,N_8062);
xor U13749 (N_13749,N_9354,N_7473);
xor U13750 (N_13750,N_9058,N_9765);
and U13751 (N_13751,N_11192,N_7418);
and U13752 (N_13752,N_8899,N_9072);
or U13753 (N_13753,N_9710,N_9436);
xnor U13754 (N_13754,N_9269,N_7557);
nor U13755 (N_13755,N_6810,N_7398);
or U13756 (N_13756,N_9653,N_8845);
and U13757 (N_13757,N_6275,N_7432);
and U13758 (N_13758,N_8513,N_8792);
xnor U13759 (N_13759,N_8614,N_7145);
and U13760 (N_13760,N_8642,N_6545);
and U13761 (N_13761,N_8889,N_6128);
xnor U13762 (N_13762,N_9777,N_8907);
and U13763 (N_13763,N_9934,N_9199);
or U13764 (N_13764,N_7181,N_11932);
nand U13765 (N_13765,N_9315,N_7758);
and U13766 (N_13766,N_9131,N_7344);
or U13767 (N_13767,N_6339,N_9869);
nand U13768 (N_13768,N_10312,N_11290);
nand U13769 (N_13769,N_11882,N_6270);
and U13770 (N_13770,N_8711,N_6318);
and U13771 (N_13771,N_9249,N_10796);
or U13772 (N_13772,N_11825,N_10583);
nor U13773 (N_13773,N_7240,N_6579);
and U13774 (N_13774,N_11535,N_9226);
xnor U13775 (N_13775,N_9372,N_9037);
or U13776 (N_13776,N_8615,N_10974);
nor U13777 (N_13777,N_9964,N_6208);
nor U13778 (N_13778,N_7266,N_7682);
nand U13779 (N_13779,N_10063,N_7149);
or U13780 (N_13780,N_6357,N_7986);
nor U13781 (N_13781,N_6800,N_10675);
xnor U13782 (N_13782,N_8870,N_7364);
and U13783 (N_13783,N_6717,N_7976);
nor U13784 (N_13784,N_11926,N_7503);
xnor U13785 (N_13785,N_11028,N_8301);
or U13786 (N_13786,N_9229,N_10513);
nor U13787 (N_13787,N_6029,N_11456);
nor U13788 (N_13788,N_8386,N_8855);
nor U13789 (N_13789,N_8535,N_8820);
nor U13790 (N_13790,N_9756,N_7532);
nand U13791 (N_13791,N_6925,N_10369);
nor U13792 (N_13792,N_6845,N_10419);
nor U13793 (N_13793,N_9398,N_11091);
nor U13794 (N_13794,N_6824,N_10893);
nor U13795 (N_13795,N_7923,N_6745);
and U13796 (N_13796,N_7305,N_6418);
nor U13797 (N_13797,N_10287,N_11011);
xor U13798 (N_13798,N_10861,N_6385);
nand U13799 (N_13799,N_7614,N_9010);
or U13800 (N_13800,N_8690,N_11714);
or U13801 (N_13801,N_7256,N_7277);
or U13802 (N_13802,N_9504,N_6642);
or U13803 (N_13803,N_10247,N_10075);
and U13804 (N_13804,N_9561,N_6148);
nor U13805 (N_13805,N_6820,N_9543);
or U13806 (N_13806,N_9021,N_11115);
xor U13807 (N_13807,N_10609,N_6269);
and U13808 (N_13808,N_10716,N_6985);
or U13809 (N_13809,N_6530,N_8232);
and U13810 (N_13810,N_9906,N_7582);
nand U13811 (N_13811,N_7745,N_9184);
xor U13812 (N_13812,N_6011,N_9965);
and U13813 (N_13813,N_8888,N_6793);
xor U13814 (N_13814,N_7378,N_9997);
xnor U13815 (N_13815,N_6622,N_9743);
and U13816 (N_13816,N_7470,N_6120);
and U13817 (N_13817,N_7436,N_9746);
nor U13818 (N_13818,N_8839,N_10641);
xnor U13819 (N_13819,N_7038,N_10106);
or U13820 (N_13820,N_6008,N_8643);
and U13821 (N_13821,N_11334,N_7722);
nor U13822 (N_13822,N_9480,N_8055);
xnor U13823 (N_13823,N_6939,N_11974);
or U13824 (N_13824,N_10726,N_9493);
nor U13825 (N_13825,N_10375,N_9941);
or U13826 (N_13826,N_10049,N_11229);
xnor U13827 (N_13827,N_9993,N_11379);
nor U13828 (N_13828,N_8434,N_8021);
xnor U13829 (N_13829,N_9799,N_6507);
xnor U13830 (N_13830,N_11986,N_9619);
xnor U13831 (N_13831,N_8158,N_7881);
and U13832 (N_13832,N_11760,N_9165);
nand U13833 (N_13833,N_11029,N_9322);
and U13834 (N_13834,N_8598,N_9747);
or U13835 (N_13835,N_11183,N_7279);
or U13836 (N_13836,N_10446,N_10028);
xor U13837 (N_13837,N_6796,N_11176);
and U13838 (N_13838,N_7732,N_9996);
or U13839 (N_13839,N_11125,N_6369);
nor U13840 (N_13840,N_10869,N_11078);
nand U13841 (N_13841,N_8393,N_10413);
nor U13842 (N_13842,N_10343,N_6681);
nand U13843 (N_13843,N_11315,N_6605);
nor U13844 (N_13844,N_7067,N_10756);
nand U13845 (N_13845,N_11041,N_9300);
nand U13846 (N_13846,N_6314,N_8284);
nor U13847 (N_13847,N_10138,N_10952);
or U13848 (N_13848,N_7187,N_11577);
or U13849 (N_13849,N_9005,N_9539);
or U13850 (N_13850,N_9647,N_9541);
nor U13851 (N_13851,N_6802,N_7231);
nor U13852 (N_13852,N_7399,N_6663);
nor U13853 (N_13853,N_10912,N_8730);
xnor U13854 (N_13854,N_11296,N_7898);
xor U13855 (N_13855,N_11016,N_9206);
nand U13856 (N_13856,N_7888,N_10887);
nand U13857 (N_13857,N_8398,N_6848);
or U13858 (N_13858,N_9815,N_10688);
nor U13859 (N_13859,N_8016,N_11359);
xor U13860 (N_13860,N_6650,N_9342);
and U13861 (N_13861,N_7652,N_11017);
or U13862 (N_13862,N_9360,N_9972);
or U13863 (N_13863,N_9484,N_9423);
and U13864 (N_13864,N_7076,N_8618);
xor U13865 (N_13865,N_9518,N_7499);
nor U13866 (N_13866,N_7814,N_10802);
nand U13867 (N_13867,N_7777,N_10200);
nor U13868 (N_13868,N_9268,N_8363);
nand U13869 (N_13869,N_9233,N_9744);
xnor U13870 (N_13870,N_9340,N_10837);
xnor U13871 (N_13871,N_7872,N_9205);
or U13872 (N_13872,N_11680,N_7847);
xnor U13873 (N_13873,N_6424,N_9530);
or U13874 (N_13874,N_10378,N_10381);
nand U13875 (N_13875,N_6329,N_11007);
nand U13876 (N_13876,N_7540,N_6772);
xnor U13877 (N_13877,N_6591,N_10169);
nor U13878 (N_13878,N_11031,N_7039);
and U13879 (N_13879,N_11127,N_10240);
or U13880 (N_13880,N_8383,N_11202);
and U13881 (N_13881,N_9059,N_8217);
nor U13882 (N_13882,N_10125,N_6634);
xnor U13883 (N_13883,N_9238,N_10810);
or U13884 (N_13884,N_8702,N_10449);
nor U13885 (N_13885,N_6030,N_10133);
and U13886 (N_13886,N_7269,N_9766);
nand U13887 (N_13887,N_11919,N_11789);
and U13888 (N_13888,N_11811,N_6819);
or U13889 (N_13889,N_10722,N_11960);
and U13890 (N_13890,N_8237,N_11538);
and U13891 (N_13891,N_6592,N_6267);
and U13892 (N_13892,N_9844,N_8135);
nand U13893 (N_13893,N_9335,N_9660);
or U13894 (N_13894,N_6946,N_7724);
xor U13895 (N_13895,N_9103,N_6254);
or U13896 (N_13896,N_8311,N_6918);
nor U13897 (N_13897,N_8065,N_8174);
nor U13898 (N_13898,N_10092,N_8656);
and U13899 (N_13899,N_10265,N_8922);
xor U13900 (N_13900,N_8429,N_11008);
and U13901 (N_13901,N_11752,N_7241);
or U13902 (N_13902,N_10290,N_6947);
nand U13903 (N_13903,N_7315,N_10438);
and U13904 (N_13904,N_9525,N_10023);
xor U13905 (N_13905,N_6277,N_8713);
nor U13906 (N_13906,N_8600,N_9375);
or U13907 (N_13907,N_11189,N_9094);
and U13908 (N_13908,N_10825,N_11111);
xnor U13909 (N_13909,N_6194,N_8457);
nor U13910 (N_13910,N_8764,N_11839);
or U13911 (N_13911,N_10551,N_6971);
xnor U13912 (N_13912,N_9096,N_6823);
nand U13913 (N_13913,N_6869,N_9512);
or U13914 (N_13914,N_6904,N_6157);
nor U13915 (N_13915,N_8512,N_7723);
nor U13916 (N_13916,N_9231,N_8826);
nand U13917 (N_13917,N_9667,N_8137);
xnor U13918 (N_13918,N_7010,N_11935);
or U13919 (N_13919,N_6374,N_7355);
nand U13920 (N_13920,N_11568,N_11174);
and U13921 (N_13921,N_8608,N_7980);
or U13922 (N_13922,N_9470,N_11543);
and U13923 (N_13923,N_8893,N_6454);
nor U13924 (N_13924,N_6978,N_7565);
or U13925 (N_13925,N_9455,N_7184);
and U13926 (N_13926,N_11305,N_9631);
or U13927 (N_13927,N_10115,N_11584);
xor U13928 (N_13928,N_6311,N_7504);
or U13929 (N_13929,N_8465,N_11989);
xor U13930 (N_13930,N_6907,N_11145);
and U13931 (N_13931,N_8565,N_8925);
nor U13932 (N_13932,N_9038,N_6450);
nand U13933 (N_13933,N_9181,N_11404);
nor U13934 (N_13934,N_7610,N_8878);
nand U13935 (N_13935,N_7159,N_9065);
xnor U13936 (N_13936,N_11598,N_10510);
nand U13937 (N_13937,N_10251,N_6104);
xor U13938 (N_13938,N_10149,N_7604);
and U13939 (N_13939,N_7313,N_9359);
xnor U13940 (N_13940,N_9203,N_11242);
nand U13941 (N_13941,N_9152,N_7026);
xnor U13942 (N_13942,N_10129,N_10185);
or U13943 (N_13943,N_10790,N_10740);
or U13944 (N_13944,N_10187,N_6328);
or U13945 (N_13945,N_10012,N_9565);
nor U13946 (N_13946,N_6838,N_8532);
and U13947 (N_13947,N_10163,N_10488);
and U13948 (N_13948,N_6649,N_9446);
xor U13949 (N_13949,N_9576,N_8570);
or U13950 (N_13950,N_6866,N_6351);
and U13951 (N_13951,N_10054,N_8561);
or U13952 (N_13952,N_11824,N_7650);
nand U13953 (N_13953,N_10404,N_10132);
and U13954 (N_13954,N_6047,N_10439);
or U13955 (N_13955,N_11525,N_11170);
nand U13956 (N_13956,N_10173,N_6167);
nor U13957 (N_13957,N_9448,N_11947);
nand U13958 (N_13958,N_10659,N_8607);
and U13959 (N_13959,N_11179,N_6474);
and U13960 (N_13960,N_8805,N_11357);
xnor U13961 (N_13961,N_6485,N_9383);
nor U13962 (N_13962,N_8807,N_10977);
or U13963 (N_13963,N_9082,N_11282);
nand U13964 (N_13964,N_8067,N_6421);
nor U13965 (N_13965,N_9081,N_7686);
and U13966 (N_13966,N_7135,N_10245);
or U13967 (N_13967,N_10524,N_6892);
and U13968 (N_13968,N_9699,N_11632);
xnor U13969 (N_13969,N_9958,N_8167);
and U13970 (N_13970,N_11113,N_6524);
xnor U13971 (N_13971,N_8639,N_11520);
xor U13972 (N_13972,N_10881,N_11795);
or U13973 (N_13973,N_8606,N_11233);
xnor U13974 (N_13974,N_8063,N_7756);
nor U13975 (N_13975,N_7245,N_8203);
xor U13976 (N_13976,N_8374,N_7632);
nand U13977 (N_13977,N_10315,N_6413);
nand U13978 (N_13978,N_11536,N_10151);
nand U13979 (N_13979,N_8545,N_6347);
or U13980 (N_13980,N_8101,N_6230);
and U13981 (N_13981,N_7867,N_11056);
nor U13982 (N_13982,N_8099,N_10748);
and U13983 (N_13983,N_6017,N_11153);
nand U13984 (N_13984,N_10642,N_6191);
xor U13985 (N_13985,N_11806,N_6861);
xnor U13986 (N_13986,N_7488,N_9672);
xor U13987 (N_13987,N_6827,N_9896);
nand U13988 (N_13988,N_8214,N_10172);
nand U13989 (N_13989,N_7014,N_11652);
and U13990 (N_13990,N_11958,N_11209);
or U13991 (N_13991,N_10340,N_7848);
or U13992 (N_13992,N_8511,N_10885);
nand U13993 (N_13993,N_11915,N_7133);
and U13994 (N_13994,N_9025,N_7554);
nand U13995 (N_13995,N_6573,N_11676);
nor U13996 (N_13996,N_10459,N_11067);
nor U13997 (N_13997,N_10389,N_7070);
or U13998 (N_13998,N_7812,N_9648);
or U13999 (N_13999,N_7037,N_7813);
nor U14000 (N_14000,N_7029,N_10100);
nor U14001 (N_14001,N_6232,N_10109);
and U14002 (N_14002,N_11450,N_7246);
and U14003 (N_14003,N_7179,N_8883);
nor U14004 (N_14004,N_9564,N_7644);
nor U14005 (N_14005,N_7866,N_8729);
xor U14006 (N_14006,N_7377,N_6130);
or U14007 (N_14007,N_10203,N_9624);
and U14008 (N_14008,N_7013,N_9039);
nor U14009 (N_14009,N_7117,N_8438);
xor U14010 (N_14010,N_8689,N_11001);
or U14011 (N_14011,N_10775,N_9886);
nand U14012 (N_14012,N_11217,N_7371);
xor U14013 (N_14013,N_9731,N_9433);
and U14014 (N_14014,N_10354,N_10199);
xnor U14015 (N_14015,N_6437,N_8344);
xor U14016 (N_14016,N_10619,N_10295);
nor U14017 (N_14017,N_7361,N_10596);
or U14018 (N_14018,N_10933,N_10733);
xnor U14019 (N_14019,N_9349,N_8283);
or U14020 (N_14020,N_8523,N_8924);
and U14021 (N_14021,N_6492,N_7228);
or U14022 (N_14022,N_11716,N_7099);
and U14023 (N_14023,N_10766,N_11589);
or U14024 (N_14024,N_10326,N_9935);
or U14025 (N_14025,N_11355,N_6272);
and U14026 (N_14026,N_10184,N_6741);
nor U14027 (N_14027,N_7725,N_7465);
and U14028 (N_14028,N_9466,N_10298);
xor U14029 (N_14029,N_8819,N_10754);
or U14030 (N_14030,N_8734,N_10044);
xor U14031 (N_14031,N_6412,N_10178);
nor U14032 (N_14032,N_9048,N_10236);
nand U14033 (N_14033,N_9155,N_8783);
xor U14034 (N_14034,N_6541,N_7708);
nor U14035 (N_14035,N_9213,N_8831);
nand U14036 (N_14036,N_9592,N_11731);
nand U14037 (N_14037,N_8934,N_6697);
nor U14038 (N_14038,N_10024,N_11797);
nand U14039 (N_14039,N_11135,N_7087);
xor U14040 (N_14040,N_9739,N_11387);
and U14041 (N_14041,N_11383,N_6999);
nand U14042 (N_14042,N_6887,N_8521);
xor U14043 (N_14043,N_7046,N_6635);
nor U14044 (N_14044,N_10874,N_7407);
xor U14045 (N_14045,N_7177,N_11792);
or U14046 (N_14046,N_7615,N_8737);
or U14047 (N_14047,N_6196,N_6806);
xnor U14048 (N_14048,N_8721,N_10559);
nand U14049 (N_14049,N_8278,N_9580);
nand U14050 (N_14050,N_7080,N_8333);
nand U14051 (N_14051,N_8507,N_9134);
or U14052 (N_14052,N_7110,N_10217);
nor U14053 (N_14053,N_9929,N_8789);
nor U14054 (N_14054,N_10175,N_6916);
xnor U14055 (N_14055,N_9696,N_8147);
nor U14056 (N_14056,N_6156,N_9827);
xnor U14057 (N_14057,N_10014,N_8694);
and U14058 (N_14058,N_11774,N_11316);
nand U14059 (N_14059,N_11923,N_7851);
or U14060 (N_14060,N_11554,N_10316);
or U14061 (N_14061,N_10473,N_8305);
or U14062 (N_14062,N_11790,N_8869);
nand U14063 (N_14063,N_11431,N_7141);
xnor U14064 (N_14064,N_6028,N_8900);
nor U14065 (N_14065,N_7651,N_9978);
nand U14066 (N_14066,N_9245,N_9177);
xnor U14067 (N_14067,N_9120,N_10156);
nand U14068 (N_14068,N_6407,N_11328);
xor U14069 (N_14069,N_7401,N_6051);
xor U14070 (N_14070,N_8972,N_10988);
or U14071 (N_14071,N_11488,N_6419);
nor U14072 (N_14072,N_10723,N_8709);
xor U14073 (N_14073,N_6473,N_8486);
xnor U14074 (N_14074,N_8660,N_6991);
nand U14075 (N_14075,N_6201,N_9575);
and U14076 (N_14076,N_8026,N_10949);
or U14077 (N_14077,N_11515,N_9585);
nor U14078 (N_14078,N_8334,N_7935);
and U14079 (N_14079,N_8510,N_7389);
nor U14080 (N_14080,N_7075,N_6716);
and U14081 (N_14081,N_9823,N_9623);
and U14082 (N_14082,N_11107,N_9524);
nor U14083 (N_14083,N_10703,N_7160);
nand U14084 (N_14084,N_10907,N_11766);
nand U14085 (N_14085,N_8321,N_7597);
xor U14086 (N_14086,N_8688,N_9718);
nand U14087 (N_14087,N_8681,N_11942);
xor U14088 (N_14088,N_11401,N_10800);
xnor U14089 (N_14089,N_10545,N_7707);
and U14090 (N_14090,N_7064,N_11968);
nor U14091 (N_14091,N_7290,N_6380);
nand U14092 (N_14092,N_8295,N_9162);
or U14093 (N_14093,N_9121,N_11292);
nor U14094 (N_14094,N_8083,N_8824);
nor U14095 (N_14095,N_7992,N_9881);
xnor U14096 (N_14096,N_8264,N_6565);
or U14097 (N_14097,N_9379,N_11638);
nor U14098 (N_14098,N_9251,N_11154);
and U14099 (N_14099,N_10097,N_11833);
xor U14100 (N_14100,N_10209,N_7955);
xor U14101 (N_14101,N_9621,N_8537);
and U14102 (N_14102,N_6689,N_9495);
nand U14103 (N_14103,N_11350,N_11876);
xor U14104 (N_14104,N_8753,N_9798);
nand U14105 (N_14105,N_6460,N_6700);
xor U14106 (N_14106,N_11542,N_7698);
xnor U14107 (N_14107,N_9256,N_8483);
nand U14108 (N_14108,N_6640,N_7619);
nor U14109 (N_14109,N_8401,N_7618);
nand U14110 (N_14110,N_6101,N_8123);
nand U14111 (N_14111,N_10767,N_8248);
xnor U14112 (N_14112,N_9760,N_6376);
and U14113 (N_14113,N_10972,N_8646);
nand U14114 (N_14114,N_11406,N_8024);
nor U14115 (N_14115,N_8107,N_11416);
nand U14116 (N_14116,N_10685,N_10951);
and U14117 (N_14117,N_6325,N_7107);
and U14118 (N_14118,N_7323,N_7852);
xor U14119 (N_14119,N_10892,N_8994);
and U14120 (N_14120,N_8230,N_7180);
and U14121 (N_14121,N_9684,N_6417);
and U14122 (N_14122,N_9320,N_8973);
and U14123 (N_14123,N_8414,N_6522);
nor U14124 (N_14124,N_9421,N_6804);
or U14125 (N_14125,N_11551,N_9507);
xnor U14126 (N_14126,N_11533,N_6995);
or U14127 (N_14127,N_11610,N_8127);
and U14128 (N_14128,N_10512,N_7974);
xnor U14129 (N_14129,N_8289,N_9821);
nor U14130 (N_14130,N_8136,N_8118);
nor U14131 (N_14131,N_7009,N_8738);
or U14132 (N_14132,N_11967,N_6543);
nor U14133 (N_14133,N_8851,N_10531);
nand U14134 (N_14134,N_9054,N_11385);
nand U14135 (N_14135,N_10877,N_6790);
nor U14136 (N_14136,N_7774,N_10769);
and U14137 (N_14137,N_10202,N_7791);
nand U14138 (N_14138,N_10319,N_7495);
and U14139 (N_14139,N_9578,N_7702);
or U14140 (N_14140,N_8187,N_7081);
nor U14141 (N_14141,N_11579,N_10153);
nor U14142 (N_14142,N_11826,N_6669);
nand U14143 (N_14143,N_11869,N_9264);
or U14144 (N_14144,N_10411,N_11917);
or U14145 (N_14145,N_7174,N_6370);
and U14146 (N_14146,N_6367,N_7242);
xor U14147 (N_14147,N_8335,N_10941);
xnor U14148 (N_14148,N_7370,N_11424);
and U14149 (N_14149,N_7826,N_9986);
xnor U14150 (N_14150,N_8786,N_10920);
and U14151 (N_14151,N_11484,N_10606);
or U14152 (N_14152,N_7464,N_9091);
nand U14153 (N_14153,N_8473,N_8542);
and U14154 (N_14154,N_6562,N_10088);
or U14155 (N_14155,N_9157,N_10915);
and U14156 (N_14156,N_11105,N_8314);
and U14157 (N_14157,N_10897,N_7828);
or U14158 (N_14158,N_8865,N_9994);
xnor U14159 (N_14159,N_10234,N_7882);
nor U14160 (N_14160,N_10947,N_8228);
nor U14161 (N_14161,N_11891,N_6175);
nand U14162 (N_14162,N_7953,N_8589);
nor U14163 (N_14163,N_7451,N_6245);
xor U14164 (N_14164,N_8126,N_7679);
and U14165 (N_14165,N_11738,N_9839);
nand U14166 (N_14166,N_11035,N_10953);
or U14167 (N_14167,N_6000,N_6659);
nor U14168 (N_14168,N_9068,N_9603);
nand U14169 (N_14169,N_11575,N_10043);
nand U14170 (N_14170,N_9600,N_9105);
nor U14171 (N_14171,N_7406,N_9078);
nor U14172 (N_14172,N_11805,N_7897);
xnor U14173 (N_14173,N_6354,N_8009);
nand U14174 (N_14174,N_6022,N_7248);
and U14175 (N_14175,N_9261,N_11251);
xnor U14176 (N_14176,N_11902,N_10614);
nor U14177 (N_14177,N_11049,N_7215);
nand U14178 (N_14178,N_10386,N_10530);
and U14179 (N_14179,N_6677,N_6026);
nor U14180 (N_14180,N_8759,N_7105);
nand U14181 (N_14181,N_6363,N_6587);
and U14182 (N_14182,N_7837,N_6317);
xor U14183 (N_14183,N_10768,N_11890);
or U14184 (N_14184,N_9957,N_6244);
nand U14185 (N_14185,N_8722,N_11037);
or U14186 (N_14186,N_11601,N_8276);
nor U14187 (N_14187,N_6151,N_7739);
xor U14188 (N_14188,N_10042,N_10399);
and U14189 (N_14189,N_7205,N_10182);
or U14190 (N_14190,N_9418,N_10582);
nor U14191 (N_14191,N_9041,N_9447);
xnor U14192 (N_14192,N_9489,N_7993);
and U14193 (N_14193,N_7124,N_9695);
nor U14194 (N_14194,N_6129,N_9434);
xnor U14195 (N_14195,N_6656,N_9380);
xor U14196 (N_14196,N_6422,N_8119);
nand U14197 (N_14197,N_11976,N_9305);
xor U14198 (N_14198,N_9257,N_10542);
and U14199 (N_14199,N_10819,N_8431);
xnor U14200 (N_14200,N_6583,N_7868);
nor U14201 (N_14201,N_7408,N_7200);
xor U14202 (N_14202,N_6739,N_9348);
or U14203 (N_14203,N_8588,N_11262);
xnor U14204 (N_14204,N_9087,N_10472);
nand U14205 (N_14205,N_7793,N_10898);
nand U14206 (N_14206,N_7507,N_10795);
and U14207 (N_14207,N_7833,N_7842);
nor U14208 (N_14208,N_8265,N_9032);
nor U14209 (N_14209,N_11464,N_6439);
or U14210 (N_14210,N_11144,N_7737);
nand U14211 (N_14211,N_9053,N_8691);
or U14212 (N_14212,N_11512,N_11707);
nand U14213 (N_14213,N_6534,N_9435);
and U14214 (N_14214,N_11686,N_11877);
xnor U14215 (N_14215,N_11021,N_8320);
nand U14216 (N_14216,N_8443,N_9668);
nand U14217 (N_14217,N_10001,N_11627);
nand U14218 (N_14218,N_10780,N_9200);
and U14219 (N_14219,N_11340,N_10372);
or U14220 (N_14220,N_7471,N_7072);
and U14221 (N_14221,N_6446,N_11906);
xor U14222 (N_14222,N_11168,N_8208);
and U14223 (N_14223,N_9506,N_8862);
nand U14224 (N_14224,N_8648,N_10760);
and U14225 (N_14225,N_10794,N_7086);
nand U14226 (N_14226,N_10141,N_10465);
nand U14227 (N_14227,N_10993,N_6685);
or U14228 (N_14228,N_10762,N_11508);
nand U14229 (N_14229,N_9532,N_8977);
and U14230 (N_14230,N_7230,N_8525);
and U14231 (N_14231,N_6706,N_9186);
xor U14232 (N_14232,N_6623,N_7932);
nor U14233 (N_14233,N_11687,N_6989);
and U14234 (N_14234,N_7862,N_9063);
nand U14235 (N_14235,N_8951,N_9627);
and U14236 (N_14236,N_11995,N_7345);
or U14237 (N_14237,N_9586,N_6393);
xnor U14238 (N_14238,N_6805,N_6281);
nand U14239 (N_14239,N_7990,N_9144);
and U14240 (N_14240,N_8463,N_9472);
nor U14241 (N_14241,N_7563,N_9202);
xnor U14242 (N_14242,N_6983,N_9003);
nor U14243 (N_14243,N_8572,N_10493);
xor U14244 (N_14244,N_9940,N_11327);
nor U14245 (N_14245,N_8822,N_8166);
nor U14246 (N_14246,N_8356,N_6038);
xor U14247 (N_14247,N_6513,N_8563);
nand U14248 (N_14248,N_8343,N_9331);
nor U14249 (N_14249,N_11830,N_10622);
nor U14250 (N_14250,N_11730,N_8712);
and U14251 (N_14251,N_9296,N_11241);
and U14252 (N_14252,N_8661,N_10499);
nand U14253 (N_14253,N_8941,N_7645);
nor U14254 (N_14254,N_6691,N_6698);
nand U14255 (N_14255,N_11063,N_7676);
xnor U14256 (N_14256,N_11875,N_7351);
and U14257 (N_14257,N_7321,N_9939);
and U14258 (N_14258,N_7922,N_9274);
nand U14259 (N_14259,N_8145,N_11171);
and U14260 (N_14260,N_9254,N_9015);
xor U14261 (N_14261,N_10759,N_10126);
nand U14262 (N_14262,N_9680,N_6769);
nand U14263 (N_14263,N_7238,N_11186);
or U14264 (N_14264,N_6027,N_11231);
nand U14265 (N_14265,N_10550,N_6250);
xor U14266 (N_14266,N_6390,N_11207);
xnor U14267 (N_14267,N_7265,N_9168);
or U14268 (N_14268,N_6864,N_6003);
nor U14269 (N_14269,N_6115,N_6846);
or U14270 (N_14270,N_6571,N_8495);
or U14271 (N_14271,N_7627,N_8195);
and U14272 (N_14272,N_8191,N_7508);
and U14273 (N_14273,N_9846,N_9384);
or U14274 (N_14274,N_10986,N_11304);
nand U14275 (N_14275,N_11003,N_11615);
and U14276 (N_14276,N_8630,N_9908);
or U14277 (N_14277,N_9691,N_6942);
and U14278 (N_14278,N_11256,N_9468);
nor U14279 (N_14279,N_7051,N_8992);
nor U14280 (N_14280,N_9243,N_10911);
nand U14281 (N_14281,N_9762,N_9463);
or U14282 (N_14282,N_7605,N_10650);
nor U14283 (N_14283,N_7529,N_7951);
or U14284 (N_14284,N_11519,N_7103);
or U14285 (N_14285,N_11724,N_7301);
nor U14286 (N_14286,N_10161,N_10724);
nor U14287 (N_14287,N_9926,N_7677);
nor U14288 (N_14288,N_8172,N_8077);
and U14289 (N_14289,N_6589,N_6395);
nand U14290 (N_14290,N_10571,N_11992);
and U14291 (N_14291,N_7982,N_11337);
nand U14292 (N_14292,N_11921,N_8448);
nand U14293 (N_14293,N_11299,N_11588);
nand U14294 (N_14294,N_9364,N_11455);
or U14295 (N_14295,N_7247,N_10677);
nor U14296 (N_14296,N_6531,N_11372);
xnor U14297 (N_14297,N_8813,N_7659);
nand U14298 (N_14298,N_8547,N_10520);
xnor U14299 (N_14299,N_6294,N_10763);
and U14300 (N_14300,N_7536,N_11576);
or U14301 (N_14301,N_6675,N_8775);
nand U14302 (N_14302,N_8945,N_9625);
and U14303 (N_14303,N_8000,N_8440);
or U14304 (N_14304,N_9046,N_10210);
nand U14305 (N_14305,N_11970,N_9006);
nor U14306 (N_14306,N_9748,N_6392);
xnor U14307 (N_14307,N_9141,N_10356);
nand U14308 (N_14308,N_6246,N_8731);
or U14309 (N_14309,N_9275,N_8493);
xnor U14310 (N_14310,N_10271,N_8029);
nand U14311 (N_14311,N_10346,N_8678);
nor U14312 (N_14312,N_7972,N_9634);
or U14313 (N_14313,N_10585,N_9106);
nand U14314 (N_14314,N_8927,N_8052);
nor U14315 (N_14315,N_9240,N_10851);
and U14316 (N_14316,N_10146,N_11747);
or U14317 (N_14317,N_7216,N_7977);
or U14318 (N_14318,N_8882,N_11329);
xnor U14319 (N_14319,N_11371,N_8433);
nor U14320 (N_14320,N_7093,N_8967);
nor U14321 (N_14321,N_9497,N_8479);
and U14322 (N_14322,N_8768,N_7544);
and U14323 (N_14323,N_7880,N_11695);
or U14324 (N_14324,N_6268,N_11859);
or U14325 (N_14325,N_6778,N_10239);
nand U14326 (N_14326,N_7126,N_9837);
xor U14327 (N_14327,N_7525,N_6009);
nand U14328 (N_14328,N_10721,N_7649);
nor U14329 (N_14329,N_8978,N_7251);
and U14330 (N_14330,N_7688,N_7819);
nor U14331 (N_14331,N_11126,N_10478);
xnor U14332 (N_14332,N_10725,N_11013);
and U14333 (N_14333,N_7271,N_11073);
nand U14334 (N_14334,N_6992,N_9676);
and U14335 (N_14335,N_6228,N_7665);
and U14336 (N_14336,N_8996,N_11740);
xnor U14337 (N_14337,N_11485,N_9386);
nand U14338 (N_14338,N_7572,N_11266);
and U14339 (N_14339,N_8428,N_8527);
and U14340 (N_14340,N_8435,N_8385);
xor U14341 (N_14341,N_9587,N_8677);
xnor U14342 (N_14342,N_6096,N_6448);
xor U14343 (N_14343,N_6106,N_11313);
xor U14344 (N_14344,N_11709,N_9324);
nand U14345 (N_14345,N_10256,N_11198);
and U14346 (N_14346,N_7222,N_9216);
nand U14347 (N_14347,N_10096,N_8159);
nand U14348 (N_14348,N_11454,N_9716);
and U14349 (N_14349,N_8348,N_10111);
and U14350 (N_14350,N_11959,N_10546);
or U14351 (N_14351,N_9991,N_6377);
or U14352 (N_14352,N_10442,N_7522);
nand U14353 (N_14353,N_10824,N_11221);
and U14354 (N_14354,N_6699,N_9761);
or U14355 (N_14355,N_10366,N_7468);
xnor U14356 (N_14356,N_8073,N_7129);
nor U14357 (N_14357,N_6922,N_6765);
xor U14358 (N_14358,N_8637,N_10332);
nor U14359 (N_14359,N_8286,N_8478);
or U14360 (N_14360,N_6366,N_11322);
nand U14361 (N_14361,N_7761,N_9197);
nand U14362 (N_14362,N_8332,N_10954);
xnor U14363 (N_14363,N_7799,N_11993);
xor U14364 (N_14364,N_9017,N_10325);
nand U14365 (N_14365,N_6043,N_9698);
nand U14366 (N_14366,N_7646,N_7114);
and U14367 (N_14367,N_9608,N_6466);
xnor U14368 (N_14368,N_9642,N_9167);
and U14369 (N_14369,N_9487,N_7957);
nor U14370 (N_14370,N_7821,N_7224);
nor U14371 (N_14371,N_6569,N_11420);
nor U14372 (N_14372,N_10603,N_9288);
nor U14373 (N_14373,N_10784,N_10301);
xnor U14374 (N_14374,N_9358,N_11191);
nand U14375 (N_14375,N_11815,N_11124);
and U14376 (N_14376,N_8244,N_7585);
and U14377 (N_14377,N_11024,N_10847);
nand U14378 (N_14378,N_8359,N_11920);
nor U14379 (N_14379,N_10170,N_10704);
xnor U14380 (N_14380,N_9904,N_8647);
nand U14381 (N_14381,N_7633,N_8829);
and U14382 (N_14382,N_9344,N_6168);
and U14383 (N_14383,N_6200,N_10868);
xnor U14384 (N_14384,N_7967,N_7041);
and U14385 (N_14385,N_11979,N_11473);
nor U14386 (N_14386,N_9270,N_10555);
nand U14387 (N_14387,N_10667,N_6770);
nand U14388 (N_14388,N_11465,N_6899);
nor U14389 (N_14389,N_6842,N_10889);
nand U14390 (N_14390,N_11684,N_6560);
or U14391 (N_14391,N_6123,N_10224);
or U14392 (N_14392,N_11867,N_11546);
and U14393 (N_14393,N_11966,N_6508);
xnor U14394 (N_14394,N_7578,N_8115);
nand U14395 (N_14395,N_8763,N_10741);
nand U14396 (N_14396,N_8179,N_7466);
nor U14397 (N_14397,N_6505,N_9500);
and U14398 (N_14398,N_7416,N_8419);
nor U14399 (N_14399,N_8748,N_10362);
xnor U14400 (N_14400,N_7074,N_11205);
and U14401 (N_14401,N_7926,N_7810);
nand U14402 (N_14402,N_9767,N_11336);
xor U14403 (N_14403,N_10308,N_9917);
and U14404 (N_14404,N_9854,N_9803);
and U14405 (N_14405,N_9027,N_8307);
nor U14406 (N_14406,N_7666,N_6321);
or U14407 (N_14407,N_8327,N_9679);
nand U14408 (N_14408,N_9629,N_10662);
or U14409 (N_14409,N_8381,N_6585);
nand U14410 (N_14410,N_9635,N_11943);
nor U14411 (N_14411,N_11635,N_9802);
nand U14412 (N_14412,N_8964,N_10538);
nor U14413 (N_14413,N_9474,N_7663);
and U14414 (N_14414,N_10745,N_6186);
and U14415 (N_14415,N_11957,N_11050);
nor U14416 (N_14416,N_10539,N_8247);
xor U14417 (N_14417,N_7030,N_10261);
xnor U14418 (N_14418,N_11631,N_9776);
xnor U14419 (N_14419,N_11384,N_8019);
xnor U14420 (N_14420,N_8799,N_10747);
nand U14421 (N_14421,N_10191,N_9159);
nor U14422 (N_14422,N_10649,N_11771);
or U14423 (N_14423,N_8251,N_10646);
xnor U14424 (N_14424,N_7958,N_9146);
nor U14425 (N_14425,N_9369,N_8259);
or U14426 (N_14426,N_6526,N_10752);
or U14427 (N_14427,N_9486,N_7581);
xnor U14428 (N_14428,N_10964,N_6404);
xnor U14429 (N_14429,N_9617,N_9284);
or U14430 (N_14430,N_10594,N_9809);
nor U14431 (N_14431,N_10518,N_7274);
nand U14432 (N_14432,N_8288,N_6274);
nand U14433 (N_14433,N_11619,N_11614);
or U14434 (N_14434,N_8188,N_10233);
nand U14435 (N_14435,N_7984,N_7524);
nand U14436 (N_14436,N_11661,N_9185);
or U14437 (N_14437,N_11514,N_11756);
nor U14438 (N_14438,N_9193,N_7052);
nand U14439 (N_14439,N_9376,N_11436);
nand U14440 (N_14440,N_8178,N_8946);
and U14441 (N_14441,N_11605,N_10155);
nand U14442 (N_14442,N_8003,N_6044);
and U14443 (N_14443,N_8707,N_9201);
or U14444 (N_14444,N_10273,N_8892);
and U14445 (N_14445,N_8963,N_9034);
or U14446 (N_14446,N_9416,N_11712);
or U14447 (N_14447,N_10194,N_9132);
or U14448 (N_14448,N_6646,N_11566);
and U14449 (N_14449,N_6209,N_6295);
xor U14450 (N_14450,N_10793,N_7558);
xor U14451 (N_14451,N_7354,N_8904);
nand U14452 (N_14452,N_9905,N_8411);
or U14453 (N_14453,N_8556,N_11840);
or U14454 (N_14454,N_11106,N_11274);
nor U14455 (N_14455,N_11594,N_10525);
and U14456 (N_14456,N_11411,N_9614);
nor U14457 (N_14457,N_9847,N_6924);
xnor U14458 (N_14458,N_8268,N_11660);
and U14459 (N_14459,N_9825,N_6540);
nor U14460 (N_14460,N_9690,N_11612);
and U14461 (N_14461,N_9085,N_7090);
nand U14462 (N_14462,N_8409,N_7430);
nor U14463 (N_14463,N_10647,N_9350);
and U14464 (N_14464,N_8128,N_10575);
nor U14465 (N_14465,N_8488,N_9652);
and U14466 (N_14466,N_10458,N_6902);
xor U14467 (N_14467,N_10654,N_10982);
and U14468 (N_14468,N_6057,N_10669);
nand U14469 (N_14469,N_11187,N_8193);
and U14470 (N_14470,N_8219,N_6113);
and U14471 (N_14471,N_7353,N_10966);
or U14472 (N_14472,N_6657,N_7750);
xnor U14473 (N_14473,N_8550,N_9107);
and U14474 (N_14474,N_9944,N_7474);
or U14475 (N_14475,N_6851,N_11718);
xor U14476 (N_14476,N_9797,N_11502);
nand U14477 (N_14477,N_10201,N_6405);
nor U14478 (N_14478,N_7840,N_6532);
nand U14479 (N_14479,N_7596,N_6116);
nor U14480 (N_14480,N_10134,N_11403);
nand U14481 (N_14481,N_6715,N_11886);
nor U14482 (N_14482,N_9641,N_7040);
and U14483 (N_14483,N_11255,N_8560);
nor U14484 (N_14484,N_7132,N_9492);
xnor U14485 (N_14485,N_10079,N_10345);
nand U14486 (N_14486,N_7098,N_10904);
or U14487 (N_14487,N_6551,N_9347);
xor U14488 (N_14488,N_6238,N_10983);
or U14489 (N_14489,N_6891,N_8061);
xor U14490 (N_14490,N_6039,N_10864);
nor U14491 (N_14491,N_7593,N_11184);
and U14492 (N_14492,N_6614,N_11778);
and U14493 (N_14493,N_10848,N_10598);
nor U14494 (N_14494,N_10213,N_10491);
or U14495 (N_14495,N_8373,N_11529);
xor U14496 (N_14496,N_10409,N_7939);
and U14497 (N_14497,N_10644,N_6158);
and U14498 (N_14498,N_8626,N_8045);
and U14499 (N_14499,N_6090,N_6653);
or U14500 (N_14500,N_11429,N_8157);
and U14501 (N_14501,N_6938,N_7386);
nand U14502 (N_14502,N_11861,N_7447);
or U14503 (N_14503,N_7553,N_8621);
or U14504 (N_14504,N_7142,N_9422);
or U14505 (N_14505,N_7170,N_6906);
nor U14506 (N_14506,N_11188,N_8584);
nor U14507 (N_14507,N_9735,N_8506);
and U14508 (N_14508,N_6705,N_7689);
nand U14509 (N_14509,N_8952,N_7482);
nand U14510 (N_14510,N_11323,N_10123);
xor U14511 (N_14511,N_9278,N_10803);
nand U14512 (N_14512,N_10421,N_10017);
and U14513 (N_14513,N_7674,N_6074);
or U14514 (N_14514,N_10009,N_8644);
nand U14515 (N_14515,N_6488,N_7588);
and U14516 (N_14516,N_7446,N_7063);
nand U14517 (N_14517,N_9412,N_10113);
nand U14518 (N_14518,N_10434,N_8509);
and U14519 (N_14519,N_10652,N_8842);
or U14520 (N_14520,N_6352,N_10336);
nor U14521 (N_14521,N_11624,N_8072);
or U14522 (N_14522,N_7714,N_11422);
xnor U14523 (N_14523,N_11433,N_9584);
and U14524 (N_14524,N_9389,N_8089);
xnor U14525 (N_14525,N_8909,N_8921);
nand U14526 (N_14526,N_10253,N_10552);
nand U14527 (N_14527,N_6817,N_9822);
nand U14528 (N_14528,N_6429,N_8051);
or U14529 (N_14529,N_6768,N_11453);
nor U14530 (N_14530,N_8751,N_7243);
nor U14531 (N_14531,N_11397,N_10204);
xor U14532 (N_14532,N_10310,N_8961);
xnor U14533 (N_14533,N_10742,N_11872);
xnor U14534 (N_14534,N_7158,N_7369);
and U14535 (N_14535,N_8186,N_10590);
nand U14536 (N_14536,N_7695,N_6161);
xnor U14537 (N_14537,N_10817,N_8182);
nor U14538 (N_14538,N_6447,N_9643);
or U14539 (N_14539,N_11953,N_7062);
and U14540 (N_14540,N_9385,N_10672);
or U14541 (N_14541,N_10888,N_7715);
and U14542 (N_14542,N_6872,N_6031);
xnor U14543 (N_14543,N_10876,N_9806);
xor U14544 (N_14544,N_7530,N_11490);
and U14545 (N_14545,N_10152,N_10168);
nand U14546 (N_14546,N_8908,N_10177);
and U14547 (N_14547,N_8890,N_8192);
nand U14548 (N_14548,N_6502,N_11244);
or U14549 (N_14549,N_8719,N_10553);
nand U14550 (N_14550,N_11857,N_6893);
nand U14551 (N_14551,N_10633,N_6176);
xnor U14552 (N_14552,N_11076,N_7227);
nor U14553 (N_14553,N_9639,N_8546);
xnor U14554 (N_14554,N_10094,N_6673);
nand U14555 (N_14555,N_7138,N_10587);
nand U14556 (N_14556,N_10508,N_7004);
xor U14557 (N_14557,N_8840,N_7413);
or U14558 (N_14558,N_8164,N_9870);
and U14559 (N_14559,N_6626,N_6093);
and U14560 (N_14560,N_7590,N_8325);
xor U14561 (N_14561,N_8986,N_10335);
or U14562 (N_14562,N_7363,N_7766);
nand U14563 (N_14563,N_11675,N_10549);
nand U14564 (N_14564,N_9989,N_9485);
and U14565 (N_14565,N_7641,N_9505);
nand U14566 (N_14566,N_7753,N_6154);
nand U14567 (N_14567,N_11626,N_11448);
nor U14568 (N_14568,N_10005,N_11862);
and U14569 (N_14569,N_8407,N_9289);
and U14570 (N_14570,N_7155,N_8706);
nand U14571 (N_14571,N_6436,N_11122);
or U14572 (N_14572,N_6080,N_11853);
or U14573 (N_14573,N_11034,N_10032);
and U14574 (N_14574,N_10826,N_11284);
or U14575 (N_14575,N_11040,N_10193);
and U14576 (N_14576,N_8092,N_8078);
and U14577 (N_14577,N_8874,N_10960);
nand U14578 (N_14578,N_7024,N_6615);
xor U14579 (N_14579,N_7510,N_7727);
nand U14580 (N_14580,N_7078,N_7579);
and U14581 (N_14581,N_8736,N_11224);
nand U14582 (N_14582,N_7687,N_11934);
xor U14583 (N_14583,N_8028,N_9501);
nand U14584 (N_14584,N_6301,N_11061);
or U14585 (N_14585,N_7448,N_9402);
nand U14586 (N_14586,N_6012,N_7780);
nand U14587 (N_14587,N_11727,N_9086);
nand U14588 (N_14588,N_6943,N_7414);
nor U14589 (N_14589,N_9545,N_7550);
and U14590 (N_14590,N_9111,N_11022);
nand U14591 (N_14591,N_7197,N_6174);
or U14592 (N_14592,N_11273,N_11451);
or U14593 (N_14593,N_11253,N_8456);
and U14594 (N_14594,N_10444,N_8828);
nor U14595 (N_14595,N_9366,N_10631);
nor U14596 (N_14596,N_11548,N_11948);
nand U14597 (N_14597,N_11246,N_8579);
or U14598 (N_14598,N_9566,N_8620);
and U14599 (N_14599,N_6383,N_6608);
nor U14600 (N_14600,N_7381,N_6762);
nor U14601 (N_14601,N_9247,N_6970);
or U14602 (N_14602,N_11137,N_7300);
nor U14603 (N_14603,N_6660,N_9898);
or U14604 (N_14604,N_9033,N_9719);
xnor U14605 (N_14605,N_8299,N_6720);
nor U14606 (N_14606,N_6069,N_11129);
xnor U14607 (N_14607,N_10221,N_8439);
or U14608 (N_14608,N_10863,N_10426);
xor U14609 (N_14609,N_11117,N_11392);
xnor U14610 (N_14610,N_10501,N_7498);
and U14611 (N_14611,N_9834,N_10431);
or U14612 (N_14612,N_9877,N_9323);
or U14613 (N_14613,N_11578,N_7907);
nand U14614 (N_14614,N_6164,N_11560);
xnor U14615 (N_14615,N_9009,N_11376);
nor U14616 (N_14616,N_11271,N_7568);
and U14617 (N_14617,N_8540,N_11480);
or U14618 (N_14618,N_9391,N_6428);
nor U14619 (N_14619,N_9330,N_9429);
nand U14620 (N_14620,N_11071,N_7918);
nor U14621 (N_14621,N_10695,N_10827);
xor U14622 (N_14622,N_9056,N_10250);
or U14623 (N_14623,N_7910,N_9573);
and U14624 (N_14624,N_8060,N_6643);
and U14625 (N_14625,N_6463,N_7250);
nand U14626 (N_14626,N_7426,N_9816);
or U14627 (N_14627,N_7157,N_11641);
nand U14628 (N_14628,N_7033,N_10612);
nand U14629 (N_14629,N_6692,N_8279);
nor U14630 (N_14630,N_8529,N_7152);
xor U14631 (N_14631,N_10671,N_7182);
and U14632 (N_14632,N_6095,N_8787);
and U14633 (N_14633,N_8516,N_11492);
nand U14634 (N_14634,N_7945,N_11788);
and U14635 (N_14635,N_10334,N_9050);
or U14636 (N_14636,N_9449,N_7055);
and U14637 (N_14637,N_7304,N_7229);
nand U14638 (N_14638,N_11764,N_8358);
or U14639 (N_14639,N_6930,N_11391);
or U14640 (N_14640,N_7551,N_9253);
xnor U14641 (N_14641,N_7816,N_9596);
nor U14642 (N_14642,N_6731,N_11759);
nand U14643 (N_14643,N_9701,N_8364);
or U14644 (N_14644,N_6742,N_9343);
nor U14645 (N_14645,N_9428,N_10683);
xor U14646 (N_14646,N_6602,N_11522);
xnor U14647 (N_14647,N_9066,N_6081);
nor U14648 (N_14648,N_10849,N_10255);
xor U14649 (N_14649,N_11332,N_6550);
or U14650 (N_14650,N_7123,N_9136);
xnor U14651 (N_14651,N_10943,N_6306);
xnor U14652 (N_14652,N_6064,N_6563);
or U14653 (N_14653,N_8377,N_10890);
and U14654 (N_14654,N_10033,N_8094);
or U14655 (N_14655,N_6260,N_9024);
nand U14656 (N_14656,N_6757,N_7220);
or U14657 (N_14657,N_11781,N_11855);
nand U14658 (N_14658,N_7512,N_7056);
and U14659 (N_14659,N_7147,N_7292);
nand U14660 (N_14660,N_11938,N_9413);
and U14661 (N_14661,N_10886,N_10415);
and U14662 (N_14662,N_11532,N_6613);
nor U14663 (N_14663,N_8867,N_10084);
nand U14664 (N_14664,N_10569,N_6948);
nor U14665 (N_14665,N_10364,N_10212);
nor U14666 (N_14666,N_9517,N_9742);
or U14667 (N_14667,N_11643,N_9551);
or U14668 (N_14668,N_8035,N_9818);
or U14669 (N_14669,N_7073,N_8034);
and U14670 (N_14670,N_11574,N_11595);
xor U14671 (N_14671,N_8405,N_8380);
and U14672 (N_14672,N_6338,N_6771);
xnor U14673 (N_14673,N_10482,N_6867);
nor U14674 (N_14674,N_8110,N_10300);
xnor U14675 (N_14675,N_7312,N_9114);
or U14676 (N_14676,N_10879,N_11571);
or U14677 (N_14677,N_11235,N_6382);
nand U14678 (N_14678,N_8756,N_8723);
xor U14679 (N_14679,N_7452,N_6553);
and U14680 (N_14680,N_8057,N_9913);
xnor U14681 (N_14681,N_7005,N_6714);
or U14682 (N_14682,N_9813,N_6909);
nand U14683 (N_14683,N_8742,N_8901);
nor U14684 (N_14684,N_11895,N_8881);
and U14685 (N_14685,N_10350,N_11312);
nor U14686 (N_14686,N_6940,N_11090);
nand U14687 (N_14687,N_8085,N_8583);
nor U14688 (N_14688,N_11955,N_11555);
or U14689 (N_14689,N_11604,N_6873);
or U14690 (N_14690,N_11079,N_6423);
nor U14691 (N_14691,N_11622,N_8965);
nand U14692 (N_14692,N_7891,N_8958);
nand U14693 (N_14693,N_11802,N_6968);
nor U14694 (N_14694,N_8240,N_11466);
nor U14695 (N_14695,N_9774,N_9796);
or U14696 (N_14696,N_11236,N_11881);
and U14697 (N_14697,N_7545,N_10368);
nor U14698 (N_14698,N_7788,N_7747);
nand U14699 (N_14699,N_9759,N_6265);
nor U14700 (N_14700,N_8566,N_10959);
and U14701 (N_14701,N_10998,N_9314);
xor U14702 (N_14702,N_8141,N_10145);
nor U14703 (N_14703,N_9140,N_10270);
nand U14704 (N_14704,N_11897,N_8852);
and U14705 (N_14705,N_6025,N_8857);
or U14706 (N_14706,N_11827,N_7289);
nand U14707 (N_14707,N_11733,N_9930);
and U14708 (N_14708,N_8985,N_10925);
or U14709 (N_14709,N_8825,N_10580);
nand U14710 (N_14710,N_7670,N_6324);
or U14711 (N_14711,N_10702,N_9711);
or U14712 (N_14712,N_8599,N_11593);
xor U14713 (N_14713,N_7895,N_8498);
nand U14714 (N_14714,N_8482,N_9805);
nand U14715 (N_14715,N_9293,N_6291);
nand U14716 (N_14716,N_9683,N_11822);
nor U14717 (N_14717,N_7239,N_9738);
and U14718 (N_14718,N_10321,N_11742);
and U14719 (N_14719,N_9610,N_9160);
xnor U14720 (N_14720,N_10992,N_9166);
nor U14721 (N_14721,N_10792,N_6457);
and U14722 (N_14722,N_10089,N_9605);
or U14723 (N_14723,N_10749,N_6481);
nand U14724 (N_14724,N_8898,N_7595);
nand U14725 (N_14725,N_8160,N_11267);
and U14726 (N_14726,N_9953,N_8937);
nor U14727 (N_14727,N_6319,N_8894);
nor U14728 (N_14728,N_7537,N_10196);
nor U14729 (N_14729,N_7617,N_6289);
nor U14730 (N_14730,N_11303,N_6795);
and U14731 (N_14731,N_11005,N_8031);
xnor U14732 (N_14732,N_9483,N_10469);
xnor U14733 (N_14733,N_9052,N_7211);
nand U14734 (N_14734,N_7629,N_10072);
nor U14735 (N_14735,N_8663,N_6335);
and U14736 (N_14736,N_9946,N_6002);
or U14737 (N_14737,N_8559,N_10613);
nand U14738 (N_14738,N_11513,N_11994);
xnor U14739 (N_14739,N_6305,N_8704);
xnor U14740 (N_14740,N_11717,N_11068);
xnor U14741 (N_14741,N_7778,N_8592);
nand U14742 (N_14742,N_8665,N_11019);
xor U14743 (N_14743,N_11352,N_9914);
nor U14744 (N_14744,N_7927,N_10940);
and U14745 (N_14745,N_7815,N_10272);
nor U14746 (N_14746,N_6193,N_6033);
or U14747 (N_14747,N_9769,N_10534);
xor U14748 (N_14748,N_8200,N_8917);
xnor U14749 (N_14749,N_10789,N_11232);
nand U14750 (N_14750,N_6664,N_11159);
and U14751 (N_14751,N_10836,N_10225);
nand U14752 (N_14752,N_11083,N_8582);
and U14753 (N_14753,N_9158,N_7785);
and U14754 (N_14754,N_9655,N_9023);
nor U14755 (N_14755,N_10648,N_7611);
nor U14756 (N_14756,N_9663,N_10678);
nand U14757 (N_14757,N_10022,N_8732);
or U14758 (N_14758,N_9574,N_9678);
and U14759 (N_14759,N_9916,N_6378);
xor U14760 (N_14760,N_6303,N_9915);
nor U14761 (N_14761,N_8919,N_10990);
nand U14762 (N_14762,N_9671,N_9745);
xnor U14763 (N_14763,N_11152,N_10870);
xor U14764 (N_14764,N_6695,N_7760);
nor U14765 (N_14765,N_7032,N_10282);
and U14766 (N_14766,N_11362,N_7429);
or U14767 (N_14767,N_9880,N_10866);
and U14768 (N_14768,N_6058,N_9080);
or U14769 (N_14769,N_10935,N_9302);
nor U14770 (N_14770,N_9899,N_11518);
nand U14771 (N_14771,N_7343,N_8076);
or U14772 (N_14772,N_9040,N_9925);
nand U14773 (N_14773,N_9651,N_10086);
xnor U14774 (N_14774,N_6198,N_7058);
nor U14775 (N_14775,N_7556,N_8100);
nor U14776 (N_14776,N_9848,N_10560);
nor U14777 (N_14777,N_6147,N_8891);
or U14778 (N_14778,N_9225,N_7865);
and U14779 (N_14779,N_6425,N_9536);
nor U14780 (N_14780,N_9425,N_8522);
or U14781 (N_14781,N_9828,N_7506);
or U14782 (N_14782,N_11506,N_9855);
or U14783 (N_14783,N_10540,N_6881);
or U14784 (N_14784,N_11596,N_6957);
xnor U14785 (N_14785,N_10243,N_7871);
and U14786 (N_14786,N_7995,N_8153);
or U14787 (N_14787,N_6340,N_7704);
nand U14788 (N_14788,N_8554,N_8697);
xor U14789 (N_14789,N_10906,N_11885);
nand U14790 (N_14790,N_7731,N_11609);
nor U14791 (N_14791,N_10918,N_9665);
and U14792 (N_14792,N_9728,N_7863);
and U14793 (N_14793,N_10158,N_11116);
and U14794 (N_14794,N_11977,N_9143);
nand U14795 (N_14795,N_10744,N_11043);
and U14796 (N_14796,N_7020,N_7943);
nor U14797 (N_14797,N_11097,N_10055);
xnor U14798 (N_14798,N_10956,N_11042);
nor U14799 (N_14799,N_6754,N_7613);
nand U14800 (N_14800,N_11234,N_8955);
and U14801 (N_14801,N_7956,N_9646);
xor U14802 (N_14802,N_7844,N_6825);
nor U14803 (N_14803,N_6498,N_8781);
or U14804 (N_14804,N_10764,N_6098);
nand U14805 (N_14805,N_7906,N_8932);
xor U14806 (N_14806,N_8423,N_6263);
xor U14807 (N_14807,N_8151,N_7146);
nor U14808 (N_14808,N_7830,N_10275);
xor U14809 (N_14809,N_10016,N_10099);
or U14810 (N_14810,N_8873,N_11297);
and U14811 (N_14811,N_7082,N_11820);
xor U14812 (N_14812,N_8470,N_6662);
and U14813 (N_14813,N_11055,N_8371);
or U14814 (N_14814,N_9872,N_7477);
nor U14815 (N_14815,N_9013,N_10574);
and U14816 (N_14816,N_11240,N_11394);
or U14817 (N_14817,N_6981,N_10991);
and U14818 (N_14818,N_7497,N_7383);
nor U14819 (N_14819,N_8680,N_10997);
nor U14820 (N_14820,N_7261,N_10021);
nor U14821 (N_14821,N_6205,N_9444);
nor U14822 (N_14822,N_7007,N_8794);
or U14823 (N_14823,N_6083,N_10494);
or U14824 (N_14824,N_9644,N_7111);
or U14825 (N_14825,N_6400,N_8408);
or U14826 (N_14826,N_10437,N_6617);
nor U14827 (N_14827,N_7874,N_11298);
nand U14828 (N_14828,N_9612,N_11702);
nand U14829 (N_14829,N_8944,N_6783);
and U14830 (N_14830,N_11201,N_6775);
or U14831 (N_14831,N_6764,N_9907);
nor U14832 (N_14832,N_7719,N_9345);
and U14833 (N_14833,N_11516,N_11104);
and U14834 (N_14834,N_11412,N_9109);
or U14835 (N_14835,N_8616,N_11677);
or U14836 (N_14836,N_10786,N_9304);
xnor U14837 (N_14837,N_6633,N_9768);
nand U14838 (N_14838,N_10238,N_6539);
and U14839 (N_14839,N_6257,N_6497);
nand U14840 (N_14840,N_10900,N_6001);
or U14841 (N_14841,N_11132,N_8216);
or U14842 (N_14842,N_6226,N_6212);
and U14843 (N_14843,N_7298,N_11374);
and U14844 (N_14844,N_10556,N_11814);
and U14845 (N_14845,N_11685,N_8318);
nor U14846 (N_14846,N_7296,N_8581);
xnor U14847 (N_14847,N_11300,N_11592);
nand U14848 (N_14848,N_11550,N_8426);
nor U14849 (N_14849,N_8084,N_11793);
nor U14850 (N_14850,N_10045,N_10772);
or U14851 (N_14851,N_8106,N_7286);
and U14852 (N_14852,N_6066,N_11109);
nor U14853 (N_14853,N_7410,N_9947);
xor U14854 (N_14854,N_8330,N_6368);
and U14855 (N_14855,N_6181,N_8983);
xor U14856 (N_14856,N_8041,N_10927);
nand U14857 (N_14857,N_7490,N_11843);
xnor U14858 (N_14858,N_7850,N_6809);
nand U14859 (N_14859,N_8180,N_6015);
xor U14860 (N_14860,N_11573,N_7150);
and U14861 (N_14861,N_11873,N_10333);
xnor U14862 (N_14862,N_11852,N_10563);
nand U14863 (N_14863,N_7288,N_10416);
and U14864 (N_14864,N_8544,N_7368);
nor U14865 (N_14865,N_11785,N_10684);
xnor U14866 (N_14866,N_8403,N_10798);
and U14867 (N_14867,N_6173,N_10978);
or U14868 (N_14868,N_11386,N_10853);
nor U14869 (N_14869,N_10400,N_11498);
nand U14870 (N_14870,N_9043,N_11269);
nor U14871 (N_14871,N_6687,N_8185);
and U14872 (N_14872,N_9092,N_9403);
and U14873 (N_14873,N_6654,N_11767);
nand U14874 (N_14874,N_10937,N_9183);
nor U14875 (N_14875,N_10081,N_6853);
nor U14876 (N_14876,N_11128,N_11779);
or U14877 (N_14877,N_11258,N_6207);
xor U14878 (N_14878,N_7091,N_8017);
xnor U14879 (N_14879,N_9633,N_6533);
nor U14880 (N_14880,N_8548,N_10923);
nor U14881 (N_14881,N_9645,N_6713);
and U14882 (N_14882,N_9849,N_8226);
or U14883 (N_14883,N_11956,N_7511);
nand U14884 (N_14884,N_8093,N_6812);
nor U14885 (N_14885,N_10816,N_10673);
or U14886 (N_14886,N_8744,N_8294);
nor U14887 (N_14887,N_10118,N_7268);
and U14888 (N_14888,N_10456,N_9548);
xnor U14889 (N_14889,N_7539,N_8312);
nor U14890 (N_14890,N_9531,N_11486);
and U14891 (N_14891,N_10743,N_9373);
nand U14892 (N_14892,N_8246,N_8928);
and U14893 (N_14893,N_8202,N_7341);
nand U14894 (N_14894,N_9176,N_11828);
nor U14895 (N_14895,N_9535,N_10532);
or U14896 (N_14896,N_11634,N_10061);
and U14897 (N_14897,N_9875,N_10268);
nor U14898 (N_14898,N_9674,N_10037);
or U14899 (N_14899,N_10289,N_10159);
nand U14900 (N_14900,N_10205,N_9955);
and U14901 (N_14901,N_11278,N_9262);
nand U14902 (N_14902,N_11892,N_7947);
nor U14903 (N_14903,N_10536,N_10127);
nand U14904 (N_14904,N_10623,N_6414);
xor U14905 (N_14905,N_8095,N_6792);
nor U14906 (N_14906,N_11799,N_6911);
nor U14907 (N_14907,N_11211,N_10878);
and U14908 (N_14908,N_9306,N_9509);
nand U14909 (N_14909,N_11794,N_6307);
and U14910 (N_14910,N_7905,N_8926);
and U14911 (N_14911,N_7287,N_11613);
or U14912 (N_14912,N_11459,N_10490);
and U14913 (N_14913,N_6859,N_6086);
and U14914 (N_14914,N_9954,N_8066);
nor U14915 (N_14915,N_7638,N_10231);
nand U14916 (N_14916,N_8088,N_8860);
xnor U14917 (N_14917,N_6159,N_7902);
xnor U14918 (N_14918,N_10838,N_6997);
and U14919 (N_14919,N_10080,N_6035);
nand U14920 (N_14920,N_6743,N_8636);
xnor U14921 (N_14921,N_10405,N_11693);
and U14922 (N_14922,N_11556,N_9207);
and U14923 (N_14923,N_8767,N_7316);
or U14924 (N_14924,N_6462,N_7195);
nor U14925 (N_14925,N_7188,N_9901);
xnor U14926 (N_14926,N_8039,N_6262);
nor U14927 (N_14927,N_6890,N_10195);
or U14928 (N_14928,N_8959,N_7284);
nor U14929 (N_14929,N_8285,N_10015);
xnor U14930 (N_14930,N_6536,N_9780);
or U14931 (N_14931,N_9290,N_6054);
or U14932 (N_14932,N_11098,N_7167);
nor U14933 (N_14933,N_7883,N_11321);
or U14934 (N_14934,N_8555,N_9171);
xor U14935 (N_14935,N_11663,N_11141);
nand U14936 (N_14936,N_6356,N_6320);
xor U14937 (N_14937,N_10412,N_6727);
and U14938 (N_14938,N_10347,N_8741);
or U14939 (N_14939,N_11504,N_7206);
xnor U14940 (N_14940,N_11701,N_10850);
nor U14941 (N_14941,N_10078,N_10645);
or U14942 (N_14942,N_8692,N_9303);
nand U14943 (N_14943,N_11796,N_8319);
or U14944 (N_14944,N_6763,N_8502);
nor U14945 (N_14945,N_10939,N_7562);
or U14946 (N_14946,N_7934,N_8766);
nor U14947 (N_14947,N_8848,N_9062);
or U14948 (N_14948,N_8990,N_9301);
and U14949 (N_14949,N_9189,N_6913);
xnor U14950 (N_14950,N_10961,N_8841);
nand U14951 (N_14951,N_6611,N_9770);
or U14952 (N_14952,N_6312,N_9723);
or U14953 (N_14953,N_11164,N_10599);
or U14954 (N_14954,N_11000,N_6590);
and U14955 (N_14955,N_6937,N_6586);
xnor U14956 (N_14956,N_6078,N_7959);
xnor U14957 (N_14957,N_8727,N_7807);
and U14958 (N_14958,N_6166,N_10981);
nor U14959 (N_14959,N_10787,N_10643);
xnor U14960 (N_14960,N_8671,N_7824);
xnor U14961 (N_14961,N_10914,N_6707);
nand U14962 (N_14962,N_7192,N_6331);
xor U14963 (N_14963,N_9677,N_6666);
nand U14964 (N_14964,N_10317,N_6155);
or U14965 (N_14965,N_6092,N_10660);
nand U14966 (N_14966,N_7478,N_11583);
and U14967 (N_14967,N_10761,N_9239);
or U14968 (N_14968,N_7971,N_9075);
nand U14969 (N_14969,N_6137,N_7173);
and U14970 (N_14970,N_11903,N_11987);
nor U14971 (N_14971,N_9891,N_8464);
and U14972 (N_14972,N_11552,N_8210);
and U14973 (N_14973,N_6189,N_10262);
nor U14974 (N_14974,N_7858,N_11277);
xnor U14975 (N_14975,N_8242,N_10813);
nand U14976 (N_14976,N_8280,N_7988);
nor U14977 (N_14977,N_6344,N_10902);
or U14978 (N_14978,N_7571,N_9217);
nand U14979 (N_14979,N_9351,N_9820);
or U14980 (N_14980,N_7694,N_6020);
or U14981 (N_14981,N_10073,N_8170);
or U14982 (N_14982,N_10846,N_6084);
and U14983 (N_14983,N_7795,N_11427);
xor U14984 (N_14984,N_11425,N_7576);
and U14985 (N_14985,N_9956,N_11708);
nor U14986 (N_14986,N_9826,N_6703);
or U14987 (N_14987,N_10462,N_6236);
nand U14988 (N_14988,N_7306,N_10263);
nor U14989 (N_14989,N_11038,N_11633);
xnor U14990 (N_14990,N_8929,N_10035);
or U14991 (N_14991,N_7500,N_7915);
and U14992 (N_14992,N_9734,N_8895);
and U14993 (N_14993,N_9014,N_6059);
nand U14994 (N_14994,N_6581,N_9579);
or U14995 (N_14995,N_6620,N_6512);
nand U14996 (N_14996,N_10865,N_7764);
and U14997 (N_14997,N_8749,N_6932);
or U14998 (N_14998,N_9462,N_9555);
nand U14999 (N_14999,N_10615,N_7622);
nand U15000 (N_15000,N_11563,N_8307);
nand U15001 (N_15001,N_6125,N_11481);
or U15002 (N_15002,N_9261,N_10360);
nand U15003 (N_15003,N_10118,N_9894);
nand U15004 (N_15004,N_11299,N_9643);
or U15005 (N_15005,N_6791,N_9812);
xor U15006 (N_15006,N_10224,N_8952);
xor U15007 (N_15007,N_6189,N_10222);
and U15008 (N_15008,N_7777,N_8937);
nand U15009 (N_15009,N_6215,N_7650);
nand U15010 (N_15010,N_10524,N_6698);
or U15011 (N_15011,N_10304,N_7446);
nor U15012 (N_15012,N_8638,N_10771);
xnor U15013 (N_15013,N_9057,N_10679);
xnor U15014 (N_15014,N_7669,N_10121);
or U15015 (N_15015,N_7517,N_9529);
nor U15016 (N_15016,N_10932,N_6497);
nand U15017 (N_15017,N_6395,N_7060);
xnor U15018 (N_15018,N_8006,N_8571);
xor U15019 (N_15019,N_7699,N_7617);
nand U15020 (N_15020,N_7644,N_6420);
nand U15021 (N_15021,N_9017,N_11425);
xor U15022 (N_15022,N_7793,N_9721);
xnor U15023 (N_15023,N_10217,N_10653);
or U15024 (N_15024,N_8428,N_7744);
xnor U15025 (N_15025,N_11530,N_11809);
or U15026 (N_15026,N_9608,N_8015);
or U15027 (N_15027,N_9921,N_10004);
and U15028 (N_15028,N_7969,N_9218);
and U15029 (N_15029,N_10648,N_11439);
or U15030 (N_15030,N_11255,N_10528);
xor U15031 (N_15031,N_8233,N_9749);
nand U15032 (N_15032,N_10798,N_10448);
nand U15033 (N_15033,N_11660,N_8391);
or U15034 (N_15034,N_9273,N_6060);
nand U15035 (N_15035,N_7068,N_10750);
xor U15036 (N_15036,N_8038,N_10906);
nand U15037 (N_15037,N_9391,N_8258);
or U15038 (N_15038,N_7798,N_11704);
xor U15039 (N_15039,N_11589,N_11662);
xor U15040 (N_15040,N_7503,N_10069);
or U15041 (N_15041,N_11496,N_7653);
and U15042 (N_15042,N_11885,N_10556);
or U15043 (N_15043,N_10789,N_7885);
or U15044 (N_15044,N_8822,N_11608);
xnor U15045 (N_15045,N_7661,N_11028);
nand U15046 (N_15046,N_8631,N_6533);
nor U15047 (N_15047,N_9031,N_6520);
or U15048 (N_15048,N_7082,N_10048);
and U15049 (N_15049,N_11259,N_8592);
xnor U15050 (N_15050,N_11391,N_6233);
nand U15051 (N_15051,N_10920,N_7212);
and U15052 (N_15052,N_6568,N_11448);
and U15053 (N_15053,N_6809,N_11573);
xnor U15054 (N_15054,N_6449,N_11255);
nor U15055 (N_15055,N_7371,N_7513);
and U15056 (N_15056,N_11909,N_9812);
and U15057 (N_15057,N_6954,N_10096);
xor U15058 (N_15058,N_11280,N_10637);
or U15059 (N_15059,N_7055,N_6499);
or U15060 (N_15060,N_10022,N_8981);
and U15061 (N_15061,N_9832,N_10208);
nor U15062 (N_15062,N_9619,N_11620);
nor U15063 (N_15063,N_9753,N_7981);
and U15064 (N_15064,N_9657,N_11374);
nand U15065 (N_15065,N_9786,N_11431);
xnor U15066 (N_15066,N_7563,N_8415);
and U15067 (N_15067,N_8332,N_7837);
xnor U15068 (N_15068,N_6413,N_10985);
nor U15069 (N_15069,N_7053,N_6766);
nand U15070 (N_15070,N_6434,N_11718);
or U15071 (N_15071,N_9064,N_6551);
and U15072 (N_15072,N_6996,N_10743);
nand U15073 (N_15073,N_10648,N_6162);
or U15074 (N_15074,N_8955,N_8577);
or U15075 (N_15075,N_8597,N_6140);
nor U15076 (N_15076,N_10659,N_10697);
nor U15077 (N_15077,N_6429,N_8171);
xnor U15078 (N_15078,N_7157,N_6261);
and U15079 (N_15079,N_10856,N_6734);
nand U15080 (N_15080,N_10524,N_6749);
nand U15081 (N_15081,N_6912,N_11078);
nand U15082 (N_15082,N_6896,N_9662);
xor U15083 (N_15083,N_9986,N_11367);
or U15084 (N_15084,N_6991,N_9675);
and U15085 (N_15085,N_8938,N_10084);
nor U15086 (N_15086,N_8691,N_8122);
xor U15087 (N_15087,N_8359,N_10394);
xnor U15088 (N_15088,N_9046,N_11315);
xor U15089 (N_15089,N_6639,N_9545);
or U15090 (N_15090,N_7059,N_11676);
nand U15091 (N_15091,N_8022,N_10556);
nor U15092 (N_15092,N_9416,N_7587);
or U15093 (N_15093,N_11342,N_6355);
nand U15094 (N_15094,N_10629,N_7640);
or U15095 (N_15095,N_6945,N_6081);
nand U15096 (N_15096,N_11856,N_10850);
and U15097 (N_15097,N_6395,N_7325);
nand U15098 (N_15098,N_6448,N_8500);
and U15099 (N_15099,N_6475,N_11094);
or U15100 (N_15100,N_7010,N_10245);
nor U15101 (N_15101,N_9714,N_9168);
xor U15102 (N_15102,N_9414,N_8466);
and U15103 (N_15103,N_6662,N_9024);
or U15104 (N_15104,N_8910,N_10215);
xnor U15105 (N_15105,N_8349,N_8900);
or U15106 (N_15106,N_10550,N_11749);
or U15107 (N_15107,N_11178,N_7182);
nor U15108 (N_15108,N_10387,N_11462);
xnor U15109 (N_15109,N_10350,N_6525);
xnor U15110 (N_15110,N_8969,N_11308);
nor U15111 (N_15111,N_6527,N_6150);
nand U15112 (N_15112,N_11825,N_6090);
nor U15113 (N_15113,N_6107,N_10326);
xor U15114 (N_15114,N_7075,N_10940);
or U15115 (N_15115,N_10083,N_7029);
and U15116 (N_15116,N_8705,N_7294);
or U15117 (N_15117,N_8047,N_9943);
or U15118 (N_15118,N_9439,N_6455);
and U15119 (N_15119,N_6552,N_9409);
nor U15120 (N_15120,N_10901,N_11483);
nor U15121 (N_15121,N_11016,N_9439);
nand U15122 (N_15122,N_9254,N_8222);
xnor U15123 (N_15123,N_8661,N_8426);
nor U15124 (N_15124,N_9810,N_11683);
and U15125 (N_15125,N_6647,N_10461);
or U15126 (N_15126,N_8364,N_11692);
or U15127 (N_15127,N_6223,N_9954);
xnor U15128 (N_15128,N_6527,N_11612);
xor U15129 (N_15129,N_10309,N_10770);
nor U15130 (N_15130,N_9320,N_9149);
and U15131 (N_15131,N_11025,N_7764);
and U15132 (N_15132,N_10399,N_8184);
and U15133 (N_15133,N_8424,N_11496);
and U15134 (N_15134,N_11500,N_7103);
or U15135 (N_15135,N_7731,N_7983);
nor U15136 (N_15136,N_8686,N_8538);
nor U15137 (N_15137,N_11632,N_9611);
or U15138 (N_15138,N_6254,N_6061);
nor U15139 (N_15139,N_7389,N_6712);
and U15140 (N_15140,N_10574,N_9776);
and U15141 (N_15141,N_9558,N_11546);
nand U15142 (N_15142,N_10704,N_10269);
xor U15143 (N_15143,N_9696,N_8817);
and U15144 (N_15144,N_6063,N_11771);
or U15145 (N_15145,N_9084,N_9607);
nand U15146 (N_15146,N_10926,N_8749);
xor U15147 (N_15147,N_6798,N_6692);
and U15148 (N_15148,N_8027,N_7178);
nor U15149 (N_15149,N_8669,N_10358);
nand U15150 (N_15150,N_9516,N_11248);
nor U15151 (N_15151,N_9476,N_7104);
xor U15152 (N_15152,N_8373,N_7392);
nor U15153 (N_15153,N_10934,N_8770);
and U15154 (N_15154,N_11072,N_7942);
nand U15155 (N_15155,N_7610,N_11279);
and U15156 (N_15156,N_11083,N_9468);
or U15157 (N_15157,N_6574,N_10067);
or U15158 (N_15158,N_7307,N_6179);
xor U15159 (N_15159,N_7727,N_10618);
nand U15160 (N_15160,N_6258,N_9589);
or U15161 (N_15161,N_6348,N_7033);
nor U15162 (N_15162,N_6581,N_7390);
nand U15163 (N_15163,N_7899,N_10477);
xor U15164 (N_15164,N_6339,N_11710);
nor U15165 (N_15165,N_8658,N_8172);
and U15166 (N_15166,N_8962,N_7883);
nand U15167 (N_15167,N_9071,N_8167);
or U15168 (N_15168,N_8384,N_9060);
nor U15169 (N_15169,N_8453,N_6808);
xor U15170 (N_15170,N_9626,N_7192);
and U15171 (N_15171,N_9494,N_6503);
or U15172 (N_15172,N_7736,N_11295);
or U15173 (N_15173,N_8197,N_8299);
nor U15174 (N_15174,N_10261,N_6158);
or U15175 (N_15175,N_10808,N_6864);
and U15176 (N_15176,N_6074,N_9449);
nor U15177 (N_15177,N_9427,N_8876);
xnor U15178 (N_15178,N_7858,N_6876);
nand U15179 (N_15179,N_6664,N_9217);
xnor U15180 (N_15180,N_8395,N_10870);
xor U15181 (N_15181,N_7054,N_11822);
nand U15182 (N_15182,N_11788,N_10960);
xnor U15183 (N_15183,N_8264,N_10274);
nand U15184 (N_15184,N_7508,N_6913);
and U15185 (N_15185,N_8847,N_9344);
xor U15186 (N_15186,N_9759,N_11527);
xor U15187 (N_15187,N_7191,N_11738);
nand U15188 (N_15188,N_6192,N_7237);
or U15189 (N_15189,N_8562,N_7065);
nor U15190 (N_15190,N_11089,N_7939);
or U15191 (N_15191,N_7015,N_6722);
or U15192 (N_15192,N_7497,N_6875);
and U15193 (N_15193,N_8784,N_9887);
and U15194 (N_15194,N_8428,N_10983);
or U15195 (N_15195,N_7341,N_7641);
xor U15196 (N_15196,N_8566,N_11900);
xnor U15197 (N_15197,N_8733,N_9202);
or U15198 (N_15198,N_11025,N_11869);
and U15199 (N_15199,N_6868,N_9541);
and U15200 (N_15200,N_9188,N_6749);
or U15201 (N_15201,N_6464,N_7134);
or U15202 (N_15202,N_7772,N_9039);
or U15203 (N_15203,N_8517,N_7140);
xnor U15204 (N_15204,N_9434,N_7475);
nor U15205 (N_15205,N_9443,N_10035);
nor U15206 (N_15206,N_6011,N_10629);
and U15207 (N_15207,N_6325,N_6340);
and U15208 (N_15208,N_10987,N_11274);
nor U15209 (N_15209,N_11709,N_9612);
nor U15210 (N_15210,N_10795,N_7775);
xnor U15211 (N_15211,N_7922,N_9857);
nor U15212 (N_15212,N_6030,N_11729);
nor U15213 (N_15213,N_11866,N_7229);
xnor U15214 (N_15214,N_7556,N_8771);
and U15215 (N_15215,N_7092,N_10056);
xnor U15216 (N_15216,N_7339,N_7879);
or U15217 (N_15217,N_9620,N_7034);
or U15218 (N_15218,N_7946,N_8458);
or U15219 (N_15219,N_7440,N_9685);
xor U15220 (N_15220,N_11664,N_11400);
nor U15221 (N_15221,N_9575,N_11050);
and U15222 (N_15222,N_11738,N_10948);
or U15223 (N_15223,N_8916,N_10513);
xnor U15224 (N_15224,N_11523,N_8929);
and U15225 (N_15225,N_10161,N_6232);
and U15226 (N_15226,N_8654,N_10524);
nand U15227 (N_15227,N_8977,N_6704);
nand U15228 (N_15228,N_10729,N_11380);
nand U15229 (N_15229,N_6417,N_7099);
or U15230 (N_15230,N_8584,N_9061);
nand U15231 (N_15231,N_11095,N_8852);
nand U15232 (N_15232,N_11403,N_10280);
xnor U15233 (N_15233,N_6780,N_9423);
nor U15234 (N_15234,N_7038,N_6703);
nor U15235 (N_15235,N_11399,N_9391);
or U15236 (N_15236,N_6324,N_9190);
xor U15237 (N_15237,N_7478,N_6725);
xnor U15238 (N_15238,N_10599,N_11119);
xor U15239 (N_15239,N_6517,N_7808);
nand U15240 (N_15240,N_11061,N_7715);
and U15241 (N_15241,N_6861,N_9521);
xnor U15242 (N_15242,N_11669,N_7471);
nand U15243 (N_15243,N_7258,N_10022);
nor U15244 (N_15244,N_10464,N_8118);
or U15245 (N_15245,N_8392,N_7087);
xnor U15246 (N_15246,N_7229,N_6369);
and U15247 (N_15247,N_7718,N_7858);
and U15248 (N_15248,N_9496,N_6377);
xor U15249 (N_15249,N_8152,N_9498);
nor U15250 (N_15250,N_7737,N_8044);
and U15251 (N_15251,N_7382,N_9058);
or U15252 (N_15252,N_10824,N_8516);
or U15253 (N_15253,N_6494,N_7307);
nand U15254 (N_15254,N_7305,N_8792);
nand U15255 (N_15255,N_10093,N_8184);
nor U15256 (N_15256,N_6827,N_8588);
nor U15257 (N_15257,N_9180,N_11237);
nor U15258 (N_15258,N_9444,N_7774);
or U15259 (N_15259,N_10872,N_9740);
and U15260 (N_15260,N_10207,N_6092);
nor U15261 (N_15261,N_11811,N_11283);
and U15262 (N_15262,N_10688,N_7750);
or U15263 (N_15263,N_7331,N_10879);
xor U15264 (N_15264,N_10892,N_11368);
or U15265 (N_15265,N_10295,N_11412);
or U15266 (N_15266,N_10165,N_11557);
and U15267 (N_15267,N_10462,N_8115);
xor U15268 (N_15268,N_10102,N_10802);
or U15269 (N_15269,N_8627,N_7096);
nor U15270 (N_15270,N_7051,N_7764);
nand U15271 (N_15271,N_11227,N_10311);
nand U15272 (N_15272,N_8566,N_7182);
nand U15273 (N_15273,N_9265,N_7513);
or U15274 (N_15274,N_6967,N_6148);
or U15275 (N_15275,N_10956,N_9444);
nor U15276 (N_15276,N_10624,N_8231);
or U15277 (N_15277,N_7636,N_8535);
nand U15278 (N_15278,N_6978,N_8905);
and U15279 (N_15279,N_9569,N_11661);
and U15280 (N_15280,N_11116,N_9482);
xnor U15281 (N_15281,N_7838,N_6866);
or U15282 (N_15282,N_11238,N_9498);
or U15283 (N_15283,N_6284,N_8299);
nor U15284 (N_15284,N_9213,N_8846);
and U15285 (N_15285,N_11037,N_7164);
nand U15286 (N_15286,N_11153,N_11797);
xnor U15287 (N_15287,N_10360,N_11442);
or U15288 (N_15288,N_8630,N_9551);
or U15289 (N_15289,N_9748,N_6181);
or U15290 (N_15290,N_6294,N_7175);
nand U15291 (N_15291,N_10413,N_6319);
nor U15292 (N_15292,N_8286,N_8058);
xnor U15293 (N_15293,N_7618,N_9870);
nor U15294 (N_15294,N_9097,N_8382);
and U15295 (N_15295,N_11386,N_7909);
or U15296 (N_15296,N_6127,N_11178);
nor U15297 (N_15297,N_8736,N_10370);
or U15298 (N_15298,N_11789,N_8296);
xor U15299 (N_15299,N_9044,N_8610);
nor U15300 (N_15300,N_10042,N_9080);
and U15301 (N_15301,N_7194,N_7465);
nor U15302 (N_15302,N_8360,N_9707);
nand U15303 (N_15303,N_11030,N_6763);
nor U15304 (N_15304,N_11796,N_9348);
nand U15305 (N_15305,N_9020,N_9799);
nor U15306 (N_15306,N_11461,N_9731);
xnor U15307 (N_15307,N_9011,N_11777);
xnor U15308 (N_15308,N_10542,N_10807);
nor U15309 (N_15309,N_11140,N_7676);
or U15310 (N_15310,N_6472,N_10971);
nor U15311 (N_15311,N_9022,N_8086);
or U15312 (N_15312,N_10071,N_10790);
and U15313 (N_15313,N_8651,N_7813);
and U15314 (N_15314,N_10173,N_6333);
xnor U15315 (N_15315,N_6854,N_9759);
or U15316 (N_15316,N_10131,N_9130);
nor U15317 (N_15317,N_11824,N_8900);
or U15318 (N_15318,N_7711,N_6332);
and U15319 (N_15319,N_9792,N_6368);
or U15320 (N_15320,N_11550,N_10078);
nand U15321 (N_15321,N_7386,N_7435);
or U15322 (N_15322,N_11493,N_8085);
and U15323 (N_15323,N_11098,N_11739);
and U15324 (N_15324,N_9326,N_7107);
or U15325 (N_15325,N_7639,N_9693);
or U15326 (N_15326,N_9401,N_6316);
nand U15327 (N_15327,N_7894,N_11768);
nand U15328 (N_15328,N_6235,N_8208);
or U15329 (N_15329,N_9766,N_8469);
nor U15330 (N_15330,N_7815,N_10137);
and U15331 (N_15331,N_11307,N_7959);
nand U15332 (N_15332,N_11380,N_9041);
xnor U15333 (N_15333,N_6658,N_11740);
nand U15334 (N_15334,N_8606,N_11818);
or U15335 (N_15335,N_8331,N_9236);
nand U15336 (N_15336,N_7271,N_9311);
or U15337 (N_15337,N_10387,N_7274);
or U15338 (N_15338,N_9763,N_10504);
nor U15339 (N_15339,N_8432,N_10821);
nand U15340 (N_15340,N_10326,N_8006);
xor U15341 (N_15341,N_9654,N_10623);
nor U15342 (N_15342,N_8014,N_10317);
or U15343 (N_15343,N_8055,N_7534);
and U15344 (N_15344,N_11782,N_8102);
nand U15345 (N_15345,N_10276,N_10169);
or U15346 (N_15346,N_9256,N_6135);
nand U15347 (N_15347,N_11860,N_9424);
xnor U15348 (N_15348,N_11538,N_8981);
and U15349 (N_15349,N_10375,N_8382);
or U15350 (N_15350,N_10033,N_10462);
nor U15351 (N_15351,N_11514,N_11851);
nor U15352 (N_15352,N_8256,N_6381);
and U15353 (N_15353,N_9990,N_9762);
nor U15354 (N_15354,N_11327,N_9460);
nand U15355 (N_15355,N_6931,N_11416);
or U15356 (N_15356,N_9236,N_9606);
nand U15357 (N_15357,N_8534,N_7055);
or U15358 (N_15358,N_9831,N_6735);
and U15359 (N_15359,N_6666,N_8355);
nand U15360 (N_15360,N_9185,N_11023);
nand U15361 (N_15361,N_11373,N_7819);
nand U15362 (N_15362,N_8396,N_11973);
nand U15363 (N_15363,N_6329,N_6810);
and U15364 (N_15364,N_9390,N_10983);
and U15365 (N_15365,N_7837,N_6537);
or U15366 (N_15366,N_6689,N_6332);
or U15367 (N_15367,N_9102,N_9311);
nor U15368 (N_15368,N_8125,N_9372);
nor U15369 (N_15369,N_8576,N_11699);
nor U15370 (N_15370,N_11142,N_9986);
nor U15371 (N_15371,N_10181,N_8205);
or U15372 (N_15372,N_6250,N_11976);
and U15373 (N_15373,N_10104,N_11924);
or U15374 (N_15374,N_11443,N_11297);
and U15375 (N_15375,N_11922,N_11956);
or U15376 (N_15376,N_8908,N_7119);
or U15377 (N_15377,N_8977,N_7365);
nand U15378 (N_15378,N_6271,N_7720);
nand U15379 (N_15379,N_8074,N_6698);
nand U15380 (N_15380,N_10092,N_8565);
or U15381 (N_15381,N_11737,N_7232);
or U15382 (N_15382,N_8554,N_8095);
nor U15383 (N_15383,N_11883,N_8730);
and U15384 (N_15384,N_11585,N_7912);
xnor U15385 (N_15385,N_9754,N_6697);
nor U15386 (N_15386,N_10490,N_8974);
xnor U15387 (N_15387,N_6383,N_7253);
xnor U15388 (N_15388,N_6861,N_8005);
and U15389 (N_15389,N_6453,N_10332);
nand U15390 (N_15390,N_11917,N_6027);
and U15391 (N_15391,N_9476,N_11480);
xnor U15392 (N_15392,N_9402,N_10679);
xor U15393 (N_15393,N_10972,N_6079);
or U15394 (N_15394,N_7571,N_6569);
or U15395 (N_15395,N_8067,N_9015);
xnor U15396 (N_15396,N_9207,N_10842);
or U15397 (N_15397,N_6571,N_10019);
and U15398 (N_15398,N_11771,N_11823);
nand U15399 (N_15399,N_9543,N_11647);
nor U15400 (N_15400,N_7355,N_10884);
and U15401 (N_15401,N_11981,N_8849);
nor U15402 (N_15402,N_6008,N_9588);
and U15403 (N_15403,N_8122,N_10649);
xor U15404 (N_15404,N_10296,N_9936);
nand U15405 (N_15405,N_11488,N_10444);
nand U15406 (N_15406,N_10061,N_10831);
and U15407 (N_15407,N_7213,N_7256);
or U15408 (N_15408,N_7223,N_11629);
xor U15409 (N_15409,N_11305,N_8850);
nand U15410 (N_15410,N_8560,N_10912);
nand U15411 (N_15411,N_10056,N_11569);
and U15412 (N_15412,N_7509,N_7050);
nor U15413 (N_15413,N_11333,N_6794);
xnor U15414 (N_15414,N_7520,N_11024);
nand U15415 (N_15415,N_8132,N_7429);
xor U15416 (N_15416,N_10200,N_8970);
or U15417 (N_15417,N_9079,N_8410);
xnor U15418 (N_15418,N_9051,N_10318);
or U15419 (N_15419,N_10568,N_11355);
xnor U15420 (N_15420,N_8667,N_11820);
nand U15421 (N_15421,N_9514,N_6684);
nor U15422 (N_15422,N_9868,N_10400);
nand U15423 (N_15423,N_7423,N_8392);
nand U15424 (N_15424,N_6830,N_9447);
and U15425 (N_15425,N_8820,N_10017);
or U15426 (N_15426,N_8991,N_10586);
or U15427 (N_15427,N_11919,N_9018);
nor U15428 (N_15428,N_6657,N_8084);
and U15429 (N_15429,N_8395,N_9678);
or U15430 (N_15430,N_7463,N_8209);
xor U15431 (N_15431,N_6689,N_9051);
and U15432 (N_15432,N_8520,N_9725);
xnor U15433 (N_15433,N_11356,N_10675);
nor U15434 (N_15434,N_9621,N_11096);
xnor U15435 (N_15435,N_10688,N_7898);
nor U15436 (N_15436,N_8041,N_10333);
or U15437 (N_15437,N_9129,N_9726);
or U15438 (N_15438,N_9575,N_8422);
nor U15439 (N_15439,N_11469,N_8306);
xnor U15440 (N_15440,N_10895,N_9242);
nor U15441 (N_15441,N_8615,N_8662);
xor U15442 (N_15442,N_7369,N_8546);
or U15443 (N_15443,N_8160,N_9819);
nand U15444 (N_15444,N_8640,N_11475);
nand U15445 (N_15445,N_7402,N_8179);
and U15446 (N_15446,N_7665,N_10765);
and U15447 (N_15447,N_9254,N_9040);
and U15448 (N_15448,N_7138,N_11916);
or U15449 (N_15449,N_11105,N_11944);
nor U15450 (N_15450,N_7795,N_6051);
nor U15451 (N_15451,N_6157,N_9772);
and U15452 (N_15452,N_10117,N_9771);
nand U15453 (N_15453,N_7144,N_8067);
or U15454 (N_15454,N_10370,N_11767);
nand U15455 (N_15455,N_8351,N_7262);
nand U15456 (N_15456,N_11584,N_7510);
or U15457 (N_15457,N_11650,N_11100);
or U15458 (N_15458,N_7492,N_11938);
and U15459 (N_15459,N_9768,N_9531);
nor U15460 (N_15460,N_11354,N_10196);
nor U15461 (N_15461,N_7621,N_11334);
nor U15462 (N_15462,N_7121,N_6602);
or U15463 (N_15463,N_10133,N_8531);
or U15464 (N_15464,N_8910,N_6837);
or U15465 (N_15465,N_9673,N_9830);
or U15466 (N_15466,N_7980,N_10457);
and U15467 (N_15467,N_11874,N_11610);
nand U15468 (N_15468,N_11716,N_9932);
and U15469 (N_15469,N_10709,N_9761);
nand U15470 (N_15470,N_10523,N_8095);
xor U15471 (N_15471,N_6421,N_11741);
or U15472 (N_15472,N_8847,N_6402);
xor U15473 (N_15473,N_10501,N_9056);
nand U15474 (N_15474,N_10872,N_9995);
or U15475 (N_15475,N_6591,N_10119);
nor U15476 (N_15476,N_6379,N_6045);
xnor U15477 (N_15477,N_7164,N_10838);
xor U15478 (N_15478,N_6877,N_11366);
nand U15479 (N_15479,N_10088,N_7530);
and U15480 (N_15480,N_9318,N_7557);
xor U15481 (N_15481,N_7864,N_9883);
xor U15482 (N_15482,N_7831,N_6587);
xor U15483 (N_15483,N_9865,N_11009);
and U15484 (N_15484,N_6880,N_11607);
nor U15485 (N_15485,N_8773,N_10085);
nor U15486 (N_15486,N_7550,N_8697);
nand U15487 (N_15487,N_11315,N_8913);
xnor U15488 (N_15488,N_7422,N_10012);
xnor U15489 (N_15489,N_6594,N_10845);
xor U15490 (N_15490,N_10346,N_8227);
or U15491 (N_15491,N_7133,N_6556);
and U15492 (N_15492,N_9677,N_11478);
xnor U15493 (N_15493,N_6023,N_6828);
nand U15494 (N_15494,N_11067,N_11418);
nor U15495 (N_15495,N_7426,N_8858);
nor U15496 (N_15496,N_7736,N_10117);
xor U15497 (N_15497,N_11154,N_8181);
nand U15498 (N_15498,N_11379,N_7283);
and U15499 (N_15499,N_6112,N_11859);
or U15500 (N_15500,N_9184,N_7763);
xor U15501 (N_15501,N_7859,N_7519);
nand U15502 (N_15502,N_7713,N_11559);
xor U15503 (N_15503,N_6611,N_10849);
nand U15504 (N_15504,N_7065,N_11053);
nand U15505 (N_15505,N_10152,N_7849);
and U15506 (N_15506,N_8335,N_11461);
and U15507 (N_15507,N_8004,N_7479);
nand U15508 (N_15508,N_8332,N_10816);
xnor U15509 (N_15509,N_10315,N_11850);
nand U15510 (N_15510,N_6936,N_6462);
or U15511 (N_15511,N_11043,N_8417);
and U15512 (N_15512,N_8027,N_7936);
or U15513 (N_15513,N_9392,N_10532);
or U15514 (N_15514,N_8297,N_11653);
nand U15515 (N_15515,N_9491,N_10363);
nor U15516 (N_15516,N_7846,N_8724);
or U15517 (N_15517,N_8540,N_7763);
xor U15518 (N_15518,N_9223,N_11611);
nand U15519 (N_15519,N_7027,N_9486);
and U15520 (N_15520,N_9274,N_6131);
and U15521 (N_15521,N_9928,N_6740);
nor U15522 (N_15522,N_11247,N_7214);
nor U15523 (N_15523,N_10054,N_9412);
or U15524 (N_15524,N_6918,N_9683);
nand U15525 (N_15525,N_7684,N_6339);
or U15526 (N_15526,N_9340,N_6677);
nand U15527 (N_15527,N_11596,N_8751);
nand U15528 (N_15528,N_11588,N_11467);
nand U15529 (N_15529,N_10715,N_7628);
xnor U15530 (N_15530,N_6892,N_8759);
nor U15531 (N_15531,N_7291,N_10584);
nor U15532 (N_15532,N_6369,N_9126);
xnor U15533 (N_15533,N_10446,N_11075);
and U15534 (N_15534,N_11388,N_11579);
or U15535 (N_15535,N_6457,N_8135);
or U15536 (N_15536,N_9521,N_8831);
nor U15537 (N_15537,N_6331,N_6746);
or U15538 (N_15538,N_7849,N_10141);
xor U15539 (N_15539,N_10264,N_9569);
and U15540 (N_15540,N_10092,N_6492);
xor U15541 (N_15541,N_8137,N_7667);
nor U15542 (N_15542,N_8894,N_6665);
or U15543 (N_15543,N_8776,N_6678);
or U15544 (N_15544,N_8603,N_8509);
or U15545 (N_15545,N_10212,N_6643);
nor U15546 (N_15546,N_6467,N_6875);
nor U15547 (N_15547,N_6550,N_8437);
xor U15548 (N_15548,N_10137,N_6176);
xnor U15549 (N_15549,N_7656,N_9361);
and U15550 (N_15550,N_9721,N_6067);
nand U15551 (N_15551,N_8589,N_7680);
or U15552 (N_15552,N_10505,N_7876);
xor U15553 (N_15553,N_7996,N_7825);
or U15554 (N_15554,N_7686,N_9249);
xnor U15555 (N_15555,N_6322,N_9090);
and U15556 (N_15556,N_8780,N_7859);
xnor U15557 (N_15557,N_7745,N_10726);
or U15558 (N_15558,N_7647,N_10318);
nor U15559 (N_15559,N_10700,N_6178);
and U15560 (N_15560,N_6759,N_7638);
nor U15561 (N_15561,N_9588,N_10574);
or U15562 (N_15562,N_7926,N_9931);
nor U15563 (N_15563,N_8603,N_11101);
and U15564 (N_15564,N_7426,N_10081);
nand U15565 (N_15565,N_8598,N_8463);
nor U15566 (N_15566,N_8862,N_8542);
and U15567 (N_15567,N_9682,N_6019);
or U15568 (N_15568,N_11276,N_6174);
xor U15569 (N_15569,N_11627,N_10433);
xor U15570 (N_15570,N_8782,N_9034);
nor U15571 (N_15571,N_9523,N_9020);
or U15572 (N_15572,N_7600,N_6354);
nor U15573 (N_15573,N_8047,N_6840);
and U15574 (N_15574,N_11615,N_7076);
nand U15575 (N_15575,N_6845,N_7957);
and U15576 (N_15576,N_11529,N_6448);
nand U15577 (N_15577,N_8562,N_7339);
or U15578 (N_15578,N_9292,N_8505);
or U15579 (N_15579,N_6599,N_11549);
nand U15580 (N_15580,N_9105,N_10320);
nor U15581 (N_15581,N_10672,N_6725);
xnor U15582 (N_15582,N_8123,N_9843);
or U15583 (N_15583,N_9789,N_11462);
nor U15584 (N_15584,N_9789,N_6334);
nand U15585 (N_15585,N_11290,N_8031);
nor U15586 (N_15586,N_8868,N_6944);
or U15587 (N_15587,N_8165,N_10431);
and U15588 (N_15588,N_7007,N_7931);
nor U15589 (N_15589,N_10266,N_8306);
nor U15590 (N_15590,N_7261,N_9072);
nand U15591 (N_15591,N_10847,N_7143);
xor U15592 (N_15592,N_11038,N_10050);
nand U15593 (N_15593,N_11419,N_11338);
xor U15594 (N_15594,N_8830,N_8309);
nor U15595 (N_15595,N_8554,N_7162);
xor U15596 (N_15596,N_8611,N_10063);
xnor U15597 (N_15597,N_7212,N_10498);
and U15598 (N_15598,N_6408,N_7715);
and U15599 (N_15599,N_8307,N_6087);
nor U15600 (N_15600,N_7270,N_7981);
and U15601 (N_15601,N_8798,N_11226);
or U15602 (N_15602,N_11252,N_6744);
nor U15603 (N_15603,N_8190,N_8897);
nand U15604 (N_15604,N_10359,N_9647);
nand U15605 (N_15605,N_7370,N_9486);
xor U15606 (N_15606,N_10334,N_9698);
nor U15607 (N_15607,N_11372,N_11289);
or U15608 (N_15608,N_7209,N_9615);
nand U15609 (N_15609,N_7151,N_11499);
and U15610 (N_15610,N_7596,N_7174);
or U15611 (N_15611,N_10519,N_10217);
or U15612 (N_15612,N_6545,N_6089);
or U15613 (N_15613,N_8369,N_7386);
or U15614 (N_15614,N_9710,N_8618);
and U15615 (N_15615,N_7667,N_9728);
nand U15616 (N_15616,N_8993,N_7493);
nor U15617 (N_15617,N_10124,N_6329);
nor U15618 (N_15618,N_8521,N_6701);
or U15619 (N_15619,N_7287,N_9354);
or U15620 (N_15620,N_8546,N_6386);
nor U15621 (N_15621,N_6838,N_6903);
nand U15622 (N_15622,N_7126,N_10704);
xnor U15623 (N_15623,N_8909,N_9883);
nor U15624 (N_15624,N_6636,N_8044);
or U15625 (N_15625,N_7175,N_7359);
nor U15626 (N_15626,N_9653,N_9394);
or U15627 (N_15627,N_7991,N_7465);
xnor U15628 (N_15628,N_10994,N_9615);
nand U15629 (N_15629,N_7948,N_11768);
or U15630 (N_15630,N_9828,N_10836);
or U15631 (N_15631,N_7142,N_11531);
nand U15632 (N_15632,N_6777,N_10252);
nor U15633 (N_15633,N_10856,N_6177);
nor U15634 (N_15634,N_11682,N_7758);
or U15635 (N_15635,N_8998,N_8104);
and U15636 (N_15636,N_8647,N_11745);
nor U15637 (N_15637,N_6799,N_11601);
or U15638 (N_15638,N_9459,N_7290);
and U15639 (N_15639,N_9692,N_10265);
nand U15640 (N_15640,N_8986,N_6073);
and U15641 (N_15641,N_6660,N_6671);
nand U15642 (N_15642,N_10865,N_9672);
nand U15643 (N_15643,N_7694,N_8341);
or U15644 (N_15644,N_6145,N_10855);
and U15645 (N_15645,N_6073,N_8040);
or U15646 (N_15646,N_11325,N_9113);
nand U15647 (N_15647,N_11713,N_9420);
nand U15648 (N_15648,N_10237,N_9226);
and U15649 (N_15649,N_7854,N_7442);
xor U15650 (N_15650,N_11517,N_11349);
and U15651 (N_15651,N_10835,N_7249);
or U15652 (N_15652,N_8469,N_6148);
nor U15653 (N_15653,N_8619,N_11663);
xnor U15654 (N_15654,N_7241,N_8188);
and U15655 (N_15655,N_7884,N_9855);
or U15656 (N_15656,N_7330,N_10510);
and U15657 (N_15657,N_7948,N_7323);
xor U15658 (N_15658,N_7469,N_7329);
nand U15659 (N_15659,N_7524,N_9735);
nor U15660 (N_15660,N_8672,N_7317);
and U15661 (N_15661,N_10455,N_9238);
or U15662 (N_15662,N_11239,N_8678);
xor U15663 (N_15663,N_8045,N_10679);
or U15664 (N_15664,N_8242,N_6301);
nand U15665 (N_15665,N_11748,N_9307);
or U15666 (N_15666,N_8717,N_8906);
nand U15667 (N_15667,N_6242,N_10791);
xor U15668 (N_15668,N_10247,N_9110);
and U15669 (N_15669,N_10512,N_10706);
xnor U15670 (N_15670,N_10532,N_6985);
xnor U15671 (N_15671,N_11261,N_7597);
and U15672 (N_15672,N_8111,N_8313);
nor U15673 (N_15673,N_11525,N_8484);
xnor U15674 (N_15674,N_8261,N_7625);
or U15675 (N_15675,N_11669,N_6587);
nand U15676 (N_15676,N_6904,N_6480);
xor U15677 (N_15677,N_11355,N_6102);
or U15678 (N_15678,N_7947,N_9542);
xnor U15679 (N_15679,N_10972,N_6666);
nor U15680 (N_15680,N_6167,N_10654);
nor U15681 (N_15681,N_11019,N_11850);
and U15682 (N_15682,N_11829,N_10079);
and U15683 (N_15683,N_7374,N_11131);
or U15684 (N_15684,N_10804,N_6135);
nor U15685 (N_15685,N_8040,N_6872);
nor U15686 (N_15686,N_9830,N_8649);
nand U15687 (N_15687,N_7434,N_10952);
and U15688 (N_15688,N_10940,N_8030);
and U15689 (N_15689,N_8828,N_7312);
nor U15690 (N_15690,N_11693,N_6083);
and U15691 (N_15691,N_9912,N_6228);
or U15692 (N_15692,N_11510,N_6380);
nand U15693 (N_15693,N_9764,N_7287);
xnor U15694 (N_15694,N_6044,N_9711);
nor U15695 (N_15695,N_10469,N_11587);
and U15696 (N_15696,N_7826,N_10419);
or U15697 (N_15697,N_7423,N_7384);
xnor U15698 (N_15698,N_8170,N_9709);
nand U15699 (N_15699,N_6467,N_11542);
or U15700 (N_15700,N_8169,N_6344);
nor U15701 (N_15701,N_7917,N_9308);
and U15702 (N_15702,N_7024,N_6318);
xnor U15703 (N_15703,N_10891,N_7296);
or U15704 (N_15704,N_10805,N_11864);
or U15705 (N_15705,N_8896,N_11531);
or U15706 (N_15706,N_11267,N_10161);
nor U15707 (N_15707,N_7639,N_7368);
or U15708 (N_15708,N_8625,N_11710);
and U15709 (N_15709,N_7701,N_10711);
or U15710 (N_15710,N_7921,N_9714);
nor U15711 (N_15711,N_11556,N_7913);
or U15712 (N_15712,N_9234,N_9475);
or U15713 (N_15713,N_7653,N_11665);
and U15714 (N_15714,N_6041,N_7914);
nand U15715 (N_15715,N_8028,N_9496);
or U15716 (N_15716,N_7792,N_6741);
xnor U15717 (N_15717,N_11246,N_8770);
or U15718 (N_15718,N_11089,N_11860);
or U15719 (N_15719,N_7004,N_7862);
nand U15720 (N_15720,N_8823,N_10199);
nor U15721 (N_15721,N_9112,N_7815);
and U15722 (N_15722,N_8401,N_9030);
xor U15723 (N_15723,N_9150,N_8015);
and U15724 (N_15724,N_9192,N_7925);
nand U15725 (N_15725,N_10881,N_9144);
nand U15726 (N_15726,N_6408,N_8020);
xnor U15727 (N_15727,N_8527,N_6369);
and U15728 (N_15728,N_11210,N_10827);
nor U15729 (N_15729,N_6556,N_6396);
and U15730 (N_15730,N_7017,N_10538);
xnor U15731 (N_15731,N_7562,N_10510);
nor U15732 (N_15732,N_7054,N_6033);
xor U15733 (N_15733,N_11414,N_9030);
nand U15734 (N_15734,N_8017,N_6887);
nand U15735 (N_15735,N_9045,N_11441);
or U15736 (N_15736,N_9749,N_11354);
nor U15737 (N_15737,N_8537,N_6046);
and U15738 (N_15738,N_6770,N_11806);
nand U15739 (N_15739,N_11557,N_10681);
xnor U15740 (N_15740,N_10872,N_11317);
nand U15741 (N_15741,N_9916,N_8128);
nand U15742 (N_15742,N_6696,N_7174);
nor U15743 (N_15743,N_8677,N_10272);
or U15744 (N_15744,N_9213,N_8827);
nor U15745 (N_15745,N_8205,N_6981);
xnor U15746 (N_15746,N_8543,N_9191);
xnor U15747 (N_15747,N_6729,N_7719);
and U15748 (N_15748,N_9722,N_8389);
xnor U15749 (N_15749,N_9442,N_6772);
or U15750 (N_15750,N_10687,N_7355);
nand U15751 (N_15751,N_11077,N_11218);
or U15752 (N_15752,N_8037,N_10518);
nand U15753 (N_15753,N_8152,N_10980);
nor U15754 (N_15754,N_9397,N_10085);
xor U15755 (N_15755,N_6079,N_9633);
or U15756 (N_15756,N_9884,N_8860);
and U15757 (N_15757,N_6463,N_11053);
and U15758 (N_15758,N_7407,N_6599);
nand U15759 (N_15759,N_8235,N_11085);
or U15760 (N_15760,N_7426,N_8170);
nand U15761 (N_15761,N_9120,N_10559);
and U15762 (N_15762,N_6160,N_9589);
xor U15763 (N_15763,N_6734,N_11249);
and U15764 (N_15764,N_11843,N_10138);
or U15765 (N_15765,N_6209,N_9799);
or U15766 (N_15766,N_6956,N_8565);
xnor U15767 (N_15767,N_8455,N_8027);
xnor U15768 (N_15768,N_11991,N_9343);
or U15769 (N_15769,N_9509,N_7692);
and U15770 (N_15770,N_9952,N_10203);
xnor U15771 (N_15771,N_10240,N_7614);
and U15772 (N_15772,N_11116,N_9871);
and U15773 (N_15773,N_8497,N_6019);
or U15774 (N_15774,N_10570,N_6840);
and U15775 (N_15775,N_10186,N_6661);
xor U15776 (N_15776,N_10592,N_7133);
nor U15777 (N_15777,N_11705,N_7410);
nor U15778 (N_15778,N_10447,N_11793);
and U15779 (N_15779,N_11620,N_6742);
and U15780 (N_15780,N_11039,N_6678);
nor U15781 (N_15781,N_11350,N_10656);
and U15782 (N_15782,N_9329,N_11719);
xnor U15783 (N_15783,N_6376,N_11708);
nor U15784 (N_15784,N_10512,N_6435);
and U15785 (N_15785,N_8011,N_9027);
xor U15786 (N_15786,N_9218,N_8787);
nand U15787 (N_15787,N_9582,N_8622);
nand U15788 (N_15788,N_11948,N_11986);
or U15789 (N_15789,N_6219,N_11832);
nand U15790 (N_15790,N_7634,N_6030);
xor U15791 (N_15791,N_9384,N_8590);
and U15792 (N_15792,N_10492,N_11016);
nand U15793 (N_15793,N_11982,N_6015);
nor U15794 (N_15794,N_7915,N_6823);
nand U15795 (N_15795,N_7181,N_9314);
xor U15796 (N_15796,N_6958,N_11865);
nor U15797 (N_15797,N_6398,N_11432);
nand U15798 (N_15798,N_11948,N_10527);
nand U15799 (N_15799,N_7571,N_8777);
nand U15800 (N_15800,N_7238,N_10249);
and U15801 (N_15801,N_7581,N_6580);
or U15802 (N_15802,N_10263,N_7007);
nor U15803 (N_15803,N_11904,N_7092);
nand U15804 (N_15804,N_11704,N_10252);
nor U15805 (N_15805,N_8253,N_7559);
or U15806 (N_15806,N_9041,N_10096);
nor U15807 (N_15807,N_7316,N_10647);
and U15808 (N_15808,N_10985,N_6047);
nor U15809 (N_15809,N_11700,N_10750);
or U15810 (N_15810,N_10601,N_11533);
xnor U15811 (N_15811,N_7532,N_10542);
nor U15812 (N_15812,N_6430,N_6703);
nor U15813 (N_15813,N_10470,N_9788);
xnor U15814 (N_15814,N_11287,N_7363);
nor U15815 (N_15815,N_6470,N_6409);
and U15816 (N_15816,N_11036,N_7702);
and U15817 (N_15817,N_11601,N_9770);
xnor U15818 (N_15818,N_9921,N_9728);
nor U15819 (N_15819,N_10295,N_11191);
xor U15820 (N_15820,N_11502,N_10977);
xnor U15821 (N_15821,N_8660,N_8582);
and U15822 (N_15822,N_8873,N_8631);
and U15823 (N_15823,N_11592,N_11543);
or U15824 (N_15824,N_11480,N_7289);
or U15825 (N_15825,N_9253,N_10300);
or U15826 (N_15826,N_7672,N_7736);
or U15827 (N_15827,N_7981,N_9446);
nand U15828 (N_15828,N_10398,N_7759);
and U15829 (N_15829,N_8460,N_11767);
xnor U15830 (N_15830,N_10512,N_11844);
nand U15831 (N_15831,N_9682,N_9412);
and U15832 (N_15832,N_7666,N_11965);
or U15833 (N_15833,N_8853,N_7667);
nand U15834 (N_15834,N_6060,N_7475);
xor U15835 (N_15835,N_6422,N_9408);
nand U15836 (N_15836,N_7553,N_9268);
or U15837 (N_15837,N_11853,N_11681);
nand U15838 (N_15838,N_6271,N_10687);
nor U15839 (N_15839,N_9140,N_6379);
and U15840 (N_15840,N_11045,N_7561);
and U15841 (N_15841,N_9544,N_8039);
or U15842 (N_15842,N_10424,N_6524);
or U15843 (N_15843,N_9858,N_7787);
nand U15844 (N_15844,N_6734,N_9816);
or U15845 (N_15845,N_8499,N_11398);
nor U15846 (N_15846,N_9854,N_9371);
nor U15847 (N_15847,N_9684,N_10283);
nor U15848 (N_15848,N_11981,N_8179);
and U15849 (N_15849,N_7943,N_11370);
and U15850 (N_15850,N_6320,N_10428);
xnor U15851 (N_15851,N_11661,N_6960);
nor U15852 (N_15852,N_7604,N_9488);
xnor U15853 (N_15853,N_11968,N_10168);
or U15854 (N_15854,N_9109,N_7024);
xnor U15855 (N_15855,N_6909,N_9671);
and U15856 (N_15856,N_10149,N_7836);
or U15857 (N_15857,N_6707,N_7338);
xor U15858 (N_15858,N_6644,N_8826);
and U15859 (N_15859,N_11641,N_8335);
and U15860 (N_15860,N_7140,N_6037);
or U15861 (N_15861,N_11674,N_11897);
nor U15862 (N_15862,N_8029,N_6867);
and U15863 (N_15863,N_11258,N_7142);
and U15864 (N_15864,N_7205,N_11012);
and U15865 (N_15865,N_11557,N_11993);
nor U15866 (N_15866,N_6613,N_9948);
and U15867 (N_15867,N_8167,N_10512);
xnor U15868 (N_15868,N_8602,N_11733);
xnor U15869 (N_15869,N_8732,N_8794);
xor U15870 (N_15870,N_10697,N_6106);
and U15871 (N_15871,N_10654,N_9870);
and U15872 (N_15872,N_7207,N_11437);
nor U15873 (N_15873,N_6688,N_11955);
nand U15874 (N_15874,N_11652,N_10947);
xnor U15875 (N_15875,N_8417,N_10987);
nand U15876 (N_15876,N_10856,N_9392);
or U15877 (N_15877,N_6114,N_11491);
or U15878 (N_15878,N_7856,N_7795);
xnor U15879 (N_15879,N_9911,N_6713);
nor U15880 (N_15880,N_8131,N_8001);
xnor U15881 (N_15881,N_8393,N_8242);
nor U15882 (N_15882,N_11953,N_7441);
nor U15883 (N_15883,N_7753,N_7156);
nor U15884 (N_15884,N_9772,N_8695);
and U15885 (N_15885,N_10476,N_8847);
xor U15886 (N_15886,N_9388,N_6654);
xnor U15887 (N_15887,N_10584,N_9511);
xor U15888 (N_15888,N_10122,N_8290);
or U15889 (N_15889,N_9253,N_11313);
nor U15890 (N_15890,N_7714,N_11142);
and U15891 (N_15891,N_9904,N_8687);
xnor U15892 (N_15892,N_8181,N_10319);
or U15893 (N_15893,N_6496,N_6599);
and U15894 (N_15894,N_7613,N_10814);
nor U15895 (N_15895,N_9508,N_6207);
xnor U15896 (N_15896,N_6012,N_6510);
or U15897 (N_15897,N_8026,N_8145);
xnor U15898 (N_15898,N_6764,N_10331);
nor U15899 (N_15899,N_6220,N_11543);
xor U15900 (N_15900,N_7232,N_6364);
or U15901 (N_15901,N_9076,N_10946);
nor U15902 (N_15902,N_7755,N_7013);
or U15903 (N_15903,N_10022,N_6143);
nand U15904 (N_15904,N_7102,N_9669);
xnor U15905 (N_15905,N_9446,N_9896);
or U15906 (N_15906,N_10686,N_7232);
nor U15907 (N_15907,N_6922,N_8509);
and U15908 (N_15908,N_9827,N_10851);
and U15909 (N_15909,N_9283,N_7052);
nor U15910 (N_15910,N_8408,N_8269);
xnor U15911 (N_15911,N_7413,N_6481);
nand U15912 (N_15912,N_11861,N_7011);
nand U15913 (N_15913,N_9208,N_11594);
nand U15914 (N_15914,N_9000,N_8816);
xor U15915 (N_15915,N_9150,N_7197);
xor U15916 (N_15916,N_11675,N_6106);
and U15917 (N_15917,N_6062,N_7766);
or U15918 (N_15918,N_6435,N_10854);
xor U15919 (N_15919,N_7179,N_8461);
xor U15920 (N_15920,N_10072,N_9978);
and U15921 (N_15921,N_8242,N_11790);
nand U15922 (N_15922,N_8657,N_10851);
xnor U15923 (N_15923,N_11432,N_11637);
xor U15924 (N_15924,N_9303,N_8031);
nand U15925 (N_15925,N_10186,N_8773);
nand U15926 (N_15926,N_10193,N_7175);
nand U15927 (N_15927,N_6758,N_7277);
nor U15928 (N_15928,N_9894,N_10196);
or U15929 (N_15929,N_11735,N_11436);
and U15930 (N_15930,N_7157,N_10744);
nor U15931 (N_15931,N_7810,N_8928);
nand U15932 (N_15932,N_10862,N_9285);
nand U15933 (N_15933,N_6942,N_6341);
nor U15934 (N_15934,N_8063,N_11543);
and U15935 (N_15935,N_6213,N_9914);
nand U15936 (N_15936,N_8187,N_9217);
nor U15937 (N_15937,N_6667,N_11419);
nor U15938 (N_15938,N_9879,N_10455);
xnor U15939 (N_15939,N_7073,N_7110);
or U15940 (N_15940,N_6521,N_9463);
xor U15941 (N_15941,N_6468,N_10155);
or U15942 (N_15942,N_11750,N_6485);
nand U15943 (N_15943,N_11939,N_9795);
xor U15944 (N_15944,N_10972,N_6902);
and U15945 (N_15945,N_10752,N_7315);
nor U15946 (N_15946,N_8776,N_7359);
nor U15947 (N_15947,N_6280,N_6457);
xnor U15948 (N_15948,N_6671,N_6081);
nor U15949 (N_15949,N_6208,N_8757);
and U15950 (N_15950,N_11455,N_6796);
nor U15951 (N_15951,N_8907,N_10432);
nor U15952 (N_15952,N_8771,N_6593);
nor U15953 (N_15953,N_9625,N_7715);
or U15954 (N_15954,N_11792,N_9568);
xor U15955 (N_15955,N_9958,N_10634);
or U15956 (N_15956,N_10992,N_10393);
nor U15957 (N_15957,N_6937,N_9499);
nor U15958 (N_15958,N_9497,N_6820);
xnor U15959 (N_15959,N_11204,N_7899);
xnor U15960 (N_15960,N_10643,N_9748);
nand U15961 (N_15961,N_9841,N_6691);
xor U15962 (N_15962,N_10004,N_8999);
or U15963 (N_15963,N_10177,N_10918);
and U15964 (N_15964,N_7317,N_7837);
nor U15965 (N_15965,N_9311,N_11460);
xor U15966 (N_15966,N_8933,N_9811);
or U15967 (N_15967,N_8142,N_6793);
nand U15968 (N_15968,N_6782,N_7692);
and U15969 (N_15969,N_9557,N_8067);
nor U15970 (N_15970,N_7463,N_6079);
nand U15971 (N_15971,N_11801,N_10985);
xnor U15972 (N_15972,N_6397,N_10007);
xnor U15973 (N_15973,N_11017,N_11057);
xor U15974 (N_15974,N_11406,N_8401);
xor U15975 (N_15975,N_10496,N_10953);
nand U15976 (N_15976,N_9009,N_8964);
xnor U15977 (N_15977,N_9642,N_7564);
nor U15978 (N_15978,N_8601,N_6154);
xnor U15979 (N_15979,N_7258,N_8484);
and U15980 (N_15980,N_6962,N_9295);
nor U15981 (N_15981,N_9158,N_7796);
xor U15982 (N_15982,N_7325,N_6975);
nand U15983 (N_15983,N_8455,N_10702);
nor U15984 (N_15984,N_11818,N_8075);
nor U15985 (N_15985,N_7584,N_8610);
and U15986 (N_15986,N_9190,N_9133);
xnor U15987 (N_15987,N_11008,N_7310);
and U15988 (N_15988,N_11464,N_7525);
and U15989 (N_15989,N_7155,N_8906);
xnor U15990 (N_15990,N_10005,N_7941);
nand U15991 (N_15991,N_9085,N_8268);
nand U15992 (N_15992,N_7195,N_6978);
nand U15993 (N_15993,N_6454,N_9770);
or U15994 (N_15994,N_10691,N_8131);
nor U15995 (N_15995,N_6153,N_9736);
nor U15996 (N_15996,N_9213,N_6000);
and U15997 (N_15997,N_10009,N_7406);
nor U15998 (N_15998,N_9299,N_7127);
nand U15999 (N_15999,N_8917,N_10802);
nand U16000 (N_16000,N_11813,N_8879);
xnor U16001 (N_16001,N_10146,N_6702);
xnor U16002 (N_16002,N_11221,N_6130);
or U16003 (N_16003,N_7548,N_6821);
xnor U16004 (N_16004,N_9689,N_10042);
or U16005 (N_16005,N_7533,N_7097);
nor U16006 (N_16006,N_10675,N_8870);
or U16007 (N_16007,N_11881,N_9081);
xnor U16008 (N_16008,N_8843,N_7675);
and U16009 (N_16009,N_8233,N_9664);
and U16010 (N_16010,N_8541,N_6541);
xor U16011 (N_16011,N_8341,N_9220);
nand U16012 (N_16012,N_6472,N_8833);
nand U16013 (N_16013,N_8421,N_11253);
or U16014 (N_16014,N_8520,N_6911);
nor U16015 (N_16015,N_8808,N_10368);
xor U16016 (N_16016,N_9124,N_10278);
or U16017 (N_16017,N_6501,N_9702);
or U16018 (N_16018,N_9407,N_9064);
and U16019 (N_16019,N_8161,N_7533);
or U16020 (N_16020,N_11629,N_9261);
or U16021 (N_16021,N_7344,N_10721);
and U16022 (N_16022,N_11077,N_9020);
or U16023 (N_16023,N_8217,N_10062);
nor U16024 (N_16024,N_7457,N_8013);
or U16025 (N_16025,N_9250,N_7106);
or U16026 (N_16026,N_7683,N_10270);
or U16027 (N_16027,N_6276,N_11082);
xor U16028 (N_16028,N_7075,N_6378);
xor U16029 (N_16029,N_6389,N_10423);
and U16030 (N_16030,N_6709,N_9098);
and U16031 (N_16031,N_11891,N_8443);
and U16032 (N_16032,N_6481,N_7058);
and U16033 (N_16033,N_11302,N_7922);
or U16034 (N_16034,N_10240,N_6016);
and U16035 (N_16035,N_6172,N_8563);
xor U16036 (N_16036,N_9258,N_9047);
nand U16037 (N_16037,N_7012,N_6713);
and U16038 (N_16038,N_11139,N_8740);
nand U16039 (N_16039,N_7211,N_7911);
and U16040 (N_16040,N_8719,N_8679);
and U16041 (N_16041,N_8132,N_11409);
nand U16042 (N_16042,N_6878,N_10949);
or U16043 (N_16043,N_6938,N_10299);
xnor U16044 (N_16044,N_7765,N_8827);
nor U16045 (N_16045,N_11981,N_6133);
xor U16046 (N_16046,N_8469,N_6626);
xnor U16047 (N_16047,N_9064,N_10947);
nand U16048 (N_16048,N_9094,N_9128);
and U16049 (N_16049,N_8675,N_7224);
nor U16050 (N_16050,N_7719,N_8412);
nand U16051 (N_16051,N_6900,N_8338);
and U16052 (N_16052,N_7247,N_8865);
nor U16053 (N_16053,N_6299,N_6974);
nand U16054 (N_16054,N_6498,N_6839);
and U16055 (N_16055,N_6868,N_6159);
or U16056 (N_16056,N_11196,N_9706);
xor U16057 (N_16057,N_8335,N_9572);
xnor U16058 (N_16058,N_10984,N_10439);
xnor U16059 (N_16059,N_9127,N_11118);
nor U16060 (N_16060,N_7536,N_8466);
and U16061 (N_16061,N_6005,N_8705);
and U16062 (N_16062,N_8562,N_6358);
nor U16063 (N_16063,N_6262,N_10537);
and U16064 (N_16064,N_7593,N_7097);
and U16065 (N_16065,N_6031,N_10855);
nor U16066 (N_16066,N_8837,N_11844);
nand U16067 (N_16067,N_11722,N_11267);
nor U16068 (N_16068,N_8991,N_6037);
nor U16069 (N_16069,N_10395,N_6919);
and U16070 (N_16070,N_11176,N_8142);
nand U16071 (N_16071,N_7043,N_6879);
and U16072 (N_16072,N_8940,N_9967);
nand U16073 (N_16073,N_7475,N_8856);
xor U16074 (N_16074,N_8418,N_11660);
or U16075 (N_16075,N_6491,N_8037);
or U16076 (N_16076,N_11366,N_9609);
nor U16077 (N_16077,N_11698,N_8813);
and U16078 (N_16078,N_8193,N_11336);
nand U16079 (N_16079,N_6345,N_11592);
and U16080 (N_16080,N_6837,N_7831);
xnor U16081 (N_16081,N_8058,N_8607);
or U16082 (N_16082,N_9936,N_7885);
nand U16083 (N_16083,N_7841,N_8346);
nor U16084 (N_16084,N_10429,N_8904);
nand U16085 (N_16085,N_6761,N_9947);
nor U16086 (N_16086,N_6468,N_11257);
nand U16087 (N_16087,N_11698,N_6806);
and U16088 (N_16088,N_10685,N_6403);
nor U16089 (N_16089,N_6605,N_7078);
xnor U16090 (N_16090,N_11496,N_9336);
nor U16091 (N_16091,N_6970,N_6015);
or U16092 (N_16092,N_7923,N_10150);
xnor U16093 (N_16093,N_6013,N_6190);
and U16094 (N_16094,N_7362,N_8234);
nor U16095 (N_16095,N_6297,N_10494);
nor U16096 (N_16096,N_8907,N_10116);
or U16097 (N_16097,N_6296,N_7259);
nand U16098 (N_16098,N_10067,N_6907);
or U16099 (N_16099,N_8820,N_7370);
and U16100 (N_16100,N_11795,N_6770);
nor U16101 (N_16101,N_11561,N_8078);
xnor U16102 (N_16102,N_8110,N_7329);
nor U16103 (N_16103,N_6149,N_8699);
nor U16104 (N_16104,N_7226,N_11868);
nand U16105 (N_16105,N_8645,N_10240);
or U16106 (N_16106,N_6927,N_7554);
or U16107 (N_16107,N_10962,N_7742);
nor U16108 (N_16108,N_10820,N_8261);
nand U16109 (N_16109,N_6851,N_10029);
or U16110 (N_16110,N_11102,N_11867);
and U16111 (N_16111,N_6363,N_7215);
and U16112 (N_16112,N_6135,N_7326);
and U16113 (N_16113,N_7085,N_10902);
nor U16114 (N_16114,N_6861,N_7019);
nand U16115 (N_16115,N_7327,N_9053);
or U16116 (N_16116,N_6467,N_11544);
nand U16117 (N_16117,N_7966,N_6461);
or U16118 (N_16118,N_10264,N_7706);
nor U16119 (N_16119,N_10349,N_9270);
nand U16120 (N_16120,N_6182,N_11749);
xnor U16121 (N_16121,N_6619,N_11259);
xnor U16122 (N_16122,N_9965,N_6905);
nand U16123 (N_16123,N_11814,N_6932);
nor U16124 (N_16124,N_11813,N_9842);
or U16125 (N_16125,N_10059,N_9534);
nor U16126 (N_16126,N_11391,N_11581);
and U16127 (N_16127,N_11554,N_11031);
and U16128 (N_16128,N_6370,N_10396);
xnor U16129 (N_16129,N_7396,N_11847);
xnor U16130 (N_16130,N_11881,N_6448);
or U16131 (N_16131,N_8867,N_9842);
xnor U16132 (N_16132,N_10236,N_10486);
xnor U16133 (N_16133,N_11773,N_11962);
xor U16134 (N_16134,N_7440,N_10596);
nor U16135 (N_16135,N_9486,N_10824);
xnor U16136 (N_16136,N_9446,N_9916);
xor U16137 (N_16137,N_8881,N_6092);
nand U16138 (N_16138,N_7440,N_10570);
nand U16139 (N_16139,N_9062,N_7876);
or U16140 (N_16140,N_10924,N_9598);
nor U16141 (N_16141,N_11142,N_8041);
and U16142 (N_16142,N_6934,N_6678);
and U16143 (N_16143,N_10476,N_11997);
and U16144 (N_16144,N_11076,N_7126);
nand U16145 (N_16145,N_9035,N_11574);
nand U16146 (N_16146,N_8996,N_8104);
or U16147 (N_16147,N_6940,N_10859);
and U16148 (N_16148,N_10480,N_11952);
and U16149 (N_16149,N_7387,N_7311);
nand U16150 (N_16150,N_6591,N_10216);
and U16151 (N_16151,N_7835,N_11664);
xnor U16152 (N_16152,N_10933,N_6715);
or U16153 (N_16153,N_6756,N_9621);
nand U16154 (N_16154,N_10540,N_6781);
or U16155 (N_16155,N_6852,N_8079);
nand U16156 (N_16156,N_9351,N_6451);
or U16157 (N_16157,N_8377,N_11255);
nor U16158 (N_16158,N_8284,N_7885);
nor U16159 (N_16159,N_9268,N_9829);
nand U16160 (N_16160,N_6889,N_7921);
xnor U16161 (N_16161,N_11909,N_9641);
and U16162 (N_16162,N_11940,N_9730);
xor U16163 (N_16163,N_10795,N_10748);
nand U16164 (N_16164,N_7395,N_7693);
and U16165 (N_16165,N_6552,N_9523);
and U16166 (N_16166,N_8359,N_9647);
nor U16167 (N_16167,N_9499,N_7965);
and U16168 (N_16168,N_11716,N_11534);
or U16169 (N_16169,N_6893,N_8276);
and U16170 (N_16170,N_10094,N_9727);
nand U16171 (N_16171,N_6824,N_9426);
nand U16172 (N_16172,N_9973,N_11342);
xnor U16173 (N_16173,N_8591,N_7620);
nor U16174 (N_16174,N_9978,N_10919);
xnor U16175 (N_16175,N_9527,N_11653);
nor U16176 (N_16176,N_8794,N_8866);
or U16177 (N_16177,N_6573,N_10534);
or U16178 (N_16178,N_6835,N_6828);
xnor U16179 (N_16179,N_7996,N_10991);
xor U16180 (N_16180,N_9317,N_8245);
and U16181 (N_16181,N_10391,N_7478);
nand U16182 (N_16182,N_7877,N_7442);
and U16183 (N_16183,N_7378,N_6302);
or U16184 (N_16184,N_10945,N_8636);
xnor U16185 (N_16185,N_10412,N_10569);
or U16186 (N_16186,N_7144,N_11790);
xor U16187 (N_16187,N_7048,N_10898);
nand U16188 (N_16188,N_6225,N_11215);
and U16189 (N_16189,N_9960,N_9662);
or U16190 (N_16190,N_6276,N_9257);
or U16191 (N_16191,N_9645,N_10303);
or U16192 (N_16192,N_8595,N_7569);
or U16193 (N_16193,N_7851,N_9980);
nand U16194 (N_16194,N_10025,N_6836);
and U16195 (N_16195,N_7062,N_8176);
nand U16196 (N_16196,N_7076,N_7888);
nand U16197 (N_16197,N_8332,N_6609);
and U16198 (N_16198,N_6840,N_8184);
nor U16199 (N_16199,N_8942,N_11693);
or U16200 (N_16200,N_7361,N_8580);
and U16201 (N_16201,N_10880,N_6640);
xnor U16202 (N_16202,N_10845,N_11602);
and U16203 (N_16203,N_9109,N_10294);
or U16204 (N_16204,N_6084,N_8824);
or U16205 (N_16205,N_10021,N_9078);
nand U16206 (N_16206,N_11639,N_8462);
nand U16207 (N_16207,N_6221,N_8404);
nor U16208 (N_16208,N_9853,N_7786);
nand U16209 (N_16209,N_11808,N_9993);
and U16210 (N_16210,N_11931,N_8833);
or U16211 (N_16211,N_11466,N_6951);
or U16212 (N_16212,N_7781,N_6883);
xnor U16213 (N_16213,N_9460,N_7129);
xor U16214 (N_16214,N_7401,N_10597);
nand U16215 (N_16215,N_9575,N_11144);
nand U16216 (N_16216,N_8159,N_11635);
nor U16217 (N_16217,N_6337,N_6572);
or U16218 (N_16218,N_7487,N_7403);
nand U16219 (N_16219,N_6697,N_6015);
xnor U16220 (N_16220,N_11936,N_11488);
xor U16221 (N_16221,N_7238,N_10290);
xor U16222 (N_16222,N_11003,N_10908);
nor U16223 (N_16223,N_11579,N_8827);
nor U16224 (N_16224,N_8546,N_11304);
xnor U16225 (N_16225,N_8549,N_9582);
or U16226 (N_16226,N_9064,N_11886);
nor U16227 (N_16227,N_8116,N_8728);
nor U16228 (N_16228,N_11847,N_6038);
nor U16229 (N_16229,N_10107,N_10345);
xor U16230 (N_16230,N_7248,N_9571);
or U16231 (N_16231,N_11535,N_9603);
nor U16232 (N_16232,N_11154,N_9262);
and U16233 (N_16233,N_7298,N_7610);
xor U16234 (N_16234,N_8217,N_9657);
nand U16235 (N_16235,N_11206,N_9779);
xor U16236 (N_16236,N_8020,N_7687);
or U16237 (N_16237,N_9346,N_9602);
nand U16238 (N_16238,N_10786,N_6925);
nand U16239 (N_16239,N_11211,N_7040);
nand U16240 (N_16240,N_9728,N_6616);
and U16241 (N_16241,N_9198,N_7507);
xor U16242 (N_16242,N_11254,N_8261);
and U16243 (N_16243,N_9931,N_10350);
nand U16244 (N_16244,N_8410,N_9892);
nand U16245 (N_16245,N_9686,N_8934);
and U16246 (N_16246,N_6475,N_6278);
nand U16247 (N_16247,N_6455,N_6605);
nor U16248 (N_16248,N_8044,N_6326);
and U16249 (N_16249,N_10479,N_10492);
xnor U16250 (N_16250,N_10565,N_9416);
xor U16251 (N_16251,N_8840,N_7603);
nor U16252 (N_16252,N_11808,N_9603);
xor U16253 (N_16253,N_8342,N_6534);
nand U16254 (N_16254,N_6284,N_10686);
xnor U16255 (N_16255,N_8001,N_11767);
and U16256 (N_16256,N_7224,N_8339);
nor U16257 (N_16257,N_8722,N_7090);
or U16258 (N_16258,N_11716,N_8153);
xor U16259 (N_16259,N_7208,N_11146);
and U16260 (N_16260,N_7779,N_11752);
nor U16261 (N_16261,N_9421,N_7435);
xor U16262 (N_16262,N_8953,N_9154);
nor U16263 (N_16263,N_9225,N_6166);
xor U16264 (N_16264,N_7914,N_8289);
nor U16265 (N_16265,N_8982,N_7933);
and U16266 (N_16266,N_6936,N_7267);
xnor U16267 (N_16267,N_10793,N_10964);
nor U16268 (N_16268,N_6032,N_9204);
or U16269 (N_16269,N_6155,N_7518);
nand U16270 (N_16270,N_7758,N_11254);
xnor U16271 (N_16271,N_8667,N_6559);
nand U16272 (N_16272,N_9905,N_6525);
xnor U16273 (N_16273,N_10011,N_9400);
and U16274 (N_16274,N_10163,N_8272);
or U16275 (N_16275,N_7835,N_8752);
or U16276 (N_16276,N_7757,N_10556);
and U16277 (N_16277,N_7813,N_8535);
and U16278 (N_16278,N_8835,N_7770);
nor U16279 (N_16279,N_11081,N_11720);
or U16280 (N_16280,N_6861,N_6811);
nor U16281 (N_16281,N_10293,N_10382);
nor U16282 (N_16282,N_8252,N_11977);
nand U16283 (N_16283,N_6707,N_6842);
nand U16284 (N_16284,N_10272,N_7301);
and U16285 (N_16285,N_9424,N_7727);
xor U16286 (N_16286,N_7268,N_11449);
xnor U16287 (N_16287,N_10420,N_10127);
xnor U16288 (N_16288,N_11062,N_6097);
nor U16289 (N_16289,N_11104,N_11277);
nand U16290 (N_16290,N_11115,N_11834);
or U16291 (N_16291,N_8882,N_9987);
nor U16292 (N_16292,N_10273,N_8607);
xnor U16293 (N_16293,N_6127,N_11995);
or U16294 (N_16294,N_6505,N_7250);
nand U16295 (N_16295,N_7898,N_8972);
or U16296 (N_16296,N_10456,N_9030);
nor U16297 (N_16297,N_6481,N_9756);
nand U16298 (N_16298,N_7276,N_6901);
nand U16299 (N_16299,N_11713,N_6434);
or U16300 (N_16300,N_8912,N_10586);
xor U16301 (N_16301,N_8750,N_6208);
nor U16302 (N_16302,N_8418,N_6029);
or U16303 (N_16303,N_11753,N_10001);
and U16304 (N_16304,N_9728,N_8859);
xnor U16305 (N_16305,N_9110,N_7942);
or U16306 (N_16306,N_10141,N_9033);
and U16307 (N_16307,N_8134,N_8518);
nand U16308 (N_16308,N_8113,N_9188);
nor U16309 (N_16309,N_9816,N_7006);
nand U16310 (N_16310,N_8714,N_8005);
xor U16311 (N_16311,N_10666,N_6144);
or U16312 (N_16312,N_8348,N_9728);
xor U16313 (N_16313,N_10112,N_11864);
xor U16314 (N_16314,N_8920,N_7381);
nor U16315 (N_16315,N_11212,N_11011);
xnor U16316 (N_16316,N_9602,N_7269);
or U16317 (N_16317,N_10673,N_10814);
nand U16318 (N_16318,N_10298,N_6049);
nor U16319 (N_16319,N_8154,N_11264);
nor U16320 (N_16320,N_8573,N_8353);
xnor U16321 (N_16321,N_10108,N_8552);
and U16322 (N_16322,N_8096,N_9549);
or U16323 (N_16323,N_11383,N_10496);
and U16324 (N_16324,N_8751,N_7642);
nor U16325 (N_16325,N_8468,N_11821);
nor U16326 (N_16326,N_8718,N_9849);
nand U16327 (N_16327,N_6253,N_9831);
or U16328 (N_16328,N_11115,N_10456);
and U16329 (N_16329,N_11800,N_11838);
nand U16330 (N_16330,N_9008,N_8703);
nand U16331 (N_16331,N_6411,N_8485);
nand U16332 (N_16332,N_8576,N_8905);
nor U16333 (N_16333,N_6802,N_9644);
nor U16334 (N_16334,N_7255,N_8470);
nor U16335 (N_16335,N_9937,N_9524);
xor U16336 (N_16336,N_9391,N_7247);
nor U16337 (N_16337,N_9923,N_6320);
and U16338 (N_16338,N_8115,N_10400);
nand U16339 (N_16339,N_7859,N_11347);
and U16340 (N_16340,N_10784,N_8472);
xor U16341 (N_16341,N_6695,N_9707);
xor U16342 (N_16342,N_9837,N_6172);
or U16343 (N_16343,N_8519,N_6681);
or U16344 (N_16344,N_9554,N_7259);
and U16345 (N_16345,N_7157,N_7656);
nor U16346 (N_16346,N_7157,N_7365);
nor U16347 (N_16347,N_8742,N_11623);
nor U16348 (N_16348,N_6117,N_8364);
or U16349 (N_16349,N_10289,N_9211);
nor U16350 (N_16350,N_7647,N_10152);
xor U16351 (N_16351,N_7376,N_6389);
and U16352 (N_16352,N_9661,N_7676);
nand U16353 (N_16353,N_6841,N_6600);
or U16354 (N_16354,N_11560,N_9410);
or U16355 (N_16355,N_6422,N_7234);
and U16356 (N_16356,N_10595,N_9420);
nand U16357 (N_16357,N_6056,N_11837);
or U16358 (N_16358,N_6572,N_7110);
nor U16359 (N_16359,N_11572,N_10635);
nand U16360 (N_16360,N_9798,N_7746);
or U16361 (N_16361,N_11110,N_7252);
or U16362 (N_16362,N_8161,N_6410);
xnor U16363 (N_16363,N_10538,N_9394);
or U16364 (N_16364,N_8802,N_7136);
nand U16365 (N_16365,N_6639,N_8590);
nand U16366 (N_16366,N_6569,N_6286);
nand U16367 (N_16367,N_9573,N_9343);
xnor U16368 (N_16368,N_6524,N_9921);
and U16369 (N_16369,N_11959,N_8052);
nand U16370 (N_16370,N_7151,N_11053);
and U16371 (N_16371,N_7170,N_11412);
and U16372 (N_16372,N_6523,N_10242);
nor U16373 (N_16373,N_7883,N_11408);
nor U16374 (N_16374,N_10559,N_9034);
and U16375 (N_16375,N_9693,N_7622);
and U16376 (N_16376,N_8881,N_7719);
and U16377 (N_16377,N_9556,N_11656);
nor U16378 (N_16378,N_8513,N_8861);
nand U16379 (N_16379,N_6814,N_11654);
nor U16380 (N_16380,N_8845,N_8661);
nand U16381 (N_16381,N_6759,N_10744);
nand U16382 (N_16382,N_10629,N_6936);
nand U16383 (N_16383,N_8671,N_7367);
and U16384 (N_16384,N_10078,N_10234);
nor U16385 (N_16385,N_10922,N_6461);
nand U16386 (N_16386,N_9400,N_6587);
or U16387 (N_16387,N_6727,N_9976);
or U16388 (N_16388,N_9007,N_7543);
xor U16389 (N_16389,N_9135,N_10948);
and U16390 (N_16390,N_8398,N_9869);
nor U16391 (N_16391,N_11653,N_6887);
xnor U16392 (N_16392,N_6930,N_9590);
and U16393 (N_16393,N_7283,N_8505);
and U16394 (N_16394,N_9070,N_10736);
or U16395 (N_16395,N_7856,N_11844);
xor U16396 (N_16396,N_7707,N_8437);
xnor U16397 (N_16397,N_7929,N_10070);
and U16398 (N_16398,N_11258,N_6690);
xor U16399 (N_16399,N_10129,N_11969);
and U16400 (N_16400,N_11572,N_6635);
and U16401 (N_16401,N_8577,N_6776);
nor U16402 (N_16402,N_9423,N_7408);
xor U16403 (N_16403,N_7331,N_8363);
nand U16404 (N_16404,N_10231,N_9056);
or U16405 (N_16405,N_11163,N_10248);
and U16406 (N_16406,N_6650,N_10822);
xnor U16407 (N_16407,N_9438,N_9335);
or U16408 (N_16408,N_7338,N_9849);
and U16409 (N_16409,N_9909,N_11283);
xor U16410 (N_16410,N_9973,N_10192);
and U16411 (N_16411,N_9394,N_9085);
and U16412 (N_16412,N_8105,N_11174);
nor U16413 (N_16413,N_7745,N_7070);
nor U16414 (N_16414,N_7978,N_11680);
xor U16415 (N_16415,N_7665,N_10346);
or U16416 (N_16416,N_6423,N_6485);
nor U16417 (N_16417,N_6220,N_8046);
xnor U16418 (N_16418,N_8221,N_6898);
nor U16419 (N_16419,N_7210,N_10368);
or U16420 (N_16420,N_6402,N_7779);
nand U16421 (N_16421,N_6194,N_6870);
xor U16422 (N_16422,N_7456,N_11174);
and U16423 (N_16423,N_6896,N_7701);
xnor U16424 (N_16424,N_11306,N_8545);
and U16425 (N_16425,N_10426,N_6769);
xor U16426 (N_16426,N_7869,N_8960);
or U16427 (N_16427,N_7993,N_6077);
and U16428 (N_16428,N_8181,N_11980);
or U16429 (N_16429,N_9592,N_9169);
xor U16430 (N_16430,N_8961,N_6988);
and U16431 (N_16431,N_7994,N_7624);
or U16432 (N_16432,N_6567,N_6435);
nor U16433 (N_16433,N_7755,N_8115);
xor U16434 (N_16434,N_9134,N_8246);
nand U16435 (N_16435,N_7298,N_7647);
nor U16436 (N_16436,N_6904,N_9312);
or U16437 (N_16437,N_9845,N_9146);
nor U16438 (N_16438,N_6926,N_7281);
nand U16439 (N_16439,N_10239,N_6580);
xnor U16440 (N_16440,N_9850,N_7881);
nor U16441 (N_16441,N_6682,N_7263);
nor U16442 (N_16442,N_7977,N_9316);
xor U16443 (N_16443,N_7738,N_11734);
or U16444 (N_16444,N_7567,N_7089);
or U16445 (N_16445,N_11565,N_9641);
nor U16446 (N_16446,N_11090,N_8798);
xor U16447 (N_16447,N_10454,N_10415);
or U16448 (N_16448,N_10128,N_7913);
and U16449 (N_16449,N_7416,N_10316);
nor U16450 (N_16450,N_9996,N_8030);
nor U16451 (N_16451,N_10034,N_7237);
and U16452 (N_16452,N_6828,N_11604);
and U16453 (N_16453,N_8154,N_8931);
and U16454 (N_16454,N_10094,N_11634);
nor U16455 (N_16455,N_9013,N_7729);
or U16456 (N_16456,N_7355,N_7399);
or U16457 (N_16457,N_11909,N_7348);
and U16458 (N_16458,N_11168,N_7037);
nand U16459 (N_16459,N_9917,N_6040);
nor U16460 (N_16460,N_7273,N_11851);
or U16461 (N_16461,N_8529,N_7252);
or U16462 (N_16462,N_7031,N_6599);
and U16463 (N_16463,N_8262,N_10021);
and U16464 (N_16464,N_6144,N_10633);
and U16465 (N_16465,N_10465,N_7326);
and U16466 (N_16466,N_8854,N_7155);
xnor U16467 (N_16467,N_8762,N_7918);
nor U16468 (N_16468,N_10046,N_11936);
xnor U16469 (N_16469,N_10906,N_8384);
and U16470 (N_16470,N_6073,N_6368);
and U16471 (N_16471,N_10264,N_6256);
xor U16472 (N_16472,N_6017,N_9680);
nand U16473 (N_16473,N_10083,N_7091);
or U16474 (N_16474,N_6187,N_7375);
and U16475 (N_16475,N_7909,N_10179);
nor U16476 (N_16476,N_8715,N_11017);
or U16477 (N_16477,N_7604,N_9353);
xnor U16478 (N_16478,N_8394,N_9901);
nand U16479 (N_16479,N_9008,N_7694);
nor U16480 (N_16480,N_11153,N_10939);
nor U16481 (N_16481,N_11445,N_6435);
nand U16482 (N_16482,N_10639,N_10721);
and U16483 (N_16483,N_7322,N_9164);
nor U16484 (N_16484,N_8689,N_6360);
nand U16485 (N_16485,N_6318,N_8678);
or U16486 (N_16486,N_6679,N_7857);
and U16487 (N_16487,N_10926,N_10436);
xnor U16488 (N_16488,N_11090,N_9554);
nor U16489 (N_16489,N_10590,N_6726);
or U16490 (N_16490,N_9479,N_6642);
or U16491 (N_16491,N_9583,N_7817);
nor U16492 (N_16492,N_9044,N_7330);
nand U16493 (N_16493,N_11156,N_11839);
nand U16494 (N_16494,N_9523,N_7517);
xor U16495 (N_16495,N_11394,N_6876);
and U16496 (N_16496,N_11463,N_6442);
nand U16497 (N_16497,N_7783,N_10292);
xnor U16498 (N_16498,N_6624,N_9976);
nand U16499 (N_16499,N_10628,N_11698);
nor U16500 (N_16500,N_9503,N_6829);
and U16501 (N_16501,N_9712,N_6918);
nand U16502 (N_16502,N_7687,N_6175);
and U16503 (N_16503,N_7039,N_7214);
and U16504 (N_16504,N_11611,N_7186);
and U16505 (N_16505,N_10432,N_7482);
nor U16506 (N_16506,N_10188,N_11549);
and U16507 (N_16507,N_10693,N_10410);
and U16508 (N_16508,N_10394,N_11780);
nor U16509 (N_16509,N_10158,N_6559);
nor U16510 (N_16510,N_7432,N_10574);
and U16511 (N_16511,N_9124,N_11684);
nor U16512 (N_16512,N_10741,N_9727);
or U16513 (N_16513,N_11675,N_10055);
or U16514 (N_16514,N_7296,N_6950);
or U16515 (N_16515,N_7584,N_11594);
nand U16516 (N_16516,N_9134,N_10253);
nor U16517 (N_16517,N_6388,N_11180);
nand U16518 (N_16518,N_8717,N_8732);
nor U16519 (N_16519,N_10855,N_9455);
and U16520 (N_16520,N_8898,N_6827);
xnor U16521 (N_16521,N_9407,N_6727);
nor U16522 (N_16522,N_6486,N_10071);
xor U16523 (N_16523,N_10465,N_9145);
and U16524 (N_16524,N_6565,N_7802);
nor U16525 (N_16525,N_10668,N_7519);
nand U16526 (N_16526,N_11337,N_10079);
nand U16527 (N_16527,N_6692,N_9518);
xnor U16528 (N_16528,N_9688,N_9678);
xnor U16529 (N_16529,N_10464,N_6050);
nor U16530 (N_16530,N_11167,N_8458);
or U16531 (N_16531,N_8410,N_6351);
or U16532 (N_16532,N_10585,N_6615);
or U16533 (N_16533,N_10606,N_7964);
or U16534 (N_16534,N_11961,N_8690);
and U16535 (N_16535,N_10009,N_6970);
and U16536 (N_16536,N_11216,N_10118);
nand U16537 (N_16537,N_9155,N_6298);
xnor U16538 (N_16538,N_8275,N_6266);
nand U16539 (N_16539,N_11990,N_7423);
nand U16540 (N_16540,N_9119,N_7507);
or U16541 (N_16541,N_9985,N_6143);
xor U16542 (N_16542,N_10840,N_8015);
nand U16543 (N_16543,N_8413,N_11778);
or U16544 (N_16544,N_9552,N_6602);
or U16545 (N_16545,N_10742,N_6697);
and U16546 (N_16546,N_8372,N_8386);
xnor U16547 (N_16547,N_11080,N_8168);
xor U16548 (N_16548,N_11315,N_8253);
and U16549 (N_16549,N_9193,N_6017);
or U16550 (N_16550,N_6421,N_10873);
nand U16551 (N_16551,N_7856,N_6539);
nor U16552 (N_16552,N_8607,N_11743);
nor U16553 (N_16553,N_10946,N_9898);
xor U16554 (N_16554,N_9187,N_11063);
xnor U16555 (N_16555,N_6575,N_10599);
and U16556 (N_16556,N_6381,N_7852);
and U16557 (N_16557,N_11316,N_10112);
or U16558 (N_16558,N_8373,N_9742);
nand U16559 (N_16559,N_11204,N_6628);
nand U16560 (N_16560,N_8117,N_6236);
xnor U16561 (N_16561,N_6378,N_9894);
nand U16562 (N_16562,N_10281,N_6801);
nand U16563 (N_16563,N_6344,N_8341);
nor U16564 (N_16564,N_9623,N_8804);
nor U16565 (N_16565,N_9033,N_9319);
or U16566 (N_16566,N_6670,N_7145);
or U16567 (N_16567,N_11478,N_9567);
xor U16568 (N_16568,N_7127,N_6360);
nand U16569 (N_16569,N_7143,N_10294);
nand U16570 (N_16570,N_6035,N_7650);
nor U16571 (N_16571,N_7741,N_8071);
and U16572 (N_16572,N_10399,N_6989);
nor U16573 (N_16573,N_11198,N_8518);
and U16574 (N_16574,N_8771,N_8846);
nand U16575 (N_16575,N_7422,N_8667);
and U16576 (N_16576,N_11581,N_7508);
and U16577 (N_16577,N_8338,N_10848);
or U16578 (N_16578,N_7349,N_6851);
and U16579 (N_16579,N_9800,N_11743);
nor U16580 (N_16580,N_11090,N_9480);
xor U16581 (N_16581,N_7948,N_6394);
xor U16582 (N_16582,N_6974,N_9351);
nor U16583 (N_16583,N_11468,N_11295);
and U16584 (N_16584,N_7946,N_10270);
xor U16585 (N_16585,N_6998,N_9850);
and U16586 (N_16586,N_7945,N_9065);
nor U16587 (N_16587,N_6707,N_10197);
and U16588 (N_16588,N_6449,N_10813);
xor U16589 (N_16589,N_8713,N_11116);
and U16590 (N_16590,N_9827,N_7133);
nand U16591 (N_16591,N_7728,N_11918);
and U16592 (N_16592,N_11736,N_11518);
and U16593 (N_16593,N_6036,N_9753);
nand U16594 (N_16594,N_7280,N_10824);
nand U16595 (N_16595,N_9698,N_9638);
or U16596 (N_16596,N_10802,N_10300);
nor U16597 (N_16597,N_9682,N_11137);
nor U16598 (N_16598,N_6793,N_8092);
or U16599 (N_16599,N_6590,N_10310);
xnor U16600 (N_16600,N_11726,N_8915);
nor U16601 (N_16601,N_7039,N_9324);
or U16602 (N_16602,N_11540,N_8268);
xor U16603 (N_16603,N_9698,N_9198);
nand U16604 (N_16604,N_9914,N_10441);
xnor U16605 (N_16605,N_7071,N_8315);
nand U16606 (N_16606,N_9873,N_6496);
and U16607 (N_16607,N_6626,N_9870);
xnor U16608 (N_16608,N_10964,N_7166);
and U16609 (N_16609,N_9172,N_8947);
nand U16610 (N_16610,N_7073,N_11627);
or U16611 (N_16611,N_10981,N_6756);
nand U16612 (N_16612,N_7064,N_11920);
xnor U16613 (N_16613,N_8957,N_9756);
xor U16614 (N_16614,N_8338,N_11453);
and U16615 (N_16615,N_11675,N_7983);
nand U16616 (N_16616,N_7232,N_8798);
or U16617 (N_16617,N_6681,N_7830);
and U16618 (N_16618,N_6532,N_8332);
nand U16619 (N_16619,N_7197,N_7587);
nand U16620 (N_16620,N_6234,N_9791);
nor U16621 (N_16621,N_7281,N_9645);
and U16622 (N_16622,N_9215,N_11347);
or U16623 (N_16623,N_6686,N_8524);
or U16624 (N_16624,N_8679,N_6553);
xnor U16625 (N_16625,N_9588,N_9059);
nand U16626 (N_16626,N_8652,N_11008);
and U16627 (N_16627,N_6220,N_10235);
and U16628 (N_16628,N_11717,N_9257);
xor U16629 (N_16629,N_10550,N_10523);
nor U16630 (N_16630,N_8012,N_7142);
nand U16631 (N_16631,N_6546,N_11536);
or U16632 (N_16632,N_8717,N_7134);
xnor U16633 (N_16633,N_11296,N_9145);
or U16634 (N_16634,N_7998,N_7413);
xnor U16635 (N_16635,N_7091,N_7210);
nand U16636 (N_16636,N_8257,N_7902);
nor U16637 (N_16637,N_11721,N_9558);
xnor U16638 (N_16638,N_11783,N_8528);
and U16639 (N_16639,N_8399,N_10171);
xnor U16640 (N_16640,N_7085,N_10881);
xor U16641 (N_16641,N_9520,N_11917);
or U16642 (N_16642,N_7773,N_6670);
nor U16643 (N_16643,N_6032,N_10688);
nand U16644 (N_16644,N_6576,N_7083);
nor U16645 (N_16645,N_8176,N_10173);
nand U16646 (N_16646,N_7466,N_11475);
xor U16647 (N_16647,N_9985,N_11765);
nand U16648 (N_16648,N_9181,N_7037);
and U16649 (N_16649,N_10633,N_8040);
and U16650 (N_16650,N_8290,N_6145);
and U16651 (N_16651,N_8511,N_9272);
xnor U16652 (N_16652,N_8416,N_6035);
and U16653 (N_16653,N_8096,N_10998);
or U16654 (N_16654,N_8797,N_9859);
nand U16655 (N_16655,N_6936,N_10008);
nor U16656 (N_16656,N_6647,N_7422);
and U16657 (N_16657,N_6389,N_6484);
and U16658 (N_16658,N_9747,N_8514);
nand U16659 (N_16659,N_7385,N_10613);
and U16660 (N_16660,N_7335,N_7428);
nand U16661 (N_16661,N_11078,N_9780);
nand U16662 (N_16662,N_8617,N_11748);
nor U16663 (N_16663,N_10025,N_7085);
and U16664 (N_16664,N_6640,N_10642);
xnor U16665 (N_16665,N_10589,N_10418);
xnor U16666 (N_16666,N_11934,N_11145);
or U16667 (N_16667,N_10106,N_8154);
nor U16668 (N_16668,N_9589,N_8349);
nor U16669 (N_16669,N_8694,N_9152);
nor U16670 (N_16670,N_7984,N_7402);
xor U16671 (N_16671,N_9370,N_6610);
or U16672 (N_16672,N_8239,N_7458);
nor U16673 (N_16673,N_10543,N_11149);
nor U16674 (N_16674,N_7352,N_7225);
and U16675 (N_16675,N_6363,N_8779);
nand U16676 (N_16676,N_8840,N_6402);
and U16677 (N_16677,N_8425,N_11403);
and U16678 (N_16678,N_7487,N_8492);
nor U16679 (N_16679,N_9826,N_6451);
or U16680 (N_16680,N_9955,N_8533);
or U16681 (N_16681,N_7541,N_8563);
nor U16682 (N_16682,N_8080,N_8104);
and U16683 (N_16683,N_9723,N_8462);
xnor U16684 (N_16684,N_10912,N_6282);
nand U16685 (N_16685,N_8277,N_8321);
nor U16686 (N_16686,N_10083,N_10007);
nand U16687 (N_16687,N_7329,N_10204);
and U16688 (N_16688,N_6668,N_11554);
and U16689 (N_16689,N_8471,N_10254);
nor U16690 (N_16690,N_8117,N_6443);
and U16691 (N_16691,N_9276,N_6685);
nor U16692 (N_16692,N_11609,N_9526);
nor U16693 (N_16693,N_11797,N_11605);
nand U16694 (N_16694,N_10742,N_8347);
and U16695 (N_16695,N_10448,N_11674);
or U16696 (N_16696,N_10794,N_8279);
nand U16697 (N_16697,N_10837,N_7394);
or U16698 (N_16698,N_8489,N_7092);
nand U16699 (N_16699,N_10480,N_11498);
and U16700 (N_16700,N_6924,N_6034);
nand U16701 (N_16701,N_6586,N_9147);
or U16702 (N_16702,N_9377,N_8458);
xor U16703 (N_16703,N_7275,N_6656);
or U16704 (N_16704,N_9243,N_10809);
and U16705 (N_16705,N_8326,N_9864);
and U16706 (N_16706,N_11884,N_7773);
and U16707 (N_16707,N_6302,N_6864);
and U16708 (N_16708,N_6930,N_11445);
xor U16709 (N_16709,N_11991,N_10662);
nor U16710 (N_16710,N_10605,N_6494);
or U16711 (N_16711,N_7895,N_10030);
nor U16712 (N_16712,N_10288,N_6608);
nor U16713 (N_16713,N_11511,N_8192);
nor U16714 (N_16714,N_6490,N_10769);
and U16715 (N_16715,N_7834,N_9056);
nand U16716 (N_16716,N_11787,N_10487);
and U16717 (N_16717,N_8808,N_9897);
nand U16718 (N_16718,N_10041,N_6179);
or U16719 (N_16719,N_11480,N_9970);
nand U16720 (N_16720,N_9071,N_10277);
nor U16721 (N_16721,N_9909,N_6512);
or U16722 (N_16722,N_8912,N_8298);
and U16723 (N_16723,N_9999,N_6500);
nand U16724 (N_16724,N_6790,N_7713);
and U16725 (N_16725,N_6405,N_6509);
nor U16726 (N_16726,N_6430,N_8288);
nor U16727 (N_16727,N_9342,N_11350);
nand U16728 (N_16728,N_10878,N_6091);
xnor U16729 (N_16729,N_8058,N_8584);
or U16730 (N_16730,N_11349,N_7439);
nor U16731 (N_16731,N_8012,N_11431);
xor U16732 (N_16732,N_10299,N_11587);
nand U16733 (N_16733,N_7656,N_8612);
nand U16734 (N_16734,N_7381,N_8496);
and U16735 (N_16735,N_9816,N_7317);
and U16736 (N_16736,N_6223,N_10874);
nor U16737 (N_16737,N_8898,N_10361);
xor U16738 (N_16738,N_11622,N_11479);
and U16739 (N_16739,N_8262,N_10364);
nand U16740 (N_16740,N_7883,N_11458);
nand U16741 (N_16741,N_11735,N_6673);
or U16742 (N_16742,N_6353,N_11666);
nor U16743 (N_16743,N_9516,N_8971);
xnor U16744 (N_16744,N_10141,N_8878);
xnor U16745 (N_16745,N_10836,N_6570);
nand U16746 (N_16746,N_6356,N_6512);
nor U16747 (N_16747,N_8552,N_9744);
or U16748 (N_16748,N_6119,N_10060);
or U16749 (N_16749,N_11676,N_6081);
nand U16750 (N_16750,N_11331,N_6140);
and U16751 (N_16751,N_11983,N_11348);
nand U16752 (N_16752,N_8034,N_7690);
nand U16753 (N_16753,N_10018,N_6214);
nand U16754 (N_16754,N_8294,N_6802);
nor U16755 (N_16755,N_10235,N_7785);
and U16756 (N_16756,N_10441,N_10809);
or U16757 (N_16757,N_11244,N_8326);
and U16758 (N_16758,N_9317,N_7624);
nor U16759 (N_16759,N_9883,N_7805);
nor U16760 (N_16760,N_6619,N_6273);
and U16761 (N_16761,N_6655,N_7280);
or U16762 (N_16762,N_11006,N_10833);
nand U16763 (N_16763,N_7229,N_10073);
xor U16764 (N_16764,N_9372,N_6250);
xor U16765 (N_16765,N_11048,N_11677);
and U16766 (N_16766,N_7947,N_11449);
nand U16767 (N_16767,N_6147,N_9280);
nand U16768 (N_16768,N_10903,N_8890);
xnor U16769 (N_16769,N_6971,N_6878);
and U16770 (N_16770,N_9819,N_10430);
nor U16771 (N_16771,N_8515,N_9908);
nor U16772 (N_16772,N_11963,N_9673);
nand U16773 (N_16773,N_7425,N_8532);
or U16774 (N_16774,N_11050,N_10274);
nor U16775 (N_16775,N_9993,N_6541);
xor U16776 (N_16776,N_10440,N_9395);
nor U16777 (N_16777,N_6759,N_10136);
xor U16778 (N_16778,N_10257,N_9520);
nand U16779 (N_16779,N_6541,N_6081);
nand U16780 (N_16780,N_7836,N_9710);
and U16781 (N_16781,N_9551,N_11508);
xor U16782 (N_16782,N_6436,N_6750);
xor U16783 (N_16783,N_8637,N_7257);
nand U16784 (N_16784,N_6365,N_6191);
nand U16785 (N_16785,N_11778,N_9888);
and U16786 (N_16786,N_7081,N_7723);
and U16787 (N_16787,N_9113,N_6930);
or U16788 (N_16788,N_7494,N_11687);
xor U16789 (N_16789,N_6191,N_10156);
xnor U16790 (N_16790,N_11895,N_11354);
nand U16791 (N_16791,N_10485,N_8240);
xnor U16792 (N_16792,N_11963,N_10850);
and U16793 (N_16793,N_6489,N_10395);
nand U16794 (N_16794,N_8332,N_8467);
nand U16795 (N_16795,N_11193,N_10509);
nor U16796 (N_16796,N_9972,N_6335);
xnor U16797 (N_16797,N_6863,N_8425);
nor U16798 (N_16798,N_11357,N_11798);
and U16799 (N_16799,N_7610,N_10859);
and U16800 (N_16800,N_11085,N_10242);
nand U16801 (N_16801,N_11775,N_7657);
and U16802 (N_16802,N_6398,N_6555);
xnor U16803 (N_16803,N_7286,N_6956);
nand U16804 (N_16804,N_8146,N_7806);
and U16805 (N_16805,N_11420,N_9508);
and U16806 (N_16806,N_9290,N_7193);
nor U16807 (N_16807,N_6765,N_10347);
nor U16808 (N_16808,N_11998,N_6024);
and U16809 (N_16809,N_7893,N_6441);
or U16810 (N_16810,N_9631,N_9890);
or U16811 (N_16811,N_10714,N_9565);
or U16812 (N_16812,N_9500,N_7663);
nor U16813 (N_16813,N_9758,N_8393);
nor U16814 (N_16814,N_8257,N_6312);
xnor U16815 (N_16815,N_9145,N_7369);
nand U16816 (N_16816,N_9315,N_11282);
or U16817 (N_16817,N_6260,N_10317);
or U16818 (N_16818,N_11665,N_9170);
xnor U16819 (N_16819,N_9253,N_9773);
or U16820 (N_16820,N_8832,N_11594);
xor U16821 (N_16821,N_8721,N_6602);
or U16822 (N_16822,N_8214,N_8688);
nor U16823 (N_16823,N_6947,N_6712);
nand U16824 (N_16824,N_6122,N_10078);
xnor U16825 (N_16825,N_7924,N_6065);
nand U16826 (N_16826,N_7837,N_7554);
nor U16827 (N_16827,N_9376,N_6498);
and U16828 (N_16828,N_7041,N_9787);
and U16829 (N_16829,N_9437,N_11401);
nand U16830 (N_16830,N_10903,N_6214);
xnor U16831 (N_16831,N_6053,N_9102);
nor U16832 (N_16832,N_9090,N_9725);
nor U16833 (N_16833,N_6627,N_8649);
xnor U16834 (N_16834,N_8317,N_11181);
and U16835 (N_16835,N_7739,N_7064);
and U16836 (N_16836,N_9739,N_9967);
nand U16837 (N_16837,N_6839,N_6856);
xnor U16838 (N_16838,N_8227,N_8880);
nor U16839 (N_16839,N_10073,N_9921);
nand U16840 (N_16840,N_7067,N_11858);
nand U16841 (N_16841,N_8118,N_11591);
or U16842 (N_16842,N_8316,N_10089);
nand U16843 (N_16843,N_10258,N_6222);
xor U16844 (N_16844,N_8779,N_6589);
nand U16845 (N_16845,N_11803,N_6840);
xor U16846 (N_16846,N_9121,N_8050);
or U16847 (N_16847,N_7028,N_11148);
or U16848 (N_16848,N_6394,N_6511);
and U16849 (N_16849,N_6797,N_6774);
or U16850 (N_16850,N_11719,N_11347);
nand U16851 (N_16851,N_7837,N_7497);
nor U16852 (N_16852,N_10012,N_9837);
xnor U16853 (N_16853,N_9862,N_10805);
and U16854 (N_16854,N_9973,N_8051);
nor U16855 (N_16855,N_9726,N_8832);
nand U16856 (N_16856,N_11150,N_6717);
and U16857 (N_16857,N_8491,N_9312);
nor U16858 (N_16858,N_11247,N_7425);
nor U16859 (N_16859,N_7515,N_8803);
and U16860 (N_16860,N_11206,N_6445);
nand U16861 (N_16861,N_10854,N_6825);
and U16862 (N_16862,N_6843,N_11960);
xnor U16863 (N_16863,N_7116,N_7449);
nor U16864 (N_16864,N_8329,N_7614);
or U16865 (N_16865,N_8964,N_7525);
nand U16866 (N_16866,N_7530,N_10530);
nor U16867 (N_16867,N_6763,N_9661);
nor U16868 (N_16868,N_8381,N_6623);
xor U16869 (N_16869,N_6490,N_11097);
nand U16870 (N_16870,N_9047,N_9950);
and U16871 (N_16871,N_7734,N_8840);
xnor U16872 (N_16872,N_8836,N_6564);
or U16873 (N_16873,N_6216,N_6998);
and U16874 (N_16874,N_10761,N_8097);
and U16875 (N_16875,N_6389,N_6496);
or U16876 (N_16876,N_10872,N_11311);
nand U16877 (N_16877,N_10252,N_7142);
xor U16878 (N_16878,N_7018,N_8346);
xnor U16879 (N_16879,N_6545,N_8001);
nor U16880 (N_16880,N_11057,N_7273);
or U16881 (N_16881,N_11032,N_7281);
nand U16882 (N_16882,N_9422,N_7582);
nand U16883 (N_16883,N_11491,N_8298);
nor U16884 (N_16884,N_6278,N_10928);
nand U16885 (N_16885,N_11805,N_6808);
nor U16886 (N_16886,N_6981,N_6638);
nor U16887 (N_16887,N_10553,N_6049);
nand U16888 (N_16888,N_11253,N_9846);
and U16889 (N_16889,N_7311,N_11942);
and U16890 (N_16890,N_11346,N_6701);
nand U16891 (N_16891,N_9847,N_7884);
and U16892 (N_16892,N_8683,N_10052);
nor U16893 (N_16893,N_6997,N_10625);
and U16894 (N_16894,N_6085,N_10259);
nor U16895 (N_16895,N_8733,N_11765);
xnor U16896 (N_16896,N_11700,N_6398);
xnor U16897 (N_16897,N_10061,N_7048);
and U16898 (N_16898,N_11232,N_7440);
and U16899 (N_16899,N_9854,N_10636);
nand U16900 (N_16900,N_8950,N_10278);
and U16901 (N_16901,N_9555,N_6568);
and U16902 (N_16902,N_8947,N_10980);
xnor U16903 (N_16903,N_9351,N_9390);
or U16904 (N_16904,N_8019,N_10183);
or U16905 (N_16905,N_9583,N_10604);
nand U16906 (N_16906,N_10481,N_8311);
xor U16907 (N_16907,N_9025,N_6800);
nor U16908 (N_16908,N_6581,N_6392);
or U16909 (N_16909,N_9836,N_11448);
nor U16910 (N_16910,N_8376,N_7822);
nor U16911 (N_16911,N_11054,N_8666);
and U16912 (N_16912,N_10551,N_9070);
nor U16913 (N_16913,N_11021,N_11034);
xnor U16914 (N_16914,N_10000,N_10605);
nor U16915 (N_16915,N_7436,N_11290);
xnor U16916 (N_16916,N_11006,N_10265);
and U16917 (N_16917,N_7962,N_9421);
and U16918 (N_16918,N_7137,N_11374);
xnor U16919 (N_16919,N_6899,N_6293);
or U16920 (N_16920,N_9959,N_10608);
nor U16921 (N_16921,N_11279,N_10321);
and U16922 (N_16922,N_7227,N_11618);
nand U16923 (N_16923,N_8757,N_8190);
or U16924 (N_16924,N_7437,N_11355);
nand U16925 (N_16925,N_8898,N_7131);
xor U16926 (N_16926,N_10797,N_6486);
xnor U16927 (N_16927,N_11341,N_6280);
nor U16928 (N_16928,N_9104,N_11112);
or U16929 (N_16929,N_11038,N_11583);
or U16930 (N_16930,N_9181,N_10835);
or U16931 (N_16931,N_9065,N_9148);
or U16932 (N_16932,N_11003,N_8306);
xor U16933 (N_16933,N_6383,N_8992);
nand U16934 (N_16934,N_10179,N_10234);
or U16935 (N_16935,N_11927,N_8695);
nor U16936 (N_16936,N_7723,N_10087);
xor U16937 (N_16937,N_6704,N_10898);
and U16938 (N_16938,N_10724,N_9787);
nor U16939 (N_16939,N_8661,N_11678);
xnor U16940 (N_16940,N_7592,N_11867);
xor U16941 (N_16941,N_11826,N_9396);
nand U16942 (N_16942,N_6114,N_9460);
nor U16943 (N_16943,N_8146,N_8790);
and U16944 (N_16944,N_11667,N_8413);
nor U16945 (N_16945,N_11761,N_8222);
or U16946 (N_16946,N_8898,N_11690);
nand U16947 (N_16947,N_10368,N_9296);
nand U16948 (N_16948,N_11365,N_6503);
nor U16949 (N_16949,N_6497,N_7736);
xnor U16950 (N_16950,N_8388,N_10367);
nand U16951 (N_16951,N_10419,N_11524);
and U16952 (N_16952,N_6941,N_6238);
or U16953 (N_16953,N_9759,N_11602);
nand U16954 (N_16954,N_7876,N_6590);
nand U16955 (N_16955,N_10963,N_9338);
xor U16956 (N_16956,N_8892,N_8119);
nor U16957 (N_16957,N_8881,N_6641);
and U16958 (N_16958,N_6468,N_9439);
nand U16959 (N_16959,N_6141,N_9743);
nand U16960 (N_16960,N_11757,N_7483);
nor U16961 (N_16961,N_9159,N_8857);
nand U16962 (N_16962,N_10053,N_8083);
nand U16963 (N_16963,N_11391,N_11074);
xnor U16964 (N_16964,N_6158,N_7752);
xnor U16965 (N_16965,N_10770,N_8580);
and U16966 (N_16966,N_9407,N_6668);
xnor U16967 (N_16967,N_7344,N_8601);
nand U16968 (N_16968,N_10596,N_8413);
nor U16969 (N_16969,N_11111,N_7874);
xnor U16970 (N_16970,N_6793,N_11131);
nor U16971 (N_16971,N_6109,N_9045);
xor U16972 (N_16972,N_9142,N_11562);
or U16973 (N_16973,N_8076,N_9206);
nand U16974 (N_16974,N_8478,N_8867);
nor U16975 (N_16975,N_7774,N_6668);
and U16976 (N_16976,N_7163,N_7087);
nand U16977 (N_16977,N_9665,N_11732);
or U16978 (N_16978,N_6279,N_11068);
nor U16979 (N_16979,N_6665,N_9368);
or U16980 (N_16980,N_8378,N_8114);
or U16981 (N_16981,N_9667,N_11191);
or U16982 (N_16982,N_10723,N_8958);
nand U16983 (N_16983,N_11370,N_6596);
nand U16984 (N_16984,N_8459,N_9545);
and U16985 (N_16985,N_6758,N_11178);
nand U16986 (N_16986,N_9143,N_10928);
nand U16987 (N_16987,N_10288,N_6469);
nor U16988 (N_16988,N_10457,N_10630);
nor U16989 (N_16989,N_10077,N_9673);
and U16990 (N_16990,N_8548,N_9907);
and U16991 (N_16991,N_9869,N_11802);
or U16992 (N_16992,N_8125,N_6537);
and U16993 (N_16993,N_10277,N_8990);
or U16994 (N_16994,N_9772,N_10705);
nand U16995 (N_16995,N_6277,N_9802);
nor U16996 (N_16996,N_6997,N_10233);
xor U16997 (N_16997,N_11647,N_6273);
nand U16998 (N_16998,N_8308,N_9155);
xor U16999 (N_16999,N_9667,N_9857);
and U17000 (N_17000,N_11515,N_9488);
and U17001 (N_17001,N_6530,N_8469);
xnor U17002 (N_17002,N_11893,N_10740);
and U17003 (N_17003,N_11381,N_8229);
xnor U17004 (N_17004,N_8942,N_7076);
nor U17005 (N_17005,N_6427,N_10117);
or U17006 (N_17006,N_9356,N_6017);
xor U17007 (N_17007,N_8501,N_11018);
xor U17008 (N_17008,N_9272,N_10048);
and U17009 (N_17009,N_8386,N_8201);
xnor U17010 (N_17010,N_7747,N_6835);
nand U17011 (N_17011,N_11273,N_6457);
xor U17012 (N_17012,N_11144,N_7778);
xor U17013 (N_17013,N_6319,N_11168);
and U17014 (N_17014,N_10441,N_11361);
xor U17015 (N_17015,N_7838,N_6642);
xnor U17016 (N_17016,N_11773,N_9480);
or U17017 (N_17017,N_11106,N_10462);
nand U17018 (N_17018,N_6248,N_11191);
and U17019 (N_17019,N_6109,N_11313);
nor U17020 (N_17020,N_11802,N_11754);
nand U17021 (N_17021,N_9222,N_9395);
nand U17022 (N_17022,N_6454,N_6707);
xor U17023 (N_17023,N_6928,N_9668);
and U17024 (N_17024,N_11561,N_9654);
or U17025 (N_17025,N_10254,N_11525);
xnor U17026 (N_17026,N_10751,N_6207);
nor U17027 (N_17027,N_7345,N_6649);
or U17028 (N_17028,N_8889,N_8905);
xor U17029 (N_17029,N_10813,N_8279);
xnor U17030 (N_17030,N_8980,N_10981);
nor U17031 (N_17031,N_7077,N_6321);
or U17032 (N_17032,N_11074,N_8137);
or U17033 (N_17033,N_6896,N_7542);
nand U17034 (N_17034,N_8588,N_9275);
xor U17035 (N_17035,N_9810,N_11031);
xnor U17036 (N_17036,N_6812,N_8583);
or U17037 (N_17037,N_11474,N_9481);
nand U17038 (N_17038,N_10394,N_11065);
nor U17039 (N_17039,N_11845,N_7509);
or U17040 (N_17040,N_10195,N_8625);
nor U17041 (N_17041,N_11209,N_8655);
or U17042 (N_17042,N_11376,N_8898);
and U17043 (N_17043,N_8011,N_11894);
and U17044 (N_17044,N_7561,N_10059);
and U17045 (N_17045,N_9195,N_7874);
nor U17046 (N_17046,N_6965,N_9102);
or U17047 (N_17047,N_9352,N_7666);
nor U17048 (N_17048,N_9140,N_8105);
nand U17049 (N_17049,N_6865,N_8672);
or U17050 (N_17050,N_10801,N_9865);
nor U17051 (N_17051,N_10485,N_9983);
nor U17052 (N_17052,N_6870,N_9699);
and U17053 (N_17053,N_6225,N_8874);
nor U17054 (N_17054,N_10081,N_9221);
and U17055 (N_17055,N_9263,N_8738);
nand U17056 (N_17056,N_10273,N_6204);
nor U17057 (N_17057,N_7033,N_9871);
or U17058 (N_17058,N_11491,N_11449);
and U17059 (N_17059,N_7480,N_7898);
xnor U17060 (N_17060,N_7593,N_9873);
and U17061 (N_17061,N_8881,N_10935);
and U17062 (N_17062,N_10206,N_8817);
xnor U17063 (N_17063,N_8165,N_7207);
nand U17064 (N_17064,N_11876,N_9582);
and U17065 (N_17065,N_8352,N_11297);
and U17066 (N_17066,N_9176,N_7297);
and U17067 (N_17067,N_10810,N_6500);
xnor U17068 (N_17068,N_11916,N_7001);
xnor U17069 (N_17069,N_11576,N_8938);
nand U17070 (N_17070,N_10808,N_6322);
and U17071 (N_17071,N_7001,N_9048);
or U17072 (N_17072,N_9231,N_8216);
nand U17073 (N_17073,N_10903,N_6470);
and U17074 (N_17074,N_6521,N_6706);
nor U17075 (N_17075,N_6850,N_10663);
or U17076 (N_17076,N_6357,N_6928);
nand U17077 (N_17077,N_9815,N_8504);
nor U17078 (N_17078,N_8412,N_9305);
nor U17079 (N_17079,N_9768,N_11471);
and U17080 (N_17080,N_6773,N_9137);
xor U17081 (N_17081,N_11556,N_9359);
nand U17082 (N_17082,N_11763,N_11393);
nand U17083 (N_17083,N_7680,N_11011);
and U17084 (N_17084,N_9533,N_11511);
nand U17085 (N_17085,N_7055,N_10554);
and U17086 (N_17086,N_11674,N_6607);
or U17087 (N_17087,N_7703,N_11142);
nand U17088 (N_17088,N_7257,N_11154);
nor U17089 (N_17089,N_7088,N_9319);
or U17090 (N_17090,N_9262,N_10344);
or U17091 (N_17091,N_6739,N_6290);
and U17092 (N_17092,N_8020,N_6243);
xnor U17093 (N_17093,N_9985,N_8144);
nand U17094 (N_17094,N_9952,N_7116);
xor U17095 (N_17095,N_7898,N_7055);
nand U17096 (N_17096,N_10164,N_7296);
nor U17097 (N_17097,N_10259,N_11655);
and U17098 (N_17098,N_9274,N_8771);
nand U17099 (N_17099,N_9252,N_9908);
or U17100 (N_17100,N_7107,N_11755);
and U17101 (N_17101,N_10630,N_6520);
nand U17102 (N_17102,N_11709,N_7640);
nand U17103 (N_17103,N_9180,N_11252);
xor U17104 (N_17104,N_11523,N_7108);
and U17105 (N_17105,N_9640,N_8889);
or U17106 (N_17106,N_11049,N_7064);
nor U17107 (N_17107,N_6773,N_11120);
and U17108 (N_17108,N_7982,N_7483);
nand U17109 (N_17109,N_9999,N_6739);
and U17110 (N_17110,N_6816,N_9754);
xor U17111 (N_17111,N_6657,N_7546);
nor U17112 (N_17112,N_7130,N_9311);
or U17113 (N_17113,N_9497,N_8250);
nand U17114 (N_17114,N_11749,N_9323);
or U17115 (N_17115,N_10342,N_11707);
and U17116 (N_17116,N_6235,N_10574);
nand U17117 (N_17117,N_7304,N_9288);
nand U17118 (N_17118,N_9254,N_10958);
nand U17119 (N_17119,N_7940,N_8392);
nor U17120 (N_17120,N_7478,N_9446);
or U17121 (N_17121,N_8070,N_7115);
and U17122 (N_17122,N_8461,N_6531);
and U17123 (N_17123,N_8338,N_10765);
and U17124 (N_17124,N_10449,N_6614);
or U17125 (N_17125,N_11535,N_6154);
nor U17126 (N_17126,N_8340,N_9031);
and U17127 (N_17127,N_11589,N_10200);
nor U17128 (N_17128,N_8998,N_9272);
nand U17129 (N_17129,N_6102,N_6516);
and U17130 (N_17130,N_7209,N_7607);
xor U17131 (N_17131,N_8519,N_10540);
xnor U17132 (N_17132,N_6204,N_6975);
or U17133 (N_17133,N_11206,N_11398);
nor U17134 (N_17134,N_11782,N_7253);
nand U17135 (N_17135,N_11317,N_7989);
nand U17136 (N_17136,N_6603,N_7345);
nand U17137 (N_17137,N_10294,N_7604);
nor U17138 (N_17138,N_6157,N_6984);
or U17139 (N_17139,N_10507,N_10451);
and U17140 (N_17140,N_8791,N_10592);
xor U17141 (N_17141,N_9232,N_6505);
and U17142 (N_17142,N_6833,N_8202);
nor U17143 (N_17143,N_9076,N_11378);
nand U17144 (N_17144,N_11984,N_8792);
or U17145 (N_17145,N_11075,N_7410);
and U17146 (N_17146,N_7033,N_10752);
xor U17147 (N_17147,N_11505,N_10505);
nand U17148 (N_17148,N_11518,N_8040);
and U17149 (N_17149,N_10017,N_8772);
and U17150 (N_17150,N_11862,N_11863);
nor U17151 (N_17151,N_10988,N_9103);
and U17152 (N_17152,N_11042,N_11467);
xor U17153 (N_17153,N_10693,N_6116);
and U17154 (N_17154,N_10064,N_9330);
xnor U17155 (N_17155,N_7334,N_7360);
or U17156 (N_17156,N_9288,N_9559);
and U17157 (N_17157,N_11102,N_8751);
xnor U17158 (N_17158,N_10859,N_10249);
nand U17159 (N_17159,N_9215,N_10264);
nand U17160 (N_17160,N_7658,N_8353);
and U17161 (N_17161,N_7833,N_8077);
or U17162 (N_17162,N_10968,N_8993);
or U17163 (N_17163,N_8800,N_11883);
and U17164 (N_17164,N_8461,N_9911);
nor U17165 (N_17165,N_7768,N_11008);
nand U17166 (N_17166,N_6740,N_9626);
nor U17167 (N_17167,N_7207,N_11645);
xor U17168 (N_17168,N_6325,N_9137);
nand U17169 (N_17169,N_6358,N_8968);
nor U17170 (N_17170,N_8218,N_8541);
and U17171 (N_17171,N_6165,N_8508);
and U17172 (N_17172,N_8289,N_10419);
nand U17173 (N_17173,N_11486,N_11993);
and U17174 (N_17174,N_10462,N_8336);
nand U17175 (N_17175,N_9120,N_6198);
xor U17176 (N_17176,N_11435,N_9800);
and U17177 (N_17177,N_8829,N_6274);
nand U17178 (N_17178,N_11471,N_6509);
xnor U17179 (N_17179,N_8022,N_11785);
and U17180 (N_17180,N_11447,N_7211);
xor U17181 (N_17181,N_7258,N_9606);
or U17182 (N_17182,N_9610,N_9466);
or U17183 (N_17183,N_10028,N_11855);
nor U17184 (N_17184,N_7378,N_7260);
or U17185 (N_17185,N_7619,N_7665);
or U17186 (N_17186,N_10047,N_9878);
and U17187 (N_17187,N_11149,N_10132);
and U17188 (N_17188,N_11634,N_6429);
nand U17189 (N_17189,N_7129,N_7928);
or U17190 (N_17190,N_6223,N_8432);
xnor U17191 (N_17191,N_11589,N_7375);
nand U17192 (N_17192,N_9679,N_6903);
nand U17193 (N_17193,N_8535,N_6734);
nor U17194 (N_17194,N_10382,N_10136);
or U17195 (N_17195,N_9448,N_9806);
or U17196 (N_17196,N_9607,N_6768);
xnor U17197 (N_17197,N_10694,N_9668);
or U17198 (N_17198,N_11540,N_7165);
nor U17199 (N_17199,N_7129,N_7879);
xnor U17200 (N_17200,N_10219,N_6512);
xor U17201 (N_17201,N_10789,N_9831);
or U17202 (N_17202,N_11932,N_9151);
or U17203 (N_17203,N_10288,N_7056);
nand U17204 (N_17204,N_6774,N_8042);
and U17205 (N_17205,N_6086,N_8340);
xnor U17206 (N_17206,N_8326,N_6726);
xnor U17207 (N_17207,N_6024,N_8535);
xor U17208 (N_17208,N_10197,N_10877);
or U17209 (N_17209,N_10529,N_9622);
xnor U17210 (N_17210,N_6368,N_6197);
nor U17211 (N_17211,N_8892,N_9332);
nor U17212 (N_17212,N_7193,N_7345);
or U17213 (N_17213,N_11667,N_7614);
xor U17214 (N_17214,N_11650,N_11926);
nand U17215 (N_17215,N_11767,N_6531);
or U17216 (N_17216,N_8515,N_10815);
or U17217 (N_17217,N_7782,N_8795);
xor U17218 (N_17218,N_8568,N_10029);
or U17219 (N_17219,N_8170,N_7846);
xnor U17220 (N_17220,N_7811,N_11087);
or U17221 (N_17221,N_8278,N_8736);
or U17222 (N_17222,N_6282,N_10305);
or U17223 (N_17223,N_11551,N_11947);
or U17224 (N_17224,N_9423,N_10725);
xor U17225 (N_17225,N_6411,N_9658);
or U17226 (N_17226,N_11340,N_9466);
xor U17227 (N_17227,N_9025,N_11788);
nor U17228 (N_17228,N_9933,N_6680);
and U17229 (N_17229,N_10015,N_6277);
nor U17230 (N_17230,N_10014,N_9166);
and U17231 (N_17231,N_7374,N_9586);
nand U17232 (N_17232,N_6090,N_6349);
nand U17233 (N_17233,N_10664,N_11227);
xnor U17234 (N_17234,N_8437,N_7321);
xnor U17235 (N_17235,N_10532,N_11752);
nor U17236 (N_17236,N_9526,N_8194);
xnor U17237 (N_17237,N_7522,N_11739);
nand U17238 (N_17238,N_9347,N_11777);
xor U17239 (N_17239,N_10891,N_6116);
xor U17240 (N_17240,N_8127,N_11347);
nand U17241 (N_17241,N_9758,N_7687);
and U17242 (N_17242,N_10119,N_6673);
and U17243 (N_17243,N_6504,N_10087);
nand U17244 (N_17244,N_7724,N_10048);
nand U17245 (N_17245,N_10573,N_7723);
or U17246 (N_17246,N_9162,N_7080);
and U17247 (N_17247,N_10574,N_11566);
nor U17248 (N_17248,N_8429,N_7025);
nand U17249 (N_17249,N_9109,N_8481);
nor U17250 (N_17250,N_7082,N_7902);
or U17251 (N_17251,N_8582,N_8552);
and U17252 (N_17252,N_7613,N_6437);
and U17253 (N_17253,N_8706,N_10460);
or U17254 (N_17254,N_7313,N_6549);
xnor U17255 (N_17255,N_8725,N_7778);
xnor U17256 (N_17256,N_6465,N_8869);
xnor U17257 (N_17257,N_6741,N_7861);
or U17258 (N_17258,N_10665,N_9184);
nand U17259 (N_17259,N_9821,N_8800);
nand U17260 (N_17260,N_7267,N_8104);
nand U17261 (N_17261,N_6439,N_11349);
nand U17262 (N_17262,N_6807,N_7940);
xnor U17263 (N_17263,N_6739,N_6847);
and U17264 (N_17264,N_8591,N_7943);
xnor U17265 (N_17265,N_8989,N_11696);
xor U17266 (N_17266,N_6237,N_11127);
nand U17267 (N_17267,N_7354,N_8821);
and U17268 (N_17268,N_6968,N_9852);
or U17269 (N_17269,N_7002,N_10377);
or U17270 (N_17270,N_8318,N_10972);
nor U17271 (N_17271,N_11568,N_10864);
and U17272 (N_17272,N_7827,N_9033);
nand U17273 (N_17273,N_8001,N_8927);
nor U17274 (N_17274,N_8525,N_6709);
nand U17275 (N_17275,N_9247,N_6190);
and U17276 (N_17276,N_7775,N_7668);
xor U17277 (N_17277,N_10606,N_7532);
and U17278 (N_17278,N_8025,N_8930);
nand U17279 (N_17279,N_8016,N_7565);
xnor U17280 (N_17280,N_8393,N_11621);
nor U17281 (N_17281,N_9953,N_10529);
and U17282 (N_17282,N_7783,N_10064);
nand U17283 (N_17283,N_11470,N_10855);
nor U17284 (N_17284,N_9261,N_10018);
xnor U17285 (N_17285,N_10395,N_9734);
nor U17286 (N_17286,N_9596,N_6256);
nand U17287 (N_17287,N_8320,N_8336);
xnor U17288 (N_17288,N_7111,N_8733);
nor U17289 (N_17289,N_10645,N_7376);
and U17290 (N_17290,N_9212,N_10684);
nor U17291 (N_17291,N_7373,N_11720);
and U17292 (N_17292,N_7923,N_6286);
or U17293 (N_17293,N_9770,N_9547);
nor U17294 (N_17294,N_8497,N_6135);
and U17295 (N_17295,N_11645,N_7748);
nor U17296 (N_17296,N_11195,N_9148);
or U17297 (N_17297,N_9678,N_10110);
nand U17298 (N_17298,N_11477,N_8913);
nor U17299 (N_17299,N_11597,N_7439);
or U17300 (N_17300,N_8898,N_10797);
nand U17301 (N_17301,N_6188,N_8077);
or U17302 (N_17302,N_8531,N_6904);
nand U17303 (N_17303,N_11080,N_9447);
nand U17304 (N_17304,N_6259,N_10179);
nor U17305 (N_17305,N_9758,N_11316);
or U17306 (N_17306,N_8604,N_11334);
and U17307 (N_17307,N_10920,N_6818);
nand U17308 (N_17308,N_8678,N_8829);
or U17309 (N_17309,N_11085,N_7193);
or U17310 (N_17310,N_10577,N_11461);
or U17311 (N_17311,N_6184,N_11161);
nand U17312 (N_17312,N_11386,N_8915);
and U17313 (N_17313,N_10139,N_6394);
or U17314 (N_17314,N_11863,N_9388);
or U17315 (N_17315,N_10070,N_9138);
xnor U17316 (N_17316,N_11012,N_7841);
xnor U17317 (N_17317,N_11467,N_6381);
nand U17318 (N_17318,N_8094,N_8022);
nor U17319 (N_17319,N_9833,N_11765);
xnor U17320 (N_17320,N_9194,N_6842);
and U17321 (N_17321,N_9731,N_8880);
nor U17322 (N_17322,N_9806,N_6878);
xnor U17323 (N_17323,N_10310,N_10647);
and U17324 (N_17324,N_9713,N_6571);
and U17325 (N_17325,N_7557,N_8366);
and U17326 (N_17326,N_6761,N_7379);
xnor U17327 (N_17327,N_7564,N_7674);
xnor U17328 (N_17328,N_11724,N_9205);
or U17329 (N_17329,N_7417,N_11333);
and U17330 (N_17330,N_7026,N_10328);
xor U17331 (N_17331,N_7920,N_11188);
and U17332 (N_17332,N_11584,N_9540);
or U17333 (N_17333,N_8180,N_10336);
and U17334 (N_17334,N_8909,N_6619);
nor U17335 (N_17335,N_10698,N_9879);
or U17336 (N_17336,N_10377,N_9367);
nor U17337 (N_17337,N_7397,N_11942);
xor U17338 (N_17338,N_6680,N_8208);
nand U17339 (N_17339,N_9030,N_11451);
nand U17340 (N_17340,N_8627,N_9893);
and U17341 (N_17341,N_11890,N_9073);
and U17342 (N_17342,N_9781,N_8392);
or U17343 (N_17343,N_9413,N_10241);
or U17344 (N_17344,N_10271,N_10193);
nor U17345 (N_17345,N_8040,N_6549);
nor U17346 (N_17346,N_10834,N_6403);
or U17347 (N_17347,N_10365,N_10114);
or U17348 (N_17348,N_6773,N_7049);
nor U17349 (N_17349,N_7112,N_11463);
and U17350 (N_17350,N_8831,N_11986);
nand U17351 (N_17351,N_8878,N_10549);
nor U17352 (N_17352,N_7624,N_9125);
and U17353 (N_17353,N_9754,N_10245);
nor U17354 (N_17354,N_7659,N_9948);
and U17355 (N_17355,N_10603,N_7141);
xnor U17356 (N_17356,N_6377,N_11347);
and U17357 (N_17357,N_8357,N_8511);
and U17358 (N_17358,N_10919,N_11270);
nand U17359 (N_17359,N_8018,N_7789);
and U17360 (N_17360,N_8852,N_10276);
nand U17361 (N_17361,N_11040,N_8875);
nor U17362 (N_17362,N_8470,N_9976);
xnor U17363 (N_17363,N_11046,N_6055);
and U17364 (N_17364,N_8411,N_7454);
nand U17365 (N_17365,N_8236,N_8468);
xnor U17366 (N_17366,N_10582,N_10116);
nand U17367 (N_17367,N_8734,N_6722);
nor U17368 (N_17368,N_8000,N_11895);
nor U17369 (N_17369,N_10257,N_7449);
and U17370 (N_17370,N_10024,N_11335);
xnor U17371 (N_17371,N_11369,N_11380);
and U17372 (N_17372,N_7740,N_11063);
and U17373 (N_17373,N_6349,N_10146);
or U17374 (N_17374,N_10874,N_8950);
nor U17375 (N_17375,N_7940,N_11242);
nor U17376 (N_17376,N_6374,N_11640);
nand U17377 (N_17377,N_10761,N_7737);
nand U17378 (N_17378,N_7313,N_9828);
nor U17379 (N_17379,N_10073,N_9378);
and U17380 (N_17380,N_9543,N_8562);
nor U17381 (N_17381,N_11401,N_9265);
nand U17382 (N_17382,N_7540,N_8504);
xor U17383 (N_17383,N_7280,N_9699);
xor U17384 (N_17384,N_8251,N_11722);
or U17385 (N_17385,N_10781,N_8858);
nand U17386 (N_17386,N_8022,N_10477);
nor U17387 (N_17387,N_8717,N_6353);
or U17388 (N_17388,N_9850,N_9619);
and U17389 (N_17389,N_10570,N_9406);
or U17390 (N_17390,N_10162,N_6302);
xor U17391 (N_17391,N_8031,N_7133);
xnor U17392 (N_17392,N_8508,N_7023);
xnor U17393 (N_17393,N_9097,N_8917);
xor U17394 (N_17394,N_11302,N_8410);
nor U17395 (N_17395,N_10924,N_6640);
xor U17396 (N_17396,N_7315,N_9759);
nor U17397 (N_17397,N_11418,N_10419);
or U17398 (N_17398,N_9406,N_9246);
xnor U17399 (N_17399,N_6681,N_11008);
xor U17400 (N_17400,N_8920,N_10837);
nor U17401 (N_17401,N_7745,N_9515);
nor U17402 (N_17402,N_8476,N_10533);
nand U17403 (N_17403,N_8598,N_9170);
or U17404 (N_17404,N_11033,N_6559);
and U17405 (N_17405,N_11691,N_7789);
xnor U17406 (N_17406,N_11613,N_10714);
nand U17407 (N_17407,N_6179,N_8971);
and U17408 (N_17408,N_6343,N_9423);
xor U17409 (N_17409,N_9116,N_6416);
xnor U17410 (N_17410,N_10121,N_6942);
or U17411 (N_17411,N_9362,N_8412);
nand U17412 (N_17412,N_6031,N_7523);
nor U17413 (N_17413,N_10097,N_8312);
nand U17414 (N_17414,N_9426,N_11351);
nand U17415 (N_17415,N_6817,N_9895);
xnor U17416 (N_17416,N_8730,N_9943);
xor U17417 (N_17417,N_6094,N_7467);
xor U17418 (N_17418,N_10169,N_11618);
or U17419 (N_17419,N_7132,N_8541);
and U17420 (N_17420,N_11064,N_8695);
and U17421 (N_17421,N_8220,N_11759);
or U17422 (N_17422,N_11407,N_6414);
or U17423 (N_17423,N_7160,N_9391);
xor U17424 (N_17424,N_8708,N_10207);
xor U17425 (N_17425,N_8266,N_8589);
nor U17426 (N_17426,N_7415,N_11184);
and U17427 (N_17427,N_10948,N_8630);
nand U17428 (N_17428,N_6653,N_9250);
or U17429 (N_17429,N_10655,N_8817);
xor U17430 (N_17430,N_7839,N_9621);
nor U17431 (N_17431,N_7669,N_7779);
xnor U17432 (N_17432,N_10512,N_10710);
and U17433 (N_17433,N_11401,N_10137);
nand U17434 (N_17434,N_6193,N_9429);
or U17435 (N_17435,N_9392,N_9887);
nor U17436 (N_17436,N_9941,N_8494);
nor U17437 (N_17437,N_8554,N_10555);
nor U17438 (N_17438,N_6385,N_9356);
and U17439 (N_17439,N_10984,N_7775);
or U17440 (N_17440,N_7974,N_10364);
and U17441 (N_17441,N_6994,N_9986);
and U17442 (N_17442,N_6680,N_11089);
and U17443 (N_17443,N_6483,N_11064);
and U17444 (N_17444,N_8048,N_8667);
and U17445 (N_17445,N_11984,N_6245);
or U17446 (N_17446,N_11258,N_6143);
or U17447 (N_17447,N_8576,N_10843);
and U17448 (N_17448,N_9465,N_7608);
or U17449 (N_17449,N_7437,N_10291);
xnor U17450 (N_17450,N_9821,N_6362);
nor U17451 (N_17451,N_10574,N_8575);
or U17452 (N_17452,N_6268,N_6670);
xnor U17453 (N_17453,N_7274,N_7865);
xnor U17454 (N_17454,N_11506,N_9879);
or U17455 (N_17455,N_7934,N_6106);
xor U17456 (N_17456,N_9555,N_6056);
nand U17457 (N_17457,N_6357,N_7314);
nand U17458 (N_17458,N_10484,N_11861);
xor U17459 (N_17459,N_7691,N_6539);
nor U17460 (N_17460,N_10214,N_10124);
and U17461 (N_17461,N_9217,N_11627);
nor U17462 (N_17462,N_9617,N_7966);
and U17463 (N_17463,N_9885,N_11602);
nand U17464 (N_17464,N_7775,N_11444);
nor U17465 (N_17465,N_6264,N_11893);
xnor U17466 (N_17466,N_11213,N_6561);
and U17467 (N_17467,N_6107,N_11682);
nand U17468 (N_17468,N_7372,N_10367);
nor U17469 (N_17469,N_10768,N_7631);
nand U17470 (N_17470,N_9933,N_10227);
and U17471 (N_17471,N_6256,N_10827);
nor U17472 (N_17472,N_9994,N_8160);
or U17473 (N_17473,N_6699,N_8113);
and U17474 (N_17474,N_10495,N_9054);
and U17475 (N_17475,N_11296,N_8847);
or U17476 (N_17476,N_7423,N_9215);
or U17477 (N_17477,N_7761,N_11987);
nor U17478 (N_17478,N_11037,N_11260);
nand U17479 (N_17479,N_10814,N_7889);
or U17480 (N_17480,N_8053,N_10463);
or U17481 (N_17481,N_9827,N_11836);
or U17482 (N_17482,N_11478,N_8292);
or U17483 (N_17483,N_6819,N_8257);
nand U17484 (N_17484,N_6328,N_9631);
xor U17485 (N_17485,N_6956,N_8024);
nand U17486 (N_17486,N_11762,N_10366);
or U17487 (N_17487,N_10001,N_7026);
or U17488 (N_17488,N_8995,N_6904);
and U17489 (N_17489,N_11211,N_7770);
and U17490 (N_17490,N_6100,N_11047);
or U17491 (N_17491,N_6147,N_11163);
xnor U17492 (N_17492,N_6338,N_7174);
nand U17493 (N_17493,N_7338,N_8004);
xor U17494 (N_17494,N_8286,N_10856);
and U17495 (N_17495,N_11209,N_11503);
xnor U17496 (N_17496,N_7573,N_6209);
xnor U17497 (N_17497,N_10673,N_10026);
and U17498 (N_17498,N_10657,N_10575);
or U17499 (N_17499,N_8103,N_8069);
nand U17500 (N_17500,N_11023,N_7863);
nand U17501 (N_17501,N_6360,N_10801);
nor U17502 (N_17502,N_8822,N_7130);
nand U17503 (N_17503,N_10272,N_8097);
nor U17504 (N_17504,N_7721,N_7247);
nor U17505 (N_17505,N_9172,N_10484);
and U17506 (N_17506,N_10833,N_11920);
and U17507 (N_17507,N_10354,N_7324);
or U17508 (N_17508,N_7437,N_11930);
and U17509 (N_17509,N_9600,N_7687);
and U17510 (N_17510,N_10973,N_7151);
nand U17511 (N_17511,N_9882,N_8831);
nand U17512 (N_17512,N_10215,N_11638);
xnor U17513 (N_17513,N_8132,N_6432);
xor U17514 (N_17514,N_9246,N_8087);
or U17515 (N_17515,N_7854,N_7884);
or U17516 (N_17516,N_9512,N_7984);
xor U17517 (N_17517,N_6119,N_6444);
or U17518 (N_17518,N_8825,N_6848);
and U17519 (N_17519,N_11520,N_8992);
and U17520 (N_17520,N_9155,N_10800);
xnor U17521 (N_17521,N_10011,N_8109);
nor U17522 (N_17522,N_11063,N_7550);
nand U17523 (N_17523,N_8696,N_11235);
xor U17524 (N_17524,N_7276,N_8318);
and U17525 (N_17525,N_11280,N_11519);
nand U17526 (N_17526,N_11865,N_9544);
xnor U17527 (N_17527,N_6771,N_6192);
nor U17528 (N_17528,N_11281,N_8138);
or U17529 (N_17529,N_8016,N_8195);
nor U17530 (N_17530,N_8131,N_6376);
and U17531 (N_17531,N_11466,N_8036);
nand U17532 (N_17532,N_11244,N_6382);
nor U17533 (N_17533,N_9735,N_11707);
or U17534 (N_17534,N_7369,N_10390);
or U17535 (N_17535,N_11141,N_6188);
nor U17536 (N_17536,N_9939,N_10798);
nor U17537 (N_17537,N_6046,N_11411);
nor U17538 (N_17538,N_9995,N_9861);
or U17539 (N_17539,N_11950,N_7512);
nand U17540 (N_17540,N_6486,N_9715);
or U17541 (N_17541,N_9285,N_6555);
and U17542 (N_17542,N_7248,N_10141);
and U17543 (N_17543,N_7181,N_8317);
xor U17544 (N_17544,N_10378,N_7718);
nand U17545 (N_17545,N_11116,N_6908);
and U17546 (N_17546,N_10118,N_6710);
and U17547 (N_17547,N_8924,N_9757);
and U17548 (N_17548,N_6892,N_9819);
nor U17549 (N_17549,N_9920,N_8794);
and U17550 (N_17550,N_10504,N_11196);
and U17551 (N_17551,N_8298,N_10102);
nand U17552 (N_17552,N_8596,N_6769);
xnor U17553 (N_17553,N_6508,N_7728);
nand U17554 (N_17554,N_10882,N_6670);
or U17555 (N_17555,N_7087,N_11982);
or U17556 (N_17556,N_6882,N_8349);
or U17557 (N_17557,N_7978,N_9661);
nand U17558 (N_17558,N_7419,N_9996);
nor U17559 (N_17559,N_7325,N_11666);
and U17560 (N_17560,N_9849,N_7563);
xor U17561 (N_17561,N_10623,N_8238);
nor U17562 (N_17562,N_9857,N_10171);
nor U17563 (N_17563,N_7366,N_9376);
xnor U17564 (N_17564,N_7925,N_11437);
and U17565 (N_17565,N_10885,N_10267);
or U17566 (N_17566,N_8144,N_6648);
xor U17567 (N_17567,N_8228,N_8901);
nand U17568 (N_17568,N_8089,N_11380);
or U17569 (N_17569,N_10366,N_10664);
and U17570 (N_17570,N_9527,N_6697);
or U17571 (N_17571,N_6187,N_11546);
nor U17572 (N_17572,N_7166,N_10901);
nor U17573 (N_17573,N_8464,N_8872);
and U17574 (N_17574,N_8451,N_7020);
or U17575 (N_17575,N_6100,N_6364);
and U17576 (N_17576,N_8801,N_8032);
nor U17577 (N_17577,N_8054,N_7939);
xor U17578 (N_17578,N_8515,N_10128);
or U17579 (N_17579,N_6456,N_9723);
and U17580 (N_17580,N_6155,N_6126);
nor U17581 (N_17581,N_11292,N_11904);
xor U17582 (N_17582,N_7344,N_10555);
nor U17583 (N_17583,N_6940,N_6810);
nand U17584 (N_17584,N_10162,N_9567);
or U17585 (N_17585,N_11050,N_6954);
xnor U17586 (N_17586,N_9246,N_9142);
xor U17587 (N_17587,N_6015,N_8412);
nand U17588 (N_17588,N_11827,N_9916);
nand U17589 (N_17589,N_7815,N_7137);
or U17590 (N_17590,N_8788,N_8942);
xnor U17591 (N_17591,N_7025,N_9476);
nand U17592 (N_17592,N_6475,N_8612);
nor U17593 (N_17593,N_11713,N_11528);
and U17594 (N_17594,N_9965,N_8801);
and U17595 (N_17595,N_10081,N_10112);
xnor U17596 (N_17596,N_9319,N_11480);
nand U17597 (N_17597,N_9308,N_8168);
and U17598 (N_17598,N_8893,N_10107);
and U17599 (N_17599,N_6538,N_7694);
nor U17600 (N_17600,N_10006,N_10092);
and U17601 (N_17601,N_11542,N_6458);
and U17602 (N_17602,N_10179,N_9600);
xor U17603 (N_17603,N_8870,N_10713);
and U17604 (N_17604,N_10264,N_10375);
nor U17605 (N_17605,N_8045,N_6928);
and U17606 (N_17606,N_6973,N_11035);
nor U17607 (N_17607,N_9448,N_11562);
and U17608 (N_17608,N_9369,N_10700);
nor U17609 (N_17609,N_7023,N_8217);
and U17610 (N_17610,N_9865,N_10363);
nor U17611 (N_17611,N_8027,N_7920);
xor U17612 (N_17612,N_11275,N_8898);
nor U17613 (N_17613,N_11674,N_6138);
nand U17614 (N_17614,N_9193,N_9897);
and U17615 (N_17615,N_10724,N_9770);
and U17616 (N_17616,N_7172,N_10622);
xnor U17617 (N_17617,N_9843,N_7513);
and U17618 (N_17618,N_7559,N_11195);
and U17619 (N_17619,N_9308,N_10757);
nand U17620 (N_17620,N_6115,N_6866);
nand U17621 (N_17621,N_6705,N_8510);
nand U17622 (N_17622,N_9168,N_6705);
or U17623 (N_17623,N_7702,N_8321);
xnor U17624 (N_17624,N_7631,N_6883);
nor U17625 (N_17625,N_11733,N_7835);
nor U17626 (N_17626,N_10304,N_9450);
nor U17627 (N_17627,N_9831,N_11003);
nor U17628 (N_17628,N_8765,N_11252);
or U17629 (N_17629,N_6478,N_10651);
nor U17630 (N_17630,N_10391,N_8330);
xor U17631 (N_17631,N_9423,N_8216);
nor U17632 (N_17632,N_8926,N_7155);
or U17633 (N_17633,N_11453,N_7268);
xnor U17634 (N_17634,N_7602,N_8720);
nand U17635 (N_17635,N_11642,N_8608);
and U17636 (N_17636,N_7125,N_7594);
and U17637 (N_17637,N_8491,N_7665);
or U17638 (N_17638,N_6839,N_6263);
or U17639 (N_17639,N_6480,N_6047);
and U17640 (N_17640,N_10980,N_7265);
and U17641 (N_17641,N_7843,N_11285);
nand U17642 (N_17642,N_6819,N_9362);
nand U17643 (N_17643,N_8330,N_9727);
or U17644 (N_17644,N_7584,N_8574);
and U17645 (N_17645,N_10132,N_11717);
xor U17646 (N_17646,N_10255,N_10238);
and U17647 (N_17647,N_6111,N_8207);
or U17648 (N_17648,N_8357,N_7849);
or U17649 (N_17649,N_6818,N_10626);
or U17650 (N_17650,N_10765,N_9331);
nor U17651 (N_17651,N_6842,N_9819);
or U17652 (N_17652,N_7080,N_10303);
xnor U17653 (N_17653,N_8323,N_8596);
nand U17654 (N_17654,N_7850,N_10645);
nor U17655 (N_17655,N_11505,N_6601);
or U17656 (N_17656,N_8899,N_7916);
or U17657 (N_17657,N_9081,N_11068);
nand U17658 (N_17658,N_10034,N_10231);
and U17659 (N_17659,N_11188,N_7466);
or U17660 (N_17660,N_8037,N_10120);
nand U17661 (N_17661,N_9548,N_6176);
xnor U17662 (N_17662,N_10653,N_11916);
nor U17663 (N_17663,N_6921,N_10376);
nor U17664 (N_17664,N_9411,N_11524);
and U17665 (N_17665,N_7252,N_8859);
or U17666 (N_17666,N_6012,N_11811);
nand U17667 (N_17667,N_10271,N_11253);
or U17668 (N_17668,N_8744,N_7910);
nand U17669 (N_17669,N_7614,N_7904);
nand U17670 (N_17670,N_8008,N_8917);
xnor U17671 (N_17671,N_8237,N_7831);
nand U17672 (N_17672,N_7563,N_6735);
nand U17673 (N_17673,N_10082,N_7347);
xor U17674 (N_17674,N_11317,N_10423);
xnor U17675 (N_17675,N_6274,N_7007);
or U17676 (N_17676,N_6981,N_9570);
nor U17677 (N_17677,N_10466,N_10222);
nor U17678 (N_17678,N_11941,N_7396);
xor U17679 (N_17679,N_7814,N_11669);
xor U17680 (N_17680,N_10884,N_8343);
and U17681 (N_17681,N_6763,N_9762);
and U17682 (N_17682,N_10050,N_10917);
nand U17683 (N_17683,N_7008,N_6734);
and U17684 (N_17684,N_8685,N_8473);
or U17685 (N_17685,N_9744,N_11574);
nand U17686 (N_17686,N_9770,N_8714);
xnor U17687 (N_17687,N_10899,N_10053);
or U17688 (N_17688,N_7298,N_9609);
xnor U17689 (N_17689,N_6049,N_6016);
and U17690 (N_17690,N_7961,N_10088);
and U17691 (N_17691,N_10696,N_11056);
nand U17692 (N_17692,N_11144,N_10440);
nor U17693 (N_17693,N_7160,N_7213);
nand U17694 (N_17694,N_7545,N_10084);
xor U17695 (N_17695,N_9517,N_8945);
nor U17696 (N_17696,N_10931,N_7341);
nand U17697 (N_17697,N_6443,N_7448);
nand U17698 (N_17698,N_8986,N_6257);
nor U17699 (N_17699,N_6734,N_6044);
nor U17700 (N_17700,N_9600,N_7190);
nand U17701 (N_17701,N_11312,N_6917);
xor U17702 (N_17702,N_8915,N_7960);
nand U17703 (N_17703,N_11101,N_8896);
and U17704 (N_17704,N_8731,N_10935);
and U17705 (N_17705,N_10812,N_6709);
nand U17706 (N_17706,N_6400,N_6512);
and U17707 (N_17707,N_11404,N_10913);
xnor U17708 (N_17708,N_7542,N_7455);
xor U17709 (N_17709,N_7135,N_8011);
nor U17710 (N_17710,N_10615,N_7391);
nand U17711 (N_17711,N_9432,N_9603);
or U17712 (N_17712,N_6878,N_10714);
and U17713 (N_17713,N_10601,N_6511);
nor U17714 (N_17714,N_6678,N_8898);
nand U17715 (N_17715,N_8423,N_8154);
and U17716 (N_17716,N_8006,N_8369);
nand U17717 (N_17717,N_11408,N_9402);
nor U17718 (N_17718,N_7097,N_7742);
and U17719 (N_17719,N_6620,N_9172);
or U17720 (N_17720,N_8865,N_10548);
nor U17721 (N_17721,N_11193,N_8134);
nor U17722 (N_17722,N_8326,N_9671);
nor U17723 (N_17723,N_10750,N_9168);
xor U17724 (N_17724,N_10029,N_9999);
or U17725 (N_17725,N_10991,N_6566);
nor U17726 (N_17726,N_7568,N_6894);
or U17727 (N_17727,N_6180,N_9247);
or U17728 (N_17728,N_11145,N_11774);
and U17729 (N_17729,N_6227,N_6730);
xor U17730 (N_17730,N_10429,N_7860);
nand U17731 (N_17731,N_11402,N_10722);
or U17732 (N_17732,N_8418,N_11942);
nand U17733 (N_17733,N_11542,N_6728);
and U17734 (N_17734,N_6403,N_7502);
nand U17735 (N_17735,N_7635,N_10209);
nor U17736 (N_17736,N_7971,N_9519);
nor U17737 (N_17737,N_7404,N_6536);
nand U17738 (N_17738,N_7719,N_8518);
nor U17739 (N_17739,N_11697,N_7899);
or U17740 (N_17740,N_11770,N_8319);
nand U17741 (N_17741,N_6263,N_9842);
nand U17742 (N_17742,N_7459,N_7706);
xor U17743 (N_17743,N_10769,N_11150);
nand U17744 (N_17744,N_7228,N_9348);
nand U17745 (N_17745,N_10358,N_11937);
and U17746 (N_17746,N_11075,N_6344);
nand U17747 (N_17747,N_10985,N_8795);
xnor U17748 (N_17748,N_11665,N_7387);
nand U17749 (N_17749,N_10627,N_9941);
nand U17750 (N_17750,N_10983,N_7190);
or U17751 (N_17751,N_9900,N_6675);
xor U17752 (N_17752,N_11823,N_8827);
nand U17753 (N_17753,N_8497,N_9767);
nand U17754 (N_17754,N_9535,N_8147);
or U17755 (N_17755,N_6746,N_8994);
and U17756 (N_17756,N_6550,N_6615);
nor U17757 (N_17757,N_11275,N_8822);
and U17758 (N_17758,N_9858,N_9374);
or U17759 (N_17759,N_8500,N_6092);
and U17760 (N_17760,N_10672,N_10062);
nand U17761 (N_17761,N_6752,N_11225);
nor U17762 (N_17762,N_9736,N_11964);
or U17763 (N_17763,N_11113,N_6460);
or U17764 (N_17764,N_9671,N_7367);
nor U17765 (N_17765,N_11780,N_6016);
and U17766 (N_17766,N_7023,N_10024);
xor U17767 (N_17767,N_6657,N_10410);
nor U17768 (N_17768,N_9326,N_9451);
or U17769 (N_17769,N_8970,N_8585);
nand U17770 (N_17770,N_8644,N_8933);
xnor U17771 (N_17771,N_6967,N_6989);
xor U17772 (N_17772,N_6631,N_7818);
nor U17773 (N_17773,N_9300,N_9167);
and U17774 (N_17774,N_6149,N_11768);
nand U17775 (N_17775,N_6199,N_8257);
nor U17776 (N_17776,N_9225,N_7451);
xnor U17777 (N_17777,N_11849,N_10969);
or U17778 (N_17778,N_8159,N_11634);
xor U17779 (N_17779,N_11603,N_9907);
and U17780 (N_17780,N_9634,N_11679);
nand U17781 (N_17781,N_9870,N_6792);
or U17782 (N_17782,N_8809,N_10411);
nand U17783 (N_17783,N_10486,N_9507);
and U17784 (N_17784,N_8219,N_11129);
and U17785 (N_17785,N_6264,N_6585);
xnor U17786 (N_17786,N_6529,N_6395);
nand U17787 (N_17787,N_7749,N_11620);
and U17788 (N_17788,N_6044,N_11178);
nand U17789 (N_17789,N_6033,N_6216);
xor U17790 (N_17790,N_11676,N_10564);
xor U17791 (N_17791,N_10286,N_10016);
or U17792 (N_17792,N_7330,N_7530);
nor U17793 (N_17793,N_6163,N_9683);
or U17794 (N_17794,N_7358,N_7151);
and U17795 (N_17795,N_7610,N_9423);
xnor U17796 (N_17796,N_9987,N_9594);
xor U17797 (N_17797,N_10343,N_9336);
or U17798 (N_17798,N_9564,N_9048);
and U17799 (N_17799,N_7031,N_10974);
and U17800 (N_17800,N_9867,N_8222);
or U17801 (N_17801,N_7783,N_9585);
or U17802 (N_17802,N_8961,N_9931);
and U17803 (N_17803,N_9804,N_9042);
xor U17804 (N_17804,N_11772,N_9452);
xor U17805 (N_17805,N_7635,N_6917);
nor U17806 (N_17806,N_11955,N_6599);
nand U17807 (N_17807,N_7379,N_7102);
nor U17808 (N_17808,N_7796,N_8095);
nand U17809 (N_17809,N_7907,N_7792);
and U17810 (N_17810,N_10360,N_9050);
nor U17811 (N_17811,N_11278,N_7947);
nor U17812 (N_17812,N_10350,N_11403);
nand U17813 (N_17813,N_10698,N_10758);
or U17814 (N_17814,N_7052,N_8802);
or U17815 (N_17815,N_11403,N_10451);
or U17816 (N_17816,N_11077,N_6999);
or U17817 (N_17817,N_10244,N_10039);
xor U17818 (N_17818,N_6063,N_9999);
nor U17819 (N_17819,N_7208,N_8314);
and U17820 (N_17820,N_7879,N_10633);
nor U17821 (N_17821,N_8630,N_11828);
nor U17822 (N_17822,N_9297,N_7913);
or U17823 (N_17823,N_8211,N_7479);
xor U17824 (N_17824,N_11990,N_11617);
nor U17825 (N_17825,N_6340,N_10775);
xor U17826 (N_17826,N_8623,N_7374);
and U17827 (N_17827,N_10642,N_7730);
xnor U17828 (N_17828,N_9642,N_6951);
and U17829 (N_17829,N_11305,N_8943);
and U17830 (N_17830,N_9870,N_11261);
xor U17831 (N_17831,N_8806,N_8918);
or U17832 (N_17832,N_10736,N_6500);
and U17833 (N_17833,N_7049,N_8290);
xor U17834 (N_17834,N_7475,N_10185);
xnor U17835 (N_17835,N_10700,N_10640);
xor U17836 (N_17836,N_8507,N_10682);
nand U17837 (N_17837,N_9154,N_8008);
xor U17838 (N_17838,N_9470,N_11333);
and U17839 (N_17839,N_6178,N_6023);
nor U17840 (N_17840,N_8039,N_9380);
nor U17841 (N_17841,N_10349,N_9432);
and U17842 (N_17842,N_10248,N_8236);
nand U17843 (N_17843,N_6193,N_10422);
and U17844 (N_17844,N_7618,N_9852);
or U17845 (N_17845,N_7005,N_8514);
and U17846 (N_17846,N_11846,N_11308);
nand U17847 (N_17847,N_7904,N_7396);
or U17848 (N_17848,N_11638,N_8637);
xor U17849 (N_17849,N_9661,N_6777);
nor U17850 (N_17850,N_10543,N_10126);
nor U17851 (N_17851,N_10225,N_10091);
nor U17852 (N_17852,N_9693,N_10872);
xor U17853 (N_17853,N_6599,N_7089);
nor U17854 (N_17854,N_7824,N_6607);
and U17855 (N_17855,N_8607,N_8259);
and U17856 (N_17856,N_8286,N_11416);
or U17857 (N_17857,N_7540,N_11833);
and U17858 (N_17858,N_6836,N_11654);
nand U17859 (N_17859,N_11125,N_10887);
and U17860 (N_17860,N_7184,N_7685);
xor U17861 (N_17861,N_7193,N_10047);
or U17862 (N_17862,N_8403,N_11403);
and U17863 (N_17863,N_10357,N_6562);
and U17864 (N_17864,N_8342,N_7135);
and U17865 (N_17865,N_9505,N_8087);
nor U17866 (N_17866,N_7929,N_8639);
nand U17867 (N_17867,N_7979,N_11280);
xnor U17868 (N_17868,N_11716,N_9559);
or U17869 (N_17869,N_7247,N_9085);
nand U17870 (N_17870,N_9136,N_7475);
xor U17871 (N_17871,N_7821,N_7773);
and U17872 (N_17872,N_9521,N_9648);
or U17873 (N_17873,N_6548,N_9247);
and U17874 (N_17874,N_9571,N_6756);
nand U17875 (N_17875,N_8515,N_7122);
xnor U17876 (N_17876,N_8514,N_10732);
nor U17877 (N_17877,N_10935,N_9621);
xnor U17878 (N_17878,N_11178,N_10891);
nand U17879 (N_17879,N_6378,N_9930);
xnor U17880 (N_17880,N_11730,N_8052);
or U17881 (N_17881,N_10089,N_10291);
and U17882 (N_17882,N_9391,N_9375);
nor U17883 (N_17883,N_10207,N_9204);
nor U17884 (N_17884,N_11944,N_10438);
nand U17885 (N_17885,N_11288,N_11329);
or U17886 (N_17886,N_9590,N_7838);
or U17887 (N_17887,N_9062,N_9930);
nand U17888 (N_17888,N_11289,N_10182);
or U17889 (N_17889,N_9393,N_10999);
and U17890 (N_17890,N_6602,N_8174);
xor U17891 (N_17891,N_7527,N_7350);
nand U17892 (N_17892,N_10361,N_10153);
xor U17893 (N_17893,N_6835,N_7141);
or U17894 (N_17894,N_8786,N_10302);
nand U17895 (N_17895,N_11029,N_7169);
or U17896 (N_17896,N_10323,N_6539);
and U17897 (N_17897,N_8287,N_11193);
or U17898 (N_17898,N_11820,N_10764);
nor U17899 (N_17899,N_7788,N_7154);
xor U17900 (N_17900,N_7749,N_6857);
and U17901 (N_17901,N_11807,N_11325);
nor U17902 (N_17902,N_11563,N_10448);
or U17903 (N_17903,N_9814,N_9429);
nand U17904 (N_17904,N_8745,N_8903);
nand U17905 (N_17905,N_6949,N_8240);
and U17906 (N_17906,N_9512,N_6306);
or U17907 (N_17907,N_11674,N_9454);
or U17908 (N_17908,N_10080,N_8095);
and U17909 (N_17909,N_7133,N_7507);
and U17910 (N_17910,N_11830,N_9794);
nor U17911 (N_17911,N_6300,N_7805);
nor U17912 (N_17912,N_11998,N_11222);
or U17913 (N_17913,N_9632,N_9241);
xor U17914 (N_17914,N_10966,N_11116);
nor U17915 (N_17915,N_8085,N_7948);
nand U17916 (N_17916,N_8460,N_7879);
nand U17917 (N_17917,N_6689,N_10105);
nor U17918 (N_17918,N_11695,N_6335);
nor U17919 (N_17919,N_6682,N_7154);
and U17920 (N_17920,N_9507,N_6374);
or U17921 (N_17921,N_11325,N_11522);
xor U17922 (N_17922,N_8949,N_8397);
nand U17923 (N_17923,N_6118,N_9710);
and U17924 (N_17924,N_6462,N_6458);
nand U17925 (N_17925,N_10253,N_9918);
nand U17926 (N_17926,N_11502,N_10902);
xnor U17927 (N_17927,N_9315,N_6489);
nor U17928 (N_17928,N_6601,N_7474);
nor U17929 (N_17929,N_6819,N_9999);
xnor U17930 (N_17930,N_10444,N_10174);
or U17931 (N_17931,N_8400,N_6639);
nand U17932 (N_17932,N_7230,N_11725);
and U17933 (N_17933,N_7505,N_11723);
and U17934 (N_17934,N_11180,N_6301);
nand U17935 (N_17935,N_11801,N_6834);
nor U17936 (N_17936,N_8124,N_9511);
or U17937 (N_17937,N_10488,N_7802);
xor U17938 (N_17938,N_8605,N_7482);
or U17939 (N_17939,N_8136,N_11128);
nor U17940 (N_17940,N_7780,N_7168);
xor U17941 (N_17941,N_8769,N_11019);
or U17942 (N_17942,N_10508,N_6344);
or U17943 (N_17943,N_9115,N_9075);
nor U17944 (N_17944,N_9853,N_10617);
or U17945 (N_17945,N_6121,N_7576);
xor U17946 (N_17946,N_10904,N_9199);
and U17947 (N_17947,N_9064,N_8800);
nand U17948 (N_17948,N_6080,N_8012);
nor U17949 (N_17949,N_8767,N_7491);
nand U17950 (N_17950,N_9610,N_8520);
nand U17951 (N_17951,N_8643,N_8360);
xor U17952 (N_17952,N_11800,N_11904);
nor U17953 (N_17953,N_9714,N_8670);
nand U17954 (N_17954,N_8782,N_11734);
and U17955 (N_17955,N_6205,N_9109);
nand U17956 (N_17956,N_7499,N_9506);
nor U17957 (N_17957,N_7423,N_7015);
and U17958 (N_17958,N_6592,N_7636);
nand U17959 (N_17959,N_7000,N_11122);
xnor U17960 (N_17960,N_6582,N_7023);
and U17961 (N_17961,N_8574,N_8086);
or U17962 (N_17962,N_7892,N_6494);
xor U17963 (N_17963,N_8694,N_7742);
or U17964 (N_17964,N_11815,N_7822);
nand U17965 (N_17965,N_8817,N_10114);
xnor U17966 (N_17966,N_8610,N_8658);
nor U17967 (N_17967,N_11076,N_7630);
xnor U17968 (N_17968,N_10457,N_7592);
nand U17969 (N_17969,N_8601,N_10642);
nor U17970 (N_17970,N_9329,N_10052);
nor U17971 (N_17971,N_10646,N_7008);
nor U17972 (N_17972,N_11465,N_11750);
nand U17973 (N_17973,N_10419,N_8504);
xor U17974 (N_17974,N_10525,N_9149);
and U17975 (N_17975,N_6091,N_11762);
or U17976 (N_17976,N_7758,N_8861);
nor U17977 (N_17977,N_10564,N_10697);
or U17978 (N_17978,N_7891,N_8720);
or U17979 (N_17979,N_6825,N_8592);
xnor U17980 (N_17980,N_11025,N_9341);
nand U17981 (N_17981,N_10704,N_8568);
nand U17982 (N_17982,N_11903,N_11151);
or U17983 (N_17983,N_7980,N_10407);
nand U17984 (N_17984,N_11147,N_9485);
xor U17985 (N_17985,N_8364,N_11691);
nor U17986 (N_17986,N_11856,N_6018);
nand U17987 (N_17987,N_10854,N_8356);
or U17988 (N_17988,N_9188,N_9226);
nor U17989 (N_17989,N_11481,N_11801);
nor U17990 (N_17990,N_6776,N_11819);
and U17991 (N_17991,N_6162,N_9152);
nand U17992 (N_17992,N_9968,N_7873);
nand U17993 (N_17993,N_7862,N_11249);
nand U17994 (N_17994,N_8060,N_7569);
and U17995 (N_17995,N_6688,N_7842);
xor U17996 (N_17996,N_10334,N_11843);
nor U17997 (N_17997,N_10502,N_6963);
nand U17998 (N_17998,N_8505,N_7759);
xor U17999 (N_17999,N_10787,N_9341);
xnor U18000 (N_18000,N_15329,N_12020);
xor U18001 (N_18001,N_16540,N_12721);
nor U18002 (N_18002,N_12654,N_13237);
xor U18003 (N_18003,N_13482,N_14581);
nand U18004 (N_18004,N_12480,N_13557);
or U18005 (N_18005,N_12334,N_16419);
xor U18006 (N_18006,N_17597,N_13930);
or U18007 (N_18007,N_14478,N_15318);
nor U18008 (N_18008,N_13585,N_16581);
or U18009 (N_18009,N_17767,N_17157);
or U18010 (N_18010,N_15139,N_15458);
nand U18011 (N_18011,N_14976,N_17579);
or U18012 (N_18012,N_13380,N_12813);
nand U18013 (N_18013,N_15400,N_17081);
nor U18014 (N_18014,N_12143,N_12380);
or U18015 (N_18015,N_13906,N_17771);
and U18016 (N_18016,N_17168,N_15200);
and U18017 (N_18017,N_12984,N_16049);
xnor U18018 (N_18018,N_15846,N_15390);
xor U18019 (N_18019,N_16727,N_17970);
or U18020 (N_18020,N_14786,N_12521);
nor U18021 (N_18021,N_12478,N_12118);
nand U18022 (N_18022,N_15960,N_17919);
and U18023 (N_18023,N_17093,N_13866);
and U18024 (N_18024,N_12648,N_16552);
and U18025 (N_18025,N_17339,N_17867);
xnor U18026 (N_18026,N_17050,N_12421);
nor U18027 (N_18027,N_16123,N_13497);
xor U18028 (N_18028,N_15504,N_17089);
xnor U18029 (N_18029,N_17301,N_13843);
or U18030 (N_18030,N_12616,N_13057);
and U18031 (N_18031,N_17054,N_14963);
or U18032 (N_18032,N_15288,N_15822);
or U18033 (N_18033,N_17197,N_12790);
nor U18034 (N_18034,N_16221,N_16172);
nor U18035 (N_18035,N_14547,N_14638);
nor U18036 (N_18036,N_13871,N_13261);
and U18037 (N_18037,N_12829,N_14022);
or U18038 (N_18038,N_15793,N_17030);
and U18039 (N_18039,N_16779,N_13978);
nand U18040 (N_18040,N_16020,N_13891);
xor U18041 (N_18041,N_12361,N_12882);
and U18042 (N_18042,N_13727,N_16306);
or U18043 (N_18043,N_14929,N_17956);
nor U18044 (N_18044,N_12774,N_13718);
xor U18045 (N_18045,N_15298,N_14082);
xnor U18046 (N_18046,N_17260,N_15280);
or U18047 (N_18047,N_14999,N_12915);
xor U18048 (N_18048,N_13505,N_17110);
xor U18049 (N_18049,N_14118,N_15014);
or U18050 (N_18050,N_12910,N_14117);
and U18051 (N_18051,N_12195,N_17566);
and U18052 (N_18052,N_12538,N_15007);
and U18053 (N_18053,N_14243,N_15627);
and U18054 (N_18054,N_17856,N_16802);
nand U18055 (N_18055,N_14564,N_15522);
or U18056 (N_18056,N_13244,N_14842);
and U18057 (N_18057,N_15872,N_16403);
nand U18058 (N_18058,N_13699,N_14385);
and U18059 (N_18059,N_14126,N_12893);
and U18060 (N_18060,N_15763,N_15454);
nor U18061 (N_18061,N_17673,N_14709);
xnor U18062 (N_18062,N_13946,N_16447);
or U18063 (N_18063,N_16492,N_13535);
nor U18064 (N_18064,N_12506,N_13013);
nand U18065 (N_18065,N_14031,N_16255);
xor U18066 (N_18066,N_12233,N_13043);
or U18067 (N_18067,N_12043,N_13001);
and U18068 (N_18068,N_13007,N_14701);
nand U18069 (N_18069,N_16128,N_16658);
nand U18070 (N_18070,N_15203,N_12198);
nand U18071 (N_18071,N_17154,N_13822);
nand U18072 (N_18072,N_15144,N_17291);
and U18073 (N_18073,N_15398,N_12185);
nor U18074 (N_18074,N_12901,N_15302);
nand U18075 (N_18075,N_14891,N_13446);
nand U18076 (N_18076,N_12962,N_12932);
or U18077 (N_18077,N_13778,N_13426);
nand U18078 (N_18078,N_17368,N_14358);
and U18079 (N_18079,N_15669,N_17978);
xor U18080 (N_18080,N_12812,N_15017);
xor U18081 (N_18081,N_17506,N_13500);
nor U18082 (N_18082,N_12465,N_13274);
xor U18083 (N_18083,N_17290,N_17418);
nand U18084 (N_18084,N_13227,N_12713);
nand U18085 (N_18085,N_12898,N_14053);
xor U18086 (N_18086,N_14503,N_12035);
or U18087 (N_18087,N_17721,N_17865);
and U18088 (N_18088,N_13732,N_14067);
and U18089 (N_18089,N_13677,N_14710);
xnor U18090 (N_18090,N_15141,N_16914);
nand U18091 (N_18091,N_16074,N_12922);
and U18092 (N_18092,N_17058,N_15730);
or U18093 (N_18093,N_13472,N_13966);
nand U18094 (N_18094,N_15900,N_16973);
and U18095 (N_18095,N_13079,N_14696);
and U18096 (N_18096,N_14860,N_12665);
or U18097 (N_18097,N_13422,N_15577);
nand U18098 (N_18098,N_14239,N_12571);
and U18099 (N_18099,N_13743,N_16901);
and U18100 (N_18100,N_17468,N_13507);
or U18101 (N_18101,N_13076,N_17790);
xnor U18102 (N_18102,N_16240,N_16896);
nand U18103 (N_18103,N_15852,N_14937);
and U18104 (N_18104,N_17554,N_16147);
or U18105 (N_18105,N_12947,N_15119);
xor U18106 (N_18106,N_12096,N_12306);
or U18107 (N_18107,N_16398,N_12941);
xnor U18108 (N_18108,N_13471,N_14602);
or U18109 (N_18109,N_17769,N_12766);
or U18110 (N_18110,N_15500,N_17213);
xnor U18111 (N_18111,N_12823,N_13265);
and U18112 (N_18112,N_14674,N_17041);
xor U18113 (N_18113,N_13243,N_12447);
xnor U18114 (N_18114,N_13335,N_13002);
or U18115 (N_18115,N_13772,N_13492);
nor U18116 (N_18116,N_16558,N_14331);
or U18117 (N_18117,N_15999,N_17442);
nand U18118 (N_18118,N_15523,N_13728);
nor U18119 (N_18119,N_15132,N_17890);
nor U18120 (N_18120,N_15131,N_16620);
xnor U18121 (N_18121,N_12073,N_15216);
and U18122 (N_18122,N_17845,N_14107);
nand U18123 (N_18123,N_15968,N_12754);
nand U18124 (N_18124,N_13617,N_13150);
or U18125 (N_18125,N_17766,N_17895);
and U18126 (N_18126,N_17859,N_17492);
nor U18127 (N_18127,N_17539,N_17922);
or U18128 (N_18128,N_12290,N_15875);
xnor U18129 (N_18129,N_16728,N_16676);
xnor U18130 (N_18130,N_16585,N_16905);
nor U18131 (N_18131,N_13347,N_16757);
or U18132 (N_18132,N_15713,N_16265);
nor U18133 (N_18133,N_17355,N_14689);
xnor U18134 (N_18134,N_13986,N_14938);
or U18135 (N_18135,N_15210,N_15902);
nand U18136 (N_18136,N_16180,N_15704);
and U18137 (N_18137,N_15898,N_15981);
nor U18138 (N_18138,N_13449,N_16774);
nand U18139 (N_18139,N_15987,N_16030);
xnor U18140 (N_18140,N_15939,N_16890);
or U18141 (N_18141,N_14227,N_13551);
or U18142 (N_18142,N_17312,N_17774);
xor U18143 (N_18143,N_14327,N_17651);
nand U18144 (N_18144,N_12113,N_16379);
nand U18145 (N_18145,N_17403,N_15374);
nand U18146 (N_18146,N_12404,N_14723);
xor U18147 (N_18147,N_15440,N_17551);
xor U18148 (N_18148,N_13631,N_14868);
and U18149 (N_18149,N_16281,N_17122);
and U18150 (N_18150,N_15663,N_12800);
or U18151 (N_18151,N_12623,N_16959);
nand U18152 (N_18152,N_15516,N_16232);
and U18153 (N_18153,N_13559,N_16010);
and U18154 (N_18154,N_15641,N_14761);
nor U18155 (N_18155,N_13663,N_16640);
nor U18156 (N_18156,N_14182,N_17155);
and U18157 (N_18157,N_16149,N_12379);
nand U18158 (N_18158,N_16308,N_17594);
and U18159 (N_18159,N_14014,N_15287);
nand U18160 (N_18160,N_16148,N_16073);
nor U18161 (N_18161,N_13339,N_14017);
nand U18162 (N_18162,N_15559,N_12843);
or U18163 (N_18163,N_14647,N_17520);
nor U18164 (N_18164,N_12191,N_14831);
or U18165 (N_18165,N_15346,N_14065);
nor U18166 (N_18166,N_15137,N_13836);
xnor U18167 (N_18167,N_14936,N_15316);
and U18168 (N_18168,N_14718,N_12117);
and U18169 (N_18169,N_13488,N_17798);
nor U18170 (N_18170,N_17920,N_14822);
or U18171 (N_18171,N_12865,N_12111);
nor U18172 (N_18172,N_13165,N_15451);
or U18173 (N_18173,N_12406,N_14977);
nor U18174 (N_18174,N_16314,N_15493);
and U18175 (N_18175,N_14998,N_14747);
nand U18176 (N_18176,N_13712,N_16819);
and U18177 (N_18177,N_13287,N_14524);
and U18178 (N_18178,N_15134,N_12219);
xnor U18179 (N_18179,N_13795,N_16223);
and U18180 (N_18180,N_14857,N_15776);
nand U18181 (N_18181,N_12493,N_17815);
and U18182 (N_18182,N_15407,N_15575);
nand U18183 (N_18183,N_14802,N_15979);
nand U18184 (N_18184,N_15226,N_12220);
or U18185 (N_18185,N_12489,N_14071);
nor U18186 (N_18186,N_13538,N_15172);
and U18187 (N_18187,N_13383,N_14667);
and U18188 (N_18188,N_16818,N_12006);
nand U18189 (N_18189,N_17908,N_16786);
or U18190 (N_18190,N_16654,N_15300);
nand U18191 (N_18191,N_14979,N_15045);
nand U18192 (N_18192,N_14203,N_15702);
nand U18193 (N_18193,N_13562,N_15608);
xor U18194 (N_18194,N_17360,N_13575);
nand U18195 (N_18195,N_15734,N_14001);
xor U18196 (N_18196,N_16674,N_13140);
xor U18197 (N_18197,N_16072,N_14537);
xnor U18198 (N_18198,N_15353,N_15239);
or U18199 (N_18199,N_16424,N_14749);
nand U18200 (N_18200,N_16246,N_17346);
and U18201 (N_18201,N_12778,N_14233);
xor U18202 (N_18202,N_14721,N_13481);
nand U18203 (N_18203,N_16462,N_17036);
or U18204 (N_18204,N_13547,N_12779);
or U18205 (N_18205,N_17563,N_17838);
xnor U18206 (N_18206,N_14297,N_12253);
and U18207 (N_18207,N_15892,N_14294);
xor U18208 (N_18208,N_15117,N_14401);
or U18209 (N_18209,N_15418,N_17354);
nand U18210 (N_18210,N_17522,N_13511);
nand U18211 (N_18211,N_12783,N_16706);
and U18212 (N_18212,N_15061,N_12719);
xor U18213 (N_18213,N_16166,N_12419);
nand U18214 (N_18214,N_16086,N_15967);
or U18215 (N_18215,N_13916,N_12628);
nor U18216 (N_18216,N_15835,N_12609);
and U18217 (N_18217,N_14738,N_13026);
and U18218 (N_18218,N_15020,N_17319);
xor U18219 (N_18219,N_16893,N_12044);
nor U18220 (N_18220,N_14733,N_15364);
nor U18221 (N_18221,N_13868,N_14049);
or U18222 (N_18222,N_14634,N_16022);
or U18223 (N_18223,N_13030,N_12343);
and U18224 (N_18224,N_14279,N_14585);
and U18225 (N_18225,N_12633,N_12630);
nor U18226 (N_18226,N_14422,N_15715);
nor U18227 (N_18227,N_14905,N_15343);
xnor U18228 (N_18228,N_13284,N_17208);
or U18229 (N_18229,N_14811,N_16029);
nor U18230 (N_18230,N_15312,N_14984);
xnor U18231 (N_18231,N_17807,N_13006);
nor U18232 (N_18232,N_17705,N_15947);
or U18233 (N_18233,N_17869,N_14463);
and U18234 (N_18234,N_17479,N_12425);
and U18235 (N_18235,N_17040,N_15774);
and U18236 (N_18236,N_15915,N_13167);
and U18237 (N_18237,N_14997,N_15076);
and U18238 (N_18238,N_14715,N_17562);
or U18239 (N_18239,N_13501,N_12482);
xor U18240 (N_18240,N_17678,N_12816);
xor U18241 (N_18241,N_12422,N_12332);
or U18242 (N_18242,N_13073,N_12651);
and U18243 (N_18243,N_13642,N_13402);
nand U18244 (N_18244,N_12758,N_14791);
nor U18245 (N_18245,N_17156,N_14743);
nor U18246 (N_18246,N_13206,N_12617);
nor U18247 (N_18247,N_15211,N_13632);
or U18248 (N_18248,N_17475,N_13907);
or U18249 (N_18249,N_12179,N_12511);
nand U18250 (N_18250,N_14508,N_15140);
nor U18251 (N_18251,N_16603,N_15464);
or U18252 (N_18252,N_15263,N_15457);
nor U18253 (N_18253,N_15854,N_12102);
xnor U18254 (N_18254,N_15416,N_16465);
or U18255 (N_18255,N_17073,N_12632);
and U18256 (N_18256,N_13236,N_17938);
nor U18257 (N_18257,N_14063,N_14466);
nor U18258 (N_18258,N_17187,N_14804);
xnor U18259 (N_18259,N_15820,N_16487);
xnor U18260 (N_18260,N_16047,N_16236);
xnor U18261 (N_18261,N_13389,N_17407);
nor U18262 (N_18262,N_17799,N_15387);
xnor U18263 (N_18263,N_14105,N_15022);
or U18264 (N_18264,N_14788,N_16821);
or U18265 (N_18265,N_14044,N_17204);
and U18266 (N_18266,N_13619,N_13198);
xor U18267 (N_18267,N_14348,N_12833);
nor U18268 (N_18268,N_13845,N_13055);
xnor U18269 (N_18269,N_17698,N_16602);
nor U18270 (N_18270,N_12640,N_16118);
or U18271 (N_18271,N_16368,N_16121);
nor U18272 (N_18272,N_12652,N_14341);
nor U18273 (N_18273,N_13103,N_12729);
xor U18274 (N_18274,N_15204,N_13021);
and U18275 (N_18275,N_12256,N_13626);
nor U18276 (N_18276,N_15728,N_15642);
and U18277 (N_18277,N_17744,N_17979);
nor U18278 (N_18278,N_13613,N_14588);
nand U18279 (N_18279,N_16241,N_15578);
nor U18280 (N_18280,N_12749,N_15354);
xor U18281 (N_18281,N_16099,N_17458);
or U18282 (N_18282,N_12352,N_13141);
or U18283 (N_18283,N_15638,N_17413);
nand U18284 (N_18284,N_12858,N_14187);
xor U18285 (N_18285,N_15135,N_13148);
xnor U18286 (N_18286,N_12810,N_13860);
or U18287 (N_18287,N_17382,N_16171);
nor U18288 (N_18288,N_17939,N_17128);
nor U18289 (N_18289,N_15264,N_15518);
nand U18290 (N_18290,N_17294,N_17203);
xnor U18291 (N_18291,N_15762,N_12786);
nand U18292 (N_18292,N_15754,N_14384);
nand U18293 (N_18293,N_15616,N_12580);
nand U18294 (N_18294,N_16413,N_14343);
nor U18295 (N_18295,N_14366,N_17366);
xnor U18296 (N_18296,N_15631,N_15471);
nand U18297 (N_18297,N_12751,N_14878);
and U18298 (N_18298,N_16437,N_12299);
xor U18299 (N_18299,N_14812,N_15348);
or U18300 (N_18300,N_13071,N_16870);
or U18301 (N_18301,N_12196,N_17210);
or U18302 (N_18302,N_12275,N_17848);
or U18303 (N_18303,N_14093,N_17246);
xor U18304 (N_18304,N_15360,N_15115);
and U18305 (N_18305,N_14516,N_14283);
xnor U18306 (N_18306,N_16993,N_16094);
and U18307 (N_18307,N_14259,N_15191);
xor U18308 (N_18308,N_13661,N_12273);
or U18309 (N_18309,N_17336,N_14406);
xnor U18310 (N_18310,N_15572,N_12838);
nor U18311 (N_18311,N_17523,N_13480);
xnor U18312 (N_18312,N_16434,N_12803);
xor U18313 (N_18313,N_17102,N_16430);
or U18314 (N_18314,N_12663,N_16527);
or U18315 (N_18315,N_13356,N_12791);
or U18316 (N_18316,N_15549,N_12587);
and U18317 (N_18317,N_14928,N_14894);
and U18318 (N_18318,N_17737,N_15103);
nand U18319 (N_18319,N_16835,N_13963);
nor U18320 (N_18320,N_17345,N_16997);
xnor U18321 (N_18321,N_13201,N_14112);
or U18322 (N_18322,N_14476,N_12936);
or U18323 (N_18323,N_17127,N_17020);
nand U18324 (N_18324,N_13144,N_16860);
xor U18325 (N_18325,N_14443,N_12576);
nand U18326 (N_18326,N_15447,N_13936);
and U18327 (N_18327,N_13693,N_16544);
and U18328 (N_18328,N_15168,N_16956);
nor U18329 (N_18329,N_15806,N_12894);
or U18330 (N_18330,N_14572,N_16333);
or U18331 (N_18331,N_17851,N_14940);
and U18332 (N_18332,N_12818,N_13968);
nor U18333 (N_18333,N_15456,N_17820);
and U18334 (N_18334,N_12579,N_16117);
or U18335 (N_18335,N_13827,N_12378);
nor U18336 (N_18336,N_12518,N_16653);
nand U18337 (N_18337,N_13257,N_13278);
xnor U18338 (N_18338,N_16883,N_12028);
nor U18339 (N_18339,N_12624,N_16725);
nand U18340 (N_18340,N_17677,N_14240);
nor U18341 (N_18341,N_14663,N_12946);
or U18342 (N_18342,N_12451,N_14950);
and U18343 (N_18343,N_14414,N_17198);
and U18344 (N_18344,N_12091,N_17192);
or U18345 (N_18345,N_15258,N_12954);
nand U18346 (N_18346,N_14630,N_16946);
nor U18347 (N_18347,N_16978,N_16197);
xor U18348 (N_18348,N_12496,N_15992);
nand U18349 (N_18349,N_12737,N_15689);
nand U18350 (N_18350,N_13735,N_12891);
or U18351 (N_18351,N_12885,N_16234);
nor U18352 (N_18352,N_16775,N_12329);
and U18353 (N_18353,N_16735,N_15536);
xnor U18354 (N_18354,N_14713,N_14897);
nor U18355 (N_18355,N_12921,N_12750);
and U18356 (N_18356,N_15817,N_16803);
nand U18357 (N_18357,N_14859,N_14392);
and U18358 (N_18358,N_16650,N_17349);
and U18359 (N_18359,N_13706,N_13410);
xor U18360 (N_18360,N_17758,N_17231);
nor U18361 (N_18361,N_13159,N_15830);
nor U18362 (N_18362,N_15121,N_16302);
xnor U18363 (N_18363,N_14218,N_12669);
and U18364 (N_18364,N_17704,N_14826);
nor U18365 (N_18365,N_17921,N_16388);
nand U18366 (N_18366,N_12627,N_17789);
or U18367 (N_18367,N_14924,N_17796);
or U18368 (N_18368,N_16460,N_13724);
or U18369 (N_18369,N_16509,N_17505);
and U18370 (N_18370,N_16903,N_13049);
and U18371 (N_18371,N_14691,N_16091);
or U18372 (N_18372,N_17502,N_13542);
xnor U18373 (N_18373,N_17605,N_14355);
and U18374 (N_18374,N_16528,N_14595);
nor U18375 (N_18375,N_12205,N_17663);
xor U18376 (N_18376,N_17745,N_16854);
or U18377 (N_18377,N_13399,N_13367);
nand U18378 (N_18378,N_16466,N_16387);
nor U18379 (N_18379,N_14367,N_17843);
xnor U18380 (N_18380,N_17607,N_16078);
or U18381 (N_18381,N_15778,N_14919);
nand U18382 (N_18382,N_17201,N_14149);
nor U18383 (N_18383,N_15664,N_17794);
or U18384 (N_18384,N_17317,N_14995);
nor U18385 (N_18385,N_12712,N_13222);
xor U18386 (N_18386,N_16731,N_17941);
nand U18387 (N_18387,N_14573,N_15041);
and U18388 (N_18388,N_14574,N_16168);
nor U18389 (N_18389,N_15444,N_15805);
nand U18390 (N_18390,N_17912,N_12672);
xor U18391 (N_18391,N_15871,N_16192);
nor U18392 (N_18392,N_13854,N_12667);
nor U18393 (N_18393,N_14321,N_15313);
or U18394 (N_18394,N_12218,N_14120);
nor U18395 (N_18395,N_12978,N_16369);
nor U18396 (N_18396,N_16406,N_12434);
xnor U18397 (N_18397,N_13969,N_13363);
nand U18398 (N_18398,N_17543,N_15335);
and U18399 (N_18399,N_16844,N_15604);
or U18400 (N_18400,N_16385,N_16810);
nand U18401 (N_18401,N_17269,N_14123);
xor U18402 (N_18402,N_17278,N_17292);
nand U18403 (N_18403,N_16962,N_13207);
nand U18404 (N_18404,N_13696,N_12702);
xor U18405 (N_18405,N_12949,N_15613);
nor U18406 (N_18406,N_14925,N_14908);
and U18407 (N_18407,N_12030,N_17793);
and U18408 (N_18408,N_15544,N_16887);
and U18409 (N_18409,N_12845,N_17824);
xnor U18410 (N_18410,N_16888,N_12528);
or U18411 (N_18411,N_14542,N_16346);
and U18412 (N_18412,N_16320,N_13685);
xor U18413 (N_18413,N_13490,N_17962);
nor U18414 (N_18414,N_13676,N_17747);
nand U18415 (N_18415,N_15413,N_16484);
xor U18416 (N_18416,N_12261,N_16547);
and U18417 (N_18417,N_12645,N_13246);
or U18418 (N_18418,N_15735,N_17332);
nand U18419 (N_18419,N_16652,N_15290);
nor U18420 (N_18420,N_15410,N_16337);
xnor U18421 (N_18421,N_15256,N_14464);
or U18422 (N_18422,N_16111,N_12358);
or U18423 (N_18423,N_12621,N_16181);
xnor U18424 (N_18424,N_13586,N_16451);
nand U18425 (N_18425,N_16056,N_17665);
or U18426 (N_18426,N_16549,N_13483);
or U18427 (N_18427,N_13396,N_16318);
and U18428 (N_18428,N_16812,N_12436);
xnor U18429 (N_18429,N_13042,N_17289);
xor U18430 (N_18430,N_15834,N_15986);
xnor U18431 (N_18431,N_17658,N_13419);
xor U18432 (N_18432,N_14262,N_15870);
and U18433 (N_18433,N_16167,N_16377);
and U18434 (N_18434,N_13835,N_15356);
nor U18435 (N_18435,N_15196,N_17258);
and U18436 (N_18436,N_13606,N_13545);
and U18437 (N_18437,N_14830,N_16729);
nor U18438 (N_18438,N_16630,N_16394);
nand U18439 (N_18439,N_16873,N_14193);
xor U18440 (N_18440,N_12155,N_17117);
or U18441 (N_18441,N_15988,N_15635);
nor U18442 (N_18442,N_14418,N_12190);
nor U18443 (N_18443,N_14800,N_12594);
xor U18444 (N_18444,N_17104,N_17171);
xnor U18445 (N_18445,N_13373,N_13997);
xor U18446 (N_18446,N_14697,N_16127);
nand U18447 (N_18447,N_14135,N_17280);
and U18448 (N_18448,N_16513,N_14681);
and U18449 (N_18449,N_17714,N_16294);
xor U18450 (N_18450,N_16651,N_17091);
nor U18451 (N_18451,N_17021,N_14395);
or U18452 (N_18452,N_17860,N_14412);
and U18453 (N_18453,N_17323,N_13185);
or U18454 (N_18454,N_17151,N_17372);
or U18455 (N_18455,N_13405,N_12367);
nor U18456 (N_18456,N_16726,N_13645);
or U18457 (N_18457,N_13698,N_13334);
xor U18458 (N_18458,N_14851,N_16421);
nand U18459 (N_18459,N_13168,N_12679);
xor U18460 (N_18460,N_14277,N_13734);
and U18461 (N_18461,N_15956,N_14612);
xor U18462 (N_18462,N_13149,N_13163);
and U18463 (N_18463,N_13248,N_17840);
xnor U18464 (N_18464,N_12026,N_16263);
or U18465 (N_18465,N_12806,N_13468);
or U18466 (N_18466,N_16065,N_16983);
and U18467 (N_18467,N_13579,N_14823);
nand U18468 (N_18468,N_17694,N_16305);
nor U18469 (N_18469,N_14329,N_16708);
or U18470 (N_18470,N_13832,N_12144);
nor U18471 (N_18471,N_12386,N_17619);
xor U18472 (N_18472,N_15467,N_16865);
nand U18473 (N_18473,N_13192,N_13543);
nand U18474 (N_18474,N_14521,N_15185);
and U18475 (N_18475,N_17286,N_14408);
and U18476 (N_18476,N_15512,N_16124);
or U18477 (N_18477,N_14382,N_16218);
or U18478 (N_18478,N_17875,N_14835);
nor U18479 (N_18479,N_13258,N_12064);
and U18480 (N_18480,N_16845,N_15099);
xnor U18481 (N_18481,N_13679,N_15063);
nor U18482 (N_18482,N_14030,N_15882);
xor U18483 (N_18483,N_17247,N_13106);
or U18484 (N_18484,N_13762,N_15640);
nand U18485 (N_18485,N_12323,N_14388);
xor U18486 (N_18486,N_14456,N_17584);
nand U18487 (N_18487,N_17486,N_16678);
nor U18488 (N_18488,N_13918,N_12126);
xor U18489 (N_18489,N_13417,N_17441);
or U18490 (N_18490,N_16741,N_15505);
nand U18491 (N_18491,N_13295,N_13173);
and U18492 (N_18492,N_12900,N_15486);
xnor U18493 (N_18493,N_12883,N_12105);
nand U18494 (N_18494,N_14509,N_14352);
and U18495 (N_18495,N_14679,N_12765);
or U18496 (N_18496,N_17402,N_13708);
and U18497 (N_18497,N_13444,N_16514);
nor U18498 (N_18498,N_16384,N_12339);
and U18499 (N_18499,N_13397,N_13960);
xor U18500 (N_18500,N_16429,N_13175);
and U18501 (N_18501,N_12961,N_16449);
nand U18502 (N_18502,N_17017,N_12509);
nor U18503 (N_18503,N_12271,N_17008);
xor U18504 (N_18504,N_16737,N_12120);
or U18505 (N_18505,N_13571,N_16321);
nor U18506 (N_18506,N_13528,N_14720);
nor U18507 (N_18507,N_14363,N_16064);
xor U18508 (N_18508,N_13443,N_17412);
xor U18509 (N_18509,N_17748,N_17733);
and U18510 (N_18510,N_17683,N_15420);
nor U18511 (N_18511,N_16505,N_16407);
and U18512 (N_18512,N_17915,N_14441);
xnor U18513 (N_18513,N_13567,N_16894);
nand U18514 (N_18514,N_15133,N_17533);
nand U18515 (N_18515,N_12532,N_15425);
nor U18516 (N_18516,N_12065,N_13731);
or U18517 (N_18517,N_14332,N_17193);
or U18518 (N_18518,N_15738,N_16601);
xor U18519 (N_18519,N_12055,N_14973);
nand U18520 (N_18520,N_14196,N_15427);
and U18521 (N_18521,N_17273,N_12267);
nor U18522 (N_18522,N_14312,N_13193);
nor U18523 (N_18523,N_16027,N_15673);
or U18524 (N_18524,N_12701,N_12068);
xor U18525 (N_18525,N_12658,N_12305);
xor U18526 (N_18526,N_17334,N_17501);
nor U18527 (N_18527,N_14903,N_12745);
nand U18528 (N_18528,N_16247,N_17559);
or U18529 (N_18529,N_16612,N_17649);
and U18530 (N_18530,N_16014,N_13271);
xnor U18531 (N_18531,N_14672,N_17066);
nor U18532 (N_18532,N_17929,N_17906);
nor U18533 (N_18533,N_16663,N_16762);
or U18534 (N_18534,N_17549,N_13223);
or U18535 (N_18535,N_17792,N_15795);
nand U18536 (N_18536,N_16291,N_16736);
xnor U18537 (N_18537,N_14344,N_16910);
or U18538 (N_18538,N_14038,N_13647);
nand U18539 (N_18539,N_13028,N_17148);
nor U18540 (N_18540,N_13067,N_12398);
and U18541 (N_18541,N_16617,N_17062);
and U18542 (N_18542,N_16992,N_14276);
xnor U18543 (N_18543,N_16567,N_12551);
nor U18544 (N_18544,N_17827,N_14242);
nor U18545 (N_18545,N_12966,N_16202);
and U18546 (N_18546,N_14350,N_13498);
xnor U18547 (N_18547,N_17923,N_16089);
nand U18548 (N_18548,N_15804,N_14028);
nand U18549 (N_18549,N_15917,N_13796);
nand U18550 (N_18550,N_17469,N_16782);
xnor U18551 (N_18551,N_16938,N_12995);
or U18552 (N_18552,N_17177,N_13518);
and U18553 (N_18553,N_16112,N_17917);
and U18554 (N_18554,N_14250,N_13840);
xnor U18555 (N_18555,N_13178,N_12093);
nor U18556 (N_18556,N_14169,N_12184);
nor U18557 (N_18557,N_15537,N_13653);
or U18558 (N_18558,N_17245,N_17045);
nand U18559 (N_18559,N_14616,N_15201);
and U18560 (N_18560,N_16771,N_15712);
and U18561 (N_18561,N_13061,N_17049);
xnor U18562 (N_18562,N_15351,N_15932);
or U18563 (N_18563,N_13099,N_17266);
xor U18564 (N_18564,N_12924,N_14039);
or U18565 (N_18565,N_15905,N_13687);
or U18566 (N_18566,N_16330,N_15180);
and U18567 (N_18567,N_15271,N_14357);
xor U18568 (N_18568,N_12938,N_16061);
or U18569 (N_18569,N_12502,N_12411);
nand U18570 (N_18570,N_15970,N_17257);
nor U18571 (N_18571,N_17988,N_16525);
nand U18572 (N_18572,N_14267,N_15181);
nor U18573 (N_18573,N_12897,N_15377);
nand U18574 (N_18574,N_13069,N_15644);
or U18575 (N_18575,N_14942,N_15474);
or U18576 (N_18576,N_13065,N_13374);
and U18577 (N_18577,N_16208,N_14618);
xnor U18578 (N_18578,N_15307,N_12606);
and U18579 (N_18579,N_17031,N_17847);
nand U18580 (N_18580,N_16904,N_16669);
xnor U18581 (N_18581,N_17119,N_15573);
or U18582 (N_18582,N_12836,N_13873);
nor U18583 (N_18583,N_14460,N_16042);
and U18584 (N_18584,N_12384,N_14445);
nor U18585 (N_18585,N_14870,N_12320);
nor U18586 (N_18586,N_16115,N_14496);
or U18587 (N_18587,N_17079,N_16960);
xor U18588 (N_18588,N_16309,N_14056);
nor U18589 (N_18589,N_17216,N_15202);
nand U18590 (N_18590,N_16559,N_15977);
nand U18591 (N_18591,N_12280,N_12867);
nand U18592 (N_18592,N_17139,N_12776);
or U18593 (N_18593,N_16574,N_14142);
xor U18594 (N_18594,N_17876,N_14251);
or U18595 (N_18595,N_17684,N_13225);
nor U18596 (N_18596,N_16051,N_12714);
xnor U18597 (N_18597,N_13924,N_12792);
and U18598 (N_18598,N_15249,N_12601);
nor U18599 (N_18599,N_17277,N_16343);
xnor U18600 (N_18600,N_17320,N_17397);
xnor U18601 (N_18601,N_15836,N_17880);
xnor U18602 (N_18602,N_16216,N_17039);
nor U18603 (N_18603,N_15029,N_12515);
and U18604 (N_18604,N_16046,N_13517);
xnor U18605 (N_18605,N_13142,N_15897);
nor U18606 (N_18606,N_15405,N_13755);
and U18607 (N_18607,N_17484,N_16342);
xor U18608 (N_18608,N_17751,N_12321);
xor U18609 (N_18609,N_17414,N_12631);
nor U18610 (N_18610,N_16215,N_14676);
xnor U18611 (N_18611,N_13387,N_12659);
or U18612 (N_18612,N_17433,N_13467);
nand U18613 (N_18613,N_12124,N_14532);
and U18614 (N_18614,N_12443,N_17467);
and U18615 (N_18615,N_12123,N_13370);
xnor U18616 (N_18616,N_17411,N_16842);
nor U18617 (N_18617,N_13814,N_15580);
xor U18618 (N_18618,N_17275,N_15533);
and U18619 (N_18619,N_13572,N_16209);
xnor U18620 (N_18620,N_16104,N_14387);
xnor U18621 (N_18621,N_12389,N_14622);
or U18622 (N_18622,N_13039,N_12178);
nor U18623 (N_18623,N_14225,N_16432);
xor U18624 (N_18624,N_13060,N_15862);
and U18625 (N_18625,N_14941,N_12839);
nand U18626 (N_18626,N_15401,N_14610);
or U18627 (N_18627,N_12084,N_15483);
and U18628 (N_18628,N_17318,N_12945);
or U18629 (N_18629,N_16587,N_15920);
xor U18630 (N_18630,N_14971,N_17830);
or U18631 (N_18631,N_15424,N_16286);
nand U18632 (N_18632,N_16995,N_16332);
or U18633 (N_18633,N_15961,N_17696);
and U18634 (N_18634,N_17446,N_13780);
or U18635 (N_18635,N_15792,N_16705);
or U18636 (N_18636,N_13436,N_16632);
and U18637 (N_18637,N_16195,N_14046);
xor U18638 (N_18638,N_17114,N_17652);
xnor U18639 (N_18639,N_17106,N_15525);
nor U18640 (N_18640,N_16068,N_13031);
or U18641 (N_18641,N_16753,N_15694);
xnor U18642 (N_18642,N_15362,N_16295);
or U18643 (N_18643,N_13066,N_17147);
nand U18644 (N_18644,N_12724,N_14773);
xnor U18645 (N_18645,N_13953,N_17517);
and U18646 (N_18646,N_16400,N_13648);
nand U18647 (N_18647,N_13292,N_13250);
or U18648 (N_18648,N_13896,N_16642);
and U18649 (N_18649,N_15665,N_16198);
or U18650 (N_18650,N_15607,N_14390);
xor U18651 (N_18651,N_17217,N_13920);
and U18652 (N_18652,N_13669,N_15724);
and U18653 (N_18653,N_17907,N_17973);
and U18654 (N_18654,N_14596,N_12114);
or U18655 (N_18655,N_13128,N_17136);
nor U18656 (N_18656,N_14625,N_12365);
or U18657 (N_18657,N_16675,N_12590);
nor U18658 (N_18658,N_17027,N_16826);
and U18659 (N_18659,N_14945,N_12637);
and U18660 (N_18660,N_12435,N_13782);
xor U18661 (N_18661,N_14400,N_13504);
nor U18662 (N_18662,N_17276,N_17916);
xnor U18663 (N_18663,N_14744,N_17440);
and U18664 (N_18664,N_17103,N_15916);
nand U18665 (N_18665,N_15611,N_15680);
xnor U18666 (N_18666,N_14007,N_16954);
xor U18667 (N_18667,N_16359,N_14889);
xnor U18668 (N_18668,N_16571,N_16442);
nand U18669 (N_18669,N_13458,N_13878);
nand U18670 (N_18670,N_17329,N_14615);
nor U18671 (N_18671,N_13381,N_16092);
xor U18672 (N_18672,N_14536,N_16785);
nand U18673 (N_18673,N_15350,N_14969);
or U18674 (N_18674,N_12689,N_15039);
nand U18675 (N_18675,N_12007,N_15031);
and U18676 (N_18676,N_16110,N_13083);
and U18677 (N_18677,N_13667,N_14768);
and U18678 (N_18678,N_17572,N_16336);
nand U18679 (N_18679,N_14862,N_14703);
nor U18680 (N_18680,N_13070,N_17034);
xnor U18681 (N_18681,N_16392,N_16698);
nand U18682 (N_18682,N_14221,N_16133);
nand U18683 (N_18683,N_12249,N_15955);
nor U18684 (N_18684,N_16832,N_14220);
or U18685 (N_18685,N_17244,N_17377);
and U18686 (N_18686,N_13546,N_13776);
nor U18687 (N_18687,N_17612,N_15110);
nand U18688 (N_18688,N_16183,N_17005);
nand U18689 (N_18689,N_16576,N_15855);
xnor U18690 (N_18690,N_14130,N_15701);
nor U18691 (N_18691,N_12804,N_14650);
or U18692 (N_18692,N_13470,N_16055);
nor U18693 (N_18693,N_15944,N_15906);
xnor U18694 (N_18694,N_12234,N_16949);
and U18695 (N_18695,N_13794,N_15408);
or U18696 (N_18696,N_17762,N_14956);
or U18697 (N_18697,N_12420,N_12523);
xor U18698 (N_18698,N_16493,N_12828);
and U18699 (N_18699,N_14646,N_13075);
nand U18700 (N_18700,N_12716,N_12958);
or U18701 (N_18701,N_12154,N_14922);
nand U18702 (N_18702,N_13789,N_17808);
and U18703 (N_18703,N_13804,N_13862);
and U18704 (N_18704,N_15047,N_13429);
nand U18705 (N_18705,N_12668,N_14064);
and U18706 (N_18706,N_17989,N_12063);
nand U18707 (N_18707,N_16436,N_14389);
and U18708 (N_18708,N_17987,N_12908);
nand U18709 (N_18709,N_12643,N_12024);
xor U18710 (N_18710,N_16416,N_17703);
nor U18711 (N_18711,N_13226,N_16756);
xor U18712 (N_18712,N_12244,N_16494);
xor U18713 (N_18713,N_16244,N_16554);
or U18714 (N_18714,N_16713,N_16150);
or U18715 (N_18715,N_12298,N_12794);
or U18716 (N_18716,N_15489,N_14798);
or U18717 (N_18717,N_12232,N_15659);
and U18718 (N_18718,N_14852,N_16524);
xor U18719 (N_18719,N_12066,N_14068);
or U18720 (N_18720,N_13714,N_14917);
nand U18721 (N_18721,N_17076,N_16701);
or U18722 (N_18722,N_12822,N_13981);
and U18723 (N_18723,N_14361,N_14469);
nand U18724 (N_18724,N_17109,N_15766);
xnor U18725 (N_18725,N_17029,N_15589);
nand U18726 (N_18726,N_14141,N_15831);
and U18727 (N_18727,N_14066,N_15938);
and U18728 (N_18728,N_16296,N_13331);
nor U18729 (N_18729,N_14944,N_13768);
and U18730 (N_18730,N_14967,N_15301);
xor U18731 (N_18731,N_12458,N_14892);
or U18732 (N_18732,N_14690,N_12834);
nand U18733 (N_18733,N_16508,N_16600);
xnor U18734 (N_18734,N_15866,N_15639);
xnor U18735 (N_18735,N_14004,N_13394);
and U18736 (N_18736,N_12855,N_17010);
and U18737 (N_18737,N_16825,N_13253);
nor U18738 (N_18738,N_13786,N_17352);
or U18739 (N_18739,N_15618,N_15219);
nor U18740 (N_18740,N_15048,N_17780);
or U18741 (N_18741,N_12394,N_16766);
and U18742 (N_18742,N_12204,N_13717);
nand U18743 (N_18743,N_17296,N_14311);
nand U18744 (N_18744,N_13496,N_12519);
and U18745 (N_18745,N_12974,N_13652);
nor U18746 (N_18746,N_13927,N_12023);
xnor U18747 (N_18747,N_16059,N_17381);
and U18748 (N_18748,N_15587,N_15560);
or U18749 (N_18749,N_16228,N_16217);
nand U18750 (N_18750,N_16546,N_13447);
xor U18751 (N_18751,N_16098,N_12678);
nand U18752 (N_18752,N_14310,N_12071);
nor U18753 (N_18753,N_13153,N_17012);
nor U18754 (N_18754,N_12597,N_13027);
or U18755 (N_18755,N_13462,N_14497);
nor U18756 (N_18756,N_16152,N_14753);
or U18757 (N_18757,N_16765,N_15297);
and U18758 (N_18758,N_14827,N_16201);
xnor U18759 (N_18759,N_14752,N_13255);
nor U18760 (N_18760,N_12477,N_17690);
or U18761 (N_18761,N_17219,N_17124);
nand U18762 (N_18762,N_15946,N_13346);
nand U18763 (N_18763,N_14589,N_17328);
and U18764 (N_18764,N_13884,N_17833);
nand U18765 (N_18765,N_13700,N_13306);
or U18766 (N_18766,N_14305,N_16572);
nand U18767 (N_18767,N_15901,N_12241);
xnor U18768 (N_18768,N_16886,N_12541);
or U18769 (N_18769,N_16031,N_14795);
and U18770 (N_18770,N_14677,N_14356);
and U18771 (N_18771,N_15654,N_16583);
and U18772 (N_18772,N_17300,N_15919);
or U18773 (N_18773,N_17461,N_15698);
or U18774 (N_18774,N_15379,N_14556);
or U18775 (N_18775,N_16339,N_13959);
nand U18776 (N_18776,N_16533,N_13208);
and U18777 (N_18777,N_17998,N_16366);
or U18778 (N_18778,N_12462,N_14241);
xor U18779 (N_18779,N_14134,N_13994);
nor U18780 (N_18780,N_16936,N_14597);
and U18781 (N_18781,N_17451,N_16807);
nand U18782 (N_18782,N_12871,N_17325);
xor U18783 (N_18783,N_17421,N_15334);
nand U18784 (N_18784,N_16352,N_12257);
or U18785 (N_18785,N_13995,N_16898);
or U18786 (N_18786,N_15237,N_13202);
xnor U18787 (N_18787,N_12363,N_14191);
and U18788 (N_18788,N_15026,N_13894);
xnor U18789 (N_18789,N_14560,N_13656);
nand U18790 (N_18790,N_12131,N_15106);
nand U18791 (N_18791,N_17432,N_14528);
and U18792 (N_18792,N_14248,N_12875);
and U18793 (N_18793,N_12505,N_12308);
or U18794 (N_18794,N_13848,N_16820);
nor U18795 (N_18795,N_16789,N_15238);
nor U18796 (N_18796,N_16951,N_14824);
nand U18797 (N_18797,N_17617,N_12206);
nor U18798 (N_18798,N_16441,N_17850);
nand U18799 (N_18799,N_14008,N_14467);
or U18800 (N_18800,N_12821,N_15429);
xnor U18801 (N_18801,N_14895,N_15620);
or U18802 (N_18802,N_14421,N_17868);
or U18803 (N_18803,N_16670,N_13304);
xnor U18804 (N_18804,N_16227,N_17558);
and U18805 (N_18805,N_14165,N_15019);
nand U18806 (N_18806,N_13365,N_12904);
xnor U18807 (N_18807,N_16358,N_14512);
and U18808 (N_18808,N_14340,N_16439);
and U18809 (N_18809,N_15937,N_13146);
or U18810 (N_18810,N_14902,N_14050);
or U18811 (N_18811,N_17709,N_12004);
xor U18812 (N_18812,N_13325,N_15279);
and U18813 (N_18813,N_16458,N_15164);
and U18814 (N_18814,N_15093,N_16231);
xnor U18815 (N_18815,N_14420,N_14249);
nor U18816 (N_18816,N_15554,N_12619);
nand U18817 (N_18817,N_16354,N_12015);
or U18818 (N_18818,N_14631,N_12876);
nor U18819 (N_18819,N_14728,N_16848);
or U18820 (N_18820,N_16169,N_12346);
nand U18821 (N_18821,N_14438,N_17316);
nand U18822 (N_18822,N_14090,N_14323);
nand U18823 (N_18823,N_14170,N_14683);
or U18824 (N_18824,N_16132,N_15503);
and U18825 (N_18825,N_12222,N_12387);
nand U18826 (N_18826,N_13293,N_15161);
and U18827 (N_18827,N_14033,N_12289);
or U18828 (N_18828,N_13883,N_15628);
or U18829 (N_18829,N_13903,N_13811);
xnor U18830 (N_18830,N_13442,N_12578);
xor U18831 (N_18831,N_12101,N_14180);
or U18832 (N_18832,N_16847,N_16428);
nor U18833 (N_18833,N_13270,N_17503);
nor U18834 (N_18834,N_16536,N_12666);
or U18835 (N_18835,N_14236,N_13961);
and U18836 (N_18836,N_16692,N_15562);
or U18837 (N_18837,N_13692,N_14119);
nand U18838 (N_18838,N_15478,N_13520);
xor U18839 (N_18839,N_16953,N_16019);
and U18840 (N_18840,N_16969,N_15825);
or U18841 (N_18841,N_17977,N_15720);
nand U18842 (N_18842,N_12438,N_13116);
nand U18843 (N_18843,N_15904,N_14304);
or U18844 (N_18844,N_17340,N_12360);
and U18845 (N_18845,N_14060,N_15760);
or U18846 (N_18846,N_15199,N_16637);
nor U18847 (N_18847,N_12809,N_13286);
or U18848 (N_18848,N_17060,N_17307);
or U18849 (N_18849,N_13578,N_12793);
and U18850 (N_18850,N_14655,N_13787);
or U18851 (N_18851,N_12802,N_13964);
and U18852 (N_18852,N_17384,N_13872);
or U18853 (N_18853,N_12918,N_14522);
or U18854 (N_18854,N_12798,N_17760);
or U18855 (N_18855,N_13047,N_17448);
or U18856 (N_18856,N_15843,N_16143);
and U18857 (N_18857,N_14865,N_16474);
nor U18858 (N_18858,N_17024,N_17033);
and U18859 (N_18859,N_13908,N_13131);
or U18860 (N_18860,N_15397,N_17633);
or U18861 (N_18861,N_15716,N_15685);
nand U18862 (N_18862,N_13625,N_17359);
nor U18863 (N_18863,N_17729,N_15332);
xnor U18864 (N_18864,N_16634,N_15233);
nand U18865 (N_18865,N_16878,N_13074);
nand U18866 (N_18866,N_16746,N_14034);
xnor U18867 (N_18867,N_17811,N_16136);
nor U18868 (N_18868,N_14162,N_14306);
xnor U18869 (N_18869,N_14568,N_17944);
nor U18870 (N_18870,N_14483,N_12074);
xor U18871 (N_18871,N_16799,N_15714);
or U18872 (N_18872,N_16656,N_16710);
xnor U18873 (N_18873,N_16945,N_16560);
xnor U18874 (N_18874,N_12112,N_15609);
and U18875 (N_18875,N_17872,N_13853);
and U18876 (N_18876,N_12741,N_12832);
nor U18877 (N_18877,N_15842,N_16261);
nand U18878 (N_18878,N_16390,N_16084);
nor U18879 (N_18879,N_16446,N_16130);
nand U18880 (N_18880,N_14565,N_17874);
nand U18881 (N_18881,N_12564,N_13837);
nor U18882 (N_18882,N_15182,N_17200);
xnor U18883 (N_18883,N_13090,N_16050);
xor U18884 (N_18884,N_15908,N_12861);
or U18885 (N_18885,N_17548,N_15773);
nor U18886 (N_18886,N_12345,N_15240);
and U18887 (N_18887,N_14527,N_13785);
and U18888 (N_18888,N_16176,N_14855);
and U18889 (N_18889,N_14533,N_16165);
xor U18890 (N_18890,N_15145,N_13182);
or U18891 (N_18891,N_15441,N_16284);
nor U18892 (N_18892,N_14453,N_14948);
nor U18893 (N_18893,N_15687,N_15677);
nor U18894 (N_18894,N_17664,N_17163);
or U18895 (N_18895,N_14666,N_15395);
and U18896 (N_18896,N_16360,N_15756);
xnor U18897 (N_18897,N_13733,N_14300);
nand U18898 (N_18898,N_15167,N_12730);
nor U18899 (N_18899,N_12122,N_14146);
and U18900 (N_18900,N_13320,N_12830);
or U18901 (N_18901,N_13338,N_12174);
nor U18902 (N_18902,N_12906,N_17866);
xor U18903 (N_18903,N_17756,N_13983);
and U18904 (N_18904,N_16570,N_17009);
and U18905 (N_18905,N_12495,N_13247);
or U18906 (N_18906,N_15190,N_12703);
nor U18907 (N_18907,N_17770,N_13328);
nor U18908 (N_18908,N_15585,N_16975);
and U18909 (N_18909,N_17560,N_13943);
nand U18910 (N_18910,N_15719,N_12159);
nand U18911 (N_18911,N_16517,N_12448);
and U18912 (N_18912,N_16809,N_15257);
nor U18913 (N_18913,N_16159,N_15118);
xor U18914 (N_18914,N_15520,N_15746);
and U18915 (N_18915,N_15059,N_16912);
or U18916 (N_18916,N_13819,N_17504);
and U18917 (N_18917,N_15557,N_15526);
nor U18918 (N_18918,N_15891,N_17395);
and U18919 (N_18919,N_12335,N_12250);
or U18920 (N_18920,N_17858,N_17693);
nor U18921 (N_18921,N_15584,N_16037);
or U18922 (N_18922,N_17075,N_16974);
nand U18923 (N_18923,N_16913,N_12767);
xnor U18924 (N_18924,N_16239,N_12338);
or U18925 (N_18925,N_12075,N_14874);
nand U18926 (N_18926,N_17942,N_15949);
nor U18927 (N_18927,N_12182,N_15291);
nand U18928 (N_18928,N_17001,N_16070);
nand U18929 (N_18929,N_16024,N_13045);
or U18930 (N_18930,N_17519,N_14083);
nand U18931 (N_18931,N_14793,N_12520);
or U18932 (N_18932,N_12811,N_15314);
nor U18933 (N_18933,N_12516,N_15220);
and U18934 (N_18934,N_17613,N_14500);
or U18935 (N_18935,N_12304,N_17002);
and U18936 (N_18936,N_13276,N_17426);
nor U18937 (N_18937,N_17087,N_16327);
or U18938 (N_18938,N_14214,N_12022);
nor U18939 (N_18939,N_14490,N_13034);
and U18940 (N_18940,N_12990,N_15636);
nand U18941 (N_18941,N_15529,N_14434);
nor U18942 (N_18942,N_15186,N_12229);
nor U18943 (N_18943,N_16947,N_15023);
or U18944 (N_18944,N_16256,N_12322);
xor U18945 (N_18945,N_17357,N_15384);
and U18946 (N_18946,N_15653,N_16749);
or U18947 (N_18947,N_17285,N_12295);
nand U18948 (N_18948,N_15727,N_15993);
xor U18949 (N_18949,N_17555,N_14981);
or U18950 (N_18950,N_16568,N_16404);
or U18951 (N_18951,N_13563,N_12753);
xnor U18952 (N_18952,N_12180,N_16264);
or U18953 (N_18953,N_16412,N_12755);
and U18954 (N_18954,N_15268,N_13984);
nor U18955 (N_18955,N_15452,N_13158);
or U18956 (N_18956,N_15422,N_15612);
and U18957 (N_18957,N_17226,N_12291);
or U18958 (N_18958,N_14688,N_17783);
nor U18959 (N_18959,N_13783,N_14019);
or U18960 (N_18960,N_14641,N_14353);
nor U18961 (N_18961,N_13110,N_17248);
and U18962 (N_18962,N_17281,N_12925);
xor U18963 (N_18963,N_14347,N_12296);
and U18964 (N_18964,N_15838,N_13503);
nor U18965 (N_18965,N_12670,N_16137);
nor U18966 (N_18966,N_16875,N_14805);
nand U18967 (N_18967,N_14765,N_13748);
or U18968 (N_18968,N_12086,N_16718);
and U18969 (N_18969,N_16395,N_17202);
nor U18970 (N_18970,N_16119,N_15923);
nor U18971 (N_18971,N_16422,N_13157);
nor U18972 (N_18972,N_13566,N_17631);
xnor U18973 (N_18973,N_12600,N_16823);
nor U18974 (N_18974,N_17734,N_14148);
nand U18975 (N_18975,N_15545,N_14699);
and U18976 (N_18976,N_12487,N_17982);
and U18977 (N_18977,N_17849,N_15428);
nor U18978 (N_18978,N_17101,N_12760);
xor U18979 (N_18979,N_17972,N_12251);
xor U18980 (N_18980,N_17648,N_16874);
or U18981 (N_18981,N_17803,N_15078);
nand U18982 (N_18982,N_12999,N_12274);
nand U18983 (N_18983,N_17406,N_15095);
nand U18984 (N_18984,N_15455,N_13716);
xor U18985 (N_18985,N_13430,N_17070);
nand U18986 (N_18986,N_17568,N_14686);
xor U18987 (N_18987,N_14286,N_15042);
xnor U18988 (N_18988,N_14970,N_13123);
and U18989 (N_18989,N_15435,N_15524);
nor U18990 (N_18990,N_12087,N_12468);
or U18991 (N_18991,N_15684,N_15890);
xnor U18992 (N_18992,N_16105,N_17436);
xor U18993 (N_18993,N_12485,N_13059);
and U18994 (N_18994,N_14575,N_17781);
and U18995 (N_18995,N_15209,N_15248);
nor U18996 (N_18996,N_12555,N_12359);
xor U18997 (N_18997,N_14296,N_15927);
nand U18998 (N_18998,N_15592,N_17741);
or U18999 (N_18999,N_15841,N_16999);
xor U19000 (N_19000,N_13495,N_12302);
nor U19001 (N_19001,N_14336,N_14157);
xnor U19002 (N_19002,N_13771,N_12780);
nor U19003 (N_19003,N_17363,N_14047);
and U19004 (N_19004,N_12340,N_13280);
and U19005 (N_19005,N_12175,N_16397);
nor U19006 (N_19006,N_14108,N_12569);
and U19007 (N_19007,N_14633,N_14635);
or U19008 (N_19008,N_15881,N_12403);
or U19009 (N_19009,N_17170,N_12466);
or U19010 (N_19010,N_14949,N_12848);
nor U19011 (N_19011,N_13766,N_13324);
nand U19012 (N_19012,N_13933,N_12787);
xor U19013 (N_19013,N_12919,N_14029);
nand U19014 (N_19014,N_17239,N_15951);
and U19015 (N_19015,N_14554,N_15985);
and U19016 (N_19016,N_13989,N_15396);
xor U19017 (N_19017,N_15033,N_13285);
nand U19018 (N_19018,N_13437,N_17477);
xor U19019 (N_19019,N_16468,N_13939);
and U19020 (N_19020,N_16088,N_14763);
nand U19021 (N_19021,N_13438,N_13875);
nand U19022 (N_19022,N_14444,N_14911);
or U19023 (N_19023,N_15796,N_12077);
xnor U19024 (N_19024,N_14051,N_16341);
and U19025 (N_19025,N_12230,N_12864);
nand U19026 (N_19026,N_15581,N_12070);
and U19027 (N_19027,N_15189,N_17063);
xnor U19028 (N_19028,N_12381,N_17378);
xnor U19029 (N_19029,N_16661,N_17521);
and U19030 (N_19030,N_17788,N_16252);
nand U19031 (N_19031,N_12099,N_12009);
or U19032 (N_19032,N_17220,N_16538);
nand U19033 (N_19033,N_12396,N_15675);
and U19034 (N_19034,N_14692,N_15832);
nand U19035 (N_19035,N_17530,N_14627);
xnor U19036 (N_19036,N_17943,N_13213);
and U19037 (N_19037,N_14173,N_13705);
or U19038 (N_19038,N_16066,N_13965);
or U19039 (N_19039,N_12757,N_17702);
xor U19040 (N_19040,N_17074,N_13972);
or U19041 (N_19041,N_16793,N_14114);
nor U19042 (N_19042,N_13602,N_15688);
xnor U19043 (N_19043,N_12342,N_16783);
xnor U19044 (N_19044,N_13751,N_13666);
nor U19045 (N_19045,N_15574,N_16797);
nor U19046 (N_19046,N_15661,N_15973);
and U19047 (N_19047,N_14735,N_13212);
xor U19048 (N_19048,N_15231,N_13214);
xnor U19049 (N_19049,N_17425,N_12119);
or U19050 (N_19050,N_14449,N_17481);
nand U19051 (N_19051,N_12586,N_14144);
and U19052 (N_19052,N_13234,N_15593);
nand U19053 (N_19053,N_15887,N_16937);
nand U19054 (N_19054,N_15333,N_17353);
nand U19055 (N_19055,N_13464,N_16102);
or U19056 (N_19056,N_16859,N_14160);
xnor U19057 (N_19057,N_17666,N_15856);
xnor U19058 (N_19058,N_12169,N_14102);
or U19059 (N_19059,N_16310,N_13627);
nand U19060 (N_19060,N_12414,N_14619);
and U19061 (N_19061,N_13890,N_17249);
nor U19062 (N_19062,N_13478,N_16929);
nand U19063 (N_19063,N_14062,N_16114);
xnor U19064 (N_19064,N_15622,N_17347);
and U19065 (N_19065,N_17775,N_13816);
nand U19066 (N_19066,N_17614,N_14293);
or U19067 (N_19067,N_14750,N_15043);
and U19068 (N_19068,N_13612,N_12573);
or U19069 (N_19069,N_14603,N_16981);
or U19070 (N_19070,N_13220,N_16751);
nand U19071 (N_19071,N_15169,N_15965);
and U19072 (N_19072,N_12676,N_13094);
or U19073 (N_19073,N_14651,N_12857);
and U19074 (N_19074,N_14724,N_13900);
xor U19075 (N_19075,N_15515,N_12815);
xnor U19076 (N_19076,N_12531,N_14015);
and U19077 (N_19077,N_17640,N_13659);
xnor U19078 (N_19078,N_16276,N_12534);
nor U19079 (N_19079,N_12368,N_17080);
nand U19080 (N_19080,N_13830,N_12472);
nand U19081 (N_19081,N_12337,N_15011);
and U19082 (N_19082,N_17835,N_14529);
nand U19083 (N_19083,N_14006,N_15341);
nor U19084 (N_19084,N_16754,N_14613);
nand U19085 (N_19085,N_15122,N_12293);
or U19086 (N_19086,N_14073,N_12142);
nor U19087 (N_19087,N_13638,N_15381);
and U19088 (N_19088,N_16288,N_16053);
or U19089 (N_19089,N_13726,N_15885);
nor U19090 (N_19090,N_12369,N_12413);
xor U19091 (N_19091,N_16322,N_16834);
and U19092 (N_19092,N_17067,N_16550);
and U19093 (N_19093,N_16622,N_14481);
or U19094 (N_19094,N_15088,N_17162);
and U19095 (N_19095,N_13668,N_13846);
xnor U19096 (N_19096,N_17500,N_12596);
xor U19097 (N_19097,N_12366,N_15789);
nand U19098 (N_19098,N_13272,N_17172);
and U19099 (N_19099,N_12740,N_15550);
and U19100 (N_19100,N_17176,N_14442);
nor U19101 (N_19101,N_12653,N_13052);
nand U19102 (N_19102,N_14659,N_12193);
or U19103 (N_19103,N_17146,N_15406);
or U19104 (N_19104,N_17052,N_16006);
or U19105 (N_19105,N_13615,N_13817);
nand U19106 (N_19106,N_14803,N_13919);
or U19107 (N_19107,N_15255,N_13414);
nor U19108 (N_19108,N_16381,N_17265);
nand U19109 (N_19109,N_17814,N_15015);
nand U19110 (N_19110,N_12912,N_15598);
or U19111 (N_19111,N_13336,N_12545);
or U19112 (N_19112,N_13368,N_14354);
nand U19113 (N_19113,N_12430,N_14403);
or U19114 (N_19114,N_15075,N_16138);
nor U19115 (N_19115,N_17423,N_12503);
xor U19116 (N_19116,N_14571,N_15283);
xor U19117 (N_19117,N_14372,N_15053);
or U19118 (N_19118,N_14947,N_17405);
nand U19119 (N_19119,N_16702,N_15543);
or U19120 (N_19120,N_16624,N_12223);
or U19121 (N_19121,N_14057,N_16145);
xor U19122 (N_19122,N_12177,N_16463);
nor U19123 (N_19123,N_17123,N_15251);
or U19124 (N_19124,N_12138,N_15564);
or U19125 (N_19125,N_13643,N_13407);
and U19126 (N_19126,N_16021,N_16039);
nand U19127 (N_19127,N_12835,N_14212);
or U19128 (N_19128,N_12330,N_14985);
xor U19129 (N_19129,N_17284,N_17299);
xnor U19130 (N_19130,N_12870,N_13524);
xor U19131 (N_19131,N_13760,N_16519);
xor U19132 (N_19132,N_17773,N_16467);
or U19133 (N_19133,N_15649,N_15506);
xnor U19134 (N_19134,N_14190,N_13952);
and U19135 (N_19135,N_14586,N_17512);
xnor U19136 (N_19136,N_17369,N_16205);
xnor U19137 (N_19137,N_14645,N_13268);
and U19138 (N_19138,N_17654,N_14459);
xnor U19139 (N_19139,N_17738,N_14607);
or U19140 (N_19140,N_15195,N_14591);
nor U19141 (N_19141,N_17950,N_14583);
or U19142 (N_19142,N_17985,N_13147);
and U19143 (N_19143,N_15439,N_13799);
nor U19144 (N_19144,N_12955,N_12061);
xor U19145 (N_19145,N_15380,N_12557);
or U19146 (N_19146,N_17601,N_15289);
nor U19147 (N_19147,N_14711,N_16915);
nor U19148 (N_19148,N_17727,N_16146);
nor U19149 (N_19149,N_13298,N_15848);
xnor U19150 (N_19150,N_17574,N_15241);
nand U19151 (N_19151,N_13527,N_17373);
or U19152 (N_19152,N_16555,N_17945);
and U19153 (N_19153,N_13357,N_15035);
xor U19154 (N_19154,N_12620,N_13400);
or U19155 (N_19155,N_16156,N_15857);
or U19156 (N_19156,N_16290,N_14045);
or U19157 (N_19157,N_13801,N_15925);
and U19158 (N_19158,N_16952,N_17298);
nand U19159 (N_19159,N_14349,N_12704);
nand U19160 (N_19160,N_15934,N_17940);
xnor U19161 (N_19161,N_17565,N_12008);
and U19162 (N_19162,N_17453,N_14461);
and U19163 (N_19163,N_13056,N_17809);
xor U19164 (N_19164,N_14990,N_14732);
and U19165 (N_19165,N_12675,N_12265);
nand U19166 (N_19166,N_14601,N_13020);
nand U19167 (N_19167,N_12526,N_12276);
xor U19168 (N_19168,N_12948,N_13318);
xnor U19169 (N_19169,N_13064,N_14026);
xor U19170 (N_19170,N_15040,N_13170);
and U19171 (N_19171,N_17724,N_16907);
nor U19172 (N_19172,N_14185,N_15814);
nor U19173 (N_19173,N_16001,N_13046);
or U19174 (N_19174,N_12069,N_15104);
nor U19175 (N_19175,N_14514,N_13145);
nand U19176 (N_19176,N_14656,N_17331);
nor U19177 (N_19177,N_17007,N_13096);
and U19178 (N_19178,N_12975,N_14813);
nor U19179 (N_19179,N_15647,N_13980);
nor U19180 (N_19180,N_16972,N_12053);
and U19181 (N_19181,N_15373,N_17164);
or U19182 (N_19182,N_13489,N_13536);
and U19183 (N_19183,N_13366,N_16607);
or U19184 (N_19184,N_16876,N_17971);
nand U19185 (N_19185,N_17831,N_16386);
nor U19186 (N_19186,N_14178,N_13779);
nand U19187 (N_19187,N_14817,N_12552);
or U19188 (N_19188,N_12050,N_16307);
or U19189 (N_19189,N_15785,N_13999);
nand U19190 (N_19190,N_17862,N_14407);
nor U19191 (N_19191,N_15748,N_13525);
xnor U19192 (N_19192,N_13221,N_14077);
and U19193 (N_19193,N_14654,N_12933);
xor U19194 (N_19194,N_15127,N_13863);
nor U19195 (N_19195,N_14210,N_15309);
nand U19196 (N_19196,N_16562,N_17061);
xnor U19197 (N_19197,N_12405,N_14133);
nor U19198 (N_19198,N_13254,N_17957);
nor U19199 (N_19199,N_12504,N_16274);
xnor U19200 (N_19200,N_17443,N_14432);
nand U19201 (N_19201,N_12415,N_12046);
or U19202 (N_19202,N_14100,N_14197);
nor U19203 (N_19203,N_14465,N_16902);
nor U19204 (N_19204,N_13673,N_17679);
or U19205 (N_19205,N_15496,N_17967);
or U19206 (N_19206,N_14958,N_13303);
and U19207 (N_19207,N_14433,N_17489);
nand U19208 (N_19208,N_15402,N_12664);
nor U19209 (N_19209,N_13273,N_13160);
nand U19210 (N_19210,N_15953,N_13388);
nor U19211 (N_19211,N_16096,N_15767);
and U19212 (N_19212,N_16687,N_17905);
nor U19213 (N_19213,N_15952,N_13024);
nand U19214 (N_19214,N_15415,N_15926);
xor U19215 (N_19215,N_13441,N_15305);
and U19216 (N_19216,N_17234,N_13614);
and U19217 (N_19217,N_16621,N_14986);
xor U19218 (N_19218,N_13097,N_15347);
and U19219 (N_19219,N_17304,N_15098);
xor U19220 (N_19220,N_14861,N_12392);
and U19221 (N_19221,N_16496,N_15177);
nor U19222 (N_19222,N_12723,N_17650);
nand U19223 (N_19223,N_16748,N_13113);
xnor U19224 (N_19224,N_12270,N_14880);
nand U19225 (N_19225,N_14726,N_17687);
or U19226 (N_19226,N_16529,N_14110);
and U19227 (N_19227,N_15157,N_12611);
and U19228 (N_19228,N_14362,N_12176);
and U19229 (N_19229,N_17750,N_14098);
and U19230 (N_19230,N_14371,N_14579);
and U19231 (N_19231,N_14605,N_13181);
xnor U19232 (N_19232,N_14657,N_15403);
xnor U19233 (N_19233,N_12269,N_13473);
xnor U19234 (N_19234,N_14468,N_14506);
or U19235 (N_19235,N_17778,N_14072);
nand U19236 (N_19236,N_17930,N_17055);
xnor U19237 (N_19237,N_14632,N_17825);
xor U19238 (N_19238,N_15463,N_15044);
xor U19239 (N_19239,N_12151,N_16350);
and U19240 (N_19240,N_15296,N_15060);
xnor U19241 (N_19241,N_12896,N_15148);
and U19242 (N_19242,N_12243,N_15565);
and U19243 (N_19243,N_16362,N_15321);
xnor U19244 (N_19244,N_13805,N_17897);
xnor U19245 (N_19245,N_16023,N_15690);
nor U19246 (N_19246,N_15431,N_15812);
nor U19247 (N_19247,N_17065,N_13455);
nor U19248 (N_19248,N_14907,N_13196);
nor U19249 (N_19249,N_15151,N_16503);
or U19250 (N_19250,N_16594,N_17542);
xnor U19251 (N_19251,N_16292,N_12018);
and U19252 (N_19252,N_17428,N_16551);
nor U19253 (N_19253,N_16920,N_14996);
nor U19254 (N_19254,N_17167,N_13512);
nand U19255 (N_19255,N_16482,N_14326);
and U19256 (N_19256,N_14345,N_16016);
and U19257 (N_19257,N_13539,N_14139);
or U19258 (N_19258,N_16194,N_12574);
xor U19259 (N_19259,N_16373,N_14714);
nor U19260 (N_19260,N_17602,N_15519);
or U19261 (N_19261,N_12639,N_12382);
xnor U19262 (N_19262,N_12866,N_14843);
nor U19263 (N_19263,N_13309,N_16134);
xnor U19264 (N_19264,N_15829,N_15775);
xnor U19265 (N_19265,N_15989,N_15448);
or U19266 (N_19266,N_15409,N_17626);
and U19267 (N_19267,N_12441,N_15818);
and U19268 (N_19268,N_13912,N_15018);
xnor U19269 (N_19269,N_14436,N_13296);
nand U19270 (N_19270,N_12762,N_13791);
or U19271 (N_19271,N_17184,N_16827);
xor U19272 (N_19272,N_15062,N_14729);
or U19273 (N_19273,N_17044,N_14993);
and U19274 (N_19274,N_15540,N_17482);
nand U19275 (N_19275,N_15911,N_16349);
nand U19276 (N_19276,N_14896,N_15591);
or U19277 (N_19277,N_12567,N_14010);
xnor U19278 (N_19278,N_17682,N_12697);
and U19279 (N_19279,N_12614,N_14337);
or U19280 (N_19280,N_14491,N_12937);
and U19281 (N_19281,N_17802,N_15779);
and U19282 (N_19282,N_17137,N_16187);
or U19283 (N_19283,N_13345,N_17185);
nor U19284 (N_19284,N_14155,N_12869);
nor U19285 (N_19285,N_16928,N_16182);
nand U19286 (N_19286,N_15470,N_13151);
and U19287 (N_19287,N_17812,N_16778);
or U19288 (N_19288,N_15178,N_13456);
or U19289 (N_19289,N_15788,N_12317);
nand U19290 (N_19290,N_13479,N_16013);
or U19291 (N_19291,N_16220,N_12150);
nor U19292 (N_19292,N_13263,N_16646);
nand U19293 (N_19293,N_12166,N_13934);
nand U19294 (N_19294,N_12393,N_13349);
nand U19295 (N_19295,N_17818,N_16881);
xor U19296 (N_19296,N_17909,N_14275);
xor U19297 (N_19297,N_17013,N_16730);
or U19298 (N_19298,N_12942,N_12965);
nand U19299 (N_19299,N_13857,N_12711);
or U19300 (N_19300,N_17984,N_17237);
nor U19301 (N_19301,N_16541,N_16957);
nand U19302 (N_19302,N_13812,N_17255);
xor U19303 (N_19303,N_14543,N_14520);
nor U19304 (N_19304,N_12467,N_14909);
and U19305 (N_19305,N_15568,N_12772);
or U19306 (N_19306,N_14978,N_13874);
or U19307 (N_19307,N_13510,N_16000);
or U19308 (N_19308,N_17333,N_16668);
nor U19309 (N_19309,N_15259,N_15232);
and U19310 (N_19310,N_17722,N_16408);
and U19311 (N_19311,N_16235,N_16100);
nor U19312 (N_19312,N_12494,N_14906);
and U19313 (N_19313,N_12348,N_12025);
and U19314 (N_19314,N_12980,N_17228);
xor U19315 (N_19315,N_14617,N_13372);
or U19316 (N_19316,N_16003,N_13688);
or U19317 (N_19317,N_14552,N_13183);
nor U19318 (N_19318,N_16323,N_15621);
xnor U19319 (N_19319,N_16804,N_14590);
and U19320 (N_19320,N_17206,N_14324);
or U19321 (N_19321,N_13051,N_12856);
and U19322 (N_19322,N_13486,N_13730);
xor U19323 (N_19323,N_12408,N_12824);
xor U19324 (N_19324,N_17846,N_14254);
nor U19325 (N_19325,N_12998,N_12089);
nor U19326 (N_19326,N_17107,N_16325);
and U19327 (N_19327,N_16822,N_17152);
xor U19328 (N_19328,N_13915,N_16671);
nor U19329 (N_19329,N_12535,N_16520);
nor U19330 (N_19330,N_14614,N_15626);
and U19331 (N_19331,N_13802,N_14881);
nand U19332 (N_19332,N_17250,N_14470);
xor U19333 (N_19333,N_17791,N_13111);
xnor U19334 (N_19334,N_13901,N_13108);
nor U19335 (N_19335,N_13654,N_16324);
xor U19336 (N_19336,N_12041,N_16480);
nor U19337 (N_19337,N_17315,N_17344);
or U19338 (N_19338,N_16017,N_17784);
xnor U19339 (N_19339,N_12585,N_13048);
nor U19340 (N_19340,N_17174,N_13465);
and U19341 (N_19341,N_17887,N_12992);
nand U19342 (N_19342,N_12575,N_17356);
or U19343 (N_19343,N_12371,N_12692);
nor U19344 (N_19344,N_17038,N_16769);
nand U19345 (N_19345,N_13690,N_14176);
and U19346 (N_19346,N_15079,N_15513);
nor U19347 (N_19347,N_14244,N_12728);
or U19348 (N_19348,N_13582,N_17085);
or U19349 (N_19349,N_16444,N_17455);
nand U19350 (N_19350,N_13130,N_16836);
xnor U19351 (N_19351,N_14359,N_17786);
xnor U19352 (N_19352,N_17509,N_15272);
nor U19353 (N_19353,N_13301,N_12336);
nand U19354 (N_19354,N_16986,N_14487);
or U19355 (N_19355,N_17059,N_17757);
nor U19356 (N_19356,N_17595,N_12228);
and U19357 (N_19357,N_14205,N_15430);
nand U19358 (N_19358,N_17472,N_17183);
and U19359 (N_19359,N_13671,N_14036);
or U19360 (N_19360,N_15013,N_17588);
nor U19361 (N_19361,N_16965,N_16897);
xor U19362 (N_19362,N_17535,N_17699);
xnor U19363 (N_19363,N_17330,N_15907);
nand U19364 (N_19364,N_14955,N_14404);
nor U19365 (N_19365,N_15978,N_17524);
xor U19366 (N_19366,N_15531,N_12116);
nand U19367 (N_19367,N_13725,N_13758);
xor U19368 (N_19368,N_17637,N_13283);
and U19369 (N_19369,N_13828,N_16409);
nand U19370 (N_19370,N_16062,N_17232);
xor U19371 (N_19371,N_15670,N_16643);
xnor U19372 (N_19372,N_15813,N_15731);
nand U19373 (N_19373,N_12161,N_12326);
xor U19374 (N_19374,N_17035,N_16335);
and U19375 (N_19375,N_14675,N_16700);
and U19376 (N_19376,N_15389,N_14845);
and U19377 (N_19377,N_17251,N_14517);
xor U19378 (N_19378,N_13379,N_17293);
nor U19379 (N_19379,N_12235,N_12577);
xnor U19380 (N_19380,N_14338,N_14954);
nand U19381 (N_19381,N_14179,N_12825);
nor U19382 (N_19382,N_12682,N_13622);
xnor U19383 (N_19383,N_12588,N_15080);
xor U19384 (N_19384,N_15394,N_17625);
or U19385 (N_19385,N_17681,N_13477);
nor U19386 (N_19386,N_12104,N_16824);
xnor U19387 (N_19387,N_12860,N_14189);
and U19388 (N_19388,N_17308,N_16684);
nor U19389 (N_19389,N_16932,N_14335);
and U19390 (N_19390,N_13560,N_13378);
xor U19391 (N_19391,N_15903,N_17927);
nand U19392 (N_19392,N_17056,N_12903);
nor U19393 (N_19393,N_13955,N_17544);
and U19394 (N_19394,N_14104,N_15600);
or U19395 (N_19395,N_12722,N_13977);
nor U19396 (N_19396,N_12372,N_12423);
nor U19397 (N_19397,N_15532,N_13844);
or U19398 (N_19398,N_14809,N_17178);
and U19399 (N_19399,N_15722,N_13133);
and U19400 (N_19400,N_16414,N_17647);
or U19401 (N_19401,N_16140,N_17003);
nand U19402 (N_19402,N_13833,N_13155);
or U19403 (N_19403,N_14216,N_15466);
nand U19404 (N_19404,N_13115,N_15697);
and U19405 (N_19405,N_17946,N_14829);
nand U19406 (N_19406,N_17955,N_17755);
nand U19407 (N_19407,N_16573,N_15003);
nor U19408 (N_19408,N_13119,N_14783);
xor U19409 (N_19409,N_14217,N_13117);
or U19410 (N_19410,N_17822,N_16351);
and U19411 (N_19411,N_13839,N_16557);
nor U19412 (N_19412,N_17314,N_13948);
xor U19413 (N_19413,N_16340,N_16097);
and U19414 (N_19414,N_13694,N_14594);
nand U19415 (N_19415,N_15998,N_17516);
nand U19416 (N_19416,N_17826,N_16151);
xor U19417 (N_19417,N_13240,N_16919);
nor U19418 (N_19418,N_13861,N_14317);
nor U19419 (N_19419,N_16877,N_15963);
and U19420 (N_19420,N_13604,N_14642);
xor U19421 (N_19421,N_15556,N_17431);
xor U19422 (N_19422,N_13084,N_16082);
nand U19423 (N_19423,N_14003,N_13124);
nor U19424 (N_19424,N_17393,N_12167);
or U19425 (N_19425,N_13740,N_12592);
or U19426 (N_19426,N_14649,N_14580);
and U19427 (N_19427,N_17303,N_13330);
or U19428 (N_19428,N_12221,N_13595);
or U19429 (N_19429,N_15058,N_16457);
xnor U19430 (N_19430,N_16278,N_14127);
nor U19431 (N_19431,N_14424,N_14946);
nor U19432 (N_19432,N_14931,N_12486);
and U19433 (N_19433,N_14561,N_16933);
and U19434 (N_19434,N_13552,N_13821);
nand U19435 (N_19435,N_14425,N_16363);
nand U19436 (N_19436,N_14992,N_15726);
or U19437 (N_19437,N_15941,N_17149);
xor U19438 (N_19438,N_13722,N_14643);
nor U19439 (N_19439,N_12134,N_15768);
nand U19440 (N_19440,N_13993,N_13440);
nor U19441 (N_19441,N_17462,N_14365);
xnor U19442 (N_19442,N_12982,N_15783);
or U19443 (N_19443,N_16107,N_12547);
nand U19444 (N_19444,N_15112,N_13797);
nor U19445 (N_19445,N_17072,N_13132);
or U19446 (N_19446,N_16139,N_12446);
nand U19447 (N_19447,N_15546,N_14128);
xor U19448 (N_19448,N_17685,N_14838);
and U19449 (N_19449,N_17186,N_14792);
or U19450 (N_19450,N_14325,N_15386);
nand U19451 (N_19451,N_17903,N_12445);
or U19452 (N_19452,N_13009,N_17697);
nor U19453 (N_19453,N_15376,N_13025);
or U19454 (N_19454,N_12706,N_15671);
or U19455 (N_19455,N_13935,N_16811);
nor U19456 (N_19456,N_15124,N_15176);
nand U19457 (N_19457,N_12171,N_14719);
or U19458 (N_19458,N_16272,N_13594);
or U19459 (N_19459,N_13194,N_12067);
and U19460 (N_19460,N_16331,N_13416);
nand U19461 (N_19461,N_17966,N_17580);
or U19462 (N_19462,N_16889,N_13911);
or U19463 (N_19463,N_12595,N_13970);
or U19464 (N_19464,N_17891,N_12964);
and U19465 (N_19465,N_17305,N_17380);
nor U19466 (N_19466,N_15747,N_14866);
or U19467 (N_19467,N_13624,N_14132);
or U19468 (N_19468,N_14136,N_14471);
nand U19469 (N_19469,N_16631,N_12453);
or U19470 (N_19470,N_16499,N_17736);
xnor U19471 (N_19471,N_17754,N_13433);
nand U19472 (N_19472,N_13596,N_14935);
or U19473 (N_19473,N_15006,N_13348);
or U19474 (N_19474,N_15918,N_15358);
nor U19475 (N_19475,N_13102,N_14725);
xnor U19476 (N_19476,N_16864,N_12525);
and U19477 (N_19477,N_16537,N_14450);
nand U19478 (N_19478,N_15498,N_15874);
xor U19479 (N_19479,N_14887,N_17410);
and U19480 (N_19480,N_16185,N_13752);
nor U19481 (N_19481,N_14489,N_14640);
nor U19482 (N_19482,N_15046,N_12199);
xor U19483 (N_19483,N_13322,N_16695);
nor U19484 (N_19484,N_17526,N_12972);
nor U19485 (N_19485,N_15150,N_15499);
and U19486 (N_19486,N_13463,N_17569);
nand U19487 (N_19487,N_16608,N_17508);
nand U19488 (N_19488,N_17361,N_17603);
or U19489 (N_19489,N_13395,N_13038);
and U19490 (N_19490,N_17483,N_13815);
nor U19491 (N_19491,N_14005,N_15847);
xnor U19492 (N_19492,N_17236,N_16759);
xnor U19493 (N_19493,N_12033,N_17048);
nor U19494 (N_19494,N_14758,N_16531);
nor U19495 (N_19495,N_13569,N_17224);
or U19496 (N_19496,N_12349,N_15143);
and U19497 (N_19497,N_14693,N_17199);
xnor U19498 (N_19498,N_17324,N_15149);
xor U19499 (N_19499,N_13275,N_15816);
nand U19500 (N_19500,N_16934,N_14684);
and U19501 (N_19501,N_14548,N_12483);
xnor U19502 (N_19502,N_14712,N_17622);
and U19503 (N_19503,N_14202,N_12612);
nand U19504 (N_19504,N_15250,N_13312);
nor U19505 (N_19505,N_15184,N_16850);
nor U19506 (N_19506,N_17473,N_17457);
nand U19507 (N_19507,N_17525,N_12078);
nand U19508 (N_19508,N_12442,N_12356);
and U19509 (N_19509,N_12681,N_15894);
and U19510 (N_19510,N_16399,N_16917);
nor U19511 (N_19511,N_16984,N_13974);
nand U19512 (N_19512,N_15566,N_15579);
xor U19513 (N_19513,N_14285,N_15603);
xor U19514 (N_19514,N_12272,N_13152);
xnor U19515 (N_19515,N_17889,N_13403);
xor U19516 (N_19516,N_17870,N_14291);
or U19517 (N_19517,N_13460,N_14078);
nand U19518 (N_19518,N_12572,N_13063);
xor U19519 (N_19519,N_12157,N_15266);
xnor U19520 (N_19520,N_12537,N_16506);
or U19521 (N_19521,N_13548,N_17011);
and U19522 (N_19522,N_15392,N_14245);
nor U19523 (N_19523,N_16035,N_13516);
xnor U19524 (N_19524,N_14876,N_13990);
nand U19525 (N_19525,N_12255,N_13686);
nor U19526 (N_19526,N_17609,N_16518);
or U19527 (N_19527,N_16923,N_17656);
nand U19528 (N_19528,N_15096,N_13633);
xor U19529 (N_19529,N_16963,N_15893);
nor U19530 (N_19530,N_13807,N_13580);
nor U19531 (N_19531,N_16122,N_16791);
nand U19532 (N_19532,N_15235,N_13590);
and U19533 (N_19533,N_17752,N_13898);
nor U19534 (N_19534,N_17209,N_17094);
or U19535 (N_19535,N_16103,N_16456);
nor U19536 (N_19536,N_14184,N_17813);
or U19537 (N_19537,N_15436,N_12085);
or U19538 (N_19538,N_15969,N_14061);
or U19539 (N_19539,N_17801,N_15630);
nand U19540 (N_19540,N_12935,N_16504);
nor U19541 (N_19541,N_14505,N_12501);
and U19542 (N_19542,N_13573,N_13945);
xnor U19543 (N_19543,N_16857,N_13281);
nor U19544 (N_19544,N_13100,N_15528);
nor U19545 (N_19545,N_12254,N_14756);
or U19546 (N_19546,N_16109,N_14271);
and U19547 (N_19547,N_16170,N_14558);
and U19548 (N_19548,N_13558,N_17188);
and U19549 (N_19549,N_15790,N_12542);
and U19550 (N_19550,N_12977,N_14578);
nand U19551 (N_19551,N_13461,N_12973);
xor U19552 (N_19552,N_14660,N_13299);
nor U19553 (N_19553,N_15310,N_13317);
xor U19554 (N_19554,N_15699,N_14777);
nor U19555 (N_19555,N_13218,N_14519);
and U19556 (N_19556,N_17873,N_16211);
nand U19557 (N_19557,N_12895,N_16526);
xor U19558 (N_19558,N_16861,N_12920);
or U19559 (N_19559,N_13393,N_16711);
xnor U19560 (N_19560,N_14177,N_17969);
and U19561 (N_19561,N_16899,N_14391);
xnor U19562 (N_19562,N_17926,N_13210);
and U19563 (N_19563,N_17242,N_16233);
nor U19564 (N_19564,N_12801,N_12347);
or U19565 (N_19565,N_16841,N_13005);
and U19566 (N_19566,N_15563,N_13424);
xnor U19567 (N_19567,N_16250,N_15784);
nand U19568 (N_19568,N_15668,N_16742);
and U19569 (N_19569,N_13913,N_17112);
and U19570 (N_19570,N_13937,N_14397);
and U19571 (N_19571,N_14009,N_14351);
and U19572 (N_19572,N_12530,N_12687);
xor U19573 (N_19573,N_13665,N_14394);
or U19574 (N_19574,N_12710,N_12062);
or U19575 (N_19575,N_17892,N_17229);
or U19576 (N_19576,N_17765,N_15087);
xnor U19577 (N_19577,N_15886,N_16357);
xor U19578 (N_19578,N_12993,N_16471);
xnor U19579 (N_19579,N_12031,N_15328);
nand U19580 (N_19580,N_14166,N_17604);
and U19581 (N_19581,N_17068,N_17740);
nor U19582 (N_19582,N_13382,N_15293);
nand U19583 (N_19583,N_15777,N_13126);
nor U19584 (N_19584,N_13162,N_12899);
nand U19585 (N_19585,N_12037,N_16389);
xnor U19586 (N_19586,N_12662,N_17952);
or U19587 (N_19587,N_15275,N_15940);
nor U19588 (N_19588,N_15465,N_14111);
nand U19589 (N_19589,N_12395,N_12058);
or U19590 (N_19590,N_13114,N_17189);
nor U19591 (N_19591,N_14988,N_13592);
nor U19592 (N_19592,N_16543,N_14680);
nor U19593 (N_19593,N_13105,N_13252);
nand U19594 (N_19594,N_16106,N_13340);
nand U19595 (N_19595,N_13313,N_12005);
or U19596 (N_19596,N_17593,N_13390);
and U19597 (N_19597,N_16469,N_16237);
xor U19598 (N_19598,N_17212,N_17528);
xor U19599 (N_19599,N_12383,N_13342);
xnor U19600 (N_19600,N_16101,N_15267);
nor U19601 (N_19601,N_12717,N_15750);
nor U19602 (N_19602,N_14106,N_14577);
nand U19603 (N_19603,N_13139,N_15509);
nor U19604 (N_19604,N_16690,N_16345);
xor U19605 (N_19605,N_17662,N_12563);
nor U19606 (N_19606,N_14211,N_14716);
nor U19607 (N_19607,N_12130,N_12881);
or U19608 (N_19608,N_16539,N_17829);
xnor U19609 (N_19609,N_15170,N_16685);
nor U19610 (N_19610,N_13019,N_16939);
or U19611 (N_19611,N_16317,N_16694);
and U19612 (N_19612,N_14901,N_15495);
or U19613 (N_19613,N_13775,N_13088);
xnor U19614 (N_19614,N_16849,N_15725);
or U19615 (N_19615,N_12344,N_12853);
nor U19616 (N_19616,N_15962,N_14550);
nor U19617 (N_19617,N_13409,N_13371);
nand U19618 (N_19618,N_17464,N_16763);
xor U19619 (N_19619,N_15086,N_17864);
or U19620 (N_19620,N_12546,N_17427);
nor U19621 (N_19621,N_14741,N_13011);
or U19622 (N_19622,N_14417,N_13125);
nand U19623 (N_19623,N_16926,N_12264);
and U19624 (N_19624,N_16478,N_13000);
and U19625 (N_19625,N_16664,N_12837);
nand U19626 (N_19626,N_12362,N_13229);
and U19627 (N_19627,N_12997,N_13769);
nor U19628 (N_19628,N_16625,N_13601);
or U19629 (N_19629,N_16925,N_17254);
nand U19630 (N_19630,N_12677,N_17531);
xnor U19631 (N_19631,N_15437,N_15739);
nand U19632 (N_19632,N_15049,N_14377);
and U19633 (N_19633,N_16829,N_14188);
nand U19634 (N_19634,N_13664,N_17288);
nand U19635 (N_19635,N_14828,N_16275);
nor U19636 (N_19636,N_15179,N_15648);
nor U19637 (N_19637,N_17980,N_13881);
nor U19638 (N_19638,N_12660,N_15372);
xnor U19639 (N_19639,N_15772,N_13137);
xnor U19640 (N_19640,N_13869,N_15128);
xnor U19641 (N_19641,N_15001,N_15244);
nor U19642 (N_19642,N_14898,N_14370);
xnor U19643 (N_19643,N_12374,N_12341);
nand U19644 (N_19644,N_12775,N_17180);
nand U19645 (N_19645,N_13662,N_16657);
or U19646 (N_19646,N_12029,N_15782);
or U19647 (N_19647,N_13062,N_12377);
nand U19648 (N_19648,N_15337,N_17051);
xnor U19649 (N_19649,N_17321,N_13469);
nor U19650 (N_19650,N_15411,N_13154);
or U19651 (N_19651,N_16566,N_15803);
or U19652 (N_19652,N_17145,N_17855);
nand U19653 (N_19653,N_14207,N_12183);
or U19654 (N_19654,N_17230,N_12764);
nand U19655 (N_19655,N_17981,N_12850);
nor U19656 (N_19656,N_14934,N_15586);
xnor U19657 (N_19657,N_14629,N_16126);
and U19658 (N_19658,N_13651,N_14582);
or U19659 (N_19659,N_12540,N_14628);
and U19660 (N_19660,N_15336,N_17195);
and U19661 (N_19661,N_13991,N_13682);
xor U19662 (N_19662,N_15551,N_14447);
and U19663 (N_19663,N_12522,N_15005);
and U19664 (N_19664,N_14611,N_14192);
nor U19665 (N_19665,N_14069,N_12375);
and U19666 (N_19666,N_13540,N_17130);
nand U19667 (N_19667,N_14226,N_16230);
and U19668 (N_19668,N_12125,N_15837);
xnor U19669 (N_19669,N_16081,N_15617);
and U19670 (N_19670,N_14181,N_12726);
or U19671 (N_19671,N_13852,N_12497);
nor U19672 (N_19672,N_16491,N_13127);
nor U19673 (N_19673,N_14760,N_16328);
nand U19674 (N_19674,N_12926,N_14872);
xnor U19675 (N_19675,N_15243,N_17578);
nand U19676 (N_19676,N_12752,N_17115);
or U19677 (N_19677,N_15067,N_14152);
nor U19678 (N_19678,N_17327,N_14853);
nor U19679 (N_19679,N_13231,N_15004);
and U19680 (N_19680,N_12967,N_17322);
nor U19681 (N_19681,N_15629,N_13744);
nor U19682 (N_19682,N_12132,N_12604);
nand U19683 (N_19683,N_17179,N_12988);
and U19684 (N_19684,N_17556,N_17306);
and U19685 (N_19685,N_17878,N_12490);
and U19686 (N_19686,N_15481,N_17415);
and U19687 (N_19687,N_14570,N_17686);
or U19688 (N_19688,N_17416,N_12282);
nand U19689 (N_19689,N_14153,N_13892);
and U19690 (N_19690,N_12127,N_16497);
or U19691 (N_19691,N_14375,N_16856);
nor U19692 (N_19692,N_15378,N_17175);
xnor U19693 (N_19693,N_12602,N_16076);
xnor U19694 (N_19694,N_16040,N_14137);
or U19695 (N_19695,N_12771,N_16840);
nand U19696 (N_19696,N_14199,N_14124);
nor U19697 (N_19697,N_16747,N_14278);
nand U19698 (N_19698,N_17636,N_15065);
xor U19699 (N_19699,N_12214,N_14369);
nor U19700 (N_19700,N_14648,N_14419);
nor U19701 (N_19701,N_16378,N_14687);
or U19702 (N_19702,N_16707,N_17422);
and U19703 (N_19703,N_12727,N_16279);
nand U19704 (N_19704,N_15366,N_12868);
nand U19705 (N_19705,N_16254,N_17348);
and U19706 (N_19706,N_15753,N_12464);
nand U19707 (N_19707,N_14058,N_13310);
nand U19708 (N_19708,N_14208,N_13549);
and U19709 (N_19709,N_17452,N_17078);
nand U19710 (N_19710,N_12768,N_13747);
or U19711 (N_19711,N_14174,N_12456);
or U19712 (N_19712,N_13672,N_13529);
nand U19713 (N_19713,N_17629,N_12603);
nand U19714 (N_19714,N_15787,N_13940);
nand U19715 (N_19715,N_16033,N_15851);
or U19716 (N_19716,N_15827,N_16647);
and U19717 (N_19717,N_14498,N_14769);
and U19718 (N_19718,N_13713,N_14260);
and U19719 (N_19719,N_12364,N_15745);
and U19720 (N_19720,N_12641,N_14546);
nand U19721 (N_19721,N_13199,N_13453);
xnor U19722 (N_19722,N_16892,N_16994);
nand U19723 (N_19723,N_17043,N_13531);
nand U19724 (N_19724,N_14926,N_17487);
or U19725 (N_19725,N_12854,N_15682);
nand U19726 (N_19726,N_14270,N_16693);
xor U19727 (N_19727,N_16715,N_17947);
xnor U19728 (N_19728,N_16206,N_17365);
nor U19729 (N_19729,N_16931,N_17026);
and U19730 (N_19730,N_14042,N_12215);
or U19731 (N_19731,N_17806,N_15281);
or U19732 (N_19732,N_17768,N_12121);
or U19733 (N_19733,N_15224,N_17583);
nand U19734 (N_19734,N_14553,N_15971);
xor U19735 (N_19735,N_13781,N_12558);
nand U19736 (N_19736,N_12657,N_15650);
and U19737 (N_19737,N_13675,N_17975);
nand U19738 (N_19738,N_14888,N_15278);
nor U19739 (N_19739,N_16815,N_14592);
nor U19740 (N_19740,N_14000,N_12287);
and U19741 (N_19741,N_13343,N_14748);
or U19742 (N_19742,N_13932,N_17646);
or U19743 (N_19743,N_15227,N_15651);
and U19744 (N_19744,N_17635,N_17337);
nand U19745 (N_19745,N_13351,N_16382);
nor U19746 (N_19746,N_12186,N_13770);
nand U19747 (N_19747,N_15085,N_17728);
xnor U19748 (N_19748,N_13591,N_16628);
nor U19749 (N_19749,N_13820,N_15363);
or U19750 (N_19750,N_13851,N_13017);
xnor U19751 (N_19751,N_13777,N_17645);
nor U19752 (N_19752,N_17538,N_15442);
or U19753 (N_19753,N_15326,N_17513);
nand U19754 (N_19754,N_16852,N_14593);
xnor U19755 (N_19755,N_16680,N_14959);
and U19756 (N_19756,N_16178,N_15213);
xnor U19757 (N_19757,N_16355,N_14545);
xnor U19758 (N_19758,N_16614,N_17261);
or U19759 (N_19759,N_13216,N_12963);
xor U19760 (N_19760,N_12890,N_15472);
and U19761 (N_19761,N_13684,N_17016);
and U19762 (N_19762,N_16011,N_17726);
nand U19763 (N_19763,N_15741,N_12914);
xnor U19764 (N_19764,N_16673,N_14482);
xnor U19765 (N_19765,N_14759,N_13323);
and U19766 (N_19766,N_14994,N_16200);
xnor U19767 (N_19767,N_17616,N_16287);
and U19768 (N_19768,N_12769,N_12194);
xnor U19769 (N_19769,N_16052,N_16376);
and U19770 (N_19770,N_16989,N_12873);
nand U19771 (N_19771,N_13988,N_12418);
nand U19772 (N_19772,N_17019,N_12820);
nand U19773 (N_19773,N_17976,N_17279);
nand U19774 (N_19774,N_13219,N_14559);
nor U19775 (N_19775,N_12985,N_15108);
or U19776 (N_19776,N_15710,N_17610);
or U19777 (N_19777,N_15576,N_13589);
nand U19778 (N_19778,N_16768,N_16370);
or U19779 (N_19779,N_17095,N_15294);
xor U19780 (N_19780,N_14982,N_14535);
and U19781 (N_19781,N_12562,N_12279);
nand U19782 (N_19782,N_15514,N_16511);
or U19783 (N_19783,N_12510,N_12457);
or U19784 (N_19784,N_12217,N_17924);
xnor U19785 (N_19785,N_17379,N_15214);
nor U19786 (N_19786,N_16299,N_17623);
nand U19787 (N_19787,N_14513,N_16716);
xnor U19788 (N_19788,N_16616,N_13838);
xor U19789 (N_19789,N_14766,N_16367);
nor U19790 (N_19790,N_16998,N_13121);
and U19791 (N_19791,N_15320,N_12158);
or U19792 (N_19792,N_16090,N_16794);
nor U19793 (N_19793,N_16486,N_16833);
xor U19794 (N_19794,N_12874,N_17882);
xnor U19795 (N_19795,N_13691,N_12690);
nand U19796 (N_19796,N_12076,N_12488);
nand U19797 (N_19797,N_12248,N_16839);
and U19798 (N_19798,N_14771,N_17536);
nand U19799 (N_19799,N_14413,N_14837);
and U19800 (N_19800,N_13864,N_13842);
or U19801 (N_19801,N_15097,N_14972);
nor U19802 (N_19802,N_14796,N_17954);
nor U19803 (N_19803,N_17585,N_13818);
and U19804 (N_19804,N_12307,N_14544);
nor U19805 (N_19805,N_16597,N_12517);
nand U19806 (N_19806,N_15706,N_15028);
nand U19807 (N_19807,N_15666,N_14965);
nor U19808 (N_19808,N_15071,N_17739);
nor U19809 (N_19809,N_12819,N_14819);
and U19810 (N_19810,N_17992,N_15809);
nor U19811 (N_19811,N_13077,N_14623);
nor U19812 (N_19812,N_16990,N_14757);
or U19813 (N_19813,N_12983,N_17692);
and U19814 (N_19814,N_16067,N_17990);
and U19815 (N_19815,N_17839,N_15443);
xnor U19816 (N_19816,N_15693,N_12688);
nor U19817 (N_19817,N_15385,N_16732);
nor U19818 (N_19818,N_16459,N_15084);
or U19819 (N_19819,N_15365,N_16372);
xnor U19820 (N_19820,N_17928,N_17689);
nand U19821 (N_19821,N_15982,N_16801);
xor U19822 (N_19822,N_17570,N_16311);
nand U19823 (N_19823,N_15469,N_13010);
nor U19824 (N_19824,N_17547,N_12357);
or U19825 (N_19825,N_13641,N_12471);
nand U19826 (N_19826,N_13485,N_12315);
and U19827 (N_19827,N_17023,N_12370);
nand U19828 (N_19828,N_13750,N_16582);
or U19829 (N_19829,N_17342,N_12410);
nand U19830 (N_19830,N_12097,N_15123);
nand U19831 (N_19831,N_15357,N_15610);
and U19832 (N_19832,N_17991,N_14863);
xor U19833 (N_19833,N_14040,N_15163);
nor U19834 (N_19834,N_13858,N_17511);
nand U19835 (N_19835,N_15010,N_14501);
nand U19836 (N_19836,N_17388,N_17022);
or U19837 (N_19837,N_14280,N_14525);
nor U19838 (N_19838,N_16071,N_17958);
or U19839 (N_19839,N_16204,N_13893);
and U19840 (N_19840,N_17731,N_16681);
and U19841 (N_19841,N_13205,N_12152);
nand U19842 (N_19842,N_16927,N_15606);
nor U19843 (N_19843,N_13723,N_15487);
nand U19844 (N_19844,N_17611,N_15815);
nand U19845 (N_19845,N_15643,N_14230);
and U19846 (N_19846,N_12258,N_15034);
or U19847 (N_19847,N_15102,N_13581);
xor U19848 (N_19848,N_15527,N_15130);
xor U19849 (N_19849,N_14315,N_12238);
and U19850 (N_19850,N_14378,N_13905);
nor U19851 (N_19851,N_15632,N_15352);
nor U19852 (N_19852,N_14927,N_14499);
nand U19853 (N_19853,N_13023,N_14621);
and U19854 (N_19854,N_13241,N_12107);
nand U19855 (N_19855,N_16563,N_13808);
or U19856 (N_19856,N_17099,N_14079);
nor U19857 (N_19857,N_16396,N_16667);
and U19858 (N_19858,N_15582,N_17214);
and U19859 (N_19859,N_15497,N_13634);
xnor U19860 (N_19860,N_12427,N_13314);
and U19861 (N_19861,N_16584,N_13176);
nand U19862 (N_19862,N_12591,N_16773);
xor U19863 (N_19863,N_17779,N_17863);
xnor U19864 (N_19864,N_17712,N_17225);
nand U19865 (N_19865,N_17534,N_15742);
nand U19866 (N_19866,N_16598,N_15057);
or U19867 (N_19867,N_16589,N_16212);
nor U19868 (N_19868,N_16679,N_15521);
or U19869 (N_19869,N_13289,N_13754);
nand U19870 (N_19870,N_12048,N_12484);
or U19871 (N_19871,N_12136,N_17621);
and U19872 (N_19872,N_16298,N_14175);
xnor U19873 (N_19873,N_13384,N_15008);
xnor U19874 (N_19874,N_12409,N_16828);
and U19875 (N_19875,N_13635,N_15173);
nor U19876 (N_19876,N_12951,N_13008);
nand U19877 (N_19877,N_17111,N_16916);
nor U19878 (N_19878,N_15198,N_16450);
or U19879 (N_19879,N_12428,N_16009);
nor U19880 (N_19880,N_12593,N_13352);
xnor U19881 (N_19881,N_15175,N_14751);
nand U19882 (N_19882,N_12092,N_16135);
xnor U19883 (N_19883,N_13239,N_15229);
nor U19884 (N_19884,N_16724,N_12355);
and U19885 (N_19885,N_12429,N_16805);
nor U19886 (N_19886,N_14921,N_12252);
nand U19887 (N_19887,N_16443,N_16516);
xnor U19888 (N_19888,N_17420,N_14620);
xnor U19889 (N_19889,N_14682,N_13565);
nand U19890 (N_19890,N_12081,N_13514);
or U19891 (N_19891,N_12475,N_14274);
nand U19892 (N_19892,N_15936,N_14088);
nor U19893 (N_19893,N_12088,N_12636);
nor U19894 (N_19894,N_17064,N_16155);
nand U19895 (N_19895,N_12000,N_16996);
nand U19896 (N_19896,N_13361,N_16417);
nor U19897 (N_19897,N_17401,N_12543);
xor U19898 (N_19898,N_17606,N_15286);
xor U19899 (N_19899,N_12003,N_17615);
or U19900 (N_19900,N_15845,N_14779);
xnor U19901 (N_19901,N_16788,N_16942);
or U19902 (N_19902,N_17444,N_14983);
nand U19903 (N_19903,N_17937,N_15480);
xor U19904 (N_19904,N_16481,N_15056);
xor U19905 (N_19905,N_13759,N_13909);
nand U19906 (N_19906,N_13885,N_16776);
and U19907 (N_19907,N_14292,N_13658);
or U19908 (N_19908,N_13987,N_15399);
or U19909 (N_19909,N_13584,N_12634);
and U19910 (N_19910,N_13532,N_14235);
nand U19911 (N_19911,N_16613,N_15230);
nand U19912 (N_19912,N_13277,N_17392);
xnor U19913 (N_19913,N_13200,N_15729);
nor U19914 (N_19914,N_12032,N_13889);
xnor U19915 (N_19915,N_17680,N_17854);
nand U19916 (N_19916,N_14943,N_16057);
and U19917 (N_19917,N_16344,N_16709);
and U19918 (N_19918,N_14252,N_15811);
or U19919 (N_19919,N_15207,N_16686);
xor U19920 (N_19920,N_13888,N_17627);
nor U19921 (N_19921,N_13767,N_17158);
nor U19922 (N_19922,N_16796,N_12756);
and U19923 (N_19923,N_15340,N_17515);
and U19924 (N_19924,N_12426,N_16129);
xor U19925 (N_19925,N_16626,N_17190);
xor U19926 (N_19926,N_12550,N_15304);
nand U19927 (N_19927,N_13519,N_15324);
nand U19928 (N_19928,N_15922,N_15672);
nand U19929 (N_19929,N_17471,N_14807);
or U19930 (N_19930,N_13502,N_15696);
nand U19931 (N_19931,N_14780,N_17262);
xnor U19932 (N_19932,N_13587,N_15174);
xnor U19933 (N_19933,N_13556,N_12892);
nor U19934 (N_19934,N_13515,N_12292);
or U19935 (N_19935,N_14364,N_17564);
xnor U19936 (N_19936,N_13951,N_16808);
xor U19937 (N_19937,N_12923,N_16093);
and U19938 (N_19938,N_14704,N_13044);
and U19939 (N_19939,N_12732,N_12433);
xor U19940 (N_19940,N_16846,N_17396);
nand U19941 (N_19941,N_15152,N_12953);
nor U19942 (N_19942,N_16222,N_17834);
or U19943 (N_19943,N_17653,N_15511);
and U19944 (N_19944,N_12748,N_12695);
and U19945 (N_19945,N_15050,N_12674);
nor U19946 (N_19946,N_12613,N_15082);
or U19947 (N_19947,N_16069,N_14539);
nand U19948 (N_19948,N_13197,N_17514);
or U19949 (N_19949,N_13541,N_12544);
xnor U19950 (N_19950,N_15711,N_12283);
and U19951 (N_19951,N_12583,N_16609);
nor U19952 (N_19952,N_16371,N_15319);
nand U19953 (N_19953,N_17644,N_12224);
or U19954 (N_19954,N_15867,N_17983);
xor U19955 (N_19955,N_17098,N_15658);
and U19956 (N_19956,N_14213,N_16243);
nand U19957 (N_19957,N_14884,N_17108);
or U19958 (N_19958,N_13377,N_17287);
xnor U19959 (N_19959,N_13593,N_12459);
or U19960 (N_19960,N_13506,N_17491);
nor U19961 (N_19961,N_16113,N_12944);
and U19962 (N_19962,N_17267,N_13856);
nand U19963 (N_19963,N_16203,N_17437);
or U19964 (N_19964,N_13876,N_13344);
nand U19965 (N_19965,N_16483,N_12310);
nor U19966 (N_19966,N_14138,N_15434);
or U19967 (N_19967,N_13087,N_12294);
nand U19968 (N_19968,N_13138,N_12673);
or U19969 (N_19969,N_14980,N_15974);
nand U19970 (N_19970,N_16285,N_12098);
or U19971 (N_19971,N_13674,N_16038);
xnor U19972 (N_19972,N_12994,N_13773);
nor U19973 (N_19973,N_13792,N_15462);
nand U19974 (N_19974,N_16909,N_13260);
nor U19975 (N_19975,N_14439,N_17540);
xor U19976 (N_19976,N_13385,N_12852);
or U19977 (N_19977,N_14116,N_16605);
and U19978 (N_19978,N_14405,N_15136);
or U19979 (N_19979,N_14815,N_15850);
and U19980 (N_19980,N_12842,N_13493);
xor U19981 (N_19981,N_14873,N_14818);
nand U19982 (N_19982,N_15553,N_16752);
nor U19983 (N_19983,N_14101,N_14518);
and U19984 (N_19984,N_15475,N_12556);
nor U19985 (N_19985,N_12245,N_15928);
and U19986 (N_19986,N_15090,N_13054);
xnor U19987 (N_19987,N_14308,N_17398);
nor U19988 (N_19988,N_13947,N_12909);
or U19989 (N_19989,N_16207,N_16184);
xnor U19990 (N_19990,N_14671,N_15355);
nand U19991 (N_19991,N_17787,N_13954);
or U19992 (N_19992,N_12049,N_12491);
nand U19993 (N_19993,N_12203,N_13015);
xnor U19994 (N_19994,N_12582,N_17445);
nand U19995 (N_19995,N_16542,N_13630);
nor U19996 (N_19996,N_16976,N_14850);
or U19997 (N_19997,N_12083,N_13829);
nor U19998 (N_19998,N_16334,N_17879);
xnor U19999 (N_19999,N_14939,N_13040);
nor U20000 (N_20000,N_16955,N_16015);
xor U20001 (N_20001,N_12108,N_14232);
nand U20002 (N_20002,N_16177,N_13143);
nor U20003 (N_20003,N_13914,N_13925);
xor U20004 (N_20004,N_15120,N_15468);
nor U20005 (N_20005,N_16633,N_17600);
nor U20006 (N_20006,N_14298,N_16777);
nor U20007 (N_20007,N_12826,N_17577);
nand U20008 (N_20008,N_12960,N_12146);
and U20009 (N_20009,N_13877,N_12052);
and U20010 (N_20010,N_17730,N_17271);
xnor U20011 (N_20011,N_12211,N_17925);
nor U20012 (N_20012,N_15840,N_15218);
xnor U20013 (N_20013,N_13729,N_13376);
and U20014 (N_20014,N_16838,N_17661);
nand U20015 (N_20015,N_13605,N_15421);
nand U20016 (N_20016,N_12303,N_16591);
xnor U20017 (N_20017,N_13412,N_13603);
nor U20018 (N_20018,N_12807,N_15222);
or U20019 (N_20019,N_17343,N_16495);
nand U20020 (N_20020,N_13423,N_12470);
or U20021 (N_20021,N_12094,N_17918);
xor U20022 (N_20022,N_13942,N_14183);
and U20023 (N_20023,N_14266,N_13944);
nand U20024 (N_20024,N_16790,N_13600);
nor U20025 (N_20025,N_12110,N_12735);
or U20026 (N_20026,N_16045,N_17160);
xor U20027 (N_20027,N_13491,N_16083);
nor U20028 (N_20028,N_16940,N_13086);
nand U20029 (N_20029,N_12911,N_13353);
xnor U20030 (N_20030,N_15083,N_15997);
nand U20031 (N_20031,N_12589,N_17823);
nand U20032 (N_20032,N_17053,N_14268);
xnor U20033 (N_20033,N_13640,N_14238);
xnor U20034 (N_20034,N_13093,N_15718);
and U20035 (N_20035,N_15791,N_13711);
or U20036 (N_20036,N_15691,N_13710);
and U20037 (N_20037,N_16606,N_16498);
nor U20038 (N_20038,N_13068,N_14234);
or U20039 (N_20039,N_16189,N_12513);
nor U20040 (N_20040,N_16365,N_16662);
xor U20041 (N_20041,N_16224,N_17270);
nor U20042 (N_20042,N_15964,N_14373);
xnor U20043 (N_20043,N_12140,N_13784);
nand U20044 (N_20044,N_14504,N_14801);
nand U20045 (N_20045,N_17816,N_15073);
and U20046 (N_20046,N_17723,N_13975);
or U20047 (N_20047,N_17302,N_14746);
nor U20048 (N_20048,N_13928,N_12463);
xor U20049 (N_20049,N_15983,N_12399);
nand U20050 (N_20050,N_15051,N_15542);
xnor U20051 (N_20051,N_17782,N_15507);
and U20052 (N_20052,N_14745,N_15036);
nand U20053 (N_20053,N_15138,N_17668);
xor U20054 (N_20054,N_13190,N_14316);
nor U20055 (N_20055,N_12162,N_13032);
nor U20056 (N_20056,N_12968,N_14962);
and U20057 (N_20057,N_16455,N_16426);
or U20058 (N_20058,N_17832,N_15433);
or U20059 (N_20059,N_13831,N_17391);
xnor U20060 (N_20060,N_15769,N_12461);
nand U20061 (N_20061,N_17642,N_16863);
or U20062 (N_20062,N_13166,N_13534);
and U20063 (N_20063,N_13316,N_17819);
xnor U20064 (N_20064,N_17545,N_12789);
or U20065 (N_20065,N_12707,N_13484);
and U20066 (N_20066,N_14231,N_14423);
xnor U20067 (N_20067,N_14912,N_17028);
xnor U20068 (N_20068,N_12444,N_15975);
and U20069 (N_20069,N_12135,N_13262);
and U20070 (N_20070,N_17893,N_14156);
or U20071 (N_20071,N_13689,N_12685);
xnor U20072 (N_20072,N_13971,N_12879);
or U20073 (N_20073,N_14209,N_14910);
nand U20074 (N_20074,N_15828,N_15274);
nand U20075 (N_20075,N_14705,N_12019);
and U20076 (N_20076,N_17842,N_16041);
and U20077 (N_20077,N_15700,N_14820);
and U20078 (N_20078,N_17914,N_13553);
xor U20079 (N_20079,N_17904,N_12137);
nand U20080 (N_20080,N_12785,N_13715);
and U20081 (N_20081,N_12309,N_17223);
nand U20082 (N_20082,N_16248,N_15459);
and U20083 (N_20083,N_13865,N_16792);
nor U20084 (N_20084,N_15656,N_13136);
or U20085 (N_20085,N_15717,N_12661);
and U20086 (N_20086,N_16879,N_12743);
xnor U20087 (N_20087,N_17259,N_16018);
or U20088 (N_20088,N_15801,N_17888);
nand U20089 (N_20089,N_13800,N_13029);
xnor U20090 (N_20090,N_17968,N_14776);
or U20091 (N_20091,N_13326,N_17599);
nor U20092 (N_20092,N_17235,N_15736);
nand U20093 (N_20093,N_14523,N_15306);
xnor U20094 (N_20094,N_17672,N_17221);
xor U20095 (N_20095,N_12034,N_12054);
xnor U20096 (N_20096,N_12581,N_12763);
and U20097 (N_20097,N_12481,N_13973);
xnor U20098 (N_20098,N_12996,N_16293);
or U20099 (N_20099,N_17959,N_13095);
nand U20100 (N_20100,N_16853,N_15749);
and U20101 (N_20101,N_15657,N_15860);
nor U20102 (N_20102,N_12646,N_15849);
or U20103 (N_20103,N_17573,N_14706);
nand U20104 (N_20104,N_16280,N_13177);
nand U20105 (N_20105,N_14263,N_15889);
nand U20106 (N_20106,N_13358,N_13228);
xnor U20107 (N_20107,N_15208,N_14360);
nand U20108 (N_20108,N_13452,N_16641);
nor U20109 (N_20109,N_16289,N_16025);
xnor U20110 (N_20110,N_16144,N_12548);
nand U20111 (N_20111,N_14707,N_13188);
and U20112 (N_20112,N_17449,N_15315);
xnor U20113 (N_20113,N_17272,N_13521);
nand U20114 (N_20114,N_12324,N_14839);
nor U20115 (N_20115,N_13749,N_14368);
or U20116 (N_20116,N_17386,N_15853);
and U20117 (N_20117,N_13996,N_16561);
nand U20118 (N_20118,N_16629,N_14849);
nand U20119 (N_20119,N_14074,N_17480);
and U20120 (N_20120,N_14790,N_17764);
and U20121 (N_20121,N_14576,N_17805);
nor U20122 (N_20122,N_14273,N_16510);
or U20123 (N_20123,N_15072,N_17450);
nand U20124 (N_20124,N_13976,N_17131);
or U20125 (N_20125,N_12950,N_17032);
xor U20126 (N_20126,N_16238,N_15212);
nand U20127 (N_20127,N_12133,N_13112);
xor U20128 (N_20128,N_17592,N_17463);
and U20129 (N_20129,N_13957,N_13719);
nand U20130 (N_20130,N_14952,N_13950);
and U20131 (N_20131,N_15074,N_12889);
and U20132 (N_20132,N_14380,N_12507);
or U20133 (N_20133,N_13608,N_13411);
or U20134 (N_20134,N_14608,N_14932);
or U20135 (N_20135,N_17857,N_16980);
nor U20136 (N_20136,N_14883,N_13810);
nand U20137 (N_20137,N_15265,N_16415);
nand U20138 (N_20138,N_14115,N_15914);
or U20139 (N_20139,N_13704,N_17086);
nand U20140 (N_20140,N_15705,N_13375);
xor U20141 (N_20141,N_13702,N_15764);
and U20142 (N_20142,N_14288,N_17499);
or U20143 (N_20143,N_14957,N_17218);
nor U20144 (N_20144,N_15910,N_12301);
xor U20145 (N_20145,N_14885,N_17297);
nand U20146 (N_20146,N_17046,N_17676);
nor U20147 (N_20147,N_12554,N_12109);
xnor U20148 (N_20148,N_14604,N_13058);
xnor U20149 (N_20149,N_15966,N_12959);
xor U20150 (N_20150,N_15371,N_12351);
nand U20151 (N_20151,N_16744,N_17641);
and U20152 (N_20152,N_12452,N_12971);
nand U20153 (N_20153,N_16002,N_14534);
or U20154 (N_20154,N_12147,N_14600);
and U20155 (N_20155,N_16610,N_15277);
nor U20156 (N_20156,N_12407,N_13475);
and U20157 (N_20157,N_15707,N_16586);
and U20158 (N_20158,N_16154,N_17795);
xor U20159 (N_20159,N_12246,N_13660);
nor U20160 (N_20160,N_13867,N_16028);
xnor U20161 (N_20161,N_14229,N_12598);
nand U20162 (N_20162,N_17986,N_13135);
nand U20163 (N_20163,N_13880,N_17632);
and U20164 (N_20164,N_14402,N_13620);
nand U20165 (N_20165,N_16431,N_12450);
nor U20166 (N_20166,N_15623,N_16402);
nor U20167 (N_20167,N_14319,N_17935);
nand U20168 (N_20168,N_15692,N_14782);
nand U20169 (N_20169,N_16548,N_17708);
nand U20170 (N_20170,N_15012,N_12886);
nand U20171 (N_20171,N_16063,N_16908);
nand U20172 (N_20172,N_15404,N_12957);
nand U20173 (N_20173,N_15541,N_13186);
and U20174 (N_20174,N_17963,N_14099);
or U20175 (N_20175,N_14737,N_15948);
xnor U20176 (N_20176,N_12625,N_17153);
xnor U20177 (N_20177,N_17362,N_13681);
nor U20178 (N_20178,N_14272,N_13561);
nand U20179 (N_20179,N_13004,N_13118);
nand U20180 (N_20180,N_13701,N_12788);
nand U20181 (N_20181,N_14448,N_16262);
nor U20182 (N_20182,N_15016,N_16814);
nor U20183 (N_20183,N_12225,N_12880);
xnor U20184 (N_20184,N_12991,N_14094);
nor U20185 (N_20185,N_16871,N_14215);
and U20186 (N_20186,N_14869,N_13709);
xor U20187 (N_20187,N_17776,N_15930);
nor U20188 (N_20188,N_12286,N_13813);
xor U20189 (N_20189,N_12216,N_17997);
or U20190 (N_20190,N_17478,N_15375);
xnor U20191 (N_20191,N_13962,N_15223);
nor U20192 (N_20192,N_12529,N_12691);
nor U20193 (N_20193,N_16599,N_12777);
and U20194 (N_20194,N_14609,N_12391);
nor U20195 (N_20195,N_16977,N_15844);
xnor U20196 (N_20196,N_16157,N_14799);
and U20197 (N_20197,N_13161,N_14435);
or U20198 (N_20198,N_12160,N_12618);
nor U20199 (N_20199,N_16648,N_17785);
xnor U20200 (N_20200,N_15758,N_16712);
and U20201 (N_20201,N_15833,N_12072);
nand U20202 (N_20202,N_14427,N_16627);
or U20203 (N_20203,N_16472,N_14258);
or U20204 (N_20204,N_17000,N_17871);
or U20205 (N_20205,N_13457,N_16043);
nand U20206 (N_20206,N_15361,N_16935);
or U20207 (N_20207,N_15759,N_13408);
nand U20208 (N_20208,N_17700,N_14833);
or U20209 (N_20209,N_16987,N_12095);
and U20210 (N_20210,N_15273,N_14103);
or U20211 (N_20211,N_14624,N_16080);
nand U20212 (N_20212,N_15303,N_16490);
or U20213 (N_20213,N_17670,N_17088);
xnor U20214 (N_20214,N_13315,N_15308);
or U20215 (N_20215,N_13588,N_12455);
nor U20216 (N_20216,N_12189,N_16423);
and U20217 (N_20217,N_16319,N_14836);
nor U20218 (N_20218,N_12492,N_16885);
nand U20219 (N_20219,N_14966,N_12969);
xor U20220 (N_20220,N_12565,N_13636);
nor U20221 (N_20221,N_12734,N_15037);
nand U20222 (N_20222,N_16464,N_15154);
and U20223 (N_20223,N_17169,N_17181);
nand U20224 (N_20224,N_17138,N_13544);
xnor U20225 (N_20225,N_15160,N_12647);
nor U20226 (N_20226,N_16991,N_16418);
xor U20227 (N_20227,N_12500,N_16162);
or U20228 (N_20228,N_16270,N_15228);
nand U20229 (N_20229,N_13415,N_14158);
xnor U20230 (N_20230,N_15678,N_13018);
nand U20231 (N_20231,N_15325,N_17394);
nor U20232 (N_20232,N_17274,N_17120);
xnor U20233 (N_20233,N_13847,N_15645);
and U20234 (N_20234,N_15676,N_14151);
xnor U20235 (N_20235,N_16475,N_16911);
and U20236 (N_20236,N_17934,N_16719);
nor U20237 (N_20237,N_17222,N_17490);
or U20238 (N_20238,N_12805,N_12559);
or U20239 (N_20239,N_12629,N_12934);
nand U20240 (N_20240,N_13646,N_12952);
nor U20241 (N_20241,N_17701,N_16179);
nor U20242 (N_20242,N_17129,N_15781);
and U20243 (N_20243,N_16868,N_13035);
xnor U20244 (N_20244,N_17510,N_16930);
nor U20245 (N_20245,N_16660,N_12956);
or U20246 (N_20246,N_14806,N_16433);
and U20247 (N_20247,N_17586,N_15417);
nor U20248 (N_20248,N_15821,N_13302);
xnor U20249 (N_20249,N_14847,N_16588);
nand U20250 (N_20250,N_13834,N_14452);
or U20251 (N_20251,N_17537,N_17113);
and U20252 (N_20252,N_15646,N_12192);
nand U20253 (N_20253,N_15253,N_16489);
or U20254 (N_20254,N_16682,N_17810);
xnor U20255 (N_20255,N_14302,N_13887);
xor U20256 (N_20256,N_14991,N_14346);
nor U20257 (N_20257,N_15052,N_12917);
xor U20258 (N_20258,N_14330,N_17804);
nor U20259 (N_20259,N_16461,N_14694);
and U20260 (N_20260,N_16569,N_17465);
xor U20261 (N_20261,N_12987,N_12202);
and U20262 (N_20262,N_17527,N_15703);
nand U20263 (N_20263,N_17590,N_15924);
nand U20264 (N_20264,N_17674,N_12736);
nand U20265 (N_20265,N_12859,N_14877);
and U20266 (N_20266,N_13742,N_16950);
or U20267 (N_20267,N_13870,N_16918);
xnor U20268 (N_20268,N_12316,N_17624);
nand U20269 (N_20269,N_15234,N_13174);
nand U20270 (N_20270,N_17132,N_15571);
and U20271 (N_20271,N_14700,N_14013);
nand U20272 (N_20272,N_15193,N_14473);
nor U20273 (N_20273,N_17821,N_15166);
and U20274 (N_20274,N_16872,N_14562);
nor U20275 (N_20275,N_17252,N_12213);
and U20276 (N_20276,N_12474,N_17310);
and U20277 (N_20277,N_14043,N_16312);
and U20278 (N_20278,N_15393,N_17268);
xor U20279 (N_20279,N_14526,N_13420);
or U20280 (N_20280,N_14549,N_16645);
nand U20281 (N_20281,N_16553,N_15619);
and U20282 (N_20282,N_12051,N_15146);
and U20283 (N_20283,N_17951,N_12239);
xor U20284 (N_20284,N_17974,N_13169);
nor U20285 (N_20285,N_17389,N_16639);
nor U20286 (N_20286,N_15322,N_17746);
or U20287 (N_20287,N_16545,N_13941);
and U20288 (N_20288,N_15492,N_14289);
xor U20289 (N_20289,N_14636,N_13129);
nand U20290 (N_20290,N_16361,N_16077);
nor U20291 (N_20291,N_13171,N_12902);
or U20292 (N_20292,N_13078,N_17638);
nor U20293 (N_20293,N_14563,N_13120);
and U20294 (N_20294,N_12181,N_17885);
nor U20295 (N_20295,N_13072,N_17434);
xnor U20296 (N_20296,N_15824,N_16282);
xnor U20297 (N_20297,N_17243,N_12680);
and U20298 (N_20298,N_15114,N_12263);
nand U20299 (N_20299,N_12642,N_15797);
nand U20300 (N_20300,N_15205,N_12432);
nor U20301 (N_20301,N_14257,N_12208);
nand U20302 (N_20302,N_16734,N_16649);
nand U20303 (N_20303,N_17910,N_15501);
nand U20304 (N_20304,N_15242,N_16427);
and U20305 (N_20305,N_17576,N_15686);
xor U20306 (N_20306,N_14474,N_17841);
nor U20307 (N_20307,N_12170,N_17628);
nand U20308 (N_20308,N_12524,N_13279);
and U20309 (N_20309,N_15339,N_16173);
or U20310 (N_20310,N_14143,N_12872);
xnor U20311 (N_20311,N_17720,N_13982);
and U20312 (N_20312,N_15877,N_12001);
xor U20313 (N_20313,N_15740,N_13583);
nor U20314 (N_20314,N_17800,N_13249);
xor U20315 (N_20315,N_17660,N_14637);
or U20316 (N_20316,N_17844,N_17518);
and U20317 (N_20317,N_16717,N_15188);
nand U20318 (N_20318,N_12042,N_16556);
or U20319 (N_20319,N_17742,N_13793);
nor U20320 (N_20320,N_14186,N_17735);
nand U20321 (N_20321,N_17655,N_14206);
or U20322 (N_20322,N_15129,N_13637);
or U20323 (N_20323,N_17494,N_13826);
nor U20324 (N_20324,N_17561,N_16882);
nand U20325 (N_20325,N_16851,N_12747);
or U20326 (N_20326,N_16266,N_14584);
or U20327 (N_20327,N_16619,N_16884);
and U20328 (N_20328,N_12846,N_14109);
and U20329 (N_20329,N_13564,N_14301);
and U20330 (N_20330,N_13753,N_17541);
nor U20331 (N_20331,N_13466,N_13109);
and U20332 (N_20332,N_16672,N_17582);
xor U20333 (N_20333,N_17553,N_12539);
or U20334 (N_20334,N_14740,N_17459);
and U20335 (N_20335,N_16075,N_12057);
nand U20336 (N_20336,N_13016,N_13841);
nand U20337 (N_20337,N_14507,N_14840);
nor U20338 (N_20338,N_12584,N_16590);
xnor U20339 (N_20339,N_15883,N_16579);
or U20340 (N_20340,N_16900,N_12021);
nor U20341 (N_20341,N_14314,N_14415);
nand U20342 (N_20342,N_15367,N_12284);
or U20343 (N_20343,N_14393,N_13697);
nand U20344 (N_20344,N_13195,N_12655);
xnor U20345 (N_20345,N_14041,N_17732);
xnor U20346 (N_20346,N_12172,N_15349);
xnor U20347 (N_20347,N_16196,N_16677);
xor U20348 (N_20348,N_17777,N_14411);
or U20349 (N_20349,N_14848,N_15535);
or U20350 (N_20350,N_13180,N_13956);
or U20351 (N_20351,N_13354,N_14048);
nor U20352 (N_20352,N_14307,N_12731);
nor U20353 (N_20353,N_16636,N_13736);
or U20354 (N_20354,N_15590,N_16831);
nand U20355 (N_20355,N_16219,N_12281);
or U20356 (N_20356,N_12080,N_15771);
nand U20357 (N_20357,N_13607,N_15552);
nor U20358 (N_20358,N_17691,N_13577);
nand U20359 (N_20359,N_14054,N_16535);
and U20360 (N_20360,N_17456,N_14290);
nor U20361 (N_20361,N_17596,N_13041);
or U20362 (N_20362,N_12128,N_16304);
and U20363 (N_20363,N_14879,N_12040);
nand U20364 (N_20364,N_12887,N_15508);
and U20365 (N_20365,N_16315,N_13695);
nand U20366 (N_20366,N_16164,N_13555);
and U20367 (N_20367,N_14246,N_17015);
nor U20368 (N_20368,N_16095,N_13788);
or U20369 (N_20369,N_13406,N_16348);
nor U20370 (N_20370,N_15895,N_15990);
or U20371 (N_20371,N_15596,N_14121);
and U20372 (N_20372,N_16644,N_13621);
or U20373 (N_20373,N_14455,N_15502);
nand U20374 (N_20374,N_13597,N_14989);
xnor U20375 (N_20375,N_15614,N_17134);
nand U20376 (N_20376,N_14821,N_16225);
or U20377 (N_20377,N_16125,N_17215);
xor U20378 (N_20378,N_17309,N_13300);
and U20379 (N_20379,N_16393,N_15382);
nor U20380 (N_20380,N_14698,N_13922);
nor U20381 (N_20381,N_13576,N_16534);
xor U20382 (N_20382,N_14867,N_15683);
and U20383 (N_20383,N_13599,N_12607);
nor U20384 (N_20384,N_15254,N_16521);
xnor U20385 (N_20385,N_14886,N_15217);
nand U20386 (N_20386,N_13598,N_17630);
and U20387 (N_20387,N_16689,N_12694);
nand U20388 (N_20388,N_17949,N_17710);
or U20389 (N_20389,N_16843,N_16401);
nand U20390 (N_20390,N_17498,N_12718);
xor U20391 (N_20391,N_16476,N_14018);
and U20392 (N_20392,N_12460,N_13494);
or U20393 (N_20393,N_13522,N_12278);
or U20394 (N_20394,N_12242,N_12570);
and U20395 (N_20395,N_14055,N_12700);
and U20396 (N_20396,N_12841,N_15786);
and U20397 (N_20397,N_17497,N_13184);
and U20398 (N_20398,N_14333,N_15330);
xor U20399 (N_20399,N_13256,N_17350);
or U20400 (N_20400,N_14426,N_12163);
nand U20401 (N_20401,N_16153,N_16199);
xnor U20402 (N_20402,N_15299,N_12808);
nand U20403 (N_20403,N_16623,N_12312);
and U20404 (N_20404,N_16213,N_14020);
or U20405 (N_20405,N_13242,N_15192);
xor U20406 (N_20406,N_16226,N_14322);
xnor U20407 (N_20407,N_13085,N_12400);
nand U20408 (N_20408,N_12439,N_17311);
and U20409 (N_20409,N_14223,N_17470);
nand U20410 (N_20410,N_16921,N_15162);
nor U20411 (N_20411,N_13179,N_16635);
nor U20412 (N_20412,N_17241,N_12297);
and U20413 (N_20413,N_13101,N_14255);
xnor U20414 (N_20414,N_17335,N_15583);
and U20415 (N_20415,N_12313,N_17069);
nand U20416 (N_20416,N_16862,N_13550);
or U20417 (N_20417,N_17713,N_14702);
and U20418 (N_20418,N_14035,N_16869);
nor U20419 (N_20419,N_13499,N_14016);
or U20420 (N_20420,N_12512,N_14339);
or U20421 (N_20421,N_16383,N_15780);
xnor U20422 (N_20422,N_14856,N_14070);
nand U20423 (N_20423,N_17675,N_16452);
nor U20424 (N_20424,N_13267,N_16855);
nor U20425 (N_20425,N_15884,N_17671);
nor U20426 (N_20426,N_14652,N_12928);
xnor U20427 (N_20427,N_14451,N_13859);
nor U20428 (N_20428,N_13439,N_13923);
and U20429 (N_20429,N_16924,N_14987);
nand U20430 (N_20430,N_15261,N_16338);
and U20431 (N_20431,N_13809,N_14172);
nand U20432 (N_20432,N_16837,N_14515);
and U20433 (N_20433,N_15414,N_13849);
nor U20434 (N_20434,N_15101,N_15345);
or U20435 (N_20435,N_13537,N_17896);
xnor U20436 (N_20436,N_16941,N_16784);
and U20437 (N_20437,N_17591,N_17718);
xnor U20438 (N_20438,N_14541,N_15344);
nand U20439 (N_20439,N_14961,N_14328);
or U20440 (N_20440,N_15323,N_12784);
nand U20441 (N_20441,N_13763,N_13217);
and U20442 (N_20442,N_17618,N_12943);
and U20443 (N_20443,N_15510,N_13401);
nand U20444 (N_20444,N_14081,N_12635);
nand U20445 (N_20445,N_12187,N_13269);
and U20446 (N_20446,N_15359,N_14284);
or U20447 (N_20447,N_15995,N_12884);
and U20448 (N_20448,N_13282,N_12397);
xnor U20449 (N_20449,N_13211,N_13509);
xnor U20450 (N_20450,N_13386,N_16440);
xor U20451 (N_20451,N_15954,N_15030);
nand U20452 (N_20452,N_15732,N_15634);
nor U20453 (N_20453,N_14457,N_15802);
nand U20454 (N_20454,N_12354,N_17716);
nand U20455 (N_20455,N_13737,N_14882);
or U20456 (N_20456,N_12469,N_16761);
or U20457 (N_20457,N_12981,N_16158);
nor U20458 (N_20458,N_16079,N_12331);
and U20459 (N_20459,N_16895,N_15873);
nand U20460 (N_20460,N_17182,N_13033);
and U20461 (N_20461,N_12599,N_12449);
nand U20462 (N_20462,N_15737,N_17581);
nor U20463 (N_20463,N_14930,N_15943);
nor U20464 (N_20464,N_16522,N_16405);
nor U20465 (N_20465,N_17097,N_17126);
nand U20466 (N_20466,N_12164,N_16269);
and U20467 (N_20467,N_15660,N_16438);
or U20468 (N_20468,N_14717,N_16260);
or U20469 (N_20469,N_16948,N_14913);
or U20470 (N_20470,N_17295,N_12207);
and U20471 (N_20471,N_15284,N_15342);
xnor U20472 (N_20472,N_17191,N_14334);
or U20473 (N_20473,N_15913,N_12188);
nand U20474 (N_20474,N_14731,N_14495);
and U20475 (N_20475,N_16008,N_14695);
or U20476 (N_20476,N_17960,N_17759);
and U20477 (N_20477,N_17376,N_14096);
and U20478 (N_20478,N_14264,N_17996);
xor U20479 (N_20479,N_14303,N_14778);
nand U20480 (N_20480,N_16034,N_13091);
nor U20481 (N_20481,N_16721,N_15570);
or U20482 (N_20482,N_14742,N_13187);
nand U20483 (N_20483,N_13037,N_16858);
nor U20484 (N_20484,N_16723,N_15810);
nand U20485 (N_20485,N_12440,N_15490);
or U20486 (N_20486,N_17358,N_12314);
nor U20487 (N_20487,N_15595,N_14871);
xnor U20488 (N_20488,N_16943,N_17211);
and U20489 (N_20489,N_13297,N_15245);
xnor U20490 (N_20490,N_17409,N_12002);
and U20491 (N_20491,N_16142,N_17495);
and U20492 (N_20492,N_16251,N_14899);
xnor U20493 (N_20493,N_17090,N_16257);
xnor U20494 (N_20494,N_16410,N_16817);
xor U20495 (N_20495,N_17121,N_14089);
or U20496 (N_20496,N_12527,N_12059);
nor U20497 (N_20497,N_12285,N_17042);
or U20498 (N_20498,N_14237,N_14095);
or U20499 (N_20499,N_14161,N_17995);
nand U20500 (N_20500,N_17639,N_12698);
or U20501 (N_20501,N_12417,N_17695);
xnor U20502 (N_20502,N_12350,N_16026);
nand U20503 (N_20503,N_15092,N_13513);
xor U20504 (N_20504,N_12773,N_14485);
or U20505 (N_20505,N_14794,N_15383);
nor U20506 (N_20506,N_15038,N_12498);
or U20507 (N_20507,N_16578,N_14076);
nand U20508 (N_20508,N_17256,N_16595);
and U20509 (N_20509,N_17351,N_13215);
or U20510 (N_20510,N_14282,N_14386);
nor U20511 (N_20511,N_16772,N_15794);
xor U20512 (N_20512,N_16866,N_17837);
or U20513 (N_20513,N_12226,N_16720);
nor U20514 (N_20514,N_16085,N_17238);
and U20515 (N_20515,N_14195,N_16210);
nor U20516 (N_20516,N_15980,N_16604);
nor U20517 (N_20517,N_17761,N_13434);
nor U20518 (N_20518,N_14429,N_16512);
and U20519 (N_20519,N_17159,N_14808);
xnor U20520 (N_20520,N_13089,N_16005);
nor U20521 (N_20521,N_17283,N_16131);
nor U20522 (N_20522,N_15808,N_15225);
nor U20523 (N_20523,N_14085,N_16108);
nand U20524 (N_20524,N_15819,N_15859);
or U20525 (N_20525,N_13803,N_13649);
or U20526 (N_20526,N_17419,N_12782);
nand U20527 (N_20527,N_17140,N_12709);
nor U20528 (N_20528,N_17557,N_15391);
xor U20529 (N_20529,N_14951,N_16425);
nor U20530 (N_20530,N_17861,N_13418);
or U20531 (N_20531,N_15089,N_17657);
or U20532 (N_20532,N_15197,N_17092);
or U20533 (N_20533,N_17608,N_15517);
or U20534 (N_20534,N_16743,N_17057);
nand U20535 (N_20535,N_17105,N_14953);
and U20536 (N_20536,N_13392,N_16190);
or U20537 (N_20537,N_17429,N_14091);
and U20538 (N_20538,N_14511,N_16004);
nand U20539 (N_20539,N_14458,N_17496);
and U20540 (N_20540,N_15270,N_13992);
or U20541 (N_20541,N_12686,N_15206);
nand U20542 (N_20542,N_13204,N_14915);
nand U20543 (N_20543,N_12561,N_14087);
and U20544 (N_20544,N_13720,N_12878);
and U20545 (N_20545,N_12847,N_17166);
xnor U20546 (N_20546,N_15798,N_12431);
xor U20547 (N_20547,N_16420,N_15027);
nand U20548 (N_20548,N_13327,N_12328);
nor U20549 (N_20549,N_14163,N_16704);
xor U20550 (N_20550,N_13291,N_16971);
and U20551 (N_20551,N_15450,N_17006);
nor U20552 (N_20552,N_13098,N_14281);
nor U20553 (N_20553,N_16249,N_17004);
and U20554 (N_20554,N_15445,N_15155);
xor U20555 (N_20555,N_17125,N_12508);
xnor U20556 (N_20556,N_16245,N_16186);
and U20557 (N_20557,N_15888,N_14320);
and U20558 (N_20558,N_15909,N_15412);
or U20559 (N_20559,N_13172,N_17173);
and U20560 (N_20560,N_17894,N_12039);
or U20561 (N_20561,N_17233,N_16313);
nor U20562 (N_20562,N_14923,N_14739);
nor U20563 (N_20563,N_16699,N_17374);
or U20564 (N_20564,N_16867,N_16353);
or U20565 (N_20565,N_14416,N_13425);
nand U20566 (N_20566,N_14678,N_16688);
or U20567 (N_20567,N_13806,N_15555);
or U20568 (N_20568,N_12877,N_13958);
nand U20569 (N_20569,N_12626,N_14975);
or U20570 (N_20570,N_13290,N_13508);
nor U20571 (N_20571,N_15125,N_15000);
nand U20572 (N_20572,N_14342,N_14551);
nand U20573 (N_20573,N_17936,N_13855);
nor U20574 (N_20574,N_15765,N_17367);
and U20575 (N_20575,N_14168,N_17460);
and U20576 (N_20576,N_13329,N_16488);
nor U20577 (N_20577,N_13554,N_12318);
xor U20578 (N_20578,N_14770,N_15292);
xor U20579 (N_20579,N_14299,N_12795);
or U20580 (N_20580,N_16326,N_15799);
xor U20581 (N_20581,N_17143,N_17965);
nand U20582 (N_20582,N_15994,N_17772);
nand U20583 (N_20583,N_16787,N_17753);
nor U20584 (N_20584,N_13639,N_13459);
nand U20585 (N_20585,N_14437,N_16659);
nand U20586 (N_20586,N_17447,N_12027);
or U20587 (N_20587,N_15091,N_17931);
xnor U20588 (N_20588,N_16683,N_14916);
xnor U20589 (N_20589,N_14639,N_12671);
nand U20590 (N_20590,N_14154,N_12746);
and U20591 (N_20591,N_13233,N_17552);
xnor U20592 (N_20592,N_15423,N_12699);
or U20593 (N_20593,N_13224,N_15599);
or U20594 (N_20594,N_16380,N_15262);
nand U20595 (N_20595,N_15236,N_13427);
and U20596 (N_20596,N_12373,N_13824);
xnor U20597 (N_20597,N_12376,N_12149);
and U20598 (N_20598,N_13882,N_17902);
and U20599 (N_20599,N_13756,N_12649);
nor U20600 (N_20600,N_15438,N_14219);
xor U20601 (N_20601,N_12454,N_13391);
xnor U20602 (N_20602,N_15655,N_12090);
xnor U20603 (N_20603,N_16515,N_15800);
and U20604 (N_20604,N_17142,N_14374);
xnor U20605 (N_20605,N_14430,N_17326);
nand U20606 (N_20606,N_17150,N_16473);
nor U20607 (N_20607,N_12402,N_15488);
and U20608 (N_20608,N_12742,N_17390);
xor U20609 (N_20609,N_17913,N_12931);
and U20610 (N_20610,N_17424,N_14846);
nand U20611 (N_20611,N_15494,N_16048);
nor U20612 (N_20612,N_16970,N_16191);
and U20613 (N_20613,N_15569,N_16141);
nor U20614 (N_20614,N_16813,N_13232);
nand U20615 (N_20615,N_14265,N_16470);
nor U20616 (N_20616,N_15094,N_16697);
and U20617 (N_20617,N_17667,N_17817);
nor U20618 (N_20618,N_15708,N_17240);
and U20619 (N_20619,N_13683,N_15032);
and U20620 (N_20620,N_16253,N_12720);
and U20621 (N_20621,N_14462,N_17408);
xor U20622 (N_20622,N_17715,N_16258);
nand U20623 (N_20623,N_13703,N_17749);
nor U20624 (N_20624,N_17898,N_16906);
or U20625 (N_20625,N_14122,N_14428);
or U20626 (N_20626,N_17083,N_16453);
xor U20627 (N_20627,N_16303,N_12929);
nand U20628 (N_20628,N_15482,N_16982);
and U20629 (N_20629,N_12849,N_15548);
nand U20630 (N_20630,N_14662,N_15751);
and U20631 (N_20631,N_14167,N_16356);
nand U20632 (N_20632,N_17466,N_16565);
nand U20633 (N_20633,N_13230,N_16193);
or U20634 (N_20634,N_14080,N_14841);
and U20635 (N_20635,N_14784,N_13350);
nor U20636 (N_20636,N_13454,N_14665);
and U20637 (N_20637,N_12986,N_13156);
nor U20638 (N_20638,N_12499,N_16770);
xor U20639 (N_20639,N_13036,N_17370);
nand U20640 (N_20640,N_12770,N_15269);
nand U20641 (N_20641,N_16638,N_12209);
or U20642 (N_20642,N_17707,N_14147);
and U20643 (N_20643,N_12333,N_14253);
nand U20644 (N_20644,N_16830,N_15899);
xor U20645 (N_20645,N_12011,N_14904);
and U20646 (N_20646,N_14440,N_13610);
nor U20647 (N_20647,N_14261,N_12888);
xor U20648 (N_20648,N_16780,N_15957);
nand U20649 (N_20649,N_15633,N_14734);
nor U20650 (N_20650,N_17634,N_14097);
and U20651 (N_20651,N_15823,N_16655);
nand U20652 (N_20652,N_14224,N_12385);
or U20653 (N_20653,N_15935,N_12705);
and U20654 (N_20654,N_17371,N_13431);
nand U20655 (N_20655,N_12799,N_14566);
nand U20656 (N_20656,N_15327,N_16391);
nor U20657 (N_20657,N_13611,N_14606);
and U20658 (N_20658,N_13629,N_14775);
xor U20659 (N_20659,N_15558,N_12200);
and U20660 (N_20660,N_15972,N_15839);
and U20661 (N_20661,N_13364,N_16880);
xnor U20662 (N_20662,N_15567,N_16816);
xor U20663 (N_20663,N_17994,N_16523);
and U20664 (N_20664,N_13053,N_15757);
nand U20665 (N_20665,N_13929,N_17387);
or U20666 (N_20666,N_16764,N_12262);
nand U20667 (N_20667,N_16283,N_15601);
or U20668 (N_20668,N_16411,N_12708);
and U20669 (N_20669,N_13435,N_17901);
nor U20670 (N_20670,N_15116,N_15111);
nand U20671 (N_20671,N_17886,N_13355);
and U20672 (N_20672,N_14569,N_16577);
and U20673 (N_20673,N_14598,N_12259);
nor U20674 (N_20674,N_15388,N_16301);
nand U20675 (N_20675,N_15912,N_12082);
or U20676 (N_20676,N_16611,N_14653);
nand U20677 (N_20677,N_15534,N_13082);
nand U20678 (N_20678,N_16174,N_14479);
xor U20679 (N_20679,N_16116,N_15077);
xor U20680 (N_20680,N_12056,N_14755);
xnor U20681 (N_20681,N_12916,N_13657);
or U20682 (N_20682,N_15260,N_13745);
or U20683 (N_20683,N_17100,N_16961);
xor U20684 (N_20684,N_14854,N_16297);
and U20685 (N_20685,N_15311,N_13526);
xnor U20686 (N_20686,N_15674,N_12615);
nor U20687 (N_20687,N_14313,N_12038);
nand U20688 (N_20688,N_13644,N_15743);
xor U20689 (N_20689,N_13235,N_12989);
nand U20690 (N_20690,N_14480,N_14376);
nand U20691 (N_20691,N_17196,N_12840);
xnor U20692 (N_20692,N_17476,N_12401);
nand U20693 (N_20693,N_12976,N_13266);
nand U20694 (N_20694,N_17485,N_14875);
xor U20695 (N_20695,N_13949,N_13333);
nor U20696 (N_20696,N_13523,N_17025);
xnor U20697 (N_20697,N_13134,N_17932);
nand U20698 (N_20698,N_15081,N_16740);
or U20699 (N_20699,N_16806,N_15921);
or U20700 (N_20700,N_12016,N_12568);
nand U20701 (N_20701,N_14200,N_12473);
xnor U20702 (N_20702,N_13369,N_13319);
nor U20703 (N_20703,N_17071,N_12106);
nand U20704 (N_20704,N_14767,N_13680);
and U20705 (N_20705,N_14567,N_12060);
nor U20706 (N_20706,N_12744,N_14084);
xor U20707 (N_20707,N_15929,N_14858);
xor U20708 (N_20708,N_14785,N_16501);
and U20709 (N_20709,N_16922,N_13450);
nor U20710 (N_20710,N_15370,N_17948);
and U20711 (N_20711,N_12260,N_12014);
and U20712 (N_20712,N_16271,N_15681);
nand U20713 (N_20713,N_15246,N_12319);
or U20714 (N_20714,N_14893,N_12693);
nand U20715 (N_20715,N_14059,N_14171);
or U20716 (N_20716,N_16229,N_16036);
xnor U20717 (N_20717,N_15446,N_12940);
xor U20718 (N_20718,N_16188,N_13259);
and U20719 (N_20719,N_16375,N_16502);
nor U20720 (N_20720,N_16364,N_15276);
nand U20721 (N_20721,N_14024,N_15602);
nor U20722 (N_20722,N_14764,N_12566);
or U20723 (N_20723,N_15171,N_15869);
nor U20724 (N_20724,N_14673,N_15933);
or U20725 (N_20725,N_13628,N_12797);
xor U20726 (N_20726,N_12103,N_17493);
or U20727 (N_20727,N_15461,N_14125);
and U20728 (N_20728,N_16054,N_15605);
xnor U20729 (N_20729,N_17881,N_14772);
nand U20730 (N_20730,N_14492,N_17161);
nor U20731 (N_20731,N_15215,N_14021);
or U20732 (N_20732,N_14754,N_14685);
nand U20733 (N_20733,N_14002,N_14540);
or U20734 (N_20734,N_14900,N_15159);
or U20735 (N_20735,N_17417,N_14201);
nor U20736 (N_20736,N_13886,N_12684);
and U20737 (N_20737,N_13445,N_12173);
and U20738 (N_20738,N_13790,N_13570);
and U20739 (N_20739,N_12683,N_12930);
xor U20740 (N_20740,N_16175,N_16007);
or U20741 (N_20741,N_13850,N_15021);
nor U20742 (N_20742,N_12012,N_13189);
or U20743 (N_20743,N_17165,N_13003);
and U20744 (N_20744,N_15637,N_16259);
or U20745 (N_20745,N_12781,N_13122);
nand U20746 (N_20746,N_15679,N_12863);
and U20747 (N_20747,N_15755,N_15868);
or U20748 (N_20748,N_15931,N_16267);
and U20749 (N_20749,N_14844,N_14644);
nand U20750 (N_20750,N_17953,N_15876);
nor U20751 (N_20751,N_15880,N_17836);
and U20752 (N_20752,N_12013,N_14446);
xor U20753 (N_20753,N_14256,N_15723);
or U20754 (N_20754,N_14670,N_17430);
or U20755 (N_20755,N_17313,N_13321);
and U20756 (N_20756,N_15865,N_14027);
nor U20757 (N_20757,N_17598,N_12017);
nor U20758 (N_20758,N_17884,N_12300);
xnor U20759 (N_20759,N_16944,N_12416);
nand U20760 (N_20760,N_14129,N_13931);
or U20761 (N_20761,N_13294,N_15597);
xor U20762 (N_20762,N_13081,N_13080);
nor U20763 (N_20763,N_16044,N_14131);
or U20764 (N_20764,N_14075,N_15826);
nor U20765 (N_20765,N_16479,N_13574);
nand U20766 (N_20766,N_17853,N_12156);
or U20767 (N_20767,N_12650,N_15942);
or U20768 (N_20768,N_13741,N_17227);
xnor U20769 (N_20769,N_16979,N_16161);
nor U20770 (N_20770,N_16032,N_13774);
or U20771 (N_20771,N_13264,N_14204);
xnor U20772 (N_20772,N_14032,N_17964);
nand U20773 (N_20773,N_12862,N_13897);
and U20774 (N_20774,N_12605,N_13311);
xnor U20775 (N_20775,N_14228,N_13917);
xor U20776 (N_20776,N_15295,N_17264);
and U20777 (N_20777,N_14810,N_12010);
or U20778 (N_20778,N_16485,N_14555);
or U20779 (N_20779,N_15667,N_16722);
xor U20780 (N_20780,N_12145,N_13739);
and U20781 (N_20781,N_12247,N_15221);
xor U20782 (N_20782,N_15285,N_15055);
xor U20783 (N_20783,N_13360,N_14488);
nor U20784 (N_20784,N_13107,N_15538);
or U20785 (N_20785,N_12036,N_13825);
xnor U20786 (N_20786,N_12227,N_14774);
or U20787 (N_20787,N_13337,N_12288);
nand U20788 (N_20788,N_15187,N_16795);
nor U20789 (N_20789,N_12939,N_15066);
and U20790 (N_20790,N_15476,N_17364);
nor U20791 (N_20791,N_17018,N_17205);
nor U20792 (N_20792,N_13979,N_15426);
or U20793 (N_20793,N_13251,N_15282);
nor U20794 (N_20794,N_14832,N_16329);
nor U20795 (N_20795,N_12796,N_14669);
nor U20796 (N_20796,N_13738,N_12831);
xor U20797 (N_20797,N_15153,N_12656);
and U20798 (N_20798,N_14960,N_16120);
and U20799 (N_20799,N_14531,N_16012);
xnor U20800 (N_20800,N_17877,N_15477);
xnor U20801 (N_20801,N_14318,N_12139);
or U20802 (N_20802,N_15996,N_16500);
xor U20803 (N_20803,N_15317,N_13985);
or U20804 (N_20804,N_12759,N_13428);
xnor U20805 (N_20805,N_14383,N_12325);
xor U20806 (N_20806,N_14484,N_14918);
and U20807 (N_20807,N_16696,N_14494);
xor U20808 (N_20808,N_13530,N_14493);
xnor U20809 (N_20809,N_16665,N_15652);
and U20810 (N_20810,N_16277,N_15539);
xor U20811 (N_20811,N_17116,N_12514);
or U20812 (N_20812,N_15950,N_16745);
nand U20813 (N_20813,N_15109,N_14475);
and U20814 (N_20814,N_13609,N_17282);
nand U20815 (N_20815,N_16268,N_14396);
nor U20816 (N_20816,N_15807,N_17620);
xnor U20817 (N_20817,N_15453,N_12268);
nand U20818 (N_20818,N_13022,N_16347);
xor U20819 (N_20819,N_15247,N_14399);
nor U20820 (N_20820,N_13998,N_15064);
and U20821 (N_20821,N_15945,N_15107);
nand U20822 (N_20822,N_14398,N_16958);
xnor U20823 (N_20823,N_13655,N_17743);
xnor U20824 (N_20824,N_14668,N_13765);
nor U20825 (N_20825,N_14431,N_17488);
or U20826 (N_20826,N_16800,N_14834);
xnor U20827 (N_20827,N_14454,N_12814);
or U20828 (N_20828,N_14052,N_15485);
nor U20829 (N_20829,N_15025,N_12738);
or U20830 (N_20830,N_13209,N_16593);
and U20831 (N_20831,N_17341,N_14140);
nand U20832 (N_20832,N_13910,N_15984);
and U20833 (N_20833,N_13398,N_17797);
nor U20834 (N_20834,N_12115,N_12761);
or U20835 (N_20835,N_15594,N_14890);
nand U20836 (N_20836,N_15479,N_14379);
or U20837 (N_20837,N_17719,N_12479);
or U20838 (N_20838,N_16615,N_12927);
xnor U20839 (N_20839,N_15615,N_16966);
nand U20840 (N_20840,N_12266,N_15761);
nand U20841 (N_20841,N_15858,N_14730);
or U20842 (N_20842,N_13967,N_16964);
or U20843 (N_20843,N_15183,N_16580);
nor U20844 (N_20844,N_15878,N_15069);
or U20845 (N_20845,N_14914,N_13014);
nand U20846 (N_20846,N_14510,N_16758);
and U20847 (N_20847,N_15863,N_15156);
and U20848 (N_20848,N_16575,N_16739);
or U20849 (N_20849,N_14150,N_17454);
xnor U20850 (N_20850,N_12327,N_17383);
nand U20851 (N_20851,N_16781,N_16507);
or U20852 (N_20852,N_15158,N_17439);
nor U20853 (N_20853,N_14626,N_12725);
xor U20854 (N_20854,N_13104,N_12388);
nor U20855 (N_20855,N_13288,N_14164);
or U20856 (N_20856,N_15625,N_16738);
and U20857 (N_20857,N_13238,N_12533);
xor U20858 (N_20858,N_16767,N_12212);
nand U20859 (N_20859,N_13203,N_17263);
xnor U20860 (N_20860,N_17999,N_12390);
xor U20861 (N_20861,N_13332,N_14974);
xor U20862 (N_20862,N_13926,N_15252);
nand U20863 (N_20863,N_14472,N_14787);
or U20864 (N_20864,N_15752,N_13413);
nand U20865 (N_20865,N_13707,N_17725);
xnor U20866 (N_20866,N_15002,N_17717);
and U20867 (N_20867,N_17014,N_13533);
and U20868 (N_20868,N_14864,N_14557);
or U20869 (N_20869,N_15991,N_16891);
and U20870 (N_20870,N_12047,N_12608);
xnor U20871 (N_20871,N_17587,N_16666);
xor U20872 (N_20872,N_16435,N_15194);
nor U20873 (N_20873,N_14736,N_13618);
and U20874 (N_20874,N_14789,N_14247);
or U20875 (N_20875,N_12412,N_17852);
nand U20876 (N_20876,N_16760,N_16300);
or U20877 (N_20877,N_16988,N_13404);
and U20878 (N_20878,N_16733,N_14092);
nor U20879 (N_20879,N_13305,N_13432);
or U20880 (N_20880,N_14920,N_14295);
xor U20881 (N_20881,N_13012,N_12733);
or U20882 (N_20882,N_17589,N_17084);
nor U20883 (N_20883,N_14722,N_13448);
xor U20884 (N_20884,N_14222,N_16564);
nand U20885 (N_20885,N_17400,N_15368);
or U20886 (N_20886,N_13921,N_13164);
nor U20887 (N_20887,N_14477,N_14486);
or U20888 (N_20888,N_13938,N_16530);
nand U20889 (N_20889,N_15976,N_12165);
nor U20890 (N_20890,N_16592,N_14086);
or U20891 (N_20891,N_17507,N_14797);
and U20892 (N_20892,N_17571,N_14198);
nor U20893 (N_20893,N_13902,N_16445);
xor U20894 (N_20894,N_12622,N_17763);
xor U20895 (N_20895,N_13050,N_17399);
nand U20896 (N_20896,N_15331,N_17474);
xnor U20897 (N_20897,N_12168,N_16985);
and U20898 (N_20898,N_14814,N_12844);
and U20899 (N_20899,N_12153,N_12240);
or U20900 (N_20900,N_13092,N_16374);
or U20901 (N_20901,N_13895,N_12851);
xor U20902 (N_20902,N_13746,N_15744);
or U20903 (N_20903,N_14661,N_16316);
nor U20904 (N_20904,N_17133,N_15624);
or U20905 (N_20905,N_12277,N_17911);
and U20906 (N_20906,N_17532,N_13721);
or U20907 (N_20907,N_15419,N_15530);
nor U20908 (N_20908,N_12715,N_14012);
xnor U20909 (N_20909,N_16714,N_16273);
or U20910 (N_20910,N_17037,N_13670);
nand U20911 (N_20911,N_15473,N_14587);
or U20912 (N_20912,N_15709,N_14825);
nor U20913 (N_20913,N_17096,N_14269);
nor U20914 (N_20914,N_13764,N_17546);
or U20915 (N_20915,N_17933,N_17883);
nand U20916 (N_20916,N_17706,N_12231);
or U20917 (N_20917,N_12437,N_13191);
nand U20918 (N_20918,N_17435,N_12638);
and U20919 (N_20919,N_17659,N_13421);
or U20920 (N_20920,N_14381,N_15068);
nand U20921 (N_20921,N_13487,N_17669);
nor U20922 (N_20922,N_14037,N_12907);
nor U20923 (N_20923,N_12476,N_12141);
xor U20924 (N_20924,N_14933,N_13798);
and U20925 (N_20925,N_17135,N_17404);
and U20926 (N_20926,N_16532,N_17643);
and U20927 (N_20927,N_13308,N_14538);
xnor U20928 (N_20928,N_16691,N_16798);
or U20929 (N_20929,N_14159,N_14727);
nand U20930 (N_20930,N_15491,N_16596);
and U20931 (N_20931,N_14599,N_12353);
xor U20932 (N_20932,N_17575,N_15484);
and U20933 (N_20933,N_16087,N_15338);
nand U20934 (N_20934,N_12739,N_15721);
or U20935 (N_20935,N_12610,N_13623);
nand U20936 (N_20936,N_13823,N_16163);
nand U20937 (N_20937,N_17993,N_12045);
nor U20938 (N_20938,N_12236,N_15959);
nand U20939 (N_20939,N_16477,N_16750);
nor U20940 (N_20940,N_12079,N_14409);
nor U20941 (N_20941,N_14502,N_12424);
xnor U20942 (N_20942,N_17711,N_14287);
or U20943 (N_20943,N_15958,N_17141);
and U20944 (N_20944,N_15561,N_17961);
nand U20945 (N_20945,N_14781,N_14530);
xor U20946 (N_20946,N_15100,N_13678);
and U20947 (N_20947,N_12536,N_14309);
nand U20948 (N_20948,N_15142,N_13341);
or U20949 (N_20949,N_15126,N_15432);
nand U20950 (N_20950,N_12210,N_14708);
or U20951 (N_20951,N_14968,N_13359);
or U20952 (N_20952,N_14762,N_16755);
xnor U20953 (N_20953,N_12913,N_14011);
nand U20954 (N_20954,N_16967,N_13474);
nor U20955 (N_20955,N_17077,N_13451);
or U20956 (N_20956,N_13650,N_17047);
and U20957 (N_20957,N_14194,N_12905);
or U20958 (N_20958,N_17144,N_13879);
nand U20959 (N_20959,N_15896,N_15449);
nor U20960 (N_20960,N_15861,N_16242);
nor U20961 (N_20961,N_12827,N_17082);
and U20962 (N_20962,N_16214,N_14658);
nor U20963 (N_20963,N_13476,N_15460);
or U20964 (N_20964,N_12644,N_12817);
nand U20965 (N_20965,N_16968,N_17438);
or U20966 (N_20966,N_15147,N_17253);
and U20967 (N_20967,N_14410,N_14023);
and U20968 (N_20968,N_17900,N_12979);
and U20969 (N_20969,N_17529,N_12553);
nor U20970 (N_20970,N_12237,N_15009);
nand U20971 (N_20971,N_15105,N_16060);
nor U20972 (N_20972,N_16454,N_14025);
nor U20973 (N_20973,N_15733,N_16058);
and U20974 (N_20974,N_17828,N_16618);
nand U20975 (N_20975,N_17567,N_15369);
nand U20976 (N_20976,N_13757,N_12549);
and U20977 (N_20977,N_16448,N_13307);
nor U20978 (N_20978,N_12129,N_12201);
nand U20979 (N_20979,N_17375,N_14664);
nand U20980 (N_20980,N_15113,N_13899);
nor U20981 (N_20981,N_12696,N_17899);
or U20982 (N_20982,N_15662,N_17194);
nor U20983 (N_20983,N_16703,N_12970);
or U20984 (N_20984,N_13616,N_15770);
nor U20985 (N_20985,N_14113,N_17207);
and U20986 (N_20986,N_13904,N_15695);
nor U20987 (N_20987,N_13245,N_15879);
or U20988 (N_20988,N_17550,N_13761);
and U20989 (N_20989,N_15054,N_14816);
or U20990 (N_20990,N_12148,N_14964);
nor U20991 (N_20991,N_15588,N_13568);
xnor U20992 (N_20992,N_17338,N_15165);
nor U20993 (N_20993,N_13362,N_15864);
and U20994 (N_20994,N_12311,N_16160);
and U20995 (N_20995,N_15547,N_12560);
nor U20996 (N_20996,N_14145,N_17118);
nor U20997 (N_20997,N_15070,N_12100);
or U20998 (N_20998,N_12197,N_17688);
xnor U20999 (N_20999,N_17385,N_15024);
or U21000 (N_21000,N_17162,N_15123);
nor U21001 (N_21001,N_17226,N_17612);
xor U21002 (N_21002,N_16333,N_17565);
nand U21003 (N_21003,N_13275,N_16283);
and U21004 (N_21004,N_14396,N_12698);
nand U21005 (N_21005,N_16191,N_16927);
nand U21006 (N_21006,N_15478,N_13044);
and U21007 (N_21007,N_14903,N_13907);
nand U21008 (N_21008,N_13489,N_16371);
xor U21009 (N_21009,N_12495,N_17213);
and U21010 (N_21010,N_13858,N_12241);
or U21011 (N_21011,N_12720,N_16237);
or U21012 (N_21012,N_16456,N_15435);
and U21013 (N_21013,N_16446,N_14742);
and U21014 (N_21014,N_17525,N_16854);
xnor U21015 (N_21015,N_17407,N_16908);
nor U21016 (N_21016,N_17050,N_13365);
and U21017 (N_21017,N_15454,N_15686);
or U21018 (N_21018,N_14462,N_16589);
xor U21019 (N_21019,N_12755,N_15905);
nor U21020 (N_21020,N_14509,N_12028);
or U21021 (N_21021,N_12787,N_14263);
nand U21022 (N_21022,N_14411,N_15076);
and U21023 (N_21023,N_14106,N_12159);
or U21024 (N_21024,N_14686,N_13652);
or U21025 (N_21025,N_13056,N_15700);
and U21026 (N_21026,N_15159,N_13998);
xnor U21027 (N_21027,N_15333,N_14914);
nor U21028 (N_21028,N_16328,N_13114);
nor U21029 (N_21029,N_17251,N_13931);
nand U21030 (N_21030,N_17169,N_13620);
and U21031 (N_21031,N_16975,N_16503);
nand U21032 (N_21032,N_17126,N_12612);
nand U21033 (N_21033,N_17274,N_17974);
or U21034 (N_21034,N_16473,N_12886);
xor U21035 (N_21035,N_14336,N_13240);
and U21036 (N_21036,N_17195,N_14403);
nand U21037 (N_21037,N_17039,N_14948);
and U21038 (N_21038,N_14350,N_15991);
nor U21039 (N_21039,N_14770,N_13856);
nand U21040 (N_21040,N_13336,N_13565);
nor U21041 (N_21041,N_12315,N_17062);
xnor U21042 (N_21042,N_17933,N_13144);
or U21043 (N_21043,N_12717,N_13894);
or U21044 (N_21044,N_14708,N_14619);
nor U21045 (N_21045,N_16799,N_13483);
and U21046 (N_21046,N_15226,N_12386);
or U21047 (N_21047,N_16641,N_15894);
or U21048 (N_21048,N_12930,N_13342);
xor U21049 (N_21049,N_14252,N_12781);
nand U21050 (N_21050,N_14771,N_17507);
and U21051 (N_21051,N_15792,N_16188);
and U21052 (N_21052,N_16832,N_13141);
nor U21053 (N_21053,N_12032,N_15260);
nor U21054 (N_21054,N_13216,N_13820);
or U21055 (N_21055,N_12875,N_15393);
or U21056 (N_21056,N_15222,N_16742);
and U21057 (N_21057,N_17011,N_17943);
or U21058 (N_21058,N_15930,N_16371);
nand U21059 (N_21059,N_15028,N_17022);
xnor U21060 (N_21060,N_14983,N_16903);
nand U21061 (N_21061,N_14401,N_12785);
or U21062 (N_21062,N_12172,N_15735);
or U21063 (N_21063,N_14979,N_14016);
xor U21064 (N_21064,N_12007,N_15888);
or U21065 (N_21065,N_13422,N_14254);
nand U21066 (N_21066,N_12596,N_14033);
nor U21067 (N_21067,N_15586,N_12874);
nor U21068 (N_21068,N_16595,N_13411);
xor U21069 (N_21069,N_16299,N_13262);
nand U21070 (N_21070,N_17572,N_14968);
or U21071 (N_21071,N_16215,N_16116);
or U21072 (N_21072,N_12554,N_13501);
nor U21073 (N_21073,N_15687,N_17756);
nor U21074 (N_21074,N_13236,N_16424);
xor U21075 (N_21075,N_16156,N_13228);
and U21076 (N_21076,N_12267,N_12015);
xor U21077 (N_21077,N_16994,N_12303);
nor U21078 (N_21078,N_12302,N_17911);
or U21079 (N_21079,N_12606,N_15196);
nand U21080 (N_21080,N_12231,N_13680);
nand U21081 (N_21081,N_15737,N_14933);
or U21082 (N_21082,N_17480,N_12346);
xor U21083 (N_21083,N_14777,N_16754);
xnor U21084 (N_21084,N_16145,N_12747);
nand U21085 (N_21085,N_15660,N_16260);
xor U21086 (N_21086,N_17190,N_13341);
or U21087 (N_21087,N_13314,N_15202);
and U21088 (N_21088,N_16295,N_14859);
nand U21089 (N_21089,N_17151,N_14401);
or U21090 (N_21090,N_12525,N_12873);
or U21091 (N_21091,N_16739,N_14047);
and U21092 (N_21092,N_16434,N_15053);
xnor U21093 (N_21093,N_14214,N_17332);
xor U21094 (N_21094,N_12516,N_17480);
xor U21095 (N_21095,N_13776,N_16395);
xnor U21096 (N_21096,N_16825,N_14629);
xnor U21097 (N_21097,N_12124,N_17612);
nand U21098 (N_21098,N_17230,N_16876);
xnor U21099 (N_21099,N_13994,N_16051);
nor U21100 (N_21100,N_16664,N_16478);
nor U21101 (N_21101,N_16860,N_12584);
or U21102 (N_21102,N_14545,N_13134);
and U21103 (N_21103,N_14972,N_13792);
xnor U21104 (N_21104,N_14076,N_15725);
nor U21105 (N_21105,N_15636,N_16035);
nor U21106 (N_21106,N_17681,N_14588);
and U21107 (N_21107,N_14714,N_12719);
or U21108 (N_21108,N_16755,N_12004);
or U21109 (N_21109,N_12251,N_15181);
or U21110 (N_21110,N_15128,N_17729);
or U21111 (N_21111,N_17001,N_13342);
nand U21112 (N_21112,N_14215,N_16580);
nand U21113 (N_21113,N_15647,N_13447);
or U21114 (N_21114,N_16543,N_12306);
or U21115 (N_21115,N_14296,N_12850);
xnor U21116 (N_21116,N_14545,N_13504);
nor U21117 (N_21117,N_16827,N_12225);
xor U21118 (N_21118,N_16445,N_17388);
and U21119 (N_21119,N_15831,N_17243);
or U21120 (N_21120,N_12500,N_14755);
nand U21121 (N_21121,N_16868,N_12512);
nor U21122 (N_21122,N_13179,N_13911);
or U21123 (N_21123,N_12564,N_12122);
and U21124 (N_21124,N_16371,N_16603);
or U21125 (N_21125,N_17192,N_17441);
and U21126 (N_21126,N_13767,N_17456);
and U21127 (N_21127,N_16470,N_17624);
nor U21128 (N_21128,N_16752,N_12364);
xor U21129 (N_21129,N_12688,N_17426);
nand U21130 (N_21130,N_12505,N_17715);
xnor U21131 (N_21131,N_14647,N_12869);
nand U21132 (N_21132,N_15966,N_16131);
xnor U21133 (N_21133,N_14373,N_12105);
nand U21134 (N_21134,N_15509,N_16391);
or U21135 (N_21135,N_16007,N_13508);
xor U21136 (N_21136,N_12965,N_17384);
nand U21137 (N_21137,N_12791,N_14136);
and U21138 (N_21138,N_12264,N_13694);
nand U21139 (N_21139,N_12448,N_13589);
nand U21140 (N_21140,N_17805,N_16835);
xnor U21141 (N_21141,N_17792,N_14780);
or U21142 (N_21142,N_12010,N_12156);
nor U21143 (N_21143,N_12536,N_17309);
xnor U21144 (N_21144,N_16175,N_14221);
and U21145 (N_21145,N_15715,N_13285);
or U21146 (N_21146,N_15692,N_16541);
nand U21147 (N_21147,N_15400,N_17806);
or U21148 (N_21148,N_15741,N_16664);
nand U21149 (N_21149,N_15042,N_16013);
xnor U21150 (N_21150,N_17745,N_13724);
or U21151 (N_21151,N_17371,N_14160);
and U21152 (N_21152,N_16962,N_14908);
xnor U21153 (N_21153,N_17651,N_17530);
or U21154 (N_21154,N_13710,N_17489);
nand U21155 (N_21155,N_17619,N_17066);
or U21156 (N_21156,N_13605,N_13421);
nor U21157 (N_21157,N_15996,N_12756);
xnor U21158 (N_21158,N_16265,N_16163);
nor U21159 (N_21159,N_17493,N_14600);
xnor U21160 (N_21160,N_17089,N_13581);
or U21161 (N_21161,N_17666,N_14057);
and U21162 (N_21162,N_14841,N_13033);
nor U21163 (N_21163,N_17014,N_13937);
xnor U21164 (N_21164,N_17817,N_14052);
nor U21165 (N_21165,N_15916,N_16008);
or U21166 (N_21166,N_14958,N_13331);
xnor U21167 (N_21167,N_13485,N_13171);
xnor U21168 (N_21168,N_17136,N_17730);
nand U21169 (N_21169,N_16994,N_16133);
and U21170 (N_21170,N_17446,N_16859);
xnor U21171 (N_21171,N_17182,N_13296);
nand U21172 (N_21172,N_17202,N_13535);
xnor U21173 (N_21173,N_13014,N_14733);
or U21174 (N_21174,N_14802,N_12544);
and U21175 (N_21175,N_15930,N_15089);
xnor U21176 (N_21176,N_13727,N_14829);
nor U21177 (N_21177,N_16212,N_14072);
nand U21178 (N_21178,N_14901,N_15523);
nand U21179 (N_21179,N_16213,N_12297);
nor U21180 (N_21180,N_12092,N_14153);
nand U21181 (N_21181,N_16130,N_13296);
xor U21182 (N_21182,N_14831,N_13766);
or U21183 (N_21183,N_12992,N_14998);
nor U21184 (N_21184,N_14584,N_13275);
nor U21185 (N_21185,N_14948,N_15750);
or U21186 (N_21186,N_14836,N_12806);
xor U21187 (N_21187,N_17761,N_13991);
or U21188 (N_21188,N_13948,N_14986);
and U21189 (N_21189,N_13241,N_13820);
and U21190 (N_21190,N_17305,N_13222);
xnor U21191 (N_21191,N_13065,N_12164);
nor U21192 (N_21192,N_15721,N_17803);
nor U21193 (N_21193,N_16354,N_14348);
nand U21194 (N_21194,N_15022,N_17263);
nor U21195 (N_21195,N_16786,N_15427);
nand U21196 (N_21196,N_17963,N_17577);
nor U21197 (N_21197,N_14337,N_17815);
nand U21198 (N_21198,N_17752,N_12048);
xor U21199 (N_21199,N_14331,N_12265);
or U21200 (N_21200,N_13233,N_16431);
xnor U21201 (N_21201,N_15744,N_13278);
or U21202 (N_21202,N_15753,N_13640);
nor U21203 (N_21203,N_12301,N_15223);
and U21204 (N_21204,N_17344,N_13776);
nand U21205 (N_21205,N_16235,N_13728);
or U21206 (N_21206,N_17460,N_12427);
and U21207 (N_21207,N_14620,N_15725);
or U21208 (N_21208,N_16077,N_12357);
or U21209 (N_21209,N_13813,N_16597);
or U21210 (N_21210,N_17064,N_12865);
xor U21211 (N_21211,N_13453,N_12544);
nor U21212 (N_21212,N_13297,N_13035);
or U21213 (N_21213,N_12714,N_14455);
nand U21214 (N_21214,N_14788,N_17810);
nor U21215 (N_21215,N_16077,N_17358);
xor U21216 (N_21216,N_17014,N_14796);
nor U21217 (N_21217,N_14908,N_12021);
or U21218 (N_21218,N_12313,N_15211);
nor U21219 (N_21219,N_12352,N_14546);
nand U21220 (N_21220,N_16570,N_17059);
nand U21221 (N_21221,N_13974,N_17234);
and U21222 (N_21222,N_12153,N_14378);
nand U21223 (N_21223,N_14683,N_13772);
or U21224 (N_21224,N_15697,N_17342);
xor U21225 (N_21225,N_16131,N_14352);
and U21226 (N_21226,N_13416,N_17053);
nand U21227 (N_21227,N_14686,N_14621);
or U21228 (N_21228,N_14219,N_16318);
xor U21229 (N_21229,N_12442,N_13719);
xor U21230 (N_21230,N_16849,N_16868);
nand U21231 (N_21231,N_16742,N_12045);
and U21232 (N_21232,N_15939,N_12585);
or U21233 (N_21233,N_17809,N_16347);
and U21234 (N_21234,N_14182,N_12834);
and U21235 (N_21235,N_12033,N_15119);
and U21236 (N_21236,N_15390,N_12248);
nand U21237 (N_21237,N_14330,N_17895);
and U21238 (N_21238,N_13456,N_16371);
nor U21239 (N_21239,N_14273,N_14069);
nor U21240 (N_21240,N_13583,N_12128);
and U21241 (N_21241,N_15064,N_13996);
xor U21242 (N_21242,N_17038,N_17138);
xor U21243 (N_21243,N_16574,N_14751);
nor U21244 (N_21244,N_17083,N_12854);
or U21245 (N_21245,N_12356,N_13222);
or U21246 (N_21246,N_17975,N_17668);
nor U21247 (N_21247,N_17853,N_14888);
nor U21248 (N_21248,N_17152,N_13863);
and U21249 (N_21249,N_17205,N_12141);
and U21250 (N_21250,N_16154,N_12966);
and U21251 (N_21251,N_12611,N_15080);
xor U21252 (N_21252,N_13443,N_15035);
xnor U21253 (N_21253,N_14557,N_13465);
nand U21254 (N_21254,N_15332,N_17205);
or U21255 (N_21255,N_15045,N_14553);
xnor U21256 (N_21256,N_17197,N_14128);
nor U21257 (N_21257,N_16156,N_13630);
and U21258 (N_21258,N_12487,N_16182);
xor U21259 (N_21259,N_15521,N_16291);
nor U21260 (N_21260,N_17047,N_14522);
and U21261 (N_21261,N_12954,N_16455);
xor U21262 (N_21262,N_13380,N_14755);
xnor U21263 (N_21263,N_15465,N_14946);
xnor U21264 (N_21264,N_13183,N_16762);
nor U21265 (N_21265,N_16895,N_17204);
or U21266 (N_21266,N_12044,N_12423);
xnor U21267 (N_21267,N_12040,N_13917);
or U21268 (N_21268,N_15692,N_16910);
or U21269 (N_21269,N_14816,N_13883);
and U21270 (N_21270,N_17997,N_15993);
xnor U21271 (N_21271,N_15983,N_12241);
and U21272 (N_21272,N_16763,N_16706);
and U21273 (N_21273,N_17941,N_13926);
and U21274 (N_21274,N_16588,N_14336);
nand U21275 (N_21275,N_12281,N_17088);
and U21276 (N_21276,N_15466,N_13325);
xnor U21277 (N_21277,N_14034,N_16633);
nand U21278 (N_21278,N_16106,N_17988);
or U21279 (N_21279,N_16457,N_12933);
and U21280 (N_21280,N_13731,N_14027);
xor U21281 (N_21281,N_14784,N_16733);
xnor U21282 (N_21282,N_12656,N_17772);
nand U21283 (N_21283,N_14575,N_15563);
nor U21284 (N_21284,N_16676,N_15116);
nand U21285 (N_21285,N_17502,N_14052);
nand U21286 (N_21286,N_13630,N_17411);
or U21287 (N_21287,N_12907,N_16795);
nand U21288 (N_21288,N_15053,N_14275);
nor U21289 (N_21289,N_13786,N_13039);
or U21290 (N_21290,N_13242,N_13725);
or U21291 (N_21291,N_16645,N_17733);
or U21292 (N_21292,N_15720,N_12203);
nor U21293 (N_21293,N_16903,N_17281);
xor U21294 (N_21294,N_13686,N_12896);
nand U21295 (N_21295,N_15367,N_12901);
or U21296 (N_21296,N_15744,N_14470);
xnor U21297 (N_21297,N_16582,N_15172);
or U21298 (N_21298,N_13324,N_15796);
xnor U21299 (N_21299,N_16016,N_17977);
xor U21300 (N_21300,N_14163,N_12432);
nor U21301 (N_21301,N_12771,N_17394);
or U21302 (N_21302,N_12729,N_15501);
nand U21303 (N_21303,N_17850,N_16388);
nand U21304 (N_21304,N_15713,N_13422);
or U21305 (N_21305,N_15488,N_13130);
nand U21306 (N_21306,N_17435,N_12772);
xor U21307 (N_21307,N_17612,N_17531);
or U21308 (N_21308,N_16416,N_14726);
and U21309 (N_21309,N_12542,N_13529);
xnor U21310 (N_21310,N_13970,N_14747);
xor U21311 (N_21311,N_17043,N_13260);
and U21312 (N_21312,N_16181,N_17206);
nand U21313 (N_21313,N_17596,N_14781);
and U21314 (N_21314,N_16049,N_12494);
and U21315 (N_21315,N_17744,N_13900);
xnor U21316 (N_21316,N_15585,N_12373);
xor U21317 (N_21317,N_13979,N_12440);
nand U21318 (N_21318,N_14250,N_12096);
nor U21319 (N_21319,N_16757,N_13288);
nand U21320 (N_21320,N_14737,N_13473);
xor U21321 (N_21321,N_16911,N_14891);
or U21322 (N_21322,N_13584,N_17675);
or U21323 (N_21323,N_14688,N_14107);
nand U21324 (N_21324,N_12763,N_14167);
xor U21325 (N_21325,N_16699,N_17059);
or U21326 (N_21326,N_13202,N_13991);
and U21327 (N_21327,N_16437,N_15051);
xnor U21328 (N_21328,N_15352,N_17198);
nor U21329 (N_21329,N_16968,N_17856);
or U21330 (N_21330,N_12130,N_14720);
nand U21331 (N_21331,N_17884,N_13888);
nand U21332 (N_21332,N_12706,N_16027);
xnor U21333 (N_21333,N_12726,N_17090);
xnor U21334 (N_21334,N_15736,N_14594);
xor U21335 (N_21335,N_14733,N_14159);
xnor U21336 (N_21336,N_17555,N_12667);
xnor U21337 (N_21337,N_13598,N_17692);
xor U21338 (N_21338,N_13901,N_16208);
and U21339 (N_21339,N_12247,N_15357);
or U21340 (N_21340,N_17350,N_12658);
or U21341 (N_21341,N_17739,N_17664);
xnor U21342 (N_21342,N_17906,N_15468);
xnor U21343 (N_21343,N_15628,N_17587);
nand U21344 (N_21344,N_17894,N_17604);
nor U21345 (N_21345,N_14663,N_14037);
and U21346 (N_21346,N_15474,N_14088);
or U21347 (N_21347,N_17466,N_15407);
xor U21348 (N_21348,N_17947,N_14788);
nor U21349 (N_21349,N_16847,N_16127);
nand U21350 (N_21350,N_14273,N_14429);
and U21351 (N_21351,N_13669,N_13594);
and U21352 (N_21352,N_16587,N_16925);
xor U21353 (N_21353,N_15536,N_14673);
and U21354 (N_21354,N_17929,N_12057);
nor U21355 (N_21355,N_13882,N_13125);
nor U21356 (N_21356,N_13350,N_14606);
nand U21357 (N_21357,N_13781,N_12491);
or U21358 (N_21358,N_15115,N_12883);
or U21359 (N_21359,N_14703,N_13776);
and U21360 (N_21360,N_15771,N_16848);
nand U21361 (N_21361,N_12362,N_17361);
or U21362 (N_21362,N_14770,N_16726);
and U21363 (N_21363,N_16528,N_12326);
nor U21364 (N_21364,N_13016,N_13972);
or U21365 (N_21365,N_14323,N_12346);
or U21366 (N_21366,N_12768,N_12147);
or U21367 (N_21367,N_17516,N_15032);
or U21368 (N_21368,N_14205,N_12842);
or U21369 (N_21369,N_16191,N_17220);
and U21370 (N_21370,N_15529,N_15151);
and U21371 (N_21371,N_12419,N_14062);
and U21372 (N_21372,N_16558,N_15277);
or U21373 (N_21373,N_14826,N_15639);
and U21374 (N_21374,N_12502,N_15845);
xor U21375 (N_21375,N_13092,N_15415);
or U21376 (N_21376,N_14107,N_16104);
and U21377 (N_21377,N_12674,N_16039);
or U21378 (N_21378,N_14341,N_16236);
or U21379 (N_21379,N_12820,N_16946);
nand U21380 (N_21380,N_15792,N_13550);
and U21381 (N_21381,N_13025,N_13437);
nor U21382 (N_21382,N_16528,N_12242);
and U21383 (N_21383,N_17149,N_17281);
or U21384 (N_21384,N_15450,N_13652);
and U21385 (N_21385,N_15699,N_17431);
nand U21386 (N_21386,N_12705,N_13752);
nor U21387 (N_21387,N_15063,N_15954);
or U21388 (N_21388,N_16141,N_17089);
or U21389 (N_21389,N_17618,N_15227);
nor U21390 (N_21390,N_15559,N_15050);
nand U21391 (N_21391,N_17325,N_16748);
or U21392 (N_21392,N_16267,N_17649);
xor U21393 (N_21393,N_16575,N_12629);
nor U21394 (N_21394,N_17485,N_15630);
or U21395 (N_21395,N_16930,N_15140);
or U21396 (N_21396,N_14028,N_15947);
and U21397 (N_21397,N_16304,N_14583);
nand U21398 (N_21398,N_15946,N_15603);
nor U21399 (N_21399,N_12561,N_15798);
xnor U21400 (N_21400,N_13581,N_16631);
and U21401 (N_21401,N_12871,N_14966);
nand U21402 (N_21402,N_17288,N_17796);
xnor U21403 (N_21403,N_17716,N_12204);
nand U21404 (N_21404,N_16928,N_12187);
nor U21405 (N_21405,N_16861,N_13104);
nor U21406 (N_21406,N_13085,N_14971);
nor U21407 (N_21407,N_14551,N_14295);
xnor U21408 (N_21408,N_14121,N_12924);
and U21409 (N_21409,N_13869,N_17765);
xor U21410 (N_21410,N_17827,N_16115);
and U21411 (N_21411,N_16827,N_15261);
or U21412 (N_21412,N_12783,N_13607);
nand U21413 (N_21413,N_15520,N_14080);
nand U21414 (N_21414,N_16456,N_17926);
xor U21415 (N_21415,N_13676,N_15828);
or U21416 (N_21416,N_17185,N_14888);
nor U21417 (N_21417,N_16761,N_12154);
and U21418 (N_21418,N_15528,N_13917);
nor U21419 (N_21419,N_17309,N_14406);
xor U21420 (N_21420,N_12343,N_14901);
and U21421 (N_21421,N_15159,N_16339);
nor U21422 (N_21422,N_14189,N_17966);
or U21423 (N_21423,N_15739,N_16073);
nand U21424 (N_21424,N_12854,N_17591);
nor U21425 (N_21425,N_16799,N_15963);
or U21426 (N_21426,N_13678,N_16224);
xnor U21427 (N_21427,N_16900,N_17125);
nand U21428 (N_21428,N_14083,N_14674);
xnor U21429 (N_21429,N_17785,N_14378);
or U21430 (N_21430,N_14013,N_17059);
and U21431 (N_21431,N_13816,N_15017);
and U21432 (N_21432,N_13041,N_13396);
xor U21433 (N_21433,N_12779,N_12645);
and U21434 (N_21434,N_16072,N_13431);
nor U21435 (N_21435,N_12371,N_13216);
and U21436 (N_21436,N_17958,N_17002);
xnor U21437 (N_21437,N_14766,N_14939);
nand U21438 (N_21438,N_14171,N_17809);
nand U21439 (N_21439,N_16793,N_13476);
or U21440 (N_21440,N_15487,N_16382);
xor U21441 (N_21441,N_13475,N_12042);
nor U21442 (N_21442,N_15288,N_15690);
and U21443 (N_21443,N_16139,N_13546);
nand U21444 (N_21444,N_14408,N_16077);
nor U21445 (N_21445,N_15731,N_17015);
nor U21446 (N_21446,N_12168,N_17476);
nor U21447 (N_21447,N_12422,N_13109);
nor U21448 (N_21448,N_12156,N_13866);
xnor U21449 (N_21449,N_17682,N_12694);
xnor U21450 (N_21450,N_15306,N_17997);
and U21451 (N_21451,N_13235,N_17945);
and U21452 (N_21452,N_17428,N_13654);
nor U21453 (N_21453,N_16182,N_17798);
nand U21454 (N_21454,N_14448,N_16124);
and U21455 (N_21455,N_15288,N_17649);
and U21456 (N_21456,N_17588,N_17867);
xnor U21457 (N_21457,N_17073,N_13937);
and U21458 (N_21458,N_17989,N_14155);
nand U21459 (N_21459,N_14250,N_12547);
and U21460 (N_21460,N_16062,N_16956);
or U21461 (N_21461,N_15361,N_15997);
or U21462 (N_21462,N_16421,N_14691);
or U21463 (N_21463,N_13551,N_17351);
and U21464 (N_21464,N_13116,N_17658);
nor U21465 (N_21465,N_17290,N_16843);
or U21466 (N_21466,N_14233,N_14380);
nor U21467 (N_21467,N_15766,N_13370);
and U21468 (N_21468,N_16996,N_13353);
nand U21469 (N_21469,N_12076,N_12304);
nand U21470 (N_21470,N_16413,N_13818);
nand U21471 (N_21471,N_12301,N_15698);
nor U21472 (N_21472,N_17920,N_14528);
nor U21473 (N_21473,N_14057,N_12190);
or U21474 (N_21474,N_15696,N_13521);
xnor U21475 (N_21475,N_14182,N_17064);
nor U21476 (N_21476,N_12178,N_16257);
and U21477 (N_21477,N_15981,N_13775);
xnor U21478 (N_21478,N_16864,N_17717);
nor U21479 (N_21479,N_17534,N_17814);
nor U21480 (N_21480,N_16366,N_17299);
nand U21481 (N_21481,N_17464,N_17452);
nor U21482 (N_21482,N_15552,N_17395);
nor U21483 (N_21483,N_17761,N_13473);
or U21484 (N_21484,N_15197,N_14157);
xnor U21485 (N_21485,N_14722,N_14804);
or U21486 (N_21486,N_13777,N_15101);
or U21487 (N_21487,N_16356,N_13575);
nor U21488 (N_21488,N_16971,N_17738);
nor U21489 (N_21489,N_14610,N_12076);
nand U21490 (N_21490,N_17370,N_16432);
nand U21491 (N_21491,N_17734,N_15965);
nor U21492 (N_21492,N_13906,N_15068);
or U21493 (N_21493,N_13936,N_14069);
or U21494 (N_21494,N_16455,N_12763);
nor U21495 (N_21495,N_15878,N_13163);
and U21496 (N_21496,N_12704,N_12005);
or U21497 (N_21497,N_15883,N_17717);
nand U21498 (N_21498,N_13953,N_12342);
nand U21499 (N_21499,N_12781,N_13824);
or U21500 (N_21500,N_14954,N_15507);
and U21501 (N_21501,N_16745,N_13818);
nor U21502 (N_21502,N_16262,N_14705);
or U21503 (N_21503,N_12780,N_14747);
nand U21504 (N_21504,N_17360,N_17399);
and U21505 (N_21505,N_14827,N_17040);
nor U21506 (N_21506,N_12319,N_16162);
or U21507 (N_21507,N_14128,N_14463);
nand U21508 (N_21508,N_13112,N_17907);
or U21509 (N_21509,N_14015,N_17159);
xnor U21510 (N_21510,N_14127,N_13924);
or U21511 (N_21511,N_14039,N_12524);
and U21512 (N_21512,N_12537,N_13066);
and U21513 (N_21513,N_13365,N_12959);
and U21514 (N_21514,N_13430,N_16974);
or U21515 (N_21515,N_16730,N_14674);
and U21516 (N_21516,N_15702,N_17596);
nand U21517 (N_21517,N_13329,N_16426);
xor U21518 (N_21518,N_12509,N_13744);
xor U21519 (N_21519,N_17655,N_13329);
or U21520 (N_21520,N_13677,N_15146);
nor U21521 (N_21521,N_14948,N_12349);
or U21522 (N_21522,N_12269,N_14759);
nand U21523 (N_21523,N_14930,N_15295);
and U21524 (N_21524,N_12514,N_12374);
nand U21525 (N_21525,N_15570,N_17793);
or U21526 (N_21526,N_14181,N_13172);
or U21527 (N_21527,N_15570,N_14490);
and U21528 (N_21528,N_14047,N_12574);
nand U21529 (N_21529,N_14455,N_14411);
nand U21530 (N_21530,N_12513,N_17200);
and U21531 (N_21531,N_13560,N_13060);
xnor U21532 (N_21532,N_17312,N_16329);
and U21533 (N_21533,N_14391,N_14159);
nor U21534 (N_21534,N_14901,N_17364);
or U21535 (N_21535,N_12952,N_17115);
nand U21536 (N_21536,N_15355,N_15590);
or U21537 (N_21537,N_17208,N_13434);
nor U21538 (N_21538,N_16957,N_13370);
or U21539 (N_21539,N_14298,N_12509);
and U21540 (N_21540,N_16720,N_17968);
nand U21541 (N_21541,N_14625,N_16888);
xnor U21542 (N_21542,N_16415,N_12388);
nor U21543 (N_21543,N_17767,N_17473);
nand U21544 (N_21544,N_15942,N_14387);
xnor U21545 (N_21545,N_14159,N_12934);
xor U21546 (N_21546,N_16161,N_15291);
or U21547 (N_21547,N_14825,N_12676);
or U21548 (N_21548,N_12865,N_16569);
and U21549 (N_21549,N_17785,N_12385);
and U21550 (N_21550,N_17181,N_12397);
or U21551 (N_21551,N_16957,N_13511);
and U21552 (N_21552,N_15290,N_13090);
and U21553 (N_21553,N_17602,N_14471);
nor U21554 (N_21554,N_13310,N_16213);
and U21555 (N_21555,N_12341,N_16519);
nor U21556 (N_21556,N_16485,N_12060);
or U21557 (N_21557,N_12643,N_17727);
nand U21558 (N_21558,N_12155,N_13519);
or U21559 (N_21559,N_14031,N_16531);
or U21560 (N_21560,N_14647,N_12463);
nand U21561 (N_21561,N_12458,N_15095);
nor U21562 (N_21562,N_16623,N_17389);
or U21563 (N_21563,N_14639,N_15116);
nor U21564 (N_21564,N_13031,N_13178);
or U21565 (N_21565,N_15613,N_13461);
nor U21566 (N_21566,N_13450,N_14187);
xnor U21567 (N_21567,N_14892,N_16650);
xnor U21568 (N_21568,N_17678,N_14811);
and U21569 (N_21569,N_16552,N_13383);
and U21570 (N_21570,N_13156,N_13274);
or U21571 (N_21571,N_17942,N_16720);
xnor U21572 (N_21572,N_14238,N_14857);
and U21573 (N_21573,N_13789,N_16804);
or U21574 (N_21574,N_16125,N_14018);
nor U21575 (N_21575,N_17628,N_16446);
nand U21576 (N_21576,N_13130,N_14095);
and U21577 (N_21577,N_16947,N_15234);
and U21578 (N_21578,N_14442,N_16238);
nand U21579 (N_21579,N_12538,N_16389);
or U21580 (N_21580,N_17575,N_16829);
nand U21581 (N_21581,N_15451,N_15820);
xor U21582 (N_21582,N_17815,N_16766);
nor U21583 (N_21583,N_15621,N_13264);
and U21584 (N_21584,N_16822,N_16107);
or U21585 (N_21585,N_16746,N_14852);
xnor U21586 (N_21586,N_17886,N_14403);
xor U21587 (N_21587,N_17215,N_14544);
and U21588 (N_21588,N_16946,N_14299);
xor U21589 (N_21589,N_14149,N_14338);
nor U21590 (N_21590,N_14355,N_17010);
nor U21591 (N_21591,N_13380,N_13782);
xnor U21592 (N_21592,N_15738,N_17418);
nand U21593 (N_21593,N_17964,N_15146);
nand U21594 (N_21594,N_13384,N_14119);
nor U21595 (N_21595,N_17756,N_14818);
or U21596 (N_21596,N_15679,N_16181);
nor U21597 (N_21597,N_12334,N_13929);
nand U21598 (N_21598,N_16213,N_12163);
nand U21599 (N_21599,N_15524,N_15525);
xnor U21600 (N_21600,N_16946,N_12020);
and U21601 (N_21601,N_16615,N_13392);
nand U21602 (N_21602,N_16596,N_12253);
and U21603 (N_21603,N_15601,N_13513);
nand U21604 (N_21604,N_13690,N_17259);
nor U21605 (N_21605,N_13785,N_13662);
nor U21606 (N_21606,N_13872,N_14947);
nor U21607 (N_21607,N_12986,N_13254);
nand U21608 (N_21608,N_13489,N_14485);
nand U21609 (N_21609,N_14675,N_15678);
nor U21610 (N_21610,N_17135,N_14446);
xnor U21611 (N_21611,N_17011,N_17008);
nand U21612 (N_21612,N_12834,N_13487);
or U21613 (N_21613,N_15482,N_12740);
nand U21614 (N_21614,N_12664,N_13279);
nand U21615 (N_21615,N_17210,N_13324);
xor U21616 (N_21616,N_17477,N_17344);
or U21617 (N_21617,N_14734,N_13254);
and U21618 (N_21618,N_16168,N_12614);
xnor U21619 (N_21619,N_12050,N_17073);
and U21620 (N_21620,N_13367,N_13379);
or U21621 (N_21621,N_15792,N_15341);
nand U21622 (N_21622,N_14562,N_15366);
or U21623 (N_21623,N_12413,N_15914);
nand U21624 (N_21624,N_17564,N_14784);
xnor U21625 (N_21625,N_17238,N_15786);
nor U21626 (N_21626,N_17933,N_13704);
xor U21627 (N_21627,N_17551,N_15394);
nor U21628 (N_21628,N_16337,N_12548);
or U21629 (N_21629,N_17961,N_12247);
nand U21630 (N_21630,N_12216,N_15065);
nor U21631 (N_21631,N_14138,N_15580);
xor U21632 (N_21632,N_12104,N_13487);
nand U21633 (N_21633,N_14915,N_15558);
xor U21634 (N_21634,N_17055,N_12848);
nor U21635 (N_21635,N_13142,N_17969);
xnor U21636 (N_21636,N_12203,N_16616);
nand U21637 (N_21637,N_15965,N_17162);
xor U21638 (N_21638,N_12533,N_13665);
nor U21639 (N_21639,N_12427,N_17102);
or U21640 (N_21640,N_16957,N_14576);
or U21641 (N_21641,N_14861,N_13257);
and U21642 (N_21642,N_16756,N_13352);
or U21643 (N_21643,N_16071,N_12387);
nand U21644 (N_21644,N_13698,N_17432);
xnor U21645 (N_21645,N_13273,N_13396);
nor U21646 (N_21646,N_13867,N_14543);
and U21647 (N_21647,N_16293,N_13237);
nor U21648 (N_21648,N_15198,N_17020);
xor U21649 (N_21649,N_12750,N_17032);
nand U21650 (N_21650,N_17584,N_13101);
and U21651 (N_21651,N_16121,N_16034);
and U21652 (N_21652,N_17341,N_12593);
or U21653 (N_21653,N_14110,N_16137);
nand U21654 (N_21654,N_12927,N_17486);
nor U21655 (N_21655,N_15753,N_13695);
or U21656 (N_21656,N_13954,N_16803);
nor U21657 (N_21657,N_13445,N_15543);
xnor U21658 (N_21658,N_17668,N_14294);
nand U21659 (N_21659,N_12590,N_14557);
or U21660 (N_21660,N_14657,N_14540);
and U21661 (N_21661,N_12628,N_15721);
or U21662 (N_21662,N_12090,N_16561);
and U21663 (N_21663,N_15474,N_13697);
xor U21664 (N_21664,N_15733,N_14451);
nor U21665 (N_21665,N_15347,N_13121);
or U21666 (N_21666,N_12747,N_13176);
and U21667 (N_21667,N_14240,N_14386);
nand U21668 (N_21668,N_17290,N_16848);
xor U21669 (N_21669,N_12049,N_15349);
xor U21670 (N_21670,N_15257,N_12650);
and U21671 (N_21671,N_15314,N_17972);
nor U21672 (N_21672,N_15206,N_16600);
nor U21673 (N_21673,N_12599,N_17429);
nor U21674 (N_21674,N_15596,N_17866);
nand U21675 (N_21675,N_12276,N_17614);
or U21676 (N_21676,N_16191,N_12669);
and U21677 (N_21677,N_14301,N_17838);
xnor U21678 (N_21678,N_12711,N_14106);
xnor U21679 (N_21679,N_17205,N_13775);
or U21680 (N_21680,N_12865,N_15050);
xor U21681 (N_21681,N_15911,N_12176);
and U21682 (N_21682,N_16447,N_14288);
nand U21683 (N_21683,N_14437,N_15029);
and U21684 (N_21684,N_15029,N_12890);
and U21685 (N_21685,N_12423,N_12264);
nand U21686 (N_21686,N_12345,N_12395);
and U21687 (N_21687,N_14142,N_15539);
xnor U21688 (N_21688,N_15794,N_15820);
nand U21689 (N_21689,N_12034,N_12791);
or U21690 (N_21690,N_15955,N_14855);
and U21691 (N_21691,N_17458,N_13336);
xnor U21692 (N_21692,N_13880,N_17923);
nor U21693 (N_21693,N_17362,N_17531);
and U21694 (N_21694,N_12773,N_17166);
xor U21695 (N_21695,N_15094,N_17616);
or U21696 (N_21696,N_16621,N_14410);
or U21697 (N_21697,N_17566,N_13015);
nand U21698 (N_21698,N_13867,N_13520);
nand U21699 (N_21699,N_13622,N_17978);
nor U21700 (N_21700,N_15333,N_16234);
or U21701 (N_21701,N_16677,N_15730);
and U21702 (N_21702,N_15095,N_14258);
xor U21703 (N_21703,N_17234,N_16211);
and U21704 (N_21704,N_16267,N_17500);
xor U21705 (N_21705,N_16820,N_15451);
or U21706 (N_21706,N_13920,N_15407);
nor U21707 (N_21707,N_12125,N_13786);
xnor U21708 (N_21708,N_16738,N_15176);
xnor U21709 (N_21709,N_17675,N_12801);
or U21710 (N_21710,N_13739,N_12412);
nand U21711 (N_21711,N_13879,N_16362);
or U21712 (N_21712,N_15090,N_17573);
nor U21713 (N_21713,N_14014,N_12116);
xor U21714 (N_21714,N_15472,N_13229);
and U21715 (N_21715,N_16262,N_15054);
nand U21716 (N_21716,N_12827,N_12293);
nor U21717 (N_21717,N_15958,N_13886);
nor U21718 (N_21718,N_17369,N_15035);
nor U21719 (N_21719,N_14695,N_14988);
nand U21720 (N_21720,N_13169,N_14261);
nand U21721 (N_21721,N_16282,N_14130);
and U21722 (N_21722,N_12870,N_16664);
nand U21723 (N_21723,N_16083,N_14493);
nor U21724 (N_21724,N_14889,N_15447);
nand U21725 (N_21725,N_17639,N_17925);
or U21726 (N_21726,N_12214,N_17316);
nor U21727 (N_21727,N_15468,N_13295);
nand U21728 (N_21728,N_14387,N_13592);
or U21729 (N_21729,N_15481,N_14341);
xor U21730 (N_21730,N_13812,N_17343);
xnor U21731 (N_21731,N_17381,N_14674);
or U21732 (N_21732,N_12397,N_15835);
and U21733 (N_21733,N_13158,N_14190);
or U21734 (N_21734,N_15476,N_17820);
and U21735 (N_21735,N_17874,N_14552);
nor U21736 (N_21736,N_17711,N_13301);
and U21737 (N_21737,N_17635,N_15404);
nand U21738 (N_21738,N_17199,N_14088);
nand U21739 (N_21739,N_12676,N_16579);
nand U21740 (N_21740,N_14822,N_17257);
nor U21741 (N_21741,N_15263,N_12609);
and U21742 (N_21742,N_13211,N_16657);
or U21743 (N_21743,N_16636,N_15673);
xor U21744 (N_21744,N_17066,N_13038);
xor U21745 (N_21745,N_12484,N_14155);
xnor U21746 (N_21746,N_17851,N_12208);
nor U21747 (N_21747,N_17898,N_15144);
xnor U21748 (N_21748,N_16798,N_17232);
nand U21749 (N_21749,N_15059,N_17125);
nor U21750 (N_21750,N_14329,N_17187);
or U21751 (N_21751,N_12117,N_15726);
nand U21752 (N_21752,N_15820,N_17967);
or U21753 (N_21753,N_15143,N_12164);
xor U21754 (N_21754,N_16160,N_15550);
and U21755 (N_21755,N_16007,N_16607);
nand U21756 (N_21756,N_13654,N_12254);
and U21757 (N_21757,N_13396,N_14022);
or U21758 (N_21758,N_14997,N_16911);
nor U21759 (N_21759,N_17212,N_13239);
and U21760 (N_21760,N_15639,N_16617);
nor U21761 (N_21761,N_16685,N_15516);
nor U21762 (N_21762,N_17902,N_13235);
and U21763 (N_21763,N_15914,N_17016);
nor U21764 (N_21764,N_16036,N_15738);
nand U21765 (N_21765,N_17873,N_13938);
and U21766 (N_21766,N_16834,N_16984);
and U21767 (N_21767,N_15054,N_15425);
xor U21768 (N_21768,N_13605,N_12675);
or U21769 (N_21769,N_13201,N_15063);
or U21770 (N_21770,N_17637,N_15948);
nor U21771 (N_21771,N_15161,N_16562);
nand U21772 (N_21772,N_15347,N_12187);
and U21773 (N_21773,N_16991,N_13528);
xnor U21774 (N_21774,N_13574,N_13973);
nand U21775 (N_21775,N_17888,N_16675);
xor U21776 (N_21776,N_15856,N_13051);
and U21777 (N_21777,N_14964,N_16511);
nor U21778 (N_21778,N_16970,N_17593);
nand U21779 (N_21779,N_13037,N_17041);
nand U21780 (N_21780,N_15159,N_13524);
xnor U21781 (N_21781,N_15326,N_17640);
nor U21782 (N_21782,N_15852,N_12863);
nand U21783 (N_21783,N_16889,N_17366);
xor U21784 (N_21784,N_17618,N_15895);
nand U21785 (N_21785,N_17950,N_17927);
nor U21786 (N_21786,N_17891,N_15114);
xor U21787 (N_21787,N_16326,N_12935);
and U21788 (N_21788,N_17517,N_15423);
nor U21789 (N_21789,N_14822,N_15025);
xnor U21790 (N_21790,N_14969,N_12720);
nand U21791 (N_21791,N_13029,N_17340);
xor U21792 (N_21792,N_16284,N_15160);
nor U21793 (N_21793,N_17982,N_14289);
xnor U21794 (N_21794,N_14909,N_12609);
xor U21795 (N_21795,N_16636,N_13378);
and U21796 (N_21796,N_15192,N_14923);
or U21797 (N_21797,N_12310,N_16199);
or U21798 (N_21798,N_13378,N_12053);
and U21799 (N_21799,N_13675,N_17616);
nand U21800 (N_21800,N_13001,N_17807);
and U21801 (N_21801,N_12490,N_12290);
nand U21802 (N_21802,N_12896,N_13504);
or U21803 (N_21803,N_12630,N_12207);
nand U21804 (N_21804,N_17585,N_14554);
nor U21805 (N_21805,N_17995,N_16355);
xor U21806 (N_21806,N_16669,N_13482);
xnor U21807 (N_21807,N_13266,N_17439);
xnor U21808 (N_21808,N_17433,N_13718);
nor U21809 (N_21809,N_12587,N_15067);
nand U21810 (N_21810,N_13889,N_14041);
nand U21811 (N_21811,N_12140,N_14280);
and U21812 (N_21812,N_12506,N_16849);
nand U21813 (N_21813,N_15643,N_14700);
or U21814 (N_21814,N_13974,N_17340);
and U21815 (N_21815,N_15723,N_17362);
nor U21816 (N_21816,N_16738,N_17552);
or U21817 (N_21817,N_13777,N_17935);
xor U21818 (N_21818,N_15399,N_14593);
nor U21819 (N_21819,N_14599,N_15720);
nand U21820 (N_21820,N_12574,N_14304);
or U21821 (N_21821,N_16804,N_15533);
or U21822 (N_21822,N_14897,N_15203);
nor U21823 (N_21823,N_14097,N_16511);
xor U21824 (N_21824,N_12257,N_15810);
nand U21825 (N_21825,N_17065,N_14563);
or U21826 (N_21826,N_12163,N_16421);
nand U21827 (N_21827,N_12791,N_15602);
nor U21828 (N_21828,N_16192,N_13975);
nand U21829 (N_21829,N_14512,N_17854);
or U21830 (N_21830,N_12305,N_13329);
nand U21831 (N_21831,N_12744,N_16961);
xor U21832 (N_21832,N_16302,N_14487);
nor U21833 (N_21833,N_17977,N_12046);
and U21834 (N_21834,N_14017,N_14253);
nand U21835 (N_21835,N_14768,N_14783);
nor U21836 (N_21836,N_13180,N_12366);
nand U21837 (N_21837,N_14342,N_13296);
nor U21838 (N_21838,N_13440,N_12775);
nand U21839 (N_21839,N_13988,N_12275);
and U21840 (N_21840,N_14605,N_16228);
xnor U21841 (N_21841,N_14263,N_13871);
and U21842 (N_21842,N_16652,N_17491);
xnor U21843 (N_21843,N_12624,N_15639);
or U21844 (N_21844,N_16009,N_17777);
nand U21845 (N_21845,N_12520,N_12000);
nor U21846 (N_21846,N_16264,N_13873);
or U21847 (N_21847,N_13980,N_17462);
or U21848 (N_21848,N_15196,N_15143);
nor U21849 (N_21849,N_14222,N_17719);
nand U21850 (N_21850,N_12243,N_16103);
xnor U21851 (N_21851,N_15300,N_12923);
and U21852 (N_21852,N_15613,N_12648);
xor U21853 (N_21853,N_15078,N_14250);
and U21854 (N_21854,N_16528,N_17421);
or U21855 (N_21855,N_16870,N_17452);
nand U21856 (N_21856,N_16393,N_17068);
and U21857 (N_21857,N_13259,N_14412);
or U21858 (N_21858,N_15834,N_12778);
or U21859 (N_21859,N_15666,N_15282);
xnor U21860 (N_21860,N_15136,N_13697);
nor U21861 (N_21861,N_12555,N_14248);
and U21862 (N_21862,N_16416,N_17536);
nand U21863 (N_21863,N_14694,N_13692);
xor U21864 (N_21864,N_16117,N_17612);
xnor U21865 (N_21865,N_15409,N_16814);
nand U21866 (N_21866,N_16389,N_12935);
nand U21867 (N_21867,N_17867,N_15892);
nand U21868 (N_21868,N_13141,N_12038);
nand U21869 (N_21869,N_13293,N_17485);
nor U21870 (N_21870,N_17657,N_16496);
xor U21871 (N_21871,N_14270,N_16310);
xnor U21872 (N_21872,N_17700,N_17142);
or U21873 (N_21873,N_16333,N_12290);
and U21874 (N_21874,N_12775,N_14284);
or U21875 (N_21875,N_15330,N_12880);
xnor U21876 (N_21876,N_13998,N_15018);
xor U21877 (N_21877,N_17732,N_17822);
and U21878 (N_21878,N_15252,N_12116);
nand U21879 (N_21879,N_13267,N_12198);
nand U21880 (N_21880,N_17723,N_13586);
or U21881 (N_21881,N_15444,N_12303);
or U21882 (N_21882,N_12825,N_17255);
nor U21883 (N_21883,N_17029,N_16155);
nand U21884 (N_21884,N_14904,N_13083);
or U21885 (N_21885,N_14379,N_17183);
nand U21886 (N_21886,N_15453,N_17373);
xnor U21887 (N_21887,N_12158,N_12231);
xor U21888 (N_21888,N_17856,N_14353);
nor U21889 (N_21889,N_14319,N_15893);
or U21890 (N_21890,N_17095,N_16713);
nor U21891 (N_21891,N_13741,N_16902);
and U21892 (N_21892,N_12990,N_17995);
nand U21893 (N_21893,N_17469,N_15253);
and U21894 (N_21894,N_12818,N_14591);
and U21895 (N_21895,N_14950,N_14236);
and U21896 (N_21896,N_16254,N_14113);
or U21897 (N_21897,N_17211,N_12615);
or U21898 (N_21898,N_16597,N_12196);
xor U21899 (N_21899,N_13727,N_14323);
and U21900 (N_21900,N_14406,N_14318);
nor U21901 (N_21901,N_13982,N_17373);
nor U21902 (N_21902,N_12280,N_17722);
nand U21903 (N_21903,N_14139,N_15325);
or U21904 (N_21904,N_13081,N_13131);
xnor U21905 (N_21905,N_14080,N_12199);
and U21906 (N_21906,N_14316,N_16560);
xor U21907 (N_21907,N_15606,N_15651);
nand U21908 (N_21908,N_17228,N_14915);
nand U21909 (N_21909,N_14063,N_15601);
or U21910 (N_21910,N_12147,N_17586);
and U21911 (N_21911,N_12573,N_13193);
nand U21912 (N_21912,N_14749,N_17171);
nand U21913 (N_21913,N_14357,N_13493);
nand U21914 (N_21914,N_13054,N_12070);
nand U21915 (N_21915,N_14136,N_16365);
xor U21916 (N_21916,N_12733,N_16646);
or U21917 (N_21917,N_14160,N_17739);
xor U21918 (N_21918,N_14193,N_15279);
nand U21919 (N_21919,N_16996,N_17238);
xnor U21920 (N_21920,N_17722,N_15436);
nor U21921 (N_21921,N_12161,N_17510);
xor U21922 (N_21922,N_16437,N_14454);
nand U21923 (N_21923,N_12289,N_12203);
and U21924 (N_21924,N_15634,N_16598);
xor U21925 (N_21925,N_13832,N_12578);
xnor U21926 (N_21926,N_13115,N_15746);
nor U21927 (N_21927,N_17280,N_13833);
nand U21928 (N_21928,N_13598,N_13258);
or U21929 (N_21929,N_12654,N_16250);
or U21930 (N_21930,N_16732,N_16689);
nand U21931 (N_21931,N_16525,N_15110);
nor U21932 (N_21932,N_13690,N_13655);
nand U21933 (N_21933,N_15797,N_17612);
and U21934 (N_21934,N_13311,N_16500);
or U21935 (N_21935,N_15356,N_15890);
and U21936 (N_21936,N_15244,N_12891);
and U21937 (N_21937,N_14183,N_12202);
nand U21938 (N_21938,N_16087,N_16420);
nor U21939 (N_21939,N_14243,N_13518);
nor U21940 (N_21940,N_13009,N_13129);
or U21941 (N_21941,N_12096,N_16324);
xnor U21942 (N_21942,N_13426,N_15487);
and U21943 (N_21943,N_13480,N_17130);
xor U21944 (N_21944,N_16327,N_16474);
nor U21945 (N_21945,N_16908,N_12123);
nor U21946 (N_21946,N_14983,N_17748);
nand U21947 (N_21947,N_13064,N_13737);
nor U21948 (N_21948,N_17866,N_12977);
and U21949 (N_21949,N_17978,N_16486);
or U21950 (N_21950,N_17769,N_17429);
nor U21951 (N_21951,N_15777,N_13763);
or U21952 (N_21952,N_17949,N_17699);
and U21953 (N_21953,N_17985,N_13333);
or U21954 (N_21954,N_17520,N_17583);
nor U21955 (N_21955,N_14286,N_15435);
xnor U21956 (N_21956,N_16822,N_17146);
nand U21957 (N_21957,N_15279,N_15401);
xnor U21958 (N_21958,N_15780,N_16187);
xor U21959 (N_21959,N_17632,N_13428);
or U21960 (N_21960,N_12073,N_12017);
or U21961 (N_21961,N_13418,N_12598);
and U21962 (N_21962,N_12312,N_17986);
or U21963 (N_21963,N_16920,N_12599);
or U21964 (N_21964,N_17734,N_15477);
and U21965 (N_21965,N_17889,N_14952);
nor U21966 (N_21966,N_15725,N_16757);
and U21967 (N_21967,N_16343,N_16592);
nor U21968 (N_21968,N_14147,N_17647);
xnor U21969 (N_21969,N_16535,N_17903);
nand U21970 (N_21970,N_12440,N_16424);
and U21971 (N_21971,N_16747,N_17978);
nand U21972 (N_21972,N_13635,N_16376);
nand U21973 (N_21973,N_17193,N_16852);
and U21974 (N_21974,N_12016,N_17553);
or U21975 (N_21975,N_14935,N_14211);
nor U21976 (N_21976,N_16560,N_15401);
and U21977 (N_21977,N_16744,N_16003);
xnor U21978 (N_21978,N_17544,N_16953);
and U21979 (N_21979,N_17829,N_14859);
xor U21980 (N_21980,N_17085,N_16284);
or U21981 (N_21981,N_17275,N_17133);
and U21982 (N_21982,N_17586,N_16009);
or U21983 (N_21983,N_12644,N_12344);
nand U21984 (N_21984,N_15774,N_12428);
or U21985 (N_21985,N_17286,N_16926);
or U21986 (N_21986,N_14613,N_16445);
nor U21987 (N_21987,N_12008,N_13169);
nor U21988 (N_21988,N_16806,N_15395);
or U21989 (N_21989,N_16992,N_16137);
nand U21990 (N_21990,N_16661,N_14671);
and U21991 (N_21991,N_17468,N_13713);
nand U21992 (N_21992,N_15744,N_12885);
nor U21993 (N_21993,N_13252,N_13710);
xor U21994 (N_21994,N_12688,N_14850);
xnor U21995 (N_21995,N_17182,N_16037);
nand U21996 (N_21996,N_17940,N_16872);
or U21997 (N_21997,N_16588,N_12624);
nor U21998 (N_21998,N_12980,N_15594);
xnor U21999 (N_21999,N_15491,N_16272);
and U22000 (N_22000,N_13829,N_17832);
nor U22001 (N_22001,N_16125,N_12024);
nor U22002 (N_22002,N_15825,N_14681);
nand U22003 (N_22003,N_14876,N_13572);
xnor U22004 (N_22004,N_12142,N_12805);
or U22005 (N_22005,N_12810,N_14317);
and U22006 (N_22006,N_17630,N_16833);
and U22007 (N_22007,N_17661,N_16094);
nor U22008 (N_22008,N_12773,N_15555);
or U22009 (N_22009,N_14496,N_12041);
nand U22010 (N_22010,N_12400,N_16106);
xnor U22011 (N_22011,N_13473,N_14254);
nand U22012 (N_22012,N_14775,N_14365);
or U22013 (N_22013,N_13326,N_12697);
nor U22014 (N_22014,N_13640,N_17012);
and U22015 (N_22015,N_15415,N_14293);
or U22016 (N_22016,N_15301,N_13513);
xor U22017 (N_22017,N_17059,N_12137);
or U22018 (N_22018,N_15550,N_13677);
nand U22019 (N_22019,N_12285,N_15136);
nand U22020 (N_22020,N_13820,N_14901);
and U22021 (N_22021,N_13652,N_14143);
nand U22022 (N_22022,N_16385,N_12892);
nor U22023 (N_22023,N_12548,N_16509);
or U22024 (N_22024,N_14395,N_14219);
nor U22025 (N_22025,N_13809,N_16582);
xnor U22026 (N_22026,N_17740,N_12502);
nand U22027 (N_22027,N_15859,N_12860);
xor U22028 (N_22028,N_14335,N_14137);
and U22029 (N_22029,N_15148,N_17908);
xor U22030 (N_22030,N_13582,N_14706);
nand U22031 (N_22031,N_13324,N_15566);
nor U22032 (N_22032,N_12615,N_13850);
xor U22033 (N_22033,N_16520,N_17741);
nand U22034 (N_22034,N_12430,N_16276);
or U22035 (N_22035,N_15953,N_16601);
or U22036 (N_22036,N_14736,N_14395);
or U22037 (N_22037,N_17744,N_13788);
and U22038 (N_22038,N_13203,N_14769);
nand U22039 (N_22039,N_12327,N_17068);
xor U22040 (N_22040,N_15026,N_17969);
nor U22041 (N_22041,N_17413,N_14542);
or U22042 (N_22042,N_15576,N_16798);
nand U22043 (N_22043,N_13862,N_13633);
nor U22044 (N_22044,N_16318,N_13582);
nand U22045 (N_22045,N_16501,N_16198);
xnor U22046 (N_22046,N_17581,N_17986);
xnor U22047 (N_22047,N_13743,N_14807);
nor U22048 (N_22048,N_17986,N_16525);
or U22049 (N_22049,N_16929,N_13093);
and U22050 (N_22050,N_17435,N_17116);
nor U22051 (N_22051,N_14821,N_15294);
xor U22052 (N_22052,N_14892,N_13015);
and U22053 (N_22053,N_17925,N_15734);
or U22054 (N_22054,N_17308,N_13472);
nand U22055 (N_22055,N_14019,N_16117);
and U22056 (N_22056,N_14315,N_13099);
nand U22057 (N_22057,N_17490,N_12097);
nor U22058 (N_22058,N_14241,N_12263);
nor U22059 (N_22059,N_13690,N_15260);
and U22060 (N_22060,N_14258,N_14982);
and U22061 (N_22061,N_16403,N_13096);
or U22062 (N_22062,N_13381,N_14903);
or U22063 (N_22063,N_12983,N_12293);
and U22064 (N_22064,N_17476,N_14221);
and U22065 (N_22065,N_14254,N_16293);
xor U22066 (N_22066,N_12085,N_13852);
nor U22067 (N_22067,N_12647,N_16488);
nor U22068 (N_22068,N_12891,N_16860);
nand U22069 (N_22069,N_12287,N_14847);
xor U22070 (N_22070,N_13024,N_16565);
nor U22071 (N_22071,N_13362,N_15394);
or U22072 (N_22072,N_15611,N_16894);
and U22073 (N_22073,N_16205,N_17877);
nand U22074 (N_22074,N_16319,N_14240);
and U22075 (N_22075,N_16843,N_12634);
or U22076 (N_22076,N_13409,N_17282);
nor U22077 (N_22077,N_14850,N_14931);
nand U22078 (N_22078,N_15017,N_15748);
and U22079 (N_22079,N_13490,N_17120);
xnor U22080 (N_22080,N_15582,N_14620);
or U22081 (N_22081,N_16015,N_17731);
nor U22082 (N_22082,N_15365,N_16661);
nor U22083 (N_22083,N_14671,N_14687);
nor U22084 (N_22084,N_16520,N_17822);
and U22085 (N_22085,N_13086,N_12829);
xor U22086 (N_22086,N_14952,N_14307);
nand U22087 (N_22087,N_16599,N_15957);
and U22088 (N_22088,N_16787,N_12191);
and U22089 (N_22089,N_15118,N_16366);
nor U22090 (N_22090,N_13571,N_15940);
or U22091 (N_22091,N_17514,N_16119);
xnor U22092 (N_22092,N_12610,N_15156);
or U22093 (N_22093,N_13846,N_14116);
or U22094 (N_22094,N_16342,N_13758);
or U22095 (N_22095,N_16071,N_17069);
nand U22096 (N_22096,N_12808,N_12073);
and U22097 (N_22097,N_14508,N_13744);
nor U22098 (N_22098,N_15408,N_13447);
and U22099 (N_22099,N_14784,N_12468);
and U22100 (N_22100,N_16584,N_12244);
nor U22101 (N_22101,N_14341,N_12185);
nand U22102 (N_22102,N_15558,N_14749);
and U22103 (N_22103,N_12735,N_16657);
nand U22104 (N_22104,N_15541,N_14048);
xor U22105 (N_22105,N_17505,N_16695);
xnor U22106 (N_22106,N_16464,N_17579);
nor U22107 (N_22107,N_13765,N_14798);
nor U22108 (N_22108,N_13235,N_12540);
nand U22109 (N_22109,N_17347,N_13806);
or U22110 (N_22110,N_15104,N_17905);
nand U22111 (N_22111,N_14912,N_15459);
nor U22112 (N_22112,N_14084,N_15871);
xor U22113 (N_22113,N_15036,N_17002);
nand U22114 (N_22114,N_12649,N_15280);
and U22115 (N_22115,N_15830,N_16464);
or U22116 (N_22116,N_12137,N_15537);
or U22117 (N_22117,N_17622,N_16669);
nor U22118 (N_22118,N_14828,N_12714);
nand U22119 (N_22119,N_13176,N_12545);
xnor U22120 (N_22120,N_13905,N_13461);
and U22121 (N_22121,N_15870,N_17240);
xor U22122 (N_22122,N_14734,N_15491);
nand U22123 (N_22123,N_17883,N_12211);
nor U22124 (N_22124,N_14249,N_16437);
nand U22125 (N_22125,N_14266,N_14287);
and U22126 (N_22126,N_13447,N_15891);
and U22127 (N_22127,N_15827,N_14632);
or U22128 (N_22128,N_17128,N_13069);
xnor U22129 (N_22129,N_15809,N_13119);
xnor U22130 (N_22130,N_14606,N_12554);
xor U22131 (N_22131,N_14584,N_14834);
nor U22132 (N_22132,N_15525,N_15893);
and U22133 (N_22133,N_12583,N_14639);
nand U22134 (N_22134,N_14192,N_12345);
or U22135 (N_22135,N_17689,N_17950);
xnor U22136 (N_22136,N_15268,N_14028);
nor U22137 (N_22137,N_12279,N_13938);
and U22138 (N_22138,N_12205,N_17782);
nor U22139 (N_22139,N_15602,N_17910);
xnor U22140 (N_22140,N_12587,N_14868);
xnor U22141 (N_22141,N_14421,N_17025);
and U22142 (N_22142,N_13235,N_14185);
nand U22143 (N_22143,N_17594,N_13219);
nand U22144 (N_22144,N_14166,N_17129);
nor U22145 (N_22145,N_14218,N_15423);
nand U22146 (N_22146,N_13838,N_15976);
or U22147 (N_22147,N_13443,N_16381);
or U22148 (N_22148,N_14620,N_16882);
xnor U22149 (N_22149,N_17631,N_12856);
xor U22150 (N_22150,N_13167,N_17957);
nor U22151 (N_22151,N_13151,N_14876);
xnor U22152 (N_22152,N_15151,N_17020);
nor U22153 (N_22153,N_12310,N_13694);
xor U22154 (N_22154,N_17886,N_13831);
nor U22155 (N_22155,N_12980,N_12090);
nand U22156 (N_22156,N_16610,N_17856);
and U22157 (N_22157,N_13383,N_13966);
and U22158 (N_22158,N_12064,N_17712);
xnor U22159 (N_22159,N_12550,N_14089);
and U22160 (N_22160,N_16218,N_15697);
nand U22161 (N_22161,N_17729,N_14963);
and U22162 (N_22162,N_16204,N_17556);
and U22163 (N_22163,N_15728,N_14312);
nand U22164 (N_22164,N_17868,N_14017);
and U22165 (N_22165,N_15837,N_15769);
nor U22166 (N_22166,N_16451,N_13926);
nor U22167 (N_22167,N_14752,N_12563);
nor U22168 (N_22168,N_17382,N_17676);
nor U22169 (N_22169,N_13271,N_14539);
nor U22170 (N_22170,N_13309,N_12928);
nor U22171 (N_22171,N_15039,N_15827);
or U22172 (N_22172,N_13335,N_14125);
nand U22173 (N_22173,N_14330,N_12223);
or U22174 (N_22174,N_13261,N_15265);
nand U22175 (N_22175,N_12346,N_14553);
and U22176 (N_22176,N_14098,N_16240);
xnor U22177 (N_22177,N_15698,N_15153);
nor U22178 (N_22178,N_12573,N_16720);
nand U22179 (N_22179,N_17376,N_12940);
and U22180 (N_22180,N_14593,N_17408);
and U22181 (N_22181,N_17765,N_13238);
nand U22182 (N_22182,N_17282,N_17819);
or U22183 (N_22183,N_13906,N_13203);
or U22184 (N_22184,N_13469,N_12123);
and U22185 (N_22185,N_17912,N_12872);
or U22186 (N_22186,N_12254,N_15569);
and U22187 (N_22187,N_12713,N_17687);
or U22188 (N_22188,N_16033,N_12780);
and U22189 (N_22189,N_16100,N_16418);
nand U22190 (N_22190,N_14426,N_17015);
xnor U22191 (N_22191,N_13204,N_12739);
or U22192 (N_22192,N_14639,N_17442);
xor U22193 (N_22193,N_14526,N_13750);
xor U22194 (N_22194,N_16309,N_14422);
and U22195 (N_22195,N_14311,N_12839);
or U22196 (N_22196,N_16255,N_14085);
nor U22197 (N_22197,N_15327,N_14456);
and U22198 (N_22198,N_16931,N_13399);
xor U22199 (N_22199,N_15348,N_15122);
and U22200 (N_22200,N_15227,N_14911);
and U22201 (N_22201,N_14433,N_17472);
nor U22202 (N_22202,N_16770,N_15288);
xnor U22203 (N_22203,N_12922,N_14287);
xnor U22204 (N_22204,N_14884,N_14060);
nor U22205 (N_22205,N_14726,N_17024);
nand U22206 (N_22206,N_17393,N_15250);
and U22207 (N_22207,N_13639,N_12682);
or U22208 (N_22208,N_17930,N_14394);
or U22209 (N_22209,N_16723,N_13168);
xor U22210 (N_22210,N_12432,N_15104);
nand U22211 (N_22211,N_13573,N_15990);
or U22212 (N_22212,N_13153,N_14644);
nand U22213 (N_22213,N_12655,N_12970);
nor U22214 (N_22214,N_13718,N_13585);
xnor U22215 (N_22215,N_16757,N_13154);
nor U22216 (N_22216,N_16010,N_12540);
xor U22217 (N_22217,N_16728,N_12123);
nor U22218 (N_22218,N_15168,N_16572);
and U22219 (N_22219,N_15710,N_17274);
or U22220 (N_22220,N_16861,N_15490);
xor U22221 (N_22221,N_15357,N_14679);
and U22222 (N_22222,N_14422,N_15100);
nor U22223 (N_22223,N_13018,N_14256);
xnor U22224 (N_22224,N_16071,N_17576);
or U22225 (N_22225,N_13118,N_17765);
or U22226 (N_22226,N_14865,N_16260);
nand U22227 (N_22227,N_15538,N_14560);
xor U22228 (N_22228,N_15141,N_12416);
nor U22229 (N_22229,N_12074,N_16084);
and U22230 (N_22230,N_15922,N_13251);
or U22231 (N_22231,N_13038,N_16994);
nor U22232 (N_22232,N_14037,N_16322);
nand U22233 (N_22233,N_16686,N_16259);
nand U22234 (N_22234,N_17458,N_12664);
nand U22235 (N_22235,N_15877,N_16353);
or U22236 (N_22236,N_12426,N_13955);
and U22237 (N_22237,N_14154,N_12738);
xnor U22238 (N_22238,N_15292,N_13301);
and U22239 (N_22239,N_17017,N_13961);
or U22240 (N_22240,N_16619,N_13543);
nand U22241 (N_22241,N_13871,N_16807);
nand U22242 (N_22242,N_15098,N_12357);
xnor U22243 (N_22243,N_14526,N_12856);
nand U22244 (N_22244,N_14559,N_14007);
and U22245 (N_22245,N_14317,N_12128);
or U22246 (N_22246,N_17851,N_14836);
nand U22247 (N_22247,N_17441,N_14695);
xor U22248 (N_22248,N_14880,N_14652);
or U22249 (N_22249,N_12949,N_17490);
nand U22250 (N_22250,N_14909,N_14520);
nand U22251 (N_22251,N_16005,N_16135);
nand U22252 (N_22252,N_13036,N_12617);
nor U22253 (N_22253,N_14955,N_13034);
or U22254 (N_22254,N_16633,N_16378);
nand U22255 (N_22255,N_14468,N_17701);
xnor U22256 (N_22256,N_14690,N_15765);
xor U22257 (N_22257,N_17580,N_17409);
nand U22258 (N_22258,N_15031,N_17580);
xnor U22259 (N_22259,N_12048,N_15454);
and U22260 (N_22260,N_16591,N_17369);
xor U22261 (N_22261,N_16645,N_15992);
nand U22262 (N_22262,N_14773,N_16968);
nor U22263 (N_22263,N_12694,N_17668);
nor U22264 (N_22264,N_16975,N_15772);
and U22265 (N_22265,N_13064,N_13532);
nor U22266 (N_22266,N_16349,N_14432);
or U22267 (N_22267,N_12218,N_17768);
and U22268 (N_22268,N_17723,N_17678);
and U22269 (N_22269,N_12054,N_12216);
and U22270 (N_22270,N_12979,N_16736);
and U22271 (N_22271,N_13284,N_13795);
nand U22272 (N_22272,N_15215,N_17693);
nor U22273 (N_22273,N_16418,N_12857);
and U22274 (N_22274,N_17123,N_17587);
or U22275 (N_22275,N_13879,N_16290);
nor U22276 (N_22276,N_13678,N_16235);
xnor U22277 (N_22277,N_12704,N_13675);
nand U22278 (N_22278,N_16953,N_17539);
or U22279 (N_22279,N_15727,N_17133);
and U22280 (N_22280,N_12506,N_13328);
or U22281 (N_22281,N_14950,N_14778);
nor U22282 (N_22282,N_13143,N_15538);
xor U22283 (N_22283,N_14381,N_17220);
nor U22284 (N_22284,N_17592,N_12365);
or U22285 (N_22285,N_14677,N_17259);
and U22286 (N_22286,N_16528,N_16087);
xnor U22287 (N_22287,N_15090,N_13384);
xor U22288 (N_22288,N_13001,N_15349);
nor U22289 (N_22289,N_14681,N_13499);
xnor U22290 (N_22290,N_14270,N_14335);
xor U22291 (N_22291,N_15565,N_13366);
xnor U22292 (N_22292,N_12594,N_12332);
nand U22293 (N_22293,N_17587,N_14929);
nand U22294 (N_22294,N_15936,N_16281);
xnor U22295 (N_22295,N_14171,N_14514);
xor U22296 (N_22296,N_13111,N_15917);
xnor U22297 (N_22297,N_16471,N_12099);
or U22298 (N_22298,N_13545,N_13136);
xor U22299 (N_22299,N_17885,N_13742);
nand U22300 (N_22300,N_14650,N_17143);
and U22301 (N_22301,N_12459,N_12760);
or U22302 (N_22302,N_13764,N_17736);
and U22303 (N_22303,N_16485,N_13739);
nand U22304 (N_22304,N_14958,N_17983);
xnor U22305 (N_22305,N_14702,N_16359);
and U22306 (N_22306,N_13055,N_12373);
xor U22307 (N_22307,N_14884,N_16255);
nor U22308 (N_22308,N_12828,N_17066);
nor U22309 (N_22309,N_16894,N_16223);
xnor U22310 (N_22310,N_14170,N_13012);
xor U22311 (N_22311,N_15216,N_12114);
xnor U22312 (N_22312,N_13539,N_12014);
and U22313 (N_22313,N_13779,N_15502);
nand U22314 (N_22314,N_12793,N_12189);
nand U22315 (N_22315,N_14619,N_17653);
xor U22316 (N_22316,N_16942,N_13373);
nor U22317 (N_22317,N_16277,N_15138);
xnor U22318 (N_22318,N_13175,N_13718);
nor U22319 (N_22319,N_16696,N_12370);
nor U22320 (N_22320,N_15448,N_14737);
nor U22321 (N_22321,N_14111,N_13656);
nor U22322 (N_22322,N_13761,N_17323);
and U22323 (N_22323,N_16818,N_17763);
nor U22324 (N_22324,N_12891,N_12610);
or U22325 (N_22325,N_15787,N_14648);
nand U22326 (N_22326,N_14273,N_17265);
nor U22327 (N_22327,N_15336,N_17631);
or U22328 (N_22328,N_12277,N_13409);
and U22329 (N_22329,N_14385,N_14852);
and U22330 (N_22330,N_17366,N_14473);
and U22331 (N_22331,N_15637,N_13801);
xnor U22332 (N_22332,N_12120,N_14256);
nor U22333 (N_22333,N_17545,N_16866);
nand U22334 (N_22334,N_13135,N_15088);
and U22335 (N_22335,N_17697,N_15359);
or U22336 (N_22336,N_17943,N_13435);
nor U22337 (N_22337,N_14232,N_17195);
xnor U22338 (N_22338,N_13991,N_14909);
xor U22339 (N_22339,N_15919,N_17707);
nor U22340 (N_22340,N_12986,N_17641);
nor U22341 (N_22341,N_14974,N_12478);
and U22342 (N_22342,N_14808,N_17899);
or U22343 (N_22343,N_13498,N_15612);
nand U22344 (N_22344,N_12279,N_13592);
or U22345 (N_22345,N_14829,N_16722);
nor U22346 (N_22346,N_15750,N_13403);
nor U22347 (N_22347,N_13165,N_12297);
and U22348 (N_22348,N_12352,N_12526);
or U22349 (N_22349,N_13656,N_15411);
nand U22350 (N_22350,N_12681,N_14729);
nand U22351 (N_22351,N_15520,N_13546);
nor U22352 (N_22352,N_15391,N_13565);
nand U22353 (N_22353,N_12894,N_12119);
xnor U22354 (N_22354,N_12758,N_12263);
and U22355 (N_22355,N_14060,N_14585);
nand U22356 (N_22356,N_15437,N_14863);
and U22357 (N_22357,N_13224,N_17372);
and U22358 (N_22358,N_16327,N_12727);
and U22359 (N_22359,N_12457,N_13048);
or U22360 (N_22360,N_17023,N_13374);
and U22361 (N_22361,N_15597,N_14339);
nand U22362 (N_22362,N_14010,N_14497);
nor U22363 (N_22363,N_14922,N_16795);
nand U22364 (N_22364,N_12023,N_12345);
nand U22365 (N_22365,N_15152,N_14107);
xor U22366 (N_22366,N_16848,N_13266);
and U22367 (N_22367,N_14383,N_13718);
xor U22368 (N_22368,N_15106,N_17125);
nor U22369 (N_22369,N_13721,N_15974);
nand U22370 (N_22370,N_14817,N_12859);
or U22371 (N_22371,N_12089,N_13577);
and U22372 (N_22372,N_12947,N_12567);
or U22373 (N_22373,N_17720,N_17747);
or U22374 (N_22374,N_17055,N_12847);
nand U22375 (N_22375,N_16390,N_14486);
and U22376 (N_22376,N_16003,N_14678);
xnor U22377 (N_22377,N_17270,N_15868);
and U22378 (N_22378,N_15563,N_15363);
and U22379 (N_22379,N_17738,N_17816);
and U22380 (N_22380,N_13731,N_17981);
and U22381 (N_22381,N_16748,N_13082);
and U22382 (N_22382,N_16995,N_12135);
or U22383 (N_22383,N_13025,N_17942);
nor U22384 (N_22384,N_17737,N_13928);
xor U22385 (N_22385,N_15805,N_15504);
nor U22386 (N_22386,N_13423,N_15799);
xor U22387 (N_22387,N_15450,N_16265);
nor U22388 (N_22388,N_14600,N_16594);
nor U22389 (N_22389,N_16795,N_16914);
nand U22390 (N_22390,N_12654,N_12384);
and U22391 (N_22391,N_17218,N_12966);
nor U22392 (N_22392,N_17780,N_16890);
and U22393 (N_22393,N_14394,N_15311);
nand U22394 (N_22394,N_13053,N_15375);
nor U22395 (N_22395,N_17098,N_15773);
nor U22396 (N_22396,N_16875,N_13532);
xor U22397 (N_22397,N_14561,N_14750);
or U22398 (N_22398,N_14706,N_12397);
nor U22399 (N_22399,N_12895,N_14160);
nor U22400 (N_22400,N_15645,N_13782);
nand U22401 (N_22401,N_13968,N_12082);
nor U22402 (N_22402,N_13925,N_14372);
or U22403 (N_22403,N_13491,N_16394);
nor U22404 (N_22404,N_14111,N_15757);
and U22405 (N_22405,N_12092,N_12122);
nor U22406 (N_22406,N_16312,N_16139);
nor U22407 (N_22407,N_15841,N_12212);
xnor U22408 (N_22408,N_12108,N_13878);
or U22409 (N_22409,N_14819,N_14332);
xor U22410 (N_22410,N_16415,N_16792);
or U22411 (N_22411,N_12979,N_12133);
and U22412 (N_22412,N_14416,N_16855);
nand U22413 (N_22413,N_12676,N_15420);
or U22414 (N_22414,N_16711,N_13318);
and U22415 (N_22415,N_14356,N_15099);
or U22416 (N_22416,N_13624,N_14748);
nor U22417 (N_22417,N_16083,N_13787);
xor U22418 (N_22418,N_14684,N_15368);
xnor U22419 (N_22419,N_13358,N_16254);
xnor U22420 (N_22420,N_17628,N_16321);
xor U22421 (N_22421,N_16223,N_14110);
and U22422 (N_22422,N_15974,N_17825);
or U22423 (N_22423,N_12388,N_17093);
xor U22424 (N_22424,N_14848,N_13463);
nor U22425 (N_22425,N_13361,N_16941);
or U22426 (N_22426,N_13006,N_16743);
nand U22427 (N_22427,N_15900,N_14865);
and U22428 (N_22428,N_15587,N_17451);
xor U22429 (N_22429,N_14308,N_14336);
nor U22430 (N_22430,N_14031,N_15456);
nand U22431 (N_22431,N_13467,N_17042);
or U22432 (N_22432,N_12689,N_13964);
xor U22433 (N_22433,N_14116,N_16720);
xor U22434 (N_22434,N_15179,N_17986);
nand U22435 (N_22435,N_12607,N_16950);
nand U22436 (N_22436,N_12483,N_13433);
and U22437 (N_22437,N_17971,N_13156);
nor U22438 (N_22438,N_13493,N_16016);
nand U22439 (N_22439,N_14417,N_16590);
and U22440 (N_22440,N_12247,N_14709);
or U22441 (N_22441,N_16471,N_17370);
nand U22442 (N_22442,N_16117,N_14374);
or U22443 (N_22443,N_12814,N_14986);
xnor U22444 (N_22444,N_13408,N_14036);
or U22445 (N_22445,N_12839,N_16893);
and U22446 (N_22446,N_14411,N_12028);
nand U22447 (N_22447,N_16696,N_15129);
xnor U22448 (N_22448,N_16539,N_16732);
nand U22449 (N_22449,N_14748,N_12309);
xnor U22450 (N_22450,N_12727,N_12794);
and U22451 (N_22451,N_15165,N_12345);
nor U22452 (N_22452,N_14646,N_16304);
or U22453 (N_22453,N_13452,N_13194);
and U22454 (N_22454,N_14776,N_13797);
or U22455 (N_22455,N_17903,N_12860);
or U22456 (N_22456,N_13931,N_14706);
xor U22457 (N_22457,N_14540,N_16527);
xor U22458 (N_22458,N_17516,N_16564);
nor U22459 (N_22459,N_13331,N_16852);
nand U22460 (N_22460,N_17670,N_13408);
or U22461 (N_22461,N_16345,N_13664);
nor U22462 (N_22462,N_16695,N_13305);
nor U22463 (N_22463,N_14836,N_13306);
nor U22464 (N_22464,N_16935,N_17938);
nor U22465 (N_22465,N_14246,N_16887);
and U22466 (N_22466,N_15623,N_15732);
xor U22467 (N_22467,N_14854,N_13106);
and U22468 (N_22468,N_12461,N_14058);
nor U22469 (N_22469,N_12992,N_16731);
and U22470 (N_22470,N_16407,N_15281);
and U22471 (N_22471,N_17592,N_14774);
and U22472 (N_22472,N_12500,N_16215);
and U22473 (N_22473,N_15828,N_15018);
nand U22474 (N_22474,N_17600,N_17378);
or U22475 (N_22475,N_13761,N_14165);
nand U22476 (N_22476,N_12820,N_17370);
nand U22477 (N_22477,N_13811,N_15547);
and U22478 (N_22478,N_16048,N_17912);
nand U22479 (N_22479,N_16665,N_15239);
xnor U22480 (N_22480,N_15607,N_14374);
or U22481 (N_22481,N_14206,N_14107);
xor U22482 (N_22482,N_14926,N_15929);
nand U22483 (N_22483,N_17316,N_14090);
and U22484 (N_22484,N_15463,N_12640);
nand U22485 (N_22485,N_16003,N_14161);
nor U22486 (N_22486,N_14588,N_17956);
or U22487 (N_22487,N_15699,N_12678);
nand U22488 (N_22488,N_16037,N_14497);
nand U22489 (N_22489,N_14114,N_15314);
and U22490 (N_22490,N_15647,N_12367);
or U22491 (N_22491,N_17299,N_12663);
xnor U22492 (N_22492,N_17400,N_17282);
or U22493 (N_22493,N_12666,N_16241);
xnor U22494 (N_22494,N_13308,N_14344);
xnor U22495 (N_22495,N_12619,N_14718);
nor U22496 (N_22496,N_13951,N_12538);
and U22497 (N_22497,N_17045,N_12661);
xor U22498 (N_22498,N_12469,N_12069);
xnor U22499 (N_22499,N_13866,N_16508);
xnor U22500 (N_22500,N_14181,N_16710);
and U22501 (N_22501,N_14607,N_16285);
nand U22502 (N_22502,N_13275,N_15763);
or U22503 (N_22503,N_12311,N_17400);
xnor U22504 (N_22504,N_15563,N_15855);
or U22505 (N_22505,N_12122,N_15871);
nor U22506 (N_22506,N_17186,N_14029);
xnor U22507 (N_22507,N_17266,N_16057);
xor U22508 (N_22508,N_16975,N_15008);
nand U22509 (N_22509,N_17717,N_15929);
or U22510 (N_22510,N_16593,N_14836);
xnor U22511 (N_22511,N_13147,N_15102);
and U22512 (N_22512,N_14220,N_17548);
and U22513 (N_22513,N_12224,N_15834);
nand U22514 (N_22514,N_16322,N_12684);
nor U22515 (N_22515,N_16220,N_17871);
xor U22516 (N_22516,N_12235,N_17173);
nand U22517 (N_22517,N_16257,N_17505);
and U22518 (N_22518,N_15034,N_12792);
nand U22519 (N_22519,N_16909,N_13470);
and U22520 (N_22520,N_15208,N_13228);
and U22521 (N_22521,N_17252,N_17414);
or U22522 (N_22522,N_17713,N_12366);
xnor U22523 (N_22523,N_12840,N_14964);
and U22524 (N_22524,N_17994,N_17747);
and U22525 (N_22525,N_16756,N_12430);
nor U22526 (N_22526,N_17578,N_17016);
nor U22527 (N_22527,N_14734,N_15153);
nand U22528 (N_22528,N_17485,N_12074);
nor U22529 (N_22529,N_15730,N_13639);
nor U22530 (N_22530,N_16884,N_16026);
xor U22531 (N_22531,N_17846,N_16500);
and U22532 (N_22532,N_15974,N_12239);
nor U22533 (N_22533,N_14289,N_17819);
or U22534 (N_22534,N_17355,N_14969);
nor U22535 (N_22535,N_12577,N_16198);
or U22536 (N_22536,N_13737,N_15440);
nor U22537 (N_22537,N_15011,N_14432);
nand U22538 (N_22538,N_14390,N_17232);
xnor U22539 (N_22539,N_14512,N_14218);
xor U22540 (N_22540,N_15486,N_12905);
and U22541 (N_22541,N_15071,N_17685);
and U22542 (N_22542,N_15563,N_13927);
nand U22543 (N_22543,N_15247,N_14538);
or U22544 (N_22544,N_13372,N_16021);
nand U22545 (N_22545,N_14115,N_12309);
nor U22546 (N_22546,N_17253,N_16312);
nor U22547 (N_22547,N_17565,N_17494);
nand U22548 (N_22548,N_17223,N_12265);
nand U22549 (N_22549,N_15919,N_13798);
xor U22550 (N_22550,N_15699,N_17948);
or U22551 (N_22551,N_15598,N_13124);
and U22552 (N_22552,N_12283,N_17869);
and U22553 (N_22553,N_12510,N_13427);
or U22554 (N_22554,N_13293,N_14246);
and U22555 (N_22555,N_15717,N_12541);
xnor U22556 (N_22556,N_12811,N_13149);
nand U22557 (N_22557,N_17847,N_14183);
or U22558 (N_22558,N_17762,N_17492);
xor U22559 (N_22559,N_14331,N_15651);
nand U22560 (N_22560,N_13695,N_12383);
nand U22561 (N_22561,N_17785,N_16209);
and U22562 (N_22562,N_12767,N_16380);
or U22563 (N_22563,N_17287,N_17096);
nand U22564 (N_22564,N_14859,N_15484);
or U22565 (N_22565,N_17634,N_16366);
xnor U22566 (N_22566,N_17124,N_15377);
and U22567 (N_22567,N_15114,N_17588);
nand U22568 (N_22568,N_12648,N_15274);
xnor U22569 (N_22569,N_14143,N_13025);
and U22570 (N_22570,N_12765,N_16674);
xnor U22571 (N_22571,N_15030,N_13305);
nand U22572 (N_22572,N_13751,N_12110);
nand U22573 (N_22573,N_16298,N_12157);
nor U22574 (N_22574,N_12582,N_17601);
or U22575 (N_22575,N_16504,N_14046);
or U22576 (N_22576,N_16797,N_17208);
nor U22577 (N_22577,N_13452,N_15133);
nand U22578 (N_22578,N_13523,N_13727);
xnor U22579 (N_22579,N_12337,N_12314);
xnor U22580 (N_22580,N_17678,N_16192);
xnor U22581 (N_22581,N_13413,N_16535);
and U22582 (N_22582,N_16072,N_14561);
and U22583 (N_22583,N_12274,N_16205);
and U22584 (N_22584,N_17442,N_13166);
xor U22585 (N_22585,N_15831,N_17499);
xnor U22586 (N_22586,N_13382,N_14753);
or U22587 (N_22587,N_13340,N_17157);
or U22588 (N_22588,N_14770,N_16244);
nor U22589 (N_22589,N_12148,N_16000);
and U22590 (N_22590,N_12757,N_13415);
nand U22591 (N_22591,N_15243,N_16367);
nor U22592 (N_22592,N_16475,N_12894);
and U22593 (N_22593,N_12369,N_13071);
xnor U22594 (N_22594,N_17901,N_14536);
nand U22595 (N_22595,N_12485,N_15010);
or U22596 (N_22596,N_17489,N_15137);
xnor U22597 (N_22597,N_14554,N_14492);
nand U22598 (N_22598,N_17403,N_17105);
or U22599 (N_22599,N_16285,N_12704);
nand U22600 (N_22600,N_13008,N_16977);
xnor U22601 (N_22601,N_15308,N_15776);
and U22602 (N_22602,N_15671,N_16125);
and U22603 (N_22603,N_13317,N_12070);
and U22604 (N_22604,N_15532,N_13320);
and U22605 (N_22605,N_15455,N_14377);
nor U22606 (N_22606,N_13353,N_13358);
nand U22607 (N_22607,N_14451,N_12124);
nor U22608 (N_22608,N_15134,N_15345);
xnor U22609 (N_22609,N_14759,N_17105);
or U22610 (N_22610,N_17181,N_17840);
and U22611 (N_22611,N_15198,N_16415);
nor U22612 (N_22612,N_13779,N_12166);
xor U22613 (N_22613,N_13709,N_16301);
nor U22614 (N_22614,N_16200,N_16232);
or U22615 (N_22615,N_16778,N_14503);
xor U22616 (N_22616,N_13240,N_16248);
nor U22617 (N_22617,N_16788,N_14966);
and U22618 (N_22618,N_13690,N_15679);
and U22619 (N_22619,N_16229,N_12946);
nand U22620 (N_22620,N_15961,N_17929);
and U22621 (N_22621,N_15869,N_17942);
nand U22622 (N_22622,N_16709,N_14398);
nor U22623 (N_22623,N_13021,N_12136);
xnor U22624 (N_22624,N_13182,N_17706);
or U22625 (N_22625,N_12086,N_17428);
xor U22626 (N_22626,N_14025,N_16067);
nor U22627 (N_22627,N_12428,N_15575);
xnor U22628 (N_22628,N_13133,N_16000);
and U22629 (N_22629,N_12470,N_17326);
nor U22630 (N_22630,N_15018,N_13862);
nor U22631 (N_22631,N_14608,N_12441);
and U22632 (N_22632,N_15630,N_15191);
xnor U22633 (N_22633,N_17442,N_14963);
xnor U22634 (N_22634,N_17425,N_16595);
xor U22635 (N_22635,N_17455,N_13578);
and U22636 (N_22636,N_14915,N_12997);
and U22637 (N_22637,N_16255,N_15932);
nand U22638 (N_22638,N_13272,N_12975);
and U22639 (N_22639,N_17066,N_16403);
and U22640 (N_22640,N_16371,N_12231);
or U22641 (N_22641,N_15993,N_17931);
nand U22642 (N_22642,N_13785,N_12427);
nor U22643 (N_22643,N_16839,N_17478);
or U22644 (N_22644,N_12436,N_16912);
nor U22645 (N_22645,N_14259,N_14614);
xor U22646 (N_22646,N_16746,N_16500);
nand U22647 (N_22647,N_13205,N_16134);
or U22648 (N_22648,N_17241,N_15486);
and U22649 (N_22649,N_13116,N_13457);
xor U22650 (N_22650,N_16702,N_15323);
nor U22651 (N_22651,N_17403,N_14123);
nor U22652 (N_22652,N_14865,N_12907);
nor U22653 (N_22653,N_13846,N_16060);
xor U22654 (N_22654,N_17488,N_17913);
or U22655 (N_22655,N_12544,N_12796);
nor U22656 (N_22656,N_16791,N_16749);
xor U22657 (N_22657,N_17964,N_15780);
nand U22658 (N_22658,N_16025,N_15809);
or U22659 (N_22659,N_13217,N_13208);
and U22660 (N_22660,N_17221,N_17129);
nor U22661 (N_22661,N_14104,N_15872);
xor U22662 (N_22662,N_12039,N_14278);
nor U22663 (N_22663,N_14938,N_17792);
nor U22664 (N_22664,N_13932,N_16981);
nor U22665 (N_22665,N_15611,N_14886);
and U22666 (N_22666,N_16664,N_15635);
or U22667 (N_22667,N_14882,N_15337);
nor U22668 (N_22668,N_13162,N_17241);
xnor U22669 (N_22669,N_12977,N_14091);
nand U22670 (N_22670,N_15697,N_14998);
and U22671 (N_22671,N_15608,N_17154);
nand U22672 (N_22672,N_13043,N_12008);
nand U22673 (N_22673,N_12619,N_14214);
nand U22674 (N_22674,N_14543,N_13398);
xor U22675 (N_22675,N_12538,N_16025);
and U22676 (N_22676,N_14944,N_17782);
or U22677 (N_22677,N_13499,N_13828);
and U22678 (N_22678,N_13721,N_14737);
or U22679 (N_22679,N_17651,N_13834);
nor U22680 (N_22680,N_12710,N_13527);
or U22681 (N_22681,N_13250,N_17090);
nor U22682 (N_22682,N_14942,N_15140);
nand U22683 (N_22683,N_16175,N_15836);
and U22684 (N_22684,N_14988,N_14511);
xnor U22685 (N_22685,N_17595,N_16975);
nand U22686 (N_22686,N_12375,N_12066);
and U22687 (N_22687,N_16996,N_17015);
or U22688 (N_22688,N_15696,N_15420);
nor U22689 (N_22689,N_12857,N_12090);
nor U22690 (N_22690,N_15876,N_17538);
nand U22691 (N_22691,N_12409,N_16210);
xor U22692 (N_22692,N_12525,N_14829);
xor U22693 (N_22693,N_17721,N_14224);
nand U22694 (N_22694,N_14471,N_15312);
nand U22695 (N_22695,N_12807,N_17142);
xnor U22696 (N_22696,N_14698,N_17269);
xnor U22697 (N_22697,N_17547,N_13508);
nand U22698 (N_22698,N_17970,N_13551);
xnor U22699 (N_22699,N_12681,N_16860);
xnor U22700 (N_22700,N_17565,N_13705);
or U22701 (N_22701,N_14424,N_16345);
nand U22702 (N_22702,N_14880,N_15109);
nand U22703 (N_22703,N_13354,N_14820);
nand U22704 (N_22704,N_12707,N_13636);
or U22705 (N_22705,N_12513,N_14836);
nor U22706 (N_22706,N_16554,N_13482);
nor U22707 (N_22707,N_12062,N_14350);
and U22708 (N_22708,N_13812,N_12535);
or U22709 (N_22709,N_13181,N_17251);
and U22710 (N_22710,N_17255,N_17333);
xnor U22711 (N_22711,N_15451,N_14773);
nor U22712 (N_22712,N_17005,N_16721);
nand U22713 (N_22713,N_15375,N_16527);
and U22714 (N_22714,N_17203,N_16214);
xor U22715 (N_22715,N_16171,N_13597);
nor U22716 (N_22716,N_14932,N_16884);
or U22717 (N_22717,N_12369,N_17832);
and U22718 (N_22718,N_17605,N_15367);
nand U22719 (N_22719,N_16791,N_17071);
and U22720 (N_22720,N_15090,N_14786);
nand U22721 (N_22721,N_12133,N_12911);
nor U22722 (N_22722,N_15803,N_15810);
xnor U22723 (N_22723,N_16924,N_14021);
or U22724 (N_22724,N_15907,N_17090);
nor U22725 (N_22725,N_14568,N_17930);
xor U22726 (N_22726,N_15068,N_14573);
xor U22727 (N_22727,N_15399,N_17857);
and U22728 (N_22728,N_13520,N_17673);
and U22729 (N_22729,N_14007,N_12959);
and U22730 (N_22730,N_13576,N_17242);
xnor U22731 (N_22731,N_16861,N_13303);
nor U22732 (N_22732,N_13317,N_17002);
xor U22733 (N_22733,N_14579,N_16711);
and U22734 (N_22734,N_16536,N_17532);
nand U22735 (N_22735,N_16490,N_16233);
nor U22736 (N_22736,N_14997,N_17347);
and U22737 (N_22737,N_16761,N_14129);
nor U22738 (N_22738,N_14093,N_14280);
nand U22739 (N_22739,N_17654,N_12941);
nand U22740 (N_22740,N_13679,N_15231);
or U22741 (N_22741,N_16862,N_14683);
xnor U22742 (N_22742,N_16487,N_15833);
or U22743 (N_22743,N_13133,N_15293);
and U22744 (N_22744,N_15903,N_17101);
nand U22745 (N_22745,N_12359,N_12923);
xnor U22746 (N_22746,N_15175,N_12136);
and U22747 (N_22747,N_15802,N_15239);
or U22748 (N_22748,N_15055,N_12832);
nor U22749 (N_22749,N_12016,N_15903);
and U22750 (N_22750,N_12071,N_13517);
xnor U22751 (N_22751,N_15187,N_15574);
xnor U22752 (N_22752,N_14500,N_14952);
or U22753 (N_22753,N_17082,N_16293);
nand U22754 (N_22754,N_13138,N_17065);
or U22755 (N_22755,N_17564,N_12454);
nand U22756 (N_22756,N_14834,N_13917);
nand U22757 (N_22757,N_15937,N_12045);
xnor U22758 (N_22758,N_13168,N_13573);
nor U22759 (N_22759,N_14864,N_14394);
nor U22760 (N_22760,N_13922,N_17009);
and U22761 (N_22761,N_13426,N_17446);
or U22762 (N_22762,N_14811,N_15006);
xnor U22763 (N_22763,N_17782,N_15362);
xor U22764 (N_22764,N_13697,N_15123);
nand U22765 (N_22765,N_16126,N_14663);
or U22766 (N_22766,N_13817,N_15104);
or U22767 (N_22767,N_16400,N_14202);
and U22768 (N_22768,N_12947,N_17543);
and U22769 (N_22769,N_17221,N_17069);
and U22770 (N_22770,N_14433,N_17076);
nand U22771 (N_22771,N_14986,N_17308);
nor U22772 (N_22772,N_12221,N_13197);
or U22773 (N_22773,N_16716,N_16822);
xnor U22774 (N_22774,N_16284,N_17359);
nand U22775 (N_22775,N_12599,N_12780);
xnor U22776 (N_22776,N_15974,N_15925);
xor U22777 (N_22777,N_12219,N_13114);
nor U22778 (N_22778,N_16018,N_16536);
nor U22779 (N_22779,N_13629,N_17413);
nor U22780 (N_22780,N_12149,N_12920);
xnor U22781 (N_22781,N_17328,N_12601);
xnor U22782 (N_22782,N_15676,N_16239);
xor U22783 (N_22783,N_13143,N_15447);
nor U22784 (N_22784,N_14712,N_13323);
and U22785 (N_22785,N_12478,N_12407);
nand U22786 (N_22786,N_15327,N_16472);
nand U22787 (N_22787,N_17479,N_16424);
nor U22788 (N_22788,N_13934,N_17211);
or U22789 (N_22789,N_12248,N_15947);
or U22790 (N_22790,N_17096,N_13432);
nand U22791 (N_22791,N_14204,N_13457);
nand U22792 (N_22792,N_14543,N_14952);
and U22793 (N_22793,N_13433,N_13089);
xor U22794 (N_22794,N_16151,N_17369);
xor U22795 (N_22795,N_16644,N_15290);
and U22796 (N_22796,N_12988,N_16562);
and U22797 (N_22797,N_13722,N_15526);
nand U22798 (N_22798,N_13486,N_14602);
nand U22799 (N_22799,N_13021,N_17043);
or U22800 (N_22800,N_13398,N_15992);
or U22801 (N_22801,N_17506,N_15179);
nand U22802 (N_22802,N_12876,N_16530);
and U22803 (N_22803,N_17716,N_17499);
and U22804 (N_22804,N_16041,N_13968);
and U22805 (N_22805,N_15039,N_13987);
nand U22806 (N_22806,N_15193,N_15125);
xnor U22807 (N_22807,N_17948,N_13334);
nand U22808 (N_22808,N_17624,N_15450);
and U22809 (N_22809,N_13412,N_16783);
xor U22810 (N_22810,N_16211,N_16333);
or U22811 (N_22811,N_13971,N_15590);
nand U22812 (N_22812,N_16890,N_15829);
nor U22813 (N_22813,N_13928,N_16881);
or U22814 (N_22814,N_15694,N_13456);
nand U22815 (N_22815,N_17400,N_14642);
or U22816 (N_22816,N_14770,N_14267);
nand U22817 (N_22817,N_15888,N_15334);
and U22818 (N_22818,N_15734,N_13535);
or U22819 (N_22819,N_17229,N_14211);
nor U22820 (N_22820,N_13910,N_14499);
nand U22821 (N_22821,N_17827,N_14573);
and U22822 (N_22822,N_13419,N_12289);
or U22823 (N_22823,N_13367,N_16164);
or U22824 (N_22824,N_17739,N_16651);
nand U22825 (N_22825,N_17416,N_16728);
and U22826 (N_22826,N_15490,N_15893);
nor U22827 (N_22827,N_14522,N_15817);
or U22828 (N_22828,N_17817,N_13182);
and U22829 (N_22829,N_12752,N_13364);
or U22830 (N_22830,N_17433,N_12679);
nand U22831 (N_22831,N_14520,N_17835);
nand U22832 (N_22832,N_15353,N_12700);
nor U22833 (N_22833,N_13233,N_14276);
and U22834 (N_22834,N_12326,N_17569);
nand U22835 (N_22835,N_12668,N_12841);
xnor U22836 (N_22836,N_12406,N_15328);
nand U22837 (N_22837,N_15557,N_17710);
and U22838 (N_22838,N_17967,N_16628);
nand U22839 (N_22839,N_16387,N_13781);
nand U22840 (N_22840,N_17224,N_16021);
nor U22841 (N_22841,N_16120,N_16227);
nand U22842 (N_22842,N_14812,N_12883);
xor U22843 (N_22843,N_17001,N_13623);
xnor U22844 (N_22844,N_12393,N_15179);
xor U22845 (N_22845,N_12095,N_17926);
xnor U22846 (N_22846,N_14023,N_14066);
nand U22847 (N_22847,N_13494,N_16662);
xnor U22848 (N_22848,N_16667,N_16081);
and U22849 (N_22849,N_16606,N_14380);
and U22850 (N_22850,N_13366,N_12471);
xnor U22851 (N_22851,N_13803,N_12039);
nand U22852 (N_22852,N_17998,N_14692);
xor U22853 (N_22853,N_13762,N_15809);
nand U22854 (N_22854,N_16772,N_13608);
nor U22855 (N_22855,N_12825,N_13021);
xnor U22856 (N_22856,N_15522,N_12589);
and U22857 (N_22857,N_14562,N_16524);
or U22858 (N_22858,N_14181,N_13201);
or U22859 (N_22859,N_16719,N_17390);
and U22860 (N_22860,N_13979,N_17676);
xor U22861 (N_22861,N_16116,N_12330);
and U22862 (N_22862,N_12077,N_17519);
nand U22863 (N_22863,N_12700,N_12271);
and U22864 (N_22864,N_14563,N_15115);
xor U22865 (N_22865,N_13120,N_12672);
or U22866 (N_22866,N_16181,N_15825);
nand U22867 (N_22867,N_13549,N_12189);
and U22868 (N_22868,N_16812,N_14981);
nand U22869 (N_22869,N_14430,N_12435);
and U22870 (N_22870,N_13707,N_13067);
and U22871 (N_22871,N_13939,N_14161);
nand U22872 (N_22872,N_12252,N_16079);
and U22873 (N_22873,N_17715,N_14343);
nor U22874 (N_22874,N_17842,N_16124);
xnor U22875 (N_22875,N_15166,N_13704);
and U22876 (N_22876,N_15279,N_12918);
nor U22877 (N_22877,N_12134,N_12947);
xnor U22878 (N_22878,N_12618,N_16565);
nor U22879 (N_22879,N_13275,N_14844);
and U22880 (N_22880,N_13704,N_15122);
nand U22881 (N_22881,N_17890,N_13740);
and U22882 (N_22882,N_12879,N_17447);
nor U22883 (N_22883,N_14808,N_17982);
nor U22884 (N_22884,N_15514,N_14813);
xnor U22885 (N_22885,N_13151,N_15560);
nor U22886 (N_22886,N_16232,N_12568);
xnor U22887 (N_22887,N_12808,N_13513);
xnor U22888 (N_22888,N_13865,N_12433);
and U22889 (N_22889,N_12706,N_15396);
nor U22890 (N_22890,N_14183,N_16073);
and U22891 (N_22891,N_16286,N_15199);
nand U22892 (N_22892,N_17975,N_13522);
xnor U22893 (N_22893,N_14610,N_13264);
xor U22894 (N_22894,N_14192,N_12802);
nor U22895 (N_22895,N_16161,N_14039);
nand U22896 (N_22896,N_12591,N_13564);
xnor U22897 (N_22897,N_13100,N_14028);
and U22898 (N_22898,N_16707,N_13989);
or U22899 (N_22899,N_13456,N_15277);
nor U22900 (N_22900,N_16909,N_16107);
and U22901 (N_22901,N_16115,N_16045);
nand U22902 (N_22902,N_17828,N_17364);
xnor U22903 (N_22903,N_16288,N_15256);
xor U22904 (N_22904,N_14610,N_15302);
or U22905 (N_22905,N_17215,N_16549);
nor U22906 (N_22906,N_13821,N_15405);
xor U22907 (N_22907,N_16295,N_14354);
nand U22908 (N_22908,N_16446,N_17619);
nand U22909 (N_22909,N_13923,N_12123);
or U22910 (N_22910,N_17672,N_17209);
or U22911 (N_22911,N_12430,N_13473);
or U22912 (N_22912,N_17946,N_16830);
nor U22913 (N_22913,N_13173,N_12512);
or U22914 (N_22914,N_17693,N_17728);
xnor U22915 (N_22915,N_16761,N_16317);
xnor U22916 (N_22916,N_16320,N_16377);
xnor U22917 (N_22917,N_14113,N_14259);
nor U22918 (N_22918,N_15911,N_12865);
nand U22919 (N_22919,N_12237,N_17228);
nand U22920 (N_22920,N_16885,N_13574);
and U22921 (N_22921,N_15036,N_16350);
nand U22922 (N_22922,N_16187,N_14293);
nand U22923 (N_22923,N_13763,N_15968);
nor U22924 (N_22924,N_14163,N_13202);
xor U22925 (N_22925,N_17364,N_15564);
and U22926 (N_22926,N_17339,N_13058);
and U22927 (N_22927,N_14691,N_12018);
nor U22928 (N_22928,N_13249,N_13136);
nand U22929 (N_22929,N_16677,N_16945);
nor U22930 (N_22930,N_15067,N_15621);
and U22931 (N_22931,N_12111,N_12070);
and U22932 (N_22932,N_14062,N_15227);
nor U22933 (N_22933,N_14273,N_13834);
nor U22934 (N_22934,N_14004,N_13948);
nand U22935 (N_22935,N_13541,N_16212);
and U22936 (N_22936,N_15291,N_12897);
and U22937 (N_22937,N_13108,N_15132);
and U22938 (N_22938,N_12482,N_17347);
nand U22939 (N_22939,N_15665,N_17926);
or U22940 (N_22940,N_14551,N_14704);
nor U22941 (N_22941,N_17057,N_17437);
nand U22942 (N_22942,N_13743,N_15320);
xnor U22943 (N_22943,N_17022,N_16908);
or U22944 (N_22944,N_12507,N_12945);
nor U22945 (N_22945,N_16774,N_16675);
and U22946 (N_22946,N_15524,N_17268);
and U22947 (N_22947,N_14046,N_17050);
and U22948 (N_22948,N_16832,N_16925);
and U22949 (N_22949,N_12406,N_13973);
and U22950 (N_22950,N_16194,N_17154);
or U22951 (N_22951,N_13432,N_16818);
and U22952 (N_22952,N_17285,N_15898);
nor U22953 (N_22953,N_14539,N_17598);
or U22954 (N_22954,N_15639,N_14691);
nand U22955 (N_22955,N_16937,N_12486);
xor U22956 (N_22956,N_12908,N_12277);
nor U22957 (N_22957,N_15045,N_16592);
xor U22958 (N_22958,N_13823,N_12200);
xor U22959 (N_22959,N_15356,N_14072);
and U22960 (N_22960,N_12167,N_12921);
xor U22961 (N_22961,N_12935,N_13327);
xnor U22962 (N_22962,N_13840,N_12548);
xnor U22963 (N_22963,N_13041,N_14314);
nand U22964 (N_22964,N_13327,N_14172);
xor U22965 (N_22965,N_14366,N_12389);
xor U22966 (N_22966,N_17290,N_16912);
nand U22967 (N_22967,N_16777,N_14561);
nand U22968 (N_22968,N_16556,N_14972);
xnor U22969 (N_22969,N_14507,N_14349);
xnor U22970 (N_22970,N_15868,N_14843);
nand U22971 (N_22971,N_13544,N_17129);
nor U22972 (N_22972,N_12538,N_13440);
xnor U22973 (N_22973,N_16976,N_14869);
xor U22974 (N_22974,N_15441,N_15293);
nor U22975 (N_22975,N_17795,N_17063);
nand U22976 (N_22976,N_15182,N_12016);
xor U22977 (N_22977,N_15582,N_12641);
nand U22978 (N_22978,N_13431,N_17231);
and U22979 (N_22979,N_14960,N_16191);
nor U22980 (N_22980,N_14381,N_14286);
nor U22981 (N_22981,N_12055,N_13243);
and U22982 (N_22982,N_17571,N_16919);
xor U22983 (N_22983,N_14043,N_13577);
or U22984 (N_22984,N_14392,N_13368);
and U22985 (N_22985,N_16063,N_12851);
and U22986 (N_22986,N_16379,N_13120);
xor U22987 (N_22987,N_12929,N_14483);
nor U22988 (N_22988,N_13287,N_13840);
nand U22989 (N_22989,N_13147,N_15557);
or U22990 (N_22990,N_15586,N_12862);
nor U22991 (N_22991,N_17334,N_16810);
xor U22992 (N_22992,N_14720,N_16116);
and U22993 (N_22993,N_14996,N_12651);
or U22994 (N_22994,N_14914,N_12442);
xnor U22995 (N_22995,N_13434,N_15653);
nand U22996 (N_22996,N_13637,N_15635);
nand U22997 (N_22997,N_13352,N_14727);
nor U22998 (N_22998,N_17345,N_14784);
and U22999 (N_22999,N_15525,N_14680);
nor U23000 (N_23000,N_15453,N_13033);
xor U23001 (N_23001,N_15401,N_14761);
xor U23002 (N_23002,N_12476,N_12109);
and U23003 (N_23003,N_16521,N_13123);
nor U23004 (N_23004,N_12374,N_12036);
and U23005 (N_23005,N_13507,N_14392);
or U23006 (N_23006,N_17531,N_12698);
or U23007 (N_23007,N_17529,N_16158);
or U23008 (N_23008,N_13996,N_13427);
and U23009 (N_23009,N_12053,N_16249);
xnor U23010 (N_23010,N_12234,N_15318);
or U23011 (N_23011,N_17132,N_14189);
or U23012 (N_23012,N_14549,N_12071);
nand U23013 (N_23013,N_15361,N_17949);
xnor U23014 (N_23014,N_15301,N_13574);
nand U23015 (N_23015,N_13267,N_14449);
or U23016 (N_23016,N_15884,N_15206);
nor U23017 (N_23017,N_15730,N_12439);
xnor U23018 (N_23018,N_14440,N_14579);
and U23019 (N_23019,N_14649,N_14746);
or U23020 (N_23020,N_16615,N_15913);
xnor U23021 (N_23021,N_12762,N_14668);
nor U23022 (N_23022,N_12871,N_13630);
nand U23023 (N_23023,N_15273,N_13501);
or U23024 (N_23024,N_16457,N_17464);
or U23025 (N_23025,N_13594,N_14806);
nand U23026 (N_23026,N_16235,N_17861);
and U23027 (N_23027,N_14698,N_16017);
nor U23028 (N_23028,N_13874,N_17321);
or U23029 (N_23029,N_12703,N_14255);
and U23030 (N_23030,N_13045,N_14905);
or U23031 (N_23031,N_13643,N_15776);
and U23032 (N_23032,N_14287,N_16598);
nand U23033 (N_23033,N_14511,N_15021);
nor U23034 (N_23034,N_17873,N_16874);
and U23035 (N_23035,N_16480,N_16801);
nand U23036 (N_23036,N_12503,N_14404);
nor U23037 (N_23037,N_14149,N_17533);
and U23038 (N_23038,N_13973,N_14193);
and U23039 (N_23039,N_15081,N_14862);
or U23040 (N_23040,N_13463,N_13195);
nand U23041 (N_23041,N_13848,N_16254);
and U23042 (N_23042,N_12917,N_16624);
or U23043 (N_23043,N_15641,N_13412);
and U23044 (N_23044,N_17316,N_17535);
xor U23045 (N_23045,N_14393,N_16359);
xor U23046 (N_23046,N_16556,N_15533);
xor U23047 (N_23047,N_16143,N_15494);
or U23048 (N_23048,N_15578,N_16878);
or U23049 (N_23049,N_17897,N_15408);
nand U23050 (N_23050,N_14154,N_12047);
or U23051 (N_23051,N_13793,N_12763);
nor U23052 (N_23052,N_15339,N_17939);
nor U23053 (N_23053,N_12854,N_17565);
or U23054 (N_23054,N_14238,N_13491);
nand U23055 (N_23055,N_17206,N_14149);
or U23056 (N_23056,N_13901,N_14178);
nand U23057 (N_23057,N_12946,N_12227);
nor U23058 (N_23058,N_17007,N_13494);
and U23059 (N_23059,N_12456,N_14895);
and U23060 (N_23060,N_15615,N_13802);
nor U23061 (N_23061,N_16234,N_12525);
nor U23062 (N_23062,N_13957,N_12464);
xnor U23063 (N_23063,N_13149,N_16561);
or U23064 (N_23064,N_17129,N_13780);
or U23065 (N_23065,N_17845,N_17203);
nor U23066 (N_23066,N_14185,N_16528);
xor U23067 (N_23067,N_12363,N_17893);
and U23068 (N_23068,N_15139,N_12447);
and U23069 (N_23069,N_14699,N_14718);
and U23070 (N_23070,N_15754,N_15683);
or U23071 (N_23071,N_13429,N_13330);
nand U23072 (N_23072,N_14473,N_17508);
or U23073 (N_23073,N_14692,N_13096);
xnor U23074 (N_23074,N_16177,N_14876);
and U23075 (N_23075,N_12875,N_17982);
or U23076 (N_23076,N_16962,N_15894);
nor U23077 (N_23077,N_13989,N_12398);
nand U23078 (N_23078,N_15379,N_17463);
xor U23079 (N_23079,N_17576,N_14807);
and U23080 (N_23080,N_17852,N_13662);
nor U23081 (N_23081,N_15877,N_12291);
or U23082 (N_23082,N_13114,N_16542);
nand U23083 (N_23083,N_13538,N_13101);
or U23084 (N_23084,N_14890,N_13835);
xnor U23085 (N_23085,N_14448,N_12489);
and U23086 (N_23086,N_14759,N_16764);
xor U23087 (N_23087,N_16912,N_16298);
nand U23088 (N_23088,N_17214,N_14946);
and U23089 (N_23089,N_15552,N_16002);
and U23090 (N_23090,N_17191,N_12820);
and U23091 (N_23091,N_13740,N_12925);
nor U23092 (N_23092,N_12174,N_12328);
xor U23093 (N_23093,N_17008,N_13319);
and U23094 (N_23094,N_17734,N_15303);
and U23095 (N_23095,N_16050,N_16467);
or U23096 (N_23096,N_15395,N_16427);
nor U23097 (N_23097,N_13254,N_17813);
nor U23098 (N_23098,N_15241,N_13835);
and U23099 (N_23099,N_15056,N_15564);
nand U23100 (N_23100,N_12365,N_13470);
or U23101 (N_23101,N_14072,N_16608);
or U23102 (N_23102,N_13538,N_12840);
and U23103 (N_23103,N_15964,N_15646);
and U23104 (N_23104,N_13432,N_12319);
nand U23105 (N_23105,N_17189,N_17778);
and U23106 (N_23106,N_17051,N_14444);
xnor U23107 (N_23107,N_13043,N_13064);
or U23108 (N_23108,N_15063,N_16463);
or U23109 (N_23109,N_12592,N_17821);
and U23110 (N_23110,N_17377,N_17540);
nand U23111 (N_23111,N_13452,N_17307);
nor U23112 (N_23112,N_13583,N_15171);
nor U23113 (N_23113,N_15510,N_12661);
xor U23114 (N_23114,N_13451,N_14785);
and U23115 (N_23115,N_12598,N_13931);
and U23116 (N_23116,N_13099,N_13254);
nand U23117 (N_23117,N_15884,N_13841);
nor U23118 (N_23118,N_13737,N_17170);
nand U23119 (N_23119,N_14370,N_13624);
or U23120 (N_23120,N_15938,N_12774);
nor U23121 (N_23121,N_14259,N_14339);
xnor U23122 (N_23122,N_17423,N_12132);
xnor U23123 (N_23123,N_17073,N_13915);
nor U23124 (N_23124,N_17529,N_12199);
xor U23125 (N_23125,N_17648,N_13932);
nand U23126 (N_23126,N_15073,N_12087);
and U23127 (N_23127,N_13909,N_15415);
xnor U23128 (N_23128,N_16283,N_16213);
xor U23129 (N_23129,N_15668,N_16268);
and U23130 (N_23130,N_13297,N_16353);
and U23131 (N_23131,N_13418,N_14481);
nand U23132 (N_23132,N_17411,N_17247);
nand U23133 (N_23133,N_17295,N_13448);
nand U23134 (N_23134,N_13769,N_16537);
or U23135 (N_23135,N_14164,N_17252);
nor U23136 (N_23136,N_15447,N_17870);
nor U23137 (N_23137,N_14144,N_16300);
or U23138 (N_23138,N_14951,N_15415);
nor U23139 (N_23139,N_17280,N_13960);
or U23140 (N_23140,N_12848,N_15216);
nand U23141 (N_23141,N_15974,N_16761);
nor U23142 (N_23142,N_16105,N_13526);
xnor U23143 (N_23143,N_13376,N_17836);
nand U23144 (N_23144,N_14137,N_15938);
nor U23145 (N_23145,N_14922,N_13545);
or U23146 (N_23146,N_12718,N_15432);
xor U23147 (N_23147,N_17602,N_17222);
or U23148 (N_23148,N_12478,N_13916);
xnor U23149 (N_23149,N_14560,N_15797);
nand U23150 (N_23150,N_15382,N_16834);
or U23151 (N_23151,N_17498,N_16616);
nand U23152 (N_23152,N_12255,N_13278);
or U23153 (N_23153,N_12477,N_17488);
nor U23154 (N_23154,N_13568,N_13264);
or U23155 (N_23155,N_15878,N_16742);
nand U23156 (N_23156,N_13230,N_13245);
xnor U23157 (N_23157,N_13314,N_16386);
xnor U23158 (N_23158,N_17915,N_13923);
and U23159 (N_23159,N_16820,N_15521);
or U23160 (N_23160,N_15742,N_13289);
nand U23161 (N_23161,N_17382,N_15980);
or U23162 (N_23162,N_14198,N_15537);
or U23163 (N_23163,N_16067,N_13266);
and U23164 (N_23164,N_13144,N_13549);
nand U23165 (N_23165,N_13095,N_15263);
nor U23166 (N_23166,N_13522,N_12021);
or U23167 (N_23167,N_13061,N_16557);
nand U23168 (N_23168,N_17080,N_12829);
nor U23169 (N_23169,N_12395,N_17650);
and U23170 (N_23170,N_14679,N_12648);
nor U23171 (N_23171,N_13244,N_12495);
and U23172 (N_23172,N_13373,N_13109);
and U23173 (N_23173,N_12130,N_16517);
nor U23174 (N_23174,N_12530,N_13823);
and U23175 (N_23175,N_13896,N_14694);
xnor U23176 (N_23176,N_17677,N_17057);
nand U23177 (N_23177,N_12932,N_16467);
xor U23178 (N_23178,N_13133,N_12736);
nor U23179 (N_23179,N_16956,N_17989);
and U23180 (N_23180,N_14631,N_16759);
and U23181 (N_23181,N_15382,N_13462);
or U23182 (N_23182,N_16904,N_13564);
nor U23183 (N_23183,N_15644,N_16263);
xor U23184 (N_23184,N_17521,N_17047);
or U23185 (N_23185,N_16095,N_12398);
or U23186 (N_23186,N_14941,N_12786);
or U23187 (N_23187,N_16977,N_17933);
nor U23188 (N_23188,N_17911,N_16170);
and U23189 (N_23189,N_15693,N_12864);
nand U23190 (N_23190,N_14096,N_16274);
and U23191 (N_23191,N_16837,N_12953);
nor U23192 (N_23192,N_14666,N_14911);
or U23193 (N_23193,N_15871,N_15588);
nor U23194 (N_23194,N_16926,N_16623);
or U23195 (N_23195,N_12189,N_12339);
xnor U23196 (N_23196,N_16586,N_17813);
and U23197 (N_23197,N_15509,N_16021);
nor U23198 (N_23198,N_14468,N_13171);
xnor U23199 (N_23199,N_12358,N_14555);
nor U23200 (N_23200,N_16835,N_14348);
nand U23201 (N_23201,N_14314,N_13600);
and U23202 (N_23202,N_14566,N_17145);
nor U23203 (N_23203,N_14378,N_12451);
or U23204 (N_23204,N_12399,N_14734);
nor U23205 (N_23205,N_13866,N_14360);
and U23206 (N_23206,N_13205,N_14631);
or U23207 (N_23207,N_17372,N_12449);
and U23208 (N_23208,N_16916,N_12005);
nand U23209 (N_23209,N_12405,N_16114);
nand U23210 (N_23210,N_14688,N_15572);
or U23211 (N_23211,N_14244,N_16794);
or U23212 (N_23212,N_16877,N_12004);
nand U23213 (N_23213,N_15827,N_15778);
and U23214 (N_23214,N_12604,N_16871);
xnor U23215 (N_23215,N_13520,N_17851);
nor U23216 (N_23216,N_17273,N_12680);
or U23217 (N_23217,N_12327,N_14708);
xor U23218 (N_23218,N_17364,N_14932);
nand U23219 (N_23219,N_15057,N_15483);
nor U23220 (N_23220,N_13197,N_14103);
or U23221 (N_23221,N_13924,N_13503);
or U23222 (N_23222,N_13785,N_15299);
and U23223 (N_23223,N_16321,N_15258);
xor U23224 (N_23224,N_16714,N_12086);
and U23225 (N_23225,N_14161,N_12678);
or U23226 (N_23226,N_12159,N_15945);
nand U23227 (N_23227,N_16968,N_12042);
or U23228 (N_23228,N_12041,N_14895);
nand U23229 (N_23229,N_16082,N_16178);
and U23230 (N_23230,N_14151,N_12566);
or U23231 (N_23231,N_17571,N_15666);
xor U23232 (N_23232,N_15731,N_14481);
or U23233 (N_23233,N_14912,N_17576);
xnor U23234 (N_23234,N_14715,N_12522);
and U23235 (N_23235,N_14853,N_15791);
nand U23236 (N_23236,N_17037,N_13282);
nand U23237 (N_23237,N_17638,N_17327);
and U23238 (N_23238,N_17502,N_14383);
xnor U23239 (N_23239,N_16932,N_17147);
and U23240 (N_23240,N_16141,N_17619);
or U23241 (N_23241,N_15160,N_12058);
nand U23242 (N_23242,N_14888,N_16965);
nor U23243 (N_23243,N_15719,N_13037);
nor U23244 (N_23244,N_12505,N_13759);
xnor U23245 (N_23245,N_15309,N_12776);
xor U23246 (N_23246,N_17315,N_13891);
xor U23247 (N_23247,N_14849,N_17017);
and U23248 (N_23248,N_12336,N_15456);
nand U23249 (N_23249,N_12686,N_16084);
xnor U23250 (N_23250,N_15435,N_17879);
xnor U23251 (N_23251,N_14031,N_14499);
nor U23252 (N_23252,N_14463,N_17784);
and U23253 (N_23253,N_14281,N_14029);
nor U23254 (N_23254,N_12949,N_12480);
nor U23255 (N_23255,N_12503,N_12553);
xnor U23256 (N_23256,N_16686,N_14059);
and U23257 (N_23257,N_15290,N_17651);
nand U23258 (N_23258,N_17240,N_14694);
or U23259 (N_23259,N_17641,N_13976);
and U23260 (N_23260,N_16244,N_15653);
xor U23261 (N_23261,N_16951,N_12508);
nor U23262 (N_23262,N_15734,N_16659);
and U23263 (N_23263,N_17597,N_15578);
nand U23264 (N_23264,N_13022,N_16939);
or U23265 (N_23265,N_15794,N_12562);
xnor U23266 (N_23266,N_15124,N_15994);
or U23267 (N_23267,N_16508,N_14269);
nor U23268 (N_23268,N_16770,N_15375);
xor U23269 (N_23269,N_14654,N_16779);
nor U23270 (N_23270,N_17407,N_12527);
xor U23271 (N_23271,N_17364,N_17611);
nor U23272 (N_23272,N_14808,N_17937);
and U23273 (N_23273,N_16979,N_17850);
nand U23274 (N_23274,N_16210,N_15645);
and U23275 (N_23275,N_14100,N_13593);
or U23276 (N_23276,N_16655,N_14881);
or U23277 (N_23277,N_17981,N_16460);
nand U23278 (N_23278,N_17436,N_17943);
nand U23279 (N_23279,N_15586,N_17968);
xnor U23280 (N_23280,N_12936,N_16275);
xnor U23281 (N_23281,N_16701,N_15257);
xor U23282 (N_23282,N_15639,N_15754);
xnor U23283 (N_23283,N_16819,N_16113);
and U23284 (N_23284,N_16493,N_15689);
nor U23285 (N_23285,N_17706,N_16166);
nor U23286 (N_23286,N_17899,N_15236);
nor U23287 (N_23287,N_16055,N_13582);
nor U23288 (N_23288,N_14702,N_16570);
xnor U23289 (N_23289,N_17936,N_13637);
nand U23290 (N_23290,N_16815,N_12624);
nor U23291 (N_23291,N_13103,N_16678);
and U23292 (N_23292,N_13523,N_12943);
nand U23293 (N_23293,N_12396,N_16252);
xor U23294 (N_23294,N_16643,N_13443);
nor U23295 (N_23295,N_14942,N_17783);
nand U23296 (N_23296,N_17682,N_16559);
nand U23297 (N_23297,N_12465,N_14853);
xor U23298 (N_23298,N_16042,N_12724);
nand U23299 (N_23299,N_15793,N_12723);
or U23300 (N_23300,N_15807,N_13413);
nor U23301 (N_23301,N_13525,N_16438);
xor U23302 (N_23302,N_17324,N_15317);
nand U23303 (N_23303,N_17196,N_14857);
and U23304 (N_23304,N_13167,N_15117);
and U23305 (N_23305,N_13887,N_13014);
nor U23306 (N_23306,N_13739,N_15139);
nand U23307 (N_23307,N_17012,N_12229);
nand U23308 (N_23308,N_13106,N_12462);
or U23309 (N_23309,N_16772,N_13181);
xor U23310 (N_23310,N_14120,N_14560);
nand U23311 (N_23311,N_16174,N_16826);
nand U23312 (N_23312,N_12615,N_14669);
nor U23313 (N_23313,N_14507,N_12305);
nor U23314 (N_23314,N_16819,N_13570);
and U23315 (N_23315,N_14241,N_14543);
nor U23316 (N_23316,N_16463,N_14982);
and U23317 (N_23317,N_14898,N_16064);
and U23318 (N_23318,N_15521,N_17684);
nor U23319 (N_23319,N_13393,N_13827);
or U23320 (N_23320,N_14988,N_14097);
nand U23321 (N_23321,N_15922,N_13083);
or U23322 (N_23322,N_12904,N_17862);
and U23323 (N_23323,N_14331,N_12646);
and U23324 (N_23324,N_14962,N_14328);
or U23325 (N_23325,N_12073,N_16378);
nand U23326 (N_23326,N_12231,N_14926);
or U23327 (N_23327,N_12381,N_17792);
nand U23328 (N_23328,N_16876,N_17678);
nand U23329 (N_23329,N_13119,N_15848);
nor U23330 (N_23330,N_15138,N_13888);
or U23331 (N_23331,N_14943,N_16653);
and U23332 (N_23332,N_15630,N_12132);
nor U23333 (N_23333,N_13280,N_15161);
xor U23334 (N_23334,N_12133,N_13691);
xnor U23335 (N_23335,N_17820,N_13293);
nand U23336 (N_23336,N_13116,N_17482);
or U23337 (N_23337,N_15874,N_17568);
xnor U23338 (N_23338,N_17338,N_16799);
nor U23339 (N_23339,N_14418,N_12236);
nand U23340 (N_23340,N_14547,N_13351);
xor U23341 (N_23341,N_12498,N_17218);
or U23342 (N_23342,N_16929,N_14475);
or U23343 (N_23343,N_12833,N_15703);
and U23344 (N_23344,N_14050,N_16319);
or U23345 (N_23345,N_14750,N_17863);
nand U23346 (N_23346,N_12318,N_16237);
nor U23347 (N_23347,N_16673,N_15267);
nand U23348 (N_23348,N_16244,N_12482);
nor U23349 (N_23349,N_12220,N_14254);
and U23350 (N_23350,N_15447,N_14848);
or U23351 (N_23351,N_16017,N_16600);
or U23352 (N_23352,N_13700,N_17758);
and U23353 (N_23353,N_17035,N_16393);
xnor U23354 (N_23354,N_12866,N_15527);
and U23355 (N_23355,N_16375,N_12491);
or U23356 (N_23356,N_16640,N_13417);
nor U23357 (N_23357,N_13853,N_13261);
or U23358 (N_23358,N_13347,N_16680);
xor U23359 (N_23359,N_16702,N_16549);
and U23360 (N_23360,N_14257,N_12675);
and U23361 (N_23361,N_12299,N_14515);
nand U23362 (N_23362,N_16903,N_15733);
and U23363 (N_23363,N_15478,N_12209);
xor U23364 (N_23364,N_14863,N_13047);
or U23365 (N_23365,N_17308,N_17605);
and U23366 (N_23366,N_14704,N_12005);
nand U23367 (N_23367,N_17139,N_13560);
or U23368 (N_23368,N_12126,N_15006);
nand U23369 (N_23369,N_15104,N_16886);
and U23370 (N_23370,N_13247,N_15665);
xor U23371 (N_23371,N_12346,N_12914);
xnor U23372 (N_23372,N_15968,N_15765);
or U23373 (N_23373,N_15458,N_13732);
and U23374 (N_23374,N_15452,N_13135);
nand U23375 (N_23375,N_17345,N_16503);
and U23376 (N_23376,N_17784,N_13348);
xnor U23377 (N_23377,N_14938,N_13707);
xor U23378 (N_23378,N_16732,N_17374);
and U23379 (N_23379,N_12480,N_17346);
nor U23380 (N_23380,N_17190,N_14934);
or U23381 (N_23381,N_16574,N_14991);
or U23382 (N_23382,N_13399,N_17913);
nor U23383 (N_23383,N_15238,N_16085);
or U23384 (N_23384,N_16097,N_17882);
or U23385 (N_23385,N_16219,N_17904);
or U23386 (N_23386,N_13713,N_14799);
and U23387 (N_23387,N_14914,N_15161);
nor U23388 (N_23388,N_16304,N_17215);
nor U23389 (N_23389,N_15828,N_15720);
or U23390 (N_23390,N_14316,N_16491);
nand U23391 (N_23391,N_17924,N_13946);
xor U23392 (N_23392,N_14012,N_13916);
nor U23393 (N_23393,N_15810,N_14878);
or U23394 (N_23394,N_13931,N_13213);
and U23395 (N_23395,N_17638,N_16129);
nor U23396 (N_23396,N_13605,N_17579);
nor U23397 (N_23397,N_15799,N_14395);
nor U23398 (N_23398,N_12526,N_13418);
nand U23399 (N_23399,N_17709,N_16125);
nor U23400 (N_23400,N_17113,N_17578);
nor U23401 (N_23401,N_12139,N_14244);
xnor U23402 (N_23402,N_13176,N_17377);
nand U23403 (N_23403,N_17378,N_15445);
xor U23404 (N_23404,N_16383,N_15375);
xnor U23405 (N_23405,N_15226,N_12367);
xnor U23406 (N_23406,N_13347,N_14862);
or U23407 (N_23407,N_12053,N_14486);
and U23408 (N_23408,N_17287,N_13190);
nor U23409 (N_23409,N_17536,N_13218);
or U23410 (N_23410,N_17872,N_15388);
nor U23411 (N_23411,N_14024,N_12832);
nand U23412 (N_23412,N_15971,N_17151);
xnor U23413 (N_23413,N_15285,N_14431);
nor U23414 (N_23414,N_15535,N_15856);
or U23415 (N_23415,N_13949,N_13982);
xor U23416 (N_23416,N_14089,N_16402);
xor U23417 (N_23417,N_14847,N_13657);
nor U23418 (N_23418,N_12367,N_16912);
nor U23419 (N_23419,N_15425,N_16299);
and U23420 (N_23420,N_14054,N_13100);
nor U23421 (N_23421,N_15480,N_13031);
nor U23422 (N_23422,N_15981,N_16736);
xnor U23423 (N_23423,N_15484,N_12071);
nand U23424 (N_23424,N_14743,N_15654);
and U23425 (N_23425,N_13166,N_13303);
xor U23426 (N_23426,N_13247,N_15117);
nor U23427 (N_23427,N_12839,N_12507);
nor U23428 (N_23428,N_14608,N_15077);
nor U23429 (N_23429,N_17069,N_14863);
nand U23430 (N_23430,N_13285,N_16500);
nand U23431 (N_23431,N_16898,N_17514);
xnor U23432 (N_23432,N_15364,N_15172);
and U23433 (N_23433,N_17325,N_14400);
nand U23434 (N_23434,N_15334,N_16215);
nand U23435 (N_23435,N_15968,N_12398);
or U23436 (N_23436,N_16247,N_14188);
nand U23437 (N_23437,N_13248,N_12979);
or U23438 (N_23438,N_12544,N_16203);
and U23439 (N_23439,N_16555,N_15608);
nor U23440 (N_23440,N_13058,N_17675);
nor U23441 (N_23441,N_14025,N_16186);
nand U23442 (N_23442,N_15459,N_16594);
and U23443 (N_23443,N_14467,N_17865);
nor U23444 (N_23444,N_12648,N_16935);
xor U23445 (N_23445,N_12394,N_15775);
and U23446 (N_23446,N_12838,N_12652);
nor U23447 (N_23447,N_15619,N_15712);
xnor U23448 (N_23448,N_17805,N_15484);
xnor U23449 (N_23449,N_13482,N_12095);
nor U23450 (N_23450,N_16220,N_12586);
or U23451 (N_23451,N_12310,N_15821);
nand U23452 (N_23452,N_15054,N_15478);
nor U23453 (N_23453,N_17048,N_15646);
xor U23454 (N_23454,N_13951,N_13174);
xor U23455 (N_23455,N_16641,N_16455);
xnor U23456 (N_23456,N_16673,N_12339);
nor U23457 (N_23457,N_16303,N_15485);
nand U23458 (N_23458,N_17328,N_13160);
and U23459 (N_23459,N_12907,N_12487);
and U23460 (N_23460,N_16272,N_12985);
nand U23461 (N_23461,N_13254,N_13811);
nand U23462 (N_23462,N_17138,N_17329);
xnor U23463 (N_23463,N_15499,N_12072);
nand U23464 (N_23464,N_17586,N_17929);
and U23465 (N_23465,N_12101,N_14962);
nor U23466 (N_23466,N_17108,N_16548);
or U23467 (N_23467,N_13966,N_12277);
nand U23468 (N_23468,N_16689,N_12703);
nor U23469 (N_23469,N_16765,N_17418);
and U23470 (N_23470,N_13079,N_17042);
and U23471 (N_23471,N_17803,N_16300);
and U23472 (N_23472,N_12777,N_12999);
and U23473 (N_23473,N_15590,N_12442);
nor U23474 (N_23474,N_16799,N_17379);
or U23475 (N_23475,N_13127,N_17166);
xnor U23476 (N_23476,N_17236,N_17773);
nor U23477 (N_23477,N_14469,N_14768);
and U23478 (N_23478,N_14995,N_15311);
and U23479 (N_23479,N_15330,N_14953);
or U23480 (N_23480,N_14893,N_17055);
or U23481 (N_23481,N_12465,N_15852);
xor U23482 (N_23482,N_16827,N_14853);
nand U23483 (N_23483,N_14224,N_13361);
or U23484 (N_23484,N_15817,N_17251);
xnor U23485 (N_23485,N_14320,N_16903);
or U23486 (N_23486,N_14713,N_16731);
nand U23487 (N_23487,N_14987,N_12579);
xnor U23488 (N_23488,N_14157,N_16783);
nand U23489 (N_23489,N_12169,N_17990);
and U23490 (N_23490,N_14552,N_12342);
or U23491 (N_23491,N_16519,N_17565);
nor U23492 (N_23492,N_17598,N_14122);
nor U23493 (N_23493,N_13292,N_15806);
or U23494 (N_23494,N_13394,N_12902);
or U23495 (N_23495,N_17875,N_17136);
and U23496 (N_23496,N_17671,N_12503);
xnor U23497 (N_23497,N_14102,N_16730);
nand U23498 (N_23498,N_16933,N_17612);
and U23499 (N_23499,N_16324,N_17675);
or U23500 (N_23500,N_16305,N_15021);
or U23501 (N_23501,N_12302,N_17948);
nand U23502 (N_23502,N_14677,N_13584);
or U23503 (N_23503,N_13323,N_15746);
nor U23504 (N_23504,N_13936,N_16172);
and U23505 (N_23505,N_16718,N_14001);
and U23506 (N_23506,N_17905,N_13072);
and U23507 (N_23507,N_15423,N_13021);
or U23508 (N_23508,N_17485,N_14959);
or U23509 (N_23509,N_15444,N_13345);
xnor U23510 (N_23510,N_13750,N_14307);
nor U23511 (N_23511,N_12271,N_14191);
nand U23512 (N_23512,N_14043,N_17333);
xnor U23513 (N_23513,N_12297,N_15218);
xor U23514 (N_23514,N_16133,N_13993);
and U23515 (N_23515,N_13306,N_15296);
nor U23516 (N_23516,N_13444,N_16929);
nor U23517 (N_23517,N_16891,N_13998);
and U23518 (N_23518,N_17263,N_14775);
and U23519 (N_23519,N_15887,N_17026);
or U23520 (N_23520,N_13517,N_13931);
or U23521 (N_23521,N_15382,N_12419);
or U23522 (N_23522,N_17248,N_16609);
xor U23523 (N_23523,N_15385,N_16181);
or U23524 (N_23524,N_15190,N_14580);
or U23525 (N_23525,N_14701,N_13213);
nand U23526 (N_23526,N_14405,N_12060);
xor U23527 (N_23527,N_16272,N_17195);
xor U23528 (N_23528,N_12675,N_12204);
and U23529 (N_23529,N_16856,N_17453);
nor U23530 (N_23530,N_16725,N_13428);
nand U23531 (N_23531,N_17610,N_17795);
nand U23532 (N_23532,N_12805,N_12289);
xor U23533 (N_23533,N_15531,N_17902);
xnor U23534 (N_23534,N_13375,N_16849);
nor U23535 (N_23535,N_12837,N_16623);
xnor U23536 (N_23536,N_14790,N_15014);
nand U23537 (N_23537,N_13631,N_16158);
xor U23538 (N_23538,N_13413,N_16378);
nand U23539 (N_23539,N_16334,N_14068);
nand U23540 (N_23540,N_14384,N_14634);
or U23541 (N_23541,N_13826,N_16888);
nor U23542 (N_23542,N_13473,N_16653);
and U23543 (N_23543,N_14499,N_16006);
or U23544 (N_23544,N_16873,N_16948);
xnor U23545 (N_23545,N_15138,N_16257);
and U23546 (N_23546,N_14089,N_13280);
and U23547 (N_23547,N_16953,N_13867);
xor U23548 (N_23548,N_14722,N_17673);
xnor U23549 (N_23549,N_13229,N_16349);
nor U23550 (N_23550,N_12695,N_12262);
nand U23551 (N_23551,N_16782,N_14832);
and U23552 (N_23552,N_12277,N_15485);
and U23553 (N_23553,N_15584,N_17416);
nor U23554 (N_23554,N_16727,N_17216);
xnor U23555 (N_23555,N_14442,N_14012);
nor U23556 (N_23556,N_15771,N_15671);
xnor U23557 (N_23557,N_17386,N_15194);
nand U23558 (N_23558,N_13977,N_15007);
nand U23559 (N_23559,N_15152,N_17940);
xor U23560 (N_23560,N_17652,N_16770);
and U23561 (N_23561,N_14840,N_14548);
or U23562 (N_23562,N_15064,N_12493);
and U23563 (N_23563,N_13556,N_16499);
xor U23564 (N_23564,N_17329,N_12246);
xor U23565 (N_23565,N_12023,N_14237);
or U23566 (N_23566,N_17606,N_17728);
xor U23567 (N_23567,N_13847,N_12352);
and U23568 (N_23568,N_15300,N_15693);
or U23569 (N_23569,N_17860,N_15728);
and U23570 (N_23570,N_15494,N_14875);
nor U23571 (N_23571,N_12991,N_13470);
xnor U23572 (N_23572,N_12153,N_12796);
and U23573 (N_23573,N_13335,N_15911);
xnor U23574 (N_23574,N_14800,N_14933);
nor U23575 (N_23575,N_16017,N_15649);
nor U23576 (N_23576,N_13689,N_12257);
xnor U23577 (N_23577,N_12588,N_16556);
nand U23578 (N_23578,N_15533,N_13221);
xnor U23579 (N_23579,N_15283,N_12289);
or U23580 (N_23580,N_16121,N_16465);
nand U23581 (N_23581,N_13097,N_12918);
and U23582 (N_23582,N_15812,N_16138);
and U23583 (N_23583,N_14771,N_13282);
nor U23584 (N_23584,N_15086,N_14980);
nor U23585 (N_23585,N_17514,N_16244);
nor U23586 (N_23586,N_12819,N_14222);
xnor U23587 (N_23587,N_13622,N_12612);
nand U23588 (N_23588,N_14812,N_15111);
nor U23589 (N_23589,N_12976,N_15332);
nand U23590 (N_23590,N_14975,N_16105);
nor U23591 (N_23591,N_14801,N_13089);
nand U23592 (N_23592,N_14905,N_16422);
nor U23593 (N_23593,N_12053,N_14670);
nand U23594 (N_23594,N_16960,N_15251);
xnor U23595 (N_23595,N_12428,N_16888);
nand U23596 (N_23596,N_15756,N_15117);
nor U23597 (N_23597,N_16212,N_12680);
or U23598 (N_23598,N_17085,N_13596);
or U23599 (N_23599,N_15577,N_14459);
nor U23600 (N_23600,N_13984,N_15517);
nor U23601 (N_23601,N_17400,N_12020);
xor U23602 (N_23602,N_14789,N_13470);
or U23603 (N_23603,N_12172,N_12092);
nand U23604 (N_23604,N_16761,N_12205);
or U23605 (N_23605,N_12423,N_13193);
nand U23606 (N_23606,N_13663,N_15158);
or U23607 (N_23607,N_12465,N_13900);
nor U23608 (N_23608,N_16327,N_15113);
xnor U23609 (N_23609,N_13192,N_17536);
xor U23610 (N_23610,N_13729,N_14834);
xor U23611 (N_23611,N_16001,N_14948);
nor U23612 (N_23612,N_12744,N_15104);
or U23613 (N_23613,N_13816,N_12864);
xnor U23614 (N_23614,N_12609,N_14261);
and U23615 (N_23615,N_17729,N_12385);
xor U23616 (N_23616,N_14370,N_17612);
nand U23617 (N_23617,N_12892,N_16724);
nand U23618 (N_23618,N_17777,N_13922);
and U23619 (N_23619,N_12306,N_17402);
nand U23620 (N_23620,N_15346,N_12053);
and U23621 (N_23621,N_17470,N_16375);
or U23622 (N_23622,N_14465,N_16567);
or U23623 (N_23623,N_16566,N_16205);
nand U23624 (N_23624,N_13478,N_14599);
nor U23625 (N_23625,N_16330,N_15899);
or U23626 (N_23626,N_15094,N_16775);
and U23627 (N_23627,N_17962,N_15085);
and U23628 (N_23628,N_12818,N_13949);
xnor U23629 (N_23629,N_16856,N_12690);
or U23630 (N_23630,N_12345,N_17940);
nand U23631 (N_23631,N_14297,N_16417);
or U23632 (N_23632,N_15939,N_16940);
xnor U23633 (N_23633,N_15419,N_13490);
nor U23634 (N_23634,N_13351,N_15960);
and U23635 (N_23635,N_16689,N_16422);
or U23636 (N_23636,N_12597,N_12338);
and U23637 (N_23637,N_15526,N_17806);
xnor U23638 (N_23638,N_15600,N_16380);
nand U23639 (N_23639,N_15889,N_13876);
nor U23640 (N_23640,N_12720,N_16388);
nor U23641 (N_23641,N_13631,N_15634);
and U23642 (N_23642,N_13115,N_14605);
or U23643 (N_23643,N_13550,N_14913);
and U23644 (N_23644,N_17536,N_16757);
or U23645 (N_23645,N_14167,N_13153);
or U23646 (N_23646,N_12044,N_12479);
or U23647 (N_23647,N_12116,N_16620);
xnor U23648 (N_23648,N_13124,N_17408);
nand U23649 (N_23649,N_15287,N_16343);
xnor U23650 (N_23650,N_17907,N_13133);
or U23651 (N_23651,N_15056,N_13003);
and U23652 (N_23652,N_17508,N_13294);
or U23653 (N_23653,N_17252,N_17496);
and U23654 (N_23654,N_12232,N_13901);
and U23655 (N_23655,N_17668,N_14207);
or U23656 (N_23656,N_17267,N_15626);
nor U23657 (N_23657,N_14542,N_16359);
or U23658 (N_23658,N_12025,N_14469);
or U23659 (N_23659,N_14067,N_17684);
xor U23660 (N_23660,N_15732,N_12247);
nor U23661 (N_23661,N_12135,N_17746);
nor U23662 (N_23662,N_15954,N_16378);
nand U23663 (N_23663,N_12256,N_16843);
nor U23664 (N_23664,N_12777,N_13504);
nor U23665 (N_23665,N_16858,N_13706);
or U23666 (N_23666,N_12285,N_12810);
xor U23667 (N_23667,N_13369,N_13896);
xor U23668 (N_23668,N_14780,N_16178);
and U23669 (N_23669,N_16310,N_15561);
nand U23670 (N_23670,N_17891,N_15463);
or U23671 (N_23671,N_13482,N_16173);
xor U23672 (N_23672,N_13603,N_17774);
nand U23673 (N_23673,N_14715,N_12909);
nor U23674 (N_23674,N_15726,N_16620);
nor U23675 (N_23675,N_15301,N_14652);
and U23676 (N_23676,N_16467,N_12054);
or U23677 (N_23677,N_16297,N_16718);
and U23678 (N_23678,N_17619,N_16537);
nor U23679 (N_23679,N_13757,N_13375);
or U23680 (N_23680,N_17781,N_16908);
and U23681 (N_23681,N_16330,N_15262);
nor U23682 (N_23682,N_16272,N_12783);
and U23683 (N_23683,N_16138,N_16443);
nand U23684 (N_23684,N_17631,N_13300);
nand U23685 (N_23685,N_16110,N_13844);
and U23686 (N_23686,N_15426,N_12369);
nand U23687 (N_23687,N_12496,N_15821);
and U23688 (N_23688,N_14042,N_14341);
or U23689 (N_23689,N_14643,N_16172);
and U23690 (N_23690,N_17014,N_13379);
or U23691 (N_23691,N_13388,N_14716);
xnor U23692 (N_23692,N_17864,N_15011);
nand U23693 (N_23693,N_14561,N_12188);
nor U23694 (N_23694,N_12289,N_17990);
nor U23695 (N_23695,N_14394,N_17360);
and U23696 (N_23696,N_16658,N_12299);
and U23697 (N_23697,N_12375,N_17014);
nor U23698 (N_23698,N_12968,N_17486);
and U23699 (N_23699,N_17139,N_14359);
nand U23700 (N_23700,N_14690,N_13181);
nor U23701 (N_23701,N_12589,N_12560);
nor U23702 (N_23702,N_14998,N_14798);
nor U23703 (N_23703,N_12088,N_12416);
or U23704 (N_23704,N_13328,N_12802);
nor U23705 (N_23705,N_14285,N_13169);
and U23706 (N_23706,N_13354,N_16536);
nand U23707 (N_23707,N_13734,N_16614);
nand U23708 (N_23708,N_17959,N_12166);
xor U23709 (N_23709,N_15185,N_12472);
nand U23710 (N_23710,N_17233,N_12948);
nand U23711 (N_23711,N_13208,N_12285);
nor U23712 (N_23712,N_12791,N_17850);
nor U23713 (N_23713,N_13328,N_13538);
and U23714 (N_23714,N_17542,N_13362);
nor U23715 (N_23715,N_14833,N_15488);
or U23716 (N_23716,N_12393,N_14350);
and U23717 (N_23717,N_16888,N_12966);
and U23718 (N_23718,N_12175,N_15715);
and U23719 (N_23719,N_16841,N_16234);
nand U23720 (N_23720,N_16204,N_13032);
or U23721 (N_23721,N_16742,N_17525);
nor U23722 (N_23722,N_12270,N_17143);
nor U23723 (N_23723,N_14110,N_15179);
xor U23724 (N_23724,N_12397,N_15960);
xor U23725 (N_23725,N_17277,N_15607);
nor U23726 (N_23726,N_13148,N_16625);
nand U23727 (N_23727,N_13803,N_12173);
or U23728 (N_23728,N_12333,N_16292);
xnor U23729 (N_23729,N_15854,N_13967);
nand U23730 (N_23730,N_17434,N_17800);
xnor U23731 (N_23731,N_14561,N_14065);
xor U23732 (N_23732,N_16459,N_13505);
nand U23733 (N_23733,N_13817,N_16946);
xor U23734 (N_23734,N_15888,N_12025);
and U23735 (N_23735,N_16891,N_12121);
nor U23736 (N_23736,N_12185,N_16059);
and U23737 (N_23737,N_16670,N_14825);
xor U23738 (N_23738,N_13539,N_16868);
nor U23739 (N_23739,N_12207,N_13230);
nand U23740 (N_23740,N_15230,N_15241);
or U23741 (N_23741,N_12958,N_14172);
nand U23742 (N_23742,N_13068,N_14457);
nand U23743 (N_23743,N_16691,N_13181);
nor U23744 (N_23744,N_13873,N_14421);
xnor U23745 (N_23745,N_15403,N_15318);
or U23746 (N_23746,N_15264,N_12063);
and U23747 (N_23747,N_15248,N_16228);
or U23748 (N_23748,N_16857,N_12490);
or U23749 (N_23749,N_13050,N_12310);
xor U23750 (N_23750,N_15708,N_16256);
nor U23751 (N_23751,N_16886,N_15608);
and U23752 (N_23752,N_17538,N_15328);
or U23753 (N_23753,N_14574,N_13088);
or U23754 (N_23754,N_16009,N_16419);
nand U23755 (N_23755,N_16282,N_15445);
xnor U23756 (N_23756,N_13327,N_16547);
and U23757 (N_23757,N_13748,N_17623);
nor U23758 (N_23758,N_16571,N_16917);
or U23759 (N_23759,N_13480,N_13849);
or U23760 (N_23760,N_15134,N_14488);
xor U23761 (N_23761,N_13230,N_15970);
nand U23762 (N_23762,N_16521,N_15895);
or U23763 (N_23763,N_16592,N_16389);
and U23764 (N_23764,N_14058,N_13512);
nor U23765 (N_23765,N_17331,N_17505);
xnor U23766 (N_23766,N_16163,N_17455);
xnor U23767 (N_23767,N_17231,N_13353);
or U23768 (N_23768,N_16512,N_14864);
nand U23769 (N_23769,N_15434,N_14335);
nand U23770 (N_23770,N_12388,N_15738);
xnor U23771 (N_23771,N_16717,N_12749);
nand U23772 (N_23772,N_15668,N_17547);
xnor U23773 (N_23773,N_13373,N_15638);
xnor U23774 (N_23774,N_13948,N_16411);
and U23775 (N_23775,N_14789,N_13471);
or U23776 (N_23776,N_16315,N_16774);
and U23777 (N_23777,N_14909,N_17623);
and U23778 (N_23778,N_15991,N_16804);
nand U23779 (N_23779,N_17450,N_12552);
or U23780 (N_23780,N_15110,N_12995);
xnor U23781 (N_23781,N_13270,N_15288);
nor U23782 (N_23782,N_13887,N_15502);
nand U23783 (N_23783,N_16318,N_13314);
or U23784 (N_23784,N_15325,N_13204);
or U23785 (N_23785,N_15690,N_15419);
xor U23786 (N_23786,N_12133,N_15765);
nor U23787 (N_23787,N_16682,N_17154);
xor U23788 (N_23788,N_14994,N_14304);
and U23789 (N_23789,N_15043,N_17970);
xor U23790 (N_23790,N_13363,N_17449);
and U23791 (N_23791,N_12968,N_13650);
or U23792 (N_23792,N_13775,N_15222);
nand U23793 (N_23793,N_14425,N_17367);
nand U23794 (N_23794,N_17661,N_13570);
or U23795 (N_23795,N_16598,N_17696);
nand U23796 (N_23796,N_12499,N_13873);
nand U23797 (N_23797,N_16036,N_15550);
nor U23798 (N_23798,N_17802,N_17868);
and U23799 (N_23799,N_16292,N_13658);
or U23800 (N_23800,N_14601,N_16801);
and U23801 (N_23801,N_13471,N_17059);
xor U23802 (N_23802,N_16399,N_16062);
nor U23803 (N_23803,N_13017,N_16278);
nand U23804 (N_23804,N_15828,N_13475);
nand U23805 (N_23805,N_12590,N_17772);
nand U23806 (N_23806,N_17912,N_17649);
and U23807 (N_23807,N_14171,N_15799);
xnor U23808 (N_23808,N_14571,N_13545);
or U23809 (N_23809,N_15429,N_14745);
nor U23810 (N_23810,N_13664,N_16534);
xnor U23811 (N_23811,N_13506,N_13454);
xnor U23812 (N_23812,N_15894,N_13418);
nand U23813 (N_23813,N_16309,N_17398);
xor U23814 (N_23814,N_15573,N_15977);
and U23815 (N_23815,N_14432,N_17044);
nor U23816 (N_23816,N_17485,N_12236);
nor U23817 (N_23817,N_13432,N_13304);
nor U23818 (N_23818,N_12690,N_16573);
and U23819 (N_23819,N_12127,N_14754);
nand U23820 (N_23820,N_17765,N_17052);
xor U23821 (N_23821,N_13883,N_16993);
and U23822 (N_23822,N_17188,N_13620);
or U23823 (N_23823,N_14828,N_15491);
nor U23824 (N_23824,N_17348,N_16603);
nand U23825 (N_23825,N_17357,N_16570);
nor U23826 (N_23826,N_16616,N_12888);
or U23827 (N_23827,N_17268,N_13122);
and U23828 (N_23828,N_12143,N_17097);
xor U23829 (N_23829,N_15361,N_15392);
xnor U23830 (N_23830,N_16702,N_13665);
xor U23831 (N_23831,N_17631,N_15614);
nor U23832 (N_23832,N_15275,N_12916);
nand U23833 (N_23833,N_16830,N_15393);
nand U23834 (N_23834,N_15265,N_15362);
nor U23835 (N_23835,N_17397,N_16020);
or U23836 (N_23836,N_15223,N_14246);
xor U23837 (N_23837,N_12394,N_15417);
and U23838 (N_23838,N_12408,N_13219);
or U23839 (N_23839,N_17290,N_15109);
and U23840 (N_23840,N_14688,N_17330);
xor U23841 (N_23841,N_13684,N_12885);
or U23842 (N_23842,N_12698,N_17356);
or U23843 (N_23843,N_12522,N_13717);
xor U23844 (N_23844,N_16971,N_15893);
nand U23845 (N_23845,N_12642,N_15492);
xnor U23846 (N_23846,N_17899,N_12878);
xor U23847 (N_23847,N_13647,N_12444);
nand U23848 (N_23848,N_13060,N_12148);
nor U23849 (N_23849,N_16452,N_16457);
nor U23850 (N_23850,N_16339,N_16489);
xor U23851 (N_23851,N_15057,N_16151);
or U23852 (N_23852,N_13273,N_17099);
nand U23853 (N_23853,N_16918,N_15720);
or U23854 (N_23854,N_17738,N_13553);
xor U23855 (N_23855,N_15215,N_12676);
nor U23856 (N_23856,N_17135,N_12228);
or U23857 (N_23857,N_16102,N_13762);
and U23858 (N_23858,N_12567,N_13729);
xnor U23859 (N_23859,N_16163,N_15286);
and U23860 (N_23860,N_14997,N_12133);
nor U23861 (N_23861,N_14671,N_16402);
nand U23862 (N_23862,N_15019,N_13175);
or U23863 (N_23863,N_12082,N_13623);
and U23864 (N_23864,N_12432,N_12668);
and U23865 (N_23865,N_15465,N_13748);
and U23866 (N_23866,N_16129,N_13123);
and U23867 (N_23867,N_13851,N_13050);
or U23868 (N_23868,N_16160,N_12213);
xor U23869 (N_23869,N_12554,N_13762);
and U23870 (N_23870,N_14428,N_16143);
and U23871 (N_23871,N_15567,N_17084);
nand U23872 (N_23872,N_16423,N_12244);
and U23873 (N_23873,N_15168,N_17408);
xnor U23874 (N_23874,N_14745,N_16280);
nand U23875 (N_23875,N_14162,N_13640);
xnor U23876 (N_23876,N_12792,N_16417);
or U23877 (N_23877,N_12223,N_16916);
nand U23878 (N_23878,N_17299,N_12814);
and U23879 (N_23879,N_14897,N_12579);
xnor U23880 (N_23880,N_12432,N_12660);
nand U23881 (N_23881,N_16634,N_14330);
nor U23882 (N_23882,N_17101,N_12172);
nand U23883 (N_23883,N_13483,N_16209);
nor U23884 (N_23884,N_17042,N_14463);
nand U23885 (N_23885,N_17398,N_14001);
nand U23886 (N_23886,N_16571,N_17785);
nand U23887 (N_23887,N_14964,N_16472);
xor U23888 (N_23888,N_14908,N_13041);
and U23889 (N_23889,N_15953,N_14331);
and U23890 (N_23890,N_16114,N_15304);
nand U23891 (N_23891,N_16164,N_13134);
or U23892 (N_23892,N_14211,N_13800);
and U23893 (N_23893,N_12076,N_16254);
or U23894 (N_23894,N_17419,N_15995);
xnor U23895 (N_23895,N_16682,N_14852);
xor U23896 (N_23896,N_15297,N_12962);
xor U23897 (N_23897,N_14387,N_13794);
nand U23898 (N_23898,N_12574,N_16257);
and U23899 (N_23899,N_17129,N_16628);
nor U23900 (N_23900,N_14764,N_17582);
and U23901 (N_23901,N_17863,N_17867);
nor U23902 (N_23902,N_12510,N_16836);
nand U23903 (N_23903,N_15343,N_14792);
and U23904 (N_23904,N_13286,N_17612);
nand U23905 (N_23905,N_13171,N_16139);
or U23906 (N_23906,N_13896,N_15296);
nand U23907 (N_23907,N_17079,N_12274);
nand U23908 (N_23908,N_17471,N_14542);
or U23909 (N_23909,N_14974,N_17903);
or U23910 (N_23910,N_13417,N_13184);
or U23911 (N_23911,N_14542,N_12810);
nand U23912 (N_23912,N_15770,N_16958);
nand U23913 (N_23913,N_16370,N_14329);
xnor U23914 (N_23914,N_12922,N_14220);
nand U23915 (N_23915,N_14380,N_13350);
nand U23916 (N_23916,N_17223,N_14573);
or U23917 (N_23917,N_12621,N_13631);
nor U23918 (N_23918,N_17345,N_15729);
nor U23919 (N_23919,N_14656,N_13907);
nand U23920 (N_23920,N_15590,N_15617);
nand U23921 (N_23921,N_13196,N_13762);
xor U23922 (N_23922,N_15412,N_14256);
and U23923 (N_23923,N_12178,N_15971);
or U23924 (N_23924,N_15852,N_16896);
or U23925 (N_23925,N_15935,N_13875);
or U23926 (N_23926,N_12626,N_14167);
nand U23927 (N_23927,N_17290,N_17310);
or U23928 (N_23928,N_15745,N_17727);
xnor U23929 (N_23929,N_12270,N_13853);
nor U23930 (N_23930,N_15073,N_17831);
and U23931 (N_23931,N_14566,N_12966);
or U23932 (N_23932,N_16294,N_13863);
nand U23933 (N_23933,N_13205,N_13604);
nor U23934 (N_23934,N_15302,N_16239);
xor U23935 (N_23935,N_15454,N_14697);
nand U23936 (N_23936,N_14670,N_15825);
and U23937 (N_23937,N_17480,N_13288);
nand U23938 (N_23938,N_13263,N_15032);
and U23939 (N_23939,N_16391,N_17297);
and U23940 (N_23940,N_16196,N_14400);
and U23941 (N_23941,N_15473,N_14026);
nor U23942 (N_23942,N_13444,N_15381);
nand U23943 (N_23943,N_16547,N_14400);
xor U23944 (N_23944,N_16798,N_14823);
nand U23945 (N_23945,N_17101,N_13464);
nand U23946 (N_23946,N_17350,N_12975);
nor U23947 (N_23947,N_17511,N_14624);
or U23948 (N_23948,N_14111,N_17973);
nor U23949 (N_23949,N_17766,N_16451);
nor U23950 (N_23950,N_12940,N_13001);
or U23951 (N_23951,N_16452,N_15457);
xnor U23952 (N_23952,N_17561,N_15529);
nand U23953 (N_23953,N_16500,N_14577);
or U23954 (N_23954,N_15660,N_17679);
nand U23955 (N_23955,N_17252,N_12997);
xnor U23956 (N_23956,N_16842,N_15498);
nand U23957 (N_23957,N_14076,N_15944);
or U23958 (N_23958,N_12332,N_12503);
or U23959 (N_23959,N_16659,N_15898);
nor U23960 (N_23960,N_14093,N_16905);
or U23961 (N_23961,N_15416,N_15691);
xnor U23962 (N_23962,N_14672,N_14681);
and U23963 (N_23963,N_15513,N_16420);
nor U23964 (N_23964,N_12675,N_15327);
nor U23965 (N_23965,N_12857,N_15937);
and U23966 (N_23966,N_13236,N_13019);
and U23967 (N_23967,N_16867,N_13478);
or U23968 (N_23968,N_16031,N_12335);
xor U23969 (N_23969,N_15795,N_15751);
nor U23970 (N_23970,N_12460,N_15285);
nand U23971 (N_23971,N_17493,N_12573);
nand U23972 (N_23972,N_17345,N_13824);
nand U23973 (N_23973,N_17523,N_12792);
xor U23974 (N_23974,N_15290,N_17975);
and U23975 (N_23975,N_15196,N_17743);
xnor U23976 (N_23976,N_17105,N_17231);
nor U23977 (N_23977,N_13937,N_17906);
or U23978 (N_23978,N_13172,N_13443);
nor U23979 (N_23979,N_13048,N_13608);
nor U23980 (N_23980,N_15353,N_17333);
nor U23981 (N_23981,N_12740,N_12808);
and U23982 (N_23982,N_14445,N_15017);
nor U23983 (N_23983,N_12912,N_15374);
nand U23984 (N_23984,N_13877,N_12087);
nor U23985 (N_23985,N_17588,N_16550);
and U23986 (N_23986,N_12590,N_12903);
or U23987 (N_23987,N_16489,N_12237);
nor U23988 (N_23988,N_16682,N_15453);
nor U23989 (N_23989,N_15657,N_13653);
and U23990 (N_23990,N_16827,N_12187);
nand U23991 (N_23991,N_12194,N_14037);
xnor U23992 (N_23992,N_14889,N_17950);
nor U23993 (N_23993,N_16649,N_14829);
nor U23994 (N_23994,N_13152,N_15791);
xnor U23995 (N_23995,N_14505,N_15135);
nor U23996 (N_23996,N_15451,N_15158);
nor U23997 (N_23997,N_12335,N_15315);
and U23998 (N_23998,N_17423,N_15976);
or U23999 (N_23999,N_16785,N_16195);
nor U24000 (N_24000,N_18028,N_19346);
xnor U24001 (N_24001,N_18177,N_20519);
nor U24002 (N_24002,N_21980,N_21480);
and U24003 (N_24003,N_19751,N_23008);
xnor U24004 (N_24004,N_21119,N_21789);
xnor U24005 (N_24005,N_18932,N_18069);
nor U24006 (N_24006,N_18638,N_23741);
nor U24007 (N_24007,N_18574,N_20960);
nor U24008 (N_24008,N_22556,N_19587);
nand U24009 (N_24009,N_20441,N_21678);
xor U24010 (N_24010,N_22560,N_20174);
xnor U24011 (N_24011,N_21208,N_18933);
nand U24012 (N_24012,N_20828,N_19914);
and U24013 (N_24013,N_22148,N_18377);
xor U24014 (N_24014,N_22321,N_23807);
nor U24015 (N_24015,N_18919,N_20758);
xor U24016 (N_24016,N_22827,N_19195);
and U24017 (N_24017,N_18428,N_22913);
nand U24018 (N_24018,N_22265,N_23345);
nand U24019 (N_24019,N_23956,N_20840);
xor U24020 (N_24020,N_19071,N_18668);
nand U24021 (N_24021,N_21090,N_20546);
nor U24022 (N_24022,N_21532,N_19208);
nor U24023 (N_24023,N_19786,N_19633);
or U24024 (N_24024,N_21377,N_20838);
nor U24025 (N_24025,N_22676,N_22071);
nand U24026 (N_24026,N_20710,N_21194);
nand U24027 (N_24027,N_23840,N_19827);
and U24028 (N_24028,N_20647,N_21612);
nor U24029 (N_24029,N_20851,N_22668);
nor U24030 (N_24030,N_23626,N_23953);
nand U24031 (N_24031,N_21530,N_18753);
or U24032 (N_24032,N_20900,N_22538);
nand U24033 (N_24033,N_21058,N_21742);
xnor U24034 (N_24034,N_19845,N_23274);
xnor U24035 (N_24035,N_20451,N_20107);
and U24036 (N_24036,N_22667,N_20494);
xnor U24037 (N_24037,N_19520,N_20037);
and U24038 (N_24038,N_23632,N_19931);
xnor U24039 (N_24039,N_21242,N_23365);
and U24040 (N_24040,N_21125,N_19872);
xor U24041 (N_24041,N_22109,N_22795);
nand U24042 (N_24042,N_20181,N_19625);
and U24043 (N_24043,N_19732,N_23570);
nor U24044 (N_24044,N_23236,N_23998);
xor U24045 (N_24045,N_23018,N_20527);
nand U24046 (N_24046,N_19535,N_23320);
nand U24047 (N_24047,N_22914,N_21739);
or U24048 (N_24048,N_20877,N_22871);
nand U24049 (N_24049,N_23708,N_22341);
xor U24050 (N_24050,N_20613,N_23916);
nor U24051 (N_24051,N_19362,N_20742);
nand U24052 (N_24052,N_18694,N_21093);
nand U24053 (N_24053,N_19151,N_18547);
or U24054 (N_24054,N_19248,N_18221);
xor U24055 (N_24055,N_19531,N_20652);
xnor U24056 (N_24056,N_22038,N_22610);
nor U24057 (N_24057,N_20166,N_23580);
nand U24058 (N_24058,N_23891,N_23778);
and U24059 (N_24059,N_20473,N_20731);
nand U24060 (N_24060,N_23042,N_19226);
and U24061 (N_24061,N_19129,N_18640);
and U24062 (N_24062,N_23392,N_20052);
nor U24063 (N_24063,N_21636,N_23828);
nand U24064 (N_24064,N_21223,N_19558);
and U24065 (N_24065,N_20621,N_22335);
and U24066 (N_24066,N_19238,N_21914);
xor U24067 (N_24067,N_19131,N_19037);
xor U24068 (N_24068,N_19705,N_19292);
and U24069 (N_24069,N_21958,N_21176);
nor U24070 (N_24070,N_22561,N_20588);
and U24071 (N_24071,N_21178,N_20283);
or U24072 (N_24072,N_21906,N_19398);
and U24073 (N_24073,N_22380,N_18661);
and U24074 (N_24074,N_18060,N_18861);
and U24075 (N_24075,N_23813,N_23865);
nand U24076 (N_24076,N_19820,N_18037);
xnor U24077 (N_24077,N_23808,N_22672);
xnor U24078 (N_24078,N_23093,N_22831);
nor U24079 (N_24079,N_19755,N_23881);
nand U24080 (N_24080,N_18670,N_22963);
and U24081 (N_24081,N_21140,N_21057);
nand U24082 (N_24082,N_18230,N_21306);
nor U24083 (N_24083,N_18154,N_22638);
or U24084 (N_24084,N_18837,N_21590);
or U24085 (N_24085,N_22081,N_21453);
or U24086 (N_24086,N_23521,N_18762);
and U24087 (N_24087,N_20693,N_19741);
nand U24088 (N_24088,N_19024,N_19726);
and U24089 (N_24089,N_21324,N_18350);
or U24090 (N_24090,N_18906,N_20247);
or U24091 (N_24091,N_20456,N_23974);
nor U24092 (N_24092,N_21620,N_23669);
nor U24093 (N_24093,N_22619,N_18282);
nor U24094 (N_24094,N_18359,N_23935);
nand U24095 (N_24095,N_19575,N_18871);
nor U24096 (N_24096,N_19361,N_22485);
nor U24097 (N_24097,N_21450,N_18092);
or U24098 (N_24098,N_23572,N_20250);
xor U24099 (N_24099,N_20899,N_21725);
and U24100 (N_24100,N_19404,N_20909);
nand U24101 (N_24101,N_23318,N_18335);
nor U24102 (N_24102,N_21696,N_18002);
xor U24103 (N_24103,N_20740,N_20753);
or U24104 (N_24104,N_22354,N_18626);
xnor U24105 (N_24105,N_18127,N_20244);
nor U24106 (N_24106,N_21128,N_18526);
nand U24107 (N_24107,N_21086,N_19018);
or U24108 (N_24108,N_21087,N_21505);
nor U24109 (N_24109,N_22030,N_21224);
or U24110 (N_24110,N_21776,N_19819);
nor U24111 (N_24111,N_19552,N_21977);
nand U24112 (N_24112,N_22091,N_18746);
nor U24113 (N_24113,N_21603,N_23887);
nand U24114 (N_24114,N_19977,N_21999);
nor U24115 (N_24115,N_23077,N_23114);
nor U24116 (N_24116,N_19472,N_18057);
xnor U24117 (N_24117,N_20605,N_21957);
nand U24118 (N_24118,N_21832,N_21391);
nand U24119 (N_24119,N_22877,N_18490);
nor U24120 (N_24120,N_22124,N_21764);
and U24121 (N_24121,N_22257,N_23243);
xnor U24122 (N_24122,N_18858,N_20395);
nor U24123 (N_24123,N_20552,N_22208);
nor U24124 (N_24124,N_21149,N_23455);
or U24125 (N_24125,N_20104,N_19034);
or U24126 (N_24126,N_18874,N_22823);
nand U24127 (N_24127,N_23343,N_18084);
xnor U24128 (N_24128,N_19893,N_23544);
xnor U24129 (N_24129,N_20866,N_20358);
nor U24130 (N_24130,N_19714,N_21415);
or U24131 (N_24131,N_21927,N_21010);
xor U24132 (N_24132,N_20919,N_22521);
nand U24133 (N_24133,N_23364,N_20574);
or U24134 (N_24134,N_20205,N_20331);
xnor U24135 (N_24135,N_21755,N_22494);
nand U24136 (N_24136,N_23086,N_22101);
and U24137 (N_24137,N_23208,N_23715);
xor U24138 (N_24138,N_19062,N_20821);
nand U24139 (N_24139,N_20614,N_23472);
xor U24140 (N_24140,N_18778,N_20080);
or U24141 (N_24141,N_23241,N_21947);
nor U24142 (N_24142,N_18340,N_23486);
or U24143 (N_24143,N_22622,N_18466);
or U24144 (N_24144,N_19859,N_22313);
and U24145 (N_24145,N_18672,N_19501);
nor U24146 (N_24146,N_22149,N_23456);
xor U24147 (N_24147,N_23100,N_23804);
nand U24148 (N_24148,N_19916,N_21627);
and U24149 (N_24149,N_18590,N_20106);
or U24150 (N_24150,N_23032,N_20564);
xnor U24151 (N_24151,N_18710,N_23940);
nand U24152 (N_24152,N_23805,N_21676);
and U24153 (N_24153,N_21289,N_21284);
nand U24154 (N_24154,N_20362,N_23589);
and U24155 (N_24155,N_23674,N_23245);
nand U24156 (N_24156,N_20910,N_18656);
nor U24157 (N_24157,N_18051,N_21826);
or U24158 (N_24158,N_20304,N_21451);
xor U24159 (N_24159,N_23185,N_18296);
nor U24160 (N_24160,N_22477,N_18579);
and U24161 (N_24161,N_18303,N_21080);
xnor U24162 (N_24162,N_23848,N_20912);
or U24163 (N_24163,N_18006,N_18387);
or U24164 (N_24164,N_19364,N_20102);
nor U24165 (N_24165,N_20890,N_18984);
nand U24166 (N_24166,N_19387,N_21235);
and U24167 (N_24167,N_23602,N_21979);
and U24168 (N_24168,N_21707,N_22966);
nor U24169 (N_24169,N_22520,N_21268);
nor U24170 (N_24170,N_23593,N_20987);
and U24171 (N_24171,N_18469,N_20369);
or U24172 (N_24172,N_23610,N_23846);
or U24173 (N_24173,N_19706,N_20415);
xnor U24174 (N_24174,N_22411,N_22403);
nand U24175 (N_24175,N_20095,N_23955);
nand U24176 (N_24176,N_23202,N_21965);
or U24177 (N_24177,N_23428,N_21897);
nand U24178 (N_24178,N_19298,N_20506);
and U24179 (N_24179,N_21386,N_22531);
xor U24180 (N_24180,N_18815,N_23514);
and U24181 (N_24181,N_23328,N_22533);
xor U24182 (N_24182,N_21746,N_18817);
and U24183 (N_24183,N_23225,N_23322);
or U24184 (N_24184,N_22625,N_21971);
and U24185 (N_24185,N_19624,N_19172);
nor U24186 (N_24186,N_22943,N_20022);
nor U24187 (N_24187,N_21133,N_19485);
xnor U24188 (N_24188,N_22969,N_22534);
nor U24189 (N_24189,N_18491,N_21003);
xnor U24190 (N_24190,N_23092,N_19224);
nand U24191 (N_24191,N_22734,N_23983);
or U24192 (N_24192,N_20285,N_18772);
nor U24193 (N_24193,N_20974,N_21805);
or U24194 (N_24194,N_20694,N_18610);
and U24195 (N_24195,N_19773,N_21720);
and U24196 (N_24196,N_18576,N_18417);
xnor U24197 (N_24197,N_23585,N_19425);
nand U24198 (N_24198,N_22474,N_22375);
nor U24199 (N_24199,N_20269,N_19943);
or U24200 (N_24200,N_21346,N_21271);
nor U24201 (N_24201,N_21218,N_22031);
and U24202 (N_24202,N_20785,N_20776);
or U24203 (N_24203,N_20975,N_23617);
xnor U24204 (N_24204,N_23188,N_20214);
nand U24205 (N_24205,N_23864,N_19489);
nand U24206 (N_24206,N_23137,N_21020);
nand U24207 (N_24207,N_21865,N_19384);
and U24208 (N_24208,N_18947,N_21232);
nand U24209 (N_24209,N_21626,N_23566);
or U24210 (N_24210,N_23221,N_18078);
nand U24211 (N_24211,N_18774,N_23298);
or U24212 (N_24212,N_19429,N_19942);
or U24213 (N_24213,N_23761,N_21082);
or U24214 (N_24214,N_19676,N_23317);
xnor U24215 (N_24215,N_19637,N_22329);
nor U24216 (N_24216,N_18599,N_19800);
nand U24217 (N_24217,N_19185,N_22242);
nand U24218 (N_24218,N_18929,N_22764);
and U24219 (N_24219,N_20745,N_23995);
nand U24220 (N_24220,N_18106,N_20423);
nand U24221 (N_24221,N_23116,N_23760);
xor U24222 (N_24222,N_21920,N_20841);
nand U24223 (N_24223,N_21097,N_19417);
xor U24224 (N_24224,N_21555,N_20813);
nand U24225 (N_24225,N_19342,N_18075);
and U24226 (N_24226,N_18558,N_18180);
nand U24227 (N_24227,N_23378,N_19781);
xor U24228 (N_24228,N_23847,N_22488);
or U24229 (N_24229,N_23128,N_18414);
nand U24230 (N_24230,N_23681,N_22654);
nor U24231 (N_24231,N_21989,N_23721);
nand U24232 (N_24232,N_19763,N_19116);
nor U24233 (N_24233,N_22805,N_18406);
or U24234 (N_24234,N_19979,N_20452);
or U24235 (N_24235,N_21238,N_18305);
nand U24236 (N_24236,N_18446,N_19405);
or U24237 (N_24237,N_23453,N_23573);
nor U24238 (N_24238,N_20935,N_18704);
or U24239 (N_24239,N_22527,N_22597);
nor U24240 (N_24240,N_21770,N_23078);
and U24241 (N_24241,N_18872,N_22153);
xnor U24242 (N_24242,N_23301,N_19385);
xnor U24243 (N_24243,N_20780,N_23101);
nor U24244 (N_24244,N_23764,N_20077);
nand U24245 (N_24245,N_18701,N_20000);
nor U24246 (N_24246,N_22884,N_21435);
xnor U24247 (N_24247,N_23199,N_18214);
nand U24248 (N_24248,N_18429,N_23145);
and U24249 (N_24249,N_20970,N_20504);
and U24250 (N_24250,N_18512,N_20595);
nand U24251 (N_24251,N_20053,N_22199);
nand U24252 (N_24252,N_19414,N_18380);
or U24253 (N_24253,N_21602,N_19158);
nand U24254 (N_24254,N_18038,N_22739);
and U24255 (N_24255,N_22318,N_20992);
and U24256 (N_24256,N_18164,N_21073);
nor U24257 (N_24257,N_23920,N_18487);
xor U24258 (N_24258,N_19794,N_18373);
or U24259 (N_24259,N_23526,N_19210);
and U24260 (N_24260,N_20123,N_22180);
nor U24261 (N_24261,N_23506,N_23495);
nand U24262 (N_24262,N_21605,N_22054);
and U24263 (N_24263,N_18244,N_21356);
xnor U24264 (N_24264,N_19117,N_20179);
or U24265 (N_24265,N_18751,N_23105);
xnor U24266 (N_24266,N_21436,N_20528);
xnor U24267 (N_24267,N_22925,N_18993);
nor U24268 (N_24268,N_20925,N_18935);
nand U24269 (N_24269,N_22789,N_18844);
xnor U24270 (N_24270,N_19019,N_21189);
nor U24271 (N_24271,N_22506,N_22684);
or U24272 (N_24272,N_19936,N_23286);
nor U24273 (N_24273,N_20117,N_21348);
and U24274 (N_24274,N_23978,N_19402);
nor U24275 (N_24275,N_19720,N_22338);
or U24276 (N_24276,N_21181,N_21623);
nand U24277 (N_24277,N_19344,N_20183);
nor U24278 (N_24278,N_19275,N_21515);
nand U24279 (N_24279,N_20539,N_18855);
nor U24280 (N_24280,N_21582,N_23487);
xnor U24281 (N_24281,N_18012,N_22922);
nand U24282 (N_24282,N_23303,N_18344);
xor U24283 (N_24283,N_18528,N_23753);
or U24284 (N_24284,N_19834,N_23664);
or U24285 (N_24285,N_21031,N_22295);
or U24286 (N_24286,N_21477,N_19271);
or U24287 (N_24287,N_20884,N_21601);
nor U24288 (N_24288,N_22733,N_19454);
xnor U24289 (N_24289,N_23903,N_21514);
nand U24290 (N_24290,N_21823,N_21731);
or U24291 (N_24291,N_22365,N_20553);
xor U24292 (N_24292,N_22077,N_19696);
or U24293 (N_24293,N_22432,N_23996);
nand U24294 (N_24294,N_22113,N_19270);
or U24295 (N_24295,N_20701,N_21970);
and U24296 (N_24296,N_18337,N_18828);
nand U24297 (N_24297,N_19369,N_23701);
xor U24298 (N_24298,N_19747,N_21682);
nor U24299 (N_24299,N_20522,N_21196);
and U24300 (N_24300,N_22026,N_23750);
or U24301 (N_24301,N_20986,N_21323);
or U24302 (N_24302,N_21816,N_18827);
nand U24303 (N_24303,N_18111,N_19801);
nor U24304 (N_24304,N_23464,N_23704);
nor U24305 (N_24305,N_22784,N_22260);
and U24306 (N_24306,N_18684,N_20837);
or U24307 (N_24307,N_23922,N_20068);
nor U24308 (N_24308,N_23130,N_22108);
or U24309 (N_24309,N_18620,N_20435);
nor U24310 (N_24310,N_19951,N_23169);
or U24311 (N_24311,N_20825,N_19709);
nand U24312 (N_24312,N_21632,N_21597);
nor U24313 (N_24313,N_22949,N_23400);
nand U24314 (N_24314,N_21358,N_18560);
or U24315 (N_24315,N_18705,N_18980);
nand U24316 (N_24316,N_22767,N_20118);
and U24317 (N_24317,N_19086,N_22110);
and U24318 (N_24318,N_22829,N_19687);
or U24319 (N_24319,N_19016,N_21290);
and U24320 (N_24320,N_19081,N_20251);
xor U24321 (N_24321,N_19498,N_18200);
nand U24322 (N_24322,N_23494,N_21220);
xnor U24323 (N_24323,N_23280,N_21750);
nor U24324 (N_24324,N_23296,N_19320);
nand U24325 (N_24325,N_18259,N_21963);
nor U24326 (N_24326,N_18114,N_20446);
nand U24327 (N_24327,N_19874,N_22256);
and U24328 (N_24328,N_23608,N_23515);
nor U24329 (N_24329,N_19846,N_20140);
nand U24330 (N_24330,N_19043,N_22117);
and U24331 (N_24331,N_22443,N_19124);
nand U24332 (N_24332,N_21596,N_22107);
nand U24333 (N_24333,N_18866,N_18109);
and U24334 (N_24334,N_20904,N_21146);
and U24335 (N_24335,N_18464,N_22118);
nor U24336 (N_24336,N_19045,N_19412);
and U24337 (N_24337,N_20718,N_23260);
or U24338 (N_24338,N_22544,N_23888);
and U24339 (N_24339,N_18156,N_20346);
nor U24340 (N_24340,N_18407,N_18291);
nand U24341 (N_24341,N_22603,N_20071);
nand U24342 (N_24342,N_21240,N_20157);
nor U24343 (N_24343,N_22841,N_18554);
or U24344 (N_24344,N_23710,N_23174);
and U24345 (N_24345,N_20526,N_20254);
and U24346 (N_24346,N_18478,N_21966);
or U24347 (N_24347,N_22004,N_21408);
xor U24348 (N_24348,N_20803,N_21420);
or U24349 (N_24349,N_22097,N_19666);
or U24350 (N_24350,N_22919,N_18323);
nand U24351 (N_24351,N_18176,N_21649);
nor U24352 (N_24352,N_21646,N_22170);
nor U24353 (N_24353,N_20727,N_19980);
and U24354 (N_24354,N_20099,N_21318);
or U24355 (N_24355,N_21634,N_22898);
or U24356 (N_24356,N_18687,N_21428);
nand U24357 (N_24357,N_20115,N_22591);
xor U24358 (N_24358,N_22896,N_18826);
xor U24359 (N_24359,N_22349,N_18249);
and U24360 (N_24360,N_22612,N_23861);
or U24361 (N_24361,N_20228,N_18669);
nor U24362 (N_24362,N_23450,N_20062);
xor U24363 (N_24363,N_20924,N_18890);
or U24364 (N_24364,N_23779,N_20516);
nor U24365 (N_24365,N_20755,N_22950);
nor U24366 (N_24366,N_19083,N_19850);
and U24367 (N_24367,N_20902,N_19830);
or U24368 (N_24368,N_19728,N_19486);
or U24369 (N_24369,N_19659,N_21354);
nand U24370 (N_24370,N_21166,N_21831);
nand U24371 (N_24371,N_19833,N_18067);
xnor U24372 (N_24372,N_23801,N_22103);
nor U24373 (N_24373,N_23726,N_22759);
and U24374 (N_24374,N_18196,N_20592);
nand U24375 (N_24375,N_21369,N_23860);
nand U24376 (N_24376,N_22730,N_20268);
and U24377 (N_24377,N_22451,N_22195);
xor U24378 (N_24378,N_22156,N_23448);
or U24379 (N_24379,N_22053,N_20826);
or U24380 (N_24380,N_20420,N_20149);
and U24381 (N_24381,N_23393,N_21079);
xnor U24382 (N_24382,N_18227,N_20305);
nand U24383 (N_24383,N_22262,N_22027);
xnor U24384 (N_24384,N_23957,N_23478);
xnor U24385 (N_24385,N_19754,N_19099);
nor U24386 (N_24386,N_21017,N_21791);
nand U24387 (N_24387,N_22616,N_18907);
and U24388 (N_24388,N_22959,N_18723);
xor U24389 (N_24389,N_19765,N_18517);
or U24390 (N_24390,N_21987,N_21299);
and U24391 (N_24391,N_18631,N_23560);
nor U24392 (N_24392,N_19242,N_19536);
or U24393 (N_24393,N_23937,N_19592);
nand U24394 (N_24394,N_22366,N_18212);
and U24395 (N_24395,N_22300,N_20411);
nand U24396 (N_24396,N_22701,N_19388);
nand U24397 (N_24397,N_18801,N_18503);
and U24398 (N_24398,N_22674,N_20659);
or U24399 (N_24399,N_20044,N_23666);
and U24400 (N_24400,N_22742,N_18473);
nand U24401 (N_24401,N_23682,N_22441);
nand U24402 (N_24402,N_23465,N_18442);
nor U24403 (N_24403,N_20733,N_19875);
nor U24404 (N_24404,N_21004,N_20455);
or U24405 (N_24405,N_22412,N_18077);
or U24406 (N_24406,N_22413,N_19730);
nand U24407 (N_24407,N_22994,N_18880);
and U24408 (N_24408,N_21441,N_20615);
nor U24409 (N_24409,N_20543,N_18594);
xor U24410 (N_24410,N_20425,N_23789);
or U24411 (N_24411,N_22765,N_18525);
nand U24412 (N_24412,N_21007,N_23076);
nor U24413 (N_24413,N_20005,N_18535);
and U24414 (N_24414,N_18794,N_19492);
and U24415 (N_24415,N_20030,N_19574);
xnor U24416 (N_24416,N_18103,N_21661);
nor U24417 (N_24417,N_21933,N_19645);
or U24418 (N_24418,N_18636,N_20663);
xnor U24419 (N_24419,N_22137,N_18916);
or U24420 (N_24420,N_20233,N_23163);
or U24421 (N_24421,N_22279,N_21748);
nor U24422 (N_24422,N_19121,N_21278);
nor U24423 (N_24423,N_23786,N_18707);
nor U24424 (N_24424,N_19465,N_18737);
nor U24425 (N_24425,N_21468,N_18703);
nor U24426 (N_24426,N_18248,N_23177);
and U24427 (N_24427,N_22476,N_21366);
nand U24428 (N_24428,N_21098,N_23843);
and U24429 (N_24429,N_18729,N_18534);
nand U24430 (N_24430,N_18465,N_18110);
nor U24431 (N_24431,N_22897,N_20607);
nor U24432 (N_24432,N_20752,N_19608);
nor U24433 (N_24433,N_23231,N_18231);
nand U24434 (N_24434,N_19969,N_23477);
nor U24435 (N_24435,N_21263,N_19565);
and U24436 (N_24436,N_18496,N_20586);
nor U24437 (N_24437,N_20908,N_21738);
nor U24438 (N_24438,N_20790,N_19511);
or U24439 (N_24439,N_20449,N_22399);
xnor U24440 (N_24440,N_18046,N_23295);
xnor U24441 (N_24441,N_22188,N_21567);
nor U24442 (N_24442,N_22824,N_20507);
and U24443 (N_24443,N_22259,N_23915);
or U24444 (N_24444,N_22414,N_23223);
nand U24445 (N_24445,N_22992,N_22849);
xnor U24446 (N_24446,N_23201,N_19743);
or U24447 (N_24447,N_22294,N_20176);
and U24448 (N_24448,N_20532,N_22601);
xor U24449 (N_24449,N_22592,N_23745);
and U24450 (N_24450,N_20996,N_21355);
and U24451 (N_24451,N_21990,N_21206);
and U24452 (N_24452,N_23323,N_18619);
nand U24453 (N_24453,N_23905,N_19998);
and U24454 (N_24454,N_19550,N_19581);
or U24455 (N_24455,N_19601,N_22434);
and U24456 (N_24456,N_18218,N_22811);
xor U24457 (N_24457,N_23658,N_20128);
or U24458 (N_24458,N_23142,N_21295);
nor U24459 (N_24459,N_20643,N_18673);
and U24460 (N_24460,N_18008,N_21185);
xnor U24461 (N_24461,N_22198,N_19166);
and U24462 (N_24462,N_21398,N_22309);
nand U24463 (N_24463,N_23975,N_22859);
or U24464 (N_24464,N_23812,N_21138);
or U24465 (N_24465,N_22754,N_21373);
nand U24466 (N_24466,N_23548,N_20572);
and U24467 (N_24467,N_22721,N_18789);
nand U24468 (N_24468,N_21281,N_22808);
or U24469 (N_24469,N_18153,N_23149);
or U24470 (N_24470,N_22015,N_20823);
xor U24471 (N_24471,N_19988,N_19206);
and U24472 (N_24472,N_19340,N_18126);
and U24473 (N_24473,N_23562,N_22410);
xnor U24474 (N_24474,N_21875,N_18091);
and U24475 (N_24475,N_22082,N_19961);
and U24476 (N_24476,N_18531,N_22602);
nor U24477 (N_24477,N_23354,N_23001);
and U24478 (N_24478,N_20380,N_23522);
and U24479 (N_24479,N_18808,N_22007);
nand U24480 (N_24480,N_20193,N_18593);
xor U24481 (N_24481,N_22853,N_23278);
or U24482 (N_24482,N_20491,N_18299);
and U24483 (N_24483,N_23686,N_21903);
nor U24484 (N_24484,N_20016,N_19103);
nor U24485 (N_24485,N_21122,N_18210);
nor U24486 (N_24486,N_20338,N_20359);
nand U24487 (N_24487,N_21861,N_22394);
nand U24488 (N_24488,N_20301,N_22965);
xor U24489 (N_24489,N_18388,N_21615);
and U24490 (N_24490,N_21893,N_21491);
or U24491 (N_24491,N_22751,N_18199);
or U24492 (N_24492,N_21244,N_23319);
or U24493 (N_24493,N_22912,N_23230);
nand U24494 (N_24494,N_20941,N_19613);
and U24495 (N_24495,N_20299,N_21210);
nor U24496 (N_24496,N_23339,N_18327);
xnor U24497 (N_24497,N_19972,N_23061);
nand U24498 (N_24498,N_23437,N_21320);
nand U24499 (N_24499,N_22094,N_23834);
nand U24500 (N_24500,N_22356,N_19177);
and U24501 (N_24501,N_23341,N_21592);
xnor U24502 (N_24502,N_23370,N_19322);
nand U24503 (N_24503,N_20370,N_20688);
nand U24504 (N_24504,N_18168,N_22937);
xnor U24505 (N_24505,N_22726,N_20042);
or U24506 (N_24506,N_21280,N_22425);
nor U24507 (N_24507,N_19266,N_19758);
nor U24508 (N_24508,N_21810,N_18033);
nor U24509 (N_24509,N_22328,N_18149);
nand U24510 (N_24510,N_20195,N_22270);
or U24511 (N_24511,N_20843,N_20822);
xor U24512 (N_24512,N_18317,N_19904);
xnor U24513 (N_24513,N_18304,N_23979);
xnor U24514 (N_24514,N_20824,N_23820);
and U24515 (N_24515,N_23757,N_21302);
nand U24516 (N_24516,N_21099,N_22267);
or U24517 (N_24517,N_19767,N_18736);
nor U24518 (N_24518,N_23803,N_22307);
and U24519 (N_24519,N_23973,N_19047);
or U24520 (N_24520,N_23496,N_22161);
xor U24521 (N_24521,N_22090,N_21145);
nand U24522 (N_24522,N_19233,N_18765);
xnor U24523 (N_24523,N_18603,N_18097);
xor U24524 (N_24524,N_18328,N_19974);
xor U24525 (N_24525,N_21890,N_22646);
xor U24526 (N_24526,N_22910,N_18518);
xnor U24527 (N_24527,N_21454,N_21030);
nand U24528 (N_24528,N_21248,N_18957);
xor U24529 (N_24529,N_21889,N_21541);
nand U24530 (N_24530,N_22945,N_22505);
and U24531 (N_24531,N_19568,N_21873);
nand U24532 (N_24532,N_23438,N_21690);
or U24533 (N_24533,N_19029,N_23700);
nor U24534 (N_24534,N_18960,N_21591);
and U24535 (N_24535,N_23892,N_19986);
nor U24536 (N_24536,N_21011,N_21624);
nand U24537 (N_24537,N_22607,N_20121);
nand U24538 (N_24538,N_18489,N_23258);
nand U24539 (N_24539,N_21061,N_23748);
nand U24540 (N_24540,N_23615,N_18854);
nand U24541 (N_24541,N_22604,N_18454);
xnor U24542 (N_24542,N_20184,N_18974);
xor U24543 (N_24543,N_21940,N_23908);
nor U24544 (N_24544,N_19407,N_19219);
xor U24545 (N_24545,N_21719,N_18329);
and U24546 (N_24546,N_21846,N_18766);
nor U24547 (N_24547,N_19245,N_20146);
xor U24548 (N_24548,N_22814,N_19100);
nand U24549 (N_24549,N_23575,N_20559);
or U24550 (N_24550,N_23727,N_18133);
or U24551 (N_24551,N_23357,N_18612);
and U24552 (N_24552,N_20178,N_22878);
nand U24553 (N_24553,N_23129,N_19091);
nor U24554 (N_24554,N_23213,N_21884);
nand U24555 (N_24555,N_18015,N_18247);
nor U24556 (N_24556,N_22997,N_22885);
and U24557 (N_24557,N_23732,N_18194);
xnor U24558 (N_24558,N_18136,N_21536);
or U24559 (N_24559,N_22073,N_22128);
nor U24560 (N_24560,N_20063,N_20145);
and U24561 (N_24561,N_18811,N_18322);
or U24562 (N_24562,N_20073,N_19435);
and U24563 (N_24563,N_23007,N_20703);
nor U24564 (N_24564,N_22398,N_18404);
and U24565 (N_24565,N_18420,N_20798);
nand U24566 (N_24566,N_18076,N_19919);
xnor U24567 (N_24567,N_23087,N_23347);
xor U24568 (N_24568,N_21372,N_22725);
and U24569 (N_24569,N_23446,N_21419);
nor U24570 (N_24570,N_19863,N_19261);
and U24571 (N_24571,N_23556,N_23876);
nor U24572 (N_24572,N_23907,N_23108);
nor U24573 (N_24573,N_22968,N_23046);
nand U24574 (N_24574,N_18026,N_23749);
and U24575 (N_24575,N_23103,N_22496);
nor U24576 (N_24576,N_23716,N_21313);
and U24577 (N_24577,N_22722,N_19188);
nand U24578 (N_24578,N_23967,N_22327);
or U24579 (N_24579,N_21492,N_22526);
xor U24580 (N_24580,N_19842,N_21053);
nor U24581 (N_24581,N_23404,N_20982);
xor U24582 (N_24582,N_21132,N_22627);
and U24583 (N_24583,N_19354,N_22803);
and U24584 (N_24584,N_19821,N_22855);
xor U24585 (N_24585,N_21216,N_22301);
nor U24586 (N_24586,N_21766,N_18949);
xor U24587 (N_24587,N_20616,N_20445);
nand U24588 (N_24588,N_21397,N_23259);
or U24589 (N_24589,N_22500,N_21363);
and U24590 (N_24590,N_20662,N_23394);
or U24591 (N_24591,N_22344,N_20778);
xor U24592 (N_24592,N_19675,N_23667);
xnor U24593 (N_24593,N_21853,N_18839);
xnor U24594 (N_24594,N_22863,N_19964);
nand U24595 (N_24595,N_21174,N_21085);
nand U24596 (N_24596,N_18403,N_22315);
nand U24597 (N_24597,N_23889,N_19890);
and U24598 (N_24598,N_22392,N_18102);
nand U24599 (N_24599,N_18664,N_18901);
nor U24600 (N_24600,N_19949,N_20221);
and U24601 (N_24601,N_18800,N_23707);
nor U24602 (N_24602,N_18742,N_21201);
and U24603 (N_24603,N_19074,N_19693);
and U24604 (N_24604,N_19562,N_20421);
and U24605 (N_24605,N_23187,N_19391);
xnor U24606 (N_24606,N_21230,N_22450);
and U24607 (N_24607,N_22005,N_20332);
nand U24608 (N_24608,N_21411,N_22956);
and U24609 (N_24609,N_22426,N_22284);
nand U24610 (N_24610,N_18345,N_22881);
nand U24611 (N_24611,N_21301,N_21384);
xnor U24612 (N_24612,N_19522,N_22792);
nor U24613 (N_24613,N_19283,N_20460);
nor U24614 (N_24614,N_20101,N_20897);
nand U24615 (N_24615,N_20590,N_20517);
xor U24616 (N_24616,N_21055,N_23338);
nand U24617 (N_24617,N_19569,N_22570);
xor U24618 (N_24618,N_20352,N_19680);
and U24619 (N_24619,N_18274,N_18970);
and U24620 (N_24620,N_18155,N_19418);
or U24621 (N_24621,N_22858,N_18159);
nand U24622 (N_24622,N_21150,N_18927);
nand U24623 (N_24623,N_20011,N_18271);
and U24624 (N_24624,N_21692,N_19718);
nor U24625 (N_24625,N_21362,N_21467);
or U24626 (N_24626,N_19918,N_21364);
or U24627 (N_24627,N_20867,N_20886);
nor U24628 (N_24628,N_23479,N_22155);
nor U24629 (N_24629,N_21184,N_18569);
nand U24630 (N_24630,N_23449,N_19753);
or U24631 (N_24631,N_20713,N_22981);
or U24632 (N_24632,N_18883,N_21399);
nor U24633 (N_24633,N_18183,N_19220);
nor U24634 (N_24634,N_23759,N_21691);
or U24635 (N_24635,N_21629,N_18019);
and U24636 (N_24636,N_21907,N_18522);
nor U24637 (N_24637,N_23299,N_18470);
and U24638 (N_24638,N_23467,N_23968);
nand U24639 (N_24639,N_22138,N_22840);
nand U24640 (N_24640,N_19922,N_23794);
or U24641 (N_24641,N_22184,N_22483);
nor U24642 (N_24642,N_20751,N_22369);
or U24643 (N_24643,N_21833,N_19406);
and U24644 (N_24644,N_20386,N_18847);
or U24645 (N_24645,N_23567,N_19699);
and U24646 (N_24646,N_22246,N_22455);
xor U24647 (N_24647,N_23070,N_20576);
nand U24648 (N_24648,N_19189,N_19110);
or U24649 (N_24649,N_20880,N_19987);
nor U24650 (N_24650,N_22115,N_21533);
or U24651 (N_24651,N_18193,N_22554);
xor U24652 (N_24652,N_18734,N_20189);
nand U24653 (N_24653,N_21167,N_21155);
nor U24654 (N_24654,N_18910,N_22288);
or U24655 (N_24655,N_21400,N_19416);
and U24656 (N_24656,N_20217,N_22704);
or U24657 (N_24657,N_19810,N_19128);
and U24658 (N_24658,N_20271,N_18898);
nor U24659 (N_24659,N_23508,N_18860);
and U24660 (N_24660,N_23882,N_22715);
xnor U24661 (N_24661,N_23665,N_20515);
xor U24662 (N_24662,N_19307,N_20914);
or U24663 (N_24663,N_18978,N_21429);
nor U24664 (N_24664,N_21276,N_18058);
and U24665 (N_24665,N_19036,N_20671);
nand U24666 (N_24666,N_19735,N_18318);
or U24667 (N_24667,N_21665,N_20505);
or U24668 (N_24668,N_19791,N_20918);
nor U24669 (N_24669,N_21677,N_18875);
nor U24670 (N_24670,N_22633,N_18676);
nor U24671 (N_24671,N_23513,N_21034);
and U24672 (N_24672,N_19347,N_21941);
and U24673 (N_24673,N_18920,N_21382);
nand U24674 (N_24674,N_22333,N_19858);
nor U24675 (N_24675,N_20480,N_18394);
nand U24676 (N_24676,N_19304,N_22537);
nand U24677 (N_24677,N_22218,N_19328);
and U24678 (N_24678,N_21885,N_20608);
and U24679 (N_24679,N_19490,N_23057);
and U24680 (N_24680,N_19211,N_20997);
or U24681 (N_24681,N_19123,N_18879);
nand U24682 (N_24682,N_23747,N_21942);
xnor U24683 (N_24683,N_20865,N_19902);
nand U24684 (N_24684,N_18511,N_22206);
nor U24685 (N_24685,N_22221,N_18617);
and U24686 (N_24686,N_19315,N_19748);
nand U24687 (N_24687,N_20227,N_22021);
or U24688 (N_24688,N_20131,N_22942);
and U24689 (N_24689,N_23895,N_20839);
and U24690 (N_24690,N_21552,N_22193);
xor U24691 (N_24691,N_19032,N_18650);
nor U24692 (N_24692,N_22429,N_21123);
xor U24693 (N_24693,N_18205,N_19707);
nor U24694 (N_24694,N_23257,N_22144);
nor U24695 (N_24695,N_18791,N_19860);
nand U24696 (N_24696,N_22177,N_23835);
xor U24697 (N_24697,N_18792,N_19213);
or U24698 (N_24698,N_21736,N_22706);
and U24699 (N_24699,N_23498,N_20264);
and U24700 (N_24700,N_22377,N_23244);
xor U24701 (N_24701,N_21153,N_18251);
and U24702 (N_24702,N_20855,N_22179);
or U24703 (N_24703,N_22675,N_19737);
and U24704 (N_24704,N_22711,N_19638);
nand U24705 (N_24705,N_20130,N_23737);
nor U24706 (N_24706,N_18148,N_18439);
xnor U24707 (N_24707,N_22799,N_21422);
and U24708 (N_24708,N_21266,N_18530);
or U24709 (N_24709,N_18787,N_18288);
nand U24710 (N_24710,N_20397,N_23558);
or U24711 (N_24711,N_22486,N_20817);
nand U24712 (N_24712,N_18853,N_20223);
xor U24713 (N_24713,N_19255,N_20567);
and U24714 (N_24714,N_21482,N_18966);
xor U24715 (N_24715,N_18977,N_22281);
nor U24716 (N_24716,N_22475,N_20679);
and U24717 (N_24717,N_19869,N_22866);
nand U24718 (N_24718,N_20220,N_20470);
or U24719 (N_24719,N_22013,N_19857);
and U24720 (N_24720,N_22807,N_23836);
or U24721 (N_24721,N_21891,N_21430);
nor U24722 (N_24722,N_19186,N_20012);
xor U24723 (N_24723,N_20313,N_18697);
and U24724 (N_24724,N_19596,N_21250);
nand U24725 (N_24725,N_20490,N_20632);
or U24726 (N_24726,N_21745,N_20045);
nor U24727 (N_24727,N_23977,N_18059);
nand U24728 (N_24728,N_23268,N_20373);
nor U24729 (N_24729,N_23647,N_18257);
xor U24730 (N_24730,N_22655,N_19906);
nand U24731 (N_24731,N_23734,N_18688);
xor U24732 (N_24732,N_18588,N_20674);
nor U24733 (N_24733,N_20498,N_22174);
nand U24734 (N_24734,N_18198,N_23170);
xor U24735 (N_24735,N_21568,N_18877);
nand U24736 (N_24736,N_23389,N_23943);
or U24737 (N_24737,N_22162,N_20579);
and U24738 (N_24738,N_19031,N_23629);
nand U24739 (N_24739,N_20262,N_23332);
and U24740 (N_24740,N_19620,N_22692);
and U24741 (N_24741,N_20198,N_23703);
and U24742 (N_24742,N_18398,N_21863);
or U24743 (N_24743,N_22691,N_19983);
nor U24744 (N_24744,N_23773,N_21688);
nand U24745 (N_24745,N_23754,N_18743);
or U24746 (N_24746,N_21950,N_19618);
xnor U24747 (N_24747,N_18698,N_18510);
nand U24748 (N_24748,N_21304,N_23186);
nand U24749 (N_24749,N_18911,N_21587);
xor U24750 (N_24750,N_21895,N_23429);
xnor U24751 (N_24751,N_20770,N_21506);
and U24752 (N_24752,N_23926,N_20619);
nand U24753 (N_24753,N_22253,N_22034);
nand U24754 (N_24754,N_19355,N_20348);
or U24755 (N_24755,N_22551,N_23797);
and U24756 (N_24756,N_20800,N_20158);
and U24757 (N_24757,N_19816,N_20809);
xnor U24758 (N_24758,N_23194,N_20226);
and U24759 (N_24759,N_23636,N_22029);
and U24760 (N_24760,N_22543,N_19133);
and U24761 (N_24761,N_18174,N_18452);
xnor U24762 (N_24762,N_21817,N_20609);
or U24763 (N_24763,N_18041,N_23536);
nor U24764 (N_24764,N_19524,N_22009);
and U24765 (N_24765,N_19104,N_18566);
nor U24766 (N_24766,N_18754,N_19090);
or U24767 (N_24767,N_22583,N_18456);
or U24768 (N_24768,N_22480,N_19333);
xnor U24769 (N_24769,N_20029,N_21949);
or U24770 (N_24770,N_19168,N_23550);
and U24771 (N_24771,N_21417,N_20891);
nor U24772 (N_24772,N_18460,N_23997);
or U24773 (N_24773,N_22067,N_19715);
or U24774 (N_24774,N_20623,N_23413);
and U24775 (N_24775,N_21837,N_22843);
xnor U24776 (N_24776,N_21385,N_23063);
nor U24777 (N_24777,N_19779,N_21735);
nor U24778 (N_24778,N_22409,N_20635);
nand U24779 (N_24779,N_19507,N_21621);
nand U24780 (N_24780,N_20015,N_20510);
nor U24781 (N_24781,N_18175,N_23255);
nand U24782 (N_24782,N_20807,N_22016);
nor U24783 (N_24783,N_20775,N_18341);
xor U24784 (N_24784,N_19900,N_19263);
or U24785 (N_24785,N_20212,N_23796);
nor U24786 (N_24786,N_21239,N_22947);
or U24787 (N_24787,N_19973,N_20883);
nand U24788 (N_24788,N_23688,N_23021);
and U24789 (N_24789,N_23503,N_20293);
nand U24790 (N_24790,N_21813,N_23982);
xor U24791 (N_24791,N_19147,N_19360);
xnor U24792 (N_24792,N_19180,N_21352);
nor U24793 (N_24793,N_21209,N_23986);
and U24794 (N_24794,N_22139,N_23618);
or U24795 (N_24795,N_20916,N_21535);
nor U24796 (N_24796,N_22984,N_23578);
and U24797 (N_24797,N_18894,N_18628);
nor U24798 (N_24798,N_21874,N_23770);
or U24799 (N_24799,N_22615,N_21148);
and U24800 (N_24800,N_23403,N_22360);
or U24801 (N_24801,N_18505,N_21291);
or U24802 (N_24802,N_22471,N_20261);
or U24803 (N_24803,N_18731,N_18838);
and U24804 (N_24804,N_19898,N_23527);
or U24805 (N_24805,N_21074,N_22276);
xnor U24806 (N_24806,N_22647,N_20139);
or U24807 (N_24807,N_21456,N_22192);
nor U24808 (N_24808,N_18217,N_19027);
nor U24809 (N_24809,N_19957,N_20190);
nand U24810 (N_24810,N_23082,N_19997);
xnor U24811 (N_24811,N_18805,N_18598);
nand U24812 (N_24812,N_20137,N_19108);
nor U24813 (N_24813,N_23352,N_21558);
and U24814 (N_24814,N_21464,N_22908);
and U24815 (N_24815,N_22286,N_22364);
nand U24816 (N_24816,N_23219,N_22820);
nor U24817 (N_24817,N_19035,N_22347);
nor U24818 (N_24818,N_21262,N_22439);
xnor U24819 (N_24819,N_20860,N_22355);
nand U24820 (N_24820,N_22771,N_20874);
xnor U24821 (N_24821,N_21513,N_18747);
nand U24822 (N_24822,N_23633,N_21820);
nand U24823 (N_24823,N_23502,N_18497);
nand U24824 (N_24824,N_21797,N_20151);
or U24825 (N_24825,N_20169,N_20236);
or U24826 (N_24826,N_22059,N_22651);
nand U24827 (N_24827,N_23696,N_18649);
nand U24828 (N_24828,N_20013,N_21576);
and U24829 (N_24829,N_19589,N_20951);
nand U24830 (N_24830,N_18483,N_18381);
nand U24831 (N_24831,N_21159,N_18072);
nor U24832 (N_24832,N_22417,N_22158);
or U24833 (N_24833,N_23226,N_23156);
nor U24834 (N_24834,N_22268,N_23396);
xor U24835 (N_24835,N_18029,N_19139);
nor U24836 (N_24836,N_20161,N_18130);
and U24837 (N_24837,N_22043,N_19366);
nand U24838 (N_24838,N_19198,N_23099);
and U24839 (N_24839,N_21493,N_21782);
nand U24840 (N_24840,N_21215,N_19837);
and U24841 (N_24841,N_23985,N_23084);
nor U24842 (N_24842,N_18492,N_19835);
and U24843 (N_24843,N_20351,N_18975);
or U24844 (N_24844,N_19590,N_23565);
or U24845 (N_24845,N_19636,N_21642);
xnor U24846 (N_24846,N_19525,N_19382);
and U24847 (N_24847,N_22975,N_20509);
nor U24848 (N_24848,N_22982,N_23972);
or U24849 (N_24849,N_21573,N_21508);
or U24850 (N_24850,N_19650,N_18397);
nor U24851 (N_24851,N_23068,N_20644);
nand U24852 (N_24852,N_23172,N_21062);
nor U24853 (N_24853,N_23969,N_23557);
nor U24854 (N_24854,N_18504,N_19991);
xor U24855 (N_24855,N_18609,N_23981);
xnor U24856 (N_24856,N_18551,N_22991);
nor U24857 (N_24857,N_23564,N_23746);
xnor U24858 (N_24858,N_19771,N_18124);
xnor U24859 (N_24859,N_19125,N_23235);
nor U24860 (N_24860,N_23426,N_20756);
or U24861 (N_24861,N_19910,N_20938);
or U24862 (N_24862,N_21653,N_22447);
xnor U24863 (N_24863,N_23175,N_19156);
nand U24864 (N_24864,N_21469,N_21254);
or U24865 (N_24865,N_18632,N_21279);
or U24866 (N_24866,N_20281,N_23401);
xor U24867 (N_24867,N_20991,N_23432);
xor U24868 (N_24868,N_19729,N_18261);
nand U24869 (N_24869,N_23288,N_21234);
or U24870 (N_24870,N_23273,N_22572);
or U24871 (N_24871,N_23291,N_21437);
or U24872 (N_24872,N_18131,N_23962);
nor U24873 (N_24873,N_23272,N_22794);
nor U24874 (N_24874,N_19383,N_18434);
nand U24875 (N_24875,N_22497,N_19892);
nor U24876 (N_24876,N_20722,N_23736);
or U24877 (N_24877,N_18400,N_21969);
xor U24878 (N_24878,N_23081,N_20861);
nand U24879 (N_24879,N_20114,N_18824);
xor U24880 (N_24880,N_19514,N_19742);
or U24881 (N_24881,N_23980,N_23326);
and U24882 (N_24882,N_21758,N_22490);
and U24883 (N_24883,N_23509,N_18655);
and U24884 (N_24884,N_18453,N_19202);
nand U24885 (N_24885,N_22744,N_23661);
xor U24886 (N_24886,N_20669,N_21319);
xor U24887 (N_24887,N_20296,N_23520);
and U24888 (N_24888,N_19374,N_22428);
nor U24889 (N_24889,N_22879,N_23609);
and U24890 (N_24890,N_23152,N_20993);
nand U24891 (N_24891,N_18633,N_21656);
and U24892 (N_24892,N_21257,N_19394);
xor U24893 (N_24893,N_20606,N_19978);
xor U24894 (N_24894,N_19686,N_23096);
xor U24895 (N_24895,N_20372,N_19537);
or U24896 (N_24896,N_23676,N_22277);
xnor U24897 (N_24897,N_20932,N_19646);
xor U24898 (N_24898,N_23038,N_19331);
or U24899 (N_24899,N_21680,N_19829);
nor U24900 (N_24900,N_20625,N_22920);
and U24901 (N_24901,N_20468,N_22740);
or U24902 (N_24902,N_18237,N_19175);
and U24903 (N_24903,N_22890,N_21075);
or U24904 (N_24904,N_21439,N_21842);
and U24905 (N_24905,N_22011,N_22130);
and U24906 (N_24906,N_19216,N_22217);
nor U24907 (N_24907,N_21497,N_22070);
nor U24908 (N_24908,N_18413,N_23991);
and U24909 (N_24909,N_22317,N_18533);
nand U24910 (N_24910,N_22785,N_18981);
xor U24911 (N_24911,N_18963,N_21229);
and U24912 (N_24912,N_19738,N_21781);
xor U24913 (N_24913,N_19824,N_20524);
nor U24914 (N_24914,N_18475,N_23525);
nand U24915 (N_24915,N_19477,N_22463);
nand U24916 (N_24916,N_20170,N_23947);
and U24917 (N_24917,N_20654,N_21396);
xor U24918 (N_24918,N_20006,N_19795);
xnor U24919 (N_24919,N_23823,N_18378);
nand U24920 (N_24920,N_18347,N_20942);
or U24921 (N_24921,N_19703,N_23954);
nor U24922 (N_24922,N_20347,N_20802);
and U24923 (N_24923,N_18708,N_19566);
xnor U24924 (N_24924,N_22899,N_23859);
nand U24925 (N_24925,N_19867,N_23841);
and U24926 (N_24926,N_22778,N_20252);
xnor U24927 (N_24927,N_20126,N_22430);
or U24928 (N_24928,N_19504,N_18733);
nor U24929 (N_24929,N_20234,N_19966);
or U24930 (N_24930,N_20599,N_22076);
xor U24931 (N_24931,N_22816,N_19411);
nor U24932 (N_24932,N_20804,N_19349);
xor U24933 (N_24933,N_18147,N_19619);
nand U24934 (N_24934,N_20278,N_18294);
nand U24935 (N_24935,N_18188,N_21054);
or U24936 (N_24936,N_19609,N_23049);
nand U24937 (N_24937,N_18285,N_21882);
nand U24938 (N_24938,N_20458,N_22553);
or U24939 (N_24939,N_21066,N_20858);
or U24940 (N_24940,N_20994,N_23706);
nand U24941 (N_24941,N_18457,N_19309);
xor U24942 (N_24942,N_19050,N_18793);
nor U24943 (N_24943,N_22786,N_23546);
and U24944 (N_24944,N_20896,N_20556);
and U24945 (N_24945,N_20229,N_19232);
nand U24946 (N_24946,N_20469,N_20092);
or U24947 (N_24947,N_23927,N_22850);
or U24948 (N_24948,N_19480,N_20152);
nand U24949 (N_24949,N_20335,N_19368);
nand U24950 (N_24950,N_18467,N_21211);
nand U24951 (N_24951,N_18190,N_20008);
or U24952 (N_24952,N_18342,N_21542);
and U24953 (N_24953,N_22530,N_19030);
nor U24954 (N_24954,N_18266,N_18495);
nand U24955 (N_24955,N_18462,N_18252);
nor U24956 (N_24956,N_19434,N_21892);
xor U24957 (N_24957,N_18421,N_23097);
or U24958 (N_24958,N_20364,N_23089);
nand U24959 (N_24959,N_23713,N_18438);
or U24960 (N_24960,N_20967,N_22507);
and U24961 (N_24961,N_18234,N_18211);
nor U24962 (N_24962,N_23601,N_18788);
xor U24963 (N_24963,N_22516,N_19994);
nand U24964 (N_24964,N_20878,N_21470);
and U24965 (N_24965,N_18739,N_23333);
and U24966 (N_24966,N_22469,N_19150);
nor U24967 (N_24967,N_20622,N_21860);
nand U24968 (N_24968,N_23242,N_19629);
or U24969 (N_24969,N_23549,N_18870);
or U24970 (N_24970,N_21198,N_20280);
nor U24971 (N_24971,N_19111,N_21625);
xnor U24972 (N_24972,N_18396,N_23409);
and U24973 (N_24973,N_19319,N_22938);
nor U24974 (N_24974,N_22577,N_22882);
nand U24975 (N_24975,N_23368,N_19757);
nor U24976 (N_24976,N_21617,N_23936);
and U24977 (N_24977,N_22391,N_20219);
and U24978 (N_24978,N_18773,N_20735);
nor U24979 (N_24979,N_21664,N_22126);
nand U24980 (N_24980,N_18135,N_22946);
and U24981 (N_24981,N_19488,N_21855);
nor U24982 (N_24982,N_20665,N_19170);
xor U24983 (N_24983,N_18309,N_22175);
nor U24984 (N_24984,N_20591,N_23144);
nor U24985 (N_24985,N_23470,N_21780);
nor U24986 (N_24986,N_22694,N_19199);
xor U24987 (N_24987,N_23543,N_21442);
xnor U24988 (N_24988,N_22387,N_19926);
nand U24989 (N_24989,N_19264,N_22974);
and U24990 (N_24990,N_23949,N_18399);
xor U24991 (N_24991,N_18863,N_18690);
nand U24992 (N_24992,N_20485,N_19612);
and U24993 (N_24993,N_21272,N_22585);
nand U24994 (N_24994,N_18757,N_22269);
or U24995 (N_24995,N_19812,N_21338);
and U24996 (N_24996,N_19022,N_22631);
nand U24997 (N_24997,N_22003,N_22185);
and U24998 (N_24998,N_23771,N_22686);
and U24999 (N_24999,N_23507,N_20569);
or U25000 (N_25000,N_22901,N_21881);
and U25001 (N_25001,N_22834,N_18021);
and U25002 (N_25002,N_18937,N_21027);
or U25003 (N_25003,N_23646,N_23388);
and U25004 (N_25004,N_21701,N_23184);
and U25005 (N_25005,N_18151,N_22420);
nand U25006 (N_25006,N_20738,N_19948);
and U25007 (N_25007,N_23862,N_21849);
or U25008 (N_25008,N_20438,N_21565);
and U25009 (N_25009,N_22001,N_20082);
xor U25010 (N_25010,N_23483,N_23657);
xor U25011 (N_25011,N_18823,N_19467);
or U25012 (N_25012,N_18922,N_22049);
or U25013 (N_25013,N_21197,N_18843);
nor U25014 (N_25014,N_21964,N_21670);
nand U25015 (N_25015,N_18727,N_23304);
and U25016 (N_25016,N_22745,N_22573);
nand U25017 (N_25017,N_18562,N_19377);
xor U25018 (N_25018,N_23002,N_22642);
or U25019 (N_25019,N_20716,N_23112);
and U25020 (N_25020,N_19844,N_21870);
and U25021 (N_25021,N_18463,N_19378);
and U25022 (N_25022,N_19886,N_18865);
xnor U25023 (N_25023,N_19431,N_22703);
and U25024 (N_25024,N_23869,N_21529);
nor U25025 (N_25025,N_19513,N_23181);
or U25026 (N_25026,N_18436,N_19300);
nor U25027 (N_25027,N_19146,N_20396);
or U25028 (N_25028,N_19343,N_23497);
nand U25029 (N_25029,N_18129,N_22934);
xor U25030 (N_25030,N_20225,N_19097);
and U25031 (N_25031,N_22986,N_21406);
and U25032 (N_25032,N_19677,N_18419);
nand U25033 (N_25033,N_18158,N_21858);
nand U25034 (N_25034,N_18343,N_18166);
and U25035 (N_25035,N_20862,N_22735);
nor U25036 (N_25036,N_23003,N_19359);
or U25037 (N_25037,N_23381,N_18013);
nand U25038 (N_25038,N_19579,N_19237);
or U25039 (N_25039,N_21345,N_22641);
xnor U25040 (N_25040,N_20700,N_18351);
and U25041 (N_25041,N_23029,N_20026);
nand U25042 (N_25042,N_22624,N_20789);
or U25043 (N_25043,N_23033,N_23534);
xnor U25044 (N_25044,N_22903,N_18964);
or U25045 (N_25045,N_20536,N_20061);
or U25046 (N_25046,N_19471,N_21800);
nand U25047 (N_25047,N_19105,N_20450);
nor U25048 (N_25048,N_21489,N_21259);
or U25049 (N_25049,N_19815,N_19351);
or U25050 (N_25050,N_19792,N_19784);
and U25051 (N_25051,N_21049,N_19836);
xnor U25052 (N_25052,N_23227,N_20844);
xor U25053 (N_25053,N_21972,N_19704);
nor U25054 (N_25054,N_18940,N_20027);
or U25055 (N_25055,N_18369,N_23356);
and U25056 (N_25056,N_22921,N_22147);
xor U25057 (N_25057,N_23639,N_23436);
xor U25058 (N_25058,N_19447,N_21697);
nor U25059 (N_25059,N_23491,N_23547);
nor U25060 (N_25060,N_19777,N_23906);
nand U25061 (N_25061,N_19301,N_23262);
nor U25062 (N_25062,N_21311,N_22636);
xor U25063 (N_25063,N_21703,N_18262);
xnor U25064 (N_25064,N_19452,N_23031);
nand U25065 (N_25065,N_19049,N_20019);
nand U25066 (N_25066,N_18643,N_20944);
xor U25067 (N_25067,N_18682,N_21868);
xnor U25068 (N_25068,N_18086,N_21458);
and U25069 (N_25069,N_19460,N_22504);
nor U25070 (N_25070,N_19055,N_19517);
nor U25071 (N_25071,N_21859,N_19736);
or U25072 (N_25072,N_18203,N_22717);
and U25073 (N_25073,N_21614,N_19396);
and U25074 (N_25074,N_20500,N_20658);
and U25075 (N_25075,N_23072,N_20771);
and U25076 (N_25076,N_20670,N_22983);
or U25077 (N_25077,N_19716,N_20814);
nor U25078 (N_25078,N_21409,N_18821);
nor U25079 (N_25079,N_23350,N_21455);
xnor U25080 (N_25080,N_21835,N_18829);
or U25081 (N_25081,N_18182,N_20319);
and U25082 (N_25082,N_19308,N_23026);
xor U25083 (N_25083,N_21351,N_21445);
xnor U25084 (N_25084,N_21065,N_18646);
nand U25085 (N_25085,N_18775,N_18018);
nor U25086 (N_25086,N_22125,N_18999);
nor U25087 (N_25087,N_20453,N_18652);
nor U25088 (N_25088,N_23349,N_23054);
nor U25089 (N_25089,N_19276,N_23993);
xnor U25090 (N_25090,N_23482,N_23246);
nor U25091 (N_25091,N_22424,N_20339);
and U25092 (N_25092,N_18209,N_22048);
nor U25093 (N_25093,N_23239,N_22324);
nor U25094 (N_25094,N_23976,N_19495);
xor U25095 (N_25095,N_18681,N_21270);
and U25096 (N_25096,N_23758,N_19130);
or U25097 (N_25097,N_18255,N_21709);
nand U25098 (N_25098,N_22102,N_23200);
nor U25099 (N_25099,N_22045,N_19000);
or U25100 (N_25100,N_21213,N_19840);
xnor U25101 (N_25101,N_22661,N_22796);
or U25102 (N_25102,N_18748,N_21662);
nand U25103 (N_25103,N_20303,N_23009);
nor U25104 (N_25104,N_18810,N_22239);
nand U25105 (N_25105,N_21136,N_20187);
nor U25106 (N_25106,N_23228,N_20164);
xnor U25107 (N_25107,N_22671,N_23765);
or U25108 (N_25108,N_22010,N_18187);
nand U25109 (N_25109,N_18225,N_23205);
or U25110 (N_25110,N_20600,N_22663);
xor U25111 (N_25111,N_21476,N_22993);
and U25112 (N_25112,N_18745,N_19959);
nor U25113 (N_25113,N_20387,N_19921);
xor U25114 (N_25114,N_23302,N_19597);
nand U25115 (N_25115,N_20808,N_20763);
xor U25116 (N_25116,N_22748,N_19487);
or U25117 (N_25117,N_19419,N_18349);
and U25118 (N_25118,N_19529,N_22876);
nand U25119 (N_25119,N_20209,N_23382);
nor U25120 (N_25120,N_22006,N_23518);
nor U25121 (N_25121,N_18618,N_18286);
xnor U25122 (N_25122,N_23193,N_23699);
nor U25123 (N_25123,N_21610,N_20216);
nand U25124 (N_25124,N_21457,N_23662);
or U25125 (N_25125,N_23845,N_19762);
nor U25126 (N_25126,N_22873,N_22249);
nand U25127 (N_25127,N_18842,N_20482);
or U25128 (N_25128,N_19184,N_19143);
or U25129 (N_25129,N_23885,N_21836);
nand U25130 (N_25130,N_22431,N_22605);
or U25131 (N_25131,N_23372,N_21887);
or U25132 (N_25132,N_20428,N_20177);
or U25133 (N_25133,N_22541,N_23670);
nor U25134 (N_25134,N_20418,N_23574);
xor U25135 (N_25135,N_22080,N_22022);
and U25136 (N_25136,N_19848,N_22738);
xor U25137 (N_25137,N_22889,N_19907);
nor U25138 (N_25138,N_22442,N_19578);
and U25139 (N_25139,N_23334,N_21383);
nor U25140 (N_25140,N_18088,N_21967);
or U25141 (N_25141,N_20724,N_19070);
and U25142 (N_25142,N_19075,N_23490);
and U25143 (N_25143,N_22818,N_19548);
nand U25144 (N_25144,N_18157,N_22660);
nor U25145 (N_25145,N_20859,N_21894);
nor U25146 (N_25146,N_19479,N_19048);
or U25147 (N_25147,N_19877,N_22907);
or U25148 (N_25148,N_23679,N_21265);
and U25149 (N_25149,N_23946,N_21499);
nand U25150 (N_25150,N_21190,N_19203);
xor U25151 (N_25151,N_23287,N_20295);
nand U25152 (N_25152,N_23711,N_22905);
and U25153 (N_25153,N_22322,N_19337);
and U25154 (N_25154,N_21144,N_20163);
nand U25155 (N_25155,N_21753,N_18913);
xnor U25156 (N_25156,N_19674,N_23266);
or U25157 (N_25157,N_21915,N_19310);
or U25158 (N_25158,N_18785,N_20957);
and U25159 (N_25159,N_23782,N_20464);
nor U25160 (N_25160,N_23386,N_19025);
nor U25161 (N_25161,N_19134,N_22264);
xnor U25162 (N_25162,N_19476,N_23022);
and U25163 (N_25163,N_18557,N_23135);
nor U25164 (N_25164,N_23466,N_19832);
and U25165 (N_25165,N_18300,N_21147);
nand U25166 (N_25166,N_23965,N_18357);
or U25167 (N_25167,N_21909,N_23250);
nand U25168 (N_25168,N_18215,N_18909);
nand U25169 (N_25169,N_18611,N_22171);
or U25170 (N_25170,N_22645,N_22244);
or U25171 (N_25171,N_18776,N_20603);
xor U25172 (N_25172,N_18722,N_19424);
nand U25173 (N_25173,N_20601,N_19807);
or U25174 (N_25174,N_19731,N_21427);
nor U25175 (N_25175,N_23059,N_18790);
nand U25176 (N_25176,N_23673,N_21293);
xnor U25177 (N_25177,N_22705,N_18917);
or U25178 (N_25178,N_19772,N_20402);
nand U25179 (N_25179,N_18485,N_18709);
nand U25180 (N_25180,N_22594,N_18902);
nand U25181 (N_25181,N_20676,N_23649);
nand U25182 (N_25182,N_18098,N_18241);
and U25183 (N_25183,N_19064,N_21741);
and U25184 (N_25184,N_22261,N_19196);
xor U25185 (N_25185,N_22197,N_20133);
or U25186 (N_25186,N_20969,N_21795);
or U25187 (N_25187,N_23795,N_21938);
or U25188 (N_25188,N_21078,N_19560);
and U25189 (N_25189,N_18049,N_21654);
and U25190 (N_25190,N_20474,N_18025);
nor U25191 (N_25191,N_20493,N_22014);
and U25192 (N_25192,N_20764,N_23559);
nor U25193 (N_25193,N_18516,N_21747);
or U25194 (N_25194,N_21423,N_22152);
nand U25195 (N_25195,N_22673,N_20657);
and U25196 (N_25196,N_22847,N_18208);
and U25197 (N_25197,N_23234,N_23628);
and U25198 (N_25198,N_21245,N_22251);
or U25199 (N_25199,N_22123,N_21091);
nand U25200 (N_25200,N_21706,N_19370);
nand U25201 (N_25201,N_19789,N_20501);
or U25202 (N_25202,N_21494,N_22055);
xnor U25203 (N_25203,N_21945,N_19971);
and U25204 (N_25204,N_19179,N_21114);
nand U25205 (N_25205,N_23447,N_18386);
nand U25206 (N_25206,N_23058,N_23780);
xor U25207 (N_25207,N_21163,N_20620);
and U25208 (N_25208,N_19466,N_23424);
or U25209 (N_25209,N_19813,N_23151);
and U25210 (N_25210,N_20760,N_20638);
and U25211 (N_25211,N_18353,N_18476);
xor U25212 (N_25212,N_21663,N_19356);
or U25213 (N_25213,N_19249,N_18678);
nand U25214 (N_25214,N_21127,N_22275);
nor U25215 (N_25215,N_21037,N_22368);
nand U25216 (N_25216,N_19287,N_20678);
and U25217 (N_25217,N_21537,N_18651);
nand U25218 (N_25218,N_20263,N_21333);
nor U25219 (N_25219,N_21523,N_18411);
xnor U25220 (N_25220,N_22729,N_21900);
nor U25221 (N_25221,N_20384,N_21486);
nand U25222 (N_25222,N_19306,N_20487);
or U25223 (N_25223,N_22677,N_23818);
nand U25224 (N_25224,N_19655,N_23207);
or U25225 (N_25225,N_23399,N_20525);
nor U25226 (N_25226,N_19901,N_23110);
xor U25227 (N_25227,N_18047,N_20911);
or U25228 (N_25228,N_20952,N_18179);
nand U25229 (N_25229,N_20383,N_20589);
and U25230 (N_25230,N_19698,N_21773);
or U25231 (N_25231,N_19305,N_23966);
nor U25232 (N_25232,N_22465,N_19023);
xor U25233 (N_25233,N_23311,N_20353);
nor U25234 (N_25234,N_19549,N_19392);
and U25235 (N_25235,N_18630,N_19960);
nand U25236 (N_25236,N_21225,N_20964);
and U25237 (N_25237,N_21309,N_22752);
nor U25238 (N_25238,N_23220,N_22851);
or U25239 (N_25239,N_18836,N_21830);
or U25240 (N_25240,N_20426,N_21973);
xor U25241 (N_25241,N_21039,N_18967);
nand U25242 (N_25242,N_20398,N_18195);
xor U25243 (N_25243,N_20321,N_18962);
or U25244 (N_25244,N_21588,N_20125);
nor U25245 (N_25245,N_22656,N_21484);
nand U25246 (N_25246,N_22044,N_22119);
and U25247 (N_25247,N_23500,N_23066);
xnor U25248 (N_25248,N_21699,N_22696);
and U25249 (N_25249,N_20854,N_22926);
xor U25250 (N_25250,N_19838,N_20594);
or U25251 (N_25251,N_21207,N_22894);
or U25252 (N_25252,N_23073,N_18474);
or U25253 (N_25253,N_20868,N_19399);
nor U25254 (N_25254,N_22948,N_19282);
nand U25255 (N_25255,N_23541,N_18339);
and U25256 (N_25256,N_21728,N_23612);
nand U25257 (N_25257,N_22939,N_20430);
nor U25258 (N_25258,N_22181,N_20357);
nor U25259 (N_25259,N_20354,N_23576);
nand U25260 (N_25260,N_20540,N_18238);
and U25261 (N_25261,N_22134,N_21648);
nand U25262 (N_25262,N_23168,N_21771);
nand U25263 (N_25263,N_18197,N_18297);
and U25264 (N_25264,N_22116,N_18803);
or U25265 (N_25265,N_21504,N_18717);
or U25266 (N_25266,N_20330,N_18458);
or U25267 (N_25267,N_22596,N_22448);
or U25268 (N_25268,N_23488,N_20630);
or U25269 (N_25269,N_19861,N_22032);
xor U25270 (N_25270,N_20316,N_19553);
or U25271 (N_25271,N_23282,N_21644);
nand U25272 (N_25272,N_20003,N_22154);
xor U25273 (N_25273,N_19534,N_22670);
nor U25274 (N_25274,N_21819,N_23616);
and U25275 (N_25275,N_22731,N_23275);
nand U25276 (N_25276,N_18185,N_19204);
xor U25277 (N_25277,N_21392,N_19894);
xor U25278 (N_25278,N_19683,N_20604);
nand U25279 (N_25279,N_21028,N_20815);
or U25280 (N_25280,N_19598,N_18841);
xnor U25281 (N_25281,N_18220,N_18014);
nand U25282 (N_25282,N_19825,N_23249);
xnor U25283 (N_25283,N_21763,N_22644);
or U25284 (N_25284,N_21452,N_19475);
nand U25285 (N_25285,N_20656,N_21978);
or U25286 (N_25286,N_19665,N_23817);
or U25287 (N_25287,N_20239,N_21187);
and U25288 (N_25288,N_20653,N_20083);
or U25289 (N_25289,N_18889,N_18625);
and U25290 (N_25290,N_20686,N_18606);
or U25291 (N_25291,N_22357,N_23837);
or U25292 (N_25292,N_18216,N_22566);
xnor U25293 (N_25293,N_19303,N_23045);
nor U25294 (N_25294,N_19852,N_23351);
xnor U25295 (N_25295,N_23124,N_22163);
and U25296 (N_25296,N_19004,N_19990);
nand U25297 (N_25297,N_20577,N_18223);
nand U25298 (N_25298,N_22801,N_22650);
xor U25299 (N_25299,N_20431,N_19809);
nor U25300 (N_25300,N_18831,N_20105);
nor U25301 (N_25301,N_23367,N_20237);
nand U25302 (N_25302,N_20871,N_22133);
or U25303 (N_25303,N_20810,N_20111);
or U25304 (N_25304,N_22025,N_18954);
or U25305 (N_25305,N_23532,N_23641);
xnor U25306 (N_25306,N_20708,N_21922);
nand U25307 (N_25307,N_21845,N_21512);
nor U25308 (N_25308,N_22150,N_19576);
nor U25309 (N_25309,N_20715,N_19278);
or U25310 (N_25310,N_23361,N_19871);
or U25311 (N_25311,N_20414,N_23265);
and U25312 (N_25312,N_23689,N_20645);
nand U25313 (N_25313,N_18570,N_21154);
or U25314 (N_25314,N_23897,N_21698);
nor U25315 (N_25315,N_18083,N_22064);
xnor U25316 (N_25316,N_22023,N_23644);
nor U25317 (N_25317,N_22305,N_20575);
or U25318 (N_25318,N_23377,N_23499);
xnor U25319 (N_25319,N_22618,N_18107);
nand U25320 (N_25320,N_22598,N_22836);
and U25321 (N_25321,N_23261,N_19152);
nand U25322 (N_25322,N_19173,N_19358);
nor U25323 (N_25323,N_23247,N_22255);
nand U25324 (N_25324,N_18493,N_20852);
and U25325 (N_25325,N_19484,N_23852);
nor U25326 (N_25326,N_21804,N_20253);
or U25327 (N_25327,N_18715,N_22405);
nor U25328 (N_25328,N_19573,N_21472);
xnor U25329 (N_25329,N_22402,N_18284);
nor U25330 (N_25330,N_21088,N_20484);
xnor U25331 (N_25331,N_20085,N_19357);
nand U25332 (N_25332,N_21799,N_22140);
nand U25333 (N_25333,N_20270,N_20672);
nand U25334 (N_25334,N_19327,N_20832);
nor U25335 (N_25335,N_19438,N_22024);
xor U25336 (N_25336,N_19001,N_23118);
xnor U25337 (N_25337,N_18281,N_18519);
xnor U25338 (N_25338,N_22780,N_19323);
and U25339 (N_25339,N_20276,N_23461);
or U25340 (N_25340,N_18702,N_18254);
nand U25341 (N_25341,N_18930,N_22895);
xor U25342 (N_25342,N_20241,N_19102);
or U25343 (N_25343,N_22100,N_21368);
xnor U25344 (N_25344,N_21025,N_20440);
nor U25345 (N_25345,N_18094,N_20736);
or U25346 (N_25346,N_23762,N_23911);
and U25347 (N_25347,N_23035,N_21487);
nand U25348 (N_25348,N_21744,N_18514);
xor U25349 (N_25349,N_23680,N_20230);
or U25350 (N_25350,N_21729,N_23910);
xor U25351 (N_25351,N_19014,N_18521);
nor U25352 (N_25352,N_20870,N_21981);
or U25353 (N_25353,N_22575,N_23925);
nand U25354 (N_25354,N_18441,N_21006);
nand U25355 (N_25355,N_18896,N_20782);
nand U25356 (N_25356,N_23752,N_23651);
nand U25357 (N_25357,N_19065,N_19508);
xor U25358 (N_25358,N_22088,N_22263);
and U25359 (N_25359,N_22310,N_18053);
and U25360 (N_25360,N_20154,N_23329);
xor U25361 (N_25361,N_23171,N_18071);
or U25362 (N_25362,N_20089,N_18991);
nor U25363 (N_25363,N_19478,N_21712);
xnor U25364 (N_25364,N_21659,N_20291);
and U25365 (N_25365,N_21393,N_21824);
xnor U25366 (N_25366,N_18437,N_19231);
nor U25367 (N_25367,N_23635,N_23071);
nor U25368 (N_25368,N_23831,N_19112);
xor U25369 (N_25369,N_21604,N_18720);
nand U25370 (N_25370,N_23577,N_20611);
and U25371 (N_25371,N_19615,N_20120);
nand U25372 (N_25372,N_23751,N_23371);
nand U25373 (N_25373,N_19796,N_20376);
nand U25374 (N_25374,N_18145,N_19695);
and U25375 (N_25375,N_23819,N_18222);
nor U25376 (N_25376,N_22523,N_23136);
and U25377 (N_25377,N_23884,N_22204);
xnor U25378 (N_25378,N_18007,N_22510);
xnor U25379 (N_25379,N_18941,N_20113);
or U25380 (N_25380,N_23080,N_22438);
or U25381 (N_25381,N_22869,N_19644);
or U25382 (N_25382,N_19652,N_22609);
nor U25383 (N_25383,N_22515,N_22687);
nor U25384 (N_25384,N_23458,N_21151);
or U25385 (N_25385,N_21630,N_18654);
xnor U25386 (N_25386,N_20726,N_18833);
nand U25387 (N_25387,N_21496,N_19544);
nand U25388 (N_25388,N_20864,N_18928);
and U25389 (N_25389,N_21157,N_19120);
xor U25390 (N_25390,N_23433,N_18240);
nand U25391 (N_25391,N_23944,N_22226);
nand U25392 (N_25392,N_20461,N_18735);
and U25393 (N_25393,N_22491,N_21139);
nor U25394 (N_25394,N_21237,N_19140);
and U25395 (N_25395,N_19682,N_23195);
and U25396 (N_25396,N_22774,N_20923);
or U25397 (N_25397,N_21563,N_21983);
nand U25398 (N_25398,N_20966,N_20206);
and U25399 (N_25399,N_23420,N_20689);
or U25400 (N_25400,N_18553,N_19421);
and U25401 (N_25401,N_22487,N_18461);
and U25402 (N_25402,N_23083,N_18096);
nor U25403 (N_25403,N_20684,N_22842);
and U25404 (N_25404,N_22579,N_21195);
nand U25405 (N_25405,N_20483,N_18998);
nand U25406 (N_25406,N_19268,N_18635);
or U25407 (N_25407,N_19808,N_19841);
or U25408 (N_25408,N_18160,N_21841);
xnor U25409 (N_25409,N_21928,N_18003);
xnor U25410 (N_25410,N_22762,N_20256);
or U25411 (N_25411,N_18926,N_19806);
xnor U25412 (N_25412,N_21310,N_18401);
or U25413 (N_25413,N_19627,N_21120);
and U25414 (N_25414,N_19853,N_22060);
nand U25415 (N_25415,N_20086,N_21534);
or U25416 (N_25416,N_22589,N_18371);
and U25417 (N_25417,N_20066,N_18385);
nand U25418 (N_25418,N_20306,N_18468);
nand U25419 (N_25419,N_22371,N_19745);
nor U25420 (N_25420,N_23599,N_22788);
nor U25421 (N_25421,N_20035,N_22732);
and U25422 (N_25422,N_23725,N_20779);
xor U25423 (N_25423,N_19325,N_18956);
nand U25424 (N_25424,N_20545,N_21768);
xnor U25425 (N_25425,N_21161,N_22708);
or U25426 (N_25426,N_19882,N_23729);
and U25427 (N_25427,N_20885,N_19532);
or U25428 (N_25428,N_23672,N_21577);
nand U25429 (N_25429,N_21518,N_22614);
nor U25430 (N_25430,N_20036,N_23211);
or U25431 (N_25431,N_22955,N_18738);
and U25432 (N_25432,N_20079,N_23719);
nand U25433 (N_25433,N_23984,N_23019);
nand U25434 (N_25434,N_23568,N_23553);
nand U25435 (N_25435,N_20323,N_18055);
and U25436 (N_25436,N_21329,N_18017);
or U25437 (N_25437,N_22202,N_23148);
and U25438 (N_25438,N_21803,N_21613);
nand U25439 (N_25439,N_22052,N_22164);
and U25440 (N_25440,N_19546,N_22518);
nor U25441 (N_25441,N_18447,N_18989);
xnor U25442 (N_25442,N_19828,N_20943);
and U25443 (N_25443,N_22194,N_22860);
xnor U25444 (N_25444,N_23932,N_21379);
xnor U25445 (N_25445,N_18293,N_20765);
and U25446 (N_25446,N_19685,N_23591);
or U25447 (N_25447,N_20933,N_20400);
or U25448 (N_25448,N_19372,N_22083);
xnor U25449 (N_25449,N_20173,N_21759);
nor U25450 (N_25450,N_18052,N_19422);
and U25451 (N_25451,N_23237,N_18846);
xor U25452 (N_25452,N_21084,N_21249);
and U25453 (N_25453,N_22273,N_19381);
xor U25454 (N_25454,N_21717,N_19092);
nand U25455 (N_25455,N_20336,N_18543);
nand U25456 (N_25456,N_19505,N_19865);
nor U25457 (N_25457,N_18959,N_20697);
nor U25458 (N_25458,N_19451,N_23938);
nor U25459 (N_25459,N_22245,N_19386);
or U25460 (N_25460,N_21777,N_21143);
nor U25461 (N_25461,N_20573,N_23431);
nand U25462 (N_25462,N_19539,N_21403);
xor U25463 (N_25463,N_21995,N_23048);
xnor U25464 (N_25464,N_21014,N_23690);
or U25465 (N_25465,N_22190,N_23138);
xnor U25466 (N_25466,N_21371,N_21018);
nand U25467 (N_25467,N_23248,N_18971);
nand U25468 (N_25468,N_23264,N_23055);
or U25469 (N_25469,N_21867,N_22781);
nor U25470 (N_25470,N_23653,N_22272);
and U25471 (N_25471,N_22248,N_19462);
nor U25472 (N_25472,N_19200,N_20786);
and U25473 (N_25473,N_20001,N_18189);
nand U25474 (N_25474,N_20617,N_20702);
nor U25475 (N_25475,N_19253,N_23209);
and U25476 (N_25476,N_21877,N_19494);
and U25477 (N_25477,N_22069,N_23158);
or U25478 (N_25478,N_22018,N_20998);
xor U25479 (N_25479,N_20521,N_18908);
nor U25480 (N_25480,N_20320,N_18144);
and U25481 (N_25481,N_19701,N_20750);
or U25482 (N_25482,N_23359,N_18245);
and U25483 (N_25483,N_18680,N_20328);
and U25484 (N_25484,N_21173,N_20580);
and U25485 (N_25485,N_22927,N_20341);
nor U25486 (N_25486,N_22600,N_22173);
nor U25487 (N_25487,N_22511,N_19769);
nand U25488 (N_25488,N_23970,N_22207);
xnor U25489 (N_25489,N_22635,N_20472);
and U25490 (N_25490,N_23422,N_20646);
and U25491 (N_25491,N_23106,N_23132);
nor U25492 (N_25492,N_22681,N_20563);
nor U25493 (N_25493,N_23043,N_23327);
xor U25494 (N_25494,N_18559,N_18939);
or U25495 (N_25495,N_21784,N_23161);
nor U25496 (N_25496,N_20655,N_21171);
and U25497 (N_25497,N_21955,N_21019);
nor U25498 (N_25498,N_19234,N_20477);
xor U25499 (N_25499,N_18671,N_21618);
nand U25500 (N_25500,N_23867,N_23416);
nand U25501 (N_25501,N_21639,N_21668);
or U25502 (N_25502,N_21998,N_18333);
nor U25503 (N_25503,N_21616,N_21129);
xnor U25504 (N_25504,N_18696,N_23098);
nor U25505 (N_25505,N_19163,N_19426);
xor U25506 (N_25506,N_21052,N_19318);
xor U25507 (N_25507,N_23878,N_22800);
xor U25508 (N_25508,N_23640,N_21035);
or U25509 (N_25509,N_19540,N_21488);
or U25510 (N_25510,N_21554,N_22482);
or U25511 (N_25511,N_23308,N_22151);
xor U25512 (N_25512,N_19523,N_18648);
nor U25513 (N_25513,N_18418,N_22770);
and U25514 (N_25514,N_22985,N_22089);
xor U25515 (N_25515,N_21466,N_19136);
nand U25516 (N_25516,N_21060,N_20401);
xor U25517 (N_25517,N_21647,N_22136);
or U25518 (N_25518,N_19106,N_22056);
nor U25519 (N_25519,N_22078,N_19928);
or U25520 (N_25520,N_23809,N_21992);
nand U25521 (N_25521,N_18213,N_20514);
nor U25522 (N_25522,N_19551,N_22271);
or U25523 (N_25523,N_23027,N_20274);
xnor U25524 (N_25524,N_19721,N_22400);
nand U25525 (N_25525,N_18825,N_23642);
nor U25526 (N_25526,N_21274,N_22761);
and U25527 (N_25527,N_23833,N_22323);
or U25528 (N_25528,N_20081,N_20091);
xor U25529 (N_25529,N_20374,N_23963);
or U25530 (N_25530,N_19463,N_23421);
or U25531 (N_25531,N_22404,N_18045);
nand U25532 (N_25532,N_18523,N_22223);
and U25533 (N_25533,N_21059,N_19913);
nand U25534 (N_25534,N_19897,N_22166);
nor U25535 (N_25535,N_19510,N_19371);
or U25536 (N_25536,N_21798,N_19042);
nor U25537 (N_25537,N_21433,N_21815);
nor U25538 (N_25538,N_21440,N_19724);
nor U25539 (N_25539,N_18755,N_19201);
nand U25540 (N_25540,N_21702,N_22590);
or U25541 (N_25541,N_23481,N_21866);
or U25542 (N_25542,N_21669,N_23537);
or U25543 (N_25543,N_21586,N_22291);
and U25544 (N_25544,N_23113,N_20381);
nand U25545 (N_25545,N_22211,N_23625);
nor U25546 (N_25546,N_19626,N_23933);
nand U25547 (N_25547,N_18368,N_19639);
or U25548 (N_25548,N_21033,N_18336);
or U25549 (N_25549,N_23709,N_22954);
nor U25550 (N_25550,N_21103,N_20273);
xnor U25551 (N_25551,N_23856,N_18450);
nand U25552 (N_25552,N_18642,N_20312);
nor U25553 (N_25553,N_22274,N_19345);
nand U25554 (N_25554,N_19870,N_21684);
and U25555 (N_25555,N_23410,N_18914);
nor U25556 (N_25556,N_19930,N_20041);
and U25557 (N_25557,N_20279,N_19538);
nor U25558 (N_25558,N_18112,N_21917);
nand U25559 (N_25559,N_21183,N_23020);
or U25560 (N_25560,N_18724,N_22587);
xor U25561 (N_25561,N_18384,N_22502);
nand U25562 (N_25562,N_19727,N_23229);
nand U25563 (N_25563,N_22416,N_23023);
xor U25564 (N_25564,N_22200,N_20811);
nand U25565 (N_25565,N_18582,N_22804);
or U25566 (N_25566,N_20075,N_22973);
nand U25567 (N_25567,N_19430,N_22568);
and U25568 (N_25568,N_19622,N_18395);
nand U25569 (N_25569,N_22749,N_19770);
xor U25570 (N_25570,N_21424,N_19229);
nand U25571 (N_25571,N_22266,N_21811);
nor U25572 (N_25572,N_18150,N_19656);
xnor U25573 (N_25573,N_21353,N_22707);
nand U25574 (N_25574,N_21414,N_22040);
xor U25575 (N_25575,N_22972,N_18888);
and U25576 (N_25576,N_21111,N_23441);
nor U25577 (N_25577,N_21774,N_23597);
xor U25578 (N_25578,N_23621,N_19775);
xnor U25579 (N_25579,N_21869,N_18565);
xor U25580 (N_25580,N_23435,N_20057);
xnor U25581 (N_25581,N_19470,N_20557);
and U25582 (N_25582,N_20442,N_20641);
nand U25583 (N_25583,N_20342,N_21040);
nand U25584 (N_25584,N_19178,N_22461);
and U25585 (N_25585,N_23342,N_18597);
and U25586 (N_25586,N_23971,N_18270);
nor U25587 (N_25587,N_21490,N_18064);
and U25588 (N_25588,N_20023,N_19909);
or U25589 (N_25589,N_22278,N_21896);
xor U25590 (N_25590,N_20325,N_22698);
xnor U25591 (N_25591,N_22980,N_19817);
nand U25592 (N_25592,N_23603,N_18275);
or U25593 (N_25593,N_21960,N_21901);
nor U25594 (N_25594,N_20901,N_18348);
xnor U25595 (N_25595,N_23730,N_18292);
xor U25596 (N_25596,N_21556,N_19013);
and U25597 (N_25597,N_21046,N_23196);
nand U25598 (N_25598,N_22168,N_19251);
xor U25599 (N_25599,N_18918,N_19397);
xnor U25600 (N_25600,N_21652,N_23074);
or U25601 (N_25601,N_22935,N_23873);
or U25602 (N_25602,N_20634,N_18232);
xnor U25603 (N_25603,N_22766,N_23369);
and U25604 (N_25604,N_19334,N_20309);
or U25605 (N_25605,N_18501,N_20928);
xor U25606 (N_25606,N_20049,N_23638);
nand U25607 (N_25607,N_20956,N_20626);
nand U25608 (N_25608,N_19542,N_19944);
and U25609 (N_25609,N_21381,N_23197);
nand U25610 (N_25610,N_22547,N_22522);
nand U25611 (N_25611,N_18290,N_18995);
and U25612 (N_25612,N_22514,N_22621);
nand U25613 (N_25613,N_22467,N_22524);
nor U25614 (N_25614,N_23739,N_18425);
xnor U25615 (N_25615,N_23492,N_18573);
nand U25616 (N_25616,N_20375,N_23586);
nor U25617 (N_25617,N_21579,N_20961);
nor U25618 (N_25618,N_19228,N_21256);
nor U25619 (N_25619,N_20255,N_20243);
nor U25620 (N_25620,N_20754,N_21330);
or U25621 (N_25621,N_18061,N_22637);
or U25622 (N_25622,N_22033,N_18622);
nor U25623 (N_25623,N_23659,N_18355);
nor U25624 (N_25624,N_23176,N_20568);
or U25625 (N_25625,N_21991,N_19855);
or U25626 (N_25626,N_22976,N_22718);
and U25627 (N_25627,N_18228,N_18657);
or U25628 (N_25628,N_19246,N_22962);
xor U25629 (N_25629,N_22035,N_18030);
xnor U25630 (N_25630,N_18477,N_22008);
xor U25631 (N_25631,N_19449,N_23380);
nand U25632 (N_25632,N_23857,N_22046);
nor U25633 (N_25633,N_21704,N_22743);
and U25634 (N_25634,N_19603,N_23918);
nor U25635 (N_25635,N_19193,N_21635);
xnor U25636 (N_25636,N_18455,N_20980);
xor U25637 (N_25637,N_21315,N_22777);
nand U25638 (N_25638,N_21921,N_21219);
xnor U25639 (N_25639,N_23179,N_20410);
or U25640 (N_25640,N_21042,N_23538);
nor U25641 (N_25641,N_20404,N_19439);
xnor U25642 (N_25642,N_18758,N_19925);
or U25643 (N_25643,N_19135,N_22028);
nand U25644 (N_25644,N_18184,N_22433);
nand U25645 (N_25645,N_20936,N_19149);
xor U25646 (N_25646,N_20028,N_19866);
nand U25647 (N_25647,N_19876,N_19183);
nor U25648 (N_25648,N_18121,N_23964);
xor U25649 (N_25649,N_23253,N_19605);
and U25650 (N_25650,N_21048,N_18085);
xor U25651 (N_25651,N_21460,N_20612);
nand U25652 (N_25652,N_21631,N_20850);
or U25653 (N_25653,N_21243,N_21337);
nand U25654 (N_25654,N_19497,N_20872);
xor U25655 (N_25655,N_21856,N_19365);
nor U25656 (N_25656,N_19107,N_23277);
nor U25657 (N_25657,N_19688,N_19672);
xnor U25658 (N_25658,N_18513,N_20863);
nand U25659 (N_25659,N_20457,N_22787);
nor U25660 (N_25660,N_20496,N_18087);
or U25661 (N_25661,N_20103,N_22988);
and U25662 (N_25662,N_18921,N_19963);
and U25663 (N_25663,N_21349,N_21679);
xor U25664 (N_25664,N_18004,N_18571);
nand U25665 (N_25665,N_19154,N_18965);
xnor U25666 (N_25666,N_22087,N_18099);
nor U25667 (N_25667,N_22952,N_20995);
or U25668 (N_25668,N_23267,N_22212);
or U25669 (N_25669,N_18563,N_23902);
nand U25670 (N_25670,N_18695,N_21044);
nand U25671 (N_25671,N_19415,N_19956);
nand U25672 (N_25672,N_18595,N_19616);
and U25673 (N_25673,N_23459,N_23215);
xor U25674 (N_25674,N_22690,N_19063);
xnor U25675 (N_25675,N_19101,N_20031);
nand U25676 (N_25676,N_18539,N_21871);
nand U25677 (N_25677,N_20520,N_19458);
and U25678 (N_25678,N_23802,N_18857);
or U25679 (N_25679,N_20361,N_23624);
xnor U25680 (N_25680,N_23724,N_22613);
or U25681 (N_25681,N_18700,N_20920);
or U25682 (N_25682,N_22797,N_22111);
and U25683 (N_25683,N_19651,N_19197);
nand U25684 (N_25684,N_23028,N_18761);
xor U25685 (N_25685,N_19393,N_23075);
and U25686 (N_25686,N_20134,N_18268);
nor U25687 (N_25687,N_20310,N_22250);
and U25688 (N_25688,N_18486,N_20555);
nand U25689 (N_25689,N_20240,N_21134);
nand U25690 (N_25690,N_20475,N_19459);
nor U25691 (N_25691,N_20463,N_22821);
and U25692 (N_25692,N_18302,N_19667);
nand U25693 (N_25693,N_22813,N_19563);
nor U25694 (N_25694,N_22874,N_22105);
or U25695 (N_25695,N_23214,N_23395);
and U25696 (N_25696,N_23924,N_22978);
nand U25697 (N_25697,N_21913,N_22875);
xnor U25698 (N_25698,N_19205,N_19570);
and U25699 (N_25699,N_23452,N_22384);
xnor U25700 (N_25700,N_19176,N_22020);
and U25701 (N_25701,N_18444,N_19148);
xor U25702 (N_25702,N_20907,N_19464);
or U25703 (N_25703,N_19583,N_21643);
xnor U25704 (N_25704,N_21277,N_20640);
xor U25705 (N_25705,N_19269,N_23115);
or U25706 (N_25706,N_18020,N_23595);
and U25707 (N_25707,N_18948,N_19259);
xnor U25708 (N_25708,N_23160,N_22298);
and U25709 (N_25709,N_18728,N_21727);
and U25710 (N_25710,N_20881,N_20812);
xnor U25711 (N_25711,N_21012,N_23468);
nand U25712 (N_25712,N_21757,N_20112);
nor U25713 (N_25713,N_18141,N_21904);
xor U25714 (N_25714,N_20124,N_20199);
nand U25715 (N_25715,N_22169,N_22479);
nand U25716 (N_25716,N_22838,N_21628);
nand U25717 (N_25717,N_23155,N_20926);
nor U25718 (N_25718,N_18862,N_20492);
and U25719 (N_25719,N_21705,N_19455);
and U25720 (N_25720,N_18005,N_20537);
xor U25721 (N_25721,N_22093,N_23740);
nor U25722 (N_25722,N_23619,N_18665);
or U25723 (N_25723,N_18524,N_20706);
and U25724 (N_25724,N_22214,N_18679);
xnor U25725 (N_25725,N_19445,N_21544);
nand U25726 (N_25726,N_23189,N_22346);
nor U25727 (N_25727,N_23414,N_20999);
and U25728 (N_25728,N_23412,N_20371);
or U25729 (N_25729,N_21205,N_22176);
xor U25730 (N_25730,N_23692,N_20523);
xnor U25731 (N_25731,N_18602,N_19007);
nand U25732 (N_25732,N_22888,N_18577);
xnor U25733 (N_25733,N_21843,N_19312);
nor U25734 (N_25734,N_20218,N_23510);
xnor U25735 (N_25735,N_20436,N_21404);
or U25736 (N_25736,N_20443,N_19095);
nor U25737 (N_25737,N_21839,N_21951);
nand U25738 (N_25738,N_20699,N_20725);
nand U25739 (N_25739,N_20300,N_20741);
nand U25740 (N_25740,N_19277,N_23340);
xor U25741 (N_25741,N_19580,N_22135);
or U25742 (N_25742,N_20513,N_18584);
xor U25743 (N_25743,N_20033,N_20215);
and U25744 (N_25744,N_19604,N_21118);
xnor U25745 (N_25745,N_19804,N_22462);
nand U25746 (N_25746,N_22806,N_18324);
nand U25747 (N_25747,N_19244,N_18040);
or U25748 (N_25748,N_23292,N_21788);
nand U25749 (N_25749,N_19218,N_23335);
nor U25750 (N_25750,N_20692,N_19521);
nor U25751 (N_25751,N_19935,N_23594);
xor U25752 (N_25752,N_21672,N_18592);
or U25753 (N_25753,N_23683,N_18969);
xor U25754 (N_25754,N_20768,N_22289);
and U25755 (N_25755,N_23060,N_23232);
or U25756 (N_25756,N_19115,N_19793);
nand U25757 (N_25757,N_19752,N_19878);
nand U25758 (N_25758,N_21580,N_22848);
or U25759 (N_25759,N_19668,N_19518);
and U25760 (N_25760,N_22084,N_22427);
nor U25761 (N_25761,N_19256,N_20681);
or U25762 (N_25762,N_22068,N_23094);
or U25763 (N_25763,N_19209,N_18279);
nand U25764 (N_25764,N_19873,N_19021);
and U25765 (N_25765,N_18095,N_18945);
and U25766 (N_25766,N_23162,N_20533);
xor U25767 (N_25767,N_22299,N_23501);
nand U25768 (N_25768,N_21919,N_19503);
nor U25769 (N_25769,N_22121,N_23620);
nor U25770 (N_25770,N_19113,N_20503);
and U25771 (N_25771,N_21710,N_22653);
and U25772 (N_25772,N_21650,N_22809);
nor U25773 (N_25773,N_19599,N_20562);
xor U25774 (N_25774,N_22213,N_18719);
and U25775 (N_25775,N_18615,N_19187);
nor U25776 (N_25776,N_19059,N_18488);
nor U25777 (N_25777,N_21926,N_22936);
and U25778 (N_25778,N_22132,N_20593);
nand U25779 (N_25779,N_20949,N_22096);
nand U25780 (N_25780,N_22129,N_18027);
nand U25781 (N_25781,N_19352,N_22714);
or U25782 (N_25782,N_22339,N_19854);
and U25783 (N_25783,N_22440,N_21829);
nand U25784 (N_25784,N_20743,N_22157);
nor U25785 (N_25785,N_21317,N_21790);
xnor U25786 (N_25786,N_22833,N_18137);
or U25787 (N_25787,N_22987,N_18306);
or U25788 (N_25788,N_18799,N_19473);
xnor U25789 (N_25789,N_23307,N_21953);
xnor U25790 (N_25790,N_23886,N_22340);
and U25791 (N_25791,N_20393,N_19350);
or U25792 (N_25792,N_18764,N_19072);
nand U25793 (N_25793,N_20766,N_20379);
xor U25794 (N_25794,N_23111,N_21156);
or U25795 (N_25795,N_19017,N_20038);
nor U25796 (N_25796,N_20805,N_20696);
and U25797 (N_25797,N_23016,N_20259);
or U25798 (N_25798,N_23694,N_19945);
xor U25799 (N_25799,N_19376,N_18647);
nor U25800 (N_25800,N_19098,N_22419);
and U25801 (N_25801,N_20021,N_22710);
xnor U25802 (N_25802,N_20835,N_21932);
and U25803 (N_25803,N_22911,N_18498);
xnor U25804 (N_25804,N_23827,N_20064);
or U25805 (N_25805,N_18376,N_21767);
and U25806 (N_25806,N_23469,N_23014);
nor U25807 (N_25807,N_21343,N_21857);
and U25808 (N_25808,N_22374,N_23125);
or U25809 (N_25809,N_19713,N_22783);
nor U25810 (N_25810,N_19915,N_23117);
and U25811 (N_25811,N_21390,N_22472);
and U25812 (N_25812,N_20729,N_18992);
xor U25813 (N_25813,N_22571,N_23561);
xnor U25814 (N_25814,N_20637,N_23914);
xor U25815 (N_25815,N_22241,N_23067);
or U25816 (N_25816,N_23358,N_21667);
and U25817 (N_25817,N_19448,N_19005);
nor U25818 (N_25818,N_19020,N_19533);
nor U25819 (N_25819,N_20171,N_22499);
xor U25820 (N_25820,N_20598,N_18424);
xor U25821 (N_25821,N_20566,N_20355);
or U25822 (N_25822,N_18683,N_20848);
nand U25823 (N_25823,N_20417,N_18115);
nor U25824 (N_25824,N_20090,N_21335);
and U25825 (N_25825,N_20698,N_19441);
or U25826 (N_25826,N_21559,N_18081);
nor U25827 (N_25827,N_23157,N_19401);
or U25828 (N_25828,N_23607,N_20272);
xnor U25829 (N_25829,N_23143,N_21660);
and U25830 (N_25830,N_21564,N_22995);
nand U25831 (N_25831,N_18283,N_22716);
nor U25832 (N_25832,N_19985,N_18581);
nand U25833 (N_25833,N_22460,N_23123);
nor U25834 (N_25834,N_21550,N_22880);
or U25835 (N_25835,N_21502,N_23517);
or U25836 (N_25836,N_18409,N_20391);
and U25837 (N_25837,N_21261,N_19630);
nor U25838 (N_25838,N_23439,N_23868);
and U25839 (N_25839,N_18876,N_22606);
xnor U25840 (N_25840,N_23900,N_23240);
or U25841 (N_25841,N_19056,N_23702);
nor U25842 (N_25842,N_18848,N_21071);
nor U25843 (N_25843,N_20197,N_22779);
nand U25844 (N_25844,N_21047,N_19932);
xor U25845 (N_25845,N_19864,N_22525);
nand U25846 (N_25846,N_22423,N_21929);
nand U25847 (N_25847,N_18634,N_23535);
nand U25848 (N_25848,N_22331,N_23613);
nand U25849 (N_25849,N_23637,N_23178);
nand U25850 (N_25850,N_23315,N_23434);
and U25851 (N_25851,N_19481,N_20799);
nand U25852 (N_25852,N_20286,N_21081);
nor U25853 (N_25853,N_23894,N_19297);
nor U25854 (N_25854,N_23344,N_19896);
xnor U25855 (N_25855,N_18549,N_20314);
xor U25856 (N_25856,N_22883,N_20188);
and U25857 (N_25857,N_20258,N_20389);
nand U25858 (N_25858,N_20408,N_20889);
nor U25859 (N_25859,N_21131,N_20116);
or U25860 (N_25860,N_21916,N_19527);
and U25861 (N_25861,N_18408,N_18383);
xor U25862 (N_25862,N_20769,N_23539);
or U25863 (N_25863,N_18311,N_18868);
xnor U25864 (N_25864,N_23912,N_20801);
xor U25865 (N_25865,N_21051,N_23167);
nand U25866 (N_25866,N_19145,N_23270);
xor U25867 (N_25867,N_22931,N_19740);
or U25868 (N_25868,N_22979,N_23355);
or U25869 (N_25869,N_21528,N_23756);
xor U25870 (N_25870,N_19681,N_19782);
and U25871 (N_25871,N_23030,N_21500);
nor U25872 (N_25872,N_21687,N_22201);
and U25873 (N_25873,N_18832,N_20437);
nand U25874 (N_25874,N_21793,N_18138);
nor U25875 (N_25875,N_23238,N_20879);
and U25876 (N_25876,N_20642,N_20200);
or U25877 (N_25877,N_18797,N_20070);
nand U25878 (N_25878,N_21473,N_19912);
and U25879 (N_25879,N_21067,N_20345);
nand U25880 (N_25880,N_19849,N_20153);
and U25881 (N_25881,N_23931,N_22967);
nor U25882 (N_25882,N_20784,N_19003);
nand U25883 (N_25883,N_18289,N_18272);
nand U25884 (N_25884,N_18206,N_23271);
nor U25885 (N_25885,N_19078,N_19640);
nand U25886 (N_25886,N_21444,N_20204);
and U25887 (N_25887,N_20959,N_23314);
or U25888 (N_25888,N_22971,N_22178);
or U25889 (N_25889,N_21792,N_22535);
nand U25890 (N_25890,N_19887,N_21517);
xnor U25891 (N_25891,N_19068,N_22036);
and U25892 (N_25892,N_21769,N_18812);
and U25893 (N_25893,N_22314,N_21102);
nand U25894 (N_25894,N_19708,N_20405);
nand U25895 (N_25895,N_21227,N_20534);
and U25896 (N_25896,N_20649,N_18878);
xnor U25897 (N_25897,N_20249,N_23826);
and U25898 (N_25898,N_23346,N_22292);
nand U25899 (N_25899,N_22815,N_18895);
or U25900 (N_25900,N_19888,N_18804);
or U25901 (N_25901,N_21438,N_19585);
and U25902 (N_25902,N_20560,N_23102);
xor U25903 (N_25903,N_18235,N_23419);
and U25904 (N_25904,N_21160,N_22382);
nand U25905 (N_25905,N_22293,N_22776);
or U25906 (N_25906,N_20690,N_20667);
or U25907 (N_25907,N_22072,N_21807);
or U25908 (N_25908,N_21910,N_22051);
xnor U25909 (N_25909,N_20368,N_23551);
or U25910 (N_25910,N_18802,N_19241);
or U25911 (N_25911,N_18885,N_20317);
nand U25912 (N_25912,N_18307,N_23387);
nor U25913 (N_25913,N_19227,N_21905);
nand U25914 (N_25914,N_23584,N_23283);
or U25915 (N_25915,N_21387,N_18451);
nand U25916 (N_25916,N_21761,N_21510);
nor U25917 (N_25917,N_19642,N_23728);
xor U25918 (N_25918,N_18382,N_20454);
or U25919 (N_25919,N_23310,N_18139);
nor U25920 (N_25920,N_22558,N_19002);
xnor U25921 (N_25921,N_21572,N_18352);
or U25922 (N_25922,N_18073,N_20792);
nand U25923 (N_25923,N_21285,N_23423);
nand U25924 (N_25924,N_19572,N_22933);
nor U25925 (N_25925,N_18834,N_19783);
nor U25926 (N_25926,N_22683,N_18699);
nand U25927 (N_25927,N_20122,N_18726);
nor U25928 (N_25928,N_20388,N_20542);
nand U25929 (N_25929,N_20691,N_21375);
and U25930 (N_25930,N_21297,N_18587);
xnor U25931 (N_25931,N_23923,N_18320);
nand U25932 (N_25932,N_19240,N_22793);
nand U25933 (N_25933,N_18331,N_18506);
nor U25934 (N_25934,N_22458,N_20985);
xnor U25935 (N_25935,N_19648,N_18435);
and U25936 (N_25936,N_23011,N_19526);
xor U25937 (N_25937,N_21589,N_22584);
or U25938 (N_25938,N_22870,N_21021);
nor U25939 (N_25939,N_18555,N_21389);
and U25940 (N_25940,N_20002,N_21188);
nor U25941 (N_25941,N_21802,N_22406);
xnor U25942 (N_25942,N_18509,N_19953);
and U25943 (N_25943,N_20704,N_20076);
nand U25944 (N_25944,N_22039,N_19215);
xor U25945 (N_25945,N_19181,N_22302);
xnor U25946 (N_25946,N_22449,N_18996);
or U25947 (N_25947,N_20819,N_19749);
and U25948 (N_25948,N_23917,N_19884);
nor U25949 (N_25949,N_18583,N_21475);
or U25950 (N_25950,N_22378,N_20797);
and U25951 (N_25951,N_23877,N_23791);
nand U25952 (N_25952,N_18146,N_21177);
xnor U25953 (N_25953,N_21655,N_18931);
and U25954 (N_25954,N_21124,N_20059);
and U25955 (N_25955,N_21292,N_23153);
and U25956 (N_25956,N_19679,N_20794);
nand U25957 (N_25957,N_22728,N_19330);
nand U25958 (N_25958,N_21069,N_19311);
xnor U25959 (N_25959,N_20367,N_22373);
nand U25960 (N_25960,N_21993,N_18806);
and U25961 (N_25961,N_18258,N_22390);
and U25962 (N_25962,N_18856,N_23254);
and U25963 (N_25963,N_20561,N_19214);
xnor U25964 (N_25964,N_19843,N_23406);
xnor U25965 (N_25965,N_23777,N_22445);
and U25966 (N_25966,N_19530,N_21551);
or U25967 (N_25967,N_21367,N_21186);
nor U25968 (N_25968,N_23146,N_20793);
or U25969 (N_25969,N_23037,N_20141);
xor U25970 (N_25970,N_23655,N_20043);
and U25971 (N_25971,N_22258,N_23353);
or U25972 (N_25972,N_22862,N_22826);
nand U25973 (N_25973,N_20937,N_22599);
or U25974 (N_25974,N_19051,N_19968);
nand U25975 (N_25975,N_18226,N_22308);
and U25976 (N_25976,N_22565,N_19353);
or U25977 (N_25977,N_20829,N_19329);
and U25978 (N_25978,N_18256,N_19225);
or U25979 (N_25979,N_23524,N_18427);
xnor U25980 (N_25980,N_23191,N_21594);
or U25981 (N_25981,N_19671,N_19992);
and U25982 (N_25982,N_19725,N_22886);
and U25983 (N_25983,N_23806,N_20875);
xnor U25984 (N_25984,N_18716,N_21607);
and U25985 (N_25985,N_19541,N_22727);
or U25986 (N_25986,N_23685,N_18979);
or U25987 (N_25987,N_21935,N_20978);
nand U25988 (N_25988,N_19390,N_19554);
nor U25989 (N_25989,N_19079,N_22546);
or U25990 (N_25990,N_23648,N_22437);
nand U25991 (N_25991,N_22017,N_19600);
and U25992 (N_25992,N_19054,N_22835);
nand U25993 (N_25993,N_21801,N_23442);
nor U25994 (N_25994,N_21447,N_22812);
nand U25995 (N_25995,N_21671,N_18840);
nor U25996 (N_25996,N_21413,N_19631);
nor U25997 (N_25997,N_23091,N_20538);
nor U25998 (N_25998,N_18050,N_21600);
xor U25999 (N_25999,N_22041,N_21503);
or U26000 (N_26000,N_18287,N_22756);
or U26001 (N_26001,N_23069,N_20971);
xor U26002 (N_26002,N_19917,N_18721);
and U26003 (N_26003,N_22915,N_18269);
and U26004 (N_26004,N_23183,N_19252);
nand U26005 (N_26005,N_18873,N_23650);
and U26006 (N_26006,N_19965,N_19564);
or U26007 (N_26007,N_19010,N_20207);
xnor U26008 (N_26008,N_19764,N_20365);
and U26009 (N_26009,N_20419,N_21721);
xor U26010 (N_26010,N_19217,N_21751);
nor U26011 (N_26011,N_19982,N_23623);
xnor U26012 (N_26012,N_23471,N_21723);
nor U26013 (N_26013,N_19119,N_18298);
nor U26014 (N_26014,N_19946,N_18415);
xnor U26015 (N_26015,N_21511,N_19516);
nor U26016 (N_26016,N_19084,N_23036);
nor U26017 (N_26017,N_20988,N_19450);
or U26018 (N_26018,N_21974,N_20119);
xor U26019 (N_26019,N_20965,N_19373);
and U26020 (N_26020,N_21713,N_22930);
nand U26021 (N_26021,N_23141,N_23476);
or U26022 (N_26022,N_23397,N_18152);
or U26023 (N_26023,N_20065,N_23769);
and U26024 (N_26024,N_19028,N_19157);
nand U26025 (N_26025,N_20946,N_19230);
xor U26026 (N_26026,N_22464,N_21876);
nor U26027 (N_26027,N_19905,N_19432);
nor U26028 (N_26028,N_23203,N_23942);
nand U26029 (N_26029,N_20447,N_22640);
and U26030 (N_26030,N_23870,N_23606);
nand U26031 (N_26031,N_19759,N_23705);
nand U26032 (N_26032,N_23671,N_18663);
nand U26033 (N_26033,N_22550,N_20990);
nor U26034 (N_26034,N_22205,N_22941);
nand U26035 (N_26035,N_22285,N_23987);
xor U26036 (N_26036,N_19723,N_19496);
and U26037 (N_26037,N_21331,N_19039);
xor U26038 (N_26038,N_22219,N_23017);
nor U26039 (N_26039,N_23563,N_18459);
or U26040 (N_26040,N_21509,N_23959);
nand U26041 (N_26041,N_20194,N_20887);
nand U26042 (N_26042,N_23289,N_20324);
nand U26043 (N_26043,N_20495,N_18143);
xnor U26044 (N_26044,N_22669,N_19493);
or U26045 (N_26045,N_20531,N_23384);
nor U26046 (N_26046,N_18056,N_22578);
xnor U26047 (N_26047,N_19661,N_20238);
and U26048 (N_26048,N_18691,N_21962);
nor U26049 (N_26049,N_18760,N_20730);
nor U26050 (N_26050,N_23044,N_22564);
and U26051 (N_26051,N_21105,N_18585);
xnor U26052 (N_26052,N_21828,N_21095);
xor U26053 (N_26053,N_23415,N_20014);
xor U26054 (N_26054,N_18416,N_23182);
or U26055 (N_26055,N_20018,N_23457);
or U26056 (N_26056,N_22593,N_18090);
and U26057 (N_26057,N_20165,N_18567);
xor U26058 (N_26058,N_22772,N_19409);
nand U26059 (N_26059,N_23668,N_21193);
nand U26060 (N_26060,N_22517,N_19950);
nand U26061 (N_26061,N_22557,N_21526);
and U26062 (N_26062,N_18782,N_20508);
nand U26063 (N_26063,N_18813,N_23555);
and U26064 (N_26064,N_21009,N_18332);
nand U26065 (N_26065,N_21013,N_23373);
nor U26066 (N_26066,N_18167,N_19410);
and U26067 (N_26067,N_21827,N_19588);
or U26068 (N_26068,N_18507,N_21412);
nand U26069 (N_26069,N_19895,N_23062);
and U26070 (N_26070,N_19367,N_21585);
nor U26071 (N_26071,N_21421,N_23374);
nor U26072 (N_26072,N_20629,N_18552);
xnor U26073 (N_26073,N_19602,N_23723);
nand U26074 (N_26074,N_18771,N_22231);
nand U26075 (N_26075,N_23768,N_18364);
and U26076 (N_26076,N_20518,N_18713);
or U26077 (N_26077,N_19403,N_19593);
or U26078 (N_26078,N_21092,N_20479);
and U26079 (N_26079,N_23582,N_20109);
and U26080 (N_26080,N_20074,N_20050);
and U26081 (N_26081,N_21619,N_20882);
nand U26082 (N_26082,N_23290,N_20406);
and U26083 (N_26083,N_22608,N_22370);
nor U26084 (N_26084,N_22306,N_19190);
and U26085 (N_26085,N_19555,N_20392);
or U26086 (N_26086,N_21686,N_20627);
nand U26087 (N_26087,N_22542,N_19239);
or U26088 (N_26088,N_19009,N_23844);
and U26089 (N_26089,N_21732,N_19057);
or U26090 (N_26090,N_21032,N_22473);
or U26091 (N_26091,N_20922,N_19689);
and U26092 (N_26092,N_21222,N_20390);
nor U26093 (N_26093,N_21525,N_20714);
and U26094 (N_26094,N_23360,N_19611);
or U26095 (N_26095,N_21288,N_18366);
xor U26096 (N_26096,N_19610,N_22682);
nand U26097 (N_26097,N_19069,N_22893);
xor U26098 (N_26098,N_23677,N_18561);
and U26099 (N_26099,N_23256,N_18374);
nand U26100 (N_26100,N_19313,N_23811);
or U26101 (N_26101,N_20413,N_22595);
nor U26102 (N_26102,N_20648,N_20350);
nand U26103 (N_26103,N_21418,N_18616);
xor U26104 (N_26104,N_19543,N_23766);
nor U26105 (N_26105,N_19739,N_20842);
and U26106 (N_26106,N_21883,N_21765);
or U26107 (N_26107,N_23960,N_21374);
and U26108 (N_26108,N_20939,N_21465);
xnor U26109 (N_26109,N_21116,N_19127);
nor U26110 (N_26110,N_20820,N_19289);
nor U26111 (N_26111,N_23898,N_23444);
or U26112 (N_26112,N_18264,N_19778);
xnor U26113 (N_26113,N_19335,N_20403);
or U26114 (N_26114,N_21063,N_20289);
xnor U26115 (N_26115,N_19938,N_21539);
nand U26116 (N_26116,N_23198,N_21939);
or U26117 (N_26117,N_21708,N_18973);
or U26118 (N_26118,N_21107,N_18718);
and U26119 (N_26119,N_21478,N_22569);
xor U26120 (N_26120,N_21988,N_19528);
nor U26121 (N_26121,N_20138,N_21931);
or U26122 (N_26122,N_20903,N_19338);
xnor U26123 (N_26123,N_21976,N_23293);
or U26124 (N_26124,N_20581,N_22234);
xor U26125 (N_26125,N_18202,N_20172);
and U26126 (N_26126,N_22047,N_18375);
xor U26127 (N_26127,N_22865,N_22666);
nand U26128 (N_26128,N_18952,N_19766);
nor U26129 (N_26129,N_22112,N_18312);
nand U26130 (N_26130,N_22953,N_21937);
and U26131 (N_26131,N_22582,N_22828);
or U26132 (N_26132,N_23376,N_22311);
xnor U26133 (N_26133,N_19161,N_23284);
nand U26134 (N_26134,N_21724,N_23919);
nand U26135 (N_26135,N_22958,N_18390);
nor U26136 (N_26136,N_20069,N_23300);
xor U26137 (N_26137,N_20360,N_23899);
and U26138 (N_26138,N_20333,N_20548);
nand U26139 (N_26139,N_22042,N_23735);
xor U26140 (N_26140,N_20394,N_18892);
nand U26141 (N_26141,N_19934,N_20459);
nand U26142 (N_26142,N_20308,N_21984);
and U26143 (N_26143,N_21854,N_22489);
and U26144 (N_26144,N_19380,N_21236);
and U26145 (N_26145,N_18532,N_21110);
or U26146 (N_26146,N_18986,N_22104);
or U26147 (N_26147,N_22435,N_19509);
xnor U26148 (N_26148,N_20711,N_19862);
and U26149 (N_26149,N_22695,N_18101);
nand U26150 (N_26150,N_23337,N_22012);
nand U26151 (N_26151,N_20940,N_18134);
xnor U26152 (N_26152,N_21524,N_18943);
xor U26153 (N_26153,N_19443,N_22210);
and U26154 (N_26154,N_22203,N_23440);
and U26155 (N_26155,N_19702,N_19294);
nand U26156 (N_26156,N_18044,N_23529);
nand U26157 (N_26157,N_20721,N_18171);
or U26158 (N_26158,N_20315,N_21322);
and U26159 (N_26159,N_22337,N_21560);
nor U26160 (N_26160,N_21307,N_22074);
nand U26161 (N_26161,N_22657,N_23294);
nand U26162 (N_26162,N_22191,N_20048);
or U26163 (N_26163,N_18242,N_19440);
and U26164 (N_26164,N_22519,N_20511);
nor U26165 (N_26165,N_18591,N_20202);
nand U26166 (N_26166,N_19700,N_19924);
nand U26167 (N_26167,N_21689,N_18118);
and U26168 (N_26168,N_18363,N_23614);
xor U26169 (N_26169,N_19632,N_21562);
or U26170 (N_26170,N_23598,N_23712);
xor U26171 (N_26171,N_23872,N_23173);
nor U26172 (N_26172,N_22186,N_22352);
nand U26173 (N_26173,N_20816,N_20972);
nor U26174 (N_26174,N_23034,N_21316);
nand U26175 (N_26175,N_20774,N_20232);
and U26176 (N_26176,N_23800,N_21640);
nor U26177 (N_26177,N_18869,N_23717);
nor U26178 (N_26178,N_21426,N_18924);
nor U26179 (N_26179,N_19280,N_18032);
nand U26180 (N_26180,N_22000,N_22209);
or U26181 (N_26181,N_21840,N_22580);
or U26182 (N_26182,N_21911,N_20587);
or U26183 (N_26183,N_20668,N_18662);
nand U26184 (N_26184,N_19281,N_22567);
nand U26185 (N_26185,N_22758,N_23530);
nor U26186 (N_26186,N_23079,N_23375);
xnor U26187 (N_26187,N_23814,N_23252);
nor U26188 (N_26188,N_21570,N_21606);
nor U26189 (N_26189,N_20989,N_18433);
and U26190 (N_26190,N_19324,N_21520);
and U26191 (N_26191,N_21083,N_19999);
nor U26192 (N_26192,N_20651,N_20108);
xnor U26193 (N_26193,N_18316,N_22167);
and U26194 (N_26194,N_18024,N_23164);
and U26195 (N_26195,N_23047,N_18389);
and U26196 (N_26196,N_19141,N_23411);
xnor U26197 (N_26197,N_18950,N_19483);
nor U26198 (N_26198,N_18310,N_21016);
nor U26199 (N_26199,N_19212,N_22397);
nor U26200 (N_26200,N_21599,N_23312);
nor U26201 (N_26201,N_19006,N_21716);
nand U26202 (N_26202,N_23552,N_21982);
nor U26203 (N_26203,N_18711,N_23451);
nand U26204 (N_26204,N_18608,N_20150);
or U26205 (N_26205,N_20039,N_22350);
or U26206 (N_26206,N_19803,N_19066);
and U26207 (N_26207,N_18515,N_21961);
nor U26208 (N_26208,N_22196,N_18850);
nor U26209 (N_26209,N_23285,N_18125);
or U26210 (N_26210,N_21778,N_23571);
and U26211 (N_26211,N_22478,N_21312);
and U26212 (N_26212,N_21740,N_20650);
nor U26213 (N_26213,N_20927,N_23815);
nand U26214 (N_26214,N_21956,N_22215);
and U26215 (N_26215,N_22917,N_21255);
nor U26216 (N_26216,N_21461,N_19851);
and U26217 (N_26217,N_22852,N_23989);
and U26218 (N_26218,N_21072,N_21001);
nand U26219 (N_26219,N_22316,N_22563);
nand U26220 (N_26220,N_22626,N_22680);
or U26221 (N_26221,N_18484,N_22724);
nor U26222 (N_26222,N_20344,N_23605);
xnor U26223 (N_26223,N_20795,N_21008);
or U26224 (N_26224,N_19474,N_22737);
xor U26225 (N_26225,N_18022,N_19267);
nand U26226 (N_26226,N_18172,N_22143);
xor U26227 (N_26227,N_19363,N_19012);
nand U26228 (N_26228,N_18859,N_22891);
xor U26229 (N_26229,N_19933,N_23842);
xnor U26230 (N_26230,N_20009,N_19389);
and U26231 (N_26231,N_23850,N_22343);
or U26232 (N_26232,N_21267,N_20660);
nand U26233 (N_26233,N_21339,N_23015);
nor U26234 (N_26234,N_20056,N_23590);
xnor U26235 (N_26235,N_18667,N_21934);
xnor U26236 (N_26236,N_22385,N_18105);
and U26237 (N_26237,N_22379,N_23331);
xor U26238 (N_26238,N_22230,N_18250);
and U26239 (N_26239,N_19408,N_20185);
nor U26240 (N_26240,N_19559,N_21152);
and U26241 (N_26241,N_20307,N_19502);
nor U26242 (N_26242,N_20530,N_23930);
nand U26243 (N_26243,N_18276,N_22586);
or U26244 (N_26244,N_23596,N_18693);
or U26245 (N_26245,N_19375,N_18677);
xnor U26246 (N_26246,N_19235,N_18604);
nand U26247 (N_26247,N_20168,N_19011);
nand U26248 (N_26248,N_18542,N_18354);
and U26249 (N_26249,N_21344,N_18968);
nor U26250 (N_26250,N_18767,N_18170);
nand U26251 (N_26251,N_19719,N_20853);
and U26252 (N_26252,N_18472,N_18392);
or U26253 (N_26253,N_23013,N_23913);
and U26254 (N_26254,N_23039,N_18624);
and U26255 (N_26255,N_22131,N_23928);
and U26256 (N_26256,N_22120,N_21952);
and U26257 (N_26257,N_21575,N_22581);
xor U26258 (N_26258,N_19088,N_19826);
and U26259 (N_26259,N_23787,N_18578);
nor U26260 (N_26260,N_23269,N_22755);
nor U26261 (N_26261,N_19456,N_23684);
and U26262 (N_26262,N_18330,N_20427);
or U26263 (N_26263,N_23427,N_20155);
and U26264 (N_26264,N_22867,N_20088);
or U26265 (N_26265,N_21645,N_20893);
and U26266 (N_26266,N_20326,N_23718);
nand U26267 (N_26267,N_22062,N_19899);
or U26268 (N_26268,N_18614,N_20476);
or U26269 (N_26269,N_20761,N_22845);
nor U26270 (N_26270,N_18236,N_23276);
and U26271 (N_26271,N_18982,N_20017);
xor U26272 (N_26272,N_22095,N_22079);
xnor U26273 (N_26273,N_19733,N_22243);
and U26274 (N_26274,N_18685,N_22678);
nand U26275 (N_26275,N_18807,N_21501);
xor U26276 (N_26276,N_23281,N_21593);
and U26277 (N_26277,N_20732,N_18412);
nand U26278 (N_26278,N_20007,N_22057);
and U26279 (N_26279,N_20894,N_22872);
nand U26280 (N_26280,N_20720,N_21448);
nand U26281 (N_26281,N_21282,N_22532);
and U26282 (N_26282,N_23336,N_20231);
or U26283 (N_26283,N_19557,N_21880);
and U26284 (N_26284,N_19109,N_23306);
nand U26285 (N_26285,N_21252,N_22280);
xor U26286 (N_26286,N_23348,N_19595);
xnor U26287 (N_26287,N_20984,N_18572);
nor U26288 (N_26288,N_23742,N_23839);
nand U26289 (N_26289,N_18987,N_23462);
or U26290 (N_26290,N_18308,N_23697);
and U26291 (N_26291,N_18365,N_21822);
nor U26292 (N_26292,N_18479,N_19222);
nor U26293 (N_26293,N_20953,N_22768);
or U26294 (N_26294,N_19285,N_23554);
or U26295 (N_26295,N_18207,N_20796);
nor U26296 (N_26296,N_18784,N_22228);
and U26297 (N_26297,N_21179,N_23784);
xnor U26298 (N_26298,N_20685,N_21162);
nor U26299 (N_26299,N_20135,N_22085);
nand U26300 (N_26300,N_21658,N_20136);
or U26301 (N_26301,N_19087,N_20719);
or U26302 (N_26302,N_22961,N_20191);
and U26303 (N_26303,N_23875,N_20905);
nand U26304 (N_26304,N_18372,N_21130);
or U26305 (N_26305,N_20465,N_21394);
or U26306 (N_26306,N_19768,N_18905);
xnor U26307 (N_26307,N_19379,N_20558);
nand U26308 (N_26308,N_23065,N_21101);
xnor U26309 (N_26309,N_19326,N_23216);
and U26310 (N_26310,N_23714,N_22576);
xor U26311 (N_26311,N_18623,N_22611);
nor U26312 (N_26312,N_20585,N_21115);
and U26313 (N_26313,N_21545,N_18186);
nand U26314 (N_26314,N_22990,N_21241);
and U26315 (N_26315,N_19746,N_19734);
and U26316 (N_26316,N_18540,N_21462);
xnor U26317 (N_26317,N_20211,N_21681);
or U26318 (N_26318,N_21326,N_19142);
nor U26319 (N_26319,N_18686,N_23952);
or U26320 (N_26320,N_21930,N_20963);
nor U26321 (N_26321,N_19911,N_23755);
and U26322 (N_26322,N_20156,N_18499);
nand U26323 (N_26323,N_19008,N_18548);
xnor U26324 (N_26324,N_21847,N_21260);
and U26325 (N_26325,N_18079,N_22351);
or U26326 (N_26326,N_20570,N_21410);
nor U26327 (N_26327,N_23988,N_23390);
nand U26328 (N_26328,N_20448,N_21772);
or U26329 (N_26329,N_22353,N_22470);
nor U26330 (N_26330,N_23005,N_18113);
nand U26331 (N_26331,N_21538,N_23950);
and U26332 (N_26332,N_21328,N_20275);
or U26333 (N_26333,N_18822,N_20773);
nand U26334 (N_26334,N_20186,N_19814);
nor U26335 (N_26335,N_21959,N_21321);
nor U26336 (N_26336,N_20302,N_20034);
xor U26337 (N_26337,N_19649,N_18768);
nand U26338 (N_26338,N_22247,N_20277);
nand U26339 (N_26339,N_22216,N_20934);
or U26340 (N_26340,N_18845,N_23545);
nand U26341 (N_26341,N_22689,N_18882);
nor U26342 (N_26342,N_23445,N_21675);
nor U26343 (N_26343,N_22918,N_20898);
xor U26344 (N_26344,N_19258,N_22944);
xnor U26345 (N_26345,N_20529,N_20385);
and U26346 (N_26346,N_21298,N_19254);
xnor U26347 (N_26347,N_18744,N_23147);
nor U26348 (N_26348,N_23630,N_18818);
nand U26349 (N_26349,N_18123,N_20512);
nand U26350 (N_26350,N_18089,N_21026);
nor U26351 (N_26351,N_23297,N_21029);
and U26352 (N_26352,N_19273,N_21089);
nand U26353 (N_26353,N_18659,N_22723);
or U26354 (N_26354,N_18938,N_22720);
nand U26355 (N_26355,N_18903,N_20602);
nand U26356 (N_26356,N_23600,N_21365);
nor U26357 (N_26357,N_21543,N_19444);
or U26358 (N_26358,N_23511,N_20399);
nor U26359 (N_26359,N_21158,N_23313);
nor U26360 (N_26360,N_19223,N_19469);
nor U26361 (N_26361,N_19428,N_22970);
nor U26362 (N_26362,N_21431,N_23279);
nor U26363 (N_26363,N_20945,N_21199);
nor U26364 (N_26364,N_22932,N_21401);
xnor U26365 (N_26365,N_22819,N_21005);
xnor U26366 (N_26366,N_22468,N_19122);
or U26367 (N_26367,N_22348,N_20618);
xor U26368 (N_26368,N_21247,N_19257);
or U26369 (N_26369,N_22782,N_19437);
nor U26370 (N_26370,N_22303,N_20127);
xnor U26371 (N_26371,N_21726,N_18314);
or U26372 (N_26372,N_22362,N_21985);
nor U26373 (N_26373,N_21844,N_20267);
nor U26374 (N_26374,N_22235,N_23622);
nor U26375 (N_26375,N_19621,N_19144);
nand U26376 (N_26376,N_20467,N_22252);
nand U26377 (N_26377,N_19433,N_20639);
xnor U26378 (N_26378,N_19954,N_23121);
and U26379 (N_26379,N_18550,N_18887);
nand U26380 (N_26380,N_18644,N_20712);
nor U26381 (N_26381,N_22381,N_22183);
or U26382 (N_26382,N_20664,N_23473);
nor U26383 (N_26383,N_23004,N_20906);
and U26384 (N_26384,N_20213,N_19561);
nor U26385 (N_26385,N_18042,N_18605);
xor U26386 (N_26386,N_23050,N_19118);
nand U26387 (N_26387,N_23893,N_22395);
xnor U26388 (N_26388,N_21754,N_18629);
xnor U26389 (N_26389,N_18660,N_22688);
nor U26390 (N_26390,N_22061,N_18899);
nor U26391 (N_26391,N_22763,N_19155);
nand U26392 (N_26392,N_23871,N_20078);
and U26393 (N_26393,N_20382,N_20739);
xor U26394 (N_26394,N_18173,N_22159);
or U26395 (N_26395,N_19286,N_22529);
nand U26396 (N_26396,N_18835,N_22220);
xnor U26397 (N_26397,N_19491,N_19811);
nor U26398 (N_26398,N_19628,N_20757);
or U26399 (N_26399,N_23824,N_19058);
or U26400 (N_26400,N_20167,N_22165);
xnor U26401 (N_26401,N_21787,N_20981);
or U26402 (N_26402,N_19461,N_21872);
nor U26403 (N_26403,N_20954,N_19989);
xor U26404 (N_26404,N_19664,N_21918);
xor U26405 (N_26405,N_22887,N_21864);
nor U26406 (N_26406,N_21752,N_19647);
and U26407 (N_26407,N_18035,N_21141);
and U26408 (N_26408,N_23645,N_23849);
nand U26409 (N_26409,N_20337,N_20265);
and U26410 (N_26410,N_21024,N_20549);
nand U26411 (N_26411,N_22662,N_18795);
xor U26412 (N_26412,N_20977,N_22552);
and U26413 (N_26413,N_23951,N_18358);
nor U26414 (N_26414,N_21112,N_23939);
or U26415 (N_26415,N_21023,N_23743);
xnor U26416 (N_26416,N_23909,N_21135);
and U26417 (N_26417,N_18756,N_20958);
xor U26418 (N_26418,N_22837,N_21308);
or U26419 (N_26419,N_22454,N_22453);
or U26420 (N_26420,N_20046,N_22929);
or U26421 (N_26421,N_22790,N_18904);
nand U26422 (N_26422,N_19976,N_22063);
or U26423 (N_26423,N_21432,N_21760);
nor U26424 (N_26424,N_19547,N_20060);
nor U26425 (N_26425,N_20132,N_19073);
xor U26426 (N_26426,N_22802,N_19582);
or U26427 (N_26427,N_23587,N_18356);
or U26428 (N_26428,N_19250,N_19040);
and U26429 (N_26429,N_19955,N_18280);
nor U26430 (N_26430,N_19669,N_18674);
or U26431 (N_26431,N_19889,N_18544);
or U26432 (N_26432,N_23493,N_20827);
nand U26433 (N_26433,N_19207,N_21548);
and U26434 (N_26434,N_23109,N_23792);
xor U26435 (N_26435,N_23383,N_21405);
xnor U26436 (N_26436,N_21495,N_18011);
and U26437 (N_26437,N_20762,N_20783);
or U26438 (N_26438,N_22320,N_21546);
nand U26439 (N_26439,N_21350,N_22868);
nand U26440 (N_26440,N_22844,N_19413);
xnor U26441 (N_26441,N_18796,N_22741);
nor U26442 (N_26442,N_23693,N_22964);
nor U26443 (N_26443,N_23120,N_20947);
or U26444 (N_26444,N_21212,N_21734);
or U26445 (N_26445,N_20162,N_22957);
xor U26446 (N_26446,N_19085,N_21908);
nor U26447 (N_26447,N_20024,N_23816);
nand U26448 (N_26448,N_19881,N_21838);
and U26449 (N_26449,N_19962,N_22388);
and U26450 (N_26450,N_19761,N_19284);
nand U26451 (N_26451,N_20182,N_19823);
and U26452 (N_26452,N_20096,N_18080);
nand U26453 (N_26453,N_19756,N_21507);
xnor U26454 (N_26454,N_22697,N_22923);
xnor U26455 (N_26455,N_22334,N_22283);
xnor U26456 (N_26456,N_19722,N_20777);
nand U26457 (N_26457,N_19941,N_23652);
or U26458 (N_26458,N_18009,N_21821);
nor U26459 (N_26459,N_20680,N_21109);
and U26460 (N_26460,N_22099,N_22436);
or U26461 (N_26461,N_22372,N_20544);
nor U26462 (N_26462,N_21924,N_23961);
nor U26463 (N_26463,N_20744,N_21825);
and U26464 (N_26464,N_19137,N_18253);
xor U26465 (N_26465,N_22444,N_21233);
and U26466 (N_26466,N_22342,N_20683);
nand U26467 (N_26467,N_23880,N_18568);
and U26468 (N_26468,N_23134,N_23305);
nor U26469 (N_26469,N_18529,N_21674);
xnor U26470 (N_26470,N_23904,N_22719);
nor U26471 (N_26471,N_22512,N_19221);
nor U26472 (N_26472,N_19710,N_19584);
nor U26473 (N_26473,N_22864,N_23309);
nand U26474 (N_26474,N_21096,N_18714);
xnor U26475 (N_26475,N_22408,N_21303);
nand U26476 (N_26476,N_21214,N_21899);
nand U26477 (N_26477,N_21015,N_20677);
and U26478 (N_26478,N_23631,N_22330);
xor U26479 (N_26479,N_23854,N_19274);
nor U26480 (N_26480,N_23921,N_19799);
or U26481 (N_26481,N_18527,N_19556);
xnor U26482 (N_26482,N_21878,N_20409);
xnor U26483 (N_26483,N_22951,N_23512);
and U26484 (N_26484,N_19797,N_19272);
nand U26485 (N_26485,N_18867,N_23126);
nand U26486 (N_26486,N_18319,N_23206);
or U26487 (N_26487,N_18994,N_19879);
xor U26488 (N_26488,N_18770,N_20222);
and U26489 (N_26489,N_22760,N_19868);
nor U26490 (N_26490,N_23592,N_18445);
and U26491 (N_26491,N_21997,N_23855);
xnor U26492 (N_26492,N_23790,N_23883);
nor U26493 (N_26493,N_20203,N_19617);
xor U26494 (N_26494,N_18692,N_18016);
xnor U26495 (N_26495,N_18405,N_20968);
nand U26496 (N_26496,N_18961,N_18852);
and U26497 (N_26497,N_22798,N_22389);
and U26498 (N_26498,N_19880,N_19958);
or U26499 (N_26499,N_22282,N_22141);
xor U26500 (N_26500,N_19937,N_21077);
and U26501 (N_26501,N_20054,N_21557);
nor U26502 (N_26502,N_19126,N_22617);
xor U26503 (N_26503,N_18645,N_18243);
nand U26504 (N_26504,N_18066,N_19697);
and U26505 (N_26505,N_23053,N_18273);
nor U26506 (N_26506,N_22361,N_18884);
and U26507 (N_26507,N_18315,N_19262);
and U26508 (N_26508,N_21685,N_22019);
nor U26509 (N_26509,N_19192,N_20888);
and U26510 (N_26510,N_21273,N_23516);
and U26511 (N_26511,N_22383,N_18777);
nor U26512 (N_26512,N_21395,N_23776);
or U26513 (N_26513,N_20973,N_19839);
and U26514 (N_26514,N_20596,N_20290);
nor U26515 (N_26515,N_18541,N_20055);
or U26516 (N_26516,N_18575,N_21553);
nand U26517 (N_26517,N_18934,N_22222);
nor U26518 (N_26518,N_19822,N_20429);
xnor U26519 (N_26519,N_19171,N_18379);
and U26520 (N_26520,N_21283,N_23523);
or U26521 (N_26521,N_22187,N_19033);
nor U26522 (N_26522,N_21583,N_18277);
nand U26523 (N_26523,N_23634,N_20334);
nor U26524 (N_26524,N_22326,N_22924);
xnor U26525 (N_26525,N_23654,N_20551);
nor U26526 (N_26526,N_21043,N_18780);
xnor U26527 (N_26527,N_19975,N_18955);
xor U26528 (N_26528,N_18360,N_21175);
nand U26529 (N_26529,N_18783,N_22639);
nor U26530 (N_26530,N_23992,N_18321);
and U26531 (N_26531,N_22254,N_18538);
xnor U26532 (N_26532,N_19515,N_18431);
and U26533 (N_26533,N_19798,N_21113);
nor U26534 (N_26534,N_20378,N_19802);
and U26535 (N_26535,N_19690,N_23832);
or U26536 (N_26536,N_19776,N_23822);
xnor U26537 (N_26537,N_23990,N_21463);
nor U26538 (N_26538,N_18752,N_21809);
xor U26539 (N_26539,N_20100,N_18942);
and U26540 (N_26540,N_19169,N_23385);
nand U26541 (N_26541,N_22484,N_18816);
nand U26542 (N_26542,N_18034,N_23896);
or U26543 (N_26543,N_18338,N_23085);
nor U26544 (N_26544,N_20356,N_18062);
nor U26545 (N_26545,N_22960,N_19265);
nand U26546 (N_26546,N_18864,N_20892);
or U26547 (N_26547,N_22746,N_21064);
or U26548 (N_26548,N_20478,N_21108);
xnor U26549 (N_26549,N_18140,N_21341);
or U26550 (N_26550,N_20831,N_22127);
and U26551 (N_26551,N_23656,N_21521);
nor U26552 (N_26552,N_21191,N_21182);
nand U26553 (N_26553,N_20297,N_20318);
nand U26554 (N_26554,N_21137,N_20847);
or U26555 (N_26555,N_23192,N_20666);
nand U26556 (N_26556,N_21434,N_18946);
and U26557 (N_26557,N_20486,N_23731);
nand U26558 (N_26558,N_18169,N_18201);
xor U26559 (N_26559,N_22238,N_22332);
nor U26560 (N_26560,N_23330,N_20098);
nor U26561 (N_26561,N_18161,N_18023);
nor U26562 (N_26562,N_23475,N_18260);
nand U26563 (N_26563,N_23454,N_21783);
or U26564 (N_26564,N_22649,N_23821);
nor U26565 (N_26565,N_18065,N_23505);
nand U26566 (N_26566,N_20084,N_23583);
nor U26567 (N_26567,N_20895,N_20266);
nand U26568 (N_26568,N_18897,N_23218);
or U26569 (N_26569,N_22940,N_21730);
and U26570 (N_26570,N_19643,N_22906);
xnor U26571 (N_26571,N_21121,N_23643);
and U26572 (N_26572,N_22861,N_23366);
and U26573 (N_26573,N_21581,N_22817);
nand U26574 (N_26574,N_19831,N_21561);
and U26575 (N_26575,N_19082,N_21547);
nor U26576 (N_26576,N_21446,N_19094);
nor U26577 (N_26577,N_22825,N_19711);
or U26578 (N_26578,N_20748,N_20422);
nand U26579 (N_26579,N_18769,N_23744);
and U26580 (N_26580,N_20955,N_23064);
and U26581 (N_26581,N_18502,N_22904);
nand U26582 (N_26582,N_18621,N_20481);
and U26583 (N_26583,N_19634,N_20094);
or U26584 (N_26584,N_20129,N_22513);
xnor U26585 (N_26585,N_21531,N_18537);
or U26586 (N_26586,N_20488,N_20597);
xnor U26587 (N_26587,N_18391,N_20180);
nor U26588 (N_26588,N_20407,N_18142);
xnor U26589 (N_26589,N_20836,N_18809);
nor U26590 (N_26590,N_20705,N_19060);
and U26591 (N_26591,N_18410,N_21886);
xnor U26592 (N_26592,N_22002,N_23785);
nor U26593 (N_26593,N_21762,N_23489);
nor U26594 (N_26594,N_19191,N_21264);
nand U26595 (N_26595,N_21485,N_21879);
nor U26596 (N_26596,N_21332,N_19052);
and U26597 (N_26597,N_19138,N_21038);
nor U26598 (N_26598,N_21522,N_21944);
xnor U26599 (N_26599,N_22996,N_18128);
xnor U26600 (N_26600,N_23139,N_18944);
or U26601 (N_26601,N_23720,N_21948);
or U26602 (N_26602,N_23781,N_21474);
nor U26603 (N_26603,N_23695,N_22712);
or U26604 (N_26604,N_20787,N_22122);
nor U26605 (N_26605,N_18162,N_18178);
nor U26606 (N_26606,N_21569,N_22240);
or U26607 (N_26607,N_21968,N_21416);
nand U26608 (N_26608,N_19299,N_23588);
or U26609 (N_26609,N_18990,N_19694);
nand U26610 (N_26610,N_23581,N_19774);
nor U26611 (N_26611,N_23948,N_22629);
and U26612 (N_26612,N_22359,N_21794);
nand U26613 (N_26613,N_20051,N_23095);
nor U26614 (N_26614,N_20412,N_23798);
nand U26615 (N_26615,N_23425,N_22386);
and U26616 (N_26616,N_19482,N_22736);
nand U26617 (N_26617,N_23006,N_23531);
nand U26618 (N_26618,N_22628,N_22854);
xnor U26619 (N_26619,N_18613,N_18893);
and U26620 (N_26620,N_20329,N_21700);
and U26621 (N_26621,N_22287,N_20322);
nand U26622 (N_26622,N_23150,N_21300);
or U26623 (N_26623,N_22999,N_20235);
xnor U26624 (N_26624,N_21812,N_22224);
nand U26625 (N_26625,N_19247,N_21361);
nand U26626 (N_26626,N_20020,N_18546);
nand U26627 (N_26627,N_22336,N_21693);
nand U26628 (N_26628,N_21360,N_22142);
xnor U26629 (N_26629,N_23119,N_22998);
nand U26630 (N_26630,N_19038,N_23460);
nand U26631 (N_26631,N_22319,N_21246);
nand U26632 (N_26632,N_20462,N_20737);
xnor U26633 (N_26633,N_23402,N_20471);
or U26634 (N_26634,N_18165,N_23122);
nand U26635 (N_26635,N_22700,N_21050);
nor U26636 (N_26636,N_21611,N_23733);
and U26637 (N_26637,N_20550,N_23838);
or U26638 (N_26638,N_18426,N_21314);
xor U26639 (N_26639,N_18362,N_21200);
xor U26640 (N_26640,N_22588,N_18814);
xnor U26641 (N_26641,N_23788,N_20260);
and U26642 (N_26642,N_19468,N_20072);
or U26643 (N_26643,N_21912,N_22493);
xor U26644 (N_26644,N_22037,N_19436);
nand U26645 (N_26645,N_18120,N_19093);
nor U26646 (N_26646,N_22536,N_19883);
and U26647 (N_26647,N_19606,N_20287);
and U26648 (N_26648,N_18313,N_18074);
nand U26649 (N_26649,N_22227,N_21657);
nand U26650 (N_26650,N_22839,N_18181);
nor U26651 (N_26651,N_21808,N_20818);
xnor U26652 (N_26652,N_21943,N_18301);
nor U26653 (N_26653,N_19302,N_21170);
and U26654 (N_26654,N_21100,N_18239);
and U26655 (N_26655,N_23165,N_19182);
or U26656 (N_26656,N_22401,N_21104);
nand U26657 (N_26657,N_22900,N_21370);
or U26658 (N_26658,N_19885,N_23363);
nand U26659 (N_26659,N_22659,N_22290);
nor U26660 (N_26660,N_23999,N_21996);
xor U26661 (N_26661,N_19785,N_23772);
and U26662 (N_26662,N_21258,N_18545);
xor U26663 (N_26663,N_23107,N_21540);
xnor U26664 (N_26664,N_21407,N_21806);
and U26665 (N_26665,N_21036,N_21168);
xnor U26666 (N_26666,N_21595,N_21862);
xor U26667 (N_26667,N_22909,N_19348);
or U26668 (N_26668,N_18725,N_22791);
or U26669 (N_26669,N_21694,N_19673);
or U26670 (N_26670,N_21711,N_23945);
and U26671 (N_26671,N_18763,N_22086);
or U26672 (N_26672,N_21481,N_19750);
xnor U26673 (N_26673,N_20734,N_20343);
nor U26674 (N_26674,N_23678,N_23691);
nand U26675 (N_26675,N_18675,N_22345);
nand U26676 (N_26676,N_21975,N_20292);
or U26677 (N_26677,N_21443,N_20661);
and U26678 (N_26678,N_20144,N_23994);
or U26679 (N_26679,N_19317,N_23166);
nor U26680 (N_26680,N_19660,N_18246);
nor U26681 (N_26681,N_23611,N_23830);
xor U26682 (N_26682,N_23391,N_21848);
nand U26683 (N_26683,N_20087,N_18054);
and U26684 (N_26684,N_21376,N_21228);
or U26685 (N_26685,N_19787,N_21749);
xnor U26686 (N_26686,N_23012,N_21402);
nor U26687 (N_26687,N_23929,N_23104);
nor U26688 (N_26688,N_18564,N_22634);
xor U26689 (N_26689,N_21946,N_19614);
or U26690 (N_26690,N_19442,N_23210);
xor U26691 (N_26691,N_18191,N_20913);
nor U26692 (N_26692,N_20631,N_21142);
xor U26693 (N_26693,N_18104,N_18370);
and U26694 (N_26694,N_22620,N_23675);
nand U26695 (N_26695,N_23204,N_18580);
xor U26696 (N_26696,N_22396,N_22699);
nor U26697 (N_26697,N_23934,N_19194);
nor U26698 (N_26698,N_19500,N_21305);
or U26699 (N_26699,N_18346,N_20535);
xnor U26700 (N_26700,N_23533,N_23722);
nor U26701 (N_26701,N_18326,N_21718);
nor U26702 (N_26702,N_19061,N_21779);
nand U26703 (N_26703,N_19691,N_20917);
xnor U26704 (N_26704,N_23774,N_20723);
nor U26705 (N_26705,N_20416,N_19332);
and U26706 (N_26706,N_20040,N_19096);
nand U26707 (N_26707,N_20687,N_21986);
or U26708 (N_26708,N_20284,N_22709);
and U26709 (N_26709,N_18749,N_21622);
or U26710 (N_26710,N_19080,N_18100);
or U26711 (N_26711,N_19658,N_18639);
nand U26712 (N_26712,N_21641,N_18010);
xnor U26713 (N_26713,N_20110,N_19923);
nor U26714 (N_26714,N_23133,N_22750);
or U26715 (N_26715,N_21743,N_22415);
nor U26716 (N_26716,N_21002,N_20499);
nand U26717 (N_26717,N_20747,N_19641);
or U26718 (N_26718,N_23418,N_20709);
nor U26719 (N_26719,N_18000,N_22630);
or U26720 (N_26720,N_19167,N_18001);
and U26721 (N_26721,N_19662,N_18494);
and U26722 (N_26722,N_18430,N_23829);
nand U26723 (N_26723,N_18596,N_18627);
and U26724 (N_26724,N_23579,N_19717);
nand U26725 (N_26725,N_22232,N_21192);
nor U26726 (N_26726,N_22652,N_21347);
and U26727 (N_26727,N_18267,N_22856);
or U26728 (N_26728,N_20497,N_19586);
or U26729 (N_26729,N_22312,N_20695);
and U26730 (N_26730,N_19400,N_21380);
nand U26731 (N_26731,N_22559,N_19744);
and U26732 (N_26732,N_23463,N_23024);
nor U26733 (N_26733,N_18117,N_22106);
nor U26734 (N_26734,N_19805,N_22902);
nand U26735 (N_26735,N_21666,N_21269);
nor U26736 (N_26736,N_21334,N_22481);
nand U26737 (N_26737,N_23958,N_23263);
or U26738 (N_26738,N_18402,N_21231);
nand U26739 (N_26739,N_21296,N_19940);
nand U26740 (N_26740,N_19939,N_18229);
and U26741 (N_26741,N_20340,N_20175);
xnor U26742 (N_26742,N_23443,N_19457);
nor U26743 (N_26743,N_19395,N_20327);
and U26744 (N_26744,N_19891,N_20849);
nor U26745 (N_26745,N_21327,N_18482);
and U26746 (N_26746,N_20093,N_19654);
nor U26747 (N_26747,N_20097,N_19545);
or U26748 (N_26748,N_21070,N_19594);
nor U26749 (N_26749,N_20554,N_19423);
nor U26750 (N_26750,N_18423,N_23480);
xnor U26751 (N_26751,N_20363,N_22457);
nand U26752 (N_26752,N_20584,N_20377);
xnor U26753 (N_26753,N_23140,N_20208);
and U26754 (N_26754,N_21775,N_18600);
nor U26755 (N_26755,N_23874,N_23879);
or U26756 (N_26756,N_19692,N_20976);
and U26757 (N_26757,N_20915,N_19339);
and U26758 (N_26758,N_20834,N_18031);
nor U26759 (N_26759,N_20983,N_21756);
nand U26760 (N_26760,N_21673,N_21336);
nand U26761 (N_26761,N_22325,N_21571);
nand U26762 (N_26762,N_22492,N_22528);
nor U26763 (N_26763,N_21902,N_23698);
nor U26764 (N_26764,N_19089,N_20846);
or U26765 (N_26765,N_23417,N_21483);
nor U26766 (N_26766,N_23010,N_18886);
and U26767 (N_26767,N_22363,N_21045);
xor U26768 (N_26768,N_23504,N_18219);
nand U26769 (N_26769,N_21388,N_23853);
nand U26770 (N_26770,N_22810,N_22172);
nand U26771 (N_26771,N_18958,N_21722);
or U26772 (N_26772,N_19427,N_23324);
xnor U26773 (N_26773,N_19236,N_19291);
nor U26774 (N_26774,N_20010,N_18798);
or U26775 (N_26775,N_18082,N_19162);
nor U26776 (N_26776,N_22822,N_19920);
and U26777 (N_26777,N_20058,N_22233);
nor U26778 (N_26778,N_21925,N_21294);
nor U26779 (N_26779,N_19908,N_20682);
nand U26780 (N_26780,N_23321,N_22145);
and U26781 (N_26781,N_21221,N_20791);
nand U26782 (N_26782,N_20311,N_23224);
nor U26783 (N_26783,N_22456,N_23783);
nand U26784 (N_26784,N_21094,N_22664);
nand U26785 (N_26785,N_18119,N_21203);
xnor U26786 (N_26786,N_20288,N_18589);
nor U26787 (N_26787,N_21818,N_19026);
and U26788 (N_26788,N_21068,N_18500);
and U26789 (N_26789,N_18233,N_22495);
and U26790 (N_26790,N_18641,N_22773);
or U26791 (N_26791,N_20565,N_18093);
nand U26792 (N_26792,N_22830,N_20833);
or U26793 (N_26793,N_18508,N_19446);
nand U26794 (N_26794,N_21852,N_20571);
xnor U26795 (N_26795,N_19607,N_18923);
nor U26796 (N_26796,N_23405,N_18988);
and U26797 (N_26797,N_18601,N_20196);
nor U26798 (N_26798,N_18786,N_21172);
xor U26799 (N_26799,N_22623,N_20444);
nor U26800 (N_26800,N_23519,N_19453);
xor U26801 (N_26801,N_18132,N_23663);
and U26802 (N_26802,N_22679,N_19684);
nor U26803 (N_26803,N_20873,N_23362);
and U26804 (N_26804,N_18637,N_19760);
or U26805 (N_26805,N_20746,N_22685);
and U26806 (N_26806,N_18443,N_23408);
and U26807 (N_26807,N_20242,N_22977);
nand U26808 (N_26808,N_23851,N_21954);
nor U26809 (N_26809,N_23866,N_20578);
xnor U26810 (N_26810,N_23775,N_20869);
or U26811 (N_26811,N_18712,N_22098);
xor U26812 (N_26812,N_18471,N_22648);
nor U26813 (N_26813,N_18422,N_20159);
and U26814 (N_26814,N_23474,N_22393);
xor U26815 (N_26815,N_18278,N_22846);
xor U26816 (N_26816,N_23041,N_23542);
nor U26817 (N_26817,N_21498,N_22643);
nand U26818 (N_26818,N_18900,N_23131);
xor U26819 (N_26819,N_23763,N_18779);
nor U26820 (N_26820,N_18741,N_19790);
xor U26821 (N_26821,N_18039,N_18265);
nand U26822 (N_26822,N_23051,N_20047);
nor U26823 (N_26823,N_18295,N_22509);
and U26824 (N_26824,N_18653,N_21022);
nand U26825 (N_26825,N_23738,N_18586);
or U26826 (N_26826,N_18781,N_21785);
or U26827 (N_26827,N_19856,N_21287);
or U26828 (N_26828,N_18325,N_18912);
nand U26829 (N_26829,N_20767,N_20929);
xnor U26830 (N_26830,N_20201,N_18036);
xor U26831 (N_26831,N_19293,N_22466);
xor U26832 (N_26832,N_22562,N_21479);
and U26833 (N_26833,N_23212,N_23159);
and U26834 (N_26834,N_23941,N_19663);
nor U26835 (N_26835,N_20246,N_20032);
or U26836 (N_26836,N_23825,N_23858);
and U26837 (N_26837,N_18983,N_19420);
nand U26838 (N_26838,N_19260,N_18263);
nand U26839 (N_26839,N_20245,N_23767);
xnor U26840 (N_26840,N_23025,N_20930);
nand U26841 (N_26841,N_18689,N_19295);
and U26842 (N_26842,N_18819,N_18192);
or U26843 (N_26843,N_19165,N_22753);
nor U26844 (N_26844,N_22545,N_19041);
nand U26845 (N_26845,N_20583,N_18972);
nand U26846 (N_26846,N_21286,N_19577);
nor U26847 (N_26847,N_22065,N_20147);
xnor U26848 (N_26848,N_18116,N_18440);
and U26849 (N_26849,N_20004,N_22296);
and U26850 (N_26850,N_20749,N_20210);
nor U26851 (N_26851,N_21169,N_18536);
nor U26852 (N_26852,N_19067,N_22658);
nand U26853 (N_26853,N_18070,N_18048);
and U26854 (N_26854,N_18068,N_21651);
nor U26855 (N_26855,N_18985,N_18449);
xor U26856 (N_26856,N_23222,N_18851);
and U26857 (N_26857,N_21608,N_21527);
nand U26858 (N_26858,N_20806,N_22160);
or U26859 (N_26859,N_21251,N_19296);
nand U26860 (N_26860,N_20148,N_21888);
nor U26861 (N_26861,N_19046,N_22548);
nor U26862 (N_26862,N_19288,N_22358);
nor U26863 (N_26863,N_19044,N_22237);
nand U26864 (N_26864,N_20759,N_21056);
and U26865 (N_26865,N_21683,N_20921);
and U26866 (N_26866,N_22508,N_20424);
nor U26867 (N_26867,N_22832,N_18997);
xor U26868 (N_26868,N_22146,N_22058);
nor U26869 (N_26869,N_23901,N_21253);
nor U26870 (N_26870,N_18925,N_20948);
and U26871 (N_26871,N_21164,N_21637);
nand U26872 (N_26872,N_23407,N_19053);
nand U26873 (N_26873,N_23660,N_21117);
nand U26874 (N_26874,N_21737,N_20298);
nor U26875 (N_26875,N_23810,N_23217);
or U26876 (N_26876,N_19519,N_18658);
or U26877 (N_26877,N_19657,N_23799);
nand U26878 (N_26878,N_23040,N_23052);
nand U26879 (N_26879,N_20610,N_20224);
nor U26880 (N_26880,N_18953,N_22540);
or U26881 (N_26881,N_20294,N_18393);
nand U26882 (N_26882,N_22989,N_21733);
and U26883 (N_26883,N_18043,N_22452);
xor U26884 (N_26884,N_21325,N_19015);
xor U26885 (N_26885,N_22498,N_21695);
nand U26886 (N_26886,N_20582,N_21041);
nand U26887 (N_26887,N_18951,N_21449);
nand U26888 (N_26888,N_20142,N_19981);
and U26889 (N_26889,N_22857,N_22632);
and U26890 (N_26890,N_21714,N_20282);
xor U26891 (N_26891,N_22916,N_19788);
or U26892 (N_26892,N_19132,N_23379);
nor U26893 (N_26893,N_20856,N_19571);
xor U26894 (N_26894,N_20434,N_22050);
or U26895 (N_26895,N_22503,N_23687);
nor U26896 (N_26896,N_18556,N_21851);
and U26897 (N_26897,N_19164,N_23627);
and U26898 (N_26898,N_19336,N_21638);
and U26899 (N_26899,N_21180,N_20541);
nand U26900 (N_26900,N_20257,N_21633);
xor U26901 (N_26901,N_20466,N_20950);
or U26902 (N_26902,N_18730,N_22693);
nand U26903 (N_26903,N_21516,N_18224);
and U26904 (N_26904,N_18163,N_19712);
and U26905 (N_26905,N_22757,N_23793);
nor U26906 (N_26906,N_20962,N_22775);
nand U26907 (N_26907,N_20624,N_18481);
nor U26908 (N_26908,N_21340,N_18361);
xor U26909 (N_26909,N_23056,N_20979);
nor U26910 (N_26910,N_19174,N_23090);
or U26911 (N_26911,N_21106,N_19341);
or U26912 (N_26912,N_22236,N_20366);
nand U26913 (N_26913,N_19321,N_19903);
xor U26914 (N_26914,N_22189,N_23233);
nor U26915 (N_26915,N_20067,N_19847);
or U26916 (N_26916,N_21898,N_21994);
and U26917 (N_26917,N_22225,N_21598);
and U26918 (N_26918,N_19591,N_21519);
xor U26919 (N_26919,N_20628,N_20502);
nor U26920 (N_26920,N_23398,N_20788);
and U26921 (N_26921,N_23484,N_21000);
or U26922 (N_26922,N_23088,N_19316);
nand U26923 (N_26923,N_19279,N_21850);
nand U26924 (N_26924,N_19077,N_20433);
and U26925 (N_26925,N_20489,N_21217);
xor U26926 (N_26926,N_21357,N_22304);
and U26927 (N_26927,N_20160,N_19967);
xor U26928 (N_26928,N_19952,N_19076);
xor U26929 (N_26929,N_23890,N_22549);
and U26930 (N_26930,N_20192,N_21609);
or U26931 (N_26931,N_21226,N_21459);
or U26932 (N_26932,N_18759,N_18891);
xnor U26933 (N_26933,N_19970,N_21584);
and U26934 (N_26934,N_22367,N_22422);
or U26935 (N_26935,N_23190,N_20717);
and U26936 (N_26936,N_22459,N_19153);
or U26937 (N_26937,N_22376,N_18976);
xnor U26938 (N_26938,N_18520,N_19780);
or U26939 (N_26939,N_19947,N_23251);
or U26940 (N_26940,N_23528,N_23569);
or U26941 (N_26941,N_18448,N_18936);
or U26942 (N_26942,N_22418,N_19290);
or U26943 (N_26943,N_19995,N_22092);
nor U26944 (N_26944,N_19499,N_21834);
nand U26945 (N_26945,N_21786,N_22407);
or U26946 (N_26946,N_21342,N_20675);
nor U26947 (N_26947,N_23863,N_20845);
or U26948 (N_26948,N_22501,N_21204);
nand U26949 (N_26949,N_20772,N_21566);
or U26950 (N_26950,N_20781,N_20728);
or U26951 (N_26951,N_19984,N_21378);
nand U26952 (N_26952,N_21425,N_18334);
xnor U26953 (N_26953,N_18849,N_23000);
or U26954 (N_26954,N_21549,N_22539);
and U26955 (N_26955,N_20636,N_19160);
and U26956 (N_26956,N_23604,N_22229);
xnor U26957 (N_26957,N_23430,N_22075);
nor U26958 (N_26958,N_19670,N_18480);
xnor U26959 (N_26959,N_21126,N_18122);
xor U26960 (N_26960,N_23485,N_20439);
and U26961 (N_26961,N_18607,N_22182);
nor U26962 (N_26962,N_23180,N_20547);
and U26963 (N_26963,N_19314,N_22892);
or U26964 (N_26964,N_19506,N_19243);
xnor U26965 (N_26965,N_22066,N_22713);
nand U26966 (N_26966,N_20876,N_23154);
and U26967 (N_26967,N_18881,N_19114);
nand U26968 (N_26968,N_20931,N_18915);
nand U26969 (N_26969,N_19512,N_20432);
nor U26970 (N_26970,N_22665,N_23540);
and U26971 (N_26971,N_18063,N_20349);
nor U26972 (N_26972,N_18666,N_19159);
and U26973 (N_26973,N_21574,N_21076);
xnor U26974 (N_26974,N_18830,N_22769);
nand U26975 (N_26975,N_18740,N_19653);
nor U26976 (N_26976,N_19623,N_20673);
nor U26977 (N_26977,N_18367,N_21471);
or U26978 (N_26978,N_19818,N_21796);
nand U26979 (N_26979,N_22574,N_21202);
or U26980 (N_26980,N_19678,N_21923);
nand U26981 (N_26981,N_20633,N_21275);
xnor U26982 (N_26982,N_22421,N_18732);
nand U26983 (N_26983,N_20025,N_21715);
nor U26984 (N_26984,N_19929,N_22928);
xnor U26985 (N_26985,N_22747,N_22446);
nand U26986 (N_26986,N_20248,N_21936);
and U26987 (N_26987,N_22297,N_22555);
or U26988 (N_26988,N_22114,N_20830);
or U26989 (N_26989,N_18108,N_18820);
xnor U26990 (N_26990,N_23325,N_20707);
nor U26991 (N_26991,N_19993,N_19927);
nand U26992 (N_26992,N_21359,N_18204);
xnor U26993 (N_26993,N_23316,N_18750);
nand U26994 (N_26994,N_19996,N_23127);
xor U26995 (N_26995,N_22702,N_21814);
nand U26996 (N_26996,N_20857,N_19635);
nand U26997 (N_26997,N_18432,N_20143);
or U26998 (N_26998,N_21578,N_19567);
or U26999 (N_26999,N_21165,N_18706);
xnor U27000 (N_27000,N_22354,N_19847);
and U27001 (N_27001,N_20177,N_19790);
xnor U27002 (N_27002,N_22663,N_19702);
nand U27003 (N_27003,N_23566,N_23215);
and U27004 (N_27004,N_19254,N_22703);
or U27005 (N_27005,N_19370,N_23614);
xnor U27006 (N_27006,N_18831,N_23230);
nor U27007 (N_27007,N_19077,N_18513);
xor U27008 (N_27008,N_19312,N_21323);
and U27009 (N_27009,N_22644,N_20591);
and U27010 (N_27010,N_18657,N_21131);
and U27011 (N_27011,N_23943,N_20450);
nand U27012 (N_27012,N_20414,N_22354);
nand U27013 (N_27013,N_19732,N_21827);
nand U27014 (N_27014,N_21775,N_18640);
nand U27015 (N_27015,N_23760,N_20514);
nor U27016 (N_27016,N_18966,N_19495);
nor U27017 (N_27017,N_21283,N_22512);
or U27018 (N_27018,N_20647,N_18975);
nor U27019 (N_27019,N_18549,N_18314);
or U27020 (N_27020,N_20407,N_23849);
and U27021 (N_27021,N_23201,N_20995);
nand U27022 (N_27022,N_19131,N_19991);
xnor U27023 (N_27023,N_18375,N_22084);
xor U27024 (N_27024,N_23028,N_19846);
nor U27025 (N_27025,N_22880,N_18775);
xnor U27026 (N_27026,N_20781,N_22031);
or U27027 (N_27027,N_23077,N_23540);
or U27028 (N_27028,N_22977,N_22428);
nand U27029 (N_27029,N_20799,N_23504);
or U27030 (N_27030,N_20415,N_21408);
or U27031 (N_27031,N_23223,N_20411);
or U27032 (N_27032,N_19436,N_18004);
nor U27033 (N_27033,N_19167,N_22385);
xnor U27034 (N_27034,N_18655,N_23512);
nor U27035 (N_27035,N_20096,N_23909);
xnor U27036 (N_27036,N_18844,N_23083);
or U27037 (N_27037,N_18760,N_19733);
xnor U27038 (N_27038,N_20470,N_21766);
nor U27039 (N_27039,N_19780,N_22358);
nor U27040 (N_27040,N_23698,N_18057);
nand U27041 (N_27041,N_23597,N_22952);
xnor U27042 (N_27042,N_23427,N_18078);
or U27043 (N_27043,N_21626,N_23034);
xnor U27044 (N_27044,N_18969,N_22290);
nand U27045 (N_27045,N_21318,N_20707);
or U27046 (N_27046,N_20751,N_19665);
and U27047 (N_27047,N_22068,N_19476);
nor U27048 (N_27048,N_23475,N_21863);
or U27049 (N_27049,N_19698,N_23907);
or U27050 (N_27050,N_21337,N_22810);
nor U27051 (N_27051,N_22827,N_20807);
xor U27052 (N_27052,N_21179,N_20846);
nor U27053 (N_27053,N_22453,N_19678);
and U27054 (N_27054,N_19393,N_20865);
nor U27055 (N_27055,N_20957,N_18253);
or U27056 (N_27056,N_23404,N_18660);
and U27057 (N_27057,N_21855,N_19446);
and U27058 (N_27058,N_23598,N_19934);
nor U27059 (N_27059,N_19834,N_22881);
nand U27060 (N_27060,N_20533,N_20585);
and U27061 (N_27061,N_19431,N_21652);
nand U27062 (N_27062,N_23129,N_22800);
and U27063 (N_27063,N_22692,N_22779);
xor U27064 (N_27064,N_20053,N_22084);
nor U27065 (N_27065,N_19074,N_23475);
nor U27066 (N_27066,N_21874,N_18776);
and U27067 (N_27067,N_22228,N_18903);
xor U27068 (N_27068,N_20125,N_22128);
or U27069 (N_27069,N_18056,N_22789);
nand U27070 (N_27070,N_21510,N_18877);
and U27071 (N_27071,N_18127,N_18001);
nor U27072 (N_27072,N_18707,N_21268);
nand U27073 (N_27073,N_22868,N_23305);
nor U27074 (N_27074,N_20400,N_20438);
nand U27075 (N_27075,N_21019,N_22013);
xor U27076 (N_27076,N_19096,N_20755);
and U27077 (N_27077,N_21507,N_22524);
nand U27078 (N_27078,N_21214,N_23160);
xnor U27079 (N_27079,N_22154,N_21266);
or U27080 (N_27080,N_20460,N_21824);
nand U27081 (N_27081,N_22418,N_21825);
or U27082 (N_27082,N_19418,N_20687);
and U27083 (N_27083,N_21630,N_23277);
or U27084 (N_27084,N_21015,N_19516);
xnor U27085 (N_27085,N_22271,N_18992);
nand U27086 (N_27086,N_23209,N_18101);
nand U27087 (N_27087,N_20682,N_18501);
and U27088 (N_27088,N_23246,N_20706);
nand U27089 (N_27089,N_18366,N_19732);
nor U27090 (N_27090,N_18271,N_20574);
nor U27091 (N_27091,N_22493,N_19590);
or U27092 (N_27092,N_19249,N_21285);
xnor U27093 (N_27093,N_20774,N_21607);
xnor U27094 (N_27094,N_20454,N_20139);
or U27095 (N_27095,N_21671,N_22740);
nor U27096 (N_27096,N_20359,N_22924);
nand U27097 (N_27097,N_18230,N_19867);
nand U27098 (N_27098,N_19876,N_21205);
nor U27099 (N_27099,N_23678,N_20998);
xor U27100 (N_27100,N_23873,N_23679);
and U27101 (N_27101,N_19531,N_19333);
or U27102 (N_27102,N_23357,N_23647);
nand U27103 (N_27103,N_23771,N_21493);
and U27104 (N_27104,N_21039,N_22843);
nand U27105 (N_27105,N_21594,N_23474);
or U27106 (N_27106,N_20008,N_20570);
and U27107 (N_27107,N_23112,N_20818);
xnor U27108 (N_27108,N_23922,N_19408);
xor U27109 (N_27109,N_23981,N_20017);
or U27110 (N_27110,N_21614,N_21903);
or U27111 (N_27111,N_19044,N_20876);
nand U27112 (N_27112,N_20125,N_19127);
nor U27113 (N_27113,N_18307,N_19233);
nor U27114 (N_27114,N_18898,N_23007);
or U27115 (N_27115,N_18783,N_19863);
nor U27116 (N_27116,N_18632,N_19853);
or U27117 (N_27117,N_19576,N_21701);
nor U27118 (N_27118,N_19123,N_23767);
and U27119 (N_27119,N_18851,N_23048);
nor U27120 (N_27120,N_23291,N_21908);
and U27121 (N_27121,N_23237,N_20243);
or U27122 (N_27122,N_23560,N_21441);
and U27123 (N_27123,N_20993,N_21760);
nor U27124 (N_27124,N_22167,N_19952);
and U27125 (N_27125,N_21475,N_20487);
nand U27126 (N_27126,N_18940,N_22145);
or U27127 (N_27127,N_20350,N_18596);
nand U27128 (N_27128,N_23746,N_23506);
nor U27129 (N_27129,N_22645,N_23119);
xor U27130 (N_27130,N_19089,N_18373);
nand U27131 (N_27131,N_19309,N_18758);
xnor U27132 (N_27132,N_18595,N_21958);
xnor U27133 (N_27133,N_19602,N_20780);
nand U27134 (N_27134,N_18156,N_23453);
xnor U27135 (N_27135,N_18333,N_20909);
nor U27136 (N_27136,N_18969,N_23322);
nor U27137 (N_27137,N_18882,N_19717);
xor U27138 (N_27138,N_22692,N_19983);
nand U27139 (N_27139,N_19282,N_22370);
nor U27140 (N_27140,N_23215,N_20625);
or U27141 (N_27141,N_18299,N_18092);
nor U27142 (N_27142,N_21749,N_23668);
and U27143 (N_27143,N_21279,N_21992);
nand U27144 (N_27144,N_23868,N_19380);
nand U27145 (N_27145,N_18202,N_19443);
nand U27146 (N_27146,N_23819,N_19987);
xnor U27147 (N_27147,N_21924,N_23815);
and U27148 (N_27148,N_22760,N_22410);
nand U27149 (N_27149,N_22565,N_23368);
and U27150 (N_27150,N_21252,N_19613);
xnor U27151 (N_27151,N_20942,N_20217);
xnor U27152 (N_27152,N_23147,N_23208);
nand U27153 (N_27153,N_22911,N_19249);
nor U27154 (N_27154,N_21983,N_18163);
and U27155 (N_27155,N_18461,N_18245);
nand U27156 (N_27156,N_18603,N_22221);
nor U27157 (N_27157,N_22938,N_21843);
nand U27158 (N_27158,N_19588,N_20866);
nand U27159 (N_27159,N_18497,N_23403);
nor U27160 (N_27160,N_22825,N_21199);
nand U27161 (N_27161,N_20417,N_23128);
and U27162 (N_27162,N_19515,N_21369);
or U27163 (N_27163,N_21254,N_21385);
and U27164 (N_27164,N_23507,N_18394);
and U27165 (N_27165,N_23342,N_23050);
nand U27166 (N_27166,N_23085,N_23927);
and U27167 (N_27167,N_19039,N_23508);
xnor U27168 (N_27168,N_21330,N_22797);
and U27169 (N_27169,N_19215,N_21267);
nor U27170 (N_27170,N_19636,N_23902);
or U27171 (N_27171,N_18204,N_23946);
or U27172 (N_27172,N_20986,N_23563);
and U27173 (N_27173,N_19103,N_19072);
or U27174 (N_27174,N_20066,N_19988);
xor U27175 (N_27175,N_19258,N_21704);
xnor U27176 (N_27176,N_20056,N_22959);
nand U27177 (N_27177,N_22382,N_19261);
nor U27178 (N_27178,N_22728,N_23018);
nor U27179 (N_27179,N_22666,N_18838);
or U27180 (N_27180,N_23591,N_20337);
xor U27181 (N_27181,N_18088,N_21108);
nand U27182 (N_27182,N_23318,N_19675);
or U27183 (N_27183,N_23434,N_18386);
and U27184 (N_27184,N_19364,N_20781);
and U27185 (N_27185,N_21072,N_19322);
xnor U27186 (N_27186,N_20978,N_22853);
nand U27187 (N_27187,N_23397,N_20656);
xnor U27188 (N_27188,N_18779,N_19205);
xnor U27189 (N_27189,N_22597,N_23994);
and U27190 (N_27190,N_22321,N_21850);
nor U27191 (N_27191,N_21370,N_19976);
and U27192 (N_27192,N_22672,N_23626);
nor U27193 (N_27193,N_23093,N_18057);
xor U27194 (N_27194,N_18471,N_18157);
or U27195 (N_27195,N_22890,N_20137);
and U27196 (N_27196,N_18120,N_21947);
nand U27197 (N_27197,N_22657,N_19439);
or U27198 (N_27198,N_23221,N_21317);
and U27199 (N_27199,N_22430,N_23264);
xor U27200 (N_27200,N_18462,N_22118);
nand U27201 (N_27201,N_23687,N_23738);
xor U27202 (N_27202,N_23635,N_20094);
or U27203 (N_27203,N_19163,N_20494);
or U27204 (N_27204,N_20390,N_18678);
nand U27205 (N_27205,N_19380,N_22657);
nand U27206 (N_27206,N_21722,N_21432);
and U27207 (N_27207,N_23799,N_19337);
nor U27208 (N_27208,N_19892,N_22846);
nand U27209 (N_27209,N_21688,N_19003);
nand U27210 (N_27210,N_22046,N_18035);
xor U27211 (N_27211,N_18904,N_23303);
xnor U27212 (N_27212,N_19573,N_19549);
and U27213 (N_27213,N_20082,N_19203);
nand U27214 (N_27214,N_20660,N_23589);
or U27215 (N_27215,N_23052,N_23580);
nor U27216 (N_27216,N_23209,N_22871);
xor U27217 (N_27217,N_20107,N_21908);
nand U27218 (N_27218,N_22388,N_22594);
nand U27219 (N_27219,N_20972,N_18368);
or U27220 (N_27220,N_22340,N_21741);
and U27221 (N_27221,N_21427,N_18669);
nand U27222 (N_27222,N_22256,N_20621);
and U27223 (N_27223,N_18114,N_21155);
and U27224 (N_27224,N_21933,N_19977);
nor U27225 (N_27225,N_20944,N_21697);
or U27226 (N_27226,N_20496,N_20159);
nand U27227 (N_27227,N_21050,N_21481);
and U27228 (N_27228,N_18789,N_19992);
and U27229 (N_27229,N_21754,N_19118);
and U27230 (N_27230,N_22280,N_20100);
nand U27231 (N_27231,N_22611,N_21526);
xnor U27232 (N_27232,N_22077,N_23498);
or U27233 (N_27233,N_21343,N_23597);
or U27234 (N_27234,N_22331,N_18340);
and U27235 (N_27235,N_21864,N_20100);
or U27236 (N_27236,N_19009,N_21335);
xnor U27237 (N_27237,N_22132,N_18177);
and U27238 (N_27238,N_19459,N_22819);
and U27239 (N_27239,N_18255,N_19160);
or U27240 (N_27240,N_21655,N_20326);
and U27241 (N_27241,N_20968,N_23828);
nor U27242 (N_27242,N_21326,N_23375);
and U27243 (N_27243,N_18218,N_18791);
nand U27244 (N_27244,N_18564,N_22256);
nor U27245 (N_27245,N_23273,N_23738);
and U27246 (N_27246,N_23600,N_22165);
nand U27247 (N_27247,N_20051,N_23910);
nand U27248 (N_27248,N_23529,N_23626);
xnor U27249 (N_27249,N_20954,N_19708);
xor U27250 (N_27250,N_23262,N_19319);
or U27251 (N_27251,N_21268,N_23507);
xor U27252 (N_27252,N_18411,N_18672);
and U27253 (N_27253,N_23768,N_21268);
xor U27254 (N_27254,N_19603,N_21043);
nor U27255 (N_27255,N_19896,N_18069);
and U27256 (N_27256,N_21253,N_21159);
and U27257 (N_27257,N_21112,N_20211);
nor U27258 (N_27258,N_23430,N_21379);
nor U27259 (N_27259,N_18526,N_22365);
nor U27260 (N_27260,N_19681,N_20969);
or U27261 (N_27261,N_23187,N_18780);
xor U27262 (N_27262,N_21135,N_19448);
or U27263 (N_27263,N_23035,N_21697);
or U27264 (N_27264,N_18063,N_19336);
nor U27265 (N_27265,N_18547,N_23195);
or U27266 (N_27266,N_20679,N_21382);
xor U27267 (N_27267,N_20128,N_20909);
and U27268 (N_27268,N_21175,N_18843);
nand U27269 (N_27269,N_20604,N_19845);
xnor U27270 (N_27270,N_22216,N_22248);
or U27271 (N_27271,N_21506,N_23479);
and U27272 (N_27272,N_23140,N_21666);
nor U27273 (N_27273,N_23801,N_21193);
nor U27274 (N_27274,N_23271,N_22110);
and U27275 (N_27275,N_20144,N_19862);
xor U27276 (N_27276,N_20777,N_21341);
nor U27277 (N_27277,N_21268,N_18550);
or U27278 (N_27278,N_21351,N_21295);
xnor U27279 (N_27279,N_19424,N_22064);
nor U27280 (N_27280,N_20278,N_21949);
or U27281 (N_27281,N_19035,N_18590);
nand U27282 (N_27282,N_22766,N_19794);
nand U27283 (N_27283,N_19290,N_21312);
nor U27284 (N_27284,N_23076,N_20363);
nand U27285 (N_27285,N_23957,N_23927);
or U27286 (N_27286,N_20453,N_21025);
nor U27287 (N_27287,N_19460,N_20157);
nand U27288 (N_27288,N_22574,N_18416);
nand U27289 (N_27289,N_19029,N_19549);
xor U27290 (N_27290,N_21437,N_19780);
nand U27291 (N_27291,N_18727,N_18977);
xor U27292 (N_27292,N_20538,N_19504);
nand U27293 (N_27293,N_18947,N_22288);
nand U27294 (N_27294,N_19595,N_21816);
nand U27295 (N_27295,N_19266,N_21737);
xor U27296 (N_27296,N_23581,N_22051);
nor U27297 (N_27297,N_23225,N_20573);
xor U27298 (N_27298,N_23993,N_20771);
nand U27299 (N_27299,N_20829,N_23022);
nor U27300 (N_27300,N_22888,N_21431);
xnor U27301 (N_27301,N_19430,N_20505);
and U27302 (N_27302,N_23276,N_23605);
xnor U27303 (N_27303,N_22482,N_23539);
nor U27304 (N_27304,N_23606,N_20146);
or U27305 (N_27305,N_19503,N_19009);
xor U27306 (N_27306,N_22651,N_19869);
nor U27307 (N_27307,N_23005,N_21479);
nor U27308 (N_27308,N_19027,N_20154);
nor U27309 (N_27309,N_21805,N_22409);
or U27310 (N_27310,N_22435,N_21673);
and U27311 (N_27311,N_21273,N_23386);
and U27312 (N_27312,N_21592,N_21898);
or U27313 (N_27313,N_23185,N_20979);
xnor U27314 (N_27314,N_23781,N_21125);
and U27315 (N_27315,N_20983,N_21640);
nand U27316 (N_27316,N_23316,N_20875);
and U27317 (N_27317,N_18435,N_18407);
xnor U27318 (N_27318,N_19729,N_18266);
nor U27319 (N_27319,N_21205,N_19067);
and U27320 (N_27320,N_18539,N_20633);
nand U27321 (N_27321,N_21713,N_21276);
and U27322 (N_27322,N_21336,N_22800);
xnor U27323 (N_27323,N_20165,N_18326);
nand U27324 (N_27324,N_21310,N_22676);
or U27325 (N_27325,N_21694,N_22788);
or U27326 (N_27326,N_21875,N_22156);
and U27327 (N_27327,N_18462,N_18968);
and U27328 (N_27328,N_18446,N_19793);
and U27329 (N_27329,N_21979,N_18001);
or U27330 (N_27330,N_22600,N_18254);
nor U27331 (N_27331,N_22912,N_20140);
nor U27332 (N_27332,N_23903,N_23232);
nor U27333 (N_27333,N_18053,N_21626);
or U27334 (N_27334,N_21253,N_22625);
and U27335 (N_27335,N_22490,N_23827);
or U27336 (N_27336,N_19398,N_22939);
or U27337 (N_27337,N_19971,N_20477);
nand U27338 (N_27338,N_21004,N_22862);
nor U27339 (N_27339,N_23211,N_23718);
and U27340 (N_27340,N_20384,N_18973);
and U27341 (N_27341,N_19060,N_18037);
or U27342 (N_27342,N_18081,N_21440);
nor U27343 (N_27343,N_19535,N_23436);
nor U27344 (N_27344,N_23182,N_21038);
and U27345 (N_27345,N_20152,N_20906);
nor U27346 (N_27346,N_21787,N_18608);
nand U27347 (N_27347,N_22138,N_21831);
and U27348 (N_27348,N_18043,N_18023);
xnor U27349 (N_27349,N_23533,N_22335);
or U27350 (N_27350,N_20408,N_21001);
nand U27351 (N_27351,N_23664,N_21423);
xor U27352 (N_27352,N_19005,N_20161);
and U27353 (N_27353,N_21436,N_21006);
or U27354 (N_27354,N_19869,N_21539);
nor U27355 (N_27355,N_21785,N_20381);
and U27356 (N_27356,N_18891,N_23316);
and U27357 (N_27357,N_20216,N_18813);
xnor U27358 (N_27358,N_23431,N_23533);
xor U27359 (N_27359,N_23073,N_18720);
and U27360 (N_27360,N_23990,N_19681);
nand U27361 (N_27361,N_22730,N_18521);
or U27362 (N_27362,N_20194,N_22738);
nor U27363 (N_27363,N_21894,N_21854);
xor U27364 (N_27364,N_21047,N_22979);
xnor U27365 (N_27365,N_19093,N_18296);
and U27366 (N_27366,N_23875,N_21680);
xnor U27367 (N_27367,N_22911,N_23270);
nand U27368 (N_27368,N_23792,N_20668);
and U27369 (N_27369,N_20092,N_19727);
or U27370 (N_27370,N_20073,N_22359);
nor U27371 (N_27371,N_23700,N_23934);
and U27372 (N_27372,N_23201,N_21026);
nor U27373 (N_27373,N_21479,N_22805);
nand U27374 (N_27374,N_23396,N_20393);
or U27375 (N_27375,N_21624,N_18727);
xor U27376 (N_27376,N_22307,N_19673);
and U27377 (N_27377,N_20801,N_23664);
nor U27378 (N_27378,N_21646,N_21096);
nor U27379 (N_27379,N_19790,N_21043);
nand U27380 (N_27380,N_20387,N_20259);
xor U27381 (N_27381,N_21064,N_21208);
or U27382 (N_27382,N_22870,N_18948);
and U27383 (N_27383,N_21094,N_20931);
or U27384 (N_27384,N_19161,N_20376);
and U27385 (N_27385,N_20731,N_23296);
and U27386 (N_27386,N_22042,N_23336);
or U27387 (N_27387,N_20515,N_18217);
or U27388 (N_27388,N_21525,N_20170);
xnor U27389 (N_27389,N_19113,N_20693);
xor U27390 (N_27390,N_21603,N_22761);
nand U27391 (N_27391,N_21837,N_22446);
and U27392 (N_27392,N_19418,N_23371);
or U27393 (N_27393,N_19449,N_21681);
xnor U27394 (N_27394,N_19264,N_20533);
and U27395 (N_27395,N_23532,N_22213);
nand U27396 (N_27396,N_18719,N_21778);
and U27397 (N_27397,N_21757,N_18100);
and U27398 (N_27398,N_23677,N_18437);
xor U27399 (N_27399,N_18671,N_21060);
nand U27400 (N_27400,N_23988,N_19185);
xor U27401 (N_27401,N_22167,N_20999);
xnor U27402 (N_27402,N_23648,N_23737);
nand U27403 (N_27403,N_19072,N_23069);
nor U27404 (N_27404,N_19603,N_21091);
xnor U27405 (N_27405,N_23294,N_18780);
xnor U27406 (N_27406,N_22452,N_21538);
and U27407 (N_27407,N_20686,N_22531);
and U27408 (N_27408,N_23839,N_19332);
xor U27409 (N_27409,N_18130,N_19566);
nand U27410 (N_27410,N_23733,N_22035);
nor U27411 (N_27411,N_22324,N_22289);
nor U27412 (N_27412,N_19639,N_23117);
nor U27413 (N_27413,N_23180,N_18373);
and U27414 (N_27414,N_20859,N_18219);
nand U27415 (N_27415,N_19186,N_21167);
nor U27416 (N_27416,N_21157,N_19549);
nand U27417 (N_27417,N_21872,N_23415);
nor U27418 (N_27418,N_20688,N_23181);
nor U27419 (N_27419,N_21467,N_23105);
and U27420 (N_27420,N_20775,N_18956);
xnor U27421 (N_27421,N_22982,N_23491);
xnor U27422 (N_27422,N_22207,N_18339);
nand U27423 (N_27423,N_18057,N_19570);
nor U27424 (N_27424,N_18452,N_23532);
or U27425 (N_27425,N_22789,N_20267);
nand U27426 (N_27426,N_21656,N_18808);
or U27427 (N_27427,N_20396,N_18820);
and U27428 (N_27428,N_21208,N_19802);
or U27429 (N_27429,N_23065,N_19913);
or U27430 (N_27430,N_22664,N_22222);
nand U27431 (N_27431,N_21484,N_20781);
nor U27432 (N_27432,N_23345,N_18752);
nand U27433 (N_27433,N_20174,N_18299);
xnor U27434 (N_27434,N_18444,N_22161);
nand U27435 (N_27435,N_21114,N_20278);
xor U27436 (N_27436,N_21690,N_21415);
or U27437 (N_27437,N_20800,N_19373);
or U27438 (N_27438,N_20334,N_22814);
xor U27439 (N_27439,N_20475,N_19682);
nand U27440 (N_27440,N_22012,N_20153);
and U27441 (N_27441,N_22587,N_18084);
nor U27442 (N_27442,N_20709,N_23987);
nand U27443 (N_27443,N_18728,N_20760);
nand U27444 (N_27444,N_19099,N_20848);
or U27445 (N_27445,N_21075,N_23384);
or U27446 (N_27446,N_19757,N_18917);
nand U27447 (N_27447,N_23476,N_18787);
xor U27448 (N_27448,N_19975,N_21580);
xor U27449 (N_27449,N_22723,N_19669);
xor U27450 (N_27450,N_18194,N_21165);
xnor U27451 (N_27451,N_21956,N_23928);
xnor U27452 (N_27452,N_18511,N_22809);
nor U27453 (N_27453,N_20550,N_22368);
xor U27454 (N_27454,N_19509,N_20763);
or U27455 (N_27455,N_19970,N_20705);
and U27456 (N_27456,N_22380,N_18216);
nand U27457 (N_27457,N_21330,N_18591);
xor U27458 (N_27458,N_23315,N_21583);
or U27459 (N_27459,N_21001,N_22345);
xor U27460 (N_27460,N_18229,N_21716);
or U27461 (N_27461,N_19340,N_20336);
nor U27462 (N_27462,N_22564,N_23366);
and U27463 (N_27463,N_19449,N_22426);
or U27464 (N_27464,N_18285,N_23029);
and U27465 (N_27465,N_19253,N_22018);
nand U27466 (N_27466,N_19904,N_18129);
nor U27467 (N_27467,N_22667,N_23652);
and U27468 (N_27468,N_19946,N_19044);
xor U27469 (N_27469,N_18201,N_19677);
and U27470 (N_27470,N_21708,N_23708);
xor U27471 (N_27471,N_21974,N_19952);
nand U27472 (N_27472,N_19908,N_21845);
nor U27473 (N_27473,N_20876,N_20601);
nand U27474 (N_27474,N_20849,N_23987);
nor U27475 (N_27475,N_21107,N_18736);
or U27476 (N_27476,N_20662,N_23805);
and U27477 (N_27477,N_20437,N_20152);
or U27478 (N_27478,N_22030,N_20007);
and U27479 (N_27479,N_20007,N_19131);
xnor U27480 (N_27480,N_19880,N_21782);
nand U27481 (N_27481,N_19209,N_19928);
nand U27482 (N_27482,N_19850,N_18338);
xor U27483 (N_27483,N_23475,N_20503);
and U27484 (N_27484,N_21038,N_22420);
or U27485 (N_27485,N_23041,N_22458);
nand U27486 (N_27486,N_23756,N_20606);
nand U27487 (N_27487,N_23481,N_23125);
and U27488 (N_27488,N_21189,N_23687);
nor U27489 (N_27489,N_22210,N_22859);
nor U27490 (N_27490,N_19965,N_20533);
and U27491 (N_27491,N_23839,N_20296);
or U27492 (N_27492,N_21297,N_21628);
xor U27493 (N_27493,N_18798,N_20521);
and U27494 (N_27494,N_23237,N_21178);
xor U27495 (N_27495,N_18379,N_19172);
or U27496 (N_27496,N_18453,N_18704);
nor U27497 (N_27497,N_19764,N_23684);
nor U27498 (N_27498,N_21884,N_19942);
nand U27499 (N_27499,N_18670,N_21313);
or U27500 (N_27500,N_23044,N_21513);
xor U27501 (N_27501,N_19647,N_22911);
nor U27502 (N_27502,N_22790,N_18384);
nand U27503 (N_27503,N_19519,N_19760);
xnor U27504 (N_27504,N_18375,N_23151);
and U27505 (N_27505,N_22948,N_20880);
nand U27506 (N_27506,N_23615,N_18058);
and U27507 (N_27507,N_21067,N_22534);
nor U27508 (N_27508,N_21247,N_23445);
xor U27509 (N_27509,N_19947,N_23185);
or U27510 (N_27510,N_19684,N_20411);
or U27511 (N_27511,N_20236,N_22246);
and U27512 (N_27512,N_18340,N_22431);
nor U27513 (N_27513,N_19349,N_18613);
nand U27514 (N_27514,N_22067,N_20238);
nand U27515 (N_27515,N_23546,N_23534);
nor U27516 (N_27516,N_19030,N_18513);
and U27517 (N_27517,N_19386,N_20214);
nand U27518 (N_27518,N_23125,N_22174);
and U27519 (N_27519,N_20965,N_19118);
nand U27520 (N_27520,N_23366,N_22388);
nor U27521 (N_27521,N_20158,N_20646);
nand U27522 (N_27522,N_18839,N_20517);
or U27523 (N_27523,N_18620,N_18213);
nor U27524 (N_27524,N_23025,N_23135);
nor U27525 (N_27525,N_19571,N_20938);
nand U27526 (N_27526,N_18246,N_23925);
or U27527 (N_27527,N_18243,N_21246);
nor U27528 (N_27528,N_20007,N_21683);
nand U27529 (N_27529,N_20978,N_23769);
nand U27530 (N_27530,N_19671,N_21416);
or U27531 (N_27531,N_21986,N_20385);
nand U27532 (N_27532,N_19487,N_19921);
nor U27533 (N_27533,N_19163,N_21840);
xor U27534 (N_27534,N_19691,N_18188);
and U27535 (N_27535,N_19146,N_21665);
nand U27536 (N_27536,N_22132,N_21512);
and U27537 (N_27537,N_23726,N_22838);
xor U27538 (N_27538,N_20310,N_23875);
nand U27539 (N_27539,N_21384,N_19641);
nor U27540 (N_27540,N_21135,N_18497);
xnor U27541 (N_27541,N_18267,N_18426);
nor U27542 (N_27542,N_19171,N_20368);
nor U27543 (N_27543,N_19077,N_23581);
nand U27544 (N_27544,N_22117,N_21047);
nand U27545 (N_27545,N_23874,N_23862);
xnor U27546 (N_27546,N_18561,N_18614);
or U27547 (N_27547,N_18798,N_21610);
xnor U27548 (N_27548,N_19960,N_19872);
or U27549 (N_27549,N_18026,N_22654);
nor U27550 (N_27550,N_18914,N_20577);
xor U27551 (N_27551,N_22049,N_21290);
xor U27552 (N_27552,N_21681,N_18259);
nand U27553 (N_27553,N_20997,N_18074);
nand U27554 (N_27554,N_19578,N_22689);
nand U27555 (N_27555,N_23988,N_19700);
nor U27556 (N_27556,N_20805,N_22407);
xor U27557 (N_27557,N_23878,N_22213);
nand U27558 (N_27558,N_19065,N_23913);
or U27559 (N_27559,N_21777,N_21813);
or U27560 (N_27560,N_22869,N_22854);
nor U27561 (N_27561,N_23951,N_20838);
and U27562 (N_27562,N_23217,N_20859);
xnor U27563 (N_27563,N_23435,N_20682);
and U27564 (N_27564,N_21806,N_19050);
or U27565 (N_27565,N_21221,N_22892);
or U27566 (N_27566,N_19934,N_22195);
xnor U27567 (N_27567,N_18444,N_22172);
and U27568 (N_27568,N_23007,N_20296);
and U27569 (N_27569,N_19819,N_21861);
and U27570 (N_27570,N_18768,N_23417);
xnor U27571 (N_27571,N_18722,N_23312);
and U27572 (N_27572,N_21545,N_22924);
xnor U27573 (N_27573,N_18963,N_23770);
nand U27574 (N_27574,N_23416,N_19925);
xor U27575 (N_27575,N_21775,N_23714);
and U27576 (N_27576,N_22690,N_20248);
and U27577 (N_27577,N_18301,N_23713);
and U27578 (N_27578,N_23496,N_23221);
nor U27579 (N_27579,N_22607,N_21218);
xor U27580 (N_27580,N_18789,N_23360);
and U27581 (N_27581,N_22934,N_18879);
nand U27582 (N_27582,N_18996,N_22989);
xor U27583 (N_27583,N_22872,N_23740);
nor U27584 (N_27584,N_21047,N_21308);
nor U27585 (N_27585,N_18159,N_19421);
nor U27586 (N_27586,N_21278,N_21126);
and U27587 (N_27587,N_20531,N_20543);
and U27588 (N_27588,N_20126,N_22708);
and U27589 (N_27589,N_23901,N_18456);
or U27590 (N_27590,N_23813,N_23941);
nor U27591 (N_27591,N_22400,N_22592);
or U27592 (N_27592,N_21414,N_19144);
and U27593 (N_27593,N_18455,N_18566);
xor U27594 (N_27594,N_18734,N_20202);
nand U27595 (N_27595,N_22904,N_22621);
nor U27596 (N_27596,N_18387,N_23347);
xor U27597 (N_27597,N_18821,N_23947);
or U27598 (N_27598,N_19753,N_19123);
xor U27599 (N_27599,N_23594,N_23238);
and U27600 (N_27600,N_19458,N_20487);
nor U27601 (N_27601,N_20176,N_20655);
nor U27602 (N_27602,N_21405,N_21731);
xor U27603 (N_27603,N_21816,N_18061);
nor U27604 (N_27604,N_23132,N_19812);
xor U27605 (N_27605,N_23013,N_19874);
nand U27606 (N_27606,N_23949,N_20820);
and U27607 (N_27607,N_18062,N_19876);
and U27608 (N_27608,N_20088,N_21080);
or U27609 (N_27609,N_19970,N_20754);
nand U27610 (N_27610,N_21644,N_18531);
xor U27611 (N_27611,N_18059,N_20775);
nand U27612 (N_27612,N_22814,N_20679);
and U27613 (N_27613,N_20725,N_20472);
xor U27614 (N_27614,N_23081,N_19185);
nand U27615 (N_27615,N_21890,N_19850);
nor U27616 (N_27616,N_22853,N_19197);
nand U27617 (N_27617,N_19203,N_19582);
or U27618 (N_27618,N_23676,N_21466);
or U27619 (N_27619,N_20083,N_21881);
nand U27620 (N_27620,N_20896,N_18697);
nand U27621 (N_27621,N_22411,N_21359);
xnor U27622 (N_27622,N_22178,N_18849);
and U27623 (N_27623,N_21830,N_21400);
or U27624 (N_27624,N_20933,N_19596);
and U27625 (N_27625,N_22856,N_18141);
nand U27626 (N_27626,N_19881,N_23275);
xnor U27627 (N_27627,N_21543,N_19379);
nand U27628 (N_27628,N_18200,N_22746);
xor U27629 (N_27629,N_20329,N_21017);
nand U27630 (N_27630,N_20762,N_20995);
or U27631 (N_27631,N_18928,N_18396);
or U27632 (N_27632,N_23448,N_18238);
nor U27633 (N_27633,N_18156,N_18338);
and U27634 (N_27634,N_22268,N_18102);
xnor U27635 (N_27635,N_22272,N_18685);
nor U27636 (N_27636,N_22911,N_23480);
xor U27637 (N_27637,N_22696,N_20327);
nand U27638 (N_27638,N_23804,N_22400);
or U27639 (N_27639,N_19494,N_18886);
nor U27640 (N_27640,N_18054,N_21743);
and U27641 (N_27641,N_20103,N_19490);
or U27642 (N_27642,N_23599,N_19886);
nor U27643 (N_27643,N_18745,N_23240);
nand U27644 (N_27644,N_21537,N_22990);
nor U27645 (N_27645,N_19905,N_18227);
xnor U27646 (N_27646,N_18508,N_18654);
nor U27647 (N_27647,N_23837,N_18762);
xor U27648 (N_27648,N_20121,N_20649);
nor U27649 (N_27649,N_22523,N_18353);
nor U27650 (N_27650,N_23878,N_22306);
xnor U27651 (N_27651,N_20891,N_22695);
nand U27652 (N_27652,N_23487,N_18561);
xor U27653 (N_27653,N_19704,N_18039);
or U27654 (N_27654,N_18591,N_19182);
nand U27655 (N_27655,N_19394,N_22717);
xnor U27656 (N_27656,N_23666,N_18207);
or U27657 (N_27657,N_21201,N_22948);
nor U27658 (N_27658,N_21998,N_20570);
xor U27659 (N_27659,N_22842,N_21859);
or U27660 (N_27660,N_19623,N_22103);
nor U27661 (N_27661,N_23924,N_23083);
and U27662 (N_27662,N_23627,N_21732);
and U27663 (N_27663,N_23188,N_20652);
or U27664 (N_27664,N_22202,N_23354);
or U27665 (N_27665,N_18231,N_23442);
nor U27666 (N_27666,N_19602,N_23481);
nand U27667 (N_27667,N_20106,N_18434);
nor U27668 (N_27668,N_22732,N_22054);
nor U27669 (N_27669,N_23663,N_19615);
or U27670 (N_27670,N_18129,N_23104);
and U27671 (N_27671,N_18956,N_18609);
xnor U27672 (N_27672,N_22897,N_21053);
nor U27673 (N_27673,N_23973,N_19110);
and U27674 (N_27674,N_22461,N_18885);
nand U27675 (N_27675,N_23914,N_20250);
xnor U27676 (N_27676,N_18526,N_19360);
or U27677 (N_27677,N_23648,N_22979);
and U27678 (N_27678,N_20374,N_23660);
or U27679 (N_27679,N_18017,N_21938);
nor U27680 (N_27680,N_21180,N_18561);
nor U27681 (N_27681,N_23114,N_18374);
nand U27682 (N_27682,N_22052,N_20857);
xor U27683 (N_27683,N_19729,N_23786);
nor U27684 (N_27684,N_18865,N_19013);
or U27685 (N_27685,N_23708,N_20251);
xnor U27686 (N_27686,N_23129,N_18786);
and U27687 (N_27687,N_18865,N_21915);
xor U27688 (N_27688,N_22579,N_20998);
xor U27689 (N_27689,N_20140,N_21017);
nand U27690 (N_27690,N_21231,N_19881);
xor U27691 (N_27691,N_23498,N_21425);
nor U27692 (N_27692,N_23484,N_23395);
or U27693 (N_27693,N_23934,N_22851);
nor U27694 (N_27694,N_18196,N_18416);
and U27695 (N_27695,N_18476,N_22656);
xor U27696 (N_27696,N_19246,N_22161);
and U27697 (N_27697,N_19150,N_18450);
or U27698 (N_27698,N_20926,N_19882);
nand U27699 (N_27699,N_19668,N_20594);
xor U27700 (N_27700,N_21126,N_19976);
and U27701 (N_27701,N_23722,N_20692);
nand U27702 (N_27702,N_21987,N_22818);
or U27703 (N_27703,N_21602,N_23829);
and U27704 (N_27704,N_21131,N_23158);
nor U27705 (N_27705,N_19133,N_20234);
nand U27706 (N_27706,N_23147,N_23590);
xor U27707 (N_27707,N_22344,N_23993);
nor U27708 (N_27708,N_19209,N_23235);
nor U27709 (N_27709,N_19821,N_23255);
nand U27710 (N_27710,N_19210,N_21350);
nand U27711 (N_27711,N_21269,N_22947);
xor U27712 (N_27712,N_22127,N_21677);
nand U27713 (N_27713,N_20042,N_23582);
xor U27714 (N_27714,N_18961,N_22790);
nor U27715 (N_27715,N_18324,N_20631);
nor U27716 (N_27716,N_23527,N_21581);
nor U27717 (N_27717,N_18811,N_19522);
and U27718 (N_27718,N_19971,N_23519);
xor U27719 (N_27719,N_21268,N_18934);
or U27720 (N_27720,N_18899,N_19777);
and U27721 (N_27721,N_21223,N_21820);
and U27722 (N_27722,N_21622,N_23781);
nor U27723 (N_27723,N_21406,N_20685);
nand U27724 (N_27724,N_19948,N_18379);
xnor U27725 (N_27725,N_19765,N_23068);
or U27726 (N_27726,N_23301,N_18028);
xor U27727 (N_27727,N_19236,N_21249);
xnor U27728 (N_27728,N_19398,N_20292);
nor U27729 (N_27729,N_21252,N_19429);
xnor U27730 (N_27730,N_22439,N_19151);
xor U27731 (N_27731,N_19184,N_23689);
nor U27732 (N_27732,N_23055,N_20951);
or U27733 (N_27733,N_23583,N_20218);
or U27734 (N_27734,N_20112,N_22098);
xor U27735 (N_27735,N_20065,N_20294);
and U27736 (N_27736,N_19736,N_21755);
and U27737 (N_27737,N_20226,N_21561);
nor U27738 (N_27738,N_20216,N_18901);
and U27739 (N_27739,N_18305,N_22404);
and U27740 (N_27740,N_21656,N_20686);
xor U27741 (N_27741,N_22974,N_20300);
and U27742 (N_27742,N_21582,N_23737);
nor U27743 (N_27743,N_19569,N_23008);
nor U27744 (N_27744,N_23391,N_21165);
and U27745 (N_27745,N_22506,N_22402);
or U27746 (N_27746,N_18298,N_19593);
and U27747 (N_27747,N_23654,N_21151);
nand U27748 (N_27748,N_20571,N_23822);
xor U27749 (N_27749,N_18063,N_20563);
and U27750 (N_27750,N_19252,N_22616);
xor U27751 (N_27751,N_18701,N_18883);
nor U27752 (N_27752,N_21059,N_21488);
xnor U27753 (N_27753,N_22331,N_18748);
and U27754 (N_27754,N_19020,N_21647);
xnor U27755 (N_27755,N_18698,N_18661);
and U27756 (N_27756,N_19103,N_19978);
nand U27757 (N_27757,N_18099,N_19148);
and U27758 (N_27758,N_22834,N_19459);
nor U27759 (N_27759,N_21933,N_21634);
nand U27760 (N_27760,N_22430,N_22169);
nand U27761 (N_27761,N_20402,N_21255);
or U27762 (N_27762,N_20731,N_21326);
nor U27763 (N_27763,N_23043,N_18376);
or U27764 (N_27764,N_23402,N_21756);
nand U27765 (N_27765,N_20000,N_19864);
xnor U27766 (N_27766,N_21981,N_23150);
and U27767 (N_27767,N_22261,N_19842);
nand U27768 (N_27768,N_19624,N_23049);
nand U27769 (N_27769,N_23689,N_18618);
or U27770 (N_27770,N_20201,N_22779);
nor U27771 (N_27771,N_23380,N_19737);
xor U27772 (N_27772,N_22813,N_19201);
and U27773 (N_27773,N_18663,N_21975);
nor U27774 (N_27774,N_23339,N_22295);
nor U27775 (N_27775,N_23935,N_22214);
nor U27776 (N_27776,N_19978,N_20786);
nor U27777 (N_27777,N_23697,N_19907);
nand U27778 (N_27778,N_18414,N_23037);
nor U27779 (N_27779,N_18973,N_21096);
nor U27780 (N_27780,N_18776,N_20708);
or U27781 (N_27781,N_20329,N_21997);
xor U27782 (N_27782,N_20857,N_22967);
or U27783 (N_27783,N_22996,N_18012);
nor U27784 (N_27784,N_22066,N_22613);
nand U27785 (N_27785,N_18711,N_18470);
nand U27786 (N_27786,N_19749,N_23328);
xnor U27787 (N_27787,N_22270,N_19312);
and U27788 (N_27788,N_22996,N_19273);
and U27789 (N_27789,N_18373,N_23707);
nand U27790 (N_27790,N_18916,N_21131);
xnor U27791 (N_27791,N_23896,N_20346);
nand U27792 (N_27792,N_23636,N_19040);
nor U27793 (N_27793,N_18083,N_22206);
nor U27794 (N_27794,N_23087,N_18136);
xor U27795 (N_27795,N_20412,N_18116);
xor U27796 (N_27796,N_23228,N_23421);
nor U27797 (N_27797,N_21506,N_22610);
xnor U27798 (N_27798,N_18261,N_23101);
nor U27799 (N_27799,N_19677,N_18896);
nor U27800 (N_27800,N_20960,N_20025);
or U27801 (N_27801,N_18876,N_20161);
and U27802 (N_27802,N_19543,N_18985);
xnor U27803 (N_27803,N_23790,N_23143);
xor U27804 (N_27804,N_20064,N_19799);
nand U27805 (N_27805,N_19102,N_22838);
nand U27806 (N_27806,N_18893,N_20408);
or U27807 (N_27807,N_19517,N_20928);
nor U27808 (N_27808,N_22841,N_20084);
nand U27809 (N_27809,N_18346,N_23431);
xnor U27810 (N_27810,N_20207,N_18296);
and U27811 (N_27811,N_21389,N_18847);
or U27812 (N_27812,N_23002,N_23322);
nand U27813 (N_27813,N_19848,N_20518);
nand U27814 (N_27814,N_21730,N_23875);
and U27815 (N_27815,N_22874,N_20968);
nand U27816 (N_27816,N_19205,N_22263);
xnor U27817 (N_27817,N_18049,N_19397);
and U27818 (N_27818,N_22794,N_18415);
nor U27819 (N_27819,N_18720,N_19349);
nor U27820 (N_27820,N_23007,N_18086);
and U27821 (N_27821,N_21318,N_20747);
xnor U27822 (N_27822,N_18182,N_20600);
or U27823 (N_27823,N_18749,N_20526);
and U27824 (N_27824,N_20421,N_23007);
nand U27825 (N_27825,N_20493,N_20981);
and U27826 (N_27826,N_22997,N_21046);
nand U27827 (N_27827,N_20434,N_20625);
nand U27828 (N_27828,N_20500,N_19371);
nand U27829 (N_27829,N_20149,N_23250);
xor U27830 (N_27830,N_18293,N_19126);
xnor U27831 (N_27831,N_20091,N_18669);
or U27832 (N_27832,N_19095,N_23039);
xor U27833 (N_27833,N_23734,N_18657);
or U27834 (N_27834,N_22590,N_18877);
nand U27835 (N_27835,N_22064,N_23893);
and U27836 (N_27836,N_23954,N_20357);
xor U27837 (N_27837,N_20929,N_23064);
nor U27838 (N_27838,N_18754,N_23553);
and U27839 (N_27839,N_22379,N_23233);
nor U27840 (N_27840,N_23762,N_23928);
nand U27841 (N_27841,N_19025,N_20221);
xor U27842 (N_27842,N_23799,N_21295);
nor U27843 (N_27843,N_19593,N_18451);
nand U27844 (N_27844,N_19177,N_19081);
nor U27845 (N_27845,N_23791,N_19764);
and U27846 (N_27846,N_22168,N_22357);
nand U27847 (N_27847,N_23355,N_19463);
nand U27848 (N_27848,N_19742,N_23528);
and U27849 (N_27849,N_18103,N_21358);
xnor U27850 (N_27850,N_19496,N_23559);
or U27851 (N_27851,N_20833,N_21140);
nor U27852 (N_27852,N_18566,N_23593);
or U27853 (N_27853,N_18428,N_23663);
xnor U27854 (N_27854,N_23768,N_18146);
nor U27855 (N_27855,N_19759,N_21249);
nor U27856 (N_27856,N_21749,N_22899);
or U27857 (N_27857,N_20615,N_22733);
and U27858 (N_27858,N_23741,N_21134);
xor U27859 (N_27859,N_21493,N_21510);
xnor U27860 (N_27860,N_20746,N_18974);
nor U27861 (N_27861,N_22683,N_23976);
or U27862 (N_27862,N_19518,N_20725);
or U27863 (N_27863,N_20972,N_23280);
or U27864 (N_27864,N_20563,N_20725);
xnor U27865 (N_27865,N_18851,N_20684);
xor U27866 (N_27866,N_22410,N_19120);
nand U27867 (N_27867,N_22658,N_21995);
or U27868 (N_27868,N_22558,N_22172);
and U27869 (N_27869,N_21572,N_19221);
xor U27870 (N_27870,N_23779,N_21678);
nand U27871 (N_27871,N_21682,N_22980);
or U27872 (N_27872,N_23074,N_21425);
and U27873 (N_27873,N_19260,N_19764);
nor U27874 (N_27874,N_18369,N_18174);
nand U27875 (N_27875,N_20181,N_23392);
nor U27876 (N_27876,N_23454,N_23862);
nand U27877 (N_27877,N_20442,N_20656);
xnor U27878 (N_27878,N_21971,N_23788);
nor U27879 (N_27879,N_18150,N_18245);
nor U27880 (N_27880,N_21946,N_22145);
nor U27881 (N_27881,N_23653,N_18533);
and U27882 (N_27882,N_20388,N_23468);
or U27883 (N_27883,N_19515,N_21646);
or U27884 (N_27884,N_21965,N_19626);
and U27885 (N_27885,N_18509,N_22427);
xor U27886 (N_27886,N_21353,N_18531);
xor U27887 (N_27887,N_22058,N_19886);
or U27888 (N_27888,N_21658,N_20110);
and U27889 (N_27889,N_20890,N_21372);
or U27890 (N_27890,N_20039,N_22505);
or U27891 (N_27891,N_22133,N_20350);
or U27892 (N_27892,N_18359,N_23840);
nand U27893 (N_27893,N_20902,N_23383);
nor U27894 (N_27894,N_20464,N_22458);
or U27895 (N_27895,N_19623,N_21417);
or U27896 (N_27896,N_21343,N_23755);
nand U27897 (N_27897,N_20133,N_23888);
nor U27898 (N_27898,N_18388,N_19953);
nand U27899 (N_27899,N_18730,N_22778);
nor U27900 (N_27900,N_20197,N_22673);
or U27901 (N_27901,N_18904,N_19192);
and U27902 (N_27902,N_23961,N_19046);
or U27903 (N_27903,N_21280,N_20470);
and U27904 (N_27904,N_18490,N_21345);
nand U27905 (N_27905,N_19138,N_22046);
nand U27906 (N_27906,N_19356,N_18397);
or U27907 (N_27907,N_20319,N_20416);
xor U27908 (N_27908,N_18201,N_22609);
and U27909 (N_27909,N_18448,N_20820);
nor U27910 (N_27910,N_18572,N_20902);
or U27911 (N_27911,N_18496,N_21510);
xor U27912 (N_27912,N_21519,N_18140);
or U27913 (N_27913,N_19640,N_21490);
and U27914 (N_27914,N_21702,N_22258);
nand U27915 (N_27915,N_22361,N_21464);
nand U27916 (N_27916,N_22434,N_20136);
and U27917 (N_27917,N_22417,N_18581);
and U27918 (N_27918,N_23722,N_20540);
nor U27919 (N_27919,N_22045,N_21193);
nor U27920 (N_27920,N_21815,N_23922);
or U27921 (N_27921,N_18370,N_21011);
nor U27922 (N_27922,N_20430,N_21131);
or U27923 (N_27923,N_20546,N_22384);
xor U27924 (N_27924,N_22765,N_19751);
xor U27925 (N_27925,N_18218,N_19285);
and U27926 (N_27926,N_23554,N_20514);
nand U27927 (N_27927,N_21425,N_22148);
or U27928 (N_27928,N_20848,N_18778);
nor U27929 (N_27929,N_21896,N_18217);
nor U27930 (N_27930,N_21917,N_18014);
and U27931 (N_27931,N_19900,N_22117);
nand U27932 (N_27932,N_21955,N_23939);
nand U27933 (N_27933,N_21356,N_18145);
xnor U27934 (N_27934,N_20043,N_21979);
nand U27935 (N_27935,N_18262,N_23130);
nor U27936 (N_27936,N_18207,N_19202);
or U27937 (N_27937,N_18951,N_21172);
nand U27938 (N_27938,N_18016,N_20241);
xnor U27939 (N_27939,N_18780,N_20289);
xnor U27940 (N_27940,N_19816,N_18096);
xnor U27941 (N_27941,N_23243,N_22699);
or U27942 (N_27942,N_19004,N_20738);
or U27943 (N_27943,N_18106,N_23138);
or U27944 (N_27944,N_23360,N_19435);
or U27945 (N_27945,N_22643,N_22052);
and U27946 (N_27946,N_19710,N_21089);
xor U27947 (N_27947,N_18886,N_19031);
or U27948 (N_27948,N_22467,N_21326);
or U27949 (N_27949,N_20467,N_23502);
nor U27950 (N_27950,N_23172,N_19906);
or U27951 (N_27951,N_23416,N_20989);
or U27952 (N_27952,N_18126,N_22370);
nor U27953 (N_27953,N_22641,N_23135);
or U27954 (N_27954,N_18098,N_19423);
and U27955 (N_27955,N_18426,N_20544);
nand U27956 (N_27956,N_22957,N_20065);
and U27957 (N_27957,N_18449,N_20319);
nor U27958 (N_27958,N_19863,N_23288);
xnor U27959 (N_27959,N_22001,N_21715);
or U27960 (N_27960,N_23120,N_22336);
xor U27961 (N_27961,N_22326,N_22552);
nor U27962 (N_27962,N_19517,N_22930);
nor U27963 (N_27963,N_21523,N_22513);
nand U27964 (N_27964,N_18889,N_23075);
xor U27965 (N_27965,N_20535,N_22753);
nand U27966 (N_27966,N_19757,N_19759);
xnor U27967 (N_27967,N_19246,N_18571);
nor U27968 (N_27968,N_20868,N_23811);
nand U27969 (N_27969,N_23421,N_20691);
and U27970 (N_27970,N_23464,N_23972);
and U27971 (N_27971,N_20206,N_19879);
and U27972 (N_27972,N_22155,N_21680);
nor U27973 (N_27973,N_21871,N_21343);
or U27974 (N_27974,N_20036,N_18990);
nor U27975 (N_27975,N_23146,N_23455);
xnor U27976 (N_27976,N_18247,N_18035);
nor U27977 (N_27977,N_19688,N_23799);
nand U27978 (N_27978,N_21281,N_20747);
and U27979 (N_27979,N_19242,N_18703);
nand U27980 (N_27980,N_18267,N_20555);
nand U27981 (N_27981,N_22881,N_18551);
xnor U27982 (N_27982,N_22109,N_20120);
and U27983 (N_27983,N_18078,N_21367);
or U27984 (N_27984,N_23109,N_20042);
nor U27985 (N_27985,N_20579,N_22919);
and U27986 (N_27986,N_19389,N_23110);
and U27987 (N_27987,N_23657,N_20670);
and U27988 (N_27988,N_18522,N_19858);
xnor U27989 (N_27989,N_18461,N_19135);
and U27990 (N_27990,N_20355,N_19847);
nand U27991 (N_27991,N_19545,N_18308);
xor U27992 (N_27992,N_23866,N_21585);
nor U27993 (N_27993,N_21000,N_19656);
nand U27994 (N_27994,N_19917,N_23227);
xnor U27995 (N_27995,N_18025,N_21625);
nor U27996 (N_27996,N_18173,N_23325);
nor U27997 (N_27997,N_19854,N_21969);
nand U27998 (N_27998,N_21310,N_19833);
and U27999 (N_27999,N_18927,N_22069);
nand U28000 (N_28000,N_21861,N_18827);
xnor U28001 (N_28001,N_18458,N_19429);
nand U28002 (N_28002,N_18725,N_19714);
nand U28003 (N_28003,N_20360,N_22846);
xnor U28004 (N_28004,N_23843,N_18123);
xor U28005 (N_28005,N_22751,N_20804);
or U28006 (N_28006,N_19051,N_20196);
or U28007 (N_28007,N_21897,N_22181);
nor U28008 (N_28008,N_19386,N_20278);
or U28009 (N_28009,N_22102,N_21609);
nand U28010 (N_28010,N_18553,N_20031);
or U28011 (N_28011,N_21890,N_18107);
or U28012 (N_28012,N_22929,N_20984);
and U28013 (N_28013,N_22585,N_19429);
nand U28014 (N_28014,N_22937,N_21526);
nand U28015 (N_28015,N_18228,N_23801);
nand U28016 (N_28016,N_23063,N_21118);
nand U28017 (N_28017,N_22171,N_18690);
xor U28018 (N_28018,N_21385,N_18751);
xor U28019 (N_28019,N_21658,N_22600);
nand U28020 (N_28020,N_18547,N_22660);
nor U28021 (N_28021,N_19184,N_19182);
nor U28022 (N_28022,N_21143,N_18498);
and U28023 (N_28023,N_21407,N_23791);
nand U28024 (N_28024,N_19945,N_18618);
nor U28025 (N_28025,N_22040,N_20611);
nor U28026 (N_28026,N_20627,N_22028);
xnor U28027 (N_28027,N_22859,N_19153);
nand U28028 (N_28028,N_20874,N_19964);
nor U28029 (N_28029,N_22958,N_19177);
and U28030 (N_28030,N_22871,N_20798);
and U28031 (N_28031,N_18030,N_19456);
or U28032 (N_28032,N_23361,N_21263);
and U28033 (N_28033,N_21694,N_18457);
or U28034 (N_28034,N_19038,N_22015);
nor U28035 (N_28035,N_20148,N_19988);
nand U28036 (N_28036,N_19820,N_22035);
nand U28037 (N_28037,N_21623,N_22132);
or U28038 (N_28038,N_19998,N_19594);
nand U28039 (N_28039,N_21086,N_21521);
and U28040 (N_28040,N_20614,N_23835);
or U28041 (N_28041,N_18616,N_19650);
or U28042 (N_28042,N_21920,N_21676);
nor U28043 (N_28043,N_21141,N_21983);
xnor U28044 (N_28044,N_21638,N_23649);
nor U28045 (N_28045,N_21907,N_23898);
or U28046 (N_28046,N_18722,N_21170);
or U28047 (N_28047,N_18917,N_22360);
and U28048 (N_28048,N_20167,N_19699);
xnor U28049 (N_28049,N_22253,N_21927);
nand U28050 (N_28050,N_22430,N_23442);
nor U28051 (N_28051,N_22710,N_20961);
or U28052 (N_28052,N_21879,N_23929);
or U28053 (N_28053,N_23152,N_22523);
or U28054 (N_28054,N_18641,N_20888);
nor U28055 (N_28055,N_21370,N_21669);
and U28056 (N_28056,N_22141,N_23362);
nor U28057 (N_28057,N_19897,N_18361);
or U28058 (N_28058,N_23885,N_20598);
or U28059 (N_28059,N_20762,N_20041);
or U28060 (N_28060,N_22918,N_21413);
nand U28061 (N_28061,N_18777,N_21206);
nor U28062 (N_28062,N_20241,N_18591);
xor U28063 (N_28063,N_18027,N_19949);
nand U28064 (N_28064,N_18089,N_21915);
xor U28065 (N_28065,N_18559,N_23062);
and U28066 (N_28066,N_18033,N_19000);
or U28067 (N_28067,N_23405,N_20111);
and U28068 (N_28068,N_22630,N_22941);
xnor U28069 (N_28069,N_18167,N_19919);
xnor U28070 (N_28070,N_19445,N_22241);
xor U28071 (N_28071,N_19088,N_19675);
and U28072 (N_28072,N_18952,N_22793);
nand U28073 (N_28073,N_18937,N_20824);
or U28074 (N_28074,N_23968,N_19187);
nand U28075 (N_28075,N_18007,N_19334);
or U28076 (N_28076,N_23489,N_19226);
nor U28077 (N_28077,N_18486,N_20424);
and U28078 (N_28078,N_19433,N_21592);
nand U28079 (N_28079,N_19182,N_22112);
nand U28080 (N_28080,N_18438,N_18029);
nor U28081 (N_28081,N_23668,N_23856);
or U28082 (N_28082,N_19598,N_22980);
nor U28083 (N_28083,N_21603,N_20619);
or U28084 (N_28084,N_19912,N_20635);
xnor U28085 (N_28085,N_23618,N_19510);
nand U28086 (N_28086,N_19591,N_23863);
nor U28087 (N_28087,N_23280,N_23013);
nand U28088 (N_28088,N_18791,N_21996);
xor U28089 (N_28089,N_20389,N_22104);
or U28090 (N_28090,N_21802,N_19974);
and U28091 (N_28091,N_23372,N_22733);
and U28092 (N_28092,N_23040,N_23959);
or U28093 (N_28093,N_19518,N_20822);
nor U28094 (N_28094,N_19505,N_19443);
xnor U28095 (N_28095,N_19280,N_22127);
or U28096 (N_28096,N_22774,N_22299);
nor U28097 (N_28097,N_18397,N_21452);
or U28098 (N_28098,N_23965,N_20404);
nand U28099 (N_28099,N_19752,N_22052);
nand U28100 (N_28100,N_22484,N_23282);
and U28101 (N_28101,N_19341,N_21994);
and U28102 (N_28102,N_23319,N_21490);
or U28103 (N_28103,N_19676,N_21175);
xnor U28104 (N_28104,N_19516,N_19283);
nor U28105 (N_28105,N_21903,N_20567);
or U28106 (N_28106,N_20207,N_18630);
nor U28107 (N_28107,N_21640,N_20606);
or U28108 (N_28108,N_23510,N_20005);
nand U28109 (N_28109,N_22510,N_20100);
nand U28110 (N_28110,N_23854,N_21691);
xor U28111 (N_28111,N_22368,N_19304);
and U28112 (N_28112,N_23390,N_22915);
or U28113 (N_28113,N_20838,N_22594);
and U28114 (N_28114,N_18281,N_20225);
and U28115 (N_28115,N_22358,N_19822);
nand U28116 (N_28116,N_19462,N_23847);
and U28117 (N_28117,N_20750,N_21108);
nand U28118 (N_28118,N_23984,N_19951);
nand U28119 (N_28119,N_19872,N_19604);
xnor U28120 (N_28120,N_21501,N_21932);
nor U28121 (N_28121,N_23877,N_21022);
nand U28122 (N_28122,N_19543,N_18468);
and U28123 (N_28123,N_18187,N_18387);
xnor U28124 (N_28124,N_20766,N_18348);
xor U28125 (N_28125,N_21780,N_21735);
nor U28126 (N_28126,N_20890,N_22169);
and U28127 (N_28127,N_19669,N_18102);
or U28128 (N_28128,N_18917,N_18148);
nand U28129 (N_28129,N_19453,N_18411);
nor U28130 (N_28130,N_20311,N_22465);
nor U28131 (N_28131,N_21462,N_20266);
or U28132 (N_28132,N_22976,N_18838);
xnor U28133 (N_28133,N_21855,N_21730);
or U28134 (N_28134,N_20002,N_19716);
xnor U28135 (N_28135,N_21682,N_21724);
nor U28136 (N_28136,N_20847,N_20726);
nor U28137 (N_28137,N_18843,N_21740);
nand U28138 (N_28138,N_21310,N_23795);
or U28139 (N_28139,N_23519,N_22095);
nand U28140 (N_28140,N_23317,N_23607);
and U28141 (N_28141,N_19659,N_19717);
nand U28142 (N_28142,N_18720,N_22746);
and U28143 (N_28143,N_18363,N_22003);
nand U28144 (N_28144,N_19181,N_19394);
xor U28145 (N_28145,N_20404,N_22471);
xor U28146 (N_28146,N_21733,N_18675);
nor U28147 (N_28147,N_20738,N_21067);
and U28148 (N_28148,N_20497,N_22115);
nor U28149 (N_28149,N_23889,N_22736);
nand U28150 (N_28150,N_22106,N_21653);
or U28151 (N_28151,N_23576,N_22997);
nand U28152 (N_28152,N_23845,N_23471);
and U28153 (N_28153,N_22398,N_18071);
and U28154 (N_28154,N_21309,N_19562);
nor U28155 (N_28155,N_23775,N_18323);
and U28156 (N_28156,N_22737,N_23357);
and U28157 (N_28157,N_21283,N_19283);
xnor U28158 (N_28158,N_19126,N_23751);
xnor U28159 (N_28159,N_21814,N_20079);
nor U28160 (N_28160,N_21377,N_22853);
nor U28161 (N_28161,N_19828,N_21988);
nand U28162 (N_28162,N_21027,N_21059);
xnor U28163 (N_28163,N_18112,N_19183);
nor U28164 (N_28164,N_23201,N_18344);
nor U28165 (N_28165,N_23634,N_23230);
and U28166 (N_28166,N_22348,N_19812);
xnor U28167 (N_28167,N_20156,N_19473);
or U28168 (N_28168,N_18035,N_21168);
or U28169 (N_28169,N_22498,N_22554);
nor U28170 (N_28170,N_21554,N_21051);
or U28171 (N_28171,N_22064,N_18014);
or U28172 (N_28172,N_21881,N_23816);
and U28173 (N_28173,N_22225,N_23134);
nand U28174 (N_28174,N_23245,N_20363);
nand U28175 (N_28175,N_22086,N_21768);
nand U28176 (N_28176,N_22360,N_20415);
or U28177 (N_28177,N_19250,N_20030);
or U28178 (N_28178,N_19374,N_21916);
and U28179 (N_28179,N_18029,N_20025);
nand U28180 (N_28180,N_22764,N_19501);
nor U28181 (N_28181,N_19643,N_23252);
nor U28182 (N_28182,N_20458,N_19973);
xnor U28183 (N_28183,N_19137,N_22136);
and U28184 (N_28184,N_18568,N_21442);
or U28185 (N_28185,N_19553,N_20343);
nand U28186 (N_28186,N_21438,N_19046);
nand U28187 (N_28187,N_19106,N_22039);
or U28188 (N_28188,N_20779,N_21545);
nor U28189 (N_28189,N_21347,N_18633);
or U28190 (N_28190,N_18082,N_22933);
or U28191 (N_28191,N_22581,N_18156);
and U28192 (N_28192,N_22786,N_23766);
xnor U28193 (N_28193,N_21573,N_23096);
nor U28194 (N_28194,N_18111,N_18376);
or U28195 (N_28195,N_23081,N_18829);
xor U28196 (N_28196,N_18190,N_23706);
nor U28197 (N_28197,N_19612,N_22290);
xnor U28198 (N_28198,N_18087,N_22643);
nand U28199 (N_28199,N_22454,N_18455);
and U28200 (N_28200,N_22616,N_23453);
xnor U28201 (N_28201,N_19388,N_21181);
and U28202 (N_28202,N_20856,N_18690);
nand U28203 (N_28203,N_21114,N_23689);
xnor U28204 (N_28204,N_22770,N_22885);
xor U28205 (N_28205,N_22894,N_19779);
nor U28206 (N_28206,N_18327,N_19611);
nor U28207 (N_28207,N_22399,N_22773);
xor U28208 (N_28208,N_22799,N_18384);
and U28209 (N_28209,N_21185,N_18547);
nor U28210 (N_28210,N_22200,N_23706);
nand U28211 (N_28211,N_22431,N_18303);
nor U28212 (N_28212,N_22091,N_21411);
or U28213 (N_28213,N_19309,N_19345);
nor U28214 (N_28214,N_20292,N_23119);
and U28215 (N_28215,N_23435,N_21575);
nor U28216 (N_28216,N_20823,N_23313);
nand U28217 (N_28217,N_22172,N_18189);
xor U28218 (N_28218,N_18233,N_20116);
or U28219 (N_28219,N_22823,N_18652);
nand U28220 (N_28220,N_20287,N_19461);
and U28221 (N_28221,N_19448,N_21931);
or U28222 (N_28222,N_20079,N_20166);
nor U28223 (N_28223,N_19923,N_19105);
or U28224 (N_28224,N_20274,N_22790);
nor U28225 (N_28225,N_23037,N_18009);
nor U28226 (N_28226,N_21864,N_19691);
nand U28227 (N_28227,N_23385,N_21482);
nor U28228 (N_28228,N_21147,N_22754);
and U28229 (N_28229,N_18496,N_19931);
nor U28230 (N_28230,N_21985,N_19398);
and U28231 (N_28231,N_22159,N_21203);
and U28232 (N_28232,N_20531,N_23685);
nor U28233 (N_28233,N_18601,N_22171);
nand U28234 (N_28234,N_22647,N_22101);
and U28235 (N_28235,N_18641,N_22601);
xor U28236 (N_28236,N_18790,N_21915);
or U28237 (N_28237,N_19404,N_21657);
nor U28238 (N_28238,N_23964,N_22021);
nor U28239 (N_28239,N_18234,N_21396);
nor U28240 (N_28240,N_19362,N_20577);
or U28241 (N_28241,N_23121,N_23744);
nand U28242 (N_28242,N_20985,N_23363);
xnor U28243 (N_28243,N_18835,N_23231);
nand U28244 (N_28244,N_22704,N_19578);
and U28245 (N_28245,N_19829,N_23141);
nor U28246 (N_28246,N_22706,N_23848);
nand U28247 (N_28247,N_19273,N_22740);
xor U28248 (N_28248,N_20049,N_19261);
nand U28249 (N_28249,N_20951,N_18818);
xor U28250 (N_28250,N_21316,N_18444);
and U28251 (N_28251,N_20017,N_21145);
or U28252 (N_28252,N_19042,N_18977);
xor U28253 (N_28253,N_21281,N_22342);
nand U28254 (N_28254,N_19141,N_23166);
xnor U28255 (N_28255,N_20168,N_21597);
nor U28256 (N_28256,N_22611,N_20715);
xor U28257 (N_28257,N_19586,N_19469);
nand U28258 (N_28258,N_21420,N_20460);
and U28259 (N_28259,N_18310,N_21716);
xor U28260 (N_28260,N_20096,N_22664);
nand U28261 (N_28261,N_18063,N_22187);
nor U28262 (N_28262,N_21771,N_21728);
or U28263 (N_28263,N_23726,N_18067);
or U28264 (N_28264,N_22350,N_18483);
and U28265 (N_28265,N_18285,N_22436);
xnor U28266 (N_28266,N_23508,N_19997);
nand U28267 (N_28267,N_19298,N_23164);
nor U28268 (N_28268,N_22472,N_22788);
nand U28269 (N_28269,N_21543,N_23244);
or U28270 (N_28270,N_21868,N_18020);
or U28271 (N_28271,N_22793,N_19221);
and U28272 (N_28272,N_20494,N_18098);
xor U28273 (N_28273,N_23469,N_23427);
or U28274 (N_28274,N_23268,N_18406);
or U28275 (N_28275,N_22941,N_19183);
nand U28276 (N_28276,N_23547,N_21685);
nand U28277 (N_28277,N_19084,N_22779);
or U28278 (N_28278,N_20217,N_22218);
and U28279 (N_28279,N_18892,N_23283);
nor U28280 (N_28280,N_23405,N_21954);
nand U28281 (N_28281,N_22649,N_21543);
nor U28282 (N_28282,N_21359,N_22723);
nand U28283 (N_28283,N_23643,N_19939);
nand U28284 (N_28284,N_20398,N_20872);
and U28285 (N_28285,N_20110,N_23329);
nand U28286 (N_28286,N_20734,N_22556);
nor U28287 (N_28287,N_20380,N_19900);
nand U28288 (N_28288,N_23759,N_21268);
and U28289 (N_28289,N_22782,N_18756);
xor U28290 (N_28290,N_21829,N_23429);
or U28291 (N_28291,N_21957,N_21526);
xnor U28292 (N_28292,N_21868,N_20940);
xor U28293 (N_28293,N_19978,N_19151);
xor U28294 (N_28294,N_22300,N_21906);
and U28295 (N_28295,N_22688,N_18727);
nand U28296 (N_28296,N_18594,N_23921);
xor U28297 (N_28297,N_19428,N_20240);
or U28298 (N_28298,N_22251,N_18355);
nor U28299 (N_28299,N_19079,N_21651);
xnor U28300 (N_28300,N_23453,N_20934);
xnor U28301 (N_28301,N_20372,N_19713);
nand U28302 (N_28302,N_18357,N_21564);
nor U28303 (N_28303,N_18040,N_18618);
nor U28304 (N_28304,N_18692,N_19164);
xor U28305 (N_28305,N_23559,N_23217);
and U28306 (N_28306,N_23692,N_18330);
xnor U28307 (N_28307,N_23693,N_23510);
and U28308 (N_28308,N_22503,N_20434);
xor U28309 (N_28309,N_23923,N_18134);
nor U28310 (N_28310,N_22035,N_19336);
nand U28311 (N_28311,N_22054,N_21316);
and U28312 (N_28312,N_18765,N_19468);
or U28313 (N_28313,N_22291,N_18907);
and U28314 (N_28314,N_22371,N_18707);
nand U28315 (N_28315,N_18565,N_21534);
xnor U28316 (N_28316,N_22240,N_22940);
nor U28317 (N_28317,N_23875,N_23504);
xor U28318 (N_28318,N_21419,N_21328);
or U28319 (N_28319,N_22801,N_21994);
nand U28320 (N_28320,N_22955,N_22238);
or U28321 (N_28321,N_21698,N_22285);
nor U28322 (N_28322,N_20577,N_22961);
nor U28323 (N_28323,N_23420,N_19081);
nand U28324 (N_28324,N_19120,N_18167);
xnor U28325 (N_28325,N_21939,N_18506);
nor U28326 (N_28326,N_20993,N_18528);
nand U28327 (N_28327,N_19103,N_20925);
nor U28328 (N_28328,N_18655,N_23677);
or U28329 (N_28329,N_19598,N_21436);
or U28330 (N_28330,N_18579,N_18469);
nor U28331 (N_28331,N_19272,N_23559);
nor U28332 (N_28332,N_22127,N_18229);
xnor U28333 (N_28333,N_18842,N_19230);
and U28334 (N_28334,N_22151,N_21867);
or U28335 (N_28335,N_23252,N_20902);
and U28336 (N_28336,N_20122,N_20380);
nor U28337 (N_28337,N_20019,N_21350);
nand U28338 (N_28338,N_23672,N_21047);
xnor U28339 (N_28339,N_22252,N_20614);
nand U28340 (N_28340,N_23101,N_21326);
xnor U28341 (N_28341,N_23081,N_22862);
and U28342 (N_28342,N_18493,N_19352);
or U28343 (N_28343,N_22468,N_22922);
nand U28344 (N_28344,N_20007,N_23270);
and U28345 (N_28345,N_20162,N_23408);
nand U28346 (N_28346,N_19461,N_22055);
nor U28347 (N_28347,N_21205,N_23696);
and U28348 (N_28348,N_21543,N_21711);
or U28349 (N_28349,N_21176,N_22989);
and U28350 (N_28350,N_20662,N_23116);
and U28351 (N_28351,N_19397,N_21148);
nor U28352 (N_28352,N_23519,N_18184);
nor U28353 (N_28353,N_20430,N_21501);
and U28354 (N_28354,N_23603,N_22342);
xor U28355 (N_28355,N_21843,N_19891);
nor U28356 (N_28356,N_21405,N_23360);
nor U28357 (N_28357,N_22829,N_21725);
or U28358 (N_28358,N_23656,N_20979);
nand U28359 (N_28359,N_23149,N_20154);
xnor U28360 (N_28360,N_21558,N_18882);
and U28361 (N_28361,N_21169,N_19169);
nand U28362 (N_28362,N_19682,N_18827);
or U28363 (N_28363,N_20508,N_18932);
nor U28364 (N_28364,N_20193,N_19580);
and U28365 (N_28365,N_18757,N_21265);
and U28366 (N_28366,N_21656,N_20947);
nand U28367 (N_28367,N_18565,N_20864);
and U28368 (N_28368,N_22540,N_19151);
or U28369 (N_28369,N_22699,N_19706);
nor U28370 (N_28370,N_21365,N_21892);
nand U28371 (N_28371,N_18746,N_19464);
nand U28372 (N_28372,N_18319,N_20360);
nand U28373 (N_28373,N_19895,N_18031);
nor U28374 (N_28374,N_18167,N_21465);
and U28375 (N_28375,N_19635,N_23577);
or U28376 (N_28376,N_20129,N_19808);
nor U28377 (N_28377,N_20515,N_18027);
nand U28378 (N_28378,N_23027,N_19848);
and U28379 (N_28379,N_21597,N_22740);
and U28380 (N_28380,N_22885,N_19692);
and U28381 (N_28381,N_18776,N_19876);
nand U28382 (N_28382,N_19262,N_20366);
xor U28383 (N_28383,N_20482,N_23174);
nand U28384 (N_28384,N_18474,N_18085);
and U28385 (N_28385,N_22754,N_21856);
and U28386 (N_28386,N_20362,N_21356);
or U28387 (N_28387,N_23569,N_23269);
xnor U28388 (N_28388,N_22591,N_18733);
nand U28389 (N_28389,N_18911,N_22796);
and U28390 (N_28390,N_20598,N_19751);
or U28391 (N_28391,N_23887,N_21162);
nor U28392 (N_28392,N_23121,N_20132);
or U28393 (N_28393,N_23425,N_23449);
nor U28394 (N_28394,N_20157,N_22227);
nand U28395 (N_28395,N_19972,N_18920);
nand U28396 (N_28396,N_18286,N_21202);
and U28397 (N_28397,N_21002,N_19397);
or U28398 (N_28398,N_22421,N_18510);
nor U28399 (N_28399,N_22669,N_20437);
xor U28400 (N_28400,N_18299,N_19966);
xnor U28401 (N_28401,N_21536,N_18664);
nand U28402 (N_28402,N_21542,N_18050);
xor U28403 (N_28403,N_21570,N_19573);
or U28404 (N_28404,N_22170,N_21230);
nor U28405 (N_28405,N_20040,N_23273);
or U28406 (N_28406,N_23024,N_19444);
nor U28407 (N_28407,N_19849,N_18259);
xor U28408 (N_28408,N_19780,N_23160);
xnor U28409 (N_28409,N_22630,N_22162);
or U28410 (N_28410,N_23920,N_19491);
or U28411 (N_28411,N_19989,N_21823);
nand U28412 (N_28412,N_22438,N_19459);
or U28413 (N_28413,N_21756,N_23004);
and U28414 (N_28414,N_23798,N_19924);
and U28415 (N_28415,N_22978,N_20143);
and U28416 (N_28416,N_21770,N_19467);
and U28417 (N_28417,N_18170,N_22246);
nor U28418 (N_28418,N_18944,N_19006);
or U28419 (N_28419,N_18555,N_23708);
nor U28420 (N_28420,N_21199,N_20594);
or U28421 (N_28421,N_19446,N_20771);
nand U28422 (N_28422,N_21622,N_21035);
or U28423 (N_28423,N_23686,N_21103);
or U28424 (N_28424,N_23617,N_18237);
and U28425 (N_28425,N_19187,N_18268);
or U28426 (N_28426,N_22984,N_22884);
and U28427 (N_28427,N_23023,N_19405);
nand U28428 (N_28428,N_23678,N_20928);
xor U28429 (N_28429,N_22463,N_22456);
nor U28430 (N_28430,N_21957,N_19107);
and U28431 (N_28431,N_21975,N_23952);
nor U28432 (N_28432,N_22800,N_20680);
and U28433 (N_28433,N_18285,N_19259);
nand U28434 (N_28434,N_18943,N_21662);
nand U28435 (N_28435,N_22909,N_19784);
xor U28436 (N_28436,N_20770,N_22968);
or U28437 (N_28437,N_19926,N_20197);
nor U28438 (N_28438,N_18880,N_20849);
nor U28439 (N_28439,N_21031,N_23311);
or U28440 (N_28440,N_19931,N_22459);
nand U28441 (N_28441,N_20785,N_22672);
xor U28442 (N_28442,N_21051,N_22624);
or U28443 (N_28443,N_20247,N_19573);
xnor U28444 (N_28444,N_21025,N_22776);
and U28445 (N_28445,N_22429,N_21630);
and U28446 (N_28446,N_19779,N_22740);
xor U28447 (N_28447,N_22642,N_18881);
or U28448 (N_28448,N_20040,N_20681);
or U28449 (N_28449,N_19199,N_21450);
and U28450 (N_28450,N_21385,N_22864);
or U28451 (N_28451,N_23779,N_21237);
nand U28452 (N_28452,N_22471,N_22218);
nand U28453 (N_28453,N_23396,N_23509);
nor U28454 (N_28454,N_19045,N_19249);
nor U28455 (N_28455,N_19276,N_20749);
or U28456 (N_28456,N_20154,N_20412);
nor U28457 (N_28457,N_21678,N_21567);
nand U28458 (N_28458,N_21121,N_23220);
nand U28459 (N_28459,N_21567,N_21970);
nand U28460 (N_28460,N_20990,N_22878);
and U28461 (N_28461,N_22065,N_18753);
and U28462 (N_28462,N_20601,N_20284);
and U28463 (N_28463,N_18197,N_20660);
xnor U28464 (N_28464,N_23489,N_21679);
xor U28465 (N_28465,N_20985,N_19840);
or U28466 (N_28466,N_21756,N_19415);
and U28467 (N_28467,N_19365,N_18590);
or U28468 (N_28468,N_19440,N_20397);
and U28469 (N_28469,N_22744,N_18644);
or U28470 (N_28470,N_21303,N_22644);
xnor U28471 (N_28471,N_19530,N_20078);
nand U28472 (N_28472,N_23394,N_20905);
or U28473 (N_28473,N_21850,N_23813);
xnor U28474 (N_28474,N_22597,N_20106);
nor U28475 (N_28475,N_19311,N_18551);
and U28476 (N_28476,N_23163,N_23202);
and U28477 (N_28477,N_23640,N_18222);
xor U28478 (N_28478,N_18601,N_20632);
and U28479 (N_28479,N_21526,N_19537);
nor U28480 (N_28480,N_22593,N_20998);
or U28481 (N_28481,N_22042,N_20575);
and U28482 (N_28482,N_18014,N_20928);
nand U28483 (N_28483,N_22360,N_22052);
nor U28484 (N_28484,N_18839,N_23553);
and U28485 (N_28485,N_18515,N_22515);
xnor U28486 (N_28486,N_22862,N_22418);
xnor U28487 (N_28487,N_22588,N_22776);
nand U28488 (N_28488,N_22219,N_20677);
xnor U28489 (N_28489,N_20772,N_23774);
and U28490 (N_28490,N_22337,N_19402);
nand U28491 (N_28491,N_19364,N_22123);
nor U28492 (N_28492,N_18347,N_21377);
nand U28493 (N_28493,N_21551,N_19356);
and U28494 (N_28494,N_23760,N_20691);
xor U28495 (N_28495,N_22382,N_19362);
or U28496 (N_28496,N_20049,N_20198);
nor U28497 (N_28497,N_19833,N_20744);
and U28498 (N_28498,N_20112,N_18875);
nand U28499 (N_28499,N_22624,N_21302);
or U28500 (N_28500,N_19346,N_19690);
nand U28501 (N_28501,N_18633,N_19166);
xnor U28502 (N_28502,N_18685,N_19500);
nand U28503 (N_28503,N_23895,N_21624);
or U28504 (N_28504,N_19794,N_20678);
or U28505 (N_28505,N_21611,N_20830);
nor U28506 (N_28506,N_20288,N_18187);
nand U28507 (N_28507,N_20931,N_19019);
xor U28508 (N_28508,N_22484,N_20847);
nand U28509 (N_28509,N_21784,N_22667);
and U28510 (N_28510,N_21872,N_19580);
and U28511 (N_28511,N_20008,N_21949);
xor U28512 (N_28512,N_20481,N_21328);
and U28513 (N_28513,N_20476,N_22565);
nor U28514 (N_28514,N_20568,N_23474);
or U28515 (N_28515,N_18503,N_19015);
nor U28516 (N_28516,N_23025,N_20704);
and U28517 (N_28517,N_19765,N_21465);
nor U28518 (N_28518,N_20022,N_21429);
xor U28519 (N_28519,N_18986,N_18854);
nor U28520 (N_28520,N_19964,N_23581);
or U28521 (N_28521,N_23761,N_23113);
nand U28522 (N_28522,N_19394,N_18185);
nor U28523 (N_28523,N_18382,N_18943);
and U28524 (N_28524,N_23298,N_20840);
or U28525 (N_28525,N_22789,N_20767);
nand U28526 (N_28526,N_21092,N_23021);
nand U28527 (N_28527,N_21324,N_22804);
or U28528 (N_28528,N_22789,N_19735);
xnor U28529 (N_28529,N_22263,N_19084);
and U28530 (N_28530,N_21920,N_23155);
or U28531 (N_28531,N_23130,N_23652);
nor U28532 (N_28532,N_18845,N_20513);
nor U28533 (N_28533,N_18100,N_20696);
or U28534 (N_28534,N_22709,N_18908);
nor U28535 (N_28535,N_21375,N_22027);
nor U28536 (N_28536,N_18759,N_19365);
nor U28537 (N_28537,N_18021,N_22589);
or U28538 (N_28538,N_21810,N_18200);
xnor U28539 (N_28539,N_20810,N_19572);
and U28540 (N_28540,N_20686,N_18961);
xnor U28541 (N_28541,N_22083,N_18483);
or U28542 (N_28542,N_18667,N_21683);
and U28543 (N_28543,N_18778,N_18931);
or U28544 (N_28544,N_20106,N_19309);
nand U28545 (N_28545,N_22933,N_23235);
or U28546 (N_28546,N_23119,N_21613);
nand U28547 (N_28547,N_21754,N_20170);
xnor U28548 (N_28548,N_18777,N_23048);
xor U28549 (N_28549,N_19880,N_20477);
xor U28550 (N_28550,N_20914,N_20473);
and U28551 (N_28551,N_22584,N_18245);
nor U28552 (N_28552,N_20555,N_22330);
and U28553 (N_28553,N_22551,N_22894);
or U28554 (N_28554,N_18307,N_20054);
and U28555 (N_28555,N_22654,N_19384);
or U28556 (N_28556,N_21412,N_21444);
and U28557 (N_28557,N_21519,N_21429);
or U28558 (N_28558,N_22682,N_22844);
nand U28559 (N_28559,N_22758,N_19740);
nor U28560 (N_28560,N_19603,N_23817);
nor U28561 (N_28561,N_18176,N_21362);
and U28562 (N_28562,N_23480,N_18734);
xnor U28563 (N_28563,N_19224,N_18019);
and U28564 (N_28564,N_23341,N_22060);
xor U28565 (N_28565,N_23196,N_19772);
xnor U28566 (N_28566,N_18178,N_21418);
and U28567 (N_28567,N_19546,N_23405);
nand U28568 (N_28568,N_18037,N_20718);
nand U28569 (N_28569,N_23067,N_23203);
nor U28570 (N_28570,N_20387,N_19308);
and U28571 (N_28571,N_22420,N_23682);
nor U28572 (N_28572,N_21331,N_23262);
and U28573 (N_28573,N_18416,N_23994);
nand U28574 (N_28574,N_18368,N_19174);
nor U28575 (N_28575,N_18390,N_21363);
nor U28576 (N_28576,N_18984,N_19926);
and U28577 (N_28577,N_23099,N_21937);
or U28578 (N_28578,N_19734,N_18914);
nor U28579 (N_28579,N_22041,N_23497);
xnor U28580 (N_28580,N_19880,N_20084);
nand U28581 (N_28581,N_18635,N_18470);
and U28582 (N_28582,N_23982,N_19789);
nand U28583 (N_28583,N_23964,N_23845);
nand U28584 (N_28584,N_23312,N_19986);
nand U28585 (N_28585,N_20359,N_22909);
and U28586 (N_28586,N_19981,N_19583);
nor U28587 (N_28587,N_19314,N_20346);
or U28588 (N_28588,N_23098,N_21954);
nor U28589 (N_28589,N_20001,N_23352);
nor U28590 (N_28590,N_23207,N_23944);
nor U28591 (N_28591,N_21345,N_21277);
or U28592 (N_28592,N_19509,N_19322);
or U28593 (N_28593,N_20059,N_23762);
and U28594 (N_28594,N_18407,N_18133);
nand U28595 (N_28595,N_18910,N_19452);
nor U28596 (N_28596,N_23845,N_18060);
nand U28597 (N_28597,N_19204,N_20052);
nand U28598 (N_28598,N_21432,N_22743);
xor U28599 (N_28599,N_22801,N_23913);
nor U28600 (N_28600,N_19668,N_20102);
xnor U28601 (N_28601,N_19839,N_20916);
nand U28602 (N_28602,N_23158,N_21555);
xor U28603 (N_28603,N_19564,N_18831);
and U28604 (N_28604,N_21395,N_20253);
xnor U28605 (N_28605,N_23142,N_22433);
xnor U28606 (N_28606,N_22908,N_18762);
xor U28607 (N_28607,N_23642,N_20612);
nand U28608 (N_28608,N_18086,N_21028);
nand U28609 (N_28609,N_19728,N_18141);
xor U28610 (N_28610,N_19017,N_18357);
and U28611 (N_28611,N_21816,N_22335);
xor U28612 (N_28612,N_22266,N_20832);
or U28613 (N_28613,N_18953,N_20200);
xor U28614 (N_28614,N_21038,N_21161);
nand U28615 (N_28615,N_19065,N_21937);
and U28616 (N_28616,N_20703,N_22673);
nand U28617 (N_28617,N_18160,N_19077);
xor U28618 (N_28618,N_23859,N_20238);
xor U28619 (N_28619,N_22719,N_23448);
xnor U28620 (N_28620,N_20786,N_23560);
nand U28621 (N_28621,N_20019,N_23003);
xnor U28622 (N_28622,N_21153,N_18463);
and U28623 (N_28623,N_18879,N_18091);
nand U28624 (N_28624,N_22965,N_20152);
xnor U28625 (N_28625,N_20271,N_22082);
or U28626 (N_28626,N_18829,N_22198);
nor U28627 (N_28627,N_22490,N_18101);
and U28628 (N_28628,N_22228,N_19196);
and U28629 (N_28629,N_21834,N_19281);
or U28630 (N_28630,N_22341,N_23535);
nor U28631 (N_28631,N_18312,N_18423);
nand U28632 (N_28632,N_20550,N_22967);
nor U28633 (N_28633,N_20996,N_20559);
nor U28634 (N_28634,N_23320,N_22734);
xnor U28635 (N_28635,N_19612,N_22663);
xor U28636 (N_28636,N_23163,N_19248);
nor U28637 (N_28637,N_19218,N_20120);
nand U28638 (N_28638,N_22299,N_20597);
and U28639 (N_28639,N_21539,N_21197);
nor U28640 (N_28640,N_19594,N_22396);
and U28641 (N_28641,N_18851,N_18969);
nor U28642 (N_28642,N_20261,N_23080);
nor U28643 (N_28643,N_21192,N_18804);
and U28644 (N_28644,N_21808,N_20320);
or U28645 (N_28645,N_19409,N_21227);
nand U28646 (N_28646,N_22333,N_21080);
nand U28647 (N_28647,N_22028,N_18921);
nor U28648 (N_28648,N_21025,N_22875);
and U28649 (N_28649,N_18611,N_19852);
or U28650 (N_28650,N_20709,N_20755);
nand U28651 (N_28651,N_18562,N_18308);
or U28652 (N_28652,N_18506,N_22670);
or U28653 (N_28653,N_23201,N_18873);
nand U28654 (N_28654,N_22132,N_23349);
and U28655 (N_28655,N_21616,N_23856);
nand U28656 (N_28656,N_20686,N_18470);
and U28657 (N_28657,N_23852,N_19637);
nand U28658 (N_28658,N_19846,N_22422);
nor U28659 (N_28659,N_19393,N_23412);
or U28660 (N_28660,N_18470,N_22401);
nor U28661 (N_28661,N_20793,N_18589);
xor U28662 (N_28662,N_18530,N_21353);
nor U28663 (N_28663,N_23772,N_19018);
nor U28664 (N_28664,N_22604,N_19603);
nand U28665 (N_28665,N_18652,N_18995);
xnor U28666 (N_28666,N_18419,N_20163);
nand U28667 (N_28667,N_21653,N_19233);
or U28668 (N_28668,N_21654,N_21631);
nand U28669 (N_28669,N_20216,N_19388);
and U28670 (N_28670,N_20075,N_18879);
xnor U28671 (N_28671,N_22642,N_19337);
nand U28672 (N_28672,N_18339,N_23863);
nand U28673 (N_28673,N_23651,N_20985);
nor U28674 (N_28674,N_20750,N_20903);
or U28675 (N_28675,N_18712,N_21978);
xnor U28676 (N_28676,N_20332,N_22337);
and U28677 (N_28677,N_18584,N_22662);
or U28678 (N_28678,N_18044,N_18012);
xnor U28679 (N_28679,N_21214,N_21479);
nor U28680 (N_28680,N_23454,N_20248);
nor U28681 (N_28681,N_21611,N_22721);
nand U28682 (N_28682,N_20804,N_19614);
or U28683 (N_28683,N_20772,N_20357);
xnor U28684 (N_28684,N_22222,N_22408);
xor U28685 (N_28685,N_20227,N_23631);
nand U28686 (N_28686,N_18974,N_21173);
and U28687 (N_28687,N_23618,N_22378);
or U28688 (N_28688,N_19657,N_20009);
and U28689 (N_28689,N_19953,N_22488);
or U28690 (N_28690,N_23938,N_19574);
nand U28691 (N_28691,N_21037,N_19405);
nand U28692 (N_28692,N_23671,N_23279);
xnor U28693 (N_28693,N_23257,N_22892);
or U28694 (N_28694,N_21896,N_20677);
xor U28695 (N_28695,N_20554,N_19927);
or U28696 (N_28696,N_18797,N_23751);
and U28697 (N_28697,N_22481,N_19709);
xnor U28698 (N_28698,N_21645,N_21237);
xor U28699 (N_28699,N_23870,N_18815);
nor U28700 (N_28700,N_18929,N_20482);
xor U28701 (N_28701,N_21561,N_20103);
and U28702 (N_28702,N_21738,N_23572);
and U28703 (N_28703,N_22243,N_23278);
xnor U28704 (N_28704,N_22979,N_21697);
and U28705 (N_28705,N_18232,N_20385);
nand U28706 (N_28706,N_19673,N_20965);
and U28707 (N_28707,N_19610,N_18950);
xnor U28708 (N_28708,N_23869,N_23909);
nor U28709 (N_28709,N_21468,N_20279);
or U28710 (N_28710,N_21721,N_19870);
and U28711 (N_28711,N_20583,N_21857);
or U28712 (N_28712,N_19414,N_22754);
nand U28713 (N_28713,N_21314,N_23933);
nor U28714 (N_28714,N_20134,N_23976);
nand U28715 (N_28715,N_21273,N_22947);
and U28716 (N_28716,N_21211,N_22067);
nor U28717 (N_28717,N_19890,N_20296);
and U28718 (N_28718,N_23455,N_19273);
nor U28719 (N_28719,N_21394,N_20025);
nand U28720 (N_28720,N_22731,N_22798);
or U28721 (N_28721,N_19645,N_21035);
and U28722 (N_28722,N_20519,N_19516);
xor U28723 (N_28723,N_18220,N_23648);
xor U28724 (N_28724,N_20864,N_19548);
xor U28725 (N_28725,N_23859,N_20014);
and U28726 (N_28726,N_18658,N_19732);
or U28727 (N_28727,N_18425,N_19642);
or U28728 (N_28728,N_22065,N_19771);
nor U28729 (N_28729,N_19728,N_20385);
or U28730 (N_28730,N_23406,N_19127);
or U28731 (N_28731,N_23591,N_21776);
xor U28732 (N_28732,N_22300,N_21840);
nor U28733 (N_28733,N_20947,N_19558);
nor U28734 (N_28734,N_20266,N_22067);
nor U28735 (N_28735,N_19691,N_21248);
nor U28736 (N_28736,N_21147,N_23162);
nand U28737 (N_28737,N_23342,N_22870);
and U28738 (N_28738,N_22818,N_20256);
nand U28739 (N_28739,N_20569,N_18530);
nand U28740 (N_28740,N_18657,N_22918);
xor U28741 (N_28741,N_23045,N_21547);
or U28742 (N_28742,N_19901,N_20832);
nand U28743 (N_28743,N_21470,N_20088);
xor U28744 (N_28744,N_21973,N_21254);
and U28745 (N_28745,N_23605,N_21313);
or U28746 (N_28746,N_18924,N_23807);
or U28747 (N_28747,N_20745,N_18989);
nand U28748 (N_28748,N_21476,N_23253);
nor U28749 (N_28749,N_23478,N_20596);
nor U28750 (N_28750,N_20555,N_21863);
nand U28751 (N_28751,N_22309,N_18207);
xor U28752 (N_28752,N_21460,N_21668);
nand U28753 (N_28753,N_23000,N_20591);
xor U28754 (N_28754,N_23090,N_22238);
and U28755 (N_28755,N_20294,N_18317);
xnor U28756 (N_28756,N_20062,N_22869);
or U28757 (N_28757,N_18155,N_20144);
xnor U28758 (N_28758,N_18518,N_22962);
nand U28759 (N_28759,N_22365,N_21677);
nand U28760 (N_28760,N_19954,N_20666);
or U28761 (N_28761,N_20471,N_20540);
nand U28762 (N_28762,N_20498,N_23413);
and U28763 (N_28763,N_19567,N_21542);
xor U28764 (N_28764,N_23996,N_22230);
nor U28765 (N_28765,N_19981,N_20262);
or U28766 (N_28766,N_19390,N_19142);
nand U28767 (N_28767,N_23569,N_23154);
nand U28768 (N_28768,N_21455,N_18485);
nand U28769 (N_28769,N_23512,N_22695);
or U28770 (N_28770,N_19386,N_23285);
or U28771 (N_28771,N_23810,N_22835);
nor U28772 (N_28772,N_23821,N_19805);
or U28773 (N_28773,N_19019,N_18143);
and U28774 (N_28774,N_20045,N_19446);
nor U28775 (N_28775,N_19292,N_19651);
nand U28776 (N_28776,N_22934,N_19891);
nand U28777 (N_28777,N_22906,N_19254);
nand U28778 (N_28778,N_20227,N_21828);
or U28779 (N_28779,N_18951,N_19563);
or U28780 (N_28780,N_18823,N_21406);
nand U28781 (N_28781,N_18614,N_20226);
or U28782 (N_28782,N_22406,N_18484);
nor U28783 (N_28783,N_19585,N_22258);
nor U28784 (N_28784,N_18741,N_22819);
or U28785 (N_28785,N_19552,N_23820);
and U28786 (N_28786,N_19861,N_22543);
or U28787 (N_28787,N_18567,N_19870);
nor U28788 (N_28788,N_19569,N_23771);
nor U28789 (N_28789,N_21286,N_18655);
nor U28790 (N_28790,N_19460,N_18848);
xnor U28791 (N_28791,N_20949,N_19499);
or U28792 (N_28792,N_19573,N_22091);
nor U28793 (N_28793,N_20645,N_19506);
and U28794 (N_28794,N_20687,N_23215);
nor U28795 (N_28795,N_23987,N_23410);
xor U28796 (N_28796,N_19265,N_23817);
nand U28797 (N_28797,N_23682,N_21362);
or U28798 (N_28798,N_20880,N_20854);
nor U28799 (N_28799,N_23237,N_22997);
nor U28800 (N_28800,N_21250,N_19741);
nand U28801 (N_28801,N_20355,N_23780);
nand U28802 (N_28802,N_18655,N_22653);
nor U28803 (N_28803,N_19125,N_20499);
nor U28804 (N_28804,N_19147,N_23935);
nand U28805 (N_28805,N_22107,N_18415);
nor U28806 (N_28806,N_21235,N_21371);
or U28807 (N_28807,N_20203,N_21075);
nand U28808 (N_28808,N_21633,N_19863);
xnor U28809 (N_28809,N_21335,N_22455);
and U28810 (N_28810,N_23009,N_19765);
nand U28811 (N_28811,N_19843,N_18378);
nand U28812 (N_28812,N_21219,N_23131);
nor U28813 (N_28813,N_19851,N_21065);
nor U28814 (N_28814,N_22732,N_20630);
and U28815 (N_28815,N_23311,N_20872);
nand U28816 (N_28816,N_21800,N_21813);
nor U28817 (N_28817,N_22476,N_18422);
nor U28818 (N_28818,N_18988,N_21617);
nand U28819 (N_28819,N_18034,N_18197);
nor U28820 (N_28820,N_21204,N_18881);
and U28821 (N_28821,N_22750,N_23465);
nand U28822 (N_28822,N_18961,N_19466);
xnor U28823 (N_28823,N_18449,N_23820);
or U28824 (N_28824,N_20979,N_23923);
or U28825 (N_28825,N_18790,N_21798);
xnor U28826 (N_28826,N_23773,N_21066);
and U28827 (N_28827,N_22056,N_21245);
nand U28828 (N_28828,N_22861,N_20144);
xor U28829 (N_28829,N_22983,N_18763);
nand U28830 (N_28830,N_22710,N_23924);
and U28831 (N_28831,N_19786,N_22107);
xor U28832 (N_28832,N_22524,N_18835);
xnor U28833 (N_28833,N_22812,N_22970);
xor U28834 (N_28834,N_22263,N_21592);
and U28835 (N_28835,N_20952,N_22687);
nand U28836 (N_28836,N_21725,N_21184);
or U28837 (N_28837,N_22851,N_20640);
and U28838 (N_28838,N_22838,N_18554);
xor U28839 (N_28839,N_21046,N_18519);
nand U28840 (N_28840,N_23587,N_22690);
nand U28841 (N_28841,N_22024,N_18561);
nand U28842 (N_28842,N_21576,N_18144);
xor U28843 (N_28843,N_23720,N_21159);
and U28844 (N_28844,N_19349,N_20531);
and U28845 (N_28845,N_21279,N_23678);
xor U28846 (N_28846,N_19830,N_20560);
nor U28847 (N_28847,N_22240,N_23843);
nor U28848 (N_28848,N_21556,N_22135);
or U28849 (N_28849,N_18983,N_22805);
xnor U28850 (N_28850,N_19696,N_23853);
nor U28851 (N_28851,N_23038,N_18563);
nand U28852 (N_28852,N_21349,N_18676);
xor U28853 (N_28853,N_23599,N_19765);
nand U28854 (N_28854,N_20403,N_19441);
nand U28855 (N_28855,N_22650,N_18382);
nor U28856 (N_28856,N_22498,N_20467);
or U28857 (N_28857,N_20646,N_20018);
xnor U28858 (N_28858,N_21384,N_23680);
and U28859 (N_28859,N_22523,N_23008);
nor U28860 (N_28860,N_21687,N_19082);
or U28861 (N_28861,N_19938,N_19632);
nand U28862 (N_28862,N_19816,N_21848);
nand U28863 (N_28863,N_18196,N_22890);
nor U28864 (N_28864,N_20538,N_23148);
and U28865 (N_28865,N_19222,N_20969);
nand U28866 (N_28866,N_19395,N_22657);
nand U28867 (N_28867,N_23977,N_19057);
xnor U28868 (N_28868,N_22654,N_23749);
nor U28869 (N_28869,N_18544,N_22264);
nand U28870 (N_28870,N_18200,N_23830);
or U28871 (N_28871,N_22518,N_23051);
or U28872 (N_28872,N_21525,N_22192);
nor U28873 (N_28873,N_22164,N_23644);
or U28874 (N_28874,N_19089,N_20593);
or U28875 (N_28875,N_19494,N_21078);
nor U28876 (N_28876,N_19833,N_20729);
or U28877 (N_28877,N_22786,N_18434);
xor U28878 (N_28878,N_22568,N_18024);
nor U28879 (N_28879,N_22611,N_21981);
nor U28880 (N_28880,N_20706,N_23974);
nand U28881 (N_28881,N_22388,N_19203);
or U28882 (N_28882,N_21847,N_21967);
xor U28883 (N_28883,N_22671,N_23269);
and U28884 (N_28884,N_19513,N_20952);
and U28885 (N_28885,N_21672,N_21398);
nand U28886 (N_28886,N_22571,N_18376);
and U28887 (N_28887,N_19806,N_19274);
nand U28888 (N_28888,N_22451,N_21263);
or U28889 (N_28889,N_20256,N_22022);
and U28890 (N_28890,N_22352,N_19812);
nand U28891 (N_28891,N_20753,N_21325);
nand U28892 (N_28892,N_22529,N_18949);
xnor U28893 (N_28893,N_21842,N_20875);
and U28894 (N_28894,N_23788,N_21010);
or U28895 (N_28895,N_20934,N_19510);
nand U28896 (N_28896,N_20774,N_19427);
nand U28897 (N_28897,N_22855,N_22536);
xor U28898 (N_28898,N_22113,N_22854);
nand U28899 (N_28899,N_20488,N_23802);
or U28900 (N_28900,N_23054,N_21591);
nand U28901 (N_28901,N_20181,N_22683);
and U28902 (N_28902,N_21959,N_20254);
and U28903 (N_28903,N_21227,N_23700);
and U28904 (N_28904,N_23969,N_21498);
nand U28905 (N_28905,N_20593,N_21580);
or U28906 (N_28906,N_18764,N_22003);
and U28907 (N_28907,N_22092,N_20136);
and U28908 (N_28908,N_19840,N_18310);
or U28909 (N_28909,N_23659,N_22354);
xor U28910 (N_28910,N_22146,N_23464);
xor U28911 (N_28911,N_18223,N_18394);
or U28912 (N_28912,N_23930,N_19129);
xor U28913 (N_28913,N_18317,N_21492);
nand U28914 (N_28914,N_20325,N_18927);
nand U28915 (N_28915,N_22713,N_21771);
and U28916 (N_28916,N_23069,N_22839);
and U28917 (N_28917,N_21147,N_20936);
nand U28918 (N_28918,N_23163,N_23159);
and U28919 (N_28919,N_20625,N_19438);
and U28920 (N_28920,N_19529,N_18345);
nand U28921 (N_28921,N_21805,N_23925);
and U28922 (N_28922,N_23968,N_19274);
or U28923 (N_28923,N_18246,N_21896);
or U28924 (N_28924,N_18083,N_20347);
and U28925 (N_28925,N_18425,N_18400);
or U28926 (N_28926,N_18079,N_20973);
nor U28927 (N_28927,N_18459,N_22416);
and U28928 (N_28928,N_21676,N_23200);
or U28929 (N_28929,N_18880,N_23283);
nor U28930 (N_28930,N_20491,N_20580);
or U28931 (N_28931,N_21499,N_22449);
or U28932 (N_28932,N_22844,N_22772);
or U28933 (N_28933,N_22569,N_21836);
nand U28934 (N_28934,N_23530,N_18628);
and U28935 (N_28935,N_19352,N_21745);
nand U28936 (N_28936,N_19561,N_22921);
nand U28937 (N_28937,N_18470,N_22407);
xor U28938 (N_28938,N_19643,N_22730);
and U28939 (N_28939,N_21766,N_23784);
nor U28940 (N_28940,N_18197,N_21736);
or U28941 (N_28941,N_18642,N_23603);
and U28942 (N_28942,N_20244,N_22802);
nand U28943 (N_28943,N_20215,N_19488);
xnor U28944 (N_28944,N_19880,N_18479);
nand U28945 (N_28945,N_22189,N_21148);
or U28946 (N_28946,N_22943,N_19696);
nand U28947 (N_28947,N_19932,N_22667);
xnor U28948 (N_28948,N_22419,N_18334);
and U28949 (N_28949,N_19728,N_19291);
nand U28950 (N_28950,N_21248,N_18454);
and U28951 (N_28951,N_23872,N_23208);
nor U28952 (N_28952,N_21205,N_21235);
nand U28953 (N_28953,N_18026,N_22045);
or U28954 (N_28954,N_19604,N_23996);
or U28955 (N_28955,N_21763,N_23283);
nand U28956 (N_28956,N_22212,N_23961);
xor U28957 (N_28957,N_21926,N_18559);
and U28958 (N_28958,N_22549,N_23725);
nor U28959 (N_28959,N_21606,N_23052);
nand U28960 (N_28960,N_18763,N_23299);
xnor U28961 (N_28961,N_18410,N_18811);
xnor U28962 (N_28962,N_21121,N_18044);
and U28963 (N_28963,N_18910,N_22114);
and U28964 (N_28964,N_19950,N_23261);
nor U28965 (N_28965,N_19774,N_19469);
or U28966 (N_28966,N_23301,N_21563);
nand U28967 (N_28967,N_23744,N_23979);
xor U28968 (N_28968,N_21479,N_22311);
nand U28969 (N_28969,N_23812,N_20685);
and U28970 (N_28970,N_22109,N_20546);
and U28971 (N_28971,N_21153,N_20489);
nand U28972 (N_28972,N_23387,N_19370);
or U28973 (N_28973,N_22866,N_23296);
and U28974 (N_28974,N_18614,N_23230);
xnor U28975 (N_28975,N_20443,N_21764);
nor U28976 (N_28976,N_18733,N_21916);
or U28977 (N_28977,N_20936,N_20925);
or U28978 (N_28978,N_21680,N_20007);
or U28979 (N_28979,N_21566,N_18808);
and U28980 (N_28980,N_20992,N_22800);
or U28981 (N_28981,N_18034,N_19967);
nor U28982 (N_28982,N_18538,N_21370);
and U28983 (N_28983,N_19266,N_19197);
nand U28984 (N_28984,N_22245,N_18665);
or U28985 (N_28985,N_20762,N_23413);
xor U28986 (N_28986,N_18855,N_18509);
and U28987 (N_28987,N_20308,N_20257);
or U28988 (N_28988,N_18818,N_23298);
or U28989 (N_28989,N_19787,N_18559);
nor U28990 (N_28990,N_18217,N_23229);
xor U28991 (N_28991,N_21840,N_19308);
and U28992 (N_28992,N_18679,N_19828);
xor U28993 (N_28993,N_22468,N_21829);
nand U28994 (N_28994,N_21203,N_19444);
or U28995 (N_28995,N_23645,N_22863);
or U28996 (N_28996,N_21661,N_22770);
or U28997 (N_28997,N_18233,N_18771);
nand U28998 (N_28998,N_19077,N_18291);
xor U28999 (N_28999,N_22385,N_22593);
xnor U29000 (N_29000,N_23266,N_22925);
xnor U29001 (N_29001,N_22110,N_23112);
nand U29002 (N_29002,N_23917,N_18321);
or U29003 (N_29003,N_23862,N_20756);
xnor U29004 (N_29004,N_20452,N_18451);
and U29005 (N_29005,N_20966,N_19320);
xor U29006 (N_29006,N_21944,N_23268);
nand U29007 (N_29007,N_21267,N_19518);
nand U29008 (N_29008,N_21041,N_20444);
nor U29009 (N_29009,N_19670,N_21564);
nand U29010 (N_29010,N_20419,N_20223);
and U29011 (N_29011,N_20365,N_22953);
or U29012 (N_29012,N_22133,N_18332);
xnor U29013 (N_29013,N_20812,N_20202);
nand U29014 (N_29014,N_19252,N_22035);
and U29015 (N_29015,N_20114,N_22540);
nand U29016 (N_29016,N_22137,N_19548);
or U29017 (N_29017,N_22724,N_20988);
and U29018 (N_29018,N_18042,N_19980);
nor U29019 (N_29019,N_21005,N_20466);
and U29020 (N_29020,N_23609,N_23305);
nor U29021 (N_29021,N_18593,N_22002);
nand U29022 (N_29022,N_21973,N_18286);
or U29023 (N_29023,N_21216,N_21172);
or U29024 (N_29024,N_23464,N_19708);
nand U29025 (N_29025,N_21379,N_22252);
nand U29026 (N_29026,N_18515,N_21452);
xor U29027 (N_29027,N_22716,N_22192);
nor U29028 (N_29028,N_21289,N_19726);
xnor U29029 (N_29029,N_22749,N_18545);
or U29030 (N_29030,N_20685,N_21865);
xnor U29031 (N_29031,N_23215,N_22885);
nor U29032 (N_29032,N_23324,N_22679);
and U29033 (N_29033,N_22148,N_20386);
or U29034 (N_29034,N_19041,N_23656);
nand U29035 (N_29035,N_19419,N_21871);
nor U29036 (N_29036,N_23193,N_20048);
or U29037 (N_29037,N_21189,N_23564);
and U29038 (N_29038,N_23371,N_22257);
nor U29039 (N_29039,N_19229,N_18508);
nor U29040 (N_29040,N_21542,N_22675);
and U29041 (N_29041,N_23915,N_21181);
xnor U29042 (N_29042,N_21686,N_18725);
xor U29043 (N_29043,N_20817,N_19695);
nor U29044 (N_29044,N_19810,N_18392);
and U29045 (N_29045,N_20184,N_21262);
nor U29046 (N_29046,N_20743,N_18919);
xor U29047 (N_29047,N_20442,N_23888);
nor U29048 (N_29048,N_21823,N_20282);
nor U29049 (N_29049,N_20174,N_20797);
nor U29050 (N_29050,N_22014,N_20021);
xnor U29051 (N_29051,N_22566,N_19667);
nand U29052 (N_29052,N_22240,N_20261);
xor U29053 (N_29053,N_22071,N_22358);
or U29054 (N_29054,N_20981,N_18113);
xor U29055 (N_29055,N_18053,N_22180);
nor U29056 (N_29056,N_21540,N_19919);
and U29057 (N_29057,N_19973,N_23141);
and U29058 (N_29058,N_21356,N_18476);
or U29059 (N_29059,N_21614,N_19355);
nand U29060 (N_29060,N_19726,N_19428);
xor U29061 (N_29061,N_23437,N_22119);
nand U29062 (N_29062,N_21135,N_23070);
nor U29063 (N_29063,N_23614,N_19269);
nand U29064 (N_29064,N_22380,N_21222);
or U29065 (N_29065,N_20381,N_20514);
nand U29066 (N_29066,N_18222,N_19736);
nand U29067 (N_29067,N_21897,N_23860);
nand U29068 (N_29068,N_23807,N_20084);
or U29069 (N_29069,N_18830,N_19345);
nor U29070 (N_29070,N_21743,N_20224);
xor U29071 (N_29071,N_22587,N_19442);
nor U29072 (N_29072,N_22072,N_18632);
or U29073 (N_29073,N_20773,N_20327);
nand U29074 (N_29074,N_22842,N_21882);
nor U29075 (N_29075,N_23369,N_22942);
xnor U29076 (N_29076,N_18052,N_21964);
or U29077 (N_29077,N_20757,N_23940);
xnor U29078 (N_29078,N_20249,N_19829);
nor U29079 (N_29079,N_20457,N_22537);
nor U29080 (N_29080,N_18081,N_22281);
nand U29081 (N_29081,N_19384,N_19228);
nor U29082 (N_29082,N_20876,N_23097);
nor U29083 (N_29083,N_20264,N_22064);
nor U29084 (N_29084,N_18104,N_20121);
or U29085 (N_29085,N_23867,N_22849);
nand U29086 (N_29086,N_22804,N_18451);
or U29087 (N_29087,N_23992,N_22070);
or U29088 (N_29088,N_23829,N_20988);
and U29089 (N_29089,N_18469,N_23095);
and U29090 (N_29090,N_21753,N_20961);
or U29091 (N_29091,N_19187,N_23362);
nand U29092 (N_29092,N_19187,N_23708);
or U29093 (N_29093,N_19622,N_23669);
xor U29094 (N_29094,N_19787,N_20316);
xor U29095 (N_29095,N_23170,N_20371);
and U29096 (N_29096,N_20592,N_19518);
nand U29097 (N_29097,N_22883,N_22128);
nor U29098 (N_29098,N_19584,N_21744);
and U29099 (N_29099,N_18651,N_19664);
nand U29100 (N_29100,N_23409,N_19931);
nand U29101 (N_29101,N_22480,N_18744);
nand U29102 (N_29102,N_18050,N_20234);
xnor U29103 (N_29103,N_21388,N_20761);
xnor U29104 (N_29104,N_22099,N_23968);
xnor U29105 (N_29105,N_21925,N_18680);
and U29106 (N_29106,N_21792,N_19051);
or U29107 (N_29107,N_21017,N_21972);
or U29108 (N_29108,N_18876,N_19522);
or U29109 (N_29109,N_21087,N_20369);
and U29110 (N_29110,N_22076,N_22567);
or U29111 (N_29111,N_21554,N_21047);
xnor U29112 (N_29112,N_19803,N_22421);
nand U29113 (N_29113,N_23548,N_23750);
and U29114 (N_29114,N_23667,N_23650);
or U29115 (N_29115,N_22739,N_18562);
nand U29116 (N_29116,N_22037,N_22080);
nor U29117 (N_29117,N_21927,N_23479);
or U29118 (N_29118,N_20377,N_23336);
nor U29119 (N_29119,N_22275,N_20154);
nand U29120 (N_29120,N_19010,N_23776);
nor U29121 (N_29121,N_21974,N_22836);
xor U29122 (N_29122,N_18391,N_22254);
and U29123 (N_29123,N_18041,N_23357);
nor U29124 (N_29124,N_19500,N_20740);
nand U29125 (N_29125,N_18297,N_21449);
or U29126 (N_29126,N_22066,N_18472);
xor U29127 (N_29127,N_23916,N_21617);
and U29128 (N_29128,N_21921,N_19394);
or U29129 (N_29129,N_22652,N_18842);
and U29130 (N_29130,N_21484,N_19862);
nor U29131 (N_29131,N_20734,N_22958);
xnor U29132 (N_29132,N_23011,N_19579);
xnor U29133 (N_29133,N_19295,N_21115);
nand U29134 (N_29134,N_20658,N_21150);
and U29135 (N_29135,N_22092,N_20878);
nor U29136 (N_29136,N_20756,N_18625);
nor U29137 (N_29137,N_21156,N_21782);
xnor U29138 (N_29138,N_22156,N_18424);
xor U29139 (N_29139,N_18240,N_23396);
xor U29140 (N_29140,N_22296,N_20018);
or U29141 (N_29141,N_22824,N_23530);
or U29142 (N_29142,N_22292,N_23369);
or U29143 (N_29143,N_21284,N_23090);
xor U29144 (N_29144,N_23552,N_22864);
xnor U29145 (N_29145,N_22481,N_19279);
xor U29146 (N_29146,N_18989,N_18908);
and U29147 (N_29147,N_18382,N_19766);
and U29148 (N_29148,N_18512,N_22450);
nand U29149 (N_29149,N_20398,N_20941);
nor U29150 (N_29150,N_18167,N_23765);
and U29151 (N_29151,N_23229,N_22656);
or U29152 (N_29152,N_18215,N_21093);
nor U29153 (N_29153,N_20041,N_23774);
nand U29154 (N_29154,N_18349,N_18129);
or U29155 (N_29155,N_19542,N_21085);
nor U29156 (N_29156,N_23529,N_22995);
nor U29157 (N_29157,N_19973,N_18039);
or U29158 (N_29158,N_18343,N_18317);
xor U29159 (N_29159,N_22212,N_22845);
xnor U29160 (N_29160,N_20542,N_23024);
xor U29161 (N_29161,N_21123,N_20441);
nand U29162 (N_29162,N_23397,N_18892);
nand U29163 (N_29163,N_18772,N_23883);
nor U29164 (N_29164,N_20583,N_23913);
nand U29165 (N_29165,N_18882,N_23142);
xnor U29166 (N_29166,N_18348,N_20760);
xnor U29167 (N_29167,N_20591,N_21214);
nand U29168 (N_29168,N_21332,N_20919);
nor U29169 (N_29169,N_18758,N_19129);
nor U29170 (N_29170,N_21842,N_20470);
nor U29171 (N_29171,N_23774,N_21687);
nor U29172 (N_29172,N_22219,N_20454);
or U29173 (N_29173,N_20379,N_19454);
nand U29174 (N_29174,N_18874,N_18494);
nor U29175 (N_29175,N_22982,N_20794);
and U29176 (N_29176,N_23745,N_18042);
nor U29177 (N_29177,N_20110,N_19730);
xor U29178 (N_29178,N_23486,N_23264);
or U29179 (N_29179,N_19721,N_21851);
or U29180 (N_29180,N_22354,N_23266);
nor U29181 (N_29181,N_20792,N_21995);
or U29182 (N_29182,N_19471,N_19303);
or U29183 (N_29183,N_20579,N_20138);
nand U29184 (N_29184,N_18431,N_19524);
and U29185 (N_29185,N_19353,N_23928);
and U29186 (N_29186,N_19144,N_20910);
nand U29187 (N_29187,N_18427,N_23076);
or U29188 (N_29188,N_21934,N_23044);
nor U29189 (N_29189,N_18247,N_20153);
or U29190 (N_29190,N_18851,N_19832);
or U29191 (N_29191,N_21496,N_20697);
nor U29192 (N_29192,N_21614,N_20125);
or U29193 (N_29193,N_21381,N_19289);
nor U29194 (N_29194,N_18701,N_19353);
xor U29195 (N_29195,N_23835,N_21144);
xor U29196 (N_29196,N_18631,N_18214);
nor U29197 (N_29197,N_23778,N_18558);
nor U29198 (N_29198,N_20508,N_19641);
or U29199 (N_29199,N_22597,N_23604);
xnor U29200 (N_29200,N_20858,N_20726);
and U29201 (N_29201,N_21005,N_22888);
xnor U29202 (N_29202,N_21461,N_21107);
and U29203 (N_29203,N_18008,N_22995);
nand U29204 (N_29204,N_22336,N_21196);
and U29205 (N_29205,N_23337,N_18766);
or U29206 (N_29206,N_21598,N_23367);
nor U29207 (N_29207,N_23844,N_22733);
and U29208 (N_29208,N_18815,N_18486);
nor U29209 (N_29209,N_22421,N_19181);
nor U29210 (N_29210,N_20047,N_19265);
and U29211 (N_29211,N_18769,N_21124);
nand U29212 (N_29212,N_21796,N_19200);
or U29213 (N_29213,N_19546,N_19708);
nor U29214 (N_29214,N_23683,N_21334);
and U29215 (N_29215,N_20067,N_20049);
or U29216 (N_29216,N_22515,N_21519);
and U29217 (N_29217,N_23974,N_22124);
nor U29218 (N_29218,N_18614,N_21723);
nand U29219 (N_29219,N_23551,N_23800);
and U29220 (N_29220,N_21079,N_19733);
nand U29221 (N_29221,N_19025,N_22610);
xnor U29222 (N_29222,N_19134,N_21624);
and U29223 (N_29223,N_22049,N_23523);
nor U29224 (N_29224,N_18916,N_21570);
xor U29225 (N_29225,N_21644,N_19876);
nor U29226 (N_29226,N_18021,N_20021);
or U29227 (N_29227,N_22317,N_21317);
xnor U29228 (N_29228,N_20544,N_23748);
nand U29229 (N_29229,N_20904,N_19221);
xor U29230 (N_29230,N_19661,N_18879);
and U29231 (N_29231,N_20202,N_22422);
nand U29232 (N_29232,N_23475,N_23292);
or U29233 (N_29233,N_20841,N_18104);
or U29234 (N_29234,N_19370,N_19276);
and U29235 (N_29235,N_23933,N_23011);
xnor U29236 (N_29236,N_22040,N_18114);
nand U29237 (N_29237,N_18526,N_22379);
or U29238 (N_29238,N_23325,N_19132);
nand U29239 (N_29239,N_21540,N_20076);
nand U29240 (N_29240,N_22192,N_20515);
nor U29241 (N_29241,N_23396,N_18157);
and U29242 (N_29242,N_19507,N_18266);
xnor U29243 (N_29243,N_20678,N_21632);
xnor U29244 (N_29244,N_22763,N_23051);
and U29245 (N_29245,N_21124,N_20803);
and U29246 (N_29246,N_23078,N_23322);
xnor U29247 (N_29247,N_22173,N_20649);
xnor U29248 (N_29248,N_20731,N_22692);
nand U29249 (N_29249,N_19755,N_19316);
xnor U29250 (N_29250,N_21769,N_23217);
or U29251 (N_29251,N_23708,N_18739);
nand U29252 (N_29252,N_20021,N_23165);
nand U29253 (N_29253,N_19839,N_18443);
or U29254 (N_29254,N_23345,N_23283);
nand U29255 (N_29255,N_21101,N_19318);
and U29256 (N_29256,N_18913,N_19561);
nand U29257 (N_29257,N_20576,N_23230);
and U29258 (N_29258,N_18418,N_22095);
and U29259 (N_29259,N_20314,N_22631);
nand U29260 (N_29260,N_19016,N_18104);
or U29261 (N_29261,N_23878,N_22720);
nor U29262 (N_29262,N_19584,N_19733);
or U29263 (N_29263,N_21588,N_21245);
nor U29264 (N_29264,N_23388,N_19002);
nor U29265 (N_29265,N_19390,N_20156);
and U29266 (N_29266,N_19557,N_23890);
nand U29267 (N_29267,N_19177,N_23474);
or U29268 (N_29268,N_23221,N_19269);
and U29269 (N_29269,N_18065,N_18792);
nand U29270 (N_29270,N_20784,N_20040);
nand U29271 (N_29271,N_22096,N_19196);
or U29272 (N_29272,N_20527,N_22130);
xor U29273 (N_29273,N_20983,N_21323);
xor U29274 (N_29274,N_18842,N_22482);
nand U29275 (N_29275,N_19056,N_21115);
or U29276 (N_29276,N_18588,N_20072);
or U29277 (N_29277,N_22228,N_19113);
or U29278 (N_29278,N_20131,N_21279);
nand U29279 (N_29279,N_19225,N_21327);
nand U29280 (N_29280,N_20427,N_23848);
or U29281 (N_29281,N_21058,N_19489);
nor U29282 (N_29282,N_21710,N_19294);
or U29283 (N_29283,N_21121,N_18998);
xor U29284 (N_29284,N_20420,N_18012);
nor U29285 (N_29285,N_23560,N_21170);
xor U29286 (N_29286,N_21190,N_20035);
and U29287 (N_29287,N_19437,N_22534);
or U29288 (N_29288,N_18174,N_22548);
nor U29289 (N_29289,N_19266,N_22954);
and U29290 (N_29290,N_18612,N_19666);
nand U29291 (N_29291,N_18593,N_20367);
xnor U29292 (N_29292,N_22068,N_20609);
nor U29293 (N_29293,N_20517,N_21686);
or U29294 (N_29294,N_22957,N_18197);
or U29295 (N_29295,N_23945,N_18003);
nand U29296 (N_29296,N_21063,N_21924);
xor U29297 (N_29297,N_23569,N_19366);
xnor U29298 (N_29298,N_20769,N_23416);
or U29299 (N_29299,N_18915,N_18277);
or U29300 (N_29300,N_23866,N_23567);
and U29301 (N_29301,N_18720,N_18946);
nor U29302 (N_29302,N_19217,N_22225);
xor U29303 (N_29303,N_19813,N_19037);
or U29304 (N_29304,N_20766,N_19970);
and U29305 (N_29305,N_18003,N_19567);
nor U29306 (N_29306,N_23870,N_21139);
nor U29307 (N_29307,N_21859,N_19513);
nand U29308 (N_29308,N_19916,N_22762);
and U29309 (N_29309,N_20973,N_23498);
or U29310 (N_29310,N_18601,N_19103);
xnor U29311 (N_29311,N_19477,N_23774);
nand U29312 (N_29312,N_21777,N_22814);
xnor U29313 (N_29313,N_21777,N_21706);
or U29314 (N_29314,N_19696,N_23696);
nand U29315 (N_29315,N_21929,N_23588);
xnor U29316 (N_29316,N_21532,N_23165);
or U29317 (N_29317,N_22139,N_21932);
xor U29318 (N_29318,N_22500,N_18505);
and U29319 (N_29319,N_18784,N_23633);
and U29320 (N_29320,N_19203,N_23196);
nor U29321 (N_29321,N_20370,N_21061);
and U29322 (N_29322,N_23477,N_22621);
and U29323 (N_29323,N_20834,N_22336);
nor U29324 (N_29324,N_21622,N_18024);
and U29325 (N_29325,N_23932,N_19275);
and U29326 (N_29326,N_19868,N_20817);
and U29327 (N_29327,N_18240,N_18564);
nand U29328 (N_29328,N_22799,N_21263);
xnor U29329 (N_29329,N_22009,N_22978);
nor U29330 (N_29330,N_18059,N_20994);
and U29331 (N_29331,N_22578,N_20339);
xnor U29332 (N_29332,N_22389,N_22238);
xor U29333 (N_29333,N_23551,N_21263);
or U29334 (N_29334,N_20403,N_22828);
nand U29335 (N_29335,N_23839,N_21558);
nor U29336 (N_29336,N_20174,N_23585);
or U29337 (N_29337,N_20509,N_18635);
nor U29338 (N_29338,N_20544,N_22887);
nor U29339 (N_29339,N_20037,N_18531);
and U29340 (N_29340,N_18049,N_19902);
nor U29341 (N_29341,N_21527,N_22050);
and U29342 (N_29342,N_18695,N_18297);
nor U29343 (N_29343,N_21761,N_23909);
or U29344 (N_29344,N_19893,N_20124);
nand U29345 (N_29345,N_18209,N_21996);
and U29346 (N_29346,N_19553,N_22781);
nand U29347 (N_29347,N_19210,N_20981);
xor U29348 (N_29348,N_23918,N_18668);
or U29349 (N_29349,N_23963,N_22417);
or U29350 (N_29350,N_21453,N_23780);
or U29351 (N_29351,N_23663,N_22345);
nand U29352 (N_29352,N_23639,N_23892);
and U29353 (N_29353,N_18032,N_20736);
xor U29354 (N_29354,N_21335,N_22815);
xnor U29355 (N_29355,N_19209,N_22562);
nand U29356 (N_29356,N_22866,N_21353);
nand U29357 (N_29357,N_21618,N_19153);
nand U29358 (N_29358,N_21772,N_23819);
nand U29359 (N_29359,N_22284,N_21996);
nor U29360 (N_29360,N_19208,N_23590);
nor U29361 (N_29361,N_20616,N_23264);
xnor U29362 (N_29362,N_18341,N_20148);
nand U29363 (N_29363,N_18619,N_22493);
nand U29364 (N_29364,N_21855,N_22271);
nor U29365 (N_29365,N_20748,N_19399);
nor U29366 (N_29366,N_22348,N_18670);
or U29367 (N_29367,N_22360,N_18408);
xor U29368 (N_29368,N_23418,N_21874);
and U29369 (N_29369,N_20894,N_21526);
xnor U29370 (N_29370,N_21167,N_22043);
xor U29371 (N_29371,N_18850,N_23511);
nand U29372 (N_29372,N_23573,N_21713);
nand U29373 (N_29373,N_22481,N_23743);
and U29374 (N_29374,N_20682,N_22662);
and U29375 (N_29375,N_22488,N_20934);
nor U29376 (N_29376,N_21289,N_20267);
nor U29377 (N_29377,N_18456,N_21571);
and U29378 (N_29378,N_22238,N_21101);
nand U29379 (N_29379,N_23441,N_22853);
or U29380 (N_29380,N_19810,N_21868);
nand U29381 (N_29381,N_20440,N_22952);
xnor U29382 (N_29382,N_20725,N_20763);
nand U29383 (N_29383,N_18929,N_20677);
nor U29384 (N_29384,N_19900,N_19682);
and U29385 (N_29385,N_19195,N_23702);
and U29386 (N_29386,N_22223,N_19359);
nor U29387 (N_29387,N_22361,N_22726);
and U29388 (N_29388,N_22523,N_22920);
and U29389 (N_29389,N_23721,N_22384);
xor U29390 (N_29390,N_19567,N_22192);
or U29391 (N_29391,N_18104,N_22422);
nor U29392 (N_29392,N_19140,N_21752);
nand U29393 (N_29393,N_21172,N_23600);
or U29394 (N_29394,N_23659,N_22054);
xnor U29395 (N_29395,N_21283,N_18199);
and U29396 (N_29396,N_19595,N_23665);
nand U29397 (N_29397,N_21158,N_18600);
nand U29398 (N_29398,N_22015,N_19378);
or U29399 (N_29399,N_20830,N_18145);
nand U29400 (N_29400,N_22068,N_19478);
nor U29401 (N_29401,N_20147,N_18823);
xnor U29402 (N_29402,N_23502,N_22454);
nand U29403 (N_29403,N_21426,N_18136);
nand U29404 (N_29404,N_20680,N_21898);
and U29405 (N_29405,N_20114,N_18734);
nand U29406 (N_29406,N_18990,N_23011);
nand U29407 (N_29407,N_23138,N_19572);
xnor U29408 (N_29408,N_21302,N_19852);
nor U29409 (N_29409,N_19279,N_18447);
and U29410 (N_29410,N_18678,N_18738);
or U29411 (N_29411,N_19339,N_22111);
nand U29412 (N_29412,N_19663,N_23400);
xor U29413 (N_29413,N_21192,N_18784);
nor U29414 (N_29414,N_21030,N_23448);
or U29415 (N_29415,N_19145,N_20448);
xor U29416 (N_29416,N_19064,N_23340);
nand U29417 (N_29417,N_22064,N_22460);
nand U29418 (N_29418,N_20685,N_22695);
xnor U29419 (N_29419,N_18394,N_18323);
nor U29420 (N_29420,N_22463,N_19674);
nand U29421 (N_29421,N_21152,N_21703);
and U29422 (N_29422,N_19950,N_18760);
nand U29423 (N_29423,N_19972,N_23147);
and U29424 (N_29424,N_22495,N_21992);
xnor U29425 (N_29425,N_23049,N_19299);
nand U29426 (N_29426,N_18018,N_21713);
nor U29427 (N_29427,N_23830,N_19222);
nand U29428 (N_29428,N_22852,N_22448);
nand U29429 (N_29429,N_23357,N_23683);
nand U29430 (N_29430,N_23174,N_18821);
nand U29431 (N_29431,N_23815,N_21243);
nand U29432 (N_29432,N_21280,N_20568);
nor U29433 (N_29433,N_18833,N_18385);
nand U29434 (N_29434,N_19549,N_19434);
nand U29435 (N_29435,N_19533,N_23031);
or U29436 (N_29436,N_21317,N_19690);
and U29437 (N_29437,N_22796,N_22151);
nand U29438 (N_29438,N_18749,N_23302);
xnor U29439 (N_29439,N_22833,N_23608);
nor U29440 (N_29440,N_23383,N_20133);
xor U29441 (N_29441,N_19282,N_21272);
nor U29442 (N_29442,N_23541,N_23374);
xnor U29443 (N_29443,N_23246,N_23253);
or U29444 (N_29444,N_19659,N_21111);
or U29445 (N_29445,N_19058,N_18074);
xor U29446 (N_29446,N_20035,N_20691);
and U29447 (N_29447,N_22426,N_18101);
nor U29448 (N_29448,N_23121,N_23626);
nor U29449 (N_29449,N_18998,N_19178);
or U29450 (N_29450,N_19921,N_23620);
or U29451 (N_29451,N_23577,N_22253);
nand U29452 (N_29452,N_22914,N_22526);
and U29453 (N_29453,N_20014,N_22512);
or U29454 (N_29454,N_20851,N_19620);
nand U29455 (N_29455,N_21734,N_18478);
xnor U29456 (N_29456,N_20342,N_18105);
nor U29457 (N_29457,N_18714,N_20833);
and U29458 (N_29458,N_22775,N_20270);
nor U29459 (N_29459,N_22759,N_18033);
nand U29460 (N_29460,N_19452,N_23340);
or U29461 (N_29461,N_21421,N_21459);
or U29462 (N_29462,N_20601,N_19509);
nor U29463 (N_29463,N_22219,N_23782);
and U29464 (N_29464,N_19278,N_19151);
nand U29465 (N_29465,N_21207,N_20098);
nor U29466 (N_29466,N_19927,N_19845);
or U29467 (N_29467,N_18705,N_20747);
nor U29468 (N_29468,N_23152,N_19802);
xor U29469 (N_29469,N_21492,N_21101);
nand U29470 (N_29470,N_23082,N_21613);
nor U29471 (N_29471,N_20526,N_21224);
and U29472 (N_29472,N_23455,N_19916);
and U29473 (N_29473,N_20202,N_19271);
or U29474 (N_29474,N_23905,N_22585);
xor U29475 (N_29475,N_21867,N_21641);
nand U29476 (N_29476,N_18980,N_23326);
and U29477 (N_29477,N_23298,N_19966);
nand U29478 (N_29478,N_18568,N_22758);
xnor U29479 (N_29479,N_19750,N_22706);
or U29480 (N_29480,N_21297,N_18424);
nand U29481 (N_29481,N_22310,N_23995);
or U29482 (N_29482,N_20976,N_22654);
and U29483 (N_29483,N_18668,N_19927);
xor U29484 (N_29484,N_21921,N_18136);
and U29485 (N_29485,N_20288,N_20240);
or U29486 (N_29486,N_18328,N_19478);
or U29487 (N_29487,N_21037,N_21507);
nand U29488 (N_29488,N_19965,N_20008);
nor U29489 (N_29489,N_23855,N_20653);
nand U29490 (N_29490,N_21411,N_19882);
nor U29491 (N_29491,N_22259,N_23855);
and U29492 (N_29492,N_21269,N_23849);
nor U29493 (N_29493,N_22276,N_21069);
nand U29494 (N_29494,N_22468,N_20330);
and U29495 (N_29495,N_18026,N_19230);
xnor U29496 (N_29496,N_20852,N_21965);
nand U29497 (N_29497,N_21470,N_19467);
and U29498 (N_29498,N_22348,N_23209);
xnor U29499 (N_29499,N_23262,N_23130);
or U29500 (N_29500,N_18591,N_22059);
xor U29501 (N_29501,N_22165,N_18146);
xor U29502 (N_29502,N_18520,N_20803);
and U29503 (N_29503,N_22008,N_22879);
xor U29504 (N_29504,N_23843,N_20083);
nand U29505 (N_29505,N_23936,N_19734);
nand U29506 (N_29506,N_18100,N_21597);
nor U29507 (N_29507,N_23228,N_20334);
or U29508 (N_29508,N_23626,N_20889);
and U29509 (N_29509,N_22851,N_22039);
and U29510 (N_29510,N_18603,N_20748);
and U29511 (N_29511,N_22028,N_19290);
nor U29512 (N_29512,N_19353,N_22572);
nor U29513 (N_29513,N_18438,N_20941);
nor U29514 (N_29514,N_21678,N_21733);
and U29515 (N_29515,N_22776,N_23411);
nor U29516 (N_29516,N_19168,N_19163);
xor U29517 (N_29517,N_20535,N_22428);
xor U29518 (N_29518,N_18430,N_18414);
xor U29519 (N_29519,N_19742,N_23433);
or U29520 (N_29520,N_22193,N_18946);
or U29521 (N_29521,N_21588,N_20160);
nor U29522 (N_29522,N_22152,N_22742);
nor U29523 (N_29523,N_19688,N_21016);
nand U29524 (N_29524,N_18279,N_23354);
xnor U29525 (N_29525,N_21199,N_21885);
or U29526 (N_29526,N_23426,N_18576);
or U29527 (N_29527,N_18305,N_23545);
xnor U29528 (N_29528,N_18926,N_23638);
or U29529 (N_29529,N_19345,N_19061);
or U29530 (N_29530,N_19813,N_21088);
or U29531 (N_29531,N_23463,N_23805);
xor U29532 (N_29532,N_21390,N_18842);
or U29533 (N_29533,N_21250,N_21817);
and U29534 (N_29534,N_23823,N_23392);
and U29535 (N_29535,N_18670,N_19103);
nor U29536 (N_29536,N_21394,N_20300);
and U29537 (N_29537,N_20488,N_18572);
xor U29538 (N_29538,N_22542,N_22591);
or U29539 (N_29539,N_18314,N_18966);
nor U29540 (N_29540,N_22793,N_22293);
nand U29541 (N_29541,N_19968,N_23514);
nor U29542 (N_29542,N_21966,N_19063);
xnor U29543 (N_29543,N_23198,N_19137);
or U29544 (N_29544,N_18883,N_18194);
xor U29545 (N_29545,N_18316,N_22566);
or U29546 (N_29546,N_19336,N_23498);
or U29547 (N_29547,N_23485,N_21614);
nand U29548 (N_29548,N_21225,N_18179);
xnor U29549 (N_29549,N_20755,N_20838);
nand U29550 (N_29550,N_21527,N_20635);
nor U29551 (N_29551,N_18774,N_21727);
or U29552 (N_29552,N_20537,N_19075);
nor U29553 (N_29553,N_21424,N_18616);
nor U29554 (N_29554,N_21238,N_22901);
nor U29555 (N_29555,N_19675,N_21434);
nand U29556 (N_29556,N_21517,N_23350);
nor U29557 (N_29557,N_18788,N_20744);
xor U29558 (N_29558,N_18417,N_19789);
nor U29559 (N_29559,N_22654,N_19004);
and U29560 (N_29560,N_21893,N_20949);
or U29561 (N_29561,N_19585,N_22242);
xnor U29562 (N_29562,N_23758,N_18724);
xnor U29563 (N_29563,N_18038,N_19690);
nand U29564 (N_29564,N_18591,N_19973);
and U29565 (N_29565,N_18426,N_18538);
nand U29566 (N_29566,N_23316,N_19959);
or U29567 (N_29567,N_18409,N_22577);
nor U29568 (N_29568,N_19482,N_23509);
nand U29569 (N_29569,N_20030,N_22151);
nand U29570 (N_29570,N_21317,N_18724);
nand U29571 (N_29571,N_21704,N_18250);
xor U29572 (N_29572,N_21934,N_21451);
nor U29573 (N_29573,N_18292,N_22724);
or U29574 (N_29574,N_18925,N_18869);
nand U29575 (N_29575,N_21471,N_20206);
nand U29576 (N_29576,N_19747,N_23247);
nand U29577 (N_29577,N_20971,N_18357);
nor U29578 (N_29578,N_20413,N_21444);
nand U29579 (N_29579,N_20701,N_21093);
nor U29580 (N_29580,N_20328,N_23445);
xor U29581 (N_29581,N_23036,N_19261);
and U29582 (N_29582,N_20526,N_18741);
nor U29583 (N_29583,N_18332,N_18183);
nand U29584 (N_29584,N_18870,N_21239);
and U29585 (N_29585,N_23990,N_21271);
nor U29586 (N_29586,N_22851,N_22779);
and U29587 (N_29587,N_19099,N_20966);
or U29588 (N_29588,N_19289,N_19572);
or U29589 (N_29589,N_22001,N_20617);
xor U29590 (N_29590,N_22609,N_23145);
xor U29591 (N_29591,N_22769,N_21443);
or U29592 (N_29592,N_18853,N_19638);
or U29593 (N_29593,N_22670,N_18778);
nand U29594 (N_29594,N_20759,N_18914);
nor U29595 (N_29595,N_20344,N_19476);
or U29596 (N_29596,N_20895,N_19481);
and U29597 (N_29597,N_21072,N_23900);
nand U29598 (N_29598,N_20907,N_23310);
xnor U29599 (N_29599,N_20946,N_19092);
xor U29600 (N_29600,N_23531,N_21204);
and U29601 (N_29601,N_21726,N_23233);
or U29602 (N_29602,N_19381,N_19443);
nor U29603 (N_29603,N_20640,N_21848);
and U29604 (N_29604,N_21963,N_20182);
nand U29605 (N_29605,N_21265,N_20108);
or U29606 (N_29606,N_21560,N_20435);
nand U29607 (N_29607,N_18975,N_19993);
nor U29608 (N_29608,N_20845,N_20256);
nor U29609 (N_29609,N_21444,N_21171);
nor U29610 (N_29610,N_18942,N_20746);
or U29611 (N_29611,N_21138,N_20238);
nor U29612 (N_29612,N_23335,N_23823);
and U29613 (N_29613,N_22756,N_18052);
or U29614 (N_29614,N_23575,N_22979);
or U29615 (N_29615,N_18247,N_22521);
or U29616 (N_29616,N_22750,N_23410);
nor U29617 (N_29617,N_20063,N_23913);
nor U29618 (N_29618,N_22005,N_20141);
xor U29619 (N_29619,N_23817,N_23807);
or U29620 (N_29620,N_22320,N_19171);
nor U29621 (N_29621,N_19658,N_22622);
and U29622 (N_29622,N_23169,N_19797);
xnor U29623 (N_29623,N_21343,N_19707);
nor U29624 (N_29624,N_23173,N_21071);
and U29625 (N_29625,N_20302,N_21016);
xor U29626 (N_29626,N_22862,N_23225);
or U29627 (N_29627,N_23165,N_22736);
nor U29628 (N_29628,N_18346,N_20388);
and U29629 (N_29629,N_21739,N_20627);
xnor U29630 (N_29630,N_18222,N_22365);
or U29631 (N_29631,N_20503,N_22067);
nand U29632 (N_29632,N_22253,N_19040);
nand U29633 (N_29633,N_21864,N_19875);
or U29634 (N_29634,N_22561,N_23921);
nor U29635 (N_29635,N_22006,N_20655);
and U29636 (N_29636,N_22047,N_23408);
nand U29637 (N_29637,N_23232,N_19585);
nand U29638 (N_29638,N_23199,N_23715);
nor U29639 (N_29639,N_20601,N_20123);
and U29640 (N_29640,N_20580,N_20237);
xor U29641 (N_29641,N_18597,N_18676);
or U29642 (N_29642,N_22847,N_20749);
xor U29643 (N_29643,N_20245,N_23719);
nand U29644 (N_29644,N_22078,N_18436);
xnor U29645 (N_29645,N_20505,N_18243);
nor U29646 (N_29646,N_22221,N_23527);
nand U29647 (N_29647,N_22278,N_18608);
nand U29648 (N_29648,N_23007,N_23239);
and U29649 (N_29649,N_18549,N_19193);
and U29650 (N_29650,N_19835,N_19607);
or U29651 (N_29651,N_23913,N_20527);
xor U29652 (N_29652,N_23681,N_23254);
nor U29653 (N_29653,N_20036,N_21148);
or U29654 (N_29654,N_22641,N_20843);
nand U29655 (N_29655,N_21365,N_20399);
nand U29656 (N_29656,N_22330,N_22392);
xor U29657 (N_29657,N_18441,N_19090);
xnor U29658 (N_29658,N_20428,N_23524);
or U29659 (N_29659,N_22739,N_20123);
xnor U29660 (N_29660,N_21649,N_20056);
nand U29661 (N_29661,N_22855,N_20999);
xnor U29662 (N_29662,N_21898,N_22939);
xnor U29663 (N_29663,N_20587,N_18240);
nand U29664 (N_29664,N_19478,N_18131);
xor U29665 (N_29665,N_20339,N_19114);
nor U29666 (N_29666,N_18476,N_19414);
and U29667 (N_29667,N_18186,N_20584);
nand U29668 (N_29668,N_18654,N_19612);
nor U29669 (N_29669,N_20464,N_21968);
nand U29670 (N_29670,N_22400,N_20864);
nor U29671 (N_29671,N_22106,N_22689);
or U29672 (N_29672,N_22587,N_23393);
or U29673 (N_29673,N_20355,N_18369);
or U29674 (N_29674,N_21864,N_22971);
or U29675 (N_29675,N_22026,N_18512);
xor U29676 (N_29676,N_20643,N_23877);
nand U29677 (N_29677,N_20713,N_18163);
or U29678 (N_29678,N_23591,N_20495);
xor U29679 (N_29679,N_21034,N_23530);
nand U29680 (N_29680,N_19797,N_18097);
or U29681 (N_29681,N_19201,N_23079);
or U29682 (N_29682,N_18911,N_22892);
xor U29683 (N_29683,N_21299,N_18198);
nor U29684 (N_29684,N_20718,N_22501);
nand U29685 (N_29685,N_19530,N_23400);
xnor U29686 (N_29686,N_22217,N_18938);
nand U29687 (N_29687,N_19485,N_20768);
and U29688 (N_29688,N_20411,N_19186);
or U29689 (N_29689,N_23106,N_19638);
xor U29690 (N_29690,N_18648,N_18053);
nor U29691 (N_29691,N_19027,N_22430);
and U29692 (N_29692,N_19027,N_22120);
xnor U29693 (N_29693,N_20392,N_21469);
nand U29694 (N_29694,N_20696,N_18108);
nand U29695 (N_29695,N_18839,N_21665);
or U29696 (N_29696,N_23464,N_20732);
xor U29697 (N_29697,N_20477,N_23021);
nor U29698 (N_29698,N_20008,N_20497);
or U29699 (N_29699,N_19024,N_23191);
xor U29700 (N_29700,N_19755,N_21083);
nor U29701 (N_29701,N_19105,N_20532);
and U29702 (N_29702,N_23320,N_22529);
nand U29703 (N_29703,N_20311,N_20674);
nand U29704 (N_29704,N_19559,N_21977);
xor U29705 (N_29705,N_21924,N_19397);
nor U29706 (N_29706,N_18816,N_22574);
and U29707 (N_29707,N_18225,N_22883);
nor U29708 (N_29708,N_20392,N_21950);
nand U29709 (N_29709,N_21036,N_20629);
or U29710 (N_29710,N_22416,N_21254);
xor U29711 (N_29711,N_21326,N_22830);
or U29712 (N_29712,N_21755,N_21455);
nand U29713 (N_29713,N_19465,N_21261);
nor U29714 (N_29714,N_20043,N_18271);
xnor U29715 (N_29715,N_23047,N_18160);
or U29716 (N_29716,N_22238,N_21545);
and U29717 (N_29717,N_23513,N_18072);
nor U29718 (N_29718,N_19054,N_19685);
or U29719 (N_29719,N_22449,N_20138);
xnor U29720 (N_29720,N_18146,N_20660);
xnor U29721 (N_29721,N_20819,N_23464);
or U29722 (N_29722,N_19765,N_18612);
nand U29723 (N_29723,N_21099,N_21702);
xor U29724 (N_29724,N_18166,N_18765);
nor U29725 (N_29725,N_20951,N_21621);
and U29726 (N_29726,N_20752,N_22849);
nor U29727 (N_29727,N_22361,N_20018);
nor U29728 (N_29728,N_20435,N_20632);
nor U29729 (N_29729,N_22769,N_23046);
nor U29730 (N_29730,N_22776,N_19032);
and U29731 (N_29731,N_22281,N_23719);
xor U29732 (N_29732,N_20182,N_23792);
or U29733 (N_29733,N_22756,N_21877);
or U29734 (N_29734,N_19461,N_23478);
or U29735 (N_29735,N_19952,N_18116);
nand U29736 (N_29736,N_18729,N_21499);
nor U29737 (N_29737,N_22474,N_20597);
and U29738 (N_29738,N_20722,N_20969);
and U29739 (N_29739,N_19281,N_19603);
and U29740 (N_29740,N_21287,N_23639);
nor U29741 (N_29741,N_20662,N_21641);
xnor U29742 (N_29742,N_23213,N_20631);
xnor U29743 (N_29743,N_20519,N_21922);
nor U29744 (N_29744,N_23975,N_19438);
xor U29745 (N_29745,N_22693,N_23702);
or U29746 (N_29746,N_23243,N_23934);
and U29747 (N_29747,N_18791,N_23186);
and U29748 (N_29748,N_21698,N_20137);
and U29749 (N_29749,N_23380,N_19001);
and U29750 (N_29750,N_18366,N_21934);
xor U29751 (N_29751,N_18993,N_19058);
and U29752 (N_29752,N_21837,N_23642);
or U29753 (N_29753,N_18159,N_23438);
nand U29754 (N_29754,N_21555,N_21399);
or U29755 (N_29755,N_20848,N_23478);
nor U29756 (N_29756,N_19246,N_18190);
nor U29757 (N_29757,N_22369,N_19312);
or U29758 (N_29758,N_19181,N_20743);
nand U29759 (N_29759,N_19279,N_20054);
and U29760 (N_29760,N_18704,N_20453);
or U29761 (N_29761,N_19410,N_19662);
nand U29762 (N_29762,N_18693,N_19523);
xor U29763 (N_29763,N_21921,N_23434);
or U29764 (N_29764,N_21549,N_22171);
and U29765 (N_29765,N_19931,N_22800);
or U29766 (N_29766,N_20452,N_22107);
or U29767 (N_29767,N_18313,N_20089);
xnor U29768 (N_29768,N_22218,N_19222);
nor U29769 (N_29769,N_23101,N_21005);
nand U29770 (N_29770,N_18076,N_19814);
nand U29771 (N_29771,N_22665,N_23640);
nor U29772 (N_29772,N_19336,N_20533);
or U29773 (N_29773,N_18897,N_20658);
or U29774 (N_29774,N_22134,N_22568);
or U29775 (N_29775,N_18953,N_20262);
nor U29776 (N_29776,N_21113,N_20523);
xor U29777 (N_29777,N_22867,N_21362);
nor U29778 (N_29778,N_20449,N_18599);
xnor U29779 (N_29779,N_20028,N_18961);
xor U29780 (N_29780,N_21965,N_23746);
xor U29781 (N_29781,N_19102,N_20356);
or U29782 (N_29782,N_20267,N_22695);
or U29783 (N_29783,N_19685,N_23365);
or U29784 (N_29784,N_19039,N_23937);
or U29785 (N_29785,N_22401,N_18815);
and U29786 (N_29786,N_21244,N_21210);
or U29787 (N_29787,N_23531,N_19806);
nor U29788 (N_29788,N_21680,N_19789);
nor U29789 (N_29789,N_19320,N_20294);
xor U29790 (N_29790,N_23799,N_20211);
nor U29791 (N_29791,N_20965,N_20597);
nor U29792 (N_29792,N_18734,N_18280);
nand U29793 (N_29793,N_23449,N_20437);
or U29794 (N_29794,N_20654,N_19594);
xor U29795 (N_29795,N_22274,N_22003);
xor U29796 (N_29796,N_21349,N_20855);
xnor U29797 (N_29797,N_18136,N_21346);
xor U29798 (N_29798,N_18205,N_22319);
nor U29799 (N_29799,N_20031,N_19652);
and U29800 (N_29800,N_22336,N_19739);
and U29801 (N_29801,N_19757,N_22974);
nor U29802 (N_29802,N_20735,N_23004);
nor U29803 (N_29803,N_18320,N_19684);
nand U29804 (N_29804,N_18720,N_19912);
nor U29805 (N_29805,N_19645,N_23318);
and U29806 (N_29806,N_22745,N_23781);
xor U29807 (N_29807,N_21427,N_23246);
or U29808 (N_29808,N_18574,N_19503);
and U29809 (N_29809,N_22664,N_19068);
or U29810 (N_29810,N_18061,N_20061);
and U29811 (N_29811,N_21298,N_22699);
nand U29812 (N_29812,N_20716,N_18790);
xnor U29813 (N_29813,N_19866,N_22761);
nor U29814 (N_29814,N_20357,N_18469);
xor U29815 (N_29815,N_18353,N_20711);
xor U29816 (N_29816,N_21602,N_20495);
nand U29817 (N_29817,N_21095,N_22030);
nor U29818 (N_29818,N_22890,N_19075);
nor U29819 (N_29819,N_21498,N_22925);
and U29820 (N_29820,N_23970,N_23735);
xnor U29821 (N_29821,N_19094,N_23704);
nand U29822 (N_29822,N_18710,N_21873);
and U29823 (N_29823,N_23544,N_20226);
xor U29824 (N_29824,N_18779,N_19030);
and U29825 (N_29825,N_18865,N_21612);
nand U29826 (N_29826,N_23507,N_18997);
nor U29827 (N_29827,N_22201,N_18684);
nor U29828 (N_29828,N_21500,N_20960);
xor U29829 (N_29829,N_21802,N_20212);
and U29830 (N_29830,N_20758,N_18863);
and U29831 (N_29831,N_20274,N_21488);
and U29832 (N_29832,N_23977,N_23672);
nor U29833 (N_29833,N_23408,N_20988);
and U29834 (N_29834,N_22515,N_21273);
nor U29835 (N_29835,N_18547,N_21614);
nor U29836 (N_29836,N_19639,N_22733);
nor U29837 (N_29837,N_20964,N_23359);
xor U29838 (N_29838,N_21817,N_20464);
and U29839 (N_29839,N_19206,N_21138);
or U29840 (N_29840,N_19086,N_22041);
or U29841 (N_29841,N_23711,N_21467);
nor U29842 (N_29842,N_19561,N_19576);
nor U29843 (N_29843,N_20493,N_18134);
and U29844 (N_29844,N_21871,N_22065);
or U29845 (N_29845,N_23357,N_20104);
nand U29846 (N_29846,N_22625,N_23220);
or U29847 (N_29847,N_19345,N_22644);
xnor U29848 (N_29848,N_21680,N_19593);
nand U29849 (N_29849,N_19991,N_19551);
or U29850 (N_29850,N_23645,N_23186);
and U29851 (N_29851,N_20782,N_20548);
or U29852 (N_29852,N_19787,N_21856);
and U29853 (N_29853,N_19445,N_20713);
nand U29854 (N_29854,N_18211,N_19156);
xnor U29855 (N_29855,N_21795,N_20910);
nor U29856 (N_29856,N_23624,N_22723);
nand U29857 (N_29857,N_18097,N_19238);
or U29858 (N_29858,N_20620,N_20938);
nand U29859 (N_29859,N_21863,N_19597);
or U29860 (N_29860,N_20152,N_20015);
and U29861 (N_29861,N_22780,N_18896);
nand U29862 (N_29862,N_18166,N_20940);
xnor U29863 (N_29863,N_20251,N_18475);
or U29864 (N_29864,N_23836,N_21943);
nor U29865 (N_29865,N_19029,N_19897);
xor U29866 (N_29866,N_19152,N_19986);
xnor U29867 (N_29867,N_18999,N_19046);
nand U29868 (N_29868,N_20058,N_21262);
nor U29869 (N_29869,N_18001,N_21171);
or U29870 (N_29870,N_18675,N_21548);
or U29871 (N_29871,N_22230,N_22287);
nor U29872 (N_29872,N_22817,N_23224);
nor U29873 (N_29873,N_20200,N_23943);
nand U29874 (N_29874,N_23172,N_22362);
nand U29875 (N_29875,N_22335,N_21873);
xnor U29876 (N_29876,N_21867,N_23567);
xor U29877 (N_29877,N_23309,N_21020);
nand U29878 (N_29878,N_23101,N_18475);
nor U29879 (N_29879,N_23508,N_22187);
and U29880 (N_29880,N_22744,N_23438);
xor U29881 (N_29881,N_18225,N_20246);
and U29882 (N_29882,N_23565,N_21131);
or U29883 (N_29883,N_21683,N_22793);
and U29884 (N_29884,N_22997,N_19941);
and U29885 (N_29885,N_19611,N_22507);
and U29886 (N_29886,N_18178,N_21117);
and U29887 (N_29887,N_18569,N_18452);
xor U29888 (N_29888,N_18050,N_19116);
nor U29889 (N_29889,N_23277,N_23861);
xnor U29890 (N_29890,N_18994,N_22572);
nor U29891 (N_29891,N_22868,N_22569);
xor U29892 (N_29892,N_19838,N_21430);
nand U29893 (N_29893,N_22335,N_18314);
nand U29894 (N_29894,N_19545,N_20602);
nor U29895 (N_29895,N_20976,N_23975);
and U29896 (N_29896,N_22242,N_18748);
or U29897 (N_29897,N_19271,N_20841);
and U29898 (N_29898,N_20985,N_19955);
nand U29899 (N_29899,N_20904,N_21981);
and U29900 (N_29900,N_22077,N_21422);
nor U29901 (N_29901,N_20318,N_22488);
nand U29902 (N_29902,N_23374,N_18171);
and U29903 (N_29903,N_21327,N_18079);
nor U29904 (N_29904,N_23512,N_21040);
nand U29905 (N_29905,N_21964,N_22193);
xor U29906 (N_29906,N_19671,N_23840);
and U29907 (N_29907,N_22274,N_20068);
and U29908 (N_29908,N_19619,N_22240);
nand U29909 (N_29909,N_22106,N_20002);
xnor U29910 (N_29910,N_19852,N_21944);
or U29911 (N_29911,N_21768,N_18286);
xnor U29912 (N_29912,N_22503,N_19281);
xor U29913 (N_29913,N_20560,N_20645);
or U29914 (N_29914,N_22849,N_20314);
nor U29915 (N_29915,N_18125,N_22381);
nand U29916 (N_29916,N_22730,N_19119);
nor U29917 (N_29917,N_23374,N_23083);
nand U29918 (N_29918,N_22007,N_22146);
nor U29919 (N_29919,N_22173,N_18473);
or U29920 (N_29920,N_22945,N_18871);
and U29921 (N_29921,N_18458,N_19869);
or U29922 (N_29922,N_19808,N_22325);
and U29923 (N_29923,N_23323,N_21410);
nor U29924 (N_29924,N_22614,N_18893);
nand U29925 (N_29925,N_20824,N_18025);
and U29926 (N_29926,N_23811,N_23236);
nand U29927 (N_29927,N_21259,N_18372);
nor U29928 (N_29928,N_23706,N_20628);
or U29929 (N_29929,N_21192,N_22250);
nor U29930 (N_29930,N_20598,N_22170);
xor U29931 (N_29931,N_18063,N_23938);
nand U29932 (N_29932,N_21650,N_20677);
and U29933 (N_29933,N_21915,N_20951);
nor U29934 (N_29934,N_19834,N_18353);
nand U29935 (N_29935,N_19482,N_19900);
or U29936 (N_29936,N_19361,N_18768);
or U29937 (N_29937,N_21688,N_23346);
or U29938 (N_29938,N_22819,N_22339);
and U29939 (N_29939,N_18986,N_21602);
nand U29940 (N_29940,N_22964,N_21289);
and U29941 (N_29941,N_21246,N_18177);
and U29942 (N_29942,N_22897,N_21843);
or U29943 (N_29943,N_21911,N_21913);
nor U29944 (N_29944,N_19341,N_21625);
nand U29945 (N_29945,N_18952,N_23743);
nor U29946 (N_29946,N_19511,N_22418);
xnor U29947 (N_29947,N_18917,N_19427);
nand U29948 (N_29948,N_21576,N_23122);
or U29949 (N_29949,N_19529,N_21630);
or U29950 (N_29950,N_22653,N_21192);
xnor U29951 (N_29951,N_18021,N_21057);
and U29952 (N_29952,N_20468,N_23839);
xnor U29953 (N_29953,N_18419,N_21966);
and U29954 (N_29954,N_18410,N_23440);
nor U29955 (N_29955,N_18051,N_20961);
xnor U29956 (N_29956,N_22381,N_23972);
or U29957 (N_29957,N_22264,N_21481);
xnor U29958 (N_29958,N_19359,N_20667);
or U29959 (N_29959,N_22208,N_21168);
nand U29960 (N_29960,N_19617,N_21152);
nor U29961 (N_29961,N_21424,N_20528);
or U29962 (N_29962,N_19957,N_20545);
xnor U29963 (N_29963,N_22822,N_22026);
or U29964 (N_29964,N_23199,N_20218);
and U29965 (N_29965,N_20618,N_22693);
and U29966 (N_29966,N_21060,N_20756);
or U29967 (N_29967,N_19079,N_20733);
xnor U29968 (N_29968,N_19030,N_21451);
nor U29969 (N_29969,N_20404,N_23773);
nor U29970 (N_29970,N_20763,N_19989);
and U29971 (N_29971,N_22802,N_23878);
xnor U29972 (N_29972,N_20669,N_22511);
or U29973 (N_29973,N_21875,N_20162);
xnor U29974 (N_29974,N_18033,N_20331);
xor U29975 (N_29975,N_19807,N_19094);
nand U29976 (N_29976,N_18408,N_18104);
nor U29977 (N_29977,N_22799,N_23921);
nor U29978 (N_29978,N_21705,N_19343);
xnor U29979 (N_29979,N_22859,N_18130);
xnor U29980 (N_29980,N_20713,N_20031);
nor U29981 (N_29981,N_18455,N_22927);
nor U29982 (N_29982,N_18323,N_23906);
nand U29983 (N_29983,N_23956,N_21748);
and U29984 (N_29984,N_22900,N_18982);
nand U29985 (N_29985,N_18503,N_23432);
or U29986 (N_29986,N_23197,N_19140);
nand U29987 (N_29987,N_20858,N_20698);
nand U29988 (N_29988,N_20586,N_22422);
nand U29989 (N_29989,N_21071,N_20565);
nand U29990 (N_29990,N_20203,N_22839);
nor U29991 (N_29991,N_20833,N_18779);
xor U29992 (N_29992,N_22178,N_18959);
nand U29993 (N_29993,N_21094,N_22673);
and U29994 (N_29994,N_21073,N_20306);
nor U29995 (N_29995,N_20766,N_20446);
nand U29996 (N_29996,N_21305,N_20915);
or U29997 (N_29997,N_18088,N_21041);
nand U29998 (N_29998,N_18669,N_21086);
nand U29999 (N_29999,N_19985,N_22089);
and UO_0 (O_0,N_26263,N_24752);
xor UO_1 (O_1,N_26855,N_26079);
or UO_2 (O_2,N_26222,N_24607);
and UO_3 (O_3,N_27427,N_25302);
xnor UO_4 (O_4,N_28605,N_28339);
xnor UO_5 (O_5,N_25147,N_26898);
or UO_6 (O_6,N_28386,N_28259);
nor UO_7 (O_7,N_28324,N_28380);
xnor UO_8 (O_8,N_25219,N_25986);
nor UO_9 (O_9,N_24118,N_29002);
xor UO_10 (O_10,N_29418,N_28650);
or UO_11 (O_11,N_28274,N_27737);
and UO_12 (O_12,N_28319,N_25179);
nor UO_13 (O_13,N_25546,N_26832);
and UO_14 (O_14,N_25169,N_24332);
nand UO_15 (O_15,N_24512,N_26108);
xnor UO_16 (O_16,N_27595,N_26385);
xor UO_17 (O_17,N_28614,N_27443);
nor UO_18 (O_18,N_25806,N_26438);
nand UO_19 (O_19,N_29786,N_29609);
nor UO_20 (O_20,N_26609,N_27319);
or UO_21 (O_21,N_28198,N_25938);
or UO_22 (O_22,N_25790,N_25225);
and UO_23 (O_23,N_24331,N_29707);
or UO_24 (O_24,N_26631,N_26544);
xnor UO_25 (O_25,N_26602,N_25077);
and UO_26 (O_26,N_25070,N_26056);
or UO_27 (O_27,N_28766,N_24440);
or UO_28 (O_28,N_28857,N_29496);
nor UO_29 (O_29,N_28648,N_24534);
and UO_30 (O_30,N_29839,N_26261);
and UO_31 (O_31,N_24961,N_25387);
or UO_32 (O_32,N_27510,N_24031);
nor UO_33 (O_33,N_26052,N_25586);
nand UO_34 (O_34,N_25705,N_26738);
and UO_35 (O_35,N_27356,N_24564);
nand UO_36 (O_36,N_24115,N_25828);
xor UO_37 (O_37,N_26600,N_24884);
or UO_38 (O_38,N_26878,N_29508);
xnor UO_39 (O_39,N_26304,N_29924);
xor UO_40 (O_40,N_25391,N_28726);
nand UO_41 (O_41,N_26007,N_24436);
or UO_42 (O_42,N_29742,N_24806);
nand UO_43 (O_43,N_28204,N_28978);
or UO_44 (O_44,N_24342,N_28351);
and UO_45 (O_45,N_27483,N_24729);
nor UO_46 (O_46,N_28753,N_29874);
nor UO_47 (O_47,N_26861,N_28475);
and UO_48 (O_48,N_29853,N_24892);
xor UO_49 (O_49,N_25029,N_28785);
xnor UO_50 (O_50,N_29128,N_27321);
and UO_51 (O_51,N_24507,N_28244);
and UO_52 (O_52,N_26800,N_24482);
nand UO_53 (O_53,N_26650,N_27590);
xnor UO_54 (O_54,N_27948,N_26257);
nand UO_55 (O_55,N_26021,N_26732);
xnor UO_56 (O_56,N_24837,N_29708);
nor UO_57 (O_57,N_29771,N_28904);
or UO_58 (O_58,N_27451,N_28360);
and UO_59 (O_59,N_24264,N_29829);
and UO_60 (O_60,N_29628,N_28188);
or UO_61 (O_61,N_29345,N_24553);
or UO_62 (O_62,N_28910,N_27278);
or UO_63 (O_63,N_24243,N_24266);
or UO_64 (O_64,N_29437,N_27576);
nor UO_65 (O_65,N_24499,N_27612);
nand UO_66 (O_66,N_28315,N_25470);
and UO_67 (O_67,N_24084,N_27669);
or UO_68 (O_68,N_26493,N_25146);
nand UO_69 (O_69,N_25587,N_28252);
nand UO_70 (O_70,N_25492,N_25199);
and UO_71 (O_71,N_29895,N_29433);
nor UO_72 (O_72,N_28589,N_25859);
and UO_73 (O_73,N_26024,N_29166);
nand UO_74 (O_74,N_28828,N_26842);
xnor UO_75 (O_75,N_24383,N_26167);
xor UO_76 (O_76,N_29423,N_29312);
xor UO_77 (O_77,N_25092,N_26607);
and UO_78 (O_78,N_24595,N_28019);
xnor UO_79 (O_79,N_26020,N_25817);
and UO_80 (O_80,N_26423,N_26075);
or UO_81 (O_81,N_28496,N_24705);
nor UO_82 (O_82,N_24157,N_29255);
nand UO_83 (O_83,N_26319,N_27051);
xnor UO_84 (O_84,N_27268,N_29144);
and UO_85 (O_85,N_25295,N_28058);
nand UO_86 (O_86,N_24171,N_27570);
xnor UO_87 (O_87,N_27238,N_25590);
nand UO_88 (O_88,N_29751,N_28584);
or UO_89 (O_89,N_24078,N_29583);
nand UO_90 (O_90,N_28957,N_28615);
nand UO_91 (O_91,N_28302,N_25410);
nor UO_92 (O_92,N_29823,N_27432);
xor UO_93 (O_93,N_29124,N_26223);
nand UO_94 (O_94,N_26339,N_25548);
xnor UO_95 (O_95,N_27758,N_29197);
or UO_96 (O_96,N_24057,N_26403);
nor UO_97 (O_97,N_25380,N_28711);
and UO_98 (O_98,N_24307,N_24364);
and UO_99 (O_99,N_24176,N_29266);
nor UO_100 (O_100,N_27435,N_26704);
and UO_101 (O_101,N_29362,N_24346);
or UO_102 (O_102,N_27607,N_28500);
or UO_103 (O_103,N_25301,N_28378);
xnor UO_104 (O_104,N_27823,N_25687);
and UO_105 (O_105,N_24645,N_29797);
xnor UO_106 (O_106,N_27724,N_25190);
nand UO_107 (O_107,N_28119,N_26958);
nand UO_108 (O_108,N_26269,N_24460);
nand UO_109 (O_109,N_26298,N_25908);
xor UO_110 (O_110,N_28431,N_29885);
nand UO_111 (O_111,N_25918,N_27281);
nor UO_112 (O_112,N_27254,N_26286);
and UO_113 (O_113,N_26813,N_27683);
or UO_114 (O_114,N_24831,N_28757);
nor UO_115 (O_115,N_24032,N_25286);
and UO_116 (O_116,N_28945,N_25030);
nand UO_117 (O_117,N_26926,N_26457);
nor UO_118 (O_118,N_26954,N_25107);
and UO_119 (O_119,N_27888,N_27565);
xor UO_120 (O_120,N_27585,N_29059);
and UO_121 (O_121,N_25799,N_25788);
nand UO_122 (O_122,N_26164,N_24672);
or UO_123 (O_123,N_28440,N_24642);
nor UO_124 (O_124,N_29611,N_25108);
or UO_125 (O_125,N_25969,N_25171);
or UO_126 (O_126,N_25943,N_24249);
xnor UO_127 (O_127,N_24721,N_25839);
nor UO_128 (O_128,N_25671,N_27566);
nand UO_129 (O_129,N_24393,N_26012);
nor UO_130 (O_130,N_29222,N_24424);
xor UO_131 (O_131,N_24166,N_26488);
nor UO_132 (O_132,N_29101,N_27863);
or UO_133 (O_133,N_25393,N_27378);
nor UO_134 (O_134,N_25456,N_28674);
nand UO_135 (O_135,N_24636,N_27347);
nand UO_136 (O_136,N_24086,N_28989);
nand UO_137 (O_137,N_26684,N_28758);
nor UO_138 (O_138,N_24802,N_28898);
or UO_139 (O_139,N_29451,N_26072);
or UO_140 (O_140,N_29097,N_28092);
and UO_141 (O_141,N_27946,N_28133);
nor UO_142 (O_142,N_26642,N_27602);
nand UO_143 (O_143,N_26256,N_28097);
nand UO_144 (O_144,N_29023,N_25259);
nand UO_145 (O_145,N_24962,N_28503);
and UO_146 (O_146,N_29231,N_24140);
nor UO_147 (O_147,N_25751,N_28723);
nand UO_148 (O_148,N_25804,N_24849);
and UO_149 (O_149,N_24898,N_29034);
xnor UO_150 (O_150,N_24174,N_26182);
nand UO_151 (O_151,N_26985,N_24133);
or UO_152 (O_152,N_28810,N_27255);
and UO_153 (O_153,N_24594,N_24568);
xor UO_154 (O_154,N_27847,N_26919);
or UO_155 (O_155,N_27145,N_27695);
nor UO_156 (O_156,N_29663,N_24798);
nand UO_157 (O_157,N_28963,N_29090);
nor UO_158 (O_158,N_27969,N_28523);
nor UO_159 (O_159,N_27620,N_26494);
xor UO_160 (O_160,N_26165,N_27790);
or UO_161 (O_161,N_24488,N_26364);
nand UO_162 (O_162,N_24352,N_25704);
or UO_163 (O_163,N_28438,N_28173);
and UO_164 (O_164,N_24565,N_25140);
nand UO_165 (O_165,N_29893,N_29820);
and UO_166 (O_166,N_26307,N_29843);
xor UO_167 (O_167,N_26295,N_24212);
xor UO_168 (O_168,N_27606,N_25215);
and UO_169 (O_169,N_29701,N_25985);
nand UO_170 (O_170,N_24469,N_28506);
nand UO_171 (O_171,N_27926,N_26825);
nor UO_172 (O_172,N_24492,N_27008);
nand UO_173 (O_173,N_24984,N_25952);
xor UO_174 (O_174,N_26288,N_24517);
and UO_175 (O_175,N_28736,N_26094);
and UO_176 (O_176,N_26977,N_25414);
xor UO_177 (O_177,N_26915,N_29268);
or UO_178 (O_178,N_29281,N_24696);
nand UO_179 (O_179,N_25231,N_24301);
nand UO_180 (O_180,N_29043,N_28333);
and UO_181 (O_181,N_27980,N_25716);
xor UO_182 (O_182,N_25399,N_24411);
nor UO_183 (O_183,N_27588,N_29119);
xnor UO_184 (O_184,N_27225,N_25931);
or UO_185 (O_185,N_29486,N_28514);
xor UO_186 (O_186,N_27126,N_26949);
nand UO_187 (O_187,N_24567,N_28236);
xor UO_188 (O_188,N_27558,N_25981);
xnor UO_189 (O_189,N_29511,N_29572);
nor UO_190 (O_190,N_28237,N_26933);
and UO_191 (O_191,N_24280,N_28468);
nor UO_192 (O_192,N_27431,N_27809);
xor UO_193 (O_193,N_26310,N_28721);
xor UO_194 (O_194,N_24043,N_27957);
nand UO_195 (O_195,N_27404,N_26584);
nor UO_196 (O_196,N_27913,N_24256);
and UO_197 (O_197,N_28307,N_26174);
and UO_198 (O_198,N_25323,N_25723);
and UO_199 (O_199,N_26003,N_25005);
nor UO_200 (O_200,N_27346,N_28825);
or UO_201 (O_201,N_25252,N_29669);
or UO_202 (O_202,N_29997,N_24953);
xor UO_203 (O_203,N_25953,N_29921);
nor UO_204 (O_204,N_28200,N_26992);
or UO_205 (O_205,N_25529,N_27376);
or UO_206 (O_206,N_26141,N_27975);
and UO_207 (O_207,N_27793,N_27977);
nor UO_208 (O_208,N_26712,N_24551);
nor UO_209 (O_209,N_24926,N_28781);
nand UO_210 (O_210,N_27954,N_27991);
or UO_211 (O_211,N_24921,N_26880);
and UO_212 (O_212,N_27932,N_27224);
and UO_213 (O_213,N_25417,N_28365);
and UO_214 (O_214,N_27244,N_29354);
nor UO_215 (O_215,N_26260,N_24593);
and UO_216 (O_216,N_25018,N_25271);
nand UO_217 (O_217,N_25111,N_29322);
and UO_218 (O_218,N_24085,N_29988);
nand UO_219 (O_219,N_28902,N_26535);
nor UO_220 (O_220,N_29524,N_26196);
or UO_221 (O_221,N_26472,N_29803);
nand UO_222 (O_222,N_25982,N_28657);
xnor UO_223 (O_223,N_25376,N_26092);
nor UO_224 (O_224,N_25383,N_26965);
nand UO_225 (O_225,N_26848,N_28722);
xnor UO_226 (O_226,N_27139,N_29850);
nor UO_227 (O_227,N_26725,N_29242);
nor UO_228 (O_228,N_29054,N_28675);
or UO_229 (O_229,N_24799,N_24856);
and UO_230 (O_230,N_24121,N_28559);
or UO_231 (O_231,N_26785,N_25448);
nor UO_232 (O_232,N_28008,N_25877);
xor UO_233 (O_233,N_24199,N_28621);
nor UO_234 (O_234,N_24107,N_25277);
xor UO_235 (O_235,N_26900,N_26904);
nor UO_236 (O_236,N_24136,N_27189);
or UO_237 (O_237,N_25032,N_27613);
or UO_238 (O_238,N_25896,N_25400);
nor UO_239 (O_239,N_28783,N_29052);
nand UO_240 (O_240,N_25866,N_28970);
nor UO_241 (O_241,N_25506,N_26990);
or UO_242 (O_242,N_27466,N_29851);
nor UO_243 (O_243,N_28918,N_25436);
nor UO_244 (O_244,N_29728,N_27961);
nand UO_245 (O_245,N_26437,N_27052);
nand UO_246 (O_246,N_26104,N_28132);
xor UO_247 (O_247,N_26357,N_29965);
and UO_248 (O_248,N_24152,N_25876);
nor UO_249 (O_249,N_25685,N_27086);
and UO_250 (O_250,N_27677,N_28733);
nand UO_251 (O_251,N_29621,N_27955);
nand UO_252 (O_252,N_24582,N_26581);
nand UO_253 (O_253,N_29678,N_26883);
nand UO_254 (O_254,N_25308,N_25700);
xnor UO_255 (O_255,N_25939,N_25006);
xnor UO_256 (O_256,N_29681,N_25475);
and UO_257 (O_257,N_28653,N_25460);
and UO_258 (O_258,N_27235,N_26081);
and UO_259 (O_259,N_29982,N_26790);
nor UO_260 (O_260,N_24833,N_28084);
or UO_261 (O_261,N_25929,N_29349);
nand UO_262 (O_262,N_27825,N_27855);
or UO_263 (O_263,N_29382,N_26711);
or UO_264 (O_264,N_29155,N_24759);
and UO_265 (O_265,N_29537,N_28344);
or UO_266 (O_266,N_27640,N_25772);
or UO_267 (O_267,N_28455,N_28376);
and UO_268 (O_268,N_27217,N_25749);
xor UO_269 (O_269,N_27937,N_29374);
or UO_270 (O_270,N_24255,N_26666);
and UO_271 (O_271,N_29233,N_27058);
and UO_272 (O_272,N_29779,N_29236);
and UO_273 (O_273,N_29688,N_26466);
xor UO_274 (O_274,N_24028,N_25442);
and UO_275 (O_275,N_24971,N_29417);
or UO_276 (O_276,N_29864,N_24985);
xor UO_277 (O_277,N_28889,N_28914);
nor UO_278 (O_278,N_28035,N_25454);
nor UO_279 (O_279,N_29446,N_25501);
or UO_280 (O_280,N_29884,N_28743);
nand UO_281 (O_281,N_27958,N_25083);
nand UO_282 (O_282,N_27622,N_24468);
xnor UO_283 (O_283,N_27207,N_24735);
and UO_284 (O_284,N_25214,N_28537);
and UO_285 (O_285,N_26103,N_25046);
and UO_286 (O_286,N_25604,N_24135);
nand UO_287 (O_287,N_27681,N_28961);
xnor UO_288 (O_288,N_29217,N_25152);
nand UO_289 (O_289,N_28972,N_25686);
or UO_290 (O_290,N_25559,N_26957);
nand UO_291 (O_291,N_29378,N_28128);
or UO_292 (O_292,N_25395,N_24196);
nor UO_293 (O_293,N_25254,N_24033);
nand UO_294 (O_294,N_25249,N_29402);
xor UO_295 (O_295,N_29713,N_24261);
or UO_296 (O_296,N_27332,N_27384);
xnor UO_297 (O_297,N_26213,N_26585);
nor UO_298 (O_298,N_26956,N_24502);
and UO_299 (O_299,N_28491,N_26124);
nand UO_300 (O_300,N_24134,N_25033);
nand UO_301 (O_301,N_24791,N_28059);
nand UO_302 (O_302,N_27591,N_25620);
nor UO_303 (O_303,N_26080,N_26264);
xnor UO_304 (O_304,N_24008,N_25420);
and UO_305 (O_305,N_26246,N_29710);
or UO_306 (O_306,N_29332,N_25059);
and UO_307 (O_307,N_27703,N_29557);
nand UO_308 (O_308,N_29393,N_27994);
and UO_309 (O_309,N_25204,N_29313);
xor UO_310 (O_310,N_27826,N_25955);
xor UO_311 (O_311,N_26728,N_24194);
xor UO_312 (O_312,N_24357,N_24385);
or UO_313 (O_313,N_26947,N_26756);
nor UO_314 (O_314,N_26185,N_27858);
and UO_315 (O_315,N_25625,N_24302);
and UO_316 (O_316,N_28213,N_26568);
and UO_317 (O_317,N_28301,N_27779);
or UO_318 (O_318,N_28962,N_24070);
or UO_319 (O_319,N_28007,N_28212);
nor UO_320 (O_320,N_25051,N_29804);
xor UO_321 (O_321,N_24144,N_25827);
nor UO_322 (O_322,N_26446,N_24699);
xor UO_323 (O_323,N_28925,N_29290);
nand UO_324 (O_324,N_24919,N_27109);
nand UO_325 (O_325,N_24706,N_25947);
and UO_326 (O_326,N_26162,N_24844);
nor UO_327 (O_327,N_25893,N_24726);
or UO_328 (O_328,N_26123,N_24614);
nand UO_329 (O_329,N_24753,N_27871);
nor UO_330 (O_330,N_29338,N_24501);
nor UO_331 (O_331,N_28091,N_24251);
and UO_332 (O_332,N_27434,N_26896);
and UO_333 (O_333,N_24841,N_25021);
xor UO_334 (O_334,N_29685,N_24649);
nor UO_335 (O_335,N_25210,N_25912);
and UO_336 (O_336,N_26248,N_26614);
nand UO_337 (O_337,N_24093,N_25889);
nand UO_338 (O_338,N_29759,N_28966);
nand UO_339 (O_339,N_29160,N_25481);
or UO_340 (O_340,N_29178,N_25372);
and UO_341 (O_341,N_24328,N_24288);
and UO_342 (O_342,N_29186,N_27929);
or UO_343 (O_343,N_28004,N_25637);
or UO_344 (O_344,N_24972,N_24345);
nand UO_345 (O_345,N_24886,N_26850);
nor UO_346 (O_346,N_24177,N_25494);
nand UO_347 (O_347,N_26690,N_28363);
nor UO_348 (O_348,N_29311,N_28974);
nor UO_349 (O_349,N_29651,N_24524);
and UO_350 (O_350,N_26018,N_26541);
or UO_351 (O_351,N_25719,N_29088);
nand UO_352 (O_352,N_28065,N_27261);
nand UO_353 (O_353,N_26244,N_29932);
xnor UO_354 (O_354,N_24448,N_28531);
nand UO_355 (O_355,N_29021,N_28156);
and UO_356 (O_356,N_28478,N_25674);
and UO_357 (O_357,N_24125,N_27582);
and UO_358 (O_358,N_24022,N_28243);
nand UO_359 (O_359,N_26909,N_25224);
xor UO_360 (O_360,N_26941,N_26486);
nor UO_361 (O_361,N_26221,N_25792);
xor UO_362 (O_362,N_24771,N_26918);
nor UO_363 (O_363,N_26573,N_28172);
nor UO_364 (O_364,N_28374,N_26176);
or UO_365 (O_365,N_27845,N_27033);
and UO_366 (O_366,N_25415,N_24644);
nand UO_367 (O_367,N_25446,N_29276);
and UO_368 (O_368,N_27773,N_25776);
nand UO_369 (O_369,N_29750,N_29598);
nor UO_370 (O_370,N_26210,N_27410);
or UO_371 (O_371,N_29964,N_27029);
or UO_372 (O_372,N_29764,N_29623);
or UO_373 (O_373,N_25557,N_29350);
nor UO_374 (O_374,N_29879,N_29722);
nand UO_375 (O_375,N_24800,N_26492);
nor UO_376 (O_376,N_28170,N_27127);
nand UO_377 (O_377,N_29387,N_29974);
nor UO_378 (O_378,N_28501,N_28806);
and UO_379 (O_379,N_27712,N_27436);
nor UO_380 (O_380,N_27036,N_29343);
or UO_381 (O_381,N_27608,N_26531);
nand UO_382 (O_382,N_26337,N_28793);
xnor UO_383 (O_383,N_28026,N_27223);
nand UO_384 (O_384,N_27220,N_24425);
nand UO_385 (O_385,N_24077,N_29258);
and UO_386 (O_386,N_26193,N_25228);
nand UO_387 (O_387,N_27997,N_28887);
and UO_388 (O_388,N_29111,N_25125);
xor UO_389 (O_389,N_27775,N_29519);
nor UO_390 (O_390,N_29140,N_29010);
and UO_391 (O_391,N_29042,N_25669);
nor UO_392 (O_392,N_24827,N_25026);
nor UO_393 (O_393,N_27234,N_26554);
nand UO_394 (O_394,N_25596,N_27045);
nor UO_395 (O_395,N_25334,N_29541);
or UO_396 (O_396,N_26516,N_28466);
nor UO_397 (O_397,N_24178,N_24306);
nand UO_398 (O_398,N_24000,N_27993);
and UO_399 (O_399,N_28534,N_28261);
xor UO_400 (O_400,N_24957,N_25621);
or UO_401 (O_401,N_24096,N_27354);
nor UO_402 (O_402,N_28687,N_26910);
xnor UO_403 (O_403,N_29815,N_29284);
or UO_404 (O_404,N_25694,N_24375);
nand UO_405 (O_405,N_27289,N_25512);
and UO_406 (O_406,N_29250,N_26950);
nor UO_407 (O_407,N_26859,N_26101);
nand UO_408 (O_408,N_24337,N_27939);
or UO_409 (O_409,N_25619,N_26552);
nand UO_410 (O_410,N_26394,N_26480);
or UO_411 (O_411,N_24730,N_29832);
nand UO_412 (O_412,N_24012,N_28320);
xnor UO_413 (O_413,N_24579,N_24542);
nand UO_414 (O_414,N_25042,N_25511);
and UO_415 (O_415,N_28557,N_28658);
or UO_416 (O_416,N_27260,N_24903);
and UO_417 (O_417,N_28412,N_25582);
nor UO_418 (O_418,N_29655,N_27144);
xnor UO_419 (O_419,N_25008,N_26200);
nand UO_420 (O_420,N_27074,N_27200);
or UO_421 (O_421,N_25297,N_27867);
and UO_422 (O_422,N_26542,N_26287);
xor UO_423 (O_423,N_24538,N_28926);
nand UO_424 (O_424,N_25978,N_25367);
nand UO_425 (O_425,N_29676,N_29272);
xor UO_426 (O_426,N_29943,N_27394);
nand UO_427 (O_427,N_24571,N_25329);
xor UO_428 (O_428,N_25285,N_27022);
nor UO_429 (O_429,N_28416,N_26456);
xor UO_430 (O_430,N_24866,N_24430);
xnor UO_431 (O_431,N_24792,N_24058);
nand UO_432 (O_432,N_25319,N_29280);
or UO_433 (O_433,N_24518,N_24300);
nand UO_434 (O_434,N_27341,N_27350);
nor UO_435 (O_435,N_28276,N_24505);
and UO_436 (O_436,N_29102,N_24338);
or UO_437 (O_437,N_29546,N_29207);
or UO_438 (O_438,N_28022,N_27942);
and UO_439 (O_439,N_25370,N_26545);
and UO_440 (O_440,N_28710,N_27917);
nor UO_441 (O_441,N_27966,N_24023);
and UO_442 (O_442,N_28778,N_26736);
or UO_443 (O_443,N_24704,N_29979);
nand UO_444 (O_444,N_27985,N_27334);
nor UO_445 (O_445,N_25269,N_24702);
and UO_446 (O_446,N_25795,N_26181);
xor UO_447 (O_447,N_24404,N_29954);
or UO_448 (O_448,N_24228,N_26186);
nand UO_449 (O_449,N_25386,N_24225);
nand UO_450 (O_450,N_27006,N_25364);
xor UO_451 (O_451,N_29246,N_26683);
nor UO_452 (O_452,N_27073,N_24749);
or UO_453 (O_453,N_26546,N_27742);
nand UO_454 (O_454,N_26377,N_28700);
nand UO_455 (O_455,N_26211,N_28473);
nor UO_456 (O_456,N_29145,N_25802);
xnor UO_457 (O_457,N_26594,N_28211);
xnor UO_458 (O_458,N_25126,N_26460);
nand UO_459 (O_459,N_25882,N_26380);
nand UO_460 (O_460,N_24592,N_26672);
and UO_461 (O_461,N_29224,N_27069);
or UO_462 (O_462,N_26139,N_26349);
nor UO_463 (O_463,N_29522,N_24528);
or UO_464 (O_464,N_27979,N_28773);
xnor UO_465 (O_465,N_28193,N_25177);
nor UO_466 (O_466,N_27514,N_29976);
nor UO_467 (O_467,N_28317,N_29748);
or UO_468 (O_468,N_26784,N_25525);
or UO_469 (O_469,N_27699,N_25754);
nor UO_470 (O_470,N_25291,N_25536);
nor UO_471 (O_471,N_25713,N_29099);
or UO_472 (O_472,N_24560,N_27174);
and UO_473 (O_473,N_28414,N_25173);
xnor UO_474 (O_474,N_26305,N_28250);
xor UO_475 (O_475,N_28239,N_29361);
nor UO_476 (O_476,N_24283,N_26844);
nor UO_477 (O_477,N_26641,N_26077);
and UO_478 (O_478,N_29784,N_25491);
or UO_479 (O_479,N_25076,N_27201);
and UO_480 (O_480,N_25532,N_29585);
and UO_481 (O_481,N_27827,N_27209);
and UO_482 (O_482,N_25545,N_27600);
nor UO_483 (O_483,N_28121,N_27971);
or UO_484 (O_484,N_24610,N_28952);
or UO_485 (O_485,N_27328,N_27623);
and UO_486 (O_486,N_26467,N_26114);
xnor UO_487 (O_487,N_29904,N_24750);
nand UO_488 (O_488,N_25745,N_29136);
xor UO_489 (O_489,N_29846,N_27284);
and UO_490 (O_490,N_29617,N_24738);
nor UO_491 (O_491,N_29720,N_24409);
xor UO_492 (O_492,N_24935,N_27248);
and UO_493 (O_493,N_25535,N_27009);
or UO_494 (O_494,N_26562,N_29934);
nor UO_495 (O_495,N_28994,N_24494);
xnor UO_496 (O_496,N_26091,N_25944);
or UO_497 (O_497,N_29562,N_26924);
nor UO_498 (O_498,N_27567,N_27584);
or UO_499 (O_499,N_27806,N_26343);
or UO_500 (O_500,N_29060,N_27479);
or UO_501 (O_501,N_24286,N_24719);
nor UO_502 (O_502,N_25401,N_27112);
and UO_503 (O_503,N_28591,N_29176);
nand UO_504 (O_504,N_29892,N_24793);
or UO_505 (O_505,N_27723,N_26363);
nand UO_506 (O_506,N_25449,N_26061);
or UO_507 (O_507,N_26431,N_24195);
or UO_508 (O_508,N_25578,N_25468);
xor UO_509 (O_509,N_27380,N_28797);
nor UO_510 (O_510,N_28441,N_24539);
or UO_511 (O_511,N_24048,N_28127);
nor UO_512 (O_512,N_26538,N_28734);
nor UO_513 (O_513,N_28906,N_25913);
or UO_514 (O_514,N_29448,N_29113);
nor UO_515 (O_515,N_26425,N_25881);
xor UO_516 (O_516,N_24974,N_25137);
xor UO_517 (O_517,N_29502,N_26359);
nand UO_518 (O_518,N_28928,N_26434);
or UO_519 (O_519,N_25887,N_29824);
or UO_520 (O_520,N_25755,N_24525);
nand UO_521 (O_521,N_27850,N_25483);
nor UO_522 (O_522,N_28922,N_27098);
xnor UO_523 (O_523,N_25309,N_25211);
nor UO_524 (O_524,N_24004,N_29092);
nor UO_525 (O_525,N_28990,N_24526);
nor UO_526 (O_526,N_28039,N_29861);
xnor UO_527 (O_527,N_26620,N_29653);
or UO_528 (O_528,N_26578,N_27323);
nor UO_529 (O_529,N_25937,N_26234);
and UO_530 (O_530,N_28768,N_27170);
nand UO_531 (O_531,N_26057,N_24487);
or UO_532 (O_532,N_27020,N_25445);
xnor UO_533 (O_533,N_26235,N_25734);
and UO_534 (O_534,N_29143,N_24398);
and UO_535 (O_535,N_24511,N_29767);
and UO_536 (O_536,N_27489,N_24271);
nor UO_537 (O_537,N_26503,N_28072);
xnor UO_538 (O_538,N_25885,N_24390);
nand UO_539 (O_539,N_26283,N_29295);
and UO_540 (O_540,N_26441,N_26444);
xnor UO_541 (O_541,N_28425,N_28370);
nand UO_542 (O_542,N_27064,N_25624);
and UO_543 (O_543,N_29789,N_24627);
nor UO_544 (O_544,N_24311,N_27119);
and UO_545 (O_545,N_25392,N_24608);
nor UO_546 (O_546,N_27160,N_29114);
and UO_547 (O_547,N_25406,N_27387);
nand UO_548 (O_548,N_27273,N_27700);
nor UO_549 (O_549,N_25612,N_25144);
nand UO_550 (O_550,N_29770,N_24334);
xor UO_551 (O_551,N_27880,N_27540);
nor UO_552 (O_552,N_27359,N_25900);
and UO_553 (O_553,N_27054,N_28705);
and UO_554 (O_554,N_25725,N_28813);
nand UO_555 (O_555,N_25697,N_28995);
xor UO_556 (O_556,N_26588,N_28960);
or UO_557 (O_557,N_27512,N_24668);
xor UO_558 (O_558,N_24414,N_26792);
and UO_559 (O_559,N_25594,N_24558);
nand UO_560 (O_560,N_26512,N_24349);
or UO_561 (O_561,N_24954,N_29918);
or UO_562 (O_562,N_25017,N_29237);
or UO_563 (O_563,N_29299,N_29152);
or UO_564 (O_564,N_28347,N_24814);
and UO_565 (O_565,N_26206,N_27448);
nor UO_566 (O_566,N_26879,N_24964);
xor UO_567 (O_567,N_25258,N_29082);
and UO_568 (O_568,N_28556,N_29105);
xnor UO_569 (O_569,N_24698,N_27759);
nor UO_570 (O_570,N_24027,N_26135);
or UO_571 (O_571,N_28628,N_26521);
nor UO_572 (O_572,N_29961,N_29775);
or UO_573 (O_573,N_29476,N_25066);
xnor UO_574 (O_574,N_25670,N_26701);
nor UO_575 (O_575,N_29896,N_28358);
or UO_576 (O_576,N_24456,N_29027);
and UO_577 (O_577,N_25085,N_28707);
nor UO_578 (O_578,N_28866,N_27240);
or UO_579 (O_579,N_26517,N_24629);
nand UO_580 (O_580,N_28158,N_29497);
xor UO_581 (O_581,N_24211,N_25547);
or UO_582 (O_582,N_27158,N_27077);
and UO_583 (O_583,N_26328,N_25970);
xor UO_584 (O_584,N_26816,N_28411);
or UO_585 (O_585,N_24535,N_29481);
nor UO_586 (O_586,N_24029,N_29983);
nor UO_587 (O_587,N_25925,N_26688);
xnor UO_588 (O_588,N_24223,N_29203);
and UO_589 (O_589,N_27470,N_25056);
xnor UO_590 (O_590,N_26410,N_26872);
nand UO_591 (O_591,N_29894,N_25759);
nor UO_592 (O_592,N_29302,N_27945);
nand UO_593 (O_593,N_24956,N_25605);
or UO_594 (O_594,N_26657,N_28706);
or UO_595 (O_595,N_29859,N_25983);
nand UO_596 (O_596,N_29328,N_24397);
nand UO_597 (O_597,N_24060,N_28812);
nor UO_598 (O_598,N_24758,N_25666);
or UO_599 (O_599,N_28522,N_25337);
and UO_600 (O_600,N_27277,N_27252);
nand UO_601 (O_601,N_26299,N_26694);
nor UO_602 (O_602,N_28727,N_29243);
or UO_603 (O_603,N_27501,N_24683);
nor UO_604 (O_604,N_28135,N_25848);
and UO_605 (O_605,N_27487,N_25296);
xor UO_606 (O_606,N_28608,N_26571);
nand UO_607 (O_607,N_29697,N_24407);
or UO_608 (O_608,N_25658,N_29800);
xor UO_609 (O_609,N_25892,N_28131);
xnor UO_610 (O_610,N_29373,N_24103);
or UO_611 (O_611,N_24110,N_25515);
nand UO_612 (O_612,N_27784,N_27760);
nand UO_613 (O_613,N_28427,N_24433);
or UO_614 (O_614,N_25366,N_27719);
and UO_615 (O_615,N_27162,N_25579);
and UO_616 (O_616,N_26547,N_26044);
nand UO_617 (O_617,N_28481,N_26769);
and UO_618 (O_618,N_27425,N_25439);
or UO_619 (O_619,N_28551,N_29639);
and UO_620 (O_620,N_27177,N_26705);
nor UO_621 (O_621,N_28842,N_25540);
nor UO_622 (O_622,N_25087,N_24080);
nor UO_623 (O_623,N_26700,N_25155);
nand UO_624 (O_624,N_28222,N_25539);
nand UO_625 (O_625,N_24741,N_25408);
xor UO_626 (O_626,N_28920,N_29151);
and UO_627 (O_627,N_24959,N_29110);
nand UO_628 (O_628,N_24944,N_29869);
and UO_629 (O_629,N_25926,N_26969);
xnor UO_630 (O_630,N_28751,N_25691);
nor UO_631 (O_631,N_28742,N_25608);
or UO_632 (O_632,N_24293,N_24825);
or UO_633 (O_633,N_26418,N_28502);
nand UO_634 (O_634,N_25917,N_24803);
and UO_635 (O_635,N_25730,N_24613);
xnor UO_636 (O_636,N_28362,N_25236);
and UO_637 (O_637,N_28388,N_28772);
or UO_638 (O_638,N_27923,N_29838);
and UO_639 (O_639,N_27733,N_28937);
nor UO_640 (O_640,N_28521,N_28016);
nor UO_641 (O_641,N_29911,N_27943);
xor UO_642 (O_642,N_25639,N_26271);
nor UO_643 (O_643,N_27910,N_27148);
nor UO_644 (O_644,N_24279,N_25533);
nor UO_645 (O_645,N_25358,N_28566);
and UO_646 (O_646,N_26122,N_25589);
nand UO_647 (O_647,N_25936,N_26389);
and UO_648 (O_648,N_26654,N_25073);
nor UO_649 (O_649,N_28056,N_29620);
or UO_650 (O_650,N_28359,N_24262);
xnor UO_651 (O_651,N_24785,N_29799);
xor UO_652 (O_652,N_28659,N_24151);
xnor UO_653 (O_653,N_27266,N_28741);
nand UO_654 (O_654,N_26929,N_27408);
and UO_655 (O_655,N_29039,N_29856);
nand UO_656 (O_656,N_24710,N_24235);
and UO_657 (O_657,N_24068,N_27708);
and UO_658 (O_658,N_27265,N_27710);
and UO_659 (O_659,N_28180,N_28398);
nor UO_660 (O_660,N_29441,N_27118);
or UO_661 (O_661,N_29738,N_24359);
xnor UO_662 (O_662,N_27675,N_25738);
nand UO_663 (O_663,N_24438,N_25212);
or UO_664 (O_664,N_29394,N_24988);
xnor UO_665 (O_665,N_24220,N_28033);
nand UO_666 (O_666,N_24708,N_26829);
xnor UO_667 (O_667,N_29238,N_28895);
or UO_668 (O_668,N_25074,N_28539);
or UO_669 (O_669,N_25516,N_25777);
nor UO_670 (O_670,N_27865,N_27738);
xor UO_671 (O_671,N_26311,N_24908);
xor UO_672 (O_672,N_26168,N_27250);
nor UO_673 (O_673,N_25966,N_25118);
and UO_674 (O_674,N_24772,N_25681);
and UO_675 (O_675,N_24790,N_28796);
nor UO_676 (O_676,N_26384,N_27718);
xnor UO_677 (O_677,N_25537,N_25419);
nand UO_678 (O_678,N_26136,N_25325);
and UO_679 (O_679,N_28720,N_29670);
or UO_680 (O_680,N_25821,N_25720);
nor UO_681 (O_681,N_27905,N_24736);
nor UO_682 (O_682,N_26499,N_29647);
and UO_683 (O_683,N_28678,N_28988);
or UO_684 (O_684,N_26519,N_27171);
nor UO_685 (O_685,N_25999,N_26276);
nor UO_686 (O_686,N_29933,N_25932);
xnor UO_687 (O_687,N_25356,N_24324);
and UO_688 (O_688,N_25390,N_27740);
and UO_689 (O_689,N_24969,N_25517);
or UO_690 (O_690,N_27766,N_29944);
and UO_691 (O_691,N_29167,N_25835);
nand UO_692 (O_692,N_25377,N_26146);
xnor UO_693 (O_693,N_26382,N_26426);
nor UO_694 (O_694,N_26608,N_29889);
or UO_695 (O_695,N_24465,N_29292);
xor UO_696 (O_696,N_28740,N_24622);
nand UO_697 (O_697,N_25327,N_27249);
nor UO_698 (O_698,N_28247,N_29632);
and UO_699 (O_699,N_26398,N_29357);
or UO_700 (O_700,N_24197,N_26142);
nand UO_701 (O_701,N_28165,N_28196);
or UO_702 (O_702,N_28761,N_28337);
or UO_703 (O_703,N_29916,N_29360);
nor UO_704 (O_704,N_25104,N_24504);
and UO_705 (O_705,N_27463,N_28839);
xnor UO_706 (O_706,N_27482,N_27461);
or UO_707 (O_707,N_25941,N_26823);
or UO_708 (O_708,N_26644,N_24588);
xnor UO_709 (O_709,N_29831,N_25189);
nor UO_710 (O_710,N_29951,N_28923);
nor UO_711 (O_711,N_27446,N_24389);
and UO_712 (O_712,N_27391,N_25740);
xor UO_713 (O_713,N_29503,N_29424);
xor UO_714 (O_714,N_29798,N_25774);
xor UO_715 (O_715,N_25878,N_24455);
xor UO_716 (O_716,N_27017,N_25350);
nand UO_717 (O_717,N_27706,N_28759);
nand UO_718 (O_718,N_26761,N_29259);
and UO_719 (O_719,N_29073,N_29791);
nand UO_720 (O_720,N_26253,N_24883);
nand UO_721 (O_721,N_27370,N_24373);
nand UO_722 (O_722,N_26110,N_27469);
nand UO_723 (O_723,N_26945,N_26505);
or UO_724 (O_724,N_27041,N_25911);
or UO_725 (O_725,N_28214,N_25451);
nand UO_726 (O_726,N_27860,N_28093);
and UO_727 (O_727,N_28750,N_25106);
and UO_728 (O_728,N_26975,N_28544);
xnor UO_729 (O_729,N_28982,N_24185);
xor UO_730 (O_730,N_26066,N_28843);
xor UO_731 (O_731,N_24829,N_27951);
or UO_732 (O_732,N_27418,N_27214);
nor UO_733 (O_733,N_28334,N_28764);
or UO_734 (O_734,N_24053,N_29256);
or UO_735 (O_735,N_28338,N_25645);
and UO_736 (O_736,N_26764,N_25113);
nor UO_737 (O_737,N_25131,N_29644);
or UO_738 (O_738,N_24826,N_26867);
nand UO_739 (O_739,N_29740,N_28305);
and UO_740 (O_740,N_29041,N_27818);
xor UO_741 (O_741,N_29652,N_29212);
nor UO_742 (O_742,N_25797,N_26845);
and UO_743 (O_743,N_24641,N_26408);
and UO_744 (O_744,N_26341,N_24040);
nand UO_745 (O_745,N_29578,N_24679);
and UO_746 (O_746,N_25574,N_26619);
xnor UO_747 (O_747,N_29627,N_28299);
nor UO_748 (O_748,N_27199,N_27545);
and UO_749 (O_749,N_25886,N_28492);
and UO_750 (O_750,N_24213,N_28930);
and UO_751 (O_751,N_28677,N_29035);
nor UO_752 (O_752,N_28596,N_24870);
nor UO_753 (O_753,N_24295,N_29112);
nor UO_754 (O_754,N_29950,N_27861);
xor UO_755 (O_755,N_27914,N_24992);
nor UO_756 (O_756,N_24955,N_24484);
xnor UO_757 (O_757,N_29629,N_29493);
nand UO_758 (O_758,N_24201,N_28948);
and UO_759 (O_759,N_28643,N_27653);
nand UO_760 (O_760,N_27882,N_29049);
nand UO_761 (O_761,N_24687,N_25648);
nand UO_762 (O_762,N_26946,N_28077);
and UO_763 (O_763,N_26497,N_25933);
nor UO_764 (O_764,N_27605,N_27313);
nand UO_765 (O_765,N_27650,N_25634);
nand UO_766 (O_766,N_26939,N_25611);
nand UO_767 (O_767,N_26344,N_28046);
or UO_768 (O_768,N_29464,N_27722);
or UO_769 (O_769,N_28646,N_26463);
or UO_770 (O_770,N_25757,N_28281);
or UO_771 (O_771,N_25616,N_24017);
or UO_772 (O_772,N_27150,N_28401);
nand UO_773 (O_773,N_29336,N_28685);
xnor UO_774 (O_774,N_26860,N_29990);
or UO_775 (O_775,N_27627,N_25148);
xor UO_776 (O_776,N_29975,N_28991);
or UO_777 (O_777,N_24378,N_28129);
or UO_778 (O_778,N_26282,N_26612);
nand UO_779 (O_779,N_26421,N_28709);
or UO_780 (O_780,N_25141,N_28660);
nand UO_781 (O_781,N_25764,N_28032);
or UO_782 (O_782,N_27533,N_26633);
or UO_783 (O_783,N_28273,N_28513);
xnor UO_784 (O_784,N_29515,N_27810);
or UO_785 (O_785,N_27068,N_26016);
xor UO_786 (O_786,N_28219,N_28382);
nor UO_787 (O_787,N_25180,N_25998);
nand UO_788 (O_788,N_25871,N_24648);
nor UO_789 (O_789,N_26001,N_26862);
and UO_790 (O_790,N_27661,N_27713);
and UO_791 (O_791,N_26655,N_25784);
xor UO_792 (O_792,N_27222,N_25534);
and UO_793 (O_793,N_26400,N_27714);
xnor UO_794 (O_794,N_27940,N_26566);
nand UO_795 (O_795,N_26085,N_26781);
and UO_796 (O_796,N_25114,N_27386);
nor UO_797 (O_797,N_29807,N_27688);
nand UO_798 (O_798,N_28924,N_24707);
nand UO_799 (O_799,N_27464,N_26780);
nor UO_800 (O_800,N_27457,N_28583);
nand UO_801 (O_801,N_28953,N_24316);
xnor UO_802 (O_802,N_29705,N_26580);
or UO_803 (O_803,N_26968,N_28080);
or UO_804 (O_804,N_28031,N_24871);
nor UO_805 (O_805,N_28436,N_29980);
xnor UO_806 (O_806,N_25109,N_24129);
xor UO_807 (O_807,N_29157,N_24474);
nor UO_808 (O_808,N_24865,N_29747);
nor UO_809 (O_809,N_29095,N_24782);
and UO_810 (O_810,N_27579,N_28125);
or UO_811 (O_811,N_25416,N_24817);
nor UO_812 (O_812,N_25976,N_28625);
nor UO_813 (O_813,N_24285,N_24441);
nor UO_814 (O_814,N_27690,N_26534);
nor UO_815 (O_815,N_24996,N_28541);
and UO_816 (O_816,N_28822,N_25891);
nand UO_817 (O_817,N_26391,N_26490);
nor UO_818 (O_818,N_24662,N_26812);
nand UO_819 (O_819,N_25044,N_26727);
and UO_820 (O_820,N_28821,N_28867);
and UO_821 (O_821,N_26279,N_24253);
nor UO_822 (O_822,N_26599,N_24044);
or UO_823 (O_823,N_27515,N_29897);
and UO_824 (O_824,N_29958,N_25294);
and UO_825 (O_825,N_28328,N_29927);
nand UO_826 (O_826,N_29205,N_28864);
or UO_827 (O_827,N_27907,N_26523);
nand UO_828 (O_828,N_25840,N_28494);
nor UO_829 (O_829,N_27895,N_26069);
or UO_830 (O_830,N_28295,N_27206);
nand UO_831 (O_831,N_28893,N_26409);
or UO_832 (O_832,N_29643,N_24824);
nor UO_833 (O_833,N_29452,N_25664);
or UO_834 (O_834,N_27611,N_29304);
xor UO_835 (O_835,N_25647,N_24417);
or UO_836 (O_836,N_25270,N_26586);
nor UO_837 (O_837,N_27325,N_28253);
nand UO_838 (O_838,N_28456,N_26491);
nor UO_839 (O_839,N_29380,N_27476);
nor UO_840 (O_840,N_26979,N_27692);
nor UO_841 (O_841,N_26796,N_25614);
xnor UO_842 (O_842,N_28221,N_28036);
xnor UO_843 (O_843,N_29845,N_29038);
nand UO_844 (O_844,N_26901,N_25266);
nor UO_845 (O_845,N_28342,N_29057);
and UO_846 (O_846,N_29568,N_29254);
nand UO_847 (O_847,N_27500,N_28611);
xor UO_848 (O_848,N_26920,N_27433);
xor UO_849 (O_849,N_28284,N_24916);
or UO_850 (O_850,N_29244,N_25934);
nor UO_851 (O_851,N_26387,N_24203);
or UO_852 (O_852,N_24257,N_28134);
or UO_853 (O_853,N_28373,N_25054);
nand UO_854 (O_854,N_27615,N_26702);
and UO_855 (O_855,N_24632,N_28038);
or UO_856 (O_856,N_27811,N_25045);
and UO_857 (O_857,N_29570,N_25842);
xor UO_858 (O_858,N_26370,N_28599);
nand UO_859 (O_859,N_29278,N_27357);
xnor UO_860 (O_860,N_29490,N_25803);
or UO_861 (O_861,N_25464,N_25226);
or UO_862 (O_862,N_25919,N_27462);
and UO_863 (O_863,N_27454,N_29624);
or UO_864 (O_864,N_25583,N_24743);
and UO_865 (O_865,N_27746,N_27868);
nand UO_866 (O_866,N_24760,N_25722);
and UO_867 (O_867,N_28831,N_29046);
nand UO_868 (O_868,N_24120,N_28443);
nand UO_869 (O_869,N_26063,N_27191);
nor UO_870 (O_870,N_29745,N_25043);
or UO_871 (O_871,N_24904,N_28245);
xnor UO_872 (O_872,N_25654,N_27909);
xnor UO_873 (O_873,N_25815,N_25610);
and UO_874 (O_874,N_24016,N_27351);
and UO_875 (O_875,N_24628,N_29641);
and UO_876 (O_876,N_29127,N_25622);
and UO_877 (O_877,N_28896,N_26533);
and UO_878 (O_878,N_26903,N_24127);
nand UO_879 (O_879,N_25458,N_29403);
and UO_880 (O_880,N_28055,N_29734);
nor UO_881 (O_881,N_27149,N_25861);
and UO_882 (O_882,N_24724,N_25905);
nand UO_883 (O_883,N_27651,N_27541);
nand UO_884 (O_884,N_24742,N_26836);
xor UO_885 (O_885,N_28612,N_25203);
nand UO_886 (O_886,N_28076,N_25262);
and UO_887 (O_887,N_25513,N_29808);
nand UO_888 (O_888,N_24406,N_29473);
or UO_889 (O_889,N_28085,N_27215);
nor UO_890 (O_890,N_25016,N_29923);
xor UO_891 (O_891,N_29234,N_24810);
and UO_892 (O_892,N_27731,N_25830);
xnor UO_893 (O_893,N_27739,N_24240);
nand UO_894 (O_894,N_28099,N_26321);
or UO_895 (O_895,N_24394,N_28695);
or UO_896 (O_896,N_28488,N_24050);
xor UO_897 (O_897,N_29466,N_25502);
nor UO_898 (O_898,N_26774,N_29935);
nand UO_899 (O_899,N_25711,N_28424);
nand UO_900 (O_900,N_24049,N_24859);
and UO_901 (O_901,N_27333,N_24343);
or UO_902 (O_902,N_27836,N_28081);
and UO_903 (O_903,N_25178,N_28182);
or UO_904 (O_904,N_27309,N_27194);
and UO_905 (O_905,N_29069,N_26105);
nand UO_906 (O_906,N_25052,N_27256);
or UO_907 (O_907,N_27697,N_27537);
nand UO_908 (O_908,N_24327,N_24336);
nor UO_909 (O_909,N_29827,N_26008);
or UO_910 (O_910,N_24873,N_27335);
or UO_911 (O_911,N_25196,N_24496);
or UO_912 (O_912,N_28682,N_27843);
nor UO_913 (O_913,N_26717,N_29900);
or UO_914 (O_914,N_27518,N_26522);
or UO_915 (O_915,N_28900,N_28089);
nor UO_916 (O_916,N_26625,N_24658);
and UO_917 (O_917,N_28164,N_29500);
or UO_918 (O_918,N_26994,N_28971);
and UO_919 (O_919,N_28518,N_24019);
or UO_920 (O_920,N_25714,N_27066);
and UO_921 (O_921,N_29960,N_25923);
nor UO_922 (O_922,N_27485,N_25865);
nor UO_923 (O_923,N_28786,N_27318);
nand UO_924 (O_924,N_24006,N_28882);
xor UO_925 (O_925,N_26928,N_24576);
nand UO_926 (O_926,N_24162,N_25721);
xnor UO_927 (O_927,N_29540,N_28474);
and UO_928 (O_928,N_28955,N_29457);
and UO_929 (O_929,N_27287,N_26828);
xnor UO_930 (O_930,N_24351,N_24691);
nor UO_931 (O_931,N_24566,N_29429);
and UO_932 (O_932,N_26155,N_29164);
nand UO_933 (O_933,N_26993,N_29665);
xor UO_934 (O_934,N_24339,N_27460);
nor UO_935 (O_935,N_25552,N_27920);
nor UO_936 (O_936,N_28691,N_25473);
nor UO_937 (O_937,N_27456,N_24026);
and UO_938 (O_938,N_26454,N_26334);
nand UO_939 (O_939,N_29132,N_24247);
xor UO_940 (O_940,N_27108,N_24191);
nor UO_941 (O_941,N_27262,N_26143);
and UO_942 (O_942,N_25158,N_28684);
or UO_943 (O_943,N_28572,N_29248);
or UO_944 (O_944,N_26187,N_24464);
nor UO_945 (O_945,N_29064,N_24615);
or UO_946 (O_946,N_25477,N_29148);
xnor UO_947 (O_947,N_24156,N_24550);
or UO_948 (O_948,N_27093,N_24557);
or UO_949 (O_949,N_27270,N_24344);
or UO_950 (O_950,N_27542,N_26846);
and UO_951 (O_951,N_25213,N_27874);
nand UO_952 (O_952,N_24052,N_25779);
and UO_953 (O_953,N_28983,N_29219);
nor UO_954 (O_954,N_29416,N_28312);
xnor UO_955 (O_955,N_29854,N_24762);
xnor UO_956 (O_956,N_25581,N_24991);
nand UO_957 (O_957,N_28369,N_29801);
nand UO_958 (O_958,N_24200,N_28368);
nand UO_959 (O_959,N_29325,N_26237);
xor UO_960 (O_960,N_25136,N_26178);
nor UO_961 (O_961,N_24678,N_29341);
or UO_962 (O_962,N_25820,N_27575);
xor UO_963 (O_963,N_26407,N_27103);
nor UO_964 (O_964,N_26852,N_29396);
or UO_965 (O_965,N_26551,N_28242);
nor UO_966 (O_966,N_27104,N_24117);
or UO_967 (O_967,N_27496,N_24090);
nor UO_968 (O_968,N_26622,N_27568);
and UO_969 (O_969,N_25897,N_29356);
nand UO_970 (O_970,N_29196,N_26379);
nand UO_971 (O_971,N_29201,N_24981);
and UO_972 (O_972,N_24745,N_24813);
nand UO_973 (O_973,N_27227,N_27085);
xnor UO_974 (O_974,N_29855,N_26636);
nor UO_975 (O_975,N_24403,N_25197);
or UO_976 (O_976,N_26054,N_26429);
xor UO_977 (O_977,N_26995,N_27574);
nand UO_978 (O_978,N_26090,N_28294);
xnor UO_979 (O_979,N_27536,N_28235);
or UO_980 (O_980,N_25105,N_26677);
nand UO_981 (O_981,N_26163,N_24317);
nor UO_982 (O_982,N_24233,N_24855);
nand UO_983 (O_983,N_27830,N_25531);
and UO_984 (O_984,N_26043,N_26940);
xnor UO_985 (O_985,N_26479,N_27055);
or UO_986 (O_986,N_26177,N_29239);
or UO_987 (O_987,N_28997,N_26338);
nor UO_988 (O_988,N_26999,N_25857);
and UO_989 (O_989,N_29604,N_27245);
nand UO_990 (O_990,N_25304,N_26356);
and UO_991 (O_991,N_24379,N_27236);
xor UO_992 (O_992,N_27789,N_24655);
or UO_993 (O_993,N_28545,N_26473);
nand UO_994 (O_994,N_29945,N_28892);
nand UO_995 (O_995,N_28404,N_25974);
or UO_996 (O_996,N_29758,N_26917);
nor UO_997 (O_997,N_26042,N_26153);
nand UO_998 (O_998,N_27288,N_25135);
nand UO_999 (O_999,N_26367,N_29690);
nand UO_1000 (O_1000,N_28788,N_27241);
xor UO_1001 (O_1001,N_27548,N_25805);
or UO_1002 (O_1002,N_26469,N_25554);
and UO_1003 (O_1003,N_24937,N_29372);
nor UO_1004 (O_1004,N_25732,N_24823);
xnor UO_1005 (O_1005,N_27851,N_24335);
xnor UO_1006 (O_1006,N_27704,N_27684);
nand UO_1007 (O_1007,N_28167,N_29209);
xnor UO_1008 (O_1008,N_27938,N_24282);
xnor UO_1009 (O_1009,N_27414,N_26035);
or UO_1010 (O_1010,N_29020,N_29521);
nand UO_1011 (O_1011,N_25110,N_26689);
or UO_1012 (O_1012,N_27365,N_29459);
nor UO_1013 (O_1013,N_29009,N_27311);
xnor UO_1014 (O_1014,N_29181,N_24423);
nand UO_1015 (O_1015,N_25260,N_25363);
and UO_1016 (O_1016,N_28824,N_25409);
nor UO_1017 (O_1017,N_24013,N_27061);
nand UO_1018 (O_1018,N_24020,N_24647);
xnor UO_1019 (O_1019,N_24838,N_29715);
xor UO_1020 (O_1020,N_29577,N_29163);
or UO_1021 (O_1021,N_25509,N_24413);
and UO_1022 (O_1022,N_29555,N_27302);
nand UO_1023 (O_1023,N_27707,N_24552);
xnor UO_1024 (O_1024,N_24578,N_25276);
xor UO_1025 (O_1025,N_28717,N_27142);
and UO_1026 (O_1026,N_27522,N_27165);
xnor UO_1027 (O_1027,N_26358,N_28651);
or UO_1028 (O_1028,N_26392,N_29543);
nor UO_1029 (O_1029,N_24897,N_27013);
nor UO_1030 (O_1030,N_27587,N_25122);
nand UO_1031 (O_1031,N_24545,N_26893);
nor UO_1032 (O_1032,N_28185,N_29388);
or UO_1033 (O_1033,N_26648,N_28602);
nor UO_1034 (O_1034,N_29514,N_25238);
and UO_1035 (O_1035,N_27437,N_27243);
nand UO_1036 (O_1036,N_27403,N_25693);
xnor UO_1037 (O_1037,N_25663,N_27559);
nor UO_1038 (O_1038,N_24635,N_25429);
and UO_1039 (O_1039,N_24230,N_25065);
nand UO_1040 (O_1040,N_26191,N_25279);
or UO_1041 (O_1041,N_24654,N_27415);
nor UO_1042 (O_1042,N_25493,N_24646);
nor UO_1043 (O_1043,N_27131,N_25718);
or UO_1044 (O_1044,N_25541,N_27292);
or UO_1045 (O_1045,N_29857,N_24392);
nor UO_1046 (O_1046,N_25847,N_29171);
xor UO_1047 (O_1047,N_29818,N_28730);
nand UO_1048 (O_1048,N_26596,N_27002);
and UO_1049 (O_1049,N_26109,N_26451);
nor UO_1050 (O_1050,N_26324,N_29413);
or UO_1051 (O_1051,N_25928,N_29494);
or UO_1052 (O_1052,N_25187,N_27747);
or UO_1053 (O_1053,N_24723,N_26047);
nor UO_1054 (O_1054,N_28203,N_29225);
xor UO_1055 (O_1055,N_29218,N_25641);
or UO_1056 (O_1056,N_25003,N_25255);
nand UO_1057 (O_1057,N_25403,N_27375);
nor UO_1058 (O_1058,N_26510,N_29307);
nand UO_1059 (O_1059,N_26731,N_26675);
or UO_1060 (O_1060,N_29586,N_29443);
nor UO_1061 (O_1061,N_26028,N_29699);
or UO_1062 (O_1062,N_25813,N_28609);
or UO_1063 (O_1063,N_25822,N_29661);
nor UO_1064 (O_1064,N_26489,N_26938);
and UO_1065 (O_1065,N_24515,N_25229);
xnor UO_1066 (O_1066,N_27734,N_25729);
nor UO_1067 (O_1067,N_29076,N_24066);
or UO_1068 (O_1068,N_28458,N_24998);
and UO_1069 (O_1069,N_28144,N_24667);
or UO_1070 (O_1070,N_25281,N_27264);
or UO_1071 (O_1071,N_27750,N_26777);
nor UO_1072 (O_1072,N_26592,N_26322);
or UO_1073 (O_1073,N_29835,N_28593);
and UO_1074 (O_1074,N_27989,N_27968);
xnor UO_1075 (O_1075,N_26663,N_26623);
xor UO_1076 (O_1076,N_28756,N_24045);
or UO_1077 (O_1077,N_26019,N_28229);
or UO_1078 (O_1078,N_25427,N_28116);
xnor UO_1079 (O_1079,N_24940,N_27402);
nor UO_1080 (O_1080,N_29363,N_25954);
nor UO_1081 (O_1081,N_24014,N_27005);
xor UO_1082 (O_1082,N_28808,N_28130);
and UO_1083 (O_1083,N_26807,N_27981);
or UO_1084 (O_1084,N_29344,N_27101);
or UO_1085 (O_1085,N_24807,N_24242);
nand UO_1086 (O_1086,N_28634,N_28771);
nor UO_1087 (O_1087,N_28664,N_24497);
and UO_1088 (O_1088,N_24963,N_25237);
nor UO_1089 (O_1089,N_26834,N_26205);
xnor UO_1090 (O_1090,N_26258,N_26034);
nor UO_1091 (O_1091,N_24333,N_25507);
xnor UO_1092 (O_1092,N_29903,N_24863);
xnor UO_1093 (O_1093,N_27986,N_26719);
xor UO_1094 (O_1094,N_24091,N_25184);
xor UO_1095 (O_1095,N_29375,N_25461);
and UO_1096 (O_1096,N_25800,N_24218);
xor UO_1097 (O_1097,N_25318,N_24530);
nor UO_1098 (O_1098,N_28151,N_28254);
or UO_1099 (O_1099,N_28811,N_26817);
xnor UO_1100 (O_1100,N_28155,N_29190);
nand UO_1101 (O_1101,N_25990,N_28272);
nor UO_1102 (O_1102,N_25247,N_24905);
and UO_1103 (O_1103,N_28916,N_25973);
nor UO_1104 (O_1104,N_27687,N_26508);
or UO_1105 (O_1105,N_27046,N_29700);
nand UO_1106 (O_1106,N_26884,N_29079);
and UO_1107 (O_1107,N_24114,N_29736);
nand UO_1108 (O_1108,N_28287,N_24854);
or UO_1109 (O_1109,N_27601,N_29756);
and UO_1110 (O_1110,N_25096,N_27879);
or UO_1111 (O_1111,N_29531,N_26032);
and UO_1112 (O_1112,N_28850,N_26386);
and UO_1113 (O_1113,N_24443,N_29484);
or UO_1114 (O_1114,N_28421,N_28860);
xor UO_1115 (O_1115,N_29969,N_26649);
xnor UO_1116 (O_1116,N_27539,N_27368);
xnor UO_1117 (O_1117,N_29886,N_28345);
or UO_1118 (O_1118,N_28184,N_28790);
nand UO_1119 (O_1119,N_24975,N_28686);
nand UO_1120 (O_1120,N_26004,N_29277);
xor UO_1121 (O_1121,N_24711,N_26336);
xnor UO_1122 (O_1122,N_26212,N_29240);
and UO_1123 (O_1123,N_26624,N_28590);
nand UO_1124 (O_1124,N_25164,N_26083);
and UO_1125 (O_1125,N_28327,N_28423);
nand UO_1126 (O_1126,N_25628,N_27444);
nand UO_1127 (O_1127,N_25632,N_26811);
or UO_1128 (O_1128,N_25015,N_28355);
or UO_1129 (O_1129,N_28286,N_27459);
nor UO_1130 (O_1130,N_27857,N_24172);
nand UO_1131 (O_1131,N_24350,N_26306);
xnor UO_1132 (O_1132,N_26315,N_24190);
and UO_1133 (O_1133,N_26978,N_24122);
or UO_1134 (O_1134,N_24670,N_28561);
nor UO_1135 (O_1135,N_25743,N_27573);
and UO_1136 (O_1136,N_25945,N_24187);
and UO_1137 (O_1137,N_27529,N_29123);
xor UO_1138 (O_1138,N_28607,N_29018);
nor UO_1139 (O_1139,N_28012,N_24931);
xor UO_1140 (O_1140,N_27617,N_26487);
nand UO_1141 (O_1141,N_27480,N_29957);
or UO_1142 (O_1142,N_28511,N_29949);
xnor UO_1143 (O_1143,N_26158,N_27822);
and UO_1144 (O_1144,N_26416,N_26726);
nand UO_1145 (O_1145,N_29509,N_25652);
nand UO_1146 (O_1146,N_29836,N_28696);
or UO_1147 (O_1147,N_25324,N_25263);
and UO_1148 (O_1148,N_24734,N_24180);
nor UO_1149 (O_1149,N_29051,N_27555);
nand UO_1150 (O_1150,N_26278,N_28001);
xor UO_1151 (O_1151,N_25284,N_28890);
nand UO_1152 (O_1152,N_29833,N_25095);
and UO_1153 (O_1153,N_26280,N_28483);
or UO_1154 (O_1154,N_27797,N_27726);
and UO_1155 (O_1155,N_28689,N_26373);
nand UO_1156 (O_1156,N_24360,N_27924);
and UO_1157 (O_1157,N_27960,N_26152);
or UO_1158 (O_1158,N_29523,N_28018);
and UO_1159 (O_1159,N_24733,N_24700);
nand UO_1160 (O_1160,N_29096,N_24405);
or UO_1161 (O_1161,N_26395,N_24765);
nand UO_1162 (O_1162,N_25062,N_28595);
nor UO_1163 (O_1163,N_27721,N_28744);
and UO_1164 (O_1164,N_28322,N_25946);
nor UO_1165 (O_1165,N_29472,N_29210);
xor UO_1166 (O_1166,N_25100,N_28714);
nand UO_1167 (O_1167,N_28403,N_29216);
or UO_1168 (O_1168,N_29172,N_24202);
nand UO_1169 (O_1169,N_25899,N_24675);
nand UO_1170 (O_1170,N_25665,N_25575);
or UO_1171 (O_1171,N_25348,N_26771);
xor UO_1172 (O_1172,N_28068,N_25770);
or UO_1173 (O_1173,N_27547,N_26073);
nor UO_1174 (O_1174,N_29371,N_24637);
nor UO_1175 (O_1175,N_25860,N_28140);
and UO_1176 (O_1176,N_29335,N_27658);
or UO_1177 (O_1177,N_24890,N_29968);
nor UO_1178 (O_1178,N_29548,N_25957);
xnor UO_1179 (O_1179,N_25873,N_26161);
or UO_1180 (O_1180,N_24145,N_24095);
nand UO_1181 (O_1181,N_28367,N_29600);
nor UO_1182 (O_1182,N_25112,N_29122);
nand UO_1183 (O_1183,N_29817,N_25248);
xnor UO_1184 (O_1184,N_26583,N_29686);
nor UO_1185 (O_1185,N_26869,N_24858);
nand UO_1186 (O_1186,N_27636,N_27374);
xnor UO_1187 (O_1187,N_29599,N_26536);
and UO_1188 (O_1188,N_24380,N_25217);
or UO_1189 (O_1189,N_26095,N_29385);
nor UO_1190 (O_1190,N_25989,N_29138);
xnor UO_1191 (O_1191,N_25407,N_26100);
nand UO_1192 (O_1192,N_24369,N_26340);
xnor UO_1193 (O_1193,N_26537,N_27777);
nor UO_1194 (O_1194,N_25469,N_25825);
and UO_1195 (O_1195,N_27024,N_28530);
xnor UO_1196 (O_1196,N_26397,N_24570);
xnor UO_1197 (O_1197,N_29712,N_28954);
or UO_1198 (O_1198,N_24234,N_29560);
xnor UO_1199 (O_1199,N_29840,N_25695);
nand UO_1200 (O_1200,N_28049,N_29793);
or UO_1201 (O_1201,N_25129,N_29735);
nor UO_1202 (O_1202,N_28967,N_24786);
xnor UO_1203 (O_1203,N_25765,N_26188);
nand UO_1204 (O_1204,N_28266,N_29534);
xor UO_1205 (O_1205,N_29552,N_25565);
and UO_1206 (O_1206,N_25837,N_24410);
xnor UO_1207 (O_1207,N_25773,N_28153);
and UO_1208 (O_1208,N_28876,N_29442);
nor UO_1209 (O_1209,N_25530,N_24952);
and UO_1210 (O_1210,N_28627,N_27546);
nor UO_1211 (O_1211,N_28652,N_25994);
nand UO_1212 (O_1212,N_27187,N_27856);
nor UO_1213 (O_1213,N_28992,N_27520);
nor UO_1214 (O_1214,N_25201,N_26509);
or UO_1215 (O_1215,N_29684,N_26131);
nor UO_1216 (O_1216,N_29680,N_29942);
nor UO_1217 (O_1217,N_24491,N_26352);
xor UO_1218 (O_1218,N_24442,N_25549);
xnor UO_1219 (O_1219,N_25585,N_26233);
and UO_1220 (O_1220,N_26130,N_24651);
or UO_1221 (O_1221,N_28931,N_28143);
xor UO_1222 (O_1222,N_25088,N_24217);
and UO_1223 (O_1223,N_28122,N_25629);
or UO_1224 (O_1224,N_28616,N_28479);
xor UO_1225 (O_1225,N_27820,N_28298);
nor UO_1226 (O_1226,N_28732,N_29183);
xnor UO_1227 (O_1227,N_28179,N_24951);
or UO_1228 (O_1228,N_27593,N_26316);
and UO_1229 (O_1229,N_24119,N_24881);
and UO_1230 (O_1230,N_28701,N_28532);
and UO_1231 (O_1231,N_29930,N_28385);
nor UO_1232 (O_1232,N_28340,N_27901);
nor UO_1233 (O_1233,N_24325,N_24420);
nand UO_1234 (O_1234,N_27846,N_26037);
nor UO_1235 (O_1235,N_24179,N_24184);
and UO_1236 (O_1236,N_29321,N_25661);
xor UO_1237 (O_1237,N_24449,N_28542);
xnor UO_1238 (O_1238,N_28161,N_27478);
and UO_1239 (O_1239,N_25832,N_27727);
and UO_1240 (O_1240,N_29726,N_29447);
or UO_1241 (O_1241,N_24396,N_27664);
xnor UO_1242 (O_1242,N_26676,N_29695);
and UO_1243 (O_1243,N_27928,N_25746);
nor UO_1244 (O_1244,N_24748,N_25218);
and UO_1245 (O_1245,N_28480,N_28226);
xor UO_1246 (O_1246,N_26147,N_26888);
nand UO_1247 (O_1247,N_27110,N_28205);
nand UO_1248 (O_1248,N_25598,N_26983);
nand UO_1249 (O_1249,N_24064,N_29575);
nand UO_1250 (O_1250,N_29337,N_28379);
xnor UO_1251 (O_1251,N_26866,N_24148);
nand UO_1252 (O_1252,N_28079,N_25321);
or UO_1253 (O_1253,N_24444,N_27091);
and UO_1254 (O_1254,N_24756,N_24788);
xor UO_1255 (O_1255,N_27581,N_26417);
nor UO_1256 (O_1256,N_25133,N_26214);
and UO_1257 (O_1257,N_26894,N_28673);
and UO_1258 (O_1258,N_26722,N_25498);
or UO_1259 (O_1259,N_24965,N_28639);
nor UO_1260 (O_1260,N_24596,N_25072);
nand UO_1261 (O_1261,N_25396,N_28467);
nor UO_1262 (O_1262,N_24245,N_28048);
or UO_1263 (O_1263,N_27012,N_25543);
nand UO_1264 (O_1264,N_27081,N_27048);
nand UO_1265 (O_1265,N_27490,N_25698);
nor UO_1266 (O_1266,N_27614,N_26040);
nand UO_1267 (O_1267,N_28738,N_28098);
nand UO_1268 (O_1268,N_25783,N_27230);
and UO_1269 (O_1269,N_28613,N_27534);
nor UO_1270 (O_1270,N_26987,N_29194);
nand UO_1271 (O_1271,N_27163,N_29202);
xor UO_1272 (O_1272,N_29235,N_28905);
or UO_1273 (O_1273,N_28393,N_28288);
and UO_1274 (O_1274,N_25089,N_29648);
or UO_1275 (O_1275,N_26332,N_27028);
or UO_1276 (O_1276,N_29650,N_27272);
nor UO_1277 (O_1277,N_26621,N_28223);
or UO_1278 (O_1278,N_25888,N_25250);
xor UO_1279 (O_1279,N_28973,N_27269);
nand UO_1280 (O_1280,N_28552,N_29458);
or UO_1281 (O_1281,N_27259,N_25841);
nor UO_1282 (O_1282,N_24725,N_27634);
xor UO_1283 (O_1283,N_27246,N_24527);
nand UO_1284 (O_1284,N_29619,N_29488);
xnor UO_1285 (O_1285,N_27848,N_25710);
and UO_1286 (O_1286,N_24828,N_26925);
nand UO_1287 (O_1287,N_28220,N_27755);
or UO_1288 (O_1288,N_25564,N_26951);
and UO_1289 (O_1289,N_28517,N_25603);
nor UO_1290 (O_1290,N_27696,N_29450);
xor UO_1291 (O_1291,N_24009,N_24454);
or UO_1292 (O_1292,N_25766,N_28588);
and UO_1293 (O_1293,N_27307,N_27026);
nor UO_1294 (O_1294,N_28465,N_29796);
or UO_1295 (O_1295,N_26436,N_26265);
nor UO_1296 (O_1296,N_29369,N_26645);
and UO_1297 (O_1297,N_26005,N_26724);
xnor UO_1298 (O_1298,N_24727,N_26262);
nor UO_1299 (O_1299,N_28070,N_24533);
nor UO_1300 (O_1300,N_29444,N_25036);
xor UO_1301 (O_1301,N_25633,N_26559);
nor UO_1302 (O_1302,N_24276,N_28177);
nand UO_1303 (O_1303,N_28996,N_29286);
xor UO_1304 (O_1304,N_28606,N_25444);
xor UO_1305 (O_1305,N_29067,N_24716);
and UO_1306 (O_1306,N_26801,N_29654);
xor UO_1307 (O_1307,N_29474,N_24015);
nor UO_1308 (O_1308,N_24248,N_29939);
or UO_1309 (O_1309,N_28979,N_26192);
nand UO_1310 (O_1310,N_24459,N_28505);
and UO_1311 (O_1311,N_24995,N_26411);
nor UO_1312 (O_1312,N_27498,N_24787);
and UO_1313 (O_1313,N_26159,N_25748);
or UO_1314 (O_1314,N_28999,N_28154);
or UO_1315 (O_1315,N_24925,N_24372);
xnor UO_1316 (O_1316,N_27530,N_25916);
and UO_1317 (O_1317,N_25455,N_29763);
nand UO_1318 (O_1318,N_28891,N_26074);
or UO_1319 (O_1319,N_25987,N_28282);
nor UO_1320 (O_1320,N_29287,N_25278);
and UO_1321 (O_1321,N_28535,N_26524);
xor UO_1322 (O_1322,N_28152,N_27247);
and UO_1323 (O_1323,N_24933,N_24294);
and UO_1324 (O_1324,N_29788,N_26478);
nand UO_1325 (O_1325,N_28006,N_26944);
nand UO_1326 (O_1326,N_27031,N_29320);
xor UO_1327 (O_1327,N_24842,N_24391);
xnor UO_1328 (O_1328,N_29931,N_27725);
or UO_1329 (O_1329,N_25988,N_29103);
xnor UO_1330 (O_1330,N_26715,N_28563);
nand UO_1331 (O_1331,N_28377,N_26495);
xnor UO_1332 (O_1332,N_29601,N_28199);
and UO_1333 (O_1333,N_29925,N_25290);
xor UO_1334 (O_1334,N_28936,N_26360);
nor UO_1335 (O_1335,N_27455,N_28516);
nand UO_1336 (O_1336,N_28405,N_24236);
nand UO_1337 (O_1337,N_25121,N_29386);
xnor UO_1338 (O_1338,N_29615,N_27655);
xor UO_1339 (O_1339,N_27791,N_29755);
nor UO_1340 (O_1340,N_27037,N_27580);
xnor UO_1341 (O_1341,N_26111,N_28430);
and UO_1342 (O_1342,N_25659,N_29691);
or UO_1343 (O_1343,N_29077,N_28998);
nor UO_1344 (O_1344,N_27556,N_29191);
xor UO_1345 (O_1345,N_24347,N_26245);
or UO_1346 (O_1346,N_24041,N_26955);
or UO_1347 (O_1347,N_28106,N_24277);
or UO_1348 (O_1348,N_29415,N_28073);
nand UO_1349 (O_1349,N_26851,N_26776);
nand UO_1350 (O_1350,N_26476,N_25542);
and UO_1351 (O_1351,N_29772,N_29677);
nand UO_1352 (O_1352,N_27705,N_29330);
or UO_1353 (O_1353,N_29334,N_26452);
xor UO_1354 (O_1354,N_27499,N_24461);
nand UO_1355 (O_1355,N_29593,N_27544);
nand UO_1356 (O_1356,N_27412,N_25086);
and UO_1357 (O_1357,N_28350,N_28249);
xor UO_1358 (O_1358,N_26107,N_28762);
xor UO_1359 (O_1359,N_27639,N_24163);
xnor UO_1360 (O_1360,N_24848,N_28021);
xor UO_1361 (O_1361,N_27372,N_27213);
xnor UO_1362 (O_1362,N_24600,N_26871);
or UO_1363 (O_1363,N_28361,N_25684);
and UO_1364 (O_1364,N_25024,N_29091);
xor UO_1365 (O_1365,N_26699,N_29019);
xnor UO_1366 (O_1366,N_27263,N_25310);
xor UO_1367 (O_1367,N_24047,N_28118);
and UO_1368 (O_1368,N_28202,N_25818);
nand UO_1369 (O_1369,N_26890,N_24563);
and UO_1370 (O_1370,N_24780,N_29814);
nand UO_1371 (O_1371,N_26030,N_24167);
or UO_1372 (O_1372,N_26837,N_25476);
or UO_1373 (O_1373,N_29991,N_29223);
or UO_1374 (O_1374,N_24911,N_24548);
or UO_1375 (O_1375,N_24761,N_29468);
or UO_1376 (O_1376,N_25607,N_24054);
and UO_1377 (O_1377,N_29134,N_24099);
and UO_1378 (O_1378,N_28422,N_25956);
xnor UO_1379 (O_1379,N_26449,N_26902);
nand UO_1380 (O_1380,N_26972,N_27812);
xnor UO_1381 (O_1381,N_28871,N_25500);
xor UO_1382 (O_1382,N_26996,N_26670);
nand UO_1383 (O_1383,N_27963,N_26115);
xor UO_1384 (O_1384,N_27059,N_25374);
xnor UO_1385 (O_1385,N_28094,N_29908);
nand UO_1386 (O_1386,N_29428,N_29153);
and UO_1387 (O_1387,N_24941,N_27804);
xor UO_1388 (O_1388,N_28885,N_26795);
or UO_1389 (O_1389,N_26068,N_24476);
or UO_1390 (O_1390,N_26401,N_26835);
and UO_1391 (O_1391,N_29882,N_26202);
xnor UO_1392 (O_1392,N_25771,N_25012);
and UO_1393 (O_1393,N_27927,N_26891);
and UO_1394 (O_1394,N_27467,N_27889);
nor UO_1395 (O_1395,N_28381,N_27014);
and UO_1396 (O_1396,N_24312,N_25872);
or UO_1397 (O_1397,N_25584,N_28064);
nor UO_1398 (O_1398,N_24966,N_29411);
nor UO_1399 (O_1399,N_28169,N_26128);
nand UO_1400 (O_1400,N_26768,N_28587);
xnor UO_1401 (O_1401,N_29773,N_26640);
or UO_1402 (O_1402,N_29410,N_25977);
nor UO_1403 (O_1403,N_28395,N_25563);
xor UO_1404 (O_1404,N_27785,N_29743);
nand UO_1405 (O_1405,N_28297,N_26980);
nor UO_1406 (O_1406,N_29730,N_27853);
xnor UO_1407 (O_1407,N_26458,N_26006);
nand UO_1408 (O_1408,N_24896,N_29367);
xnor UO_1409 (O_1409,N_29298,N_29795);
nor UO_1410 (O_1410,N_27527,N_26023);
nand UO_1411 (O_1411,N_27854,N_26179);
or UO_1412 (O_1412,N_25090,N_24164);
nor UO_1413 (O_1413,N_29723,N_24789);
nand UO_1414 (O_1414,N_29554,N_24341);
and UO_1415 (O_1415,N_24267,N_27392);
nand UO_1416 (O_1416,N_28767,N_24100);
xor UO_1417 (O_1417,N_25200,N_28366);
nor UO_1418 (O_1418,N_26219,N_27221);
or UO_1419 (O_1419,N_28777,N_25731);
nor UO_1420 (O_1420,N_24779,N_26970);
nand UO_1421 (O_1421,N_26716,N_27080);
nand UO_1422 (O_1422,N_26617,N_25597);
xnor UO_1423 (O_1423,N_28459,N_29200);
or UO_1424 (O_1424,N_26433,N_29888);
or UO_1425 (O_1425,N_28629,N_28562);
nand UO_1426 (O_1426,N_26967,N_25851);
nand UO_1427 (O_1427,N_27505,N_25384);
nor UO_1428 (O_1428,N_29674,N_25601);
and UO_1429 (O_1429,N_27237,N_28275);
or UO_1430 (O_1430,N_26595,N_24109);
nor UO_1431 (O_1431,N_28124,N_25850);
nand UO_1432 (O_1432,N_29226,N_29989);
xnor UO_1433 (O_1433,N_26402,N_26138);
xor UO_1434 (O_1434,N_26218,N_27992);
nand UO_1435 (O_1435,N_24260,N_29608);
nor UO_1436 (O_1436,N_24318,N_29762);
xnor UO_1437 (O_1437,N_27988,N_26687);
or UO_1438 (O_1438,N_27004,N_24308);
nor UO_1439 (O_1439,N_29326,N_26088);
or UO_1440 (O_1440,N_24836,N_29093);
xor UO_1441 (O_1441,N_26255,N_27875);
nand UO_1442 (O_1442,N_25336,N_27662);
or UO_1443 (O_1443,N_24239,N_27837);
xor UO_1444 (O_1444,N_29813,N_26952);
nor UO_1445 (O_1445,N_25028,N_25246);
and UO_1446 (O_1446,N_24083,N_25521);
xor UO_1447 (O_1447,N_24997,N_26563);
nor UO_1448 (O_1448,N_28040,N_25053);
nor UO_1449 (O_1449,N_29314,N_25487);
nand UO_1450 (O_1450,N_28865,N_24682);
and UO_1451 (O_1451,N_25466,N_26576);
nor UO_1452 (O_1452,N_28246,N_27034);
or UO_1453 (O_1453,N_25063,N_24001);
xor UO_1454 (O_1454,N_27197,N_27337);
xor UO_1455 (O_1455,N_25060,N_27752);
and UO_1456 (O_1456,N_29996,N_26662);
and UO_1457 (O_1457,N_24221,N_28944);
xnor UO_1458 (O_1458,N_25438,N_25315);
nor UO_1459 (O_1459,N_24516,N_28448);
and UO_1460 (O_1460,N_25655,N_28349);
nand UO_1461 (O_1461,N_24663,N_26430);
and UO_1462 (O_1462,N_28880,N_27814);
nand UO_1463 (O_1463,N_24495,N_26396);
nand UO_1464 (O_1464,N_24305,N_26525);
xnor UO_1465 (O_1465,N_24458,N_25373);
nand UO_1466 (O_1466,N_25606,N_25739);
or UO_1467 (O_1467,N_29063,N_28163);
and UO_1468 (O_1468,N_28454,N_29267);
xor UO_1469 (O_1469,N_26814,N_25526);
or UO_1470 (O_1470,N_25316,N_28801);
nor UO_1471 (O_1471,N_26703,N_26948);
xnor UO_1472 (O_1472,N_27212,N_28688);
or UO_1473 (O_1473,N_24876,N_28208);
nand UO_1474 (O_1474,N_29118,N_26971);
and UO_1475 (O_1475,N_25573,N_26858);
xnor UO_1476 (O_1476,N_28789,N_28088);
or UO_1477 (O_1477,N_27682,N_29026);
nand UO_1478 (O_1478,N_26247,N_29826);
xor UO_1479 (O_1479,N_24081,N_24676);
and UO_1480 (O_1480,N_24263,N_26150);
xor UO_1481 (O_1481,N_25864,N_28969);
or UO_1482 (O_1482,N_29790,N_25261);
xnor UO_1483 (O_1483,N_24580,N_28934);
and UO_1484 (O_1484,N_27152,N_28139);
nand UO_1485 (O_1485,N_27592,N_24604);
xnor UO_1486 (O_1486,N_27828,N_26366);
xor UO_1487 (O_1487,N_26868,N_28576);
nand UO_1488 (O_1488,N_29711,N_28490);
nand UO_1489 (O_1489,N_28654,N_29368);
nor UO_1490 (O_1490,N_29071,N_25510);
nor UO_1491 (O_1491,N_25737,N_24432);
nor UO_1492 (O_1492,N_27930,N_26518);
xor UO_1493 (O_1493,N_28601,N_26681);
or UO_1494 (O_1494,N_27526,N_28804);
nor UO_1495 (O_1495,N_24363,N_28037);
xnor UO_1496 (O_1496,N_25360,N_27010);
nor UO_1497 (O_1497,N_26369,N_29003);
or UO_1498 (O_1498,N_25570,N_24094);
nand UO_1499 (O_1499,N_24943,N_25854);
nand UO_1500 (O_1500,N_26708,N_29106);
nand UO_1501 (O_1501,N_24500,N_26618);
and UO_1502 (O_1502,N_24210,N_28724);
and UO_1503 (O_1503,N_29133,N_24770);
xor UO_1504 (O_1504,N_24737,N_25170);
xor UO_1505 (O_1505,N_27283,N_24493);
nand UO_1506 (O_1506,N_27944,N_25702);
or UO_1507 (O_1507,N_24353,N_29806);
nor UO_1508 (O_1508,N_27475,N_27834);
nand UO_1509 (O_1509,N_26017,N_28838);
xnor UO_1510 (O_1510,N_29852,N_26140);
and UO_1511 (O_1511,N_24401,N_28901);
nand UO_1512 (O_1512,N_28277,N_29671);
xor UO_1513 (O_1513,N_25485,N_26089);
or UO_1514 (O_1514,N_29637,N_26613);
and UO_1515 (O_1515,N_28175,N_27516);
and UO_1516 (O_1516,N_26674,N_25750);
nor UO_1517 (O_1517,N_26297,N_27890);
nor UO_1518 (O_1518,N_28437,N_29081);
and UO_1519 (O_1519,N_26078,N_27794);
xnor UO_1520 (O_1520,N_28985,N_24281);
and UO_1521 (O_1521,N_24874,N_29890);
nand UO_1522 (O_1522,N_28428,N_25256);
or UO_1523 (O_1523,N_26548,N_28859);
nor UO_1524 (O_1524,N_26847,N_26022);
xnor UO_1525 (O_1525,N_28050,N_24186);
or UO_1526 (O_1526,N_28114,N_25894);
nor UO_1527 (O_1527,N_25138,N_26766);
nor UO_1528 (O_1528,N_26351,N_26744);
and UO_1529 (O_1529,N_25206,N_29282);
nor UO_1530 (O_1530,N_29597,N_26763);
nand UO_1531 (O_1531,N_26273,N_29440);
nand UO_1532 (O_1532,N_29513,N_24924);
nor UO_1533 (O_1533,N_29044,N_27282);
or UO_1534 (O_1534,N_28011,N_26892);
and UO_1535 (O_1535,N_29024,N_29724);
and UO_1536 (O_1536,N_28194,N_29873);
or UO_1537 (O_1537,N_26798,N_29141);
and UO_1538 (O_1538,N_24906,N_26629);
nand UO_1539 (O_1539,N_26593,N_25192);
and UO_1540 (O_1540,N_28832,N_27120);
or UO_1541 (O_1541,N_26557,N_26097);
xor UO_1542 (O_1542,N_24087,N_29381);
xnor UO_1543 (O_1543,N_26118,N_25810);
and UO_1544 (O_1544,N_24686,N_26296);
and UO_1545 (O_1545,N_29622,N_24226);
nand UO_1546 (O_1546,N_24612,N_27904);
and UO_1547 (O_1547,N_28913,N_29479);
and UO_1548 (O_1548,N_24757,N_27887);
xnor UO_1549 (O_1549,N_24774,N_26254);
nor UO_1550 (O_1550,N_29993,N_29510);
or UO_1551 (O_1551,N_25174,N_29455);
xor UO_1552 (O_1552,N_28816,N_28029);
nand UO_1553 (O_1553,N_28942,N_26755);
nand UO_1554 (O_1554,N_27198,N_27123);
nand UO_1555 (O_1555,N_29955,N_29072);
xnor UO_1556 (O_1556,N_25638,N_27517);
or UO_1557 (O_1557,N_25690,N_25519);
nor UO_1558 (O_1558,N_26201,N_29065);
nor UO_1559 (O_1559,N_25156,N_24227);
nor UO_1560 (O_1560,N_29264,N_29858);
or UO_1561 (O_1561,N_29606,N_29169);
xor UO_1562 (O_1562,N_24463,N_28538);
nand UO_1563 (O_1563,N_28464,N_28201);
or UO_1564 (O_1564,N_27342,N_24275);
xnor UO_1565 (O_1565,N_27097,N_25275);
or UO_1566 (O_1566,N_27629,N_24061);
or UO_1567 (O_1567,N_25216,N_25115);
xor UO_1568 (O_1568,N_24451,N_27862);
xnor UO_1569 (O_1569,N_25020,N_26669);
and UO_1570 (O_1570,N_29383,N_27411);
or UO_1571 (O_1571,N_29050,N_28968);
nand UO_1572 (O_1572,N_29392,N_28435);
xnor UO_1573 (O_1573,N_29877,N_29881);
nand UO_1574 (O_1574,N_26632,N_24326);
or UO_1575 (O_1575,N_28357,N_27286);
nor UO_1576 (O_1576,N_27698,N_26986);
or UO_1577 (O_1577,N_27102,N_26027);
and UO_1578 (O_1578,N_26465,N_29849);
or UO_1579 (O_1579,N_25351,N_25778);
nand UO_1580 (O_1580,N_27228,N_26126);
nor UO_1581 (O_1581,N_24108,N_25528);
xor UO_1582 (O_1582,N_29407,N_29717);
nand UO_1583 (O_1583,N_29187,N_24650);
nand UO_1584 (O_1584,N_25342,N_28354);
and UO_1585 (O_1585,N_27625,N_28986);
nand UO_1586 (O_1586,N_26598,N_28408);
and UO_1587 (O_1587,N_25735,N_24471);
and UO_1588 (O_1588,N_25744,N_25769);
nor UO_1589 (O_1589,N_27571,N_26347);
nand UO_1590 (O_1590,N_24764,N_24549);
or UO_1591 (O_1591,N_28044,N_26039);
nor UO_1592 (O_1592,N_24690,N_28017);
nand UO_1593 (O_1593,N_24537,N_28708);
and UO_1594 (O_1594,N_27934,N_28669);
and UO_1595 (O_1595,N_27339,N_24149);
or UO_1596 (O_1596,N_28663,N_27974);
nand UO_1597 (O_1597,N_25921,N_28146);
and UO_1598 (O_1598,N_27275,N_27344);
nand UO_1599 (O_1599,N_24864,N_25495);
nand UO_1600 (O_1600,N_28752,N_29569);
or UO_1601 (O_1601,N_26710,N_29229);
xnor UO_1602 (O_1602,N_27953,N_29998);
and UO_1603 (O_1603,N_25760,N_24003);
nand UO_1604 (O_1604,N_28959,N_27908);
nand UO_1605 (O_1605,N_29883,N_29948);
or UO_1606 (O_1606,N_25667,N_27090);
nor UO_1607 (O_1607,N_25762,N_28291);
or UO_1608 (O_1608,N_24072,N_27038);
or UO_1609 (O_1609,N_29129,N_29431);
nor UO_1610 (O_1610,N_24415,N_25041);
xnor UO_1611 (O_1611,N_27831,N_25159);
nand UO_1612 (O_1612,N_27626,N_29261);
and UO_1613 (O_1613,N_28794,N_28533);
and UO_1614 (O_1614,N_25385,N_29232);
and UO_1615 (O_1615,N_27645,N_27941);
xnor UO_1616 (O_1616,N_29104,N_27528);
nor UO_1617 (O_1617,N_29070,N_24036);
xnor UO_1618 (O_1618,N_24204,N_25130);
and UO_1619 (O_1619,N_24685,N_26329);
nor UO_1620 (O_1620,N_24320,N_24428);
and UO_1621 (O_1621,N_29397,N_26011);
nand UO_1622 (O_1622,N_29317,N_29058);
nor UO_1623 (O_1623,N_28332,N_25709);
xor UO_1624 (O_1624,N_27422,N_29482);
and UO_1625 (O_1625,N_25961,N_25651);
nor UO_1626 (O_1626,N_27452,N_27783);
xnor UO_1627 (O_1627,N_24531,N_24513);
and UO_1628 (O_1628,N_28586,N_28774);
nand UO_1629 (O_1629,N_28013,N_25422);
nand UO_1630 (O_1630,N_24146,N_28323);
xor UO_1631 (O_1631,N_28090,N_27172);
nor UO_1632 (O_1632,N_24291,N_26709);
nor UO_1633 (O_1633,N_29161,N_28460);
nor UO_1634 (O_1634,N_25037,N_25963);
xnor UO_1635 (O_1635,N_28267,N_28112);
nand UO_1636 (O_1636,N_28069,N_28977);
nand UO_1637 (O_1637,N_27770,N_26511);
nand UO_1638 (O_1638,N_24598,N_26532);
xnor UO_1639 (O_1639,N_26853,N_28486);
nor UO_1640 (O_1640,N_24296,N_26345);
and UO_1641 (O_1641,N_25550,N_27782);
and UO_1642 (O_1642,N_29679,N_27204);
nor UO_1643 (O_1643,N_25067,N_29645);
nor UO_1644 (O_1644,N_29802,N_27745);
nand UO_1645 (O_1645,N_25098,N_28858);
nand UO_1646 (O_1646,N_28775,N_27912);
or UO_1647 (O_1647,N_26190,N_25555);
xnor UO_1648 (O_1648,N_28002,N_27481);
and UO_1649 (O_1649,N_29398,N_25668);
or UO_1650 (O_1650,N_29594,N_25450);
nand UO_1651 (O_1651,N_27753,N_26754);
and UO_1652 (O_1652,N_24130,N_26002);
or UO_1653 (O_1653,N_25011,N_26874);
nand UO_1654 (O_1654,N_28075,N_24805);
xnor UO_1655 (O_1655,N_29085,N_29084);
or UO_1656 (O_1656,N_25423,N_27202);
nand UO_1657 (O_1657,N_29204,N_26746);
and UO_1658 (O_1658,N_25369,N_28568);
or UO_1659 (O_1659,N_24215,N_29878);
or UO_1660 (O_1660,N_25441,N_28649);
or UO_1661 (O_1661,N_25829,N_24562);
or UO_1662 (O_1662,N_25375,N_26062);
xor UO_1663 (O_1663,N_26215,N_25368);
xor UO_1664 (O_1664,N_26145,N_27154);
nand UO_1665 (O_1665,N_24902,N_25823);
nand UO_1666 (O_1666,N_27521,N_27007);
xor UO_1667 (O_1667,N_25181,N_26788);
and UO_1668 (O_1668,N_25424,N_28597);
nand UO_1669 (O_1669,N_28915,N_28439);
nor UO_1670 (O_1670,N_28390,N_25081);
xor UO_1671 (O_1671,N_24437,N_29994);
nand UO_1672 (O_1672,N_27155,N_29342);
nand UO_1673 (O_1673,N_27324,N_26242);
nor UO_1674 (O_1674,N_29195,N_25398);
nor UO_1675 (O_1675,N_27730,N_25682);
and UO_1676 (O_1676,N_25644,N_24188);
nor UO_1677 (O_1677,N_27787,N_27161);
nand UO_1678 (O_1678,N_25068,N_28445);
and UO_1679 (O_1679,N_26180,N_25413);
nor UO_1680 (O_1680,N_27468,N_26496);
xnor UO_1681 (O_1681,N_25736,N_24025);
or UO_1682 (O_1682,N_29704,N_28814);
nand UO_1683 (O_1683,N_27329,N_27656);
nand UO_1684 (O_1684,N_27147,N_29213);
nor UO_1685 (O_1685,N_28083,N_24715);
nand UO_1686 (O_1686,N_29721,N_25080);
nor UO_1687 (O_1687,N_27774,N_28715);
or UO_1688 (O_1688,N_24039,N_29032);
nand UO_1689 (O_1689,N_27503,N_28638);
or UO_1690 (O_1690,N_29816,N_26539);
and UO_1691 (O_1691,N_26302,N_29359);
xor UO_1692 (O_1692,N_28779,N_24987);
or UO_1693 (O_1693,N_26422,N_24065);
nor UO_1694 (O_1694,N_27397,N_25328);
xnor UO_1695 (O_1695,N_28878,N_27666);
xnor UO_1696 (O_1696,N_24722,N_28935);
nand UO_1697 (O_1697,N_27295,N_27633);
xor UO_1698 (O_1698,N_28309,N_27331);
nand UO_1699 (O_1699,N_24173,N_29596);
nand UO_1700 (O_1700,N_25577,N_27373);
and UO_1701 (O_1701,N_27096,N_29275);
or UO_1702 (O_1702,N_27239,N_24088);
nand UO_1703 (O_1703,N_24930,N_25523);
or UO_1704 (O_1704,N_28899,N_27915);
and UO_1705 (O_1705,N_28241,N_28209);
xnor UO_1706 (O_1706,N_28951,N_24878);
nand UO_1707 (O_1707,N_26281,N_24182);
xnor UO_1708 (O_1708,N_25071,N_25346);
nor UO_1709 (O_1709,N_27450,N_29471);
and UO_1710 (O_1710,N_24879,N_25335);
xor UO_1711 (O_1711,N_29787,N_26673);
nand UO_1712 (O_1712,N_26432,N_27715);
and UO_1713 (O_1713,N_26127,N_28389);
nand UO_1714 (O_1714,N_25898,N_28984);
nand UO_1715 (O_1715,N_28737,N_29739);
nor UO_1716 (O_1716,N_24522,N_27216);
and UO_1717 (O_1717,N_25580,N_28581);
nor UO_1718 (O_1718,N_28126,N_28869);
nor UO_1719 (O_1719,N_29477,N_29914);
xnor UO_1720 (O_1720,N_24809,N_27053);
or UO_1721 (O_1721,N_27728,N_26865);
or UO_1722 (O_1722,N_27362,N_29544);
or UO_1723 (O_1723,N_26870,N_27400);
nand UO_1724 (O_1724,N_25023,N_29574);
xnor UO_1725 (O_1725,N_29693,N_29355);
nand UO_1726 (O_1726,N_27798,N_29536);
xor UO_1727 (O_1727,N_27092,N_25343);
nor UO_1728 (O_1728,N_26443,N_28644);
or UO_1729 (O_1729,N_24222,N_24092);
xor UO_1730 (O_1730,N_29581,N_28300);
xnor UO_1731 (O_1731,N_28225,N_24816);
and UO_1732 (O_1732,N_27523,N_24402);
xor UO_1733 (O_1733,N_28060,N_28406);
and UO_1734 (O_1734,N_25497,N_28981);
nand UO_1735 (O_1735,N_26361,N_28318);
nand UO_1736 (O_1736,N_25761,N_28289);
nor UO_1737 (O_1737,N_27027,N_25489);
xor UO_1738 (O_1738,N_26758,N_24701);
nand UO_1739 (O_1739,N_28471,N_27043);
nor UO_1740 (O_1740,N_26543,N_29047);
or UO_1741 (O_1741,N_25920,N_24970);
nand UO_1742 (O_1742,N_25845,N_27445);
and UO_1743 (O_1743,N_27465,N_29614);
nand UO_1744 (O_1744,N_27788,N_26309);
nand UO_1745 (O_1745,N_24900,N_25984);
nor UO_1746 (O_1746,N_27050,N_24586);
or UO_1747 (O_1747,N_26046,N_24980);
and UO_1748 (O_1748,N_24623,N_25047);
xnor UO_1749 (O_1749,N_26053,N_26959);
nand UO_1750 (O_1750,N_26025,N_27019);
nand UO_1751 (O_1751,N_29785,N_28637);
nand UO_1752 (O_1752,N_28234,N_26036);
xnor UO_1753 (O_1753,N_28528,N_27643);
nor UO_1754 (O_1754,N_25326,N_27474);
xnor UO_1755 (O_1755,N_29115,N_24739);
or UO_1756 (O_1756,N_26112,N_28746);
xnor UO_1757 (O_1757,N_27764,N_25869);
nand UO_1758 (O_1758,N_26739,N_28903);
and UO_1759 (O_1759,N_28803,N_26290);
and UO_1760 (O_1760,N_25312,N_26864);
and UO_1761 (O_1761,N_26272,N_28499);
and UO_1762 (O_1762,N_26208,N_29028);
or UO_1763 (O_1763,N_27390,N_25389);
nor UO_1764 (O_1764,N_29485,N_28168);
nor UO_1765 (O_1765,N_27423,N_24062);
and UO_1766 (O_1766,N_29331,N_29737);
nor UO_1767 (O_1767,N_26822,N_25486);
nand UO_1768 (O_1768,N_27632,N_28023);
nand UO_1769 (O_1769,N_27442,N_24983);
nand UO_1770 (O_1770,N_27146,N_26610);
or UO_1771 (O_1771,N_24979,N_25280);
nor UO_1772 (O_1772,N_28626,N_25942);
nor UO_1773 (O_1773,N_27756,N_29029);
nand UO_1774 (O_1774,N_27075,N_27877);
and UO_1775 (O_1775,N_24292,N_25093);
nand UO_1776 (O_1776,N_27409,N_29316);
or UO_1777 (O_1777,N_25022,N_26587);
nor UO_1778 (O_1778,N_25244,N_25768);
nand UO_1779 (O_1779,N_27306,N_26564);
xor UO_1780 (O_1780,N_27852,N_28034);
and UO_1781 (O_1781,N_25243,N_24877);
and UO_1782 (O_1782,N_28524,N_25631);
or UO_1783 (O_1783,N_28792,N_25696);
or UO_1784 (O_1784,N_25418,N_26942);
nor UO_1785 (O_1785,N_25128,N_26474);
or UO_1786 (O_1786,N_28946,N_24131);
nand UO_1787 (O_1787,N_25853,N_26198);
nor UO_1788 (O_1788,N_29917,N_26565);
and UO_1789 (O_1789,N_26762,N_26569);
xnor UO_1790 (O_1790,N_27447,N_27671);
nand UO_1791 (O_1791,N_26502,N_24142);
and UO_1792 (O_1792,N_24259,N_24067);
and UO_1793 (O_1793,N_24994,N_27603);
nand UO_1794 (O_1794,N_28103,N_25264);
and UO_1795 (O_1795,N_26810,N_29862);
nand UO_1796 (O_1796,N_25463,N_28846);
nor UO_1797 (O_1797,N_29323,N_28620);
and UO_1798 (O_1798,N_27701,N_26483);
or UO_1799 (O_1799,N_29462,N_24388);
nand UO_1800 (O_1800,N_24720,N_27271);
xor UO_1801 (O_1801,N_29303,N_28600);
or UO_1802 (O_1802,N_25992,N_25997);
xor UO_1803 (O_1803,N_24927,N_24575);
and UO_1804 (O_1804,N_27652,N_26203);
nand UO_1805 (O_1805,N_24368,N_24477);
xor UO_1806 (O_1806,N_24123,N_29430);
or UO_1807 (O_1807,N_27099,N_29809);
and UO_1808 (O_1808,N_25636,N_27525);
xnor UO_1809 (O_1809,N_25657,N_28218);
nand UO_1810 (O_1810,N_25794,N_26818);
nand UO_1811 (O_1811,N_26291,N_27122);
nand UO_1812 (O_1812,N_24978,N_29567);
nand UO_1813 (O_1813,N_28233,N_27134);
and UO_1814 (O_1814,N_25465,N_27336);
nor UO_1815 (O_1815,N_24543,N_28142);
and UO_1816 (O_1816,N_26856,N_24161);
xnor UO_1817 (O_1817,N_28799,N_24621);
nand UO_1818 (O_1818,N_27151,N_29579);
or UO_1819 (O_1819,N_27089,N_29727);
or UO_1820 (O_1820,N_29612,N_26453);
nand UO_1821 (O_1821,N_28159,N_28027);
xor UO_1822 (O_1822,N_28585,N_26656);
nor UO_1823 (O_1823,N_29269,N_25836);
nand UO_1824 (O_1824,N_28138,N_27829);
or UO_1825 (O_1825,N_27743,N_28570);
nand UO_1826 (O_1826,N_24625,N_29182);
nor UO_1827 (O_1827,N_24755,N_27428);
or UO_1828 (O_1828,N_26840,N_27023);
nor UO_1829 (O_1829,N_28025,N_24462);
and UO_1830 (O_1830,N_29780,N_26713);
nand UO_1831 (O_1831,N_24769,N_28749);
xor UO_1832 (O_1832,N_27870,N_27657);
or UO_1833 (O_1833,N_29074,N_24887);
and UO_1834 (O_1834,N_27543,N_24446);
nor UO_1835 (O_1835,N_24467,N_26734);
or UO_1836 (O_1836,N_29683,N_27833);
nor UO_1837 (O_1837,N_29506,N_25922);
nand UO_1838 (O_1838,N_26908,N_26833);
and UO_1839 (O_1839,N_28258,N_26048);
nand UO_1840 (O_1840,N_28508,N_27735);
nand UO_1841 (O_1841,N_25635,N_29810);
and UO_1842 (O_1842,N_26204,N_25660);
nor UO_1843 (O_1843,N_29108,N_24246);
xor UO_1844 (O_1844,N_28087,N_26740);
xnor UO_1845 (O_1845,N_24098,N_26553);
xor UO_1846 (O_1846,N_28306,N_26932);
nor UO_1847 (O_1847,N_26528,N_27348);
and UO_1848 (O_1848,N_27314,N_29100);
nor UO_1849 (O_1849,N_26513,N_26889);
nor UO_1850 (O_1850,N_24252,N_25430);
or UO_1851 (O_1851,N_29970,N_25902);
xor UO_1852 (O_1852,N_26087,N_26808);
xnor UO_1853 (O_1853,N_28888,N_24811);
nand UO_1854 (O_1854,N_29427,N_29518);
nand UO_1855 (O_1855,N_26420,N_29247);
and UO_1856 (O_1856,N_28549,N_26270);
xor UO_1857 (O_1857,N_28264,N_29400);
xnor UO_1858 (O_1858,N_29782,N_24315);
nand UO_1859 (O_1859,N_29746,N_25576);
and UO_1860 (O_1860,N_26606,N_28844);
xor UO_1861 (O_1861,N_24021,N_28232);
and UO_1862 (O_1862,N_27996,N_26907);
xnor UO_1863 (O_1863,N_29483,N_25161);
or UO_1864 (O_1864,N_25787,N_26603);
and UO_1865 (O_1865,N_28255,N_27630);
nor UO_1866 (O_1866,N_29558,N_25617);
xor UO_1867 (O_1867,N_25927,N_27140);
xnor UO_1868 (O_1868,N_25340,N_26374);
xor UO_1869 (O_1869,N_29866,N_27143);
and UO_1870 (O_1870,N_27003,N_27762);
nand UO_1871 (O_1871,N_27678,N_25207);
and UO_1872 (O_1872,N_27519,N_28120);
nand UO_1873 (O_1873,N_28262,N_29283);
and UO_1874 (O_1874,N_27345,N_25102);
xnor UO_1875 (O_1875,N_26381,N_29414);
xor UO_1876 (O_1876,N_28285,N_28884);
nand UO_1877 (O_1877,N_25940,N_25240);
nand UO_1878 (O_1878,N_25538,N_28835);
or UO_1879 (O_1879,N_29001,N_27872);
nand UO_1880 (O_1880,N_25819,N_29376);
xnor UO_1881 (O_1881,N_27844,N_29956);
and UO_1882 (O_1882,N_26070,N_28819);
xnor UO_1883 (O_1883,N_26885,N_25478);
nand UO_1884 (O_1884,N_24284,N_28504);
and UO_1885 (O_1885,N_28356,N_26160);
xnor UO_1886 (O_1886,N_27242,N_27406);
or UO_1887 (O_1887,N_27839,N_24731);
and UO_1888 (O_1888,N_26098,N_25411);
xor UO_1889 (O_1889,N_29769,N_25142);
xnor UO_1890 (O_1890,N_28308,N_27716);
nand UO_1891 (O_1891,N_27835,N_28932);
nand UO_1892 (O_1892,N_24555,N_25701);
or UO_1893 (O_1893,N_29478,N_26791);
nor UO_1894 (O_1894,N_24244,N_24509);
nand UO_1895 (O_1895,N_27618,N_28509);
and UO_1896 (O_1896,N_24498,N_29899);
nor UO_1897 (O_1897,N_25435,N_24011);
nand UO_1898 (O_1898,N_26895,N_29532);
xor UO_1899 (O_1899,N_28330,N_27416);
nor UO_1900 (O_1900,N_27293,N_24193);
nand UO_1901 (O_1901,N_27440,N_29582);
and UO_1902 (O_1902,N_27060,N_28849);
nor UO_1903 (O_1903,N_25145,N_25163);
and UO_1904 (O_1904,N_27840,N_24216);
and UO_1905 (O_1905,N_29646,N_24671);
and UO_1906 (O_1906,N_24209,N_28680);
and UO_1907 (O_1907,N_25116,N_29008);
nor UO_1908 (O_1908,N_27744,N_28484);
or UO_1909 (O_1909,N_24473,N_24751);
xor UO_1910 (O_1910,N_29825,N_29208);
or UO_1911 (O_1911,N_27638,N_28656);
nand UO_1912 (O_1912,N_24421,N_28956);
nand UO_1913 (O_1913,N_27322,N_29469);
and UO_1914 (O_1914,N_26604,N_26390);
nor UO_1915 (O_1915,N_26498,N_27899);
and UO_1916 (O_1916,N_26157,N_24042);
or UO_1917 (O_1917,N_26514,N_29033);
and UO_1918 (O_1918,N_29406,N_24899);
xnor UO_1919 (O_1919,N_29638,N_24422);
and UO_1920 (O_1920,N_25188,N_28157);
or UO_1921 (O_1921,N_26714,N_29571);
nand UO_1922 (O_1922,N_26931,N_27903);
and UO_1923 (O_1923,N_28567,N_27358);
xor UO_1924 (O_1924,N_25950,N_24485);
and UO_1925 (O_1925,N_27290,N_25221);
nand UO_1926 (O_1926,N_25789,N_25479);
and UO_1927 (O_1927,N_24605,N_28109);
nor UO_1928 (O_1928,N_24665,N_26362);
nor UO_1929 (O_1929,N_24982,N_27316);
or UO_1930 (O_1930,N_29656,N_25457);
xnor UO_1931 (O_1931,N_29030,N_24356);
nor UO_1932 (O_1932,N_24365,N_26775);
or UO_1933 (O_1933,N_28364,N_24310);
or UO_1934 (O_1934,N_27136,N_27553);
nand UO_1935 (O_1935,N_29999,N_28791);
nor UO_1936 (O_1936,N_28009,N_27754);
nor UO_1937 (O_1937,N_28647,N_29016);
nor UO_1938 (O_1938,N_27458,N_26877);
or UO_1939 (O_1939,N_26320,N_29580);
xnor UO_1940 (O_1940,N_27156,N_25724);
or UO_1941 (O_1941,N_26230,N_28547);
xor UO_1942 (O_1942,N_25609,N_28515);
and UO_1943 (O_1943,N_25208,N_28873);
and UO_1944 (O_1944,N_24232,N_29635);
and UO_1945 (O_1945,N_27364,N_28041);
and UO_1946 (O_1946,N_24097,N_27299);
and UO_1947 (O_1947,N_25149,N_28745);
and UO_1948 (O_1948,N_26921,N_24229);
nor UO_1949 (O_1949,N_24258,N_29938);
nand UO_1950 (O_1950,N_26767,N_28348);
xor UO_1951 (O_1951,N_28269,N_27196);
or UO_1952 (O_1952,N_29761,N_28030);
or UO_1953 (O_1953,N_29061,N_26330);
or UO_1954 (O_1954,N_29015,N_26665);
and UO_1955 (O_1955,N_25712,N_25227);
or UO_1956 (O_1956,N_29841,N_24381);
and UO_1957 (O_1957,N_24950,N_26730);
nand UO_1958 (O_1958,N_24104,N_25120);
and UO_1959 (O_1959,N_26399,N_29563);
and UO_1960 (O_1960,N_25798,N_24126);
nor UO_1961 (O_1961,N_25069,N_27815);
nand UO_1962 (O_1962,N_26935,N_27205);
nand UO_1963 (O_1963,N_28712,N_26660);
or UO_1964 (O_1964,N_26698,N_28482);
nor UO_1965 (O_1965,N_25150,N_29959);
nor UO_1966 (O_1966,N_28429,N_26696);
nor UO_1967 (O_1967,N_26652,N_29538);
or UO_1968 (O_1968,N_29366,N_25627);
xor UO_1969 (O_1969,N_26184,N_26268);
or UO_1970 (O_1970,N_29649,N_27417);
nand UO_1971 (O_1971,N_26250,N_26350);
and UO_1972 (O_1972,N_26013,N_24479);
nand UO_1973 (O_1973,N_27842,N_28489);
or UO_1974 (O_1974,N_24830,N_24546);
xnor UO_1975 (O_1975,N_26782,N_29781);
nand UO_1976 (O_1976,N_26973,N_27900);
nand UO_1977 (O_1977,N_29752,N_28248);
nor UO_1978 (O_1978,N_26442,N_26440);
nand UO_1979 (O_1979,N_27208,N_27124);
or UO_1980 (O_1980,N_28840,N_29516);
nand UO_1981 (O_1981,N_24237,N_27193);
xor UO_1982 (O_1982,N_27886,N_24416);
and UO_1983 (O_1983,N_27918,N_26984);
and UO_1984 (O_1984,N_27647,N_24374);
and UO_1985 (O_1985,N_24639,N_25048);
and UO_1986 (O_1986,N_26059,N_24355);
xor UO_1987 (O_1987,N_27082,N_27135);
nand UO_1988 (O_1988,N_24895,N_24155);
nand UO_1989 (O_1989,N_24584,N_29438);
xnor UO_1990 (O_1990,N_29642,N_25381);
nor UO_1991 (O_1991,N_25742,N_26745);
nor UO_1992 (O_1992,N_27598,N_29664);
or UO_1993 (O_1993,N_29947,N_25027);
or UO_1994 (O_1994,N_27471,N_29214);
and UO_1995 (O_1995,N_28062,N_25191);
or UO_1996 (O_1996,N_25781,N_24297);
or UO_1997 (O_1997,N_26470,N_24918);
xnor UO_1998 (O_1998,N_28853,N_28178);
or UO_1999 (O_1999,N_25630,N_27554);
or UO_2000 (O_2000,N_24661,N_29230);
and UO_2001 (O_2001,N_27018,N_26982);
nor UO_2002 (O_2002,N_24989,N_25642);
nand UO_2003 (O_2003,N_26169,N_28662);
nand UO_2004 (O_2004,N_26231,N_28487);
nor UO_2005 (O_2005,N_25553,N_28051);
and UO_2006 (O_2006,N_27153,N_29952);
and UO_2007 (O_2007,N_27649,N_28171);
xnor UO_2008 (O_2008,N_27884,N_25079);
nor UO_2009 (O_2009,N_27648,N_27561);
or UO_2010 (O_2010,N_25234,N_26076);
nor UO_2011 (O_2011,N_24618,N_28394);
nand UO_2012 (O_2012,N_24321,N_25222);
and UO_2013 (O_2013,N_27377,N_26251);
nor UO_2014 (O_2014,N_24797,N_28874);
and UO_2015 (O_2015,N_25421,N_26857);
nand UO_2016 (O_2016,N_26772,N_24597);
nand UO_2017 (O_2017,N_27950,N_26556);
xor UO_2018 (O_2018,N_25688,N_28278);
or UO_2019 (O_2019,N_27763,N_28375);
nand UO_2020 (O_2020,N_25699,N_25257);
xor UO_2021 (O_2021,N_28550,N_27578);
xnor UO_2022 (O_2022,N_29098,N_25235);
nor UO_2023 (O_2023,N_25600,N_28704);
nor UO_2024 (O_2024,N_25345,N_25332);
nor UO_2025 (O_2025,N_27965,N_29978);
and UO_2026 (O_2026,N_27562,N_25833);
nand UO_2027 (O_2027,N_29940,N_27694);
or UO_2028 (O_2028,N_27396,N_25958);
nand UO_2029 (O_2029,N_29906,N_26236);
nand UO_2030 (O_2030,N_29605,N_26695);
xor UO_2031 (O_2031,N_29109,N_24508);
and UO_2032 (O_2032,N_29432,N_29672);
nand UO_2033 (O_2033,N_26923,N_29211);
nor UO_2034 (O_2034,N_27231,N_25311);
nor UO_2035 (O_2035,N_29329,N_24783);
xnor UO_2036 (O_2036,N_24620,N_28260);
nor UO_2037 (O_2037,N_27042,N_25242);
nor UO_2038 (O_2038,N_27449,N_29668);
nor UO_2039 (O_2039,N_24768,N_26435);
xor UO_2040 (O_2040,N_28352,N_27355);
or UO_2041 (O_2041,N_28372,N_27401);
xor UO_2042 (O_2042,N_24059,N_28304);
nor UO_2043 (O_2043,N_29489,N_27484);
nor UO_2044 (O_2044,N_24893,N_26331);
or UO_2045 (O_2045,N_25811,N_24867);
or UO_2046 (O_2046,N_28603,N_27125);
nor UO_2047 (O_2047,N_29694,N_24888);
and UO_2048 (O_2048,N_25273,N_26961);
or UO_2049 (O_2049,N_29587,N_27340);
and UO_2050 (O_2050,N_26317,N_25303);
xor UO_2051 (O_2051,N_26913,N_25101);
or UO_2052 (O_2052,N_29333,N_29006);
nor UO_2053 (O_2053,N_25183,N_25453);
nand UO_2054 (O_2054,N_28976,N_29946);
xnor UO_2055 (O_2055,N_26691,N_29660);
nor UO_2056 (O_2056,N_26375,N_29310);
and UO_2057 (O_2057,N_29309,N_27405);
nand UO_2058 (O_2058,N_28054,N_25339);
nor UO_2059 (O_2059,N_26378,N_24934);
and UO_2060 (O_2060,N_29590,N_25306);
nand UO_2061 (O_2061,N_27049,N_25378);
or UO_2062 (O_2062,N_24143,N_27056);
nor UO_2063 (O_2063,N_29130,N_25412);
nand UO_2064 (O_2064,N_29036,N_28074);
and UO_2065 (O_2065,N_27990,N_24206);
xnor UO_2066 (O_2066,N_26207,N_28592);
and UO_2067 (O_2067,N_29221,N_29941);
and UO_2068 (O_2068,N_29012,N_27188);
nor UO_2069 (O_2069,N_27597,N_26991);
and UO_2070 (O_2070,N_27429,N_27495);
and UO_2071 (O_2071,N_29811,N_28618);
nor UO_2072 (O_2072,N_27361,N_29139);
nand UO_2073 (O_2073,N_26427,N_29179);
xnor UO_2074 (O_2074,N_25379,N_28053);
nand UO_2075 (O_2075,N_26348,N_24475);
or UO_2076 (O_2076,N_27956,N_28162);
xor UO_2077 (O_2077,N_25752,N_28387);
xor UO_2078 (O_2078,N_29346,N_24358);
nor UO_2079 (O_2079,N_26504,N_24633);
and UO_2080 (O_2080,N_25480,N_28477);
and UO_2081 (O_2081,N_24510,N_29919);
nor UO_2082 (O_2082,N_27873,N_24540);
nand UO_2083 (O_2083,N_26799,N_25232);
nand UO_2084 (O_2084,N_26086,N_28231);
xor UO_2085 (O_2085,N_24183,N_25359);
nor UO_2086 (O_2086,N_29520,N_25447);
nand UO_2087 (O_2087,N_28191,N_28554);
xor UO_2088 (O_2088,N_27667,N_24695);
nand UO_2089 (O_2089,N_24808,N_25904);
xor UO_2090 (O_2090,N_29089,N_28061);
nor UO_2091 (O_2091,N_25471,N_26579);
nand UO_2092 (O_2092,N_24590,N_28071);
or UO_2093 (O_2093,N_24868,N_28939);
nand UO_2094 (O_2094,N_25948,N_26770);
or UO_2095 (O_2095,N_25402,N_26151);
xor UO_2096 (O_2096,N_29470,N_27076);
nand UO_2097 (O_2097,N_27998,N_29566);
or UO_2098 (O_2098,N_24314,N_29819);
and UO_2099 (O_2099,N_24885,N_29847);
and UO_2100 (O_2100,N_24869,N_26697);
xnor UO_2101 (O_2101,N_25353,N_27803);
or UO_2102 (O_2102,N_28110,N_26325);
nand UO_2103 (O_2103,N_29252,N_24208);
and UO_2104 (O_2104,N_26129,N_28446);
nand UO_2105 (O_2105,N_25151,N_27679);
xnor UO_2106 (O_2106,N_28800,N_29613);
xnor UO_2107 (O_2107,N_25099,N_27717);
and UO_2108 (O_2108,N_29492,N_29467);
or UO_2109 (O_2109,N_28941,N_27881);
and UO_2110 (O_2110,N_25572,N_26786);
xnor UO_2111 (O_2111,N_26647,N_26567);
nor UO_2112 (O_2112,N_27353,N_25672);
nor UO_2113 (O_2113,N_28321,N_28493);
or UO_2114 (O_2114,N_25728,N_26342);
and UO_2115 (O_2115,N_26899,N_25205);
nand UO_2116 (O_2116,N_25437,N_28699);
nor UO_2117 (O_2117,N_28067,N_24170);
or UO_2118 (O_2118,N_25656,N_29666);
nand UO_2119 (O_2119,N_27025,N_27363);
xnor UO_2120 (O_2120,N_26574,N_26353);
xor UO_2121 (O_2121,N_24544,N_28417);
nand UO_2122 (O_2122,N_27999,N_28470);
nand UO_2123 (O_2123,N_29480,N_26966);
nor UO_2124 (O_2124,N_26000,N_25490);
nor UO_2125 (O_2125,N_28815,N_26252);
nand UO_2126 (O_2126,N_24395,N_27426);
or UO_2127 (O_2127,N_24399,N_29865);
xor UO_2128 (O_2128,N_25405,N_29692);
and UO_2129 (O_2129,N_28510,N_26455);
nand UO_2130 (O_2130,N_27388,N_25812);
nor UO_2131 (O_2131,N_28564,N_27577);
nor UO_2132 (O_2132,N_24664,N_29251);
nor UO_2133 (O_2133,N_24309,N_28197);
and UO_2134 (O_2134,N_25643,N_29066);
nand UO_2135 (O_2135,N_26500,N_29603);
xnor UO_2136 (O_2136,N_25856,N_25031);
xor UO_2137 (O_2137,N_28148,N_25796);
xnor UO_2138 (O_2138,N_29783,N_24046);
nand UO_2139 (O_2139,N_24681,N_26294);
nand UO_2140 (O_2140,N_24640,N_27280);
or UO_2141 (O_2141,N_29048,N_29004);
and UO_2142 (O_2142,N_27616,N_29192);
and UO_2143 (O_2143,N_26843,N_26354);
nor UO_2144 (O_2144,N_24850,N_28497);
nand UO_2145 (O_2145,N_25035,N_27799);
nand UO_2146 (O_2146,N_25166,N_26643);
nand UO_2147 (O_2147,N_24101,N_29634);
or UO_2148 (O_2148,N_28830,N_27065);
and UO_2149 (O_2149,N_29013,N_29435);
or UO_2150 (O_2150,N_26501,N_29760);
or UO_2151 (O_2151,N_26806,N_28311);
xnor UO_2152 (O_2152,N_25117,N_29260);
nor UO_2153 (O_2153,N_28115,N_28432);
and UO_2154 (O_2154,N_24319,N_24138);
or UO_2155 (O_2155,N_28731,N_26678);
nand UO_2156 (O_2156,N_28943,N_28703);
xnor UO_2157 (O_2157,N_29588,N_29075);
nor UO_2158 (O_2158,N_29549,N_29420);
nor UO_2159 (O_2159,N_27133,N_29526);
nand UO_2160 (O_2160,N_28770,N_26824);
nand UO_2161 (O_2161,N_27680,N_27438);
or UO_2162 (O_2162,N_24541,N_26323);
or UO_2163 (O_2163,N_24181,N_29741);
or UO_2164 (O_2164,N_25558,N_27876);
nor UO_2165 (O_2165,N_28147,N_24861);
nand UO_2166 (O_2166,N_28326,N_24457);
nor UO_2167 (O_2167,N_24693,N_25650);
or UO_2168 (O_2168,N_25251,N_27686);
and UO_2169 (O_2169,N_26555,N_24089);
and UO_2170 (O_2170,N_27178,N_25428);
or UO_2171 (O_2171,N_25064,N_27970);
nand UO_2172 (O_2172,N_29498,N_28190);
nor UO_2173 (O_2173,N_26582,N_27902);
and UO_2174 (O_2174,N_27776,N_25895);
xnor UO_2175 (O_2175,N_28206,N_27210);
xnor UO_2176 (O_2176,N_24007,N_27635);
nor UO_2177 (O_2177,N_29315,N_26134);
xnor UO_2178 (O_2178,N_27935,N_24913);
and UO_2179 (O_2179,N_24418,N_25160);
and UO_2180 (O_2180,N_27619,N_28927);
nand UO_2181 (O_2181,N_26170,N_27473);
or UO_2182 (O_2182,N_25673,N_28690);
nand UO_2183 (O_2183,N_26038,N_29121);
nand UO_2184 (O_2184,N_24071,N_29630);
nand UO_2185 (O_2185,N_26779,N_26292);
nor UO_2186 (O_2186,N_27253,N_28908);
nand UO_2187 (O_2187,N_24932,N_25814);
xor UO_2188 (O_2188,N_27298,N_28003);
nand UO_2189 (O_2189,N_26096,N_28672);
xor UO_2190 (O_2190,N_27560,N_27113);
nand UO_2191 (O_2191,N_28548,N_25733);
and UO_2192 (O_2192,N_29253,N_26183);
nand UO_2193 (O_2193,N_26882,N_28739);
or UO_2194 (O_2194,N_26635,N_28447);
nand UO_2195 (O_2195,N_25292,N_25571);
and UO_2196 (O_2196,N_28760,N_24466);
nor UO_2197 (O_2197,N_24754,N_27121);
nand UO_2198 (O_2198,N_28579,N_26308);
xnor UO_2199 (O_2199,N_27557,N_26783);
nor UO_2200 (O_2200,N_28251,N_28268);
and UO_2201 (O_2201,N_24076,N_25305);
and UO_2202 (O_2202,N_28667,N_29517);
nand UO_2203 (O_2203,N_29984,N_28670);
xor UO_2204 (O_2204,N_28005,N_27972);
nor UO_2205 (O_2205,N_27371,N_29962);
and UO_2206 (O_2206,N_26664,N_24313);
or UO_2207 (O_2207,N_26289,N_28553);
nor UO_2208 (O_2208,N_24775,N_28141);
xnor UO_2209 (O_2209,N_29625,N_26974);
or UO_2210 (O_2210,N_24569,N_29953);
nand UO_2211 (O_2211,N_28047,N_28336);
and UO_2212 (O_2212,N_29487,N_29928);
xnor UO_2213 (O_2213,N_26507,N_27513);
nor UO_2214 (O_2214,N_28217,N_24812);
nand UO_2215 (O_2215,N_25785,N_26274);
xor UO_2216 (O_2216,N_24820,N_29527);
nand UO_2217 (O_2217,N_28671,N_27802);
nand UO_2218 (O_2218,N_27897,N_26197);
or UO_2219 (O_2219,N_26117,N_28238);
nor UO_2220 (O_2220,N_29995,N_29449);
or UO_2221 (O_2221,N_25909,N_29177);
xnor UO_2222 (O_2222,N_24556,N_28861);
nor UO_2223 (O_2223,N_27720,N_27748);
nand UO_2224 (O_2224,N_26327,N_26830);
or UO_2225 (O_2225,N_26520,N_27130);
nand UO_2226 (O_2226,N_25801,N_26682);
or UO_2227 (O_2227,N_26346,N_28000);
or UO_2228 (O_2228,N_27736,N_24999);
or UO_2229 (O_2229,N_29318,N_27084);
nor UO_2230 (O_2230,N_28851,N_29659);
nand UO_2231 (O_2231,N_28683,N_29188);
nor UO_2232 (O_2232,N_29193,N_28958);
and UO_2233 (O_2233,N_25831,N_29206);
xor UO_2234 (O_2234,N_28836,N_26314);
nor UO_2235 (O_2235,N_27922,N_25091);
nand UO_2236 (O_2236,N_24660,N_24603);
nor UO_2237 (O_2237,N_28883,N_28078);
nand UO_2238 (O_2238,N_24192,N_27317);
nand UO_2239 (O_2239,N_24445,N_28754);
and UO_2240 (O_2240,N_28569,N_28476);
nor UO_2241 (O_2241,N_27486,N_28558);
xnor UO_2242 (O_2242,N_29068,N_24384);
nor UO_2243 (O_2243,N_24583,N_28240);
or UO_2244 (O_2244,N_24922,N_27105);
xnor UO_2245 (O_2245,N_25175,N_24611);
xor UO_2246 (O_2246,N_26886,N_26679);
or UO_2247 (O_2247,N_26447,N_24796);
and UO_2248 (O_2248,N_29053,N_28829);
xor UO_2249 (O_2249,N_25014,N_25404);
nor UO_2250 (O_2250,N_24947,N_25055);
and UO_2251 (O_2251,N_28823,N_25599);
nand UO_2252 (O_2252,N_29241,N_24452);
xnor UO_2253 (O_2253,N_28713,N_27792);
or UO_2254 (O_2254,N_28293,N_26149);
and UO_2255 (O_2255,N_28176,N_24158);
xor UO_2256 (O_2256,N_29460,N_29618);
nand UO_2257 (O_2257,N_28442,N_25649);
xnor UO_2258 (O_2258,N_24948,N_27795);
nor UO_2259 (O_2259,N_24113,N_26753);
nand UO_2260 (O_2260,N_25843,N_25849);
xnor UO_2261 (O_2261,N_25567,N_29703);
and UO_2262 (O_2262,N_29154,N_28174);
and UO_2263 (O_2263,N_24506,N_27015);
or UO_2264 (O_2264,N_24400,N_27813);
nand UO_2265 (O_2265,N_26934,N_27800);
xor UO_2266 (O_2266,N_28837,N_29535);
and UO_2267 (O_2267,N_26277,N_28461);
nor UO_2268 (O_2268,N_25753,N_25979);
xor UO_2269 (O_2269,N_28419,N_24322);
or UO_2270 (O_2270,N_29465,N_26803);
or UO_2271 (O_2271,N_29573,N_24523);
nand UO_2272 (O_2272,N_24154,N_26368);
and UO_2273 (O_2273,N_25268,N_26881);
xnor UO_2274 (O_2274,N_28303,N_26284);
nand UO_2275 (O_2275,N_28400,N_26371);
nor UO_2276 (O_2276,N_28457,N_25314);
and UO_2277 (O_2277,N_27312,N_24111);
nor UO_2278 (O_2278,N_27995,N_26428);
xnor UO_2279 (O_2279,N_27781,N_24634);
nand UO_2280 (O_2280,N_25683,N_24382);
nor UO_2281 (O_2281,N_28028,N_25330);
nand UO_2282 (O_2282,N_28622,N_28136);
and UO_2283 (O_2283,N_24617,N_26475);
nor UO_2284 (O_2284,N_27552,N_26189);
nor UO_2285 (O_2285,N_25365,N_24289);
nor UO_2286 (O_2286,N_26572,N_28921);
nor UO_2287 (O_2287,N_29658,N_28879);
nand UO_2288 (O_2288,N_29602,N_26450);
nor UO_2289 (O_2289,N_29729,N_25361);
xor UO_2290 (O_2290,N_27167,N_29395);
or UO_2291 (O_2291,N_26106,N_26058);
xnor UO_2292 (O_2292,N_29972,N_26922);
nor UO_2293 (O_2293,N_24447,N_26482);
nor UO_2294 (O_2294,N_29907,N_27164);
or UO_2295 (O_2295,N_25556,N_26137);
nor UO_2296 (O_2296,N_25002,N_26055);
or UO_2297 (O_2297,N_24160,N_26033);
nand UO_2298 (O_2298,N_27673,N_29863);
nor UO_2299 (O_2299,N_28580,N_29227);
and UO_2300 (O_2300,N_25706,N_25223);
and UO_2301 (O_2301,N_29714,N_27175);
and UO_2302 (O_2302,N_28993,N_27819);
xnor UO_2303 (O_2303,N_25084,N_28735);
nor UO_2304 (O_2304,N_26558,N_29812);
xnor UO_2305 (O_2305,N_26471,N_26144);
and UO_2306 (O_2306,N_27751,N_27330);
nand UO_2307 (O_2307,N_27267,N_27419);
nand UO_2308 (O_2308,N_25299,N_25592);
or UO_2309 (O_2309,N_27509,N_28108);
and UO_2310 (O_2310,N_28280,N_24847);
nand UO_2311 (O_2311,N_26318,N_27257);
nor UO_2312 (O_2312,N_29126,N_25824);
nand UO_2313 (O_2313,N_29561,N_26789);
xor UO_2314 (O_2314,N_25809,N_28894);
xnor UO_2315 (O_2315,N_25883,N_27936);
and UO_2316 (O_2316,N_25162,N_26570);
nor UO_2317 (O_2317,N_25504,N_26718);
or UO_2318 (O_2318,N_29675,N_29875);
nand UO_2319 (O_2319,N_28574,N_24928);
nand UO_2320 (O_2320,N_29719,N_24977);
xor UO_2321 (O_2321,N_25949,N_24835);
nand UO_2322 (O_2322,N_28346,N_28104);
xor UO_2323 (O_2323,N_24304,N_24939);
or UO_2324 (O_2324,N_29842,N_25527);
nor UO_2325 (O_2325,N_27477,N_26927);
xnor UO_2326 (O_2326,N_26224,N_24124);
and UO_2327 (O_2327,N_26876,N_26549);
nor UO_2328 (O_2328,N_24106,N_24920);
and UO_2329 (O_2329,N_25675,N_28331);
nand UO_2330 (O_2330,N_27642,N_25274);
nor UO_2331 (O_2331,N_29891,N_27203);
nand UO_2332 (O_2332,N_24912,N_26751);
or UO_2333 (O_2333,N_27637,N_29992);
nor UO_2334 (O_2334,N_25186,N_24631);
or UO_2335 (O_2335,N_27497,N_26102);
nor UO_2336 (O_2336,N_24718,N_28526);
and UO_2337 (O_2337,N_27572,N_29262);
or UO_2338 (O_2338,N_26404,N_25626);
nand UO_2339 (O_2339,N_29005,N_29870);
nor UO_2340 (O_2340,N_24914,N_26863);
nand UO_2341 (O_2341,N_27609,N_24852);
or UO_2342 (O_2342,N_28353,N_29872);
and UO_2343 (O_2343,N_24018,N_29822);
nand UO_2344 (O_2344,N_27898,N_25165);
nor UO_2345 (O_2345,N_26749,N_26099);
and UO_2346 (O_2346,N_29689,N_25834);
and UO_2347 (O_2347,N_26550,N_27976);
nand UO_2348 (O_2348,N_28636,N_26743);
and UO_2349 (O_2349,N_26976,N_27439);
nor UO_2350 (O_2350,N_27424,N_27369);
or UO_2351 (O_2351,N_29401,N_28747);
nand UO_2352 (O_2352,N_26778,N_26173);
nor UO_2353 (O_2353,N_25560,N_28578);
or UO_2354 (O_2354,N_24889,N_29725);
and UO_2355 (O_2355,N_29055,N_28949);
nand UO_2356 (O_2356,N_25355,N_24299);
xor UO_2357 (O_2357,N_27407,N_24616);
or UO_2358 (O_2358,N_24075,N_26243);
or UO_2359 (O_2359,N_25991,N_24035);
and UO_2360 (O_2360,N_25462,N_25459);
nor UO_2361 (O_2361,N_29422,N_28863);
nand UO_2362 (O_2362,N_25198,N_24585);
xor UO_2363 (O_2363,N_24917,N_27173);
or UO_2364 (O_2364,N_29031,N_25293);
and UO_2365 (O_2365,N_27039,N_24519);
nand UO_2366 (O_2366,N_29545,N_28383);
xnor UO_2367 (O_2367,N_24481,N_26912);
or UO_2368 (O_2368,N_26217,N_28402);
nand UO_2369 (O_2369,N_24472,N_24224);
nor UO_2370 (O_2370,N_29358,N_27385);
nand UO_2371 (O_2371,N_29056,N_29556);
xor UO_2372 (O_2372,N_28676,N_25034);
xnor UO_2373 (O_2373,N_27765,N_24141);
xnor UO_2374 (O_2374,N_26821,N_27952);
or UO_2375 (O_2375,N_24486,N_27138);
nand UO_2376 (O_2376,N_28665,N_25134);
or UO_2377 (O_2377,N_24936,N_29733);
nor UO_2378 (O_2378,N_24747,N_26093);
and UO_2379 (O_2379,N_26530,N_28410);
xnor UO_2380 (O_2380,N_25176,N_27772);
and UO_2381 (O_2381,N_29696,N_28096);
xnor UO_2382 (O_2382,N_25996,N_25522);
nand UO_2383 (O_2383,N_28571,N_29215);
nand UO_2384 (O_2384,N_26916,N_26084);
nand UO_2385 (O_2385,N_24520,N_24794);
nor UO_2386 (O_2386,N_24845,N_29966);
xnor UO_2387 (O_2387,N_27808,N_27226);
nand UO_2388 (O_2388,N_27047,N_24303);
xnor UO_2389 (O_2389,N_27709,N_26026);
nand UO_2390 (O_2390,N_27807,N_24915);
nand UO_2391 (O_2391,N_26239,N_27586);
nor UO_2392 (O_2392,N_25357,N_24139);
nor UO_2393 (O_2393,N_27349,N_26071);
or UO_2394 (O_2394,N_27030,N_27493);
nand UO_2395 (O_2395,N_29640,N_26943);
and UO_2396 (O_2396,N_28224,N_24431);
xnor UO_2397 (O_2397,N_29045,N_24521);
and UO_2398 (O_2398,N_29673,N_28661);
and UO_2399 (O_2399,N_29390,N_26827);
nand UO_2400 (O_2400,N_24591,N_24529);
xnor UO_2401 (O_2401,N_28633,N_26686);
xnor UO_2402 (O_2402,N_25756,N_28145);
and UO_2403 (O_2403,N_25907,N_25767);
and UO_2404 (O_2404,N_29086,N_28102);
xnor UO_2405 (O_2405,N_24766,N_29662);
and UO_2406 (O_2406,N_29040,N_27967);
or UO_2407 (O_2407,N_24082,N_27067);
or UO_2408 (O_2408,N_26226,N_27947);
xor UO_2409 (O_2409,N_27044,N_25288);
nor UO_2410 (O_2410,N_24547,N_29636);
or UO_2411 (O_2411,N_28933,N_27757);
nand UO_2412 (O_2412,N_29306,N_27211);
nor UO_2413 (O_2413,N_29529,N_27531);
xor UO_2414 (O_2414,N_24290,N_29405);
xor UO_2415 (O_2415,N_28987,N_26199);
and UO_2416 (O_2416,N_24714,N_27711);
nor UO_2417 (O_2417,N_27021,N_26148);
xor UO_2418 (O_2418,N_26720,N_24688);
nand UO_2419 (O_2419,N_24362,N_27181);
and UO_2420 (O_2420,N_28856,N_25058);
xnor UO_2421 (O_2421,N_29439,N_28024);
and UO_2422 (O_2422,N_28575,N_27507);
and UO_2423 (O_2423,N_28817,N_24514);
nand UO_2424 (O_2424,N_28462,N_29718);
xnor UO_2425 (O_2425,N_27859,N_27116);
xnor UO_2426 (O_2426,N_29271,N_27233);
or UO_2427 (O_2427,N_28630,N_24577);
nor UO_2428 (O_2428,N_24960,N_29905);
or UO_2429 (O_2429,N_29135,N_28426);
nor UO_2430 (O_2430,N_28655,N_26560);
nor UO_2431 (O_2431,N_25855,N_28392);
nor UO_2432 (O_2432,N_27869,N_26424);
xnor UO_2433 (O_2433,N_24821,N_29848);
nand UO_2434 (O_2434,N_26831,N_25061);
or UO_2435 (O_2435,N_25562,N_27106);
or UO_2436 (O_2436,N_24740,N_24419);
nor UO_2437 (O_2437,N_28216,N_24778);
nor UO_2438 (O_2438,N_26616,N_27111);
and UO_2439 (O_2439,N_28335,N_29589);
nor UO_2440 (O_2440,N_29453,N_29174);
nand UO_2441 (O_2441,N_24434,N_26259);
or UO_2442 (O_2442,N_26802,N_25602);
and UO_2443 (O_2443,N_24626,N_24348);
and UO_2444 (O_2444,N_29270,N_29156);
and UO_2445 (O_2445,N_25388,N_29821);
or UO_2446 (O_2446,N_27382,N_29564);
nor UO_2447 (O_2447,N_29550,N_24574);
xor UO_2448 (O_2448,N_26060,N_26988);
xor UO_2449 (O_2449,N_28052,N_29080);
xor UO_2450 (O_2450,N_29340,N_25040);
nor UO_2451 (O_2451,N_26195,N_24801);
xnor UO_2452 (O_2452,N_29353,N_24503);
nand UO_2453 (O_2453,N_24024,N_26668);
or UO_2454 (O_2454,N_24005,N_29463);
and UO_2455 (O_2455,N_28452,N_25910);
nor UO_2456 (O_2456,N_25344,N_27494);
xor UO_2457 (O_2457,N_26615,N_24532);
nand UO_2458 (O_2458,N_28149,N_27232);
and UO_2459 (O_2459,N_26930,N_27078);
nand UO_2460 (O_2460,N_24536,N_29364);
xnor UO_2461 (O_2461,N_29461,N_28855);
xor UO_2462 (O_2462,N_27594,N_29525);
nand UO_2463 (O_2463,N_26875,N_26300);
nor UO_2464 (O_2464,N_25703,N_28371);
xor UO_2465 (O_2465,N_29273,N_28875);
and UO_2466 (O_2466,N_24366,N_26067);
nand UO_2467 (O_2467,N_28257,N_29291);
xor UO_2468 (O_2468,N_24063,N_25884);
nand UO_2469 (O_2469,N_24938,N_26685);
nand UO_2470 (O_2470,N_28343,N_28826);
nand UO_2471 (O_2471,N_29475,N_25971);
or UO_2472 (O_2472,N_27308,N_28748);
nand UO_2473 (O_2473,N_28313,N_25993);
nand UO_2474 (O_2474,N_25780,N_29626);
or UO_2475 (O_2475,N_28827,N_26154);
nand UO_2476 (O_2476,N_24361,N_27564);
nand UO_2477 (O_2477,N_26787,N_26692);
xnor UO_2478 (O_2478,N_24599,N_29168);
nor UO_2479 (O_2479,N_24832,N_29766);
nor UO_2480 (O_2480,N_24002,N_25482);
xnor UO_2481 (O_2481,N_25103,N_25283);
or UO_2482 (O_2482,N_29339,N_25677);
or UO_2483 (O_2483,N_27305,N_26838);
nand UO_2484 (O_2484,N_29682,N_24274);
nor UO_2485 (O_2485,N_24207,N_25640);
nor UO_2486 (O_2486,N_25443,N_28965);
nand UO_2487 (O_2487,N_25195,N_26905);
nor UO_2488 (O_2488,N_24055,N_27672);
or UO_2489 (O_2489,N_29501,N_25124);
and UO_2490 (O_2490,N_27841,N_28449);
and UO_2491 (O_2491,N_24746,N_25127);
or UO_2492 (O_2492,N_29805,N_26577);
nor UO_2493 (O_2493,N_29389,N_28325);
and UO_2494 (O_2494,N_28137,N_27117);
nor UO_2495 (O_2495,N_28668,N_25338);
nor UO_2496 (O_2496,N_28117,N_29754);
nand UO_2497 (O_2497,N_29146,N_27327);
nand UO_2498 (O_2498,N_28160,N_27157);
nand UO_2499 (O_2499,N_25167,N_24815);
or UO_2500 (O_2500,N_29454,N_24968);
nor UO_2501 (O_2501,N_24214,N_29591);
and UO_2502 (O_2502,N_24079,N_27180);
and UO_2503 (O_2503,N_29528,N_24116);
xnor UO_2504 (O_2504,N_28938,N_25613);
nor UO_2505 (O_2505,N_24377,N_25588);
xor UO_2506 (O_2506,N_29116,N_28780);
or UO_2507 (O_2507,N_29175,N_26120);
nand UO_2508 (O_2508,N_28399,N_24923);
nor UO_2509 (O_2509,N_25593,N_24958);
xor UO_2510 (O_2510,N_29289,N_24601);
or UO_2511 (O_2511,N_27079,N_28314);
xnor UO_2512 (O_2512,N_27987,N_25775);
nor UO_2513 (O_2513,N_26805,N_29794);
xor UO_2514 (O_2514,N_25782,N_26733);
nand UO_2515 (O_2515,N_27300,N_29379);
xor UO_2516 (O_2516,N_25431,N_28807);
and UO_2517 (O_2517,N_28852,N_28872);
xnor UO_2518 (O_2518,N_29657,N_28014);
and UO_2519 (O_2519,N_24657,N_26049);
nand UO_2520 (O_2520,N_24376,N_29702);
nand UO_2521 (O_2521,N_27304,N_29936);
or UO_2522 (O_2522,N_26989,N_25185);
nand UO_2523 (O_2523,N_28645,N_28577);
and UO_2524 (O_2524,N_24712,N_26748);
and UO_2525 (O_2525,N_25452,N_28113);
or UO_2526 (O_2526,N_28623,N_27624);
and UO_2527 (O_2527,N_29107,N_26630);
nand UO_2528 (O_2528,N_25472,N_24659);
xnor UO_2529 (O_2529,N_25013,N_28769);
nor UO_2530 (O_2530,N_25520,N_25914);
or UO_2531 (O_2531,N_25518,N_25968);
nand UO_2532 (O_2532,N_29926,N_25551);
nor UO_2533 (O_2533,N_24168,N_28917);
and UO_2534 (O_2534,N_26227,N_27676);
xnor UO_2535 (O_2535,N_28107,N_29301);
nand UO_2536 (O_2536,N_29757,N_26194);
xnor UO_2537 (O_2537,N_28100,N_28316);
xnor UO_2538 (O_2538,N_29709,N_24439);
and UO_2539 (O_2539,N_29434,N_25300);
nand UO_2540 (O_2540,N_29732,N_29037);
nand UO_2541 (O_2541,N_27183,N_25707);
xnor UO_2542 (O_2542,N_29014,N_28594);
xor UO_2543 (O_2543,N_28640,N_28453);
nor UO_2544 (O_2544,N_25049,N_28397);
xnor UO_2545 (O_2545,N_29319,N_26659);
nor UO_2546 (O_2546,N_27399,N_29876);
nand UO_2547 (O_2547,N_29512,N_26171);
xnor UO_2548 (O_2548,N_24976,N_29426);
or UO_2549 (O_2549,N_24819,N_25505);
nand UO_2550 (O_2550,N_25233,N_27285);
xnor UO_2551 (O_2551,N_24818,N_24882);
nor UO_2552 (O_2552,N_25747,N_25692);
xor UO_2553 (O_2553,N_24329,N_25680);
nor UO_2554 (O_2554,N_25220,N_25202);
or UO_2555 (O_2555,N_27538,N_28187);
nand UO_2556 (O_2556,N_28845,N_28560);
or UO_2557 (O_2557,N_24169,N_29421);
nor UO_2558 (O_2558,N_25382,N_29871);
xnor UO_2559 (O_2559,N_25874,N_26627);
nor UO_2560 (O_2560,N_25025,N_24744);
or UO_2561 (O_2561,N_26752,N_27000);
or UO_2562 (O_2562,N_29078,N_25352);
nor UO_2563 (O_2563,N_26132,N_25313);
xor UO_2564 (O_2564,N_27925,N_26646);
nand UO_2565 (O_2565,N_24986,N_25168);
or UO_2566 (O_2566,N_26484,N_29257);
nand UO_2567 (O_2567,N_25679,N_27057);
xnor UO_2568 (O_2568,N_29165,N_29149);
nor UO_2569 (O_2569,N_29753,N_25050);
xnor UO_2570 (O_2570,N_25139,N_24490);
and UO_2571 (O_2571,N_28444,N_28451);
nor UO_2572 (O_2572,N_29971,N_24287);
and UO_2573 (O_2573,N_24872,N_27849);
xnor UO_2574 (O_2574,N_28228,N_25347);
and UO_2575 (O_2575,N_26667,N_28693);
and UO_2576 (O_2576,N_27761,N_28384);
or UO_2577 (O_2577,N_26658,N_28919);
or UO_2578 (O_2578,N_27169,N_24606);
or UO_2579 (O_2579,N_25371,N_27420);
xor UO_2580 (O_2580,N_27128,N_25320);
nor UO_2581 (O_2581,N_25287,N_29880);
nor UO_2582 (O_2582,N_25962,N_25010);
nand UO_2583 (O_2583,N_27129,N_25282);
nor UO_2584 (O_2584,N_26819,N_25499);
and UO_2585 (O_2585,N_26529,N_26232);
and UO_2586 (O_2586,N_28265,N_25867);
nand UO_2587 (O_2587,N_24371,N_27654);
nand UO_2588 (O_2588,N_29565,N_26506);
nor UO_2589 (O_2589,N_25331,N_26729);
and UO_2590 (O_2590,N_29765,N_24219);
xor UO_2591 (O_2591,N_25618,N_24581);
or UO_2592 (O_2592,N_26166,N_25862);
xnor UO_2593 (O_2593,N_29131,N_28270);
nand UO_2594 (O_2594,N_24269,N_24105);
xor UO_2595 (O_2595,N_25082,N_27921);
and UO_2596 (O_2596,N_26220,N_28105);
and UO_2597 (O_2597,N_26793,N_28755);
or UO_2598 (O_2598,N_28507,N_24967);
nand UO_2599 (O_2599,N_29125,N_28975);
xnor UO_2600 (O_2600,N_24370,N_29731);
nand UO_2601 (O_2601,N_29377,N_27674);
nor UO_2602 (O_2602,N_27817,N_29087);
nand UO_2603 (O_2603,N_27589,N_25623);
or UO_2604 (O_2604,N_29774,N_25009);
xor UO_2605 (O_2605,N_27780,N_25514);
xnor UO_2606 (O_2606,N_25004,N_26448);
nor UO_2607 (O_2607,N_25322,N_24074);
nor UO_2608 (O_2608,N_29419,N_28947);
nor UO_2609 (O_2609,N_26355,N_25078);
nor UO_2610 (O_2610,N_24763,N_25838);
and UO_2611 (O_2611,N_24602,N_25708);
or UO_2612 (O_2612,N_26680,N_24692);
and UO_2613 (O_2613,N_24946,N_29425);
nand UO_2614 (O_2614,N_24354,N_28980);
nor UO_2615 (O_2615,N_26651,N_28063);
or UO_2616 (O_2616,N_28519,N_26121);
nand UO_2617 (O_2617,N_28624,N_24587);
and UO_2618 (O_2618,N_25879,N_24268);
nor UO_2619 (O_2619,N_29348,N_27184);
and UO_2620 (O_2620,N_26414,N_24638);
or UO_2621 (O_2621,N_25858,N_25333);
nand UO_2622 (O_2622,N_25354,N_28666);
nor UO_2623 (O_2623,N_26963,N_29083);
nor UO_2624 (O_2624,N_29834,N_27071);
or UO_2625 (O_2625,N_29308,N_27502);
or UO_2626 (O_2626,N_26742,N_24238);
nor UO_2627 (O_2627,N_26757,N_26216);
or UO_2628 (O_2628,N_24674,N_28540);
nand UO_2629 (O_2629,N_25245,N_24901);
and UO_2630 (O_2630,N_29633,N_28964);
nand UO_2631 (O_2631,N_26133,N_27962);
or UO_2632 (O_2632,N_28407,N_28525);
or UO_2633 (O_2633,N_29456,N_25715);
nor UO_2634 (O_2634,N_25397,N_29910);
nor UO_2635 (O_2635,N_26601,N_25474);
nor UO_2636 (O_2636,N_28694,N_25880);
and UO_2637 (O_2637,N_29436,N_28043);
and UO_2638 (O_2638,N_25193,N_24834);
nand UO_2639 (O_2639,N_27801,N_26383);
nor UO_2640 (O_2640,N_26671,N_26809);
nand UO_2641 (O_2641,N_24270,N_28834);
nand UO_2642 (O_2642,N_25972,N_27563);
xor UO_2643 (O_2643,N_24198,N_29094);
nand UO_2644 (O_2644,N_29915,N_28290);
and UO_2645 (O_2645,N_25317,N_29901);
nand UO_2646 (O_2646,N_27095,N_29547);
and UO_2647 (O_2647,N_26082,N_29384);
nand UO_2648 (O_2648,N_25591,N_25727);
or UO_2649 (O_2649,N_24624,N_24677);
and UO_2650 (O_2650,N_28207,N_24910);
and UO_2651 (O_2651,N_25959,N_28183);
or UO_2652 (O_2652,N_27115,N_26376);
nand UO_2653 (O_2653,N_24993,N_26737);
or UO_2654 (O_2654,N_26293,N_29913);
xnor UO_2655 (O_2655,N_25154,N_26064);
xnor UO_2656 (O_2656,N_25038,N_27659);
xor UO_2657 (O_2657,N_29288,N_28719);
nand UO_2658 (O_2658,N_24165,N_26515);
nor UO_2659 (O_2659,N_24478,N_29404);
xor UO_2660 (O_2660,N_27878,N_27959);
nand UO_2661 (O_2661,N_26540,N_26960);
or UO_2662 (O_2662,N_28546,N_29296);
and UO_2663 (O_2663,N_27472,N_24840);
or UO_2664 (O_2664,N_24330,N_28604);
nand UO_2665 (O_2665,N_24153,N_27964);
and UO_2666 (O_2666,N_28679,N_29987);
nand UO_2667 (O_2667,N_28909,N_25995);
xor UO_2668 (O_2668,N_27141,N_29173);
nor UO_2669 (O_2669,N_26275,N_25595);
xor UO_2670 (O_2670,N_27883,N_28911);
xor UO_2671 (O_2671,N_24684,N_29499);
or UO_2672 (O_2672,N_27641,N_26413);
xor UO_2673 (O_2673,N_26723,N_28818);
nor UO_2674 (O_2674,N_29137,N_27891);
nor UO_2675 (O_2675,N_27668,N_27229);
and UO_2676 (O_2676,N_25964,N_24150);
nand UO_2677 (O_2677,N_26045,N_26333);
nand UO_2678 (O_2678,N_27621,N_29616);
and UO_2679 (O_2679,N_26125,N_26653);
and UO_2680 (O_2680,N_25467,N_26998);
nor UO_2681 (O_2681,N_26794,N_26815);
or UO_2682 (O_2682,N_28802,N_28805);
nand UO_2683 (O_2683,N_29986,N_28495);
nand UO_2684 (O_2684,N_29408,N_29245);
nand UO_2685 (O_2685,N_29778,N_26936);
nor UO_2686 (O_2686,N_27893,N_29667);
nor UO_2687 (O_2687,N_29559,N_25425);
and UO_2688 (O_2688,N_26313,N_27504);
and UO_2689 (O_2689,N_27491,N_28820);
xor UO_2690 (O_2690,N_29828,N_25844);
nor UO_2691 (O_2691,N_29592,N_26405);
and UO_2692 (O_2692,N_25265,N_27906);
nor UO_2693 (O_2693,N_25863,N_28123);
nor UO_2694 (O_2694,N_29274,N_27749);
nor UO_2695 (O_2695,N_24367,N_27982);
xnor UO_2696 (O_2696,N_29117,N_27070);
or UO_2697 (O_2697,N_26365,N_28512);
or UO_2698 (O_2698,N_25678,N_28181);
nor UO_2699 (O_2699,N_28415,N_24250);
xnor UO_2700 (O_2700,N_29263,N_24273);
xnor UO_2701 (O_2701,N_25975,N_27644);
nand UO_2702 (O_2702,N_29967,N_26229);
nand UO_2703 (O_2703,N_24673,N_26412);
nor UO_2704 (O_2704,N_27040,N_29792);
nor UO_2705 (O_2705,N_29507,N_27168);
or UO_2706 (O_2706,N_26964,N_26029);
or UO_2707 (O_2707,N_28279,N_26249);
nand UO_2708 (O_2708,N_26009,N_26015);
nor UO_2709 (O_2709,N_26372,N_28635);
and UO_2710 (O_2710,N_26575,N_27689);
nor UO_2711 (O_2711,N_29294,N_29868);
and UO_2712 (O_2712,N_24656,N_26706);
or UO_2713 (O_2713,N_25960,N_28765);
nor UO_2714 (O_2714,N_28150,N_29445);
or UO_2715 (O_2715,N_25209,N_24340);
nand UO_2716 (O_2716,N_24781,N_26561);
or UO_2717 (O_2717,N_26639,N_26797);
nor UO_2718 (O_2718,N_24851,N_28870);
xor UO_2719 (O_2719,N_26526,N_29011);
xor UO_2720 (O_2720,N_24694,N_25967);
or UO_2721 (O_2721,N_29768,N_29860);
xor UO_2722 (O_2722,N_28230,N_24990);
nor UO_2723 (O_2723,N_27631,N_26415);
and UO_2724 (O_2724,N_27132,N_25965);
xor UO_2725 (O_2725,N_27083,N_24128);
and UO_2726 (O_2726,N_29120,N_29285);
and UO_2727 (O_2727,N_24010,N_28529);
nand UO_2728 (O_2728,N_27916,N_25298);
nand UO_2729 (O_2729,N_27685,N_27732);
nand UO_2730 (O_2730,N_24483,N_29189);
nand UO_2731 (O_2731,N_27166,N_25924);
and UO_2732 (O_2732,N_25484,N_25123);
or UO_2733 (O_2733,N_29391,N_26459);
and UO_2734 (O_2734,N_28015,N_29776);
or UO_2735 (O_2735,N_26388,N_27978);
xnor UO_2736 (O_2736,N_28469,N_28192);
xor UO_2737 (O_2737,N_25689,N_25870);
nand UO_2738 (O_2738,N_27665,N_28619);
or UO_2739 (O_2739,N_24408,N_25846);
and UO_2740 (O_2740,N_26693,N_28536);
xnor UO_2741 (O_2741,N_25615,N_29365);
and UO_2742 (O_2742,N_24767,N_27610);
xor UO_2743 (O_2743,N_25172,N_27393);
xnor UO_2744 (O_2744,N_25662,N_26172);
nand UO_2745 (O_2745,N_28450,N_25239);
and UO_2746 (O_2746,N_26050,N_28784);
xor UO_2747 (O_2747,N_25808,N_27398);
nor UO_2748 (O_2748,N_29142,N_29228);
nand UO_2749 (O_2749,N_26628,N_25852);
and UO_2750 (O_2750,N_27366,N_28283);
nand UO_2751 (O_2751,N_28292,N_26481);
xnor UO_2752 (O_2752,N_28256,N_29777);
nor UO_2753 (O_2753,N_25000,N_26721);
or UO_2754 (O_2754,N_25653,N_29963);
or UO_2755 (O_2755,N_25875,N_25007);
and UO_2756 (O_2756,N_27511,N_24265);
and UO_2757 (O_2757,N_26820,N_25980);
nand UO_2758 (O_2758,N_24572,N_25890);
xor UO_2759 (O_2759,N_24619,N_26041);
nand UO_2760 (O_2760,N_25094,N_27062);
or UO_2761 (O_2761,N_28642,N_24732);
xor UO_2762 (O_2762,N_28697,N_26611);
nor UO_2763 (O_2763,N_26854,N_24412);
nor UO_2764 (O_2764,N_28057,N_28907);
xnor UO_2765 (O_2765,N_24435,N_28543);
xor UO_2766 (O_2766,N_27441,N_24427);
nand UO_2767 (O_2767,N_29830,N_25440);
nand UO_2768 (O_2768,N_24051,N_28498);
xnor UO_2769 (O_2769,N_26839,N_27343);
nor UO_2770 (O_2770,N_29412,N_27192);
and UO_2771 (O_2771,N_28555,N_28082);
xor UO_2772 (O_2772,N_27182,N_27933);
or UO_2773 (O_2773,N_27911,N_29327);
nor UO_2774 (O_2774,N_28641,N_25143);
nor UO_2775 (O_2775,N_27251,N_26914);
and UO_2776 (O_2776,N_28848,N_27771);
and UO_2777 (O_2777,N_24875,N_28702);
and UO_2778 (O_2778,N_27838,N_28809);
xnor UO_2779 (O_2779,N_26393,N_26267);
nor UO_2780 (O_2780,N_28227,N_28520);
nor UO_2781 (O_2781,N_29837,N_27805);
xor UO_2782 (O_2782,N_27549,N_25496);
nor UO_2783 (O_2783,N_27159,N_26209);
xor UO_2784 (O_2784,N_28862,N_28912);
or UO_2785 (O_2785,N_28020,N_24038);
nor UO_2786 (O_2786,N_29687,N_27741);
nor UO_2787 (O_2787,N_28271,N_24853);
nand UO_2788 (O_2788,N_28463,N_24489);
nor UO_2789 (O_2789,N_27767,N_28692);
xnor UO_2790 (O_2790,N_29025,N_24429);
or UO_2791 (O_2791,N_27949,N_24450);
and UO_2792 (O_2792,N_29530,N_28485);
nor UO_2793 (O_2793,N_26116,N_27195);
xor UO_2794 (O_2794,N_29937,N_27702);
nand UO_2795 (O_2795,N_25289,N_26240);
and UO_2796 (O_2796,N_26605,N_27094);
and UO_2797 (O_2797,N_25057,N_24891);
nor UO_2798 (O_2798,N_27492,N_29867);
nor UO_2799 (O_2799,N_27551,N_25132);
nand UO_2800 (O_2800,N_25561,N_29162);
and UO_2801 (O_2801,N_27274,N_29576);
or UO_2802 (O_2802,N_25903,N_27896);
or UO_2803 (O_2803,N_25726,N_27894);
nor UO_2804 (O_2804,N_26406,N_25503);
and UO_2805 (O_2805,N_28341,N_26228);
nor UO_2806 (O_2806,N_27176,N_28263);
nor UO_2807 (O_2807,N_29607,N_25272);
or UO_2808 (O_2808,N_27524,N_24272);
or UO_2809 (O_2809,N_29007,N_29985);
and UO_2810 (O_2810,N_26014,N_24697);
and UO_2811 (O_2811,N_26760,N_25569);
and UO_2812 (O_2812,N_28565,N_28310);
nor UO_2813 (O_2813,N_29504,N_27389);
nor UO_2814 (O_2814,N_26589,N_29170);
xnor UO_2815 (O_2815,N_28610,N_24554);
nand UO_2816 (O_2816,N_26590,N_26175);
and UO_2817 (O_2817,N_29909,N_25488);
and UO_2818 (O_2818,N_29706,N_26759);
and UO_2819 (O_2819,N_29505,N_27786);
nand UO_2820 (O_2820,N_29749,N_24894);
or UO_2821 (O_2821,N_29220,N_24034);
nor UO_2822 (O_2822,N_28409,N_26461);
nor UO_2823 (O_2823,N_25019,N_29981);
nand UO_2824 (O_2824,N_28420,N_28718);
or UO_2825 (O_2825,N_28631,N_28413);
xor UO_2826 (O_2826,N_25434,N_24709);
nand UO_2827 (O_2827,N_24857,N_24669);
nand UO_2828 (O_2828,N_24822,N_28729);
nor UO_2829 (O_2829,N_27310,N_27320);
nand UO_2830 (O_2830,N_27973,N_28854);
and UO_2831 (O_2831,N_27821,N_29844);
and UO_2832 (O_2832,N_25646,N_28101);
nor UO_2833 (O_2833,N_29185,N_28833);
xor UO_2834 (O_2834,N_29744,N_27816);
and UO_2835 (O_2835,N_26527,N_27395);
or UO_2836 (O_2836,N_27032,N_24323);
nand UO_2837 (O_2837,N_26238,N_24159);
and UO_2838 (O_2838,N_26997,N_26750);
or UO_2839 (O_2839,N_28728,N_25816);
nor UO_2840 (O_2840,N_26765,N_28573);
nor UO_2841 (O_2841,N_25267,N_27919);
nor UO_2842 (O_2842,N_26031,N_24069);
nand UO_2843 (O_2843,N_29399,N_28215);
nor UO_2844 (O_2844,N_25524,N_29495);
nand UO_2845 (O_2845,N_29180,N_24839);
nand UO_2846 (O_2846,N_29265,N_27604);
or UO_2847 (O_2847,N_24609,N_28433);
or UO_2848 (O_2848,N_27072,N_25075);
and UO_2849 (O_2849,N_29922,N_27864);
xor UO_2850 (O_2850,N_25157,N_27303);
and UO_2851 (O_2851,N_24189,N_26113);
and UO_2852 (O_2852,N_28950,N_26065);
and UO_2853 (O_2853,N_25807,N_26335);
xor UO_2854 (O_2854,N_25241,N_28582);
or UO_2855 (O_2855,N_27413,N_29595);
and UO_2856 (O_2856,N_27276,N_29000);
xor UO_2857 (O_2857,N_25786,N_26804);
nand UO_2858 (O_2858,N_25930,N_28329);
or UO_2859 (O_2859,N_26010,N_24713);
xor UO_2860 (O_2860,N_29551,N_28782);
and UO_2861 (O_2861,N_24102,N_24666);
and UO_2862 (O_2862,N_29370,N_27693);
and UO_2863 (O_2863,N_24773,N_27646);
nand UO_2864 (O_2864,N_29610,N_26051);
nand UO_2865 (O_2865,N_27660,N_26873);
or UO_2866 (O_2866,N_25676,N_29347);
nand UO_2867 (O_2867,N_24073,N_26634);
nor UO_2868 (O_2868,N_29912,N_24907);
and UO_2869 (O_2869,N_26638,N_26462);
xor UO_2870 (O_2870,N_29533,N_26887);
nor UO_2871 (O_2871,N_25253,N_27179);
nor UO_2872 (O_2872,N_25362,N_25568);
nor UO_2873 (O_2873,N_27508,N_24056);
xor UO_2874 (O_2874,N_29198,N_26312);
nand UO_2875 (O_2875,N_25432,N_27583);
nand UO_2876 (O_2876,N_24973,N_24132);
nor UO_2877 (O_2877,N_27569,N_27506);
or UO_2878 (O_2878,N_28472,N_26637);
nor UO_2879 (O_2879,N_28940,N_27983);
nor UO_2880 (O_2880,N_27421,N_26626);
nand UO_2881 (O_2881,N_28725,N_29150);
and UO_2882 (O_2882,N_29022,N_25394);
nor UO_2883 (O_2883,N_24426,N_28787);
or UO_2884 (O_2884,N_25194,N_29297);
nor UO_2885 (O_2885,N_24945,N_25119);
and UO_2886 (O_2886,N_27892,N_27088);
or UO_2887 (O_2887,N_28210,N_24630);
and UO_2888 (O_2888,N_24112,N_28296);
nor UO_2889 (O_2889,N_28795,N_24231);
nor UO_2890 (O_2890,N_24254,N_29491);
xor UO_2891 (O_2891,N_29898,N_27218);
and UO_2892 (O_2892,N_28868,N_26981);
or UO_2893 (O_2893,N_26937,N_27769);
nand UO_2894 (O_2894,N_28763,N_29887);
or UO_2895 (O_2895,N_24728,N_27768);
and UO_2896 (O_2896,N_26661,N_29159);
or UO_2897 (O_2897,N_26485,N_29249);
xnor UO_2898 (O_2898,N_26741,N_29929);
or UO_2899 (O_2899,N_26841,N_25426);
nand UO_2900 (O_2900,N_24298,N_26301);
or UO_2901 (O_2901,N_28396,N_27383);
and UO_2902 (O_2902,N_27984,N_27367);
xnor UO_2903 (O_2903,N_27532,N_24559);
xnor UO_2904 (O_2904,N_29553,N_28527);
or UO_2905 (O_2905,N_28391,N_24862);
xnor UO_2906 (O_2906,N_24561,N_26953);
nor UO_2907 (O_2907,N_26597,N_27488);
and UO_2908 (O_2908,N_25901,N_24470);
and UO_2909 (O_2909,N_29300,N_27190);
nand UO_2910 (O_2910,N_28681,N_29305);
xor UO_2911 (O_2911,N_24573,N_27691);
and UO_2912 (O_2912,N_24680,N_24643);
or UO_2913 (O_2913,N_25741,N_27832);
nand UO_2914 (O_2914,N_29409,N_28166);
or UO_2915 (O_2915,N_25906,N_25230);
and UO_2916 (O_2916,N_24777,N_27315);
and UO_2917 (O_2917,N_27219,N_26326);
and UO_2918 (O_2918,N_24860,N_26464);
nand UO_2919 (O_2919,N_26849,N_26747);
or UO_2920 (O_2920,N_25566,N_27596);
xor UO_2921 (O_2921,N_24137,N_29902);
and UO_2922 (O_2922,N_29716,N_28095);
or UO_2923 (O_2923,N_24909,N_25039);
xor UO_2924 (O_2924,N_27352,N_24175);
or UO_2925 (O_2925,N_28847,N_26439);
nand UO_2926 (O_2926,N_24689,N_29062);
and UO_2927 (O_2927,N_25097,N_27381);
nand UO_2928 (O_2928,N_27379,N_29698);
and UO_2929 (O_2929,N_24205,N_28434);
nor UO_2930 (O_2930,N_28617,N_25182);
and UO_2931 (O_2931,N_27360,N_28189);
nand UO_2932 (O_2932,N_25508,N_27107);
or UO_2933 (O_2933,N_25791,N_28066);
or UO_2934 (O_2934,N_27550,N_26419);
and UO_2935 (O_2935,N_29977,N_29631);
nand UO_2936 (O_2936,N_27301,N_27663);
nor UO_2937 (O_2937,N_27291,N_28841);
and UO_2938 (O_2938,N_27087,N_27186);
xor UO_2939 (O_2939,N_26773,N_24795);
or UO_2940 (O_2940,N_28186,N_25153);
or UO_2941 (O_2941,N_29539,N_24147);
nand UO_2942 (O_2942,N_27137,N_25868);
nor UO_2943 (O_2943,N_26707,N_24653);
and UO_2944 (O_2944,N_27430,N_25307);
and UO_2945 (O_2945,N_24589,N_25001);
xor UO_2946 (O_2946,N_26826,N_24804);
or UO_2947 (O_2947,N_27297,N_26285);
nand UO_2948 (O_2948,N_25935,N_26911);
or UO_2949 (O_2949,N_27258,N_27326);
nor UO_2950 (O_2950,N_24030,N_27535);
nor UO_2951 (O_2951,N_28929,N_29542);
and UO_2952 (O_2952,N_27628,N_28886);
or UO_2953 (O_2953,N_26962,N_24480);
nor UO_2954 (O_2954,N_28195,N_27729);
and UO_2955 (O_2955,N_29351,N_26225);
xor UO_2956 (O_2956,N_27011,N_27778);
nand UO_2957 (O_2957,N_28045,N_24278);
nand UO_2958 (O_2958,N_29017,N_26477);
nand UO_2959 (O_2959,N_26445,N_28111);
or UO_2960 (O_2960,N_24037,N_27824);
nor UO_2961 (O_2961,N_27453,N_27866);
or UO_2962 (O_2962,N_26303,N_24949);
or UO_2963 (O_2963,N_29973,N_25544);
nand UO_2964 (O_2964,N_28632,N_28418);
nand UO_2965 (O_2965,N_28010,N_25717);
nor UO_2966 (O_2966,N_27796,N_24386);
nand UO_2967 (O_2967,N_29920,N_24846);
nand UO_2968 (O_2968,N_27016,N_25341);
nand UO_2969 (O_2969,N_24652,N_25826);
and UO_2970 (O_2970,N_24776,N_26241);
nand UO_2971 (O_2971,N_27114,N_24703);
xor UO_2972 (O_2972,N_24784,N_28877);
and UO_2973 (O_2973,N_27294,N_26591);
and UO_2974 (O_2974,N_29324,N_29147);
or UO_2975 (O_2975,N_26897,N_27931);
xor UO_2976 (O_2976,N_26119,N_29352);
xor UO_2977 (O_2977,N_28798,N_24880);
or UO_2978 (O_2978,N_24717,N_28042);
xnor UO_2979 (O_2979,N_25349,N_27100);
xor UO_2980 (O_2980,N_28776,N_28086);
nor UO_2981 (O_2981,N_28897,N_25793);
xor UO_2982 (O_2982,N_26156,N_27338);
and UO_2983 (O_2983,N_24942,N_27885);
or UO_2984 (O_2984,N_29184,N_27599);
and UO_2985 (O_2985,N_29293,N_27185);
nand UO_2986 (O_2986,N_24453,N_26735);
or UO_2987 (O_2987,N_27279,N_24241);
xnor UO_2988 (O_2988,N_27063,N_29158);
nor UO_2989 (O_2989,N_26266,N_25951);
nor UO_2990 (O_2990,N_27296,N_27035);
nor UO_2991 (O_2991,N_25758,N_25763);
or UO_2992 (O_2992,N_28698,N_29279);
nand UO_2993 (O_2993,N_28716,N_25433);
nor UO_2994 (O_2994,N_26468,N_28881);
nor UO_2995 (O_2995,N_27670,N_29199);
nor UO_2996 (O_2996,N_27001,N_28598);
or UO_2997 (O_2997,N_25915,N_26906);
nor UO_2998 (O_2998,N_24929,N_29584);
or UO_2999 (O_2999,N_24387,N_24843);
nand UO_3000 (O_3000,N_28169,N_24558);
nor UO_3001 (O_3001,N_26171,N_27958);
and UO_3002 (O_3002,N_27017,N_24142);
or UO_3003 (O_3003,N_27927,N_26708);
and UO_3004 (O_3004,N_28425,N_27612);
or UO_3005 (O_3005,N_28609,N_26102);
or UO_3006 (O_3006,N_24422,N_27068);
nor UO_3007 (O_3007,N_26971,N_26746);
xor UO_3008 (O_3008,N_29456,N_24474);
or UO_3009 (O_3009,N_25998,N_27585);
or UO_3010 (O_3010,N_25381,N_25083);
xor UO_3011 (O_3011,N_25072,N_24258);
nand UO_3012 (O_3012,N_24385,N_27937);
nor UO_3013 (O_3013,N_25578,N_29803);
xnor UO_3014 (O_3014,N_29234,N_26819);
and UO_3015 (O_3015,N_28181,N_27334);
or UO_3016 (O_3016,N_29896,N_29834);
nor UO_3017 (O_3017,N_24383,N_24132);
or UO_3018 (O_3018,N_24234,N_25581);
nor UO_3019 (O_3019,N_29075,N_25240);
xnor UO_3020 (O_3020,N_24103,N_26463);
and UO_3021 (O_3021,N_24480,N_25212);
xor UO_3022 (O_3022,N_27281,N_25792);
and UO_3023 (O_3023,N_29208,N_24194);
xor UO_3024 (O_3024,N_29468,N_26279);
nand UO_3025 (O_3025,N_28671,N_29097);
nor UO_3026 (O_3026,N_29293,N_29993);
xnor UO_3027 (O_3027,N_28079,N_26405);
nor UO_3028 (O_3028,N_29633,N_28564);
nor UO_3029 (O_3029,N_29985,N_28908);
or UO_3030 (O_3030,N_25810,N_24112);
nor UO_3031 (O_3031,N_24575,N_24342);
and UO_3032 (O_3032,N_29913,N_26838);
or UO_3033 (O_3033,N_26704,N_24809);
nor UO_3034 (O_3034,N_29102,N_25526);
nand UO_3035 (O_3035,N_28108,N_25811);
or UO_3036 (O_3036,N_29189,N_28651);
nor UO_3037 (O_3037,N_28186,N_25933);
xnor UO_3038 (O_3038,N_29534,N_26993);
xnor UO_3039 (O_3039,N_27313,N_28674);
nor UO_3040 (O_3040,N_24006,N_24455);
xor UO_3041 (O_3041,N_26853,N_26130);
nor UO_3042 (O_3042,N_24056,N_29096);
xnor UO_3043 (O_3043,N_27636,N_26711);
xor UO_3044 (O_3044,N_29663,N_29767);
xnor UO_3045 (O_3045,N_27311,N_29147);
xor UO_3046 (O_3046,N_24178,N_29511);
nor UO_3047 (O_3047,N_25695,N_25529);
xor UO_3048 (O_3048,N_28711,N_24560);
nand UO_3049 (O_3049,N_26619,N_26707);
nand UO_3050 (O_3050,N_25460,N_24060);
xnor UO_3051 (O_3051,N_28372,N_26096);
and UO_3052 (O_3052,N_26696,N_26063);
nand UO_3053 (O_3053,N_29241,N_28546);
or UO_3054 (O_3054,N_25956,N_27601);
nand UO_3055 (O_3055,N_26580,N_25004);
nand UO_3056 (O_3056,N_29474,N_25790);
or UO_3057 (O_3057,N_27301,N_24977);
and UO_3058 (O_3058,N_28277,N_26375);
xor UO_3059 (O_3059,N_29992,N_29731);
xor UO_3060 (O_3060,N_28441,N_26078);
and UO_3061 (O_3061,N_26094,N_27074);
or UO_3062 (O_3062,N_26731,N_27357);
nor UO_3063 (O_3063,N_29993,N_29365);
and UO_3064 (O_3064,N_26014,N_28584);
or UO_3065 (O_3065,N_27251,N_26562);
nor UO_3066 (O_3066,N_29206,N_29370);
xnor UO_3067 (O_3067,N_26460,N_27987);
or UO_3068 (O_3068,N_24010,N_29863);
nor UO_3069 (O_3069,N_29526,N_28332);
nand UO_3070 (O_3070,N_29875,N_28420);
nand UO_3071 (O_3071,N_24486,N_27222);
or UO_3072 (O_3072,N_24587,N_28345);
xor UO_3073 (O_3073,N_28289,N_25431);
or UO_3074 (O_3074,N_25516,N_25931);
or UO_3075 (O_3075,N_25652,N_28117);
nor UO_3076 (O_3076,N_24580,N_29251);
xnor UO_3077 (O_3077,N_27198,N_29594);
or UO_3078 (O_3078,N_29141,N_25000);
xor UO_3079 (O_3079,N_25500,N_28492);
xor UO_3080 (O_3080,N_27741,N_27787);
nor UO_3081 (O_3081,N_26039,N_24057);
nor UO_3082 (O_3082,N_27119,N_25130);
nor UO_3083 (O_3083,N_25164,N_28013);
nor UO_3084 (O_3084,N_26998,N_29767);
nand UO_3085 (O_3085,N_28789,N_25741);
nor UO_3086 (O_3086,N_26672,N_29349);
nor UO_3087 (O_3087,N_24485,N_26810);
nor UO_3088 (O_3088,N_24373,N_29292);
nand UO_3089 (O_3089,N_27560,N_24848);
nand UO_3090 (O_3090,N_25374,N_24404);
nand UO_3091 (O_3091,N_25166,N_29908);
or UO_3092 (O_3092,N_28914,N_27000);
or UO_3093 (O_3093,N_29410,N_29115);
or UO_3094 (O_3094,N_26400,N_26182);
and UO_3095 (O_3095,N_27600,N_25959);
and UO_3096 (O_3096,N_29467,N_29894);
xnor UO_3097 (O_3097,N_27728,N_29507);
and UO_3098 (O_3098,N_24247,N_26793);
and UO_3099 (O_3099,N_26656,N_29643);
and UO_3100 (O_3100,N_27110,N_25222);
and UO_3101 (O_3101,N_27910,N_24064);
and UO_3102 (O_3102,N_29231,N_25134);
nand UO_3103 (O_3103,N_28074,N_28052);
nor UO_3104 (O_3104,N_29613,N_25854);
and UO_3105 (O_3105,N_26196,N_28562);
and UO_3106 (O_3106,N_28530,N_27657);
nand UO_3107 (O_3107,N_24535,N_27241);
or UO_3108 (O_3108,N_25868,N_27619);
or UO_3109 (O_3109,N_25241,N_27521);
or UO_3110 (O_3110,N_27921,N_27765);
nand UO_3111 (O_3111,N_24661,N_24947);
xnor UO_3112 (O_3112,N_24029,N_29183);
or UO_3113 (O_3113,N_24239,N_26777);
nor UO_3114 (O_3114,N_29583,N_24009);
nand UO_3115 (O_3115,N_26667,N_28689);
xnor UO_3116 (O_3116,N_28067,N_28905);
nor UO_3117 (O_3117,N_25807,N_27384);
or UO_3118 (O_3118,N_25980,N_29310);
nor UO_3119 (O_3119,N_27291,N_29677);
xor UO_3120 (O_3120,N_27768,N_28168);
or UO_3121 (O_3121,N_24576,N_26088);
or UO_3122 (O_3122,N_24886,N_27140);
nand UO_3123 (O_3123,N_24466,N_24064);
or UO_3124 (O_3124,N_29739,N_26602);
nand UO_3125 (O_3125,N_27326,N_29890);
and UO_3126 (O_3126,N_26075,N_27468);
or UO_3127 (O_3127,N_24839,N_25790);
xor UO_3128 (O_3128,N_28478,N_25563);
xnor UO_3129 (O_3129,N_28982,N_26801);
or UO_3130 (O_3130,N_27115,N_28395);
or UO_3131 (O_3131,N_26577,N_28398);
or UO_3132 (O_3132,N_24466,N_27139);
xnor UO_3133 (O_3133,N_24952,N_28819);
or UO_3134 (O_3134,N_24566,N_28932);
and UO_3135 (O_3135,N_25418,N_28466);
and UO_3136 (O_3136,N_25935,N_26036);
nand UO_3137 (O_3137,N_24491,N_28478);
or UO_3138 (O_3138,N_28642,N_24025);
nor UO_3139 (O_3139,N_27181,N_25827);
xnor UO_3140 (O_3140,N_29211,N_28767);
nand UO_3141 (O_3141,N_25488,N_29244);
xor UO_3142 (O_3142,N_24592,N_26136);
nand UO_3143 (O_3143,N_28032,N_29497);
or UO_3144 (O_3144,N_27961,N_24549);
xor UO_3145 (O_3145,N_27331,N_26221);
and UO_3146 (O_3146,N_26361,N_27063);
xor UO_3147 (O_3147,N_27286,N_24712);
xor UO_3148 (O_3148,N_24260,N_27081);
nand UO_3149 (O_3149,N_24923,N_24959);
nor UO_3150 (O_3150,N_27912,N_28412);
nor UO_3151 (O_3151,N_29685,N_24427);
xnor UO_3152 (O_3152,N_24073,N_28322);
and UO_3153 (O_3153,N_27596,N_26302);
and UO_3154 (O_3154,N_25521,N_25958);
and UO_3155 (O_3155,N_26669,N_26291);
or UO_3156 (O_3156,N_26068,N_24171);
and UO_3157 (O_3157,N_25304,N_27879);
or UO_3158 (O_3158,N_28294,N_25909);
and UO_3159 (O_3159,N_26955,N_24676);
nor UO_3160 (O_3160,N_27117,N_25238);
nor UO_3161 (O_3161,N_26318,N_24895);
nand UO_3162 (O_3162,N_28609,N_28879);
and UO_3163 (O_3163,N_27569,N_29642);
nor UO_3164 (O_3164,N_24759,N_27803);
xnor UO_3165 (O_3165,N_27926,N_27369);
xor UO_3166 (O_3166,N_28865,N_27364);
xor UO_3167 (O_3167,N_29803,N_27192);
nand UO_3168 (O_3168,N_26583,N_26597);
and UO_3169 (O_3169,N_29752,N_28966);
nor UO_3170 (O_3170,N_29305,N_25015);
xnor UO_3171 (O_3171,N_24506,N_29198);
nor UO_3172 (O_3172,N_27737,N_25490);
xor UO_3173 (O_3173,N_25496,N_27477);
or UO_3174 (O_3174,N_24601,N_28939);
or UO_3175 (O_3175,N_24336,N_29313);
or UO_3176 (O_3176,N_25969,N_27562);
xnor UO_3177 (O_3177,N_27593,N_26598);
xnor UO_3178 (O_3178,N_28839,N_24245);
and UO_3179 (O_3179,N_29251,N_24852);
nor UO_3180 (O_3180,N_29536,N_29744);
nor UO_3181 (O_3181,N_24530,N_28837);
and UO_3182 (O_3182,N_25984,N_26012);
nand UO_3183 (O_3183,N_24859,N_28755);
nand UO_3184 (O_3184,N_28253,N_24099);
xor UO_3185 (O_3185,N_29100,N_24092);
nor UO_3186 (O_3186,N_26138,N_27438);
nor UO_3187 (O_3187,N_27801,N_24699);
xnor UO_3188 (O_3188,N_25414,N_27069);
or UO_3189 (O_3189,N_27197,N_29912);
and UO_3190 (O_3190,N_24713,N_29302);
and UO_3191 (O_3191,N_28714,N_26927);
or UO_3192 (O_3192,N_26880,N_27657);
and UO_3193 (O_3193,N_27554,N_25216);
nand UO_3194 (O_3194,N_27518,N_24344);
xor UO_3195 (O_3195,N_24490,N_27290);
and UO_3196 (O_3196,N_26120,N_25771);
xor UO_3197 (O_3197,N_27914,N_27518);
nand UO_3198 (O_3198,N_26948,N_25217);
or UO_3199 (O_3199,N_29100,N_29847);
xnor UO_3200 (O_3200,N_24355,N_27546);
nor UO_3201 (O_3201,N_26783,N_28033);
nand UO_3202 (O_3202,N_29233,N_24355);
or UO_3203 (O_3203,N_25940,N_26083);
nor UO_3204 (O_3204,N_29351,N_28498);
nand UO_3205 (O_3205,N_24397,N_24430);
nand UO_3206 (O_3206,N_25305,N_26872);
and UO_3207 (O_3207,N_24315,N_29475);
nor UO_3208 (O_3208,N_24570,N_29406);
and UO_3209 (O_3209,N_28214,N_24362);
nor UO_3210 (O_3210,N_27903,N_28534);
nor UO_3211 (O_3211,N_25793,N_25123);
or UO_3212 (O_3212,N_26728,N_27763);
and UO_3213 (O_3213,N_29929,N_24995);
or UO_3214 (O_3214,N_24635,N_28020);
and UO_3215 (O_3215,N_24762,N_29319);
xnor UO_3216 (O_3216,N_25774,N_29223);
nor UO_3217 (O_3217,N_25034,N_27335);
and UO_3218 (O_3218,N_28363,N_28628);
xor UO_3219 (O_3219,N_25125,N_24275);
nor UO_3220 (O_3220,N_26588,N_27679);
nand UO_3221 (O_3221,N_26374,N_28280);
nand UO_3222 (O_3222,N_29619,N_26668);
xnor UO_3223 (O_3223,N_26807,N_28551);
or UO_3224 (O_3224,N_26194,N_27347);
nor UO_3225 (O_3225,N_29673,N_29177);
nor UO_3226 (O_3226,N_28483,N_24983);
or UO_3227 (O_3227,N_24692,N_24529);
xnor UO_3228 (O_3228,N_27317,N_27179);
and UO_3229 (O_3229,N_24926,N_28177);
nor UO_3230 (O_3230,N_24292,N_28598);
nand UO_3231 (O_3231,N_28481,N_24837);
nand UO_3232 (O_3232,N_24766,N_26795);
nand UO_3233 (O_3233,N_28347,N_27661);
or UO_3234 (O_3234,N_28259,N_24626);
or UO_3235 (O_3235,N_29230,N_26571);
nor UO_3236 (O_3236,N_27723,N_25248);
nand UO_3237 (O_3237,N_24778,N_27107);
xnor UO_3238 (O_3238,N_29139,N_25775);
nand UO_3239 (O_3239,N_28678,N_28035);
or UO_3240 (O_3240,N_25179,N_28792);
nand UO_3241 (O_3241,N_29837,N_25612);
or UO_3242 (O_3242,N_24225,N_29001);
and UO_3243 (O_3243,N_27581,N_28012);
or UO_3244 (O_3244,N_28062,N_28057);
nand UO_3245 (O_3245,N_29781,N_25580);
nand UO_3246 (O_3246,N_28252,N_24664);
nand UO_3247 (O_3247,N_27763,N_29383);
or UO_3248 (O_3248,N_27070,N_28167);
nor UO_3249 (O_3249,N_29198,N_29652);
xnor UO_3250 (O_3250,N_24739,N_29087);
nor UO_3251 (O_3251,N_25936,N_29943);
or UO_3252 (O_3252,N_26653,N_29717);
and UO_3253 (O_3253,N_27356,N_26280);
or UO_3254 (O_3254,N_25725,N_29956);
xor UO_3255 (O_3255,N_29408,N_28969);
xnor UO_3256 (O_3256,N_29407,N_25046);
or UO_3257 (O_3257,N_25832,N_24781);
or UO_3258 (O_3258,N_26798,N_28466);
nand UO_3259 (O_3259,N_24541,N_25844);
nor UO_3260 (O_3260,N_25620,N_27837);
xor UO_3261 (O_3261,N_29598,N_26095);
nand UO_3262 (O_3262,N_24396,N_28388);
xor UO_3263 (O_3263,N_27256,N_24042);
nand UO_3264 (O_3264,N_24131,N_28150);
or UO_3265 (O_3265,N_28859,N_24551);
nand UO_3266 (O_3266,N_28688,N_26710);
xor UO_3267 (O_3267,N_26672,N_24071);
and UO_3268 (O_3268,N_28629,N_28547);
nand UO_3269 (O_3269,N_26676,N_28596);
and UO_3270 (O_3270,N_26026,N_28903);
or UO_3271 (O_3271,N_29029,N_29746);
nand UO_3272 (O_3272,N_27374,N_25202);
and UO_3273 (O_3273,N_28470,N_24236);
nand UO_3274 (O_3274,N_27998,N_29988);
or UO_3275 (O_3275,N_26088,N_24876);
nor UO_3276 (O_3276,N_27548,N_29180);
or UO_3277 (O_3277,N_26889,N_24671);
or UO_3278 (O_3278,N_25163,N_28503);
and UO_3279 (O_3279,N_26995,N_27115);
or UO_3280 (O_3280,N_24361,N_27713);
or UO_3281 (O_3281,N_25071,N_28820);
nor UO_3282 (O_3282,N_29047,N_29441);
and UO_3283 (O_3283,N_28585,N_25237);
nand UO_3284 (O_3284,N_27490,N_29353);
nand UO_3285 (O_3285,N_28722,N_29276);
xor UO_3286 (O_3286,N_27789,N_24732);
nand UO_3287 (O_3287,N_27577,N_29119);
xor UO_3288 (O_3288,N_24603,N_26882);
or UO_3289 (O_3289,N_25138,N_25021);
nor UO_3290 (O_3290,N_27470,N_29791);
and UO_3291 (O_3291,N_24057,N_24695);
xnor UO_3292 (O_3292,N_24875,N_25117);
or UO_3293 (O_3293,N_26084,N_24633);
and UO_3294 (O_3294,N_26623,N_24141);
nor UO_3295 (O_3295,N_29934,N_26712);
or UO_3296 (O_3296,N_29887,N_29542);
or UO_3297 (O_3297,N_26968,N_24665);
nand UO_3298 (O_3298,N_29354,N_24739);
or UO_3299 (O_3299,N_28847,N_29195);
nor UO_3300 (O_3300,N_26513,N_27343);
xnor UO_3301 (O_3301,N_28727,N_25400);
or UO_3302 (O_3302,N_25746,N_27621);
nand UO_3303 (O_3303,N_24657,N_28742);
nand UO_3304 (O_3304,N_24010,N_28393);
or UO_3305 (O_3305,N_26640,N_29167);
xor UO_3306 (O_3306,N_27043,N_24169);
nand UO_3307 (O_3307,N_25375,N_28248);
xor UO_3308 (O_3308,N_25618,N_25016);
nor UO_3309 (O_3309,N_29877,N_29984);
xor UO_3310 (O_3310,N_28560,N_26221);
and UO_3311 (O_3311,N_25193,N_26288);
or UO_3312 (O_3312,N_25546,N_25254);
nand UO_3313 (O_3313,N_28622,N_26811);
xor UO_3314 (O_3314,N_24380,N_26139);
and UO_3315 (O_3315,N_27952,N_26297);
nor UO_3316 (O_3316,N_25450,N_27074);
nand UO_3317 (O_3317,N_26703,N_28596);
xor UO_3318 (O_3318,N_28115,N_27864);
xor UO_3319 (O_3319,N_27017,N_29231);
nand UO_3320 (O_3320,N_28676,N_28281);
nand UO_3321 (O_3321,N_28432,N_26015);
nor UO_3322 (O_3322,N_26760,N_29357);
or UO_3323 (O_3323,N_27522,N_25620);
xnor UO_3324 (O_3324,N_27929,N_26038);
and UO_3325 (O_3325,N_24151,N_28733);
and UO_3326 (O_3326,N_28911,N_29385);
xnor UO_3327 (O_3327,N_27146,N_28081);
nand UO_3328 (O_3328,N_27289,N_28647);
nor UO_3329 (O_3329,N_24927,N_29762);
xnor UO_3330 (O_3330,N_29309,N_25917);
xnor UO_3331 (O_3331,N_25180,N_25686);
nor UO_3332 (O_3332,N_25841,N_24708);
or UO_3333 (O_3333,N_25311,N_29127);
or UO_3334 (O_3334,N_29513,N_27550);
and UO_3335 (O_3335,N_26731,N_27469);
and UO_3336 (O_3336,N_27753,N_28940);
or UO_3337 (O_3337,N_26856,N_28756);
nand UO_3338 (O_3338,N_27312,N_24349);
xnor UO_3339 (O_3339,N_24289,N_28434);
nor UO_3340 (O_3340,N_27342,N_28257);
or UO_3341 (O_3341,N_26736,N_29363);
or UO_3342 (O_3342,N_29481,N_28574);
or UO_3343 (O_3343,N_24724,N_28102);
nand UO_3344 (O_3344,N_27279,N_26275);
or UO_3345 (O_3345,N_27709,N_28368);
xnor UO_3346 (O_3346,N_28504,N_24044);
xor UO_3347 (O_3347,N_27489,N_24546);
xor UO_3348 (O_3348,N_24897,N_25278);
nor UO_3349 (O_3349,N_29071,N_27313);
or UO_3350 (O_3350,N_29936,N_28283);
nor UO_3351 (O_3351,N_24528,N_24987);
xnor UO_3352 (O_3352,N_26834,N_26276);
or UO_3353 (O_3353,N_29726,N_27973);
nand UO_3354 (O_3354,N_24995,N_26274);
nor UO_3355 (O_3355,N_28939,N_24267);
nor UO_3356 (O_3356,N_27752,N_28476);
xnor UO_3357 (O_3357,N_28089,N_26506);
or UO_3358 (O_3358,N_27629,N_28210);
and UO_3359 (O_3359,N_26524,N_28147);
xnor UO_3360 (O_3360,N_27664,N_29010);
xnor UO_3361 (O_3361,N_25285,N_26362);
nor UO_3362 (O_3362,N_29024,N_24174);
xor UO_3363 (O_3363,N_26634,N_24581);
or UO_3364 (O_3364,N_27384,N_29465);
nor UO_3365 (O_3365,N_25649,N_26363);
nor UO_3366 (O_3366,N_24548,N_25595);
xnor UO_3367 (O_3367,N_29437,N_27943);
and UO_3368 (O_3368,N_26845,N_24980);
nor UO_3369 (O_3369,N_27169,N_28284);
nand UO_3370 (O_3370,N_29609,N_27987);
xnor UO_3371 (O_3371,N_24047,N_27200);
and UO_3372 (O_3372,N_27791,N_26983);
nand UO_3373 (O_3373,N_24421,N_28428);
xnor UO_3374 (O_3374,N_27394,N_28830);
xnor UO_3375 (O_3375,N_26625,N_27292);
nand UO_3376 (O_3376,N_27531,N_24512);
and UO_3377 (O_3377,N_26177,N_25508);
or UO_3378 (O_3378,N_25400,N_25652);
and UO_3379 (O_3379,N_27412,N_29241);
nor UO_3380 (O_3380,N_25787,N_24587);
nor UO_3381 (O_3381,N_24020,N_29711);
nor UO_3382 (O_3382,N_29034,N_27470);
and UO_3383 (O_3383,N_25723,N_28625);
or UO_3384 (O_3384,N_26214,N_26047);
nor UO_3385 (O_3385,N_24626,N_25262);
nor UO_3386 (O_3386,N_24048,N_25603);
nor UO_3387 (O_3387,N_25988,N_25785);
or UO_3388 (O_3388,N_24112,N_28983);
nand UO_3389 (O_3389,N_25971,N_29955);
xor UO_3390 (O_3390,N_29314,N_27795);
nor UO_3391 (O_3391,N_24767,N_25835);
and UO_3392 (O_3392,N_26098,N_29398);
and UO_3393 (O_3393,N_29580,N_26030);
nor UO_3394 (O_3394,N_29941,N_28814);
nand UO_3395 (O_3395,N_24007,N_24324);
and UO_3396 (O_3396,N_29210,N_27492);
and UO_3397 (O_3397,N_27076,N_28839);
and UO_3398 (O_3398,N_27511,N_27803);
xor UO_3399 (O_3399,N_28506,N_29060);
nand UO_3400 (O_3400,N_28355,N_26570);
nor UO_3401 (O_3401,N_28199,N_27644);
nand UO_3402 (O_3402,N_29329,N_24138);
xnor UO_3403 (O_3403,N_24583,N_27253);
xnor UO_3404 (O_3404,N_26447,N_28391);
or UO_3405 (O_3405,N_25217,N_29321);
nor UO_3406 (O_3406,N_28019,N_27861);
and UO_3407 (O_3407,N_24767,N_28349);
xnor UO_3408 (O_3408,N_29540,N_24623);
nor UO_3409 (O_3409,N_26569,N_24527);
and UO_3410 (O_3410,N_29709,N_26356);
xnor UO_3411 (O_3411,N_26795,N_25145);
nand UO_3412 (O_3412,N_25420,N_28761);
and UO_3413 (O_3413,N_24842,N_29391);
nand UO_3414 (O_3414,N_25461,N_25327);
and UO_3415 (O_3415,N_25320,N_27712);
and UO_3416 (O_3416,N_26692,N_29517);
nor UO_3417 (O_3417,N_26967,N_28355);
or UO_3418 (O_3418,N_27920,N_26589);
and UO_3419 (O_3419,N_25908,N_26743);
xor UO_3420 (O_3420,N_28305,N_25895);
xnor UO_3421 (O_3421,N_26358,N_29579);
nor UO_3422 (O_3422,N_28931,N_29712);
or UO_3423 (O_3423,N_28752,N_26668);
and UO_3424 (O_3424,N_27438,N_28062);
nor UO_3425 (O_3425,N_25575,N_28559);
or UO_3426 (O_3426,N_29105,N_24815);
and UO_3427 (O_3427,N_26395,N_27675);
nor UO_3428 (O_3428,N_29075,N_26956);
nor UO_3429 (O_3429,N_29252,N_27558);
or UO_3430 (O_3430,N_27034,N_24757);
nor UO_3431 (O_3431,N_28189,N_28651);
and UO_3432 (O_3432,N_25333,N_25753);
or UO_3433 (O_3433,N_24603,N_28642);
xor UO_3434 (O_3434,N_27823,N_27470);
xnor UO_3435 (O_3435,N_24246,N_27793);
or UO_3436 (O_3436,N_24300,N_26031);
xnor UO_3437 (O_3437,N_24946,N_26625);
or UO_3438 (O_3438,N_27069,N_29246);
and UO_3439 (O_3439,N_28204,N_26393);
and UO_3440 (O_3440,N_24215,N_29536);
nand UO_3441 (O_3441,N_27481,N_28951);
nor UO_3442 (O_3442,N_26662,N_27501);
nand UO_3443 (O_3443,N_29162,N_29388);
xnor UO_3444 (O_3444,N_29345,N_24581);
nor UO_3445 (O_3445,N_29718,N_26096);
or UO_3446 (O_3446,N_29376,N_24421);
nor UO_3447 (O_3447,N_24472,N_26155);
and UO_3448 (O_3448,N_27802,N_24035);
nand UO_3449 (O_3449,N_29197,N_25695);
and UO_3450 (O_3450,N_25913,N_28085);
and UO_3451 (O_3451,N_24751,N_26748);
xnor UO_3452 (O_3452,N_28681,N_27674);
xnor UO_3453 (O_3453,N_28609,N_28529);
nor UO_3454 (O_3454,N_27457,N_26618);
nand UO_3455 (O_3455,N_26405,N_28156);
nand UO_3456 (O_3456,N_26516,N_26602);
nand UO_3457 (O_3457,N_26150,N_24793);
xnor UO_3458 (O_3458,N_24470,N_27413);
and UO_3459 (O_3459,N_29988,N_29033);
xnor UO_3460 (O_3460,N_25338,N_25747);
nor UO_3461 (O_3461,N_26283,N_26944);
and UO_3462 (O_3462,N_27180,N_25968);
nand UO_3463 (O_3463,N_28569,N_27946);
and UO_3464 (O_3464,N_24874,N_28200);
nand UO_3465 (O_3465,N_25896,N_27452);
xnor UO_3466 (O_3466,N_26024,N_27135);
nand UO_3467 (O_3467,N_27144,N_28716);
xor UO_3468 (O_3468,N_29420,N_29895);
nand UO_3469 (O_3469,N_26190,N_26624);
or UO_3470 (O_3470,N_28458,N_28432);
nor UO_3471 (O_3471,N_24992,N_26843);
nand UO_3472 (O_3472,N_26848,N_28189);
xor UO_3473 (O_3473,N_26862,N_25992);
xnor UO_3474 (O_3474,N_25676,N_29635);
nand UO_3475 (O_3475,N_29705,N_27383);
nor UO_3476 (O_3476,N_29395,N_26680);
and UO_3477 (O_3477,N_24615,N_24963);
or UO_3478 (O_3478,N_24754,N_28471);
nor UO_3479 (O_3479,N_24039,N_25666);
nand UO_3480 (O_3480,N_27318,N_24550);
xor UO_3481 (O_3481,N_25495,N_25765);
and UO_3482 (O_3482,N_28053,N_27403);
xnor UO_3483 (O_3483,N_24416,N_28738);
nor UO_3484 (O_3484,N_28266,N_27541);
and UO_3485 (O_3485,N_25623,N_28807);
nor UO_3486 (O_3486,N_27508,N_29900);
xor UO_3487 (O_3487,N_29122,N_26272);
nand UO_3488 (O_3488,N_25112,N_27891);
or UO_3489 (O_3489,N_26086,N_27696);
nor UO_3490 (O_3490,N_24679,N_29445);
nand UO_3491 (O_3491,N_29306,N_29720);
and UO_3492 (O_3492,N_29256,N_29499);
xnor UO_3493 (O_3493,N_29840,N_28687);
or UO_3494 (O_3494,N_24430,N_24964);
nor UO_3495 (O_3495,N_27618,N_25274);
or UO_3496 (O_3496,N_25991,N_25872);
nor UO_3497 (O_3497,N_29038,N_29110);
and UO_3498 (O_3498,N_29094,N_29386);
or UO_3499 (O_3499,N_28187,N_29752);
endmodule