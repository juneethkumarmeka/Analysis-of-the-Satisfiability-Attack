module basic_750_5000_1000_5_levels_10xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
and U0 (N_0,In_364,In_204);
nor U1 (N_1,In_403,In_327);
nand U2 (N_2,In_519,In_647);
nor U3 (N_3,In_676,In_578);
xnor U4 (N_4,In_379,In_474);
and U5 (N_5,In_714,In_342);
or U6 (N_6,In_84,In_555);
xnor U7 (N_7,In_596,In_92);
xnor U8 (N_8,In_457,In_160);
and U9 (N_9,In_566,In_175);
nor U10 (N_10,In_642,In_462);
nor U11 (N_11,In_664,In_299);
and U12 (N_12,In_627,In_203);
nor U13 (N_13,In_202,In_608);
nand U14 (N_14,In_214,In_530);
nor U15 (N_15,In_586,In_51);
or U16 (N_16,In_521,In_53);
xnor U17 (N_17,In_66,In_245);
xor U18 (N_18,In_70,In_511);
nand U19 (N_19,In_649,In_675);
nand U20 (N_20,In_226,In_551);
xor U21 (N_21,In_308,In_372);
nor U22 (N_22,In_728,In_142);
and U23 (N_23,In_77,In_37);
xor U24 (N_24,In_346,In_445);
xnor U25 (N_25,In_493,In_437);
nor U26 (N_26,In_148,In_580);
nor U27 (N_27,In_562,In_145);
xnor U28 (N_28,In_234,In_362);
xnor U29 (N_29,In_112,In_141);
xor U30 (N_30,In_638,In_701);
nor U31 (N_31,In_380,In_679);
or U32 (N_32,In_72,In_516);
nand U33 (N_33,In_262,In_13);
xnor U34 (N_34,In_236,In_723);
and U35 (N_35,In_206,In_375);
nor U36 (N_36,In_539,In_450);
xnor U37 (N_37,In_123,In_549);
and U38 (N_38,In_400,In_653);
nand U39 (N_39,In_528,In_600);
and U40 (N_40,In_146,In_44);
nor U41 (N_41,In_573,In_703);
and U42 (N_42,In_67,In_257);
and U43 (N_43,In_100,In_295);
or U44 (N_44,In_483,In_274);
or U45 (N_45,In_698,In_629);
nand U46 (N_46,In_315,In_136);
xor U47 (N_47,In_46,In_189);
or U48 (N_48,In_561,In_536);
nand U49 (N_49,In_416,In_275);
xor U50 (N_50,In_106,In_127);
or U51 (N_51,In_184,In_113);
xor U52 (N_52,In_232,In_572);
nor U53 (N_53,In_176,In_691);
nand U54 (N_54,In_48,In_405);
and U55 (N_55,In_495,In_122);
xor U56 (N_56,In_294,In_690);
nor U57 (N_57,In_65,In_111);
xnor U58 (N_58,In_465,In_417);
or U59 (N_59,In_497,In_150);
or U60 (N_60,In_569,In_431);
xor U61 (N_61,In_440,In_481);
nand U62 (N_62,In_25,In_291);
or U63 (N_63,In_620,In_435);
nand U64 (N_64,In_674,In_27);
xor U65 (N_65,In_745,In_339);
nor U66 (N_66,In_643,In_548);
nand U67 (N_67,In_482,In_449);
and U68 (N_68,In_470,In_397);
nor U69 (N_69,In_218,In_60);
nand U70 (N_70,In_606,In_692);
xnor U71 (N_71,In_35,In_689);
nand U72 (N_72,In_338,In_744);
or U73 (N_73,In_311,In_360);
nor U74 (N_74,In_278,In_87);
xor U75 (N_75,In_314,In_162);
nor U76 (N_76,In_115,In_731);
xnor U77 (N_77,In_505,In_394);
or U78 (N_78,In_300,In_699);
and U79 (N_79,In_742,In_211);
or U80 (N_80,In_590,In_533);
or U81 (N_81,In_614,In_373);
and U82 (N_82,In_165,In_544);
xor U83 (N_83,In_334,In_96);
or U84 (N_84,In_740,In_584);
and U85 (N_85,In_448,In_737);
or U86 (N_86,In_290,In_0);
and U87 (N_87,In_266,In_149);
nor U88 (N_88,In_560,In_556);
or U89 (N_89,In_355,In_532);
nand U90 (N_90,In_240,In_542);
xor U91 (N_91,In_14,In_237);
and U92 (N_92,In_452,In_718);
and U93 (N_93,In_194,In_395);
nor U94 (N_94,In_504,In_531);
nor U95 (N_95,In_345,In_658);
nor U96 (N_96,In_711,In_282);
nor U97 (N_97,In_7,In_591);
and U98 (N_98,In_478,In_101);
xor U99 (N_99,In_683,In_665);
or U100 (N_100,In_292,In_579);
or U101 (N_101,In_348,In_632);
nand U102 (N_102,In_49,In_201);
and U103 (N_103,In_337,In_69);
and U104 (N_104,In_215,In_678);
nor U105 (N_105,In_329,In_59);
nand U106 (N_106,In_577,In_509);
nor U107 (N_107,In_438,In_270);
nand U108 (N_108,In_9,In_29);
nand U109 (N_109,In_408,In_30);
nor U110 (N_110,In_11,In_631);
or U111 (N_111,In_120,In_534);
or U112 (N_112,In_351,In_568);
or U113 (N_113,In_419,In_81);
xor U114 (N_114,In_306,In_684);
nor U115 (N_115,In_258,In_210);
nor U116 (N_116,In_52,In_253);
nor U117 (N_117,In_143,In_62);
and U118 (N_118,In_110,In_139);
nor U119 (N_119,In_15,In_363);
nor U120 (N_120,In_97,In_490);
nand U121 (N_121,In_507,In_114);
xnor U122 (N_122,In_147,In_229);
nand U123 (N_123,In_54,In_444);
nand U124 (N_124,In_433,In_494);
nand U125 (N_125,In_209,In_280);
nand U126 (N_126,In_641,In_358);
and U127 (N_127,In_2,In_715);
nand U128 (N_128,In_354,In_694);
nand U129 (N_129,In_721,In_571);
nand U130 (N_130,In_704,In_89);
xor U131 (N_131,In_17,In_567);
nor U132 (N_132,In_654,In_19);
and U133 (N_133,In_63,In_377);
xor U134 (N_134,In_242,In_366);
nor U135 (N_135,In_381,In_276);
or U136 (N_136,In_50,In_697);
xor U137 (N_137,In_598,In_456);
nand U138 (N_138,In_124,In_3);
xor U139 (N_139,In_134,In_264);
nand U140 (N_140,In_344,In_503);
nor U141 (N_141,In_657,In_422);
xor U142 (N_142,In_79,In_582);
or U143 (N_143,In_22,In_707);
xor U144 (N_144,In_669,In_479);
xnor U145 (N_145,In_559,In_386);
xor U146 (N_146,In_732,In_547);
nand U147 (N_147,In_498,In_621);
xor U148 (N_148,In_263,In_168);
nor U149 (N_149,In_126,In_180);
nand U150 (N_150,In_563,In_57);
nand U151 (N_151,In_188,In_623);
nor U152 (N_152,In_451,In_152);
nand U153 (N_153,In_365,In_702);
xor U154 (N_154,In_288,In_182);
or U155 (N_155,In_390,In_217);
nor U156 (N_156,In_537,In_499);
nor U157 (N_157,In_619,In_475);
nor U158 (N_158,In_332,In_33);
and U159 (N_159,In_39,In_31);
or U160 (N_160,In_522,In_36);
xnor U161 (N_161,In_595,In_520);
xor U162 (N_162,In_648,In_628);
and U163 (N_163,In_615,In_538);
nand U164 (N_164,In_318,In_196);
or U165 (N_165,In_325,In_179);
or U166 (N_166,In_45,In_349);
xor U167 (N_167,In_304,In_73);
xnor U168 (N_168,In_157,In_441);
xnor U169 (N_169,In_645,In_575);
nand U170 (N_170,In_398,In_513);
and U171 (N_171,In_335,In_713);
nand U172 (N_172,In_399,In_213);
nor U173 (N_173,In_487,In_42);
or U174 (N_174,In_489,In_421);
xor U175 (N_175,In_91,In_251);
xor U176 (N_176,In_524,In_594);
or U177 (N_177,In_454,In_726);
nor U178 (N_178,In_671,In_535);
nand U179 (N_179,In_401,In_167);
and U180 (N_180,In_130,In_265);
or U181 (N_181,In_733,In_480);
nand U182 (N_182,In_191,In_287);
and U183 (N_183,In_552,In_652);
nor U184 (N_184,In_64,In_221);
or U185 (N_185,In_310,In_387);
nor U186 (N_186,In_635,In_739);
and U187 (N_187,In_404,In_166);
xnor U188 (N_188,In_8,In_611);
xor U189 (N_189,In_720,In_748);
or U190 (N_190,In_252,In_28);
nor U191 (N_191,In_576,In_249);
nand U192 (N_192,In_68,In_170);
or U193 (N_193,In_383,In_333);
xnor U194 (N_194,In_693,In_687);
and U195 (N_195,In_612,In_467);
and U196 (N_196,In_370,In_646);
nand U197 (N_197,In_105,In_564);
nand U198 (N_198,In_281,In_78);
nor U199 (N_199,In_117,In_662);
nand U200 (N_200,In_95,In_430);
nand U201 (N_201,In_722,In_393);
nor U202 (N_202,In_486,In_650);
or U203 (N_203,In_322,In_453);
nand U204 (N_204,In_410,In_545);
and U205 (N_205,In_540,In_5);
and U206 (N_206,In_216,In_369);
and U207 (N_207,In_601,In_427);
xnor U208 (N_208,In_350,In_384);
or U209 (N_209,In_446,In_668);
and U210 (N_210,In_301,In_197);
and U211 (N_211,In_599,In_121);
nand U212 (N_212,In_321,In_463);
or U213 (N_213,In_227,In_298);
nand U214 (N_214,In_220,In_198);
nand U215 (N_215,In_436,In_90);
xor U216 (N_216,In_340,In_554);
nor U217 (N_217,In_378,In_432);
nand U218 (N_218,In_407,In_207);
xor U219 (N_219,In_492,In_447);
or U220 (N_220,In_376,In_330);
nand U221 (N_221,In_735,In_6);
or U222 (N_222,In_367,In_98);
nor U223 (N_223,In_686,In_34);
nand U224 (N_224,In_391,In_94);
or U225 (N_225,In_464,In_624);
and U226 (N_226,In_233,In_592);
xnor U227 (N_227,In_38,In_75);
and U228 (N_228,In_514,In_472);
nand U229 (N_229,In_622,In_501);
nand U230 (N_230,In_734,In_268);
or U231 (N_231,In_685,In_651);
nand U232 (N_232,In_230,In_389);
xor U233 (N_233,In_4,In_717);
and U234 (N_234,In_666,In_151);
and U235 (N_235,In_428,In_71);
xnor U236 (N_236,In_86,In_107);
nand U237 (N_237,In_730,In_104);
nor U238 (N_238,In_56,In_640);
nor U239 (N_239,In_102,In_284);
nor U240 (N_240,In_593,In_637);
and U241 (N_241,In_589,In_279);
or U242 (N_242,In_382,In_272);
nand U243 (N_243,In_239,In_618);
and U244 (N_244,In_336,In_710);
xor U245 (N_245,In_546,In_357);
nand U246 (N_246,In_396,In_736);
nand U247 (N_247,In_323,In_565);
nand U248 (N_248,In_305,In_604);
xnor U249 (N_249,In_241,In_250);
nand U250 (N_250,In_40,In_244);
xnor U251 (N_251,In_247,In_103);
or U252 (N_252,In_413,In_461);
xor U253 (N_253,In_80,In_231);
nor U254 (N_254,In_585,In_420);
and U255 (N_255,In_273,In_177);
nand U256 (N_256,In_385,In_696);
xnor U257 (N_257,In_660,In_353);
nand U258 (N_258,In_429,In_708);
xnor U259 (N_259,In_469,In_259);
nand U260 (N_260,In_442,In_267);
nor U261 (N_261,In_512,In_208);
or U262 (N_262,In_137,In_125);
xor U263 (N_263,In_169,In_688);
nand U264 (N_264,In_316,In_248);
nand U265 (N_265,In_418,In_525);
or U266 (N_266,In_317,In_634);
nand U267 (N_267,In_517,In_153);
and U268 (N_268,In_476,In_293);
and U269 (N_269,In_307,In_529);
xor U270 (N_270,In_138,In_673);
and U271 (N_271,In_729,In_558);
and U272 (N_272,In_439,In_131);
nor U273 (N_273,In_200,In_523);
nor U274 (N_274,In_326,In_541);
nand U275 (N_275,In_23,In_61);
nor U276 (N_276,In_343,In_706);
and U277 (N_277,In_625,In_426);
and U278 (N_278,In_361,In_719);
xor U279 (N_279,In_24,In_459);
or U280 (N_280,In_260,In_163);
xor U281 (N_281,In_617,In_1);
nand U282 (N_282,In_144,In_741);
nand U283 (N_283,In_331,In_109);
nor U284 (N_284,In_171,In_434);
nand U285 (N_285,In_412,In_709);
xnor U286 (N_286,In_93,In_246);
or U287 (N_287,In_313,In_656);
and U288 (N_288,In_550,In_425);
and U289 (N_289,In_12,In_374);
nand U290 (N_290,In_255,In_302);
nand U291 (N_291,In_749,In_553);
nand U292 (N_292,In_727,In_271);
and U293 (N_293,In_466,In_83);
and U294 (N_294,In_473,In_661);
and U295 (N_295,In_18,In_414);
nor U296 (N_296,In_411,In_88);
and U297 (N_297,In_402,In_655);
or U298 (N_298,In_626,In_477);
and U299 (N_299,In_190,In_164);
or U300 (N_300,In_156,In_603);
or U301 (N_301,In_223,In_609);
nor U302 (N_302,In_471,In_256);
and U303 (N_303,In_633,In_43);
or U304 (N_304,In_341,In_173);
nand U305 (N_305,In_518,In_677);
xnor U306 (N_306,In_725,In_506);
nor U307 (N_307,In_133,In_468);
nor U308 (N_308,In_680,In_128);
and U309 (N_309,In_607,In_132);
xnor U310 (N_310,In_458,In_455);
and U311 (N_311,In_140,In_672);
or U312 (N_312,In_597,In_154);
nor U313 (N_313,In_10,In_118);
or U314 (N_314,In_527,In_219);
or U315 (N_315,In_283,In_222);
or U316 (N_316,In_639,In_289);
nand U317 (N_317,In_574,In_570);
xnor U318 (N_318,In_724,In_199);
nor U319 (N_319,In_174,In_235);
or U320 (N_320,In_347,In_583);
nand U321 (N_321,In_616,In_116);
nand U322 (N_322,In_712,In_630);
xor U323 (N_323,In_488,In_423);
nand U324 (N_324,In_41,In_21);
nor U325 (N_325,In_158,In_667);
nor U326 (N_326,In_663,In_324);
nand U327 (N_327,In_187,In_286);
nand U328 (N_328,In_277,In_183);
xnor U329 (N_329,In_443,In_543);
xor U330 (N_330,In_178,In_320);
and U331 (N_331,In_682,In_496);
nand U332 (N_332,In_285,In_581);
or U333 (N_333,In_356,In_20);
xnor U334 (N_334,In_502,In_681);
nor U335 (N_335,In_224,In_135);
nand U336 (N_336,In_636,In_238);
nor U337 (N_337,In_243,In_508);
nand U338 (N_338,In_491,In_352);
xnor U339 (N_339,In_82,In_32);
or U340 (N_340,In_228,In_181);
or U341 (N_341,In_716,In_700);
xor U342 (N_342,In_359,In_644);
nor U343 (N_343,In_500,In_587);
nor U344 (N_344,In_424,In_296);
xor U345 (N_345,In_705,In_74);
or U346 (N_346,In_99,In_371);
xor U347 (N_347,In_388,In_225);
xor U348 (N_348,In_610,In_261);
nand U349 (N_349,In_510,In_738);
nand U350 (N_350,In_26,In_409);
nor U351 (N_351,In_205,In_485);
nand U352 (N_352,In_55,In_319);
or U353 (N_353,In_186,In_695);
xnor U354 (N_354,In_743,In_602);
and U355 (N_355,In_392,In_312);
or U356 (N_356,In_484,In_155);
xnor U357 (N_357,In_159,In_406);
nand U358 (N_358,In_16,In_368);
nor U359 (N_359,In_193,In_515);
xnor U360 (N_360,In_670,In_328);
or U361 (N_361,In_526,In_303);
and U362 (N_362,In_605,In_254);
xnor U363 (N_363,In_557,In_47);
xnor U364 (N_364,In_76,In_58);
nor U365 (N_365,In_613,In_195);
or U366 (N_366,In_192,In_460);
nand U367 (N_367,In_746,In_172);
nor U368 (N_368,In_129,In_185);
and U369 (N_369,In_269,In_212);
xnor U370 (N_370,In_309,In_108);
nor U371 (N_371,In_85,In_161);
nand U372 (N_372,In_297,In_588);
nor U373 (N_373,In_119,In_659);
or U374 (N_374,In_747,In_415);
nand U375 (N_375,In_70,In_141);
xor U376 (N_376,In_258,In_305);
nor U377 (N_377,In_28,In_283);
nor U378 (N_378,In_272,In_260);
or U379 (N_379,In_224,In_740);
nand U380 (N_380,In_62,In_659);
nand U381 (N_381,In_389,In_560);
nor U382 (N_382,In_382,In_232);
and U383 (N_383,In_181,In_506);
or U384 (N_384,In_281,In_438);
xor U385 (N_385,In_604,In_48);
or U386 (N_386,In_230,In_419);
nor U387 (N_387,In_60,In_260);
and U388 (N_388,In_636,In_610);
xnor U389 (N_389,In_150,In_291);
xor U390 (N_390,In_595,In_641);
or U391 (N_391,In_675,In_424);
xor U392 (N_392,In_528,In_677);
xor U393 (N_393,In_230,In_724);
nand U394 (N_394,In_597,In_110);
xor U395 (N_395,In_165,In_677);
nor U396 (N_396,In_695,In_126);
xor U397 (N_397,In_128,In_14);
xor U398 (N_398,In_187,In_533);
nor U399 (N_399,In_86,In_574);
nand U400 (N_400,In_544,In_498);
and U401 (N_401,In_83,In_636);
nand U402 (N_402,In_321,In_329);
nand U403 (N_403,In_287,In_54);
nor U404 (N_404,In_596,In_339);
nor U405 (N_405,In_299,In_366);
nand U406 (N_406,In_537,In_106);
nand U407 (N_407,In_202,In_379);
nor U408 (N_408,In_338,In_652);
and U409 (N_409,In_731,In_352);
nand U410 (N_410,In_258,In_657);
nor U411 (N_411,In_96,In_739);
or U412 (N_412,In_575,In_362);
nor U413 (N_413,In_546,In_399);
nor U414 (N_414,In_688,In_150);
or U415 (N_415,In_120,In_677);
or U416 (N_416,In_496,In_294);
nor U417 (N_417,In_704,In_134);
nand U418 (N_418,In_165,In_685);
xor U419 (N_419,In_180,In_163);
nand U420 (N_420,In_597,In_670);
or U421 (N_421,In_621,In_596);
xnor U422 (N_422,In_700,In_373);
and U423 (N_423,In_276,In_161);
and U424 (N_424,In_335,In_512);
nor U425 (N_425,In_68,In_532);
and U426 (N_426,In_700,In_155);
and U427 (N_427,In_749,In_194);
and U428 (N_428,In_202,In_346);
and U429 (N_429,In_631,In_742);
or U430 (N_430,In_710,In_495);
nor U431 (N_431,In_600,In_512);
or U432 (N_432,In_108,In_431);
nand U433 (N_433,In_563,In_90);
nand U434 (N_434,In_446,In_3);
and U435 (N_435,In_179,In_632);
nor U436 (N_436,In_243,In_412);
xnor U437 (N_437,In_669,In_317);
nand U438 (N_438,In_154,In_412);
nand U439 (N_439,In_605,In_317);
or U440 (N_440,In_152,In_168);
xor U441 (N_441,In_518,In_529);
xnor U442 (N_442,In_513,In_41);
nor U443 (N_443,In_279,In_55);
nor U444 (N_444,In_327,In_401);
nand U445 (N_445,In_580,In_40);
nand U446 (N_446,In_230,In_35);
xor U447 (N_447,In_522,In_561);
nand U448 (N_448,In_581,In_193);
nand U449 (N_449,In_717,In_287);
and U450 (N_450,In_8,In_371);
or U451 (N_451,In_16,In_692);
or U452 (N_452,In_180,In_182);
xor U453 (N_453,In_370,In_207);
and U454 (N_454,In_331,In_278);
or U455 (N_455,In_599,In_618);
nor U456 (N_456,In_122,In_682);
nand U457 (N_457,In_426,In_640);
or U458 (N_458,In_94,In_678);
or U459 (N_459,In_249,In_240);
or U460 (N_460,In_92,In_322);
or U461 (N_461,In_95,In_126);
or U462 (N_462,In_27,In_171);
nand U463 (N_463,In_642,In_603);
xor U464 (N_464,In_369,In_656);
nand U465 (N_465,In_458,In_384);
and U466 (N_466,In_248,In_646);
xnor U467 (N_467,In_379,In_367);
or U468 (N_468,In_692,In_591);
xor U469 (N_469,In_329,In_601);
and U470 (N_470,In_458,In_732);
xnor U471 (N_471,In_243,In_25);
nor U472 (N_472,In_404,In_203);
nand U473 (N_473,In_322,In_1);
nand U474 (N_474,In_692,In_446);
xnor U475 (N_475,In_354,In_62);
nand U476 (N_476,In_675,In_520);
or U477 (N_477,In_502,In_236);
and U478 (N_478,In_301,In_430);
nand U479 (N_479,In_660,In_320);
nand U480 (N_480,In_98,In_159);
xor U481 (N_481,In_64,In_244);
nand U482 (N_482,In_85,In_125);
and U483 (N_483,In_99,In_657);
xor U484 (N_484,In_129,In_476);
nor U485 (N_485,In_316,In_0);
or U486 (N_486,In_101,In_465);
or U487 (N_487,In_66,In_243);
nand U488 (N_488,In_113,In_602);
nand U489 (N_489,In_56,In_744);
nand U490 (N_490,In_475,In_701);
nand U491 (N_491,In_731,In_426);
or U492 (N_492,In_256,In_680);
xnor U493 (N_493,In_625,In_211);
nor U494 (N_494,In_125,In_82);
xor U495 (N_495,In_9,In_423);
xor U496 (N_496,In_222,In_680);
nand U497 (N_497,In_66,In_564);
or U498 (N_498,In_501,In_606);
nor U499 (N_499,In_576,In_422);
and U500 (N_500,In_632,In_521);
and U501 (N_501,In_548,In_30);
xnor U502 (N_502,In_291,In_158);
nand U503 (N_503,In_32,In_292);
nand U504 (N_504,In_680,In_501);
xnor U505 (N_505,In_615,In_139);
nand U506 (N_506,In_435,In_120);
xor U507 (N_507,In_506,In_172);
or U508 (N_508,In_293,In_744);
xor U509 (N_509,In_464,In_730);
xnor U510 (N_510,In_56,In_1);
xnor U511 (N_511,In_112,In_226);
or U512 (N_512,In_104,In_439);
and U513 (N_513,In_154,In_232);
nand U514 (N_514,In_91,In_295);
nand U515 (N_515,In_156,In_568);
and U516 (N_516,In_242,In_363);
and U517 (N_517,In_154,In_580);
nor U518 (N_518,In_673,In_388);
nand U519 (N_519,In_323,In_749);
nor U520 (N_520,In_324,In_420);
and U521 (N_521,In_6,In_408);
and U522 (N_522,In_43,In_391);
nand U523 (N_523,In_84,In_214);
and U524 (N_524,In_678,In_477);
or U525 (N_525,In_91,In_101);
nor U526 (N_526,In_43,In_254);
nand U527 (N_527,In_487,In_529);
xor U528 (N_528,In_536,In_666);
and U529 (N_529,In_692,In_682);
or U530 (N_530,In_276,In_213);
xnor U531 (N_531,In_206,In_268);
nor U532 (N_532,In_682,In_253);
xor U533 (N_533,In_83,In_678);
xnor U534 (N_534,In_180,In_659);
or U535 (N_535,In_698,In_628);
or U536 (N_536,In_430,In_227);
and U537 (N_537,In_25,In_458);
nor U538 (N_538,In_263,In_265);
nor U539 (N_539,In_261,In_81);
or U540 (N_540,In_720,In_231);
xor U541 (N_541,In_686,In_500);
or U542 (N_542,In_104,In_526);
nand U543 (N_543,In_146,In_260);
or U544 (N_544,In_409,In_243);
and U545 (N_545,In_281,In_514);
and U546 (N_546,In_209,In_378);
nor U547 (N_547,In_562,In_590);
and U548 (N_548,In_209,In_59);
or U549 (N_549,In_609,In_291);
or U550 (N_550,In_614,In_702);
nor U551 (N_551,In_480,In_45);
xor U552 (N_552,In_233,In_452);
and U553 (N_553,In_81,In_524);
and U554 (N_554,In_401,In_306);
xnor U555 (N_555,In_539,In_647);
nor U556 (N_556,In_40,In_10);
xor U557 (N_557,In_200,In_412);
nor U558 (N_558,In_109,In_21);
nor U559 (N_559,In_677,In_62);
nand U560 (N_560,In_76,In_550);
xnor U561 (N_561,In_485,In_573);
xnor U562 (N_562,In_301,In_589);
xor U563 (N_563,In_457,In_638);
and U564 (N_564,In_670,In_235);
and U565 (N_565,In_696,In_40);
and U566 (N_566,In_490,In_240);
and U567 (N_567,In_338,In_685);
xnor U568 (N_568,In_700,In_374);
or U569 (N_569,In_689,In_297);
nand U570 (N_570,In_367,In_605);
and U571 (N_571,In_658,In_682);
or U572 (N_572,In_700,In_605);
nand U573 (N_573,In_195,In_503);
xor U574 (N_574,In_282,In_157);
nand U575 (N_575,In_125,In_508);
or U576 (N_576,In_127,In_534);
nor U577 (N_577,In_677,In_157);
nand U578 (N_578,In_723,In_339);
nand U579 (N_579,In_80,In_127);
nor U580 (N_580,In_195,In_389);
nand U581 (N_581,In_70,In_173);
nor U582 (N_582,In_339,In_528);
and U583 (N_583,In_441,In_411);
or U584 (N_584,In_514,In_175);
or U585 (N_585,In_398,In_521);
or U586 (N_586,In_581,In_315);
and U587 (N_587,In_45,In_713);
nor U588 (N_588,In_508,In_416);
and U589 (N_589,In_239,In_517);
xor U590 (N_590,In_336,In_650);
and U591 (N_591,In_183,In_305);
or U592 (N_592,In_355,In_591);
nand U593 (N_593,In_623,In_505);
nor U594 (N_594,In_368,In_471);
and U595 (N_595,In_506,In_555);
or U596 (N_596,In_746,In_485);
nor U597 (N_597,In_280,In_383);
nor U598 (N_598,In_387,In_376);
nand U599 (N_599,In_428,In_594);
and U600 (N_600,In_565,In_594);
nor U601 (N_601,In_164,In_728);
xor U602 (N_602,In_477,In_25);
or U603 (N_603,In_201,In_323);
and U604 (N_604,In_747,In_107);
xnor U605 (N_605,In_325,In_69);
nor U606 (N_606,In_513,In_3);
nand U607 (N_607,In_271,In_707);
nand U608 (N_608,In_313,In_515);
and U609 (N_609,In_489,In_359);
xnor U610 (N_610,In_5,In_711);
nand U611 (N_611,In_110,In_663);
or U612 (N_612,In_736,In_200);
and U613 (N_613,In_400,In_442);
or U614 (N_614,In_96,In_329);
nand U615 (N_615,In_387,In_391);
and U616 (N_616,In_220,In_533);
nor U617 (N_617,In_270,In_741);
xnor U618 (N_618,In_412,In_733);
nor U619 (N_619,In_34,In_6);
and U620 (N_620,In_462,In_128);
or U621 (N_621,In_247,In_0);
or U622 (N_622,In_266,In_242);
and U623 (N_623,In_540,In_314);
or U624 (N_624,In_708,In_579);
or U625 (N_625,In_383,In_340);
and U626 (N_626,In_434,In_622);
nor U627 (N_627,In_318,In_608);
or U628 (N_628,In_309,In_614);
and U629 (N_629,In_368,In_8);
xnor U630 (N_630,In_235,In_426);
nand U631 (N_631,In_592,In_120);
or U632 (N_632,In_312,In_12);
nand U633 (N_633,In_82,In_122);
or U634 (N_634,In_589,In_422);
nand U635 (N_635,In_290,In_562);
xnor U636 (N_636,In_250,In_288);
nand U637 (N_637,In_439,In_149);
or U638 (N_638,In_61,In_458);
nor U639 (N_639,In_288,In_173);
xor U640 (N_640,In_708,In_413);
and U641 (N_641,In_562,In_375);
and U642 (N_642,In_704,In_738);
or U643 (N_643,In_351,In_597);
and U644 (N_644,In_595,In_739);
or U645 (N_645,In_282,In_238);
nand U646 (N_646,In_629,In_111);
or U647 (N_647,In_334,In_685);
xor U648 (N_648,In_359,In_612);
and U649 (N_649,In_199,In_613);
or U650 (N_650,In_667,In_467);
or U651 (N_651,In_678,In_664);
or U652 (N_652,In_211,In_562);
and U653 (N_653,In_483,In_146);
and U654 (N_654,In_576,In_21);
nand U655 (N_655,In_230,In_356);
or U656 (N_656,In_360,In_115);
or U657 (N_657,In_227,In_296);
nor U658 (N_658,In_640,In_22);
or U659 (N_659,In_527,In_585);
xnor U660 (N_660,In_29,In_569);
nor U661 (N_661,In_497,In_416);
nand U662 (N_662,In_250,In_195);
xnor U663 (N_663,In_34,In_304);
nor U664 (N_664,In_647,In_458);
nor U665 (N_665,In_415,In_498);
nor U666 (N_666,In_735,In_212);
xor U667 (N_667,In_658,In_53);
nor U668 (N_668,In_309,In_114);
nor U669 (N_669,In_141,In_746);
or U670 (N_670,In_160,In_297);
or U671 (N_671,In_134,In_365);
and U672 (N_672,In_285,In_539);
xor U673 (N_673,In_10,In_9);
and U674 (N_674,In_84,In_112);
nand U675 (N_675,In_594,In_30);
or U676 (N_676,In_294,In_533);
xor U677 (N_677,In_638,In_656);
nand U678 (N_678,In_37,In_313);
and U679 (N_679,In_713,In_515);
and U680 (N_680,In_613,In_728);
nor U681 (N_681,In_568,In_256);
xor U682 (N_682,In_90,In_297);
and U683 (N_683,In_314,In_532);
or U684 (N_684,In_184,In_54);
or U685 (N_685,In_707,In_419);
xor U686 (N_686,In_542,In_88);
xnor U687 (N_687,In_217,In_558);
nand U688 (N_688,In_207,In_688);
and U689 (N_689,In_462,In_360);
or U690 (N_690,In_183,In_467);
and U691 (N_691,In_285,In_737);
nand U692 (N_692,In_20,In_105);
and U693 (N_693,In_611,In_11);
nor U694 (N_694,In_392,In_383);
and U695 (N_695,In_124,In_369);
nand U696 (N_696,In_705,In_417);
nand U697 (N_697,In_498,In_182);
nor U698 (N_698,In_296,In_109);
nand U699 (N_699,In_531,In_633);
or U700 (N_700,In_711,In_138);
xnor U701 (N_701,In_407,In_645);
nor U702 (N_702,In_257,In_20);
or U703 (N_703,In_170,In_743);
xor U704 (N_704,In_367,In_604);
nand U705 (N_705,In_607,In_676);
and U706 (N_706,In_160,In_209);
or U707 (N_707,In_480,In_66);
nand U708 (N_708,In_584,In_27);
or U709 (N_709,In_552,In_654);
nor U710 (N_710,In_630,In_167);
nor U711 (N_711,In_1,In_421);
nand U712 (N_712,In_486,In_247);
xor U713 (N_713,In_304,In_319);
and U714 (N_714,In_283,In_314);
xnor U715 (N_715,In_273,In_677);
and U716 (N_716,In_466,In_684);
xnor U717 (N_717,In_341,In_720);
nand U718 (N_718,In_123,In_476);
and U719 (N_719,In_440,In_550);
xor U720 (N_720,In_661,In_557);
nor U721 (N_721,In_28,In_653);
nor U722 (N_722,In_651,In_211);
or U723 (N_723,In_10,In_55);
or U724 (N_724,In_452,In_259);
nor U725 (N_725,In_534,In_617);
nor U726 (N_726,In_111,In_51);
nand U727 (N_727,In_509,In_147);
or U728 (N_728,In_22,In_543);
xnor U729 (N_729,In_444,In_656);
or U730 (N_730,In_10,In_432);
xnor U731 (N_731,In_242,In_513);
xnor U732 (N_732,In_597,In_371);
nand U733 (N_733,In_615,In_697);
or U734 (N_734,In_389,In_666);
nor U735 (N_735,In_373,In_187);
nand U736 (N_736,In_153,In_539);
xnor U737 (N_737,In_573,In_175);
nor U738 (N_738,In_375,In_589);
xor U739 (N_739,In_624,In_197);
and U740 (N_740,In_687,In_724);
nand U741 (N_741,In_125,In_96);
and U742 (N_742,In_397,In_231);
nand U743 (N_743,In_626,In_692);
or U744 (N_744,In_678,In_300);
or U745 (N_745,In_48,In_651);
or U746 (N_746,In_61,In_514);
and U747 (N_747,In_378,In_686);
and U748 (N_748,In_404,In_613);
nand U749 (N_749,In_689,In_198);
and U750 (N_750,In_403,In_385);
or U751 (N_751,In_316,In_343);
and U752 (N_752,In_721,In_654);
nand U753 (N_753,In_647,In_684);
or U754 (N_754,In_648,In_213);
nor U755 (N_755,In_705,In_377);
or U756 (N_756,In_175,In_422);
nand U757 (N_757,In_305,In_125);
nand U758 (N_758,In_7,In_538);
xnor U759 (N_759,In_12,In_469);
or U760 (N_760,In_168,In_286);
and U761 (N_761,In_195,In_730);
nand U762 (N_762,In_269,In_544);
nand U763 (N_763,In_37,In_205);
xor U764 (N_764,In_359,In_319);
nand U765 (N_765,In_151,In_601);
nor U766 (N_766,In_248,In_307);
xor U767 (N_767,In_426,In_528);
or U768 (N_768,In_370,In_72);
xnor U769 (N_769,In_716,In_62);
xnor U770 (N_770,In_178,In_196);
nor U771 (N_771,In_504,In_593);
xnor U772 (N_772,In_190,In_257);
nand U773 (N_773,In_252,In_33);
nand U774 (N_774,In_215,In_728);
xnor U775 (N_775,In_105,In_520);
nand U776 (N_776,In_647,In_514);
or U777 (N_777,In_199,In_561);
and U778 (N_778,In_28,In_456);
nor U779 (N_779,In_274,In_216);
xor U780 (N_780,In_174,In_604);
and U781 (N_781,In_65,In_652);
nor U782 (N_782,In_392,In_502);
nor U783 (N_783,In_690,In_439);
and U784 (N_784,In_319,In_574);
and U785 (N_785,In_182,In_643);
nand U786 (N_786,In_236,In_748);
and U787 (N_787,In_616,In_60);
and U788 (N_788,In_617,In_280);
or U789 (N_789,In_158,In_509);
nor U790 (N_790,In_376,In_236);
xnor U791 (N_791,In_554,In_676);
xnor U792 (N_792,In_599,In_457);
nand U793 (N_793,In_460,In_382);
xor U794 (N_794,In_13,In_592);
nand U795 (N_795,In_430,In_208);
xnor U796 (N_796,In_271,In_564);
xor U797 (N_797,In_71,In_469);
and U798 (N_798,In_446,In_529);
and U799 (N_799,In_9,In_399);
nor U800 (N_800,In_466,In_279);
xor U801 (N_801,In_441,In_356);
nand U802 (N_802,In_507,In_135);
nor U803 (N_803,In_132,In_21);
nand U804 (N_804,In_713,In_159);
nor U805 (N_805,In_425,In_175);
xnor U806 (N_806,In_690,In_307);
or U807 (N_807,In_424,In_581);
nand U808 (N_808,In_252,In_272);
nand U809 (N_809,In_13,In_474);
and U810 (N_810,In_610,In_31);
xnor U811 (N_811,In_264,In_531);
and U812 (N_812,In_64,In_106);
or U813 (N_813,In_468,In_563);
nor U814 (N_814,In_556,In_118);
nor U815 (N_815,In_614,In_602);
or U816 (N_816,In_566,In_606);
and U817 (N_817,In_581,In_1);
nor U818 (N_818,In_330,In_92);
xnor U819 (N_819,In_709,In_97);
or U820 (N_820,In_529,In_171);
nor U821 (N_821,In_406,In_503);
nand U822 (N_822,In_240,In_347);
or U823 (N_823,In_621,In_605);
nand U824 (N_824,In_229,In_748);
xnor U825 (N_825,In_117,In_737);
and U826 (N_826,In_382,In_113);
nor U827 (N_827,In_73,In_378);
or U828 (N_828,In_378,In_377);
nand U829 (N_829,In_655,In_311);
nand U830 (N_830,In_390,In_726);
nand U831 (N_831,In_687,In_288);
nand U832 (N_832,In_648,In_373);
nand U833 (N_833,In_702,In_50);
nand U834 (N_834,In_426,In_436);
xnor U835 (N_835,In_142,In_78);
nor U836 (N_836,In_624,In_272);
nor U837 (N_837,In_147,In_199);
nor U838 (N_838,In_734,In_137);
xnor U839 (N_839,In_544,In_3);
or U840 (N_840,In_701,In_195);
nor U841 (N_841,In_694,In_434);
or U842 (N_842,In_89,In_79);
nand U843 (N_843,In_85,In_717);
nand U844 (N_844,In_461,In_625);
or U845 (N_845,In_252,In_242);
and U846 (N_846,In_399,In_400);
nor U847 (N_847,In_433,In_286);
nand U848 (N_848,In_503,In_289);
nor U849 (N_849,In_142,In_180);
and U850 (N_850,In_140,In_731);
or U851 (N_851,In_572,In_49);
nand U852 (N_852,In_455,In_311);
and U853 (N_853,In_505,In_68);
nand U854 (N_854,In_266,In_81);
or U855 (N_855,In_272,In_40);
xnor U856 (N_856,In_129,In_519);
nor U857 (N_857,In_512,In_744);
or U858 (N_858,In_216,In_644);
xor U859 (N_859,In_636,In_568);
nor U860 (N_860,In_626,In_546);
or U861 (N_861,In_396,In_360);
xor U862 (N_862,In_703,In_607);
or U863 (N_863,In_82,In_701);
nand U864 (N_864,In_531,In_126);
and U865 (N_865,In_513,In_316);
and U866 (N_866,In_2,In_438);
nand U867 (N_867,In_172,In_718);
or U868 (N_868,In_232,In_635);
and U869 (N_869,In_292,In_641);
xnor U870 (N_870,In_232,In_737);
and U871 (N_871,In_485,In_437);
and U872 (N_872,In_363,In_235);
xnor U873 (N_873,In_565,In_130);
nor U874 (N_874,In_12,In_564);
nor U875 (N_875,In_398,In_566);
or U876 (N_876,In_433,In_359);
or U877 (N_877,In_514,In_629);
xnor U878 (N_878,In_727,In_639);
or U879 (N_879,In_646,In_135);
or U880 (N_880,In_658,In_72);
nand U881 (N_881,In_215,In_140);
xor U882 (N_882,In_119,In_617);
nor U883 (N_883,In_132,In_17);
xnor U884 (N_884,In_667,In_300);
and U885 (N_885,In_373,In_569);
nor U886 (N_886,In_43,In_659);
nand U887 (N_887,In_422,In_447);
xor U888 (N_888,In_457,In_271);
nor U889 (N_889,In_90,In_82);
and U890 (N_890,In_329,In_641);
xor U891 (N_891,In_109,In_43);
nor U892 (N_892,In_672,In_480);
nor U893 (N_893,In_208,In_289);
nor U894 (N_894,In_217,In_27);
or U895 (N_895,In_668,In_32);
xor U896 (N_896,In_315,In_256);
nand U897 (N_897,In_66,In_741);
nand U898 (N_898,In_740,In_69);
xnor U899 (N_899,In_112,In_648);
or U900 (N_900,In_376,In_515);
xnor U901 (N_901,In_543,In_461);
and U902 (N_902,In_638,In_292);
and U903 (N_903,In_354,In_718);
nand U904 (N_904,In_493,In_507);
xnor U905 (N_905,In_66,In_344);
nand U906 (N_906,In_151,In_570);
and U907 (N_907,In_424,In_417);
nand U908 (N_908,In_447,In_454);
nor U909 (N_909,In_633,In_708);
xor U910 (N_910,In_667,In_106);
nor U911 (N_911,In_74,In_675);
or U912 (N_912,In_481,In_135);
and U913 (N_913,In_18,In_559);
nor U914 (N_914,In_322,In_690);
nand U915 (N_915,In_201,In_387);
nand U916 (N_916,In_160,In_409);
and U917 (N_917,In_556,In_539);
xnor U918 (N_918,In_658,In_501);
xor U919 (N_919,In_20,In_690);
xnor U920 (N_920,In_18,In_39);
nor U921 (N_921,In_544,In_480);
or U922 (N_922,In_739,In_326);
or U923 (N_923,In_240,In_739);
nor U924 (N_924,In_262,In_28);
nor U925 (N_925,In_552,In_535);
or U926 (N_926,In_274,In_394);
or U927 (N_927,In_59,In_579);
xor U928 (N_928,In_272,In_192);
xor U929 (N_929,In_452,In_96);
nor U930 (N_930,In_64,In_7);
nor U931 (N_931,In_300,In_124);
xor U932 (N_932,In_23,In_686);
and U933 (N_933,In_589,In_627);
nand U934 (N_934,In_550,In_498);
nor U935 (N_935,In_519,In_423);
and U936 (N_936,In_243,In_201);
nor U937 (N_937,In_476,In_225);
xor U938 (N_938,In_638,In_565);
nor U939 (N_939,In_306,In_550);
nor U940 (N_940,In_528,In_669);
nor U941 (N_941,In_582,In_246);
nor U942 (N_942,In_415,In_103);
or U943 (N_943,In_591,In_6);
xnor U944 (N_944,In_209,In_151);
and U945 (N_945,In_385,In_39);
nor U946 (N_946,In_22,In_21);
nand U947 (N_947,In_441,In_487);
nor U948 (N_948,In_33,In_484);
xor U949 (N_949,In_380,In_410);
and U950 (N_950,In_261,In_358);
and U951 (N_951,In_609,In_640);
and U952 (N_952,In_229,In_213);
nand U953 (N_953,In_207,In_403);
nor U954 (N_954,In_139,In_535);
nor U955 (N_955,In_485,In_355);
xor U956 (N_956,In_660,In_210);
or U957 (N_957,In_624,In_230);
nor U958 (N_958,In_497,In_631);
xor U959 (N_959,In_634,In_472);
or U960 (N_960,In_201,In_648);
and U961 (N_961,In_74,In_107);
nor U962 (N_962,In_202,In_275);
and U963 (N_963,In_713,In_716);
xor U964 (N_964,In_222,In_612);
nand U965 (N_965,In_684,In_718);
nand U966 (N_966,In_693,In_585);
xnor U967 (N_967,In_191,In_215);
or U968 (N_968,In_448,In_613);
and U969 (N_969,In_5,In_112);
nor U970 (N_970,In_7,In_456);
and U971 (N_971,In_489,In_252);
or U972 (N_972,In_137,In_351);
or U973 (N_973,In_373,In_527);
nand U974 (N_974,In_378,In_464);
xnor U975 (N_975,In_604,In_200);
and U976 (N_976,In_48,In_301);
or U977 (N_977,In_586,In_3);
nor U978 (N_978,In_419,In_633);
nor U979 (N_979,In_425,In_557);
or U980 (N_980,In_326,In_248);
or U981 (N_981,In_460,In_582);
or U982 (N_982,In_386,In_526);
nand U983 (N_983,In_547,In_11);
nand U984 (N_984,In_340,In_13);
nor U985 (N_985,In_168,In_242);
or U986 (N_986,In_566,In_379);
nand U987 (N_987,In_614,In_53);
xnor U988 (N_988,In_201,In_249);
nand U989 (N_989,In_36,In_547);
nor U990 (N_990,In_587,In_282);
xor U991 (N_991,In_194,In_398);
xnor U992 (N_992,In_56,In_562);
xnor U993 (N_993,In_470,In_65);
and U994 (N_994,In_401,In_747);
nand U995 (N_995,In_655,In_208);
and U996 (N_996,In_262,In_446);
or U997 (N_997,In_430,In_645);
nand U998 (N_998,In_249,In_718);
and U999 (N_999,In_698,In_254);
nand U1000 (N_1000,N_472,N_698);
nand U1001 (N_1001,N_536,N_270);
or U1002 (N_1002,N_150,N_413);
xnor U1003 (N_1003,N_576,N_902);
nor U1004 (N_1004,N_951,N_237);
xnor U1005 (N_1005,N_399,N_329);
nor U1006 (N_1006,N_671,N_913);
xnor U1007 (N_1007,N_464,N_262);
nor U1008 (N_1008,N_597,N_622);
and U1009 (N_1009,N_455,N_208);
and U1010 (N_1010,N_44,N_965);
nand U1011 (N_1011,N_719,N_403);
nand U1012 (N_1012,N_922,N_676);
or U1013 (N_1013,N_986,N_627);
and U1014 (N_1014,N_756,N_788);
nor U1015 (N_1015,N_117,N_699);
and U1016 (N_1016,N_351,N_625);
nor U1017 (N_1017,N_566,N_791);
or U1018 (N_1018,N_710,N_907);
or U1019 (N_1019,N_129,N_84);
nand U1020 (N_1020,N_310,N_532);
nor U1021 (N_1021,N_99,N_672);
or U1022 (N_1022,N_31,N_711);
or U1023 (N_1023,N_520,N_174);
nor U1024 (N_1024,N_517,N_892);
and U1025 (N_1025,N_445,N_164);
and U1026 (N_1026,N_289,N_496);
or U1027 (N_1027,N_666,N_934);
and U1028 (N_1028,N_790,N_100);
nand U1029 (N_1029,N_513,N_957);
or U1030 (N_1030,N_964,N_848);
nand U1031 (N_1031,N_786,N_346);
or U1032 (N_1032,N_578,N_628);
and U1033 (N_1033,N_102,N_746);
xnor U1034 (N_1034,N_658,N_897);
nand U1035 (N_1035,N_168,N_21);
or U1036 (N_1036,N_405,N_126);
nand U1037 (N_1037,N_758,N_211);
nand U1038 (N_1038,N_217,N_125);
xor U1039 (N_1039,N_905,N_384);
nand U1040 (N_1040,N_140,N_368);
or U1041 (N_1041,N_89,N_130);
or U1042 (N_1042,N_94,N_475);
nor U1043 (N_1043,N_400,N_610);
or U1044 (N_1044,N_912,N_669);
or U1045 (N_1045,N_814,N_233);
and U1046 (N_1046,N_352,N_919);
nor U1047 (N_1047,N_134,N_401);
nor U1048 (N_1048,N_460,N_603);
nor U1049 (N_1049,N_454,N_693);
xor U1050 (N_1050,N_937,N_663);
and U1051 (N_1051,N_205,N_250);
or U1052 (N_1052,N_728,N_203);
or U1053 (N_1053,N_773,N_884);
and U1054 (N_1054,N_583,N_426);
nand U1055 (N_1055,N_362,N_458);
nor U1056 (N_1056,N_406,N_960);
nor U1057 (N_1057,N_56,N_969);
nand U1058 (N_1058,N_124,N_223);
nor U1059 (N_1059,N_192,N_879);
xor U1060 (N_1060,N_421,N_579);
and U1061 (N_1061,N_556,N_999);
xnor U1062 (N_1062,N_651,N_643);
and U1063 (N_1063,N_506,N_569);
nor U1064 (N_1064,N_936,N_909);
nand U1065 (N_1065,N_732,N_623);
xnor U1066 (N_1066,N_383,N_335);
nor U1067 (N_1067,N_255,N_197);
xor U1068 (N_1068,N_325,N_570);
and U1069 (N_1069,N_260,N_135);
or U1070 (N_1070,N_248,N_928);
and U1071 (N_1071,N_468,N_862);
xor U1072 (N_1072,N_883,N_62);
or U1073 (N_1073,N_704,N_678);
nor U1074 (N_1074,N_200,N_77);
xor U1075 (N_1075,N_314,N_420);
nor U1076 (N_1076,N_530,N_615);
xnor U1077 (N_1077,N_462,N_794);
xnor U1078 (N_1078,N_575,N_187);
and U1079 (N_1079,N_785,N_272);
nor U1080 (N_1080,N_37,N_253);
or U1081 (N_1081,N_280,N_846);
and U1082 (N_1082,N_179,N_59);
nand U1083 (N_1083,N_30,N_221);
nand U1084 (N_1084,N_12,N_57);
nor U1085 (N_1085,N_545,N_1);
and U1086 (N_1086,N_984,N_473);
or U1087 (N_1087,N_602,N_165);
xnor U1088 (N_1088,N_238,N_65);
xnor U1089 (N_1089,N_642,N_474);
or U1090 (N_1090,N_370,N_561);
nand U1091 (N_1091,N_844,N_730);
nand U1092 (N_1092,N_103,N_166);
xnor U1093 (N_1093,N_22,N_149);
and U1094 (N_1094,N_596,N_55);
or U1095 (N_1095,N_157,N_201);
nand U1096 (N_1096,N_144,N_820);
xnor U1097 (N_1097,N_116,N_747);
nand U1098 (N_1098,N_664,N_774);
nor U1099 (N_1099,N_754,N_595);
or U1100 (N_1100,N_618,N_921);
nor U1101 (N_1101,N_874,N_234);
and U1102 (N_1102,N_482,N_833);
and U1103 (N_1103,N_298,N_387);
nand U1104 (N_1104,N_621,N_364);
nor U1105 (N_1105,N_619,N_261);
xnor U1106 (N_1106,N_268,N_834);
nor U1107 (N_1107,N_493,N_981);
and U1108 (N_1108,N_590,N_617);
nor U1109 (N_1109,N_680,N_613);
nand U1110 (N_1110,N_654,N_751);
and U1111 (N_1111,N_489,N_151);
and U1112 (N_1112,N_818,N_558);
nor U1113 (N_1113,N_342,N_690);
nor U1114 (N_1114,N_41,N_19);
xnor U1115 (N_1115,N_216,N_956);
and U1116 (N_1116,N_373,N_374);
and U1117 (N_1117,N_191,N_859);
xnor U1118 (N_1118,N_692,N_817);
or U1119 (N_1119,N_51,N_600);
or U1120 (N_1120,N_341,N_550);
nor U1121 (N_1121,N_92,N_868);
xor U1122 (N_1122,N_313,N_772);
and U1123 (N_1123,N_273,N_224);
nand U1124 (N_1124,N_819,N_543);
nor U1125 (N_1125,N_620,N_648);
or U1126 (N_1126,N_703,N_444);
or U1127 (N_1127,N_91,N_988);
nor U1128 (N_1128,N_682,N_305);
nand U1129 (N_1129,N_229,N_733);
and U1130 (N_1130,N_968,N_837);
nand U1131 (N_1131,N_891,N_835);
nand U1132 (N_1132,N_43,N_990);
or U1133 (N_1133,N_511,N_86);
or U1134 (N_1134,N_867,N_656);
or U1135 (N_1135,N_688,N_687);
xnor U1136 (N_1136,N_955,N_152);
and U1137 (N_1137,N_283,N_170);
nand U1138 (N_1138,N_39,N_795);
and U1139 (N_1139,N_562,N_809);
and U1140 (N_1140,N_748,N_750);
and U1141 (N_1141,N_153,N_213);
nor U1142 (N_1142,N_802,N_184);
or U1143 (N_1143,N_34,N_525);
or U1144 (N_1144,N_391,N_10);
and U1145 (N_1145,N_592,N_294);
and U1146 (N_1146,N_32,N_29);
or U1147 (N_1147,N_186,N_829);
xnor U1148 (N_1148,N_207,N_198);
xnor U1149 (N_1149,N_626,N_498);
nand U1150 (N_1150,N_488,N_548);
xor U1151 (N_1151,N_549,N_243);
nor U1152 (N_1152,N_348,N_23);
xor U1153 (N_1153,N_942,N_667);
nor U1154 (N_1154,N_966,N_584);
xnor U1155 (N_1155,N_958,N_853);
nand U1156 (N_1156,N_898,N_98);
nor U1157 (N_1157,N_247,N_158);
or U1158 (N_1158,N_553,N_507);
nor U1159 (N_1159,N_587,N_755);
and U1160 (N_1160,N_202,N_641);
nor U1161 (N_1161,N_638,N_204);
or U1162 (N_1162,N_428,N_823);
xor U1163 (N_1163,N_457,N_118);
xor U1164 (N_1164,N_604,N_514);
xor U1165 (N_1165,N_78,N_895);
xnor U1166 (N_1166,N_308,N_903);
nor U1167 (N_1167,N_74,N_167);
xor U1168 (N_1168,N_175,N_48);
or U1169 (N_1169,N_718,N_299);
nor U1170 (N_1170,N_259,N_850);
xnor U1171 (N_1171,N_614,N_531);
xor U1172 (N_1172,N_822,N_736);
nand U1173 (N_1173,N_855,N_605);
nor U1174 (N_1174,N_963,N_265);
and U1175 (N_1175,N_24,N_155);
and U1176 (N_1176,N_64,N_887);
nand U1177 (N_1177,N_141,N_353);
and U1178 (N_1178,N_504,N_477);
nand U1179 (N_1179,N_251,N_431);
xor U1180 (N_1180,N_447,N_6);
or U1181 (N_1181,N_67,N_529);
or U1182 (N_1182,N_226,N_630);
nand U1183 (N_1183,N_744,N_307);
and U1184 (N_1184,N_894,N_2);
xnor U1185 (N_1185,N_63,N_696);
nor U1186 (N_1186,N_408,N_541);
nand U1187 (N_1187,N_714,N_206);
xor U1188 (N_1188,N_275,N_412);
and U1189 (N_1189,N_385,N_925);
and U1190 (N_1190,N_392,N_97);
and U1191 (N_1191,N_559,N_586);
xnor U1192 (N_1192,N_396,N_712);
or U1193 (N_1193,N_231,N_194);
nor U1194 (N_1194,N_832,N_568);
and U1195 (N_1195,N_826,N_441);
nor U1196 (N_1196,N_232,N_589);
and U1197 (N_1197,N_611,N_330);
xor U1198 (N_1198,N_560,N_297);
nand U1199 (N_1199,N_683,N_81);
or U1200 (N_1200,N_14,N_737);
and U1201 (N_1201,N_673,N_143);
or U1202 (N_1202,N_674,N_939);
and U1203 (N_1203,N_300,N_527);
xor U1204 (N_1204,N_96,N_865);
nand U1205 (N_1205,N_948,N_378);
xnor U1206 (N_1206,N_371,N_389);
nor U1207 (N_1207,N_707,N_292);
nand U1208 (N_1208,N_442,N_784);
nand U1209 (N_1209,N_776,N_222);
and U1210 (N_1210,N_872,N_847);
and U1211 (N_1211,N_881,N_128);
and U1212 (N_1212,N_524,N_974);
and U1213 (N_1213,N_176,N_775);
xnor U1214 (N_1214,N_418,N_146);
or U1215 (N_1215,N_411,N_920);
and U1216 (N_1216,N_177,N_888);
xnor U1217 (N_1217,N_899,N_662);
xnor U1218 (N_1218,N_101,N_713);
and U1219 (N_1219,N_681,N_269);
or U1220 (N_1220,N_148,N_388);
xor U1221 (N_1221,N_114,N_427);
xor U1222 (N_1222,N_950,N_311);
or U1223 (N_1223,N_398,N_293);
and U1224 (N_1224,N_246,N_691);
and U1225 (N_1225,N_528,N_321);
nor U1226 (N_1226,N_563,N_731);
nor U1227 (N_1227,N_959,N_797);
or U1228 (N_1228,N_456,N_813);
and U1229 (N_1229,N_212,N_914);
nor U1230 (N_1230,N_869,N_841);
or U1231 (N_1231,N_766,N_107);
nand U1232 (N_1232,N_734,N_769);
and U1233 (N_1233,N_432,N_616);
nor U1234 (N_1234,N_646,N_980);
xor U1235 (N_1235,N_480,N_580);
xor U1236 (N_1236,N_705,N_375);
and U1237 (N_1237,N_356,N_838);
and U1238 (N_1238,N_286,N_634);
xnor U1239 (N_1239,N_66,N_133);
and U1240 (N_1240,N_11,N_975);
nor U1241 (N_1241,N_193,N_953);
and U1242 (N_1242,N_228,N_369);
or U1243 (N_1243,N_857,N_5);
nor U1244 (N_1244,N_635,N_161);
and U1245 (N_1245,N_448,N_136);
nand U1246 (N_1246,N_180,N_303);
nand U1247 (N_1247,N_123,N_295);
and U1248 (N_1248,N_471,N_76);
nand U1249 (N_1249,N_196,N_893);
nand U1250 (N_1250,N_104,N_591);
or U1251 (N_1251,N_416,N_75);
or U1252 (N_1252,N_106,N_73);
or U1253 (N_1253,N_332,N_533);
or U1254 (N_1254,N_831,N_555);
or U1255 (N_1255,N_497,N_740);
nor U1256 (N_1256,N_17,N_915);
and U1257 (N_1257,N_808,N_320);
nor U1258 (N_1258,N_544,N_105);
nand U1259 (N_1259,N_652,N_328);
xor U1260 (N_1260,N_230,N_402);
and U1261 (N_1261,N_476,N_762);
and U1262 (N_1262,N_377,N_612);
xor U1263 (N_1263,N_876,N_924);
nand U1264 (N_1264,N_763,N_521);
or U1265 (N_1265,N_644,N_564);
or U1266 (N_1266,N_18,N_417);
nand U1267 (N_1267,N_944,N_169);
nor U1268 (N_1268,N_565,N_923);
nor U1269 (N_1269,N_20,N_410);
and U1270 (N_1270,N_429,N_885);
and U1271 (N_1271,N_875,N_910);
and U1272 (N_1272,N_787,N_749);
nand U1273 (N_1273,N_120,N_440);
nor U1274 (N_1274,N_941,N_962);
nand U1275 (N_1275,N_390,N_866);
nand U1276 (N_1276,N_677,N_985);
or U1277 (N_1277,N_350,N_800);
xor U1278 (N_1278,N_967,N_119);
and U1279 (N_1279,N_694,N_633);
xor U1280 (N_1280,N_499,N_864);
and U1281 (N_1281,N_381,N_483);
and U1282 (N_1282,N_873,N_199);
xor U1283 (N_1283,N_535,N_240);
and U1284 (N_1284,N_281,N_172);
nand U1285 (N_1285,N_121,N_154);
nand U1286 (N_1286,N_380,N_706);
or U1287 (N_1287,N_492,N_276);
and U1288 (N_1288,N_995,N_929);
nor U1289 (N_1289,N_799,N_282);
nand U1290 (N_1290,N_190,N_954);
nor U1291 (N_1291,N_552,N_82);
nand U1292 (N_1292,N_494,N_318);
nor U1293 (N_1293,N_349,N_573);
xor U1294 (N_1294,N_804,N_26);
nor U1295 (N_1295,N_113,N_52);
and U1296 (N_1296,N_998,N_434);
and U1297 (N_1297,N_162,N_509);
or U1298 (N_1298,N_340,N_111);
or U1299 (N_1299,N_856,N_469);
or U1300 (N_1300,N_395,N_979);
or U1301 (N_1301,N_721,N_365);
or U1302 (N_1302,N_145,N_242);
or U1303 (N_1303,N_931,N_854);
and U1304 (N_1304,N_779,N_650);
and U1305 (N_1305,N_970,N_996);
xnor U1306 (N_1306,N_323,N_220);
or U1307 (N_1307,N_210,N_911);
or U1308 (N_1308,N_88,N_236);
and U1309 (N_1309,N_239,N_639);
nor U1310 (N_1310,N_13,N_28);
or U1311 (N_1311,N_3,N_842);
and U1312 (N_1312,N_752,N_689);
xor U1313 (N_1313,N_816,N_79);
nor U1314 (N_1314,N_505,N_83);
nor U1315 (N_1315,N_46,N_463);
and U1316 (N_1316,N_764,N_249);
and U1317 (N_1317,N_753,N_68);
or U1318 (N_1318,N_547,N_219);
nor U1319 (N_1319,N_309,N_274);
nand U1320 (N_1320,N_852,N_685);
xor U1321 (N_1321,N_945,N_871);
nor U1322 (N_1322,N_594,N_337);
xor U1323 (N_1323,N_363,N_486);
and U1324 (N_1324,N_810,N_163);
and U1325 (N_1325,N_495,N_636);
nand U1326 (N_1326,N_306,N_424);
nand U1327 (N_1327,N_745,N_354);
nor U1328 (N_1328,N_640,N_508);
nand U1329 (N_1329,N_729,N_252);
nor U1330 (N_1330,N_423,N_726);
or U1331 (N_1331,N_93,N_132);
xor U1332 (N_1332,N_142,N_112);
or U1333 (N_1333,N_539,N_870);
or U1334 (N_1334,N_812,N_933);
and U1335 (N_1335,N_478,N_993);
nand U1336 (N_1336,N_987,N_173);
nor U1337 (N_1337,N_322,N_502);
nand U1338 (N_1338,N_782,N_256);
and U1339 (N_1339,N_4,N_684);
or U1340 (N_1340,N_279,N_244);
nand U1341 (N_1341,N_554,N_930);
nor U1342 (N_1342,N_61,N_697);
nor U1343 (N_1343,N_333,N_765);
nand U1344 (N_1344,N_339,N_843);
or U1345 (N_1345,N_830,N_304);
and U1346 (N_1346,N_245,N_708);
or U1347 (N_1347,N_302,N_572);
or U1348 (N_1348,N_459,N_357);
nand U1349 (N_1349,N_827,N_160);
and U1350 (N_1350,N_315,N_15);
nand U1351 (N_1351,N_825,N_637);
nand U1352 (N_1352,N_422,N_845);
and U1353 (N_1353,N_394,N_742);
xor U1354 (N_1354,N_336,N_404);
or U1355 (N_1355,N_451,N_479);
or U1356 (N_1356,N_901,N_860);
and U1357 (N_1357,N_811,N_465);
nor U1358 (N_1358,N_917,N_906);
and U1359 (N_1359,N_58,N_438);
and U1360 (N_1360,N_645,N_185);
or U1361 (N_1361,N_338,N_886);
nor U1362 (N_1362,N_85,N_258);
and U1363 (N_1363,N_519,N_947);
or U1364 (N_1364,N_367,N_631);
xnor U1365 (N_1365,N_889,N_271);
and U1366 (N_1366,N_598,N_110);
xor U1367 (N_1367,N_334,N_659);
nand U1368 (N_1368,N_661,N_227);
or U1369 (N_1369,N_461,N_491);
nand U1370 (N_1370,N_358,N_49);
or U1371 (N_1371,N_670,N_538);
nor U1372 (N_1372,N_436,N_481);
nor U1373 (N_1373,N_437,N_943);
xor U1374 (N_1374,N_526,N_588);
nor U1375 (N_1375,N_409,N_700);
or U1376 (N_1376,N_858,N_803);
and U1377 (N_1377,N_127,N_653);
nand U1378 (N_1378,N_296,N_137);
and U1379 (N_1379,N_815,N_977);
and U1380 (N_1380,N_880,N_382);
nand U1381 (N_1381,N_551,N_961);
or U1382 (N_1382,N_38,N_761);
and U1383 (N_1383,N_319,N_989);
or U1384 (N_1384,N_71,N_178);
nor U1385 (N_1385,N_821,N_500);
nor U1386 (N_1386,N_971,N_156);
and U1387 (N_1387,N_940,N_430);
and U1388 (N_1388,N_33,N_757);
xnor U1389 (N_1389,N_972,N_702);
or U1390 (N_1390,N_288,N_537);
or U1391 (N_1391,N_655,N_601);
nand U1392 (N_1392,N_277,N_415);
nor U1393 (N_1393,N_189,N_789);
or U1394 (N_1394,N_840,N_397);
or U1395 (N_1395,N_890,N_345);
xnor U1396 (N_1396,N_978,N_938);
nand U1397 (N_1397,N_425,N_9);
nor U1398 (N_1398,N_647,N_278);
or U1399 (N_1399,N_777,N_443);
nand U1400 (N_1400,N_379,N_376);
or U1401 (N_1401,N_87,N_466);
nor U1402 (N_1402,N_768,N_534);
and U1403 (N_1403,N_490,N_632);
nor U1404 (N_1404,N_324,N_723);
or U1405 (N_1405,N_904,N_257);
nand U1406 (N_1406,N_72,N_805);
xnor U1407 (N_1407,N_743,N_908);
or U1408 (N_1408,N_686,N_585);
nand U1409 (N_1409,N_608,N_649);
xnor U1410 (N_1410,N_824,N_188);
xnor U1411 (N_1411,N_759,N_982);
and U1412 (N_1412,N_796,N_446);
nor U1413 (N_1413,N_69,N_331);
nor U1414 (N_1414,N_53,N_781);
nor U1415 (N_1415,N_571,N_522);
nor U1416 (N_1416,N_657,N_523);
nand U1417 (N_1417,N_629,N_828);
xor U1418 (N_1418,N_992,N_209);
xor U1419 (N_1419,N_439,N_147);
nor U1420 (N_1420,N_326,N_593);
xor U1421 (N_1421,N_183,N_574);
or U1422 (N_1422,N_516,N_839);
nand U1423 (N_1423,N_806,N_717);
and U1424 (N_1424,N_582,N_878);
xor U1425 (N_1425,N_42,N_312);
nor U1426 (N_1426,N_952,N_836);
or U1427 (N_1427,N_793,N_567);
xnor U1428 (N_1428,N_433,N_360);
nor U1429 (N_1429,N_109,N_991);
or U1430 (N_1430,N_994,N_372);
nor U1431 (N_1431,N_770,N_927);
or U1432 (N_1432,N_877,N_316);
and U1433 (N_1433,N_218,N_54);
and U1434 (N_1434,N_503,N_946);
xor U1435 (N_1435,N_95,N_361);
or U1436 (N_1436,N_181,N_861);
nor U1437 (N_1437,N_679,N_435);
and U1438 (N_1438,N_918,N_414);
xor U1439 (N_1439,N_393,N_139);
or U1440 (N_1440,N_735,N_783);
nor U1441 (N_1441,N_36,N_542);
nand U1442 (N_1442,N_983,N_215);
and U1443 (N_1443,N_599,N_668);
nor U1444 (N_1444,N_449,N_171);
xnor U1445 (N_1445,N_675,N_182);
xnor U1446 (N_1446,N_863,N_16);
and U1447 (N_1447,N_290,N_467);
and U1448 (N_1448,N_267,N_347);
xor U1449 (N_1449,N_355,N_900);
nand U1450 (N_1450,N_701,N_487);
and U1451 (N_1451,N_896,N_882);
and U1452 (N_1452,N_501,N_973);
or U1453 (N_1453,N_624,N_291);
nor U1454 (N_1454,N_515,N_778);
xnor U1455 (N_1455,N_609,N_285);
xor U1456 (N_1456,N_45,N_115);
nor U1457 (N_1457,N_715,N_108);
nand U1458 (N_1458,N_518,N_716);
xnor U1459 (N_1459,N_131,N_607);
xor U1460 (N_1460,N_577,N_581);
xnor U1461 (N_1461,N_660,N_997);
nand U1462 (N_1462,N_301,N_90);
xor U1463 (N_1463,N_8,N_807);
and U1464 (N_1464,N_40,N_159);
nor U1465 (N_1465,N_709,N_725);
and U1466 (N_1466,N_47,N_540);
and U1467 (N_1467,N_485,N_738);
nand U1468 (N_1468,N_450,N_287);
or U1469 (N_1469,N_386,N_949);
xor U1470 (N_1470,N_195,N_916);
and U1471 (N_1471,N_122,N_557);
or U1472 (N_1472,N_317,N_512);
nor U1473 (N_1473,N_798,N_27);
or U1474 (N_1474,N_767,N_546);
nand U1475 (N_1475,N_80,N_727);
nor U1476 (N_1476,N_50,N_932);
or U1477 (N_1477,N_263,N_935);
nor U1478 (N_1478,N_470,N_343);
xnor U1479 (N_1479,N_35,N_254);
and U1480 (N_1480,N_771,N_695);
or U1481 (N_1481,N_484,N_366);
and U1482 (N_1482,N_926,N_722);
nor U1483 (N_1483,N_976,N_665);
nand U1484 (N_1484,N_70,N_453);
nand U1485 (N_1485,N_7,N_60);
xnor U1486 (N_1486,N_327,N_849);
and U1487 (N_1487,N_235,N_606);
or U1488 (N_1488,N_266,N_792);
nand U1489 (N_1489,N_419,N_452);
xnor U1490 (N_1490,N_214,N_760);
or U1491 (N_1491,N_284,N_225);
and U1492 (N_1492,N_241,N_739);
and U1493 (N_1493,N_780,N_138);
or U1494 (N_1494,N_720,N_344);
and U1495 (N_1495,N_25,N_359);
nor U1496 (N_1496,N_851,N_264);
nand U1497 (N_1497,N_724,N_741);
xor U1498 (N_1498,N_0,N_407);
and U1499 (N_1499,N_801,N_510);
xnor U1500 (N_1500,N_396,N_508);
nand U1501 (N_1501,N_835,N_787);
and U1502 (N_1502,N_793,N_229);
nand U1503 (N_1503,N_422,N_538);
or U1504 (N_1504,N_22,N_452);
nor U1505 (N_1505,N_327,N_195);
nor U1506 (N_1506,N_792,N_370);
nand U1507 (N_1507,N_415,N_30);
xor U1508 (N_1508,N_492,N_487);
nor U1509 (N_1509,N_336,N_436);
xnor U1510 (N_1510,N_755,N_547);
or U1511 (N_1511,N_534,N_933);
and U1512 (N_1512,N_345,N_328);
nand U1513 (N_1513,N_344,N_835);
nand U1514 (N_1514,N_124,N_588);
xnor U1515 (N_1515,N_617,N_939);
and U1516 (N_1516,N_404,N_907);
nor U1517 (N_1517,N_978,N_131);
xor U1518 (N_1518,N_550,N_717);
nand U1519 (N_1519,N_425,N_670);
nand U1520 (N_1520,N_445,N_499);
nand U1521 (N_1521,N_946,N_656);
nor U1522 (N_1522,N_898,N_767);
or U1523 (N_1523,N_138,N_812);
nor U1524 (N_1524,N_797,N_755);
nand U1525 (N_1525,N_337,N_373);
nand U1526 (N_1526,N_617,N_514);
nand U1527 (N_1527,N_218,N_52);
nand U1528 (N_1528,N_395,N_929);
and U1529 (N_1529,N_521,N_860);
nor U1530 (N_1530,N_551,N_636);
nand U1531 (N_1531,N_61,N_94);
xor U1532 (N_1532,N_43,N_772);
and U1533 (N_1533,N_500,N_631);
and U1534 (N_1534,N_593,N_798);
and U1535 (N_1535,N_456,N_514);
and U1536 (N_1536,N_977,N_244);
xor U1537 (N_1537,N_995,N_225);
nor U1538 (N_1538,N_564,N_206);
nor U1539 (N_1539,N_684,N_977);
and U1540 (N_1540,N_262,N_834);
xor U1541 (N_1541,N_533,N_24);
nand U1542 (N_1542,N_0,N_51);
nor U1543 (N_1543,N_910,N_437);
nand U1544 (N_1544,N_974,N_301);
xor U1545 (N_1545,N_855,N_599);
nor U1546 (N_1546,N_137,N_164);
and U1547 (N_1547,N_537,N_920);
xnor U1548 (N_1548,N_345,N_646);
xor U1549 (N_1549,N_821,N_258);
or U1550 (N_1550,N_610,N_593);
nand U1551 (N_1551,N_498,N_418);
nor U1552 (N_1552,N_502,N_791);
nor U1553 (N_1553,N_145,N_479);
or U1554 (N_1554,N_878,N_595);
nand U1555 (N_1555,N_114,N_47);
xor U1556 (N_1556,N_426,N_898);
nand U1557 (N_1557,N_576,N_626);
or U1558 (N_1558,N_530,N_965);
and U1559 (N_1559,N_723,N_184);
nor U1560 (N_1560,N_725,N_755);
or U1561 (N_1561,N_906,N_335);
nor U1562 (N_1562,N_846,N_140);
and U1563 (N_1563,N_156,N_798);
or U1564 (N_1564,N_93,N_175);
nand U1565 (N_1565,N_31,N_442);
xor U1566 (N_1566,N_746,N_821);
or U1567 (N_1567,N_511,N_108);
or U1568 (N_1568,N_240,N_445);
or U1569 (N_1569,N_169,N_634);
xnor U1570 (N_1570,N_605,N_506);
and U1571 (N_1571,N_316,N_675);
nor U1572 (N_1572,N_650,N_62);
and U1573 (N_1573,N_717,N_736);
or U1574 (N_1574,N_140,N_946);
nor U1575 (N_1575,N_783,N_713);
xnor U1576 (N_1576,N_371,N_802);
and U1577 (N_1577,N_482,N_363);
or U1578 (N_1578,N_173,N_853);
and U1579 (N_1579,N_948,N_143);
or U1580 (N_1580,N_455,N_476);
nand U1581 (N_1581,N_504,N_873);
or U1582 (N_1582,N_124,N_67);
nor U1583 (N_1583,N_46,N_196);
or U1584 (N_1584,N_650,N_97);
and U1585 (N_1585,N_371,N_584);
nand U1586 (N_1586,N_740,N_137);
and U1587 (N_1587,N_363,N_176);
and U1588 (N_1588,N_629,N_569);
nand U1589 (N_1589,N_69,N_966);
or U1590 (N_1590,N_24,N_651);
and U1591 (N_1591,N_153,N_940);
xor U1592 (N_1592,N_769,N_43);
and U1593 (N_1593,N_558,N_443);
or U1594 (N_1594,N_215,N_476);
nand U1595 (N_1595,N_688,N_736);
nand U1596 (N_1596,N_291,N_29);
or U1597 (N_1597,N_266,N_674);
nand U1598 (N_1598,N_592,N_675);
or U1599 (N_1599,N_682,N_386);
and U1600 (N_1600,N_644,N_841);
nand U1601 (N_1601,N_557,N_8);
and U1602 (N_1602,N_330,N_143);
nand U1603 (N_1603,N_563,N_687);
nand U1604 (N_1604,N_945,N_877);
xor U1605 (N_1605,N_693,N_498);
and U1606 (N_1606,N_48,N_998);
nand U1607 (N_1607,N_821,N_599);
xnor U1608 (N_1608,N_136,N_142);
or U1609 (N_1609,N_953,N_344);
nor U1610 (N_1610,N_478,N_989);
xnor U1611 (N_1611,N_165,N_88);
or U1612 (N_1612,N_182,N_293);
nor U1613 (N_1613,N_11,N_416);
nand U1614 (N_1614,N_3,N_708);
nand U1615 (N_1615,N_941,N_292);
nand U1616 (N_1616,N_555,N_834);
and U1617 (N_1617,N_462,N_10);
nor U1618 (N_1618,N_513,N_794);
and U1619 (N_1619,N_928,N_30);
or U1620 (N_1620,N_1,N_611);
xor U1621 (N_1621,N_714,N_274);
nor U1622 (N_1622,N_676,N_727);
nand U1623 (N_1623,N_233,N_942);
nand U1624 (N_1624,N_309,N_645);
and U1625 (N_1625,N_34,N_270);
or U1626 (N_1626,N_624,N_886);
nor U1627 (N_1627,N_57,N_296);
xnor U1628 (N_1628,N_960,N_428);
or U1629 (N_1629,N_867,N_7);
and U1630 (N_1630,N_319,N_811);
or U1631 (N_1631,N_55,N_920);
and U1632 (N_1632,N_587,N_238);
xnor U1633 (N_1633,N_740,N_736);
nor U1634 (N_1634,N_233,N_395);
nand U1635 (N_1635,N_773,N_665);
nand U1636 (N_1636,N_83,N_969);
xor U1637 (N_1637,N_940,N_884);
xnor U1638 (N_1638,N_76,N_141);
xnor U1639 (N_1639,N_791,N_116);
nor U1640 (N_1640,N_843,N_243);
nand U1641 (N_1641,N_203,N_486);
and U1642 (N_1642,N_259,N_703);
nor U1643 (N_1643,N_469,N_808);
or U1644 (N_1644,N_324,N_201);
and U1645 (N_1645,N_426,N_467);
nand U1646 (N_1646,N_363,N_615);
or U1647 (N_1647,N_834,N_579);
nand U1648 (N_1648,N_217,N_498);
nand U1649 (N_1649,N_448,N_568);
xor U1650 (N_1650,N_247,N_161);
xnor U1651 (N_1651,N_179,N_227);
xor U1652 (N_1652,N_762,N_475);
nand U1653 (N_1653,N_103,N_750);
and U1654 (N_1654,N_838,N_115);
nand U1655 (N_1655,N_592,N_953);
and U1656 (N_1656,N_138,N_329);
or U1657 (N_1657,N_678,N_951);
and U1658 (N_1658,N_2,N_183);
nand U1659 (N_1659,N_73,N_504);
nor U1660 (N_1660,N_443,N_470);
and U1661 (N_1661,N_117,N_825);
or U1662 (N_1662,N_225,N_744);
nor U1663 (N_1663,N_469,N_196);
nand U1664 (N_1664,N_511,N_759);
and U1665 (N_1665,N_256,N_550);
xor U1666 (N_1666,N_618,N_665);
nand U1667 (N_1667,N_121,N_413);
or U1668 (N_1668,N_458,N_871);
nand U1669 (N_1669,N_60,N_580);
and U1670 (N_1670,N_954,N_408);
xnor U1671 (N_1671,N_634,N_917);
xor U1672 (N_1672,N_516,N_934);
nor U1673 (N_1673,N_13,N_380);
xnor U1674 (N_1674,N_345,N_510);
or U1675 (N_1675,N_866,N_923);
or U1676 (N_1676,N_285,N_477);
xnor U1677 (N_1677,N_332,N_275);
nor U1678 (N_1678,N_547,N_618);
xor U1679 (N_1679,N_263,N_326);
or U1680 (N_1680,N_496,N_67);
nor U1681 (N_1681,N_782,N_615);
nor U1682 (N_1682,N_204,N_98);
xor U1683 (N_1683,N_643,N_352);
and U1684 (N_1684,N_648,N_211);
xnor U1685 (N_1685,N_233,N_743);
nand U1686 (N_1686,N_138,N_574);
or U1687 (N_1687,N_573,N_490);
nor U1688 (N_1688,N_552,N_180);
or U1689 (N_1689,N_607,N_115);
nor U1690 (N_1690,N_133,N_339);
or U1691 (N_1691,N_460,N_569);
xnor U1692 (N_1692,N_915,N_93);
xor U1693 (N_1693,N_350,N_836);
and U1694 (N_1694,N_995,N_229);
nand U1695 (N_1695,N_901,N_699);
nor U1696 (N_1696,N_816,N_402);
nand U1697 (N_1697,N_68,N_248);
nand U1698 (N_1698,N_90,N_316);
or U1699 (N_1699,N_784,N_128);
xor U1700 (N_1700,N_818,N_83);
nand U1701 (N_1701,N_99,N_128);
nor U1702 (N_1702,N_255,N_505);
nand U1703 (N_1703,N_478,N_258);
and U1704 (N_1704,N_573,N_24);
nor U1705 (N_1705,N_472,N_21);
xor U1706 (N_1706,N_934,N_164);
or U1707 (N_1707,N_327,N_102);
or U1708 (N_1708,N_672,N_658);
nor U1709 (N_1709,N_724,N_167);
nand U1710 (N_1710,N_560,N_574);
or U1711 (N_1711,N_138,N_560);
nand U1712 (N_1712,N_54,N_409);
nor U1713 (N_1713,N_438,N_622);
xnor U1714 (N_1714,N_573,N_597);
and U1715 (N_1715,N_362,N_618);
nand U1716 (N_1716,N_217,N_28);
nor U1717 (N_1717,N_572,N_298);
nor U1718 (N_1718,N_944,N_851);
nand U1719 (N_1719,N_888,N_603);
nor U1720 (N_1720,N_304,N_41);
nor U1721 (N_1721,N_269,N_166);
nand U1722 (N_1722,N_576,N_48);
xnor U1723 (N_1723,N_317,N_977);
or U1724 (N_1724,N_282,N_482);
and U1725 (N_1725,N_64,N_220);
and U1726 (N_1726,N_655,N_350);
nand U1727 (N_1727,N_820,N_745);
nand U1728 (N_1728,N_855,N_937);
or U1729 (N_1729,N_314,N_741);
nand U1730 (N_1730,N_488,N_506);
or U1731 (N_1731,N_731,N_652);
and U1732 (N_1732,N_768,N_245);
nor U1733 (N_1733,N_989,N_620);
nand U1734 (N_1734,N_646,N_179);
nor U1735 (N_1735,N_504,N_322);
and U1736 (N_1736,N_808,N_91);
nand U1737 (N_1737,N_621,N_338);
or U1738 (N_1738,N_975,N_406);
nand U1739 (N_1739,N_420,N_240);
and U1740 (N_1740,N_339,N_4);
nand U1741 (N_1741,N_217,N_687);
or U1742 (N_1742,N_807,N_839);
xor U1743 (N_1743,N_565,N_423);
and U1744 (N_1744,N_108,N_250);
nand U1745 (N_1745,N_456,N_848);
xnor U1746 (N_1746,N_250,N_941);
or U1747 (N_1747,N_40,N_831);
nand U1748 (N_1748,N_404,N_634);
or U1749 (N_1749,N_107,N_188);
or U1750 (N_1750,N_576,N_280);
xor U1751 (N_1751,N_706,N_903);
nor U1752 (N_1752,N_75,N_870);
or U1753 (N_1753,N_429,N_777);
nor U1754 (N_1754,N_391,N_939);
and U1755 (N_1755,N_711,N_860);
or U1756 (N_1756,N_964,N_998);
and U1757 (N_1757,N_576,N_36);
and U1758 (N_1758,N_823,N_310);
or U1759 (N_1759,N_432,N_604);
nand U1760 (N_1760,N_407,N_85);
and U1761 (N_1761,N_205,N_162);
nor U1762 (N_1762,N_948,N_380);
or U1763 (N_1763,N_637,N_722);
xnor U1764 (N_1764,N_546,N_650);
nand U1765 (N_1765,N_637,N_195);
or U1766 (N_1766,N_367,N_129);
and U1767 (N_1767,N_728,N_708);
nor U1768 (N_1768,N_941,N_455);
nor U1769 (N_1769,N_150,N_534);
or U1770 (N_1770,N_685,N_293);
nor U1771 (N_1771,N_569,N_882);
nand U1772 (N_1772,N_104,N_938);
and U1773 (N_1773,N_373,N_317);
and U1774 (N_1774,N_382,N_41);
or U1775 (N_1775,N_842,N_588);
xor U1776 (N_1776,N_957,N_145);
nand U1777 (N_1777,N_444,N_755);
and U1778 (N_1778,N_82,N_16);
and U1779 (N_1779,N_962,N_183);
or U1780 (N_1780,N_864,N_455);
nand U1781 (N_1781,N_543,N_589);
and U1782 (N_1782,N_748,N_149);
xnor U1783 (N_1783,N_523,N_763);
or U1784 (N_1784,N_360,N_532);
or U1785 (N_1785,N_730,N_533);
nand U1786 (N_1786,N_91,N_309);
or U1787 (N_1787,N_65,N_682);
or U1788 (N_1788,N_241,N_75);
nor U1789 (N_1789,N_531,N_164);
nand U1790 (N_1790,N_283,N_13);
or U1791 (N_1791,N_266,N_276);
nor U1792 (N_1792,N_729,N_505);
nand U1793 (N_1793,N_799,N_529);
nor U1794 (N_1794,N_189,N_606);
nand U1795 (N_1795,N_851,N_481);
nand U1796 (N_1796,N_390,N_102);
xor U1797 (N_1797,N_276,N_143);
or U1798 (N_1798,N_163,N_281);
nor U1799 (N_1799,N_978,N_37);
xor U1800 (N_1800,N_797,N_97);
or U1801 (N_1801,N_105,N_67);
xor U1802 (N_1802,N_616,N_811);
nand U1803 (N_1803,N_745,N_122);
nand U1804 (N_1804,N_841,N_117);
nor U1805 (N_1805,N_982,N_199);
nand U1806 (N_1806,N_413,N_215);
xor U1807 (N_1807,N_916,N_749);
nand U1808 (N_1808,N_781,N_711);
xor U1809 (N_1809,N_104,N_387);
or U1810 (N_1810,N_221,N_357);
and U1811 (N_1811,N_589,N_591);
nor U1812 (N_1812,N_596,N_38);
and U1813 (N_1813,N_978,N_982);
and U1814 (N_1814,N_337,N_627);
nor U1815 (N_1815,N_649,N_869);
xnor U1816 (N_1816,N_27,N_247);
nor U1817 (N_1817,N_952,N_311);
nor U1818 (N_1818,N_974,N_160);
xor U1819 (N_1819,N_105,N_941);
xor U1820 (N_1820,N_140,N_538);
xor U1821 (N_1821,N_982,N_50);
or U1822 (N_1822,N_139,N_291);
nand U1823 (N_1823,N_544,N_396);
nand U1824 (N_1824,N_654,N_280);
or U1825 (N_1825,N_80,N_945);
xnor U1826 (N_1826,N_189,N_209);
nor U1827 (N_1827,N_360,N_807);
nor U1828 (N_1828,N_116,N_108);
xor U1829 (N_1829,N_239,N_63);
and U1830 (N_1830,N_96,N_960);
and U1831 (N_1831,N_648,N_743);
nand U1832 (N_1832,N_134,N_615);
or U1833 (N_1833,N_306,N_345);
nand U1834 (N_1834,N_776,N_118);
or U1835 (N_1835,N_422,N_211);
and U1836 (N_1836,N_585,N_529);
and U1837 (N_1837,N_291,N_728);
nor U1838 (N_1838,N_91,N_847);
or U1839 (N_1839,N_813,N_798);
xnor U1840 (N_1840,N_458,N_694);
xnor U1841 (N_1841,N_543,N_650);
nor U1842 (N_1842,N_435,N_204);
xnor U1843 (N_1843,N_840,N_529);
and U1844 (N_1844,N_400,N_340);
nand U1845 (N_1845,N_750,N_703);
nor U1846 (N_1846,N_107,N_937);
or U1847 (N_1847,N_327,N_278);
nor U1848 (N_1848,N_175,N_538);
xnor U1849 (N_1849,N_643,N_660);
or U1850 (N_1850,N_337,N_332);
xor U1851 (N_1851,N_41,N_428);
nor U1852 (N_1852,N_33,N_579);
and U1853 (N_1853,N_68,N_233);
nand U1854 (N_1854,N_247,N_716);
xnor U1855 (N_1855,N_441,N_31);
nand U1856 (N_1856,N_904,N_558);
and U1857 (N_1857,N_170,N_262);
nor U1858 (N_1858,N_449,N_471);
nor U1859 (N_1859,N_787,N_614);
nand U1860 (N_1860,N_333,N_99);
nor U1861 (N_1861,N_587,N_638);
nand U1862 (N_1862,N_500,N_565);
nor U1863 (N_1863,N_564,N_741);
nor U1864 (N_1864,N_996,N_552);
and U1865 (N_1865,N_60,N_216);
and U1866 (N_1866,N_960,N_359);
nor U1867 (N_1867,N_474,N_918);
and U1868 (N_1868,N_578,N_659);
or U1869 (N_1869,N_481,N_599);
xor U1870 (N_1870,N_61,N_277);
xnor U1871 (N_1871,N_370,N_17);
or U1872 (N_1872,N_615,N_471);
nand U1873 (N_1873,N_677,N_352);
xnor U1874 (N_1874,N_865,N_302);
nand U1875 (N_1875,N_872,N_7);
xnor U1876 (N_1876,N_744,N_748);
and U1877 (N_1877,N_666,N_424);
nor U1878 (N_1878,N_396,N_341);
or U1879 (N_1879,N_820,N_526);
nor U1880 (N_1880,N_711,N_796);
and U1881 (N_1881,N_397,N_707);
nor U1882 (N_1882,N_637,N_826);
nand U1883 (N_1883,N_875,N_975);
xnor U1884 (N_1884,N_8,N_384);
and U1885 (N_1885,N_158,N_607);
nand U1886 (N_1886,N_466,N_942);
nand U1887 (N_1887,N_828,N_660);
and U1888 (N_1888,N_351,N_923);
or U1889 (N_1889,N_818,N_402);
or U1890 (N_1890,N_326,N_331);
and U1891 (N_1891,N_372,N_245);
nand U1892 (N_1892,N_49,N_352);
xor U1893 (N_1893,N_569,N_103);
xor U1894 (N_1894,N_334,N_563);
nor U1895 (N_1895,N_177,N_504);
nand U1896 (N_1896,N_355,N_63);
xnor U1897 (N_1897,N_764,N_2);
or U1898 (N_1898,N_924,N_198);
and U1899 (N_1899,N_321,N_752);
nor U1900 (N_1900,N_796,N_810);
and U1901 (N_1901,N_874,N_967);
nand U1902 (N_1902,N_839,N_260);
nand U1903 (N_1903,N_540,N_743);
or U1904 (N_1904,N_589,N_516);
nor U1905 (N_1905,N_594,N_295);
nand U1906 (N_1906,N_195,N_756);
xor U1907 (N_1907,N_89,N_837);
xor U1908 (N_1908,N_216,N_696);
and U1909 (N_1909,N_373,N_293);
or U1910 (N_1910,N_758,N_254);
xnor U1911 (N_1911,N_278,N_415);
or U1912 (N_1912,N_867,N_905);
or U1913 (N_1913,N_373,N_492);
nand U1914 (N_1914,N_396,N_136);
nor U1915 (N_1915,N_676,N_621);
and U1916 (N_1916,N_785,N_899);
nand U1917 (N_1917,N_740,N_677);
xnor U1918 (N_1918,N_346,N_173);
and U1919 (N_1919,N_286,N_609);
xor U1920 (N_1920,N_479,N_288);
xnor U1921 (N_1921,N_327,N_365);
nand U1922 (N_1922,N_726,N_76);
xnor U1923 (N_1923,N_860,N_659);
nand U1924 (N_1924,N_750,N_865);
nor U1925 (N_1925,N_735,N_793);
nor U1926 (N_1926,N_776,N_250);
nor U1927 (N_1927,N_224,N_95);
nor U1928 (N_1928,N_726,N_235);
xor U1929 (N_1929,N_721,N_752);
nor U1930 (N_1930,N_906,N_65);
nand U1931 (N_1931,N_506,N_409);
and U1932 (N_1932,N_344,N_523);
nor U1933 (N_1933,N_867,N_541);
nand U1934 (N_1934,N_68,N_280);
and U1935 (N_1935,N_430,N_104);
nor U1936 (N_1936,N_104,N_401);
nor U1937 (N_1937,N_563,N_846);
nand U1938 (N_1938,N_866,N_761);
nor U1939 (N_1939,N_866,N_440);
or U1940 (N_1940,N_184,N_206);
xor U1941 (N_1941,N_326,N_38);
and U1942 (N_1942,N_899,N_810);
and U1943 (N_1943,N_940,N_63);
nand U1944 (N_1944,N_753,N_459);
xor U1945 (N_1945,N_812,N_572);
nand U1946 (N_1946,N_188,N_709);
and U1947 (N_1947,N_680,N_255);
and U1948 (N_1948,N_22,N_510);
xor U1949 (N_1949,N_964,N_913);
and U1950 (N_1950,N_185,N_570);
xor U1951 (N_1951,N_452,N_458);
nor U1952 (N_1952,N_440,N_11);
and U1953 (N_1953,N_372,N_145);
nor U1954 (N_1954,N_725,N_964);
or U1955 (N_1955,N_178,N_471);
and U1956 (N_1956,N_444,N_28);
nand U1957 (N_1957,N_267,N_588);
xor U1958 (N_1958,N_829,N_612);
and U1959 (N_1959,N_45,N_485);
nor U1960 (N_1960,N_466,N_490);
and U1961 (N_1961,N_147,N_567);
xnor U1962 (N_1962,N_490,N_814);
nor U1963 (N_1963,N_947,N_862);
nand U1964 (N_1964,N_780,N_599);
nand U1965 (N_1965,N_925,N_657);
and U1966 (N_1966,N_105,N_344);
xnor U1967 (N_1967,N_117,N_550);
xor U1968 (N_1968,N_442,N_599);
nand U1969 (N_1969,N_830,N_358);
nor U1970 (N_1970,N_199,N_254);
nand U1971 (N_1971,N_109,N_38);
xnor U1972 (N_1972,N_666,N_436);
and U1973 (N_1973,N_438,N_92);
nor U1974 (N_1974,N_581,N_60);
nand U1975 (N_1975,N_367,N_429);
nor U1976 (N_1976,N_199,N_656);
nor U1977 (N_1977,N_341,N_507);
nand U1978 (N_1978,N_577,N_256);
xnor U1979 (N_1979,N_721,N_219);
xor U1980 (N_1980,N_540,N_84);
and U1981 (N_1981,N_620,N_398);
xnor U1982 (N_1982,N_32,N_899);
and U1983 (N_1983,N_222,N_619);
nor U1984 (N_1984,N_252,N_960);
or U1985 (N_1985,N_130,N_650);
or U1986 (N_1986,N_599,N_637);
nor U1987 (N_1987,N_665,N_61);
nor U1988 (N_1988,N_383,N_920);
or U1989 (N_1989,N_709,N_818);
nor U1990 (N_1990,N_95,N_764);
nor U1991 (N_1991,N_468,N_509);
nand U1992 (N_1992,N_31,N_57);
xor U1993 (N_1993,N_714,N_101);
nand U1994 (N_1994,N_722,N_808);
and U1995 (N_1995,N_931,N_482);
and U1996 (N_1996,N_920,N_904);
nand U1997 (N_1997,N_587,N_100);
and U1998 (N_1998,N_643,N_392);
or U1999 (N_1999,N_461,N_652);
xor U2000 (N_2000,N_1445,N_1602);
or U2001 (N_2001,N_1978,N_1118);
nor U2002 (N_2002,N_1912,N_1960);
nor U2003 (N_2003,N_1254,N_1493);
nor U2004 (N_2004,N_1712,N_1982);
and U2005 (N_2005,N_1010,N_1657);
or U2006 (N_2006,N_1244,N_1084);
nand U2007 (N_2007,N_1317,N_1729);
nor U2008 (N_2008,N_1311,N_1298);
and U2009 (N_2009,N_1726,N_1742);
and U2010 (N_2010,N_1461,N_1324);
nor U2011 (N_2011,N_1603,N_1123);
nand U2012 (N_2012,N_1888,N_1651);
xor U2013 (N_2013,N_1971,N_1631);
and U2014 (N_2014,N_1815,N_1558);
and U2015 (N_2015,N_1228,N_1834);
nor U2016 (N_2016,N_1377,N_1235);
nor U2017 (N_2017,N_1135,N_1483);
nor U2018 (N_2018,N_1098,N_1580);
nor U2019 (N_2019,N_1386,N_1225);
xor U2020 (N_2020,N_1796,N_1753);
nand U2021 (N_2021,N_1586,N_1102);
or U2022 (N_2022,N_1464,N_1107);
xnor U2023 (N_2023,N_1266,N_1448);
xor U2024 (N_2024,N_1049,N_1820);
nand U2025 (N_2025,N_1261,N_1637);
or U2026 (N_2026,N_1111,N_1278);
or U2027 (N_2027,N_1406,N_1515);
xor U2028 (N_2028,N_1957,N_1976);
nand U2029 (N_2029,N_1552,N_1440);
nor U2030 (N_2030,N_1025,N_1808);
nand U2031 (N_2031,N_1650,N_1217);
and U2032 (N_2032,N_1824,N_1147);
xor U2033 (N_2033,N_1661,N_1142);
or U2034 (N_2034,N_1994,N_1466);
or U2035 (N_2035,N_1194,N_1294);
nand U2036 (N_2036,N_1260,N_1685);
or U2037 (N_2037,N_1703,N_1990);
nor U2038 (N_2038,N_1349,N_1148);
nor U2039 (N_2039,N_1851,N_1044);
nor U2040 (N_2040,N_1841,N_1314);
xnor U2041 (N_2041,N_1719,N_1418);
nand U2042 (N_2042,N_1594,N_1935);
nand U2043 (N_2043,N_1894,N_1436);
or U2044 (N_2044,N_1321,N_1562);
nand U2045 (N_2045,N_1042,N_1200);
nor U2046 (N_2046,N_1598,N_1926);
nor U2047 (N_2047,N_1832,N_1407);
nor U2048 (N_2048,N_1199,N_1573);
nor U2049 (N_2049,N_1197,N_1211);
or U2050 (N_2050,N_1277,N_1952);
and U2051 (N_2051,N_1114,N_1119);
or U2052 (N_2052,N_1420,N_1969);
nand U2053 (N_2053,N_1245,N_1860);
nor U2054 (N_2054,N_1563,N_1925);
or U2055 (N_2055,N_1901,N_1900);
or U2056 (N_2056,N_1996,N_1438);
or U2057 (N_2057,N_1943,N_1737);
and U2058 (N_2058,N_1604,N_1028);
xor U2059 (N_2059,N_1450,N_1307);
nor U2060 (N_2060,N_1739,N_1187);
nor U2061 (N_2061,N_1346,N_1053);
or U2062 (N_2062,N_1209,N_1747);
nor U2063 (N_2063,N_1539,N_1428);
nand U2064 (N_2064,N_1907,N_1046);
and U2065 (N_2065,N_1584,N_1267);
xor U2066 (N_2066,N_1588,N_1746);
xnor U2067 (N_2067,N_1587,N_1340);
and U2068 (N_2068,N_1125,N_1139);
and U2069 (N_2069,N_1919,N_1797);
nor U2070 (N_2070,N_1872,N_1621);
nand U2071 (N_2071,N_1763,N_1155);
xor U2072 (N_2072,N_1227,N_1845);
xor U2073 (N_2073,N_1662,N_1030);
or U2074 (N_2074,N_1082,N_1836);
or U2075 (N_2075,N_1501,N_1092);
nor U2076 (N_2076,N_1224,N_1761);
xor U2077 (N_2077,N_1078,N_1702);
or U2078 (N_2078,N_1259,N_1786);
or U2079 (N_2079,N_1776,N_1974);
nor U2080 (N_2080,N_1560,N_1096);
nor U2081 (N_2081,N_1095,N_1452);
nor U2082 (N_2082,N_1387,N_1575);
or U2083 (N_2083,N_1997,N_1048);
or U2084 (N_2084,N_1237,N_1451);
xor U2085 (N_2085,N_1565,N_1985);
or U2086 (N_2086,N_1358,N_1889);
and U2087 (N_2087,N_1429,N_1353);
xor U2088 (N_2088,N_1868,N_1853);
nor U2089 (N_2089,N_1667,N_1638);
and U2090 (N_2090,N_1998,N_1243);
nand U2091 (N_2091,N_1364,N_1833);
or U2092 (N_2092,N_1434,N_1972);
xnor U2093 (N_2093,N_1991,N_1034);
nand U2094 (N_2094,N_1906,N_1890);
and U2095 (N_2095,N_1714,N_1019);
nand U2096 (N_2096,N_1127,N_1809);
or U2097 (N_2097,N_1433,N_1457);
nand U2098 (N_2098,N_1492,N_1359);
or U2099 (N_2099,N_1936,N_1541);
and U2100 (N_2100,N_1517,N_1137);
xor U2101 (N_2101,N_1764,N_1910);
and U2102 (N_2102,N_1361,N_1380);
xor U2103 (N_2103,N_1213,N_1533);
nand U2104 (N_2104,N_1009,N_1649);
xnor U2105 (N_2105,N_1226,N_1474);
and U2106 (N_2106,N_1758,N_1374);
and U2107 (N_2107,N_1247,N_1124);
or U2108 (N_2108,N_1877,N_1556);
xnor U2109 (N_2109,N_1167,N_1686);
or U2110 (N_2110,N_1143,N_1619);
and U2111 (N_2111,N_1502,N_1818);
nor U2112 (N_2112,N_1400,N_1842);
and U2113 (N_2113,N_1837,N_1166);
or U2114 (N_2114,N_1027,N_1415);
nand U2115 (N_2115,N_1654,N_1617);
xor U2116 (N_2116,N_1191,N_1693);
or U2117 (N_2117,N_1695,N_1062);
or U2118 (N_2118,N_1465,N_1002);
or U2119 (N_2119,N_1937,N_1819);
nand U2120 (N_2120,N_1680,N_1876);
or U2121 (N_2121,N_1196,N_1599);
nand U2122 (N_2122,N_1987,N_1945);
and U2123 (N_2123,N_1850,N_1664);
nand U2124 (N_2124,N_1655,N_1402);
xnor U2125 (N_2125,N_1891,N_1543);
and U2126 (N_2126,N_1615,N_1516);
nor U2127 (N_2127,N_1767,N_1899);
nand U2128 (N_2128,N_1270,N_1723);
nor U2129 (N_2129,N_1146,N_1319);
xor U2130 (N_2130,N_1168,N_1572);
nor U2131 (N_2131,N_1134,N_1117);
nand U2132 (N_2132,N_1376,N_1787);
and U2133 (N_2133,N_1365,N_1472);
xnor U2134 (N_2134,N_1488,N_1626);
xnor U2135 (N_2135,N_1863,N_1838);
or U2136 (N_2136,N_1902,N_1172);
nor U2137 (N_2137,N_1977,N_1005);
or U2138 (N_2138,N_1692,N_1431);
xor U2139 (N_2139,N_1789,N_1162);
and U2140 (N_2140,N_1144,N_1547);
or U2141 (N_2141,N_1338,N_1866);
or U2142 (N_2142,N_1086,N_1810);
nand U2143 (N_2143,N_1857,N_1867);
xor U2144 (N_2144,N_1934,N_1373);
xnor U2145 (N_2145,N_1322,N_1339);
nor U2146 (N_2146,N_1458,N_1233);
or U2147 (N_2147,N_1839,N_1514);
xnor U2148 (N_2148,N_1091,N_1608);
nand U2149 (N_2149,N_1577,N_1555);
nand U2150 (N_2150,N_1807,N_1491);
xor U2151 (N_2151,N_1955,N_1333);
nand U2152 (N_2152,N_1766,N_1442);
or U2153 (N_2153,N_1660,N_1846);
xor U2154 (N_2154,N_1469,N_1616);
nand U2155 (N_2155,N_1684,N_1439);
nor U2156 (N_2156,N_1700,N_1885);
xor U2157 (N_2157,N_1554,N_1534);
or U2158 (N_2158,N_1828,N_1499);
xnor U2159 (N_2159,N_1736,N_1215);
or U2160 (N_2160,N_1051,N_1132);
xor U2161 (N_2161,N_1468,N_1455);
xor U2162 (N_2162,N_1579,N_1481);
nand U2163 (N_2163,N_1122,N_1592);
and U2164 (N_2164,N_1256,N_1363);
nand U2165 (N_2165,N_1881,N_1262);
nand U2166 (N_2166,N_1264,N_1487);
xnor U2167 (N_2167,N_1816,N_1675);
nor U2168 (N_2168,N_1967,N_1989);
xor U2169 (N_2169,N_1698,N_1120);
nor U2170 (N_2170,N_1065,N_1077);
nor U2171 (N_2171,N_1043,N_1152);
nor U2172 (N_2172,N_1255,N_1372);
xor U2173 (N_2173,N_1404,N_1540);
xnor U2174 (N_2174,N_1745,N_1980);
nor U2175 (N_2175,N_1559,N_1778);
or U2176 (N_2176,N_1825,N_1038);
xor U2177 (N_2177,N_1360,N_1323);
and U2178 (N_2178,N_1180,N_1506);
or U2179 (N_2179,N_1524,N_1727);
nand U2180 (N_2180,N_1318,N_1798);
and U2181 (N_2181,N_1236,N_1682);
or U2182 (N_2182,N_1896,N_1923);
nor U2183 (N_2183,N_1371,N_1368);
and U2184 (N_2184,N_1208,N_1652);
xnor U2185 (N_2185,N_1843,N_1751);
or U2186 (N_2186,N_1239,N_1183);
and U2187 (N_2187,N_1337,N_1207);
xor U2188 (N_2188,N_1417,N_1768);
xnor U2189 (N_2189,N_1014,N_1320);
nor U2190 (N_2190,N_1918,N_1403);
and U2191 (N_2191,N_1932,N_1003);
nor U2192 (N_2192,N_1733,N_1905);
nand U2193 (N_2193,N_1179,N_1668);
nand U2194 (N_2194,N_1342,N_1618);
and U2195 (N_2195,N_1823,N_1958);
and U2196 (N_2196,N_1496,N_1583);
or U2197 (N_2197,N_1192,N_1738);
nor U2198 (N_2198,N_1701,N_1503);
xnor U2199 (N_2199,N_1272,N_1110);
nor U2200 (N_2200,N_1198,N_1800);
or U2201 (N_2201,N_1128,N_1351);
nand U2202 (N_2202,N_1813,N_1663);
or U2203 (N_2203,N_1715,N_1308);
xor U2204 (N_2204,N_1874,N_1814);
nand U2205 (N_2205,N_1697,N_1462);
and U2206 (N_2206,N_1067,N_1538);
nor U2207 (N_2207,N_1916,N_1389);
xnor U2208 (N_2208,N_1486,N_1422);
nand U2209 (N_2209,N_1047,N_1671);
or U2210 (N_2210,N_1000,N_1007);
or U2211 (N_2211,N_1691,N_1313);
nand U2212 (N_2212,N_1748,N_1201);
nand U2213 (N_2213,N_1396,N_1567);
nor U2214 (N_2214,N_1665,N_1061);
nand U2215 (N_2215,N_1018,N_1467);
nand U2216 (N_2216,N_1206,N_1688);
nand U2217 (N_2217,N_1774,N_1614);
and U2218 (N_2218,N_1793,N_1520);
or U2219 (N_2219,N_1006,N_1391);
nor U2220 (N_2220,N_1382,N_1397);
and U2221 (N_2221,N_1770,N_1394);
nand U2222 (N_2222,N_1276,N_1505);
nor U2223 (N_2223,N_1419,N_1858);
and U2224 (N_2224,N_1108,N_1089);
xnor U2225 (N_2225,N_1893,N_1151);
xnor U2226 (N_2226,N_1634,N_1844);
and U2227 (N_2227,N_1510,N_1740);
nor U2228 (N_2228,N_1571,N_1523);
nand U2229 (N_2229,N_1717,N_1178);
or U2230 (N_2230,N_1306,N_1454);
or U2231 (N_2231,N_1345,N_1988);
and U2232 (N_2232,N_1498,N_1882);
xnor U2233 (N_2233,N_1069,N_1425);
or U2234 (N_2234,N_1287,N_1348);
xnor U2235 (N_2235,N_1694,N_1385);
nand U2236 (N_2236,N_1731,N_1141);
nand U2237 (N_2237,N_1444,N_1783);
nand U2238 (N_2238,N_1352,N_1105);
nor U2239 (N_2239,N_1286,N_1288);
xnor U2240 (N_2240,N_1924,N_1230);
or U2241 (N_2241,N_1606,N_1795);
xnor U2242 (N_2242,N_1384,N_1375);
and U2243 (N_2243,N_1759,N_1161);
nor U2244 (N_2244,N_1149,N_1303);
nand U2245 (N_2245,N_1922,N_1412);
and U2246 (N_2246,N_1975,N_1852);
and U2247 (N_2247,N_1821,N_1803);
nor U2248 (N_2248,N_1164,N_1170);
or U2249 (N_2249,N_1012,N_1920);
nor U2250 (N_2250,N_1903,N_1581);
nor U2251 (N_2251,N_1176,N_1656);
nor U2252 (N_2252,N_1341,N_1897);
and U2253 (N_2253,N_1589,N_1271);
nor U2254 (N_2254,N_1706,N_1551);
nand U2255 (N_2255,N_1100,N_1302);
or U2256 (N_2256,N_1252,N_1855);
and U2257 (N_2257,N_1116,N_1248);
nor U2258 (N_2258,N_1981,N_1772);
xnor U2259 (N_2259,N_1829,N_1627);
or U2260 (N_2260,N_1421,N_1268);
nand U2261 (N_2261,N_1312,N_1090);
xnor U2262 (N_2262,N_1184,N_1623);
nand U2263 (N_2263,N_1913,N_1635);
and U2264 (N_2264,N_1544,N_1521);
or U2265 (N_2265,N_1343,N_1231);
and U2266 (N_2266,N_1909,N_1275);
nor U2267 (N_2267,N_1249,N_1355);
or U2268 (N_2268,N_1639,N_1756);
and U2269 (N_2269,N_1140,N_1518);
or U2270 (N_2270,N_1522,N_1242);
nor U2271 (N_2271,N_1088,N_1273);
nand U2272 (N_2272,N_1914,N_1743);
or U2273 (N_2273,N_1849,N_1115);
and U2274 (N_2274,N_1917,N_1525);
xnor U2275 (N_2275,N_1395,N_1328);
or U2276 (N_2276,N_1050,N_1873);
or U2277 (N_2277,N_1332,N_1875);
and U2278 (N_2278,N_1113,N_1984);
nor U2279 (N_2279,N_1659,N_1036);
and U2280 (N_2280,N_1413,N_1630);
nor U2281 (N_2281,N_1250,N_1696);
nor U2282 (N_2282,N_1362,N_1218);
or U2283 (N_2283,N_1292,N_1204);
or U2284 (N_2284,N_1754,N_1032);
xnor U2285 (N_2285,N_1709,N_1079);
or U2286 (N_2286,N_1812,N_1773);
xnor U2287 (N_2287,N_1760,N_1173);
and U2288 (N_2288,N_1854,N_1946);
and U2289 (N_2289,N_1241,N_1781);
nand U2290 (N_2290,N_1950,N_1447);
and U2291 (N_2291,N_1840,N_1378);
or U2292 (N_2292,N_1802,N_1613);
nor U2293 (N_2293,N_1966,N_1093);
or U2294 (N_2294,N_1435,N_1281);
or U2295 (N_2295,N_1195,N_1512);
nor U2296 (N_2296,N_1785,N_1367);
nand U2297 (N_2297,N_1205,N_1951);
and U2298 (N_2298,N_1721,N_1182);
or U2299 (N_2299,N_1494,N_1379);
and U2300 (N_2300,N_1507,N_1653);
nand U2301 (N_2301,N_1713,N_1478);
xnor U2302 (N_2302,N_1532,N_1535);
and U2303 (N_2303,N_1528,N_1291);
nand U2304 (N_2304,N_1557,N_1104);
and U2305 (N_2305,N_1500,N_1174);
and U2306 (N_2306,N_1263,N_1865);
xor U2307 (N_2307,N_1274,N_1940);
nand U2308 (N_2308,N_1058,N_1459);
and U2309 (N_2309,N_1040,N_1536);
nor U2310 (N_2310,N_1234,N_1056);
xnor U2311 (N_2311,N_1707,N_1610);
nand U2312 (N_2312,N_1257,N_1405);
and U2313 (N_2313,N_1060,N_1762);
or U2314 (N_2314,N_1410,N_1732);
nor U2315 (N_2315,N_1674,N_1238);
or U2316 (N_2316,N_1177,N_1677);
xor U2317 (N_2317,N_1016,N_1189);
xnor U2318 (N_2318,N_1548,N_1513);
or U2319 (N_2319,N_1640,N_1424);
or U2320 (N_2320,N_1777,N_1826);
nor U2321 (N_2321,N_1026,N_1045);
or U2322 (N_2322,N_1453,N_1871);
nor U2323 (N_2323,N_1299,N_1961);
nor U2324 (N_2324,N_1370,N_1011);
nor U2325 (N_2325,N_1568,N_1181);
or U2326 (N_2326,N_1601,N_1130);
or U2327 (N_2327,N_1670,N_1642);
and U2328 (N_2328,N_1862,N_1861);
nand U2329 (N_2329,N_1750,N_1771);
nand U2330 (N_2330,N_1356,N_1013);
nand U2331 (N_2331,N_1327,N_1432);
and U2332 (N_2332,N_1280,N_1390);
nor U2333 (N_2333,N_1956,N_1310);
or U2334 (N_2334,N_1632,N_1574);
or U2335 (N_2335,N_1411,N_1979);
xnor U2336 (N_2336,N_1553,N_1335);
xnor U2337 (N_2337,N_1791,N_1220);
or U2338 (N_2338,N_1460,N_1546);
nor U2339 (N_2339,N_1171,N_1041);
or U2340 (N_2340,N_1154,N_1190);
xor U2341 (N_2341,N_1441,N_1835);
xnor U2342 (N_2342,N_1409,N_1811);
xor U2343 (N_2343,N_1904,N_1301);
nand U2344 (N_2344,N_1549,N_1780);
nor U2345 (N_2345,N_1145,N_1624);
and U2346 (N_2346,N_1993,N_1720);
nand U2347 (N_2347,N_1954,N_1806);
and U2348 (N_2348,N_1175,N_1024);
nand U2349 (N_2349,N_1326,N_1157);
or U2350 (N_2350,N_1392,N_1689);
and U2351 (N_2351,N_1704,N_1730);
and U2352 (N_2352,N_1511,N_1240);
nor U2353 (N_2353,N_1929,N_1962);
nand U2354 (N_2354,N_1887,N_1063);
nand U2355 (N_2355,N_1672,N_1232);
and U2356 (N_2356,N_1509,N_1057);
or U2357 (N_2357,N_1071,N_1325);
xor U2358 (N_2358,N_1138,N_1879);
nand U2359 (N_2359,N_1004,N_1269);
nor U2360 (N_2360,N_1463,N_1734);
nor U2361 (N_2361,N_1039,N_1210);
nor U2362 (N_2362,N_1073,N_1953);
or U2363 (N_2363,N_1446,N_1947);
or U2364 (N_2364,N_1537,N_1595);
xor U2365 (N_2365,N_1790,N_1831);
xnor U2366 (N_2366,N_1265,N_1775);
or U2367 (N_2367,N_1188,N_1643);
xnor U2368 (N_2368,N_1576,N_1633);
nand U2369 (N_2369,N_1297,N_1927);
and U2370 (N_2370,N_1895,N_1289);
and U2371 (N_2371,N_1636,N_1430);
nand U2372 (N_2372,N_1366,N_1316);
xnor U2373 (N_2373,N_1059,N_1066);
nor U2374 (N_2374,N_1859,N_1864);
xor U2375 (N_2375,N_1687,N_1443);
and U2376 (N_2376,N_1126,N_1593);
or U2377 (N_2377,N_1473,N_1054);
and U2378 (N_2378,N_1504,N_1490);
xor U2379 (N_2379,N_1471,N_1037);
and U2380 (N_2380,N_1129,N_1221);
and U2381 (N_2381,N_1545,N_1497);
and U2382 (N_2382,N_1611,N_1561);
nand U2383 (N_2383,N_1344,N_1699);
and U2384 (N_2384,N_1749,N_1258);
xnor U2385 (N_2385,N_1892,N_1622);
and U2386 (N_2386,N_1035,N_1992);
and U2387 (N_2387,N_1015,N_1995);
nand U2388 (N_2388,N_1112,N_1570);
nor U2389 (N_2389,N_1085,N_1068);
and U2390 (N_2390,N_1856,N_1334);
or U2391 (N_2391,N_1099,N_1527);
nor U2392 (N_2392,N_1489,N_1931);
nor U2393 (N_2393,N_1109,N_1566);
nor U2394 (N_2394,N_1884,N_1282);
nor U2395 (N_2395,N_1414,N_1799);
xnor U2396 (N_2396,N_1804,N_1792);
xnor U2397 (N_2397,N_1679,N_1757);
nor U2398 (N_2398,N_1354,N_1283);
and U2399 (N_2399,N_1883,N_1304);
xnor U2400 (N_2400,N_1519,N_1596);
and U2401 (N_2401,N_1647,N_1970);
or U2402 (N_2402,N_1531,N_1315);
or U2403 (N_2403,N_1564,N_1898);
nor U2404 (N_2404,N_1886,N_1075);
nand U2405 (N_2405,N_1437,N_1331);
and U2406 (N_2406,N_1628,N_1309);
nor U2407 (N_2407,N_1949,N_1765);
xor U2408 (N_2408,N_1641,N_1716);
nand U2409 (N_2409,N_1484,N_1648);
or U2410 (N_2410,N_1133,N_1336);
nor U2411 (N_2411,N_1094,N_1165);
nand U2412 (N_2412,N_1293,N_1725);
and U2413 (N_2413,N_1921,N_1064);
nand U2414 (N_2414,N_1399,N_1482);
nand U2415 (N_2415,N_1550,N_1782);
or U2416 (N_2416,N_1156,N_1582);
nand U2417 (N_2417,N_1784,N_1222);
nor U2418 (N_2418,N_1470,N_1087);
xor U2419 (N_2419,N_1973,N_1880);
nand U2420 (N_2420,N_1052,N_1296);
or U2421 (N_2421,N_1718,N_1159);
or U2422 (N_2422,N_1081,N_1681);
nand U2423 (N_2423,N_1690,N_1017);
xnor U2424 (N_2424,N_1542,N_1944);
nor U2425 (N_2425,N_1008,N_1216);
or U2426 (N_2426,N_1948,N_1708);
xor U2427 (N_2427,N_1103,N_1569);
xor U2428 (N_2428,N_1878,N_1001);
or U2429 (N_2429,N_1965,N_1822);
nand U2430 (N_2430,N_1076,N_1449);
and U2431 (N_2431,N_1620,N_1644);
xnor U2432 (N_2432,N_1908,N_1711);
nor U2433 (N_2433,N_1938,N_1959);
and U2434 (N_2434,N_1928,N_1666);
or U2435 (N_2435,N_1279,N_1160);
nand U2436 (N_2436,N_1020,N_1131);
xor U2437 (N_2437,N_1401,N_1031);
xor U2438 (N_2438,N_1607,N_1476);
xor U2439 (N_2439,N_1529,N_1968);
or U2440 (N_2440,N_1097,N_1830);
xnor U2441 (N_2441,N_1485,N_1769);
xnor U2442 (N_2442,N_1609,N_1915);
nand U2443 (N_2443,N_1941,N_1741);
xor U2444 (N_2444,N_1779,N_1383);
xnor U2445 (N_2445,N_1848,N_1408);
and U2446 (N_2446,N_1805,N_1369);
xnor U2447 (N_2447,N_1070,N_1223);
nor U2448 (N_2448,N_1590,N_1597);
nand U2449 (N_2449,N_1074,N_1285);
nor U2450 (N_2450,N_1163,N_1153);
or U2451 (N_2451,N_1456,N_1827);
nor U2452 (N_2452,N_1801,N_1933);
xnor U2453 (N_2453,N_1479,N_1755);
xor U2454 (N_2454,N_1600,N_1710);
xor U2455 (N_2455,N_1752,N_1794);
xnor U2456 (N_2456,N_1305,N_1029);
or U2457 (N_2457,N_1253,N_1999);
xnor U2458 (N_2458,N_1388,N_1629);
or U2459 (N_2459,N_1246,N_1347);
nand U2460 (N_2460,N_1083,N_1393);
nor U2461 (N_2461,N_1625,N_1229);
and U2462 (N_2462,N_1022,N_1416);
nor U2463 (N_2463,N_1423,N_1939);
or U2464 (N_2464,N_1072,N_1475);
nand U2465 (N_2465,N_1330,N_1673);
nand U2466 (N_2466,N_1645,N_1724);
or U2467 (N_2467,N_1023,N_1219);
xnor U2468 (N_2468,N_1300,N_1963);
nor U2469 (N_2469,N_1295,N_1203);
nand U2470 (N_2470,N_1983,N_1185);
and U2471 (N_2471,N_1136,N_1678);
nor U2472 (N_2472,N_1847,N_1158);
xnor U2473 (N_2473,N_1251,N_1193);
and U2474 (N_2474,N_1676,N_1477);
xor U2475 (N_2475,N_1585,N_1986);
nand U2476 (N_2476,N_1121,N_1930);
nor U2477 (N_2477,N_1817,N_1669);
nand U2478 (N_2478,N_1202,N_1728);
nand U2479 (N_2479,N_1683,N_1055);
nand U2480 (N_2480,N_1788,N_1530);
or U2481 (N_2481,N_1033,N_1869);
xor U2482 (N_2482,N_1646,N_1605);
xor U2483 (N_2483,N_1744,N_1284);
and U2484 (N_2484,N_1578,N_1480);
and U2485 (N_2485,N_1508,N_1212);
and U2486 (N_2486,N_1021,N_1357);
xnor U2487 (N_2487,N_1722,N_1350);
nand U2488 (N_2488,N_1427,N_1381);
or U2489 (N_2489,N_1290,N_1398);
and U2490 (N_2490,N_1426,N_1106);
nor U2491 (N_2491,N_1942,N_1214);
xor U2492 (N_2492,N_1101,N_1169);
and U2493 (N_2493,N_1870,N_1964);
or U2494 (N_2494,N_1080,N_1658);
nand U2495 (N_2495,N_1150,N_1735);
xor U2496 (N_2496,N_1612,N_1911);
and U2497 (N_2497,N_1186,N_1591);
xor U2498 (N_2498,N_1495,N_1526);
nand U2499 (N_2499,N_1705,N_1329);
and U2500 (N_2500,N_1533,N_1318);
xor U2501 (N_2501,N_1291,N_1581);
nand U2502 (N_2502,N_1117,N_1482);
or U2503 (N_2503,N_1977,N_1315);
nand U2504 (N_2504,N_1892,N_1828);
or U2505 (N_2505,N_1927,N_1872);
nor U2506 (N_2506,N_1227,N_1797);
or U2507 (N_2507,N_1162,N_1400);
or U2508 (N_2508,N_1778,N_1084);
or U2509 (N_2509,N_1345,N_1584);
nand U2510 (N_2510,N_1409,N_1273);
nand U2511 (N_2511,N_1730,N_1727);
or U2512 (N_2512,N_1489,N_1289);
and U2513 (N_2513,N_1722,N_1747);
and U2514 (N_2514,N_1296,N_1608);
or U2515 (N_2515,N_1742,N_1527);
or U2516 (N_2516,N_1559,N_1867);
xnor U2517 (N_2517,N_1200,N_1488);
and U2518 (N_2518,N_1412,N_1388);
nor U2519 (N_2519,N_1366,N_1009);
and U2520 (N_2520,N_1086,N_1212);
and U2521 (N_2521,N_1836,N_1036);
nand U2522 (N_2522,N_1828,N_1135);
xnor U2523 (N_2523,N_1034,N_1866);
xnor U2524 (N_2524,N_1757,N_1739);
xnor U2525 (N_2525,N_1156,N_1231);
nand U2526 (N_2526,N_1201,N_1337);
xor U2527 (N_2527,N_1519,N_1116);
or U2528 (N_2528,N_1198,N_1326);
nand U2529 (N_2529,N_1093,N_1320);
or U2530 (N_2530,N_1897,N_1165);
xnor U2531 (N_2531,N_1315,N_1206);
and U2532 (N_2532,N_1583,N_1460);
or U2533 (N_2533,N_1821,N_1839);
or U2534 (N_2534,N_1240,N_1039);
and U2535 (N_2535,N_1050,N_1955);
xnor U2536 (N_2536,N_1622,N_1534);
or U2537 (N_2537,N_1003,N_1179);
and U2538 (N_2538,N_1490,N_1347);
nor U2539 (N_2539,N_1442,N_1123);
xnor U2540 (N_2540,N_1645,N_1731);
nor U2541 (N_2541,N_1672,N_1434);
nand U2542 (N_2542,N_1243,N_1480);
nand U2543 (N_2543,N_1973,N_1252);
xnor U2544 (N_2544,N_1429,N_1335);
and U2545 (N_2545,N_1861,N_1841);
nor U2546 (N_2546,N_1957,N_1040);
nor U2547 (N_2547,N_1599,N_1247);
nor U2548 (N_2548,N_1361,N_1830);
nor U2549 (N_2549,N_1123,N_1081);
and U2550 (N_2550,N_1107,N_1741);
or U2551 (N_2551,N_1199,N_1635);
nor U2552 (N_2552,N_1875,N_1552);
or U2553 (N_2553,N_1457,N_1142);
or U2554 (N_2554,N_1770,N_1116);
nand U2555 (N_2555,N_1171,N_1304);
nor U2556 (N_2556,N_1752,N_1193);
nand U2557 (N_2557,N_1894,N_1870);
and U2558 (N_2558,N_1911,N_1225);
nand U2559 (N_2559,N_1739,N_1307);
nand U2560 (N_2560,N_1610,N_1655);
xnor U2561 (N_2561,N_1447,N_1500);
nor U2562 (N_2562,N_1427,N_1527);
and U2563 (N_2563,N_1956,N_1160);
or U2564 (N_2564,N_1035,N_1469);
nand U2565 (N_2565,N_1784,N_1712);
or U2566 (N_2566,N_1884,N_1062);
or U2567 (N_2567,N_1568,N_1787);
nor U2568 (N_2568,N_1200,N_1132);
nor U2569 (N_2569,N_1632,N_1289);
xor U2570 (N_2570,N_1294,N_1805);
or U2571 (N_2571,N_1277,N_1127);
nand U2572 (N_2572,N_1563,N_1955);
and U2573 (N_2573,N_1532,N_1480);
and U2574 (N_2574,N_1982,N_1587);
and U2575 (N_2575,N_1971,N_1707);
nor U2576 (N_2576,N_1404,N_1467);
xnor U2577 (N_2577,N_1898,N_1689);
nand U2578 (N_2578,N_1739,N_1501);
nand U2579 (N_2579,N_1566,N_1994);
nand U2580 (N_2580,N_1050,N_1018);
xor U2581 (N_2581,N_1007,N_1804);
nand U2582 (N_2582,N_1234,N_1899);
xnor U2583 (N_2583,N_1416,N_1850);
xor U2584 (N_2584,N_1167,N_1612);
nor U2585 (N_2585,N_1155,N_1554);
nor U2586 (N_2586,N_1579,N_1417);
or U2587 (N_2587,N_1381,N_1274);
nand U2588 (N_2588,N_1893,N_1747);
nor U2589 (N_2589,N_1254,N_1068);
and U2590 (N_2590,N_1809,N_1719);
xnor U2591 (N_2591,N_1818,N_1624);
xor U2592 (N_2592,N_1883,N_1786);
nor U2593 (N_2593,N_1385,N_1479);
and U2594 (N_2594,N_1822,N_1674);
nand U2595 (N_2595,N_1563,N_1131);
xor U2596 (N_2596,N_1521,N_1025);
nand U2597 (N_2597,N_1280,N_1780);
and U2598 (N_2598,N_1091,N_1913);
or U2599 (N_2599,N_1079,N_1375);
nor U2600 (N_2600,N_1363,N_1725);
xnor U2601 (N_2601,N_1708,N_1594);
or U2602 (N_2602,N_1833,N_1629);
nand U2603 (N_2603,N_1117,N_1886);
nor U2604 (N_2604,N_1633,N_1861);
nor U2605 (N_2605,N_1002,N_1592);
and U2606 (N_2606,N_1850,N_1066);
nor U2607 (N_2607,N_1072,N_1192);
xnor U2608 (N_2608,N_1848,N_1628);
nand U2609 (N_2609,N_1187,N_1970);
or U2610 (N_2610,N_1747,N_1101);
or U2611 (N_2611,N_1007,N_1384);
xor U2612 (N_2612,N_1948,N_1896);
or U2613 (N_2613,N_1250,N_1381);
and U2614 (N_2614,N_1524,N_1800);
or U2615 (N_2615,N_1152,N_1850);
xnor U2616 (N_2616,N_1776,N_1419);
and U2617 (N_2617,N_1229,N_1332);
xor U2618 (N_2618,N_1419,N_1411);
nor U2619 (N_2619,N_1086,N_1242);
nand U2620 (N_2620,N_1632,N_1765);
or U2621 (N_2621,N_1535,N_1187);
nor U2622 (N_2622,N_1799,N_1090);
and U2623 (N_2623,N_1345,N_1454);
and U2624 (N_2624,N_1659,N_1232);
xnor U2625 (N_2625,N_1679,N_1423);
nor U2626 (N_2626,N_1079,N_1403);
or U2627 (N_2627,N_1268,N_1533);
or U2628 (N_2628,N_1382,N_1396);
nand U2629 (N_2629,N_1118,N_1657);
and U2630 (N_2630,N_1492,N_1526);
xnor U2631 (N_2631,N_1315,N_1754);
nor U2632 (N_2632,N_1997,N_1105);
nand U2633 (N_2633,N_1772,N_1009);
xor U2634 (N_2634,N_1567,N_1316);
nand U2635 (N_2635,N_1297,N_1620);
nand U2636 (N_2636,N_1183,N_1040);
or U2637 (N_2637,N_1290,N_1499);
xor U2638 (N_2638,N_1273,N_1098);
and U2639 (N_2639,N_1530,N_1431);
xnor U2640 (N_2640,N_1156,N_1203);
xor U2641 (N_2641,N_1161,N_1087);
and U2642 (N_2642,N_1075,N_1997);
xnor U2643 (N_2643,N_1391,N_1458);
nand U2644 (N_2644,N_1810,N_1222);
or U2645 (N_2645,N_1721,N_1961);
and U2646 (N_2646,N_1016,N_1600);
nand U2647 (N_2647,N_1284,N_1706);
or U2648 (N_2648,N_1792,N_1756);
xor U2649 (N_2649,N_1433,N_1546);
nor U2650 (N_2650,N_1755,N_1928);
nor U2651 (N_2651,N_1749,N_1939);
xnor U2652 (N_2652,N_1987,N_1077);
nor U2653 (N_2653,N_1291,N_1719);
or U2654 (N_2654,N_1814,N_1742);
nand U2655 (N_2655,N_1400,N_1979);
nor U2656 (N_2656,N_1802,N_1395);
and U2657 (N_2657,N_1250,N_1574);
nand U2658 (N_2658,N_1296,N_1076);
nand U2659 (N_2659,N_1852,N_1608);
xor U2660 (N_2660,N_1282,N_1777);
and U2661 (N_2661,N_1280,N_1964);
xnor U2662 (N_2662,N_1568,N_1191);
xnor U2663 (N_2663,N_1894,N_1497);
nand U2664 (N_2664,N_1960,N_1518);
and U2665 (N_2665,N_1587,N_1392);
xor U2666 (N_2666,N_1204,N_1536);
xnor U2667 (N_2667,N_1767,N_1375);
or U2668 (N_2668,N_1837,N_1377);
and U2669 (N_2669,N_1187,N_1794);
xor U2670 (N_2670,N_1752,N_1557);
nor U2671 (N_2671,N_1803,N_1555);
or U2672 (N_2672,N_1326,N_1855);
nand U2673 (N_2673,N_1299,N_1475);
nor U2674 (N_2674,N_1980,N_1729);
and U2675 (N_2675,N_1579,N_1623);
and U2676 (N_2676,N_1292,N_1762);
or U2677 (N_2677,N_1068,N_1551);
and U2678 (N_2678,N_1821,N_1746);
xnor U2679 (N_2679,N_1623,N_1198);
or U2680 (N_2680,N_1060,N_1739);
and U2681 (N_2681,N_1190,N_1111);
and U2682 (N_2682,N_1414,N_1374);
nor U2683 (N_2683,N_1342,N_1468);
nor U2684 (N_2684,N_1546,N_1606);
or U2685 (N_2685,N_1635,N_1511);
and U2686 (N_2686,N_1934,N_1720);
nand U2687 (N_2687,N_1752,N_1551);
nor U2688 (N_2688,N_1131,N_1975);
nand U2689 (N_2689,N_1994,N_1118);
and U2690 (N_2690,N_1548,N_1482);
xnor U2691 (N_2691,N_1992,N_1367);
and U2692 (N_2692,N_1418,N_1425);
nor U2693 (N_2693,N_1899,N_1645);
or U2694 (N_2694,N_1851,N_1013);
or U2695 (N_2695,N_1735,N_1520);
or U2696 (N_2696,N_1219,N_1631);
and U2697 (N_2697,N_1426,N_1472);
and U2698 (N_2698,N_1257,N_1813);
nor U2699 (N_2699,N_1495,N_1793);
nand U2700 (N_2700,N_1778,N_1942);
or U2701 (N_2701,N_1720,N_1778);
and U2702 (N_2702,N_1239,N_1189);
nand U2703 (N_2703,N_1681,N_1543);
xnor U2704 (N_2704,N_1628,N_1860);
or U2705 (N_2705,N_1634,N_1135);
nor U2706 (N_2706,N_1401,N_1109);
nor U2707 (N_2707,N_1939,N_1990);
nand U2708 (N_2708,N_1337,N_1977);
xnor U2709 (N_2709,N_1581,N_1507);
nor U2710 (N_2710,N_1530,N_1089);
nand U2711 (N_2711,N_1141,N_1636);
nor U2712 (N_2712,N_1384,N_1668);
xor U2713 (N_2713,N_1190,N_1899);
nand U2714 (N_2714,N_1505,N_1523);
nor U2715 (N_2715,N_1760,N_1411);
and U2716 (N_2716,N_1973,N_1863);
and U2717 (N_2717,N_1482,N_1924);
and U2718 (N_2718,N_1619,N_1972);
and U2719 (N_2719,N_1139,N_1447);
xnor U2720 (N_2720,N_1296,N_1952);
and U2721 (N_2721,N_1188,N_1488);
or U2722 (N_2722,N_1854,N_1667);
and U2723 (N_2723,N_1664,N_1597);
nor U2724 (N_2724,N_1579,N_1603);
xor U2725 (N_2725,N_1056,N_1507);
xnor U2726 (N_2726,N_1818,N_1724);
nand U2727 (N_2727,N_1862,N_1461);
nor U2728 (N_2728,N_1483,N_1826);
nand U2729 (N_2729,N_1491,N_1913);
and U2730 (N_2730,N_1645,N_1046);
nor U2731 (N_2731,N_1415,N_1447);
xor U2732 (N_2732,N_1182,N_1245);
xor U2733 (N_2733,N_1384,N_1984);
and U2734 (N_2734,N_1185,N_1826);
xnor U2735 (N_2735,N_1272,N_1966);
and U2736 (N_2736,N_1797,N_1286);
nor U2737 (N_2737,N_1815,N_1025);
nand U2738 (N_2738,N_1560,N_1677);
nor U2739 (N_2739,N_1760,N_1825);
and U2740 (N_2740,N_1558,N_1298);
nand U2741 (N_2741,N_1163,N_1100);
nand U2742 (N_2742,N_1751,N_1584);
or U2743 (N_2743,N_1912,N_1525);
or U2744 (N_2744,N_1514,N_1120);
and U2745 (N_2745,N_1076,N_1657);
or U2746 (N_2746,N_1239,N_1462);
or U2747 (N_2747,N_1391,N_1127);
xor U2748 (N_2748,N_1266,N_1658);
or U2749 (N_2749,N_1378,N_1207);
nor U2750 (N_2750,N_1483,N_1122);
nor U2751 (N_2751,N_1794,N_1733);
xnor U2752 (N_2752,N_1980,N_1081);
xnor U2753 (N_2753,N_1874,N_1234);
nand U2754 (N_2754,N_1831,N_1231);
xor U2755 (N_2755,N_1065,N_1638);
xor U2756 (N_2756,N_1340,N_1611);
xnor U2757 (N_2757,N_1748,N_1875);
xnor U2758 (N_2758,N_1699,N_1777);
nand U2759 (N_2759,N_1575,N_1868);
nand U2760 (N_2760,N_1773,N_1018);
nor U2761 (N_2761,N_1856,N_1008);
or U2762 (N_2762,N_1565,N_1937);
or U2763 (N_2763,N_1646,N_1597);
or U2764 (N_2764,N_1905,N_1324);
nor U2765 (N_2765,N_1659,N_1761);
nor U2766 (N_2766,N_1635,N_1503);
xor U2767 (N_2767,N_1065,N_1434);
nand U2768 (N_2768,N_1983,N_1420);
or U2769 (N_2769,N_1096,N_1111);
nand U2770 (N_2770,N_1285,N_1020);
or U2771 (N_2771,N_1631,N_1211);
and U2772 (N_2772,N_1313,N_1509);
nand U2773 (N_2773,N_1684,N_1881);
and U2774 (N_2774,N_1016,N_1640);
nor U2775 (N_2775,N_1932,N_1482);
or U2776 (N_2776,N_1751,N_1079);
xnor U2777 (N_2777,N_1334,N_1428);
and U2778 (N_2778,N_1373,N_1509);
nand U2779 (N_2779,N_1696,N_1393);
nand U2780 (N_2780,N_1864,N_1356);
or U2781 (N_2781,N_1601,N_1991);
and U2782 (N_2782,N_1681,N_1670);
nor U2783 (N_2783,N_1616,N_1676);
or U2784 (N_2784,N_1913,N_1976);
and U2785 (N_2785,N_1348,N_1711);
nor U2786 (N_2786,N_1188,N_1015);
nand U2787 (N_2787,N_1719,N_1507);
and U2788 (N_2788,N_1037,N_1330);
and U2789 (N_2789,N_1891,N_1763);
nor U2790 (N_2790,N_1769,N_1463);
nor U2791 (N_2791,N_1574,N_1646);
nand U2792 (N_2792,N_1406,N_1771);
nand U2793 (N_2793,N_1406,N_1871);
or U2794 (N_2794,N_1581,N_1306);
or U2795 (N_2795,N_1064,N_1248);
and U2796 (N_2796,N_1086,N_1259);
or U2797 (N_2797,N_1549,N_1362);
nand U2798 (N_2798,N_1095,N_1469);
xor U2799 (N_2799,N_1252,N_1391);
nand U2800 (N_2800,N_1618,N_1875);
xnor U2801 (N_2801,N_1440,N_1641);
xor U2802 (N_2802,N_1471,N_1445);
nor U2803 (N_2803,N_1383,N_1170);
xnor U2804 (N_2804,N_1494,N_1885);
and U2805 (N_2805,N_1509,N_1075);
nor U2806 (N_2806,N_1075,N_1147);
or U2807 (N_2807,N_1886,N_1709);
xnor U2808 (N_2808,N_1416,N_1880);
nor U2809 (N_2809,N_1228,N_1087);
nor U2810 (N_2810,N_1153,N_1473);
nand U2811 (N_2811,N_1310,N_1224);
or U2812 (N_2812,N_1801,N_1851);
xor U2813 (N_2813,N_1166,N_1622);
and U2814 (N_2814,N_1809,N_1844);
xor U2815 (N_2815,N_1746,N_1159);
nand U2816 (N_2816,N_1404,N_1511);
nand U2817 (N_2817,N_1593,N_1308);
xor U2818 (N_2818,N_1369,N_1158);
xnor U2819 (N_2819,N_1396,N_1443);
or U2820 (N_2820,N_1493,N_1367);
xor U2821 (N_2821,N_1043,N_1462);
or U2822 (N_2822,N_1935,N_1129);
and U2823 (N_2823,N_1853,N_1843);
nor U2824 (N_2824,N_1292,N_1138);
nand U2825 (N_2825,N_1525,N_1725);
nor U2826 (N_2826,N_1635,N_1844);
or U2827 (N_2827,N_1755,N_1540);
xnor U2828 (N_2828,N_1200,N_1209);
nand U2829 (N_2829,N_1796,N_1952);
xnor U2830 (N_2830,N_1164,N_1607);
xor U2831 (N_2831,N_1765,N_1851);
nand U2832 (N_2832,N_1119,N_1925);
and U2833 (N_2833,N_1285,N_1467);
xor U2834 (N_2834,N_1669,N_1527);
and U2835 (N_2835,N_1766,N_1571);
and U2836 (N_2836,N_1102,N_1983);
nand U2837 (N_2837,N_1290,N_1148);
or U2838 (N_2838,N_1785,N_1934);
xnor U2839 (N_2839,N_1403,N_1954);
nor U2840 (N_2840,N_1764,N_1178);
nor U2841 (N_2841,N_1931,N_1033);
and U2842 (N_2842,N_1016,N_1368);
or U2843 (N_2843,N_1930,N_1310);
nor U2844 (N_2844,N_1174,N_1849);
and U2845 (N_2845,N_1614,N_1317);
nor U2846 (N_2846,N_1585,N_1288);
xor U2847 (N_2847,N_1499,N_1442);
nand U2848 (N_2848,N_1254,N_1960);
xor U2849 (N_2849,N_1449,N_1424);
nand U2850 (N_2850,N_1491,N_1978);
and U2851 (N_2851,N_1010,N_1661);
or U2852 (N_2852,N_1333,N_1012);
xnor U2853 (N_2853,N_1260,N_1494);
nand U2854 (N_2854,N_1032,N_1373);
xor U2855 (N_2855,N_1484,N_1915);
and U2856 (N_2856,N_1761,N_1371);
xnor U2857 (N_2857,N_1669,N_1034);
xor U2858 (N_2858,N_1004,N_1091);
xnor U2859 (N_2859,N_1750,N_1575);
or U2860 (N_2860,N_1683,N_1404);
or U2861 (N_2861,N_1136,N_1443);
or U2862 (N_2862,N_1428,N_1642);
xor U2863 (N_2863,N_1324,N_1912);
nor U2864 (N_2864,N_1309,N_1806);
nor U2865 (N_2865,N_1884,N_1412);
or U2866 (N_2866,N_1965,N_1923);
xnor U2867 (N_2867,N_1080,N_1466);
and U2868 (N_2868,N_1637,N_1447);
xor U2869 (N_2869,N_1900,N_1154);
and U2870 (N_2870,N_1427,N_1685);
nor U2871 (N_2871,N_1556,N_1462);
nand U2872 (N_2872,N_1916,N_1997);
and U2873 (N_2873,N_1248,N_1135);
nor U2874 (N_2874,N_1541,N_1833);
or U2875 (N_2875,N_1664,N_1053);
xnor U2876 (N_2876,N_1573,N_1267);
or U2877 (N_2877,N_1015,N_1737);
or U2878 (N_2878,N_1797,N_1668);
and U2879 (N_2879,N_1276,N_1751);
and U2880 (N_2880,N_1959,N_1212);
xor U2881 (N_2881,N_1835,N_1665);
and U2882 (N_2882,N_1669,N_1283);
xor U2883 (N_2883,N_1955,N_1895);
xnor U2884 (N_2884,N_1292,N_1328);
nand U2885 (N_2885,N_1727,N_1684);
xnor U2886 (N_2886,N_1365,N_1979);
and U2887 (N_2887,N_1325,N_1090);
nor U2888 (N_2888,N_1105,N_1675);
and U2889 (N_2889,N_1666,N_1250);
or U2890 (N_2890,N_1217,N_1605);
nand U2891 (N_2891,N_1010,N_1272);
nand U2892 (N_2892,N_1929,N_1417);
or U2893 (N_2893,N_1750,N_1306);
nand U2894 (N_2894,N_1672,N_1836);
nor U2895 (N_2895,N_1877,N_1141);
and U2896 (N_2896,N_1975,N_1783);
xor U2897 (N_2897,N_1480,N_1617);
or U2898 (N_2898,N_1781,N_1949);
nor U2899 (N_2899,N_1828,N_1750);
xor U2900 (N_2900,N_1915,N_1287);
nor U2901 (N_2901,N_1219,N_1227);
xnor U2902 (N_2902,N_1102,N_1897);
and U2903 (N_2903,N_1423,N_1513);
nand U2904 (N_2904,N_1404,N_1178);
nor U2905 (N_2905,N_1738,N_1680);
or U2906 (N_2906,N_1432,N_1464);
xnor U2907 (N_2907,N_1742,N_1885);
or U2908 (N_2908,N_1702,N_1328);
or U2909 (N_2909,N_1020,N_1456);
or U2910 (N_2910,N_1826,N_1967);
xnor U2911 (N_2911,N_1966,N_1942);
or U2912 (N_2912,N_1049,N_1435);
nand U2913 (N_2913,N_1513,N_1404);
xor U2914 (N_2914,N_1360,N_1344);
or U2915 (N_2915,N_1468,N_1054);
nand U2916 (N_2916,N_1175,N_1076);
xor U2917 (N_2917,N_1155,N_1864);
nor U2918 (N_2918,N_1880,N_1027);
nor U2919 (N_2919,N_1834,N_1508);
nor U2920 (N_2920,N_1100,N_1292);
or U2921 (N_2921,N_1928,N_1356);
and U2922 (N_2922,N_1210,N_1088);
nor U2923 (N_2923,N_1576,N_1590);
nand U2924 (N_2924,N_1797,N_1676);
xnor U2925 (N_2925,N_1207,N_1703);
nand U2926 (N_2926,N_1913,N_1889);
and U2927 (N_2927,N_1258,N_1741);
nor U2928 (N_2928,N_1576,N_1754);
nor U2929 (N_2929,N_1830,N_1013);
nand U2930 (N_2930,N_1915,N_1053);
xor U2931 (N_2931,N_1091,N_1283);
and U2932 (N_2932,N_1120,N_1803);
and U2933 (N_2933,N_1534,N_1959);
or U2934 (N_2934,N_1701,N_1273);
nor U2935 (N_2935,N_1745,N_1734);
nor U2936 (N_2936,N_1377,N_1083);
xor U2937 (N_2937,N_1524,N_1487);
xnor U2938 (N_2938,N_1091,N_1160);
and U2939 (N_2939,N_1773,N_1752);
or U2940 (N_2940,N_1957,N_1418);
nand U2941 (N_2941,N_1697,N_1859);
and U2942 (N_2942,N_1717,N_1172);
or U2943 (N_2943,N_1766,N_1706);
or U2944 (N_2944,N_1048,N_1550);
and U2945 (N_2945,N_1128,N_1996);
and U2946 (N_2946,N_1995,N_1211);
and U2947 (N_2947,N_1669,N_1689);
xnor U2948 (N_2948,N_1292,N_1504);
nand U2949 (N_2949,N_1988,N_1685);
xor U2950 (N_2950,N_1186,N_1452);
or U2951 (N_2951,N_1131,N_1348);
xnor U2952 (N_2952,N_1970,N_1976);
and U2953 (N_2953,N_1039,N_1688);
nor U2954 (N_2954,N_1535,N_1877);
xor U2955 (N_2955,N_1024,N_1891);
and U2956 (N_2956,N_1343,N_1606);
or U2957 (N_2957,N_1671,N_1960);
xor U2958 (N_2958,N_1458,N_1958);
and U2959 (N_2959,N_1548,N_1849);
nand U2960 (N_2960,N_1048,N_1065);
xnor U2961 (N_2961,N_1942,N_1909);
and U2962 (N_2962,N_1068,N_1850);
or U2963 (N_2963,N_1075,N_1670);
nand U2964 (N_2964,N_1825,N_1181);
xor U2965 (N_2965,N_1090,N_1214);
nand U2966 (N_2966,N_1347,N_1026);
nor U2967 (N_2967,N_1450,N_1887);
and U2968 (N_2968,N_1506,N_1257);
nor U2969 (N_2969,N_1430,N_1764);
nand U2970 (N_2970,N_1766,N_1763);
xor U2971 (N_2971,N_1647,N_1107);
nand U2972 (N_2972,N_1316,N_1507);
nor U2973 (N_2973,N_1780,N_1617);
nor U2974 (N_2974,N_1052,N_1666);
nand U2975 (N_2975,N_1429,N_1836);
nand U2976 (N_2976,N_1625,N_1218);
or U2977 (N_2977,N_1444,N_1918);
xor U2978 (N_2978,N_1455,N_1205);
and U2979 (N_2979,N_1303,N_1974);
or U2980 (N_2980,N_1604,N_1922);
nand U2981 (N_2981,N_1945,N_1032);
nor U2982 (N_2982,N_1746,N_1445);
or U2983 (N_2983,N_1367,N_1958);
and U2984 (N_2984,N_1892,N_1880);
nor U2985 (N_2985,N_1694,N_1838);
or U2986 (N_2986,N_1176,N_1890);
nor U2987 (N_2987,N_1357,N_1338);
xnor U2988 (N_2988,N_1362,N_1524);
and U2989 (N_2989,N_1157,N_1645);
nand U2990 (N_2990,N_1694,N_1087);
nor U2991 (N_2991,N_1104,N_1917);
or U2992 (N_2992,N_1182,N_1228);
or U2993 (N_2993,N_1102,N_1111);
xnor U2994 (N_2994,N_1491,N_1126);
nor U2995 (N_2995,N_1034,N_1207);
or U2996 (N_2996,N_1258,N_1417);
nor U2997 (N_2997,N_1023,N_1066);
nor U2998 (N_2998,N_1232,N_1358);
or U2999 (N_2999,N_1252,N_1217);
nand U3000 (N_3000,N_2755,N_2441);
or U3001 (N_3001,N_2480,N_2879);
nor U3002 (N_3002,N_2065,N_2208);
nand U3003 (N_3003,N_2020,N_2064);
nand U3004 (N_3004,N_2865,N_2778);
or U3005 (N_3005,N_2133,N_2558);
and U3006 (N_3006,N_2867,N_2543);
nand U3007 (N_3007,N_2469,N_2583);
xor U3008 (N_3008,N_2640,N_2106);
or U3009 (N_3009,N_2123,N_2517);
or U3010 (N_3010,N_2346,N_2040);
xnor U3011 (N_3011,N_2785,N_2393);
and U3012 (N_3012,N_2807,N_2304);
or U3013 (N_3013,N_2895,N_2787);
or U3014 (N_3014,N_2137,N_2608);
and U3015 (N_3015,N_2868,N_2345);
and U3016 (N_3016,N_2662,N_2666);
nand U3017 (N_3017,N_2988,N_2170);
xnor U3018 (N_3018,N_2436,N_2426);
nor U3019 (N_3019,N_2748,N_2049);
or U3020 (N_3020,N_2761,N_2111);
xor U3021 (N_3021,N_2779,N_2474);
or U3022 (N_3022,N_2844,N_2802);
nor U3023 (N_3023,N_2401,N_2103);
nand U3024 (N_3024,N_2708,N_2042);
nor U3025 (N_3025,N_2764,N_2015);
or U3026 (N_3026,N_2570,N_2364);
xnor U3027 (N_3027,N_2655,N_2857);
nor U3028 (N_3028,N_2523,N_2860);
xnor U3029 (N_3029,N_2335,N_2855);
or U3030 (N_3030,N_2941,N_2265);
or U3031 (N_3031,N_2997,N_2925);
and U3032 (N_3032,N_2890,N_2544);
xnor U3033 (N_3033,N_2944,N_2097);
xor U3034 (N_3034,N_2035,N_2612);
and U3035 (N_3035,N_2102,N_2771);
and U3036 (N_3036,N_2502,N_2915);
nor U3037 (N_3037,N_2260,N_2278);
or U3038 (N_3038,N_2720,N_2846);
or U3039 (N_3039,N_2358,N_2383);
and U3040 (N_3040,N_2631,N_2684);
or U3041 (N_3041,N_2200,N_2812);
or U3042 (N_3042,N_2117,N_2396);
nand U3043 (N_3043,N_2786,N_2562);
xor U3044 (N_3044,N_2759,N_2829);
xor U3045 (N_3045,N_2847,N_2365);
nand U3046 (N_3046,N_2861,N_2987);
nand U3047 (N_3047,N_2242,N_2859);
or U3048 (N_3048,N_2238,N_2391);
xor U3049 (N_3049,N_2830,N_2984);
and U3050 (N_3050,N_2501,N_2023);
or U3051 (N_3051,N_2649,N_2394);
nand U3052 (N_3052,N_2813,N_2456);
nor U3053 (N_3053,N_2189,N_2642);
and U3054 (N_3054,N_2418,N_2369);
nand U3055 (N_3055,N_2176,N_2713);
nor U3056 (N_3056,N_2085,N_2164);
nor U3057 (N_3057,N_2992,N_2680);
xnor U3058 (N_3058,N_2719,N_2279);
or U3059 (N_3059,N_2076,N_2781);
xor U3060 (N_3060,N_2343,N_2109);
nand U3061 (N_3061,N_2425,N_2247);
and U3062 (N_3062,N_2810,N_2332);
or U3063 (N_3063,N_2739,N_2950);
xnor U3064 (N_3064,N_2055,N_2679);
nand U3065 (N_3065,N_2478,N_2257);
xnor U3066 (N_3066,N_2016,N_2473);
xnor U3067 (N_3067,N_2309,N_2460);
or U3068 (N_3068,N_2917,N_2653);
and U3069 (N_3069,N_2609,N_2689);
nand U3070 (N_3070,N_2591,N_2906);
and U3071 (N_3071,N_2534,N_2316);
and U3072 (N_3072,N_2096,N_2700);
nand U3073 (N_3073,N_2008,N_2734);
nand U3074 (N_3074,N_2766,N_2530);
nor U3075 (N_3075,N_2089,N_2465);
nor U3076 (N_3076,N_2047,N_2453);
or U3077 (N_3077,N_2535,N_2056);
or U3078 (N_3078,N_2281,N_2407);
or U3079 (N_3079,N_2538,N_2427);
nand U3080 (N_3080,N_2930,N_2045);
xor U3081 (N_3081,N_2409,N_2773);
or U3082 (N_3082,N_2710,N_2240);
nor U3083 (N_3083,N_2521,N_2131);
or U3084 (N_3084,N_2126,N_2792);
or U3085 (N_3085,N_2156,N_2228);
or U3086 (N_3086,N_2158,N_2754);
or U3087 (N_3087,N_2081,N_2439);
and U3088 (N_3088,N_2869,N_2485);
xnor U3089 (N_3089,N_2641,N_2326);
and U3090 (N_3090,N_2313,N_2797);
and U3091 (N_3091,N_2901,N_2337);
or U3092 (N_3092,N_2576,N_2516);
and U3093 (N_3093,N_2590,N_2034);
nor U3094 (N_3094,N_2083,N_2665);
nor U3095 (N_3095,N_2673,N_2549);
xor U3096 (N_3096,N_2408,N_2205);
nor U3097 (N_3097,N_2455,N_2490);
xor U3098 (N_3098,N_2273,N_2163);
nand U3099 (N_3099,N_2774,N_2211);
or U3100 (N_3100,N_2889,N_2522);
nor U3101 (N_3101,N_2004,N_2715);
or U3102 (N_3102,N_2765,N_2705);
nor U3103 (N_3103,N_2822,N_2723);
nor U3104 (N_3104,N_2028,N_2216);
or U3105 (N_3105,N_2139,N_2561);
or U3106 (N_3106,N_2874,N_2491);
xor U3107 (N_3107,N_2972,N_2617);
xor U3108 (N_3108,N_2448,N_2018);
and U3109 (N_3109,N_2054,N_2149);
xor U3110 (N_3110,N_2645,N_2563);
nand U3111 (N_3111,N_2373,N_2266);
xnor U3112 (N_3112,N_2237,N_2498);
nand U3113 (N_3113,N_2671,N_2864);
or U3114 (N_3114,N_2360,N_2142);
nand U3115 (N_3115,N_2185,N_2012);
nor U3116 (N_3116,N_2716,N_2721);
nor U3117 (N_3117,N_2479,N_2637);
xor U3118 (N_3118,N_2957,N_2752);
nor U3119 (N_3119,N_2610,N_2887);
and U3120 (N_3120,N_2438,N_2589);
and U3121 (N_3121,N_2294,N_2573);
xor U3122 (N_3122,N_2512,N_2132);
nor U3123 (N_3123,N_2146,N_2660);
xor U3124 (N_3124,N_2419,N_2220);
nor U3125 (N_3125,N_2134,N_2735);
xor U3126 (N_3126,N_2046,N_2392);
xor U3127 (N_3127,N_2722,N_2977);
nor U3128 (N_3128,N_2282,N_2619);
nand U3129 (N_3129,N_2504,N_2525);
nor U3130 (N_3130,N_2644,N_2935);
nand U3131 (N_3131,N_2592,N_2798);
xor U3132 (N_3132,N_2799,N_2800);
nor U3133 (N_3133,N_2330,N_2922);
nor U3134 (N_3134,N_2036,N_2875);
nand U3135 (N_3135,N_2454,N_2937);
xor U3136 (N_3136,N_2301,N_2733);
xnor U3137 (N_3137,N_2010,N_2921);
or U3138 (N_3138,N_2470,N_2809);
and U3139 (N_3139,N_2091,N_2537);
and U3140 (N_3140,N_2732,N_2528);
nand U3141 (N_3141,N_2758,N_2298);
xnor U3142 (N_3142,N_2581,N_2390);
nor U3143 (N_3143,N_2214,N_2569);
or U3144 (N_3144,N_2661,N_2577);
nand U3145 (N_3145,N_2731,N_2099);
xor U3146 (N_3146,N_2956,N_2995);
or U3147 (N_3147,N_2414,N_2753);
nand U3148 (N_3148,N_2295,N_2351);
nor U3149 (N_3149,N_2918,N_2958);
xnor U3150 (N_3150,N_2420,N_2912);
nand U3151 (N_3151,N_2746,N_2952);
and U3152 (N_3152,N_2652,N_2994);
or U3153 (N_3153,N_2635,N_2938);
nor U3154 (N_3154,N_2670,N_2724);
or U3155 (N_3155,N_2225,N_2738);
or U3156 (N_3156,N_2333,N_2587);
nand U3157 (N_3157,N_2467,N_2495);
nor U3158 (N_3158,N_2442,N_2902);
and U3159 (N_3159,N_2234,N_2325);
and U3160 (N_3160,N_2695,N_2182);
xor U3161 (N_3161,N_2384,N_2698);
and U3162 (N_3162,N_2772,N_2461);
nand U3163 (N_3163,N_2595,N_2924);
nand U3164 (N_3164,N_2511,N_2468);
or U3165 (N_3165,N_2604,N_2704);
xnor U3166 (N_3166,N_2751,N_2848);
and U3167 (N_3167,N_2388,N_2990);
or U3168 (N_3168,N_2622,N_2310);
or U3169 (N_3169,N_2775,N_2380);
xor U3170 (N_3170,N_2885,N_2639);
xor U3171 (N_3171,N_2699,N_2368);
and U3172 (N_3172,N_2566,N_2080);
nand U3173 (N_3173,N_2006,N_2709);
nor U3174 (N_3174,N_2334,N_2446);
and U3175 (N_3175,N_2614,N_2227);
nor U3176 (N_3176,N_2362,N_2066);
nor U3177 (N_3177,N_2029,N_2946);
xnor U3178 (N_3178,N_2850,N_2090);
or U3179 (N_3179,N_2411,N_2253);
or U3180 (N_3180,N_2873,N_2820);
or U3181 (N_3181,N_2296,N_2181);
or U3182 (N_3182,N_2877,N_2905);
or U3183 (N_3183,N_2967,N_2180);
nand U3184 (N_3184,N_2236,N_2808);
and U3185 (N_3185,N_2959,N_2487);
nand U3186 (N_3186,N_2472,N_2776);
nand U3187 (N_3187,N_2542,N_2389);
or U3188 (N_3188,N_2274,N_2231);
or U3189 (N_3189,N_2415,N_2361);
xor U3190 (N_3190,N_2508,N_2329);
xnor U3191 (N_3191,N_2607,N_2378);
xnor U3192 (N_3192,N_2302,N_2536);
and U3193 (N_3193,N_2352,N_2140);
nand U3194 (N_3194,N_2311,N_2038);
nor U3195 (N_3195,N_2588,N_2152);
nor U3196 (N_3196,N_2199,N_2907);
nand U3197 (N_3197,N_2062,N_2736);
and U3198 (N_3198,N_2936,N_2672);
nor U3199 (N_3199,N_2837,N_2340);
nor U3200 (N_3200,N_2806,N_2878);
or U3201 (N_3201,N_2039,N_2961);
nand U3202 (N_3202,N_2819,N_2261);
nor U3203 (N_3203,N_2688,N_2651);
or U3204 (N_3204,N_2423,N_2969);
nand U3205 (N_3205,N_2572,N_2078);
nor U3206 (N_3206,N_2048,N_2899);
xnor U3207 (N_3207,N_2694,N_2285);
or U3208 (N_3208,N_2367,N_2726);
or U3209 (N_3209,N_2175,N_2827);
and U3210 (N_3210,N_2908,N_2954);
nor U3211 (N_3211,N_2267,N_2903);
or U3212 (N_3212,N_2741,N_2965);
nor U3213 (N_3213,N_2618,N_2585);
nand U3214 (N_3214,N_2114,N_2763);
and U3215 (N_3215,N_2318,N_2292);
and U3216 (N_3216,N_2059,N_2596);
and U3217 (N_3217,N_2675,N_2186);
xnor U3218 (N_3218,N_2852,N_2603);
or U3219 (N_3219,N_2818,N_2434);
and U3220 (N_3220,N_2451,N_2219);
or U3221 (N_3221,N_2854,N_2206);
xor U3222 (N_3222,N_2832,N_2482);
xor U3223 (N_3223,N_2286,N_2744);
xor U3224 (N_3224,N_2853,N_2385);
and U3225 (N_3225,N_2658,N_2375);
nand U3226 (N_3226,N_2341,N_2061);
xor U3227 (N_3227,N_2983,N_2963);
or U3228 (N_3228,N_2239,N_2481);
nor U3229 (N_3229,N_2728,N_2223);
nand U3230 (N_3230,N_2030,N_2740);
xnor U3231 (N_3231,N_2663,N_2022);
or U3232 (N_3232,N_2322,N_2013);
nand U3233 (N_3233,N_2578,N_2410);
xor U3234 (N_3234,N_2221,N_2664);
xor U3235 (N_3235,N_2399,N_2518);
nor U3236 (N_3236,N_2226,N_2377);
xor U3237 (N_3237,N_2336,N_2998);
nand U3238 (N_3238,N_2945,N_2909);
or U3239 (N_3239,N_2043,N_2087);
nor U3240 (N_3240,N_2009,N_2307);
nand U3241 (N_3241,N_2553,N_2347);
nand U3242 (N_3242,N_2729,N_2696);
xor U3243 (N_3243,N_2898,N_2403);
nand U3244 (N_3244,N_2546,N_2510);
xnor U3245 (N_3245,N_2252,N_2489);
nand U3246 (N_3246,N_2184,N_2691);
and U3247 (N_3247,N_2193,N_2230);
nand U3248 (N_3248,N_2677,N_2027);
or U3249 (N_3249,N_2654,N_2305);
and U3250 (N_3250,N_2623,N_2058);
or U3251 (N_3251,N_2624,N_2063);
nor U3252 (N_3252,N_2835,N_2817);
nor U3253 (N_3253,N_2110,N_2801);
nand U3254 (N_3254,N_2883,N_2412);
and U3255 (N_3255,N_2217,N_2756);
or U3256 (N_3256,N_2145,N_2981);
xnor U3257 (N_3257,N_2750,N_2559);
or U3258 (N_3258,N_2505,N_2457);
xnor U3259 (N_3259,N_2191,N_2327);
and U3260 (N_3260,N_2920,N_2471);
and U3261 (N_3261,N_2506,N_2381);
nand U3262 (N_3262,N_2633,N_2284);
and U3263 (N_3263,N_2833,N_2567);
or U3264 (N_3264,N_2727,N_2440);
and U3265 (N_3265,N_2683,N_2079);
and U3266 (N_3266,N_2711,N_2795);
xnor U3267 (N_3267,N_2093,N_2975);
nand U3268 (N_3268,N_2714,N_2162);
xor U3269 (N_3269,N_2195,N_2116);
nor U3270 (N_3270,N_2843,N_2463);
xnor U3271 (N_3271,N_2355,N_2911);
nand U3272 (N_3272,N_2914,N_2507);
nor U3273 (N_3273,N_2836,N_2929);
nand U3274 (N_3274,N_2620,N_2277);
and U3275 (N_3275,N_2119,N_2449);
nand U3276 (N_3276,N_2202,N_2319);
nor U3277 (N_3277,N_2250,N_2526);
xnor U3278 (N_3278,N_2207,N_2976);
or U3279 (N_3279,N_2026,N_2953);
and U3280 (N_3280,N_2107,N_2387);
nor U3281 (N_3281,N_2628,N_2703);
or U3282 (N_3282,N_2767,N_2224);
or U3283 (N_3283,N_2057,N_2173);
and U3284 (N_3284,N_2290,N_2594);
and U3285 (N_3285,N_2514,N_2991);
and U3286 (N_3286,N_2215,N_2357);
and U3287 (N_3287,N_2031,N_2300);
or U3288 (N_3288,N_2552,N_2769);
xnor U3289 (N_3289,N_2476,N_2105);
or U3290 (N_3290,N_2303,N_2229);
and U3291 (N_3291,N_2916,N_2678);
or U3292 (N_3292,N_2007,N_2674);
nand U3293 (N_3293,N_2147,N_2749);
and U3294 (N_3294,N_2932,N_2073);
nand U3295 (N_3295,N_2101,N_2315);
nor U3296 (N_3296,N_2160,N_2893);
nand U3297 (N_3297,N_2297,N_2627);
nand U3298 (N_3298,N_2509,N_2973);
and U3299 (N_3299,N_2574,N_2762);
or U3300 (N_3300,N_2177,N_2376);
nor U3301 (N_3301,N_2520,N_2138);
nand U3302 (N_3302,N_2565,N_2086);
nand U3303 (N_3303,N_2613,N_2657);
and U3304 (N_3304,N_2095,N_2122);
nor U3305 (N_3305,N_2070,N_2112);
xor U3306 (N_3306,N_2349,N_2980);
nor U3307 (N_3307,N_2784,N_2320);
nor U3308 (N_3308,N_2494,N_2712);
xor U3309 (N_3309,N_2796,N_2169);
nand U3310 (N_3310,N_2141,N_2743);
nor U3311 (N_3311,N_2880,N_2650);
and U3312 (N_3312,N_2458,N_2165);
or U3313 (N_3313,N_2350,N_2218);
and U3314 (N_3314,N_2533,N_2584);
and U3315 (N_3315,N_2308,N_2851);
xnor U3316 (N_3316,N_2730,N_2823);
and U3317 (N_3317,N_2276,N_2582);
nor U3318 (N_3318,N_2249,N_2372);
xor U3319 (N_3319,N_2477,N_2209);
xor U3320 (N_3320,N_2702,N_2601);
nand U3321 (N_3321,N_2791,N_2725);
nand U3322 (N_3322,N_2259,N_2246);
nor U3323 (N_3323,N_2268,N_2192);
nand U3324 (N_3324,N_2269,N_2891);
and U3325 (N_3325,N_2964,N_2545);
nor U3326 (N_3326,N_2475,N_2421);
nand U3327 (N_3327,N_2747,N_2556);
nor U3328 (N_3328,N_2187,N_2328);
and U3329 (N_3329,N_2245,N_2262);
and U3330 (N_3330,N_2821,N_2519);
xnor U3331 (N_3331,N_2052,N_2154);
and U3332 (N_3332,N_2737,N_2831);
and U3333 (N_3333,N_2805,N_2032);
and U3334 (N_3334,N_2636,N_2135);
or U3335 (N_3335,N_2452,N_2148);
xor U3336 (N_3336,N_2982,N_2824);
nor U3337 (N_3337,N_2579,N_2757);
or U3338 (N_3338,N_2892,N_2264);
and U3339 (N_3339,N_2551,N_2000);
nor U3340 (N_3340,N_2586,N_2197);
nand U3341 (N_3341,N_2524,N_2499);
nor U3342 (N_3342,N_2210,N_2804);
nor U3343 (N_3343,N_2171,N_2212);
and U3344 (N_3344,N_2437,N_2190);
or U3345 (N_3345,N_2404,N_2430);
xnor U3346 (N_3346,N_2493,N_2842);
xnor U3347 (N_3347,N_2069,N_2539);
nand U3348 (N_3348,N_2621,N_2232);
xnor U3349 (N_3349,N_2659,N_2996);
or U3350 (N_3350,N_2400,N_2803);
xor U3351 (N_3351,N_2428,N_2356);
xor U3352 (N_3352,N_2024,N_2872);
xnor U3353 (N_3353,N_2432,N_2940);
and U3354 (N_3354,N_2926,N_2834);
xnor U3355 (N_3355,N_2235,N_2483);
xnor U3356 (N_3356,N_2331,N_2939);
nor U3357 (N_3357,N_2782,N_2989);
nand U3358 (N_3358,N_2575,N_2841);
and U3359 (N_3359,N_2615,N_2629);
xor U3360 (N_3360,N_2971,N_2179);
or U3361 (N_3361,N_2422,N_2166);
or U3362 (N_3362,N_2405,N_2011);
and U3363 (N_3363,N_2100,N_2815);
nand U3364 (N_3364,N_2198,N_2488);
nand U3365 (N_3365,N_2094,N_2993);
and U3366 (N_3366,N_2634,N_2985);
or U3367 (N_3367,N_2676,N_2910);
nor U3368 (N_3368,N_2406,N_2204);
nand U3369 (N_3369,N_2287,N_2697);
xor U3370 (N_3370,N_2363,N_2760);
or U3371 (N_3371,N_2072,N_2560);
or U3372 (N_3372,N_2129,N_2717);
nor U3373 (N_3373,N_2647,N_2339);
nor U3374 (N_3374,N_2690,N_2338);
and U3375 (N_3375,N_2082,N_2681);
nand U3376 (N_3376,N_2611,N_2194);
xor U3377 (N_3377,N_2433,N_2075);
nor U3378 (N_3378,N_2682,N_2839);
or U3379 (N_3379,N_2118,N_2547);
xnor U3380 (N_3380,N_2793,N_2386);
or U3381 (N_3381,N_2243,N_2923);
nor U3382 (N_3382,N_2395,N_2770);
and U3383 (N_3383,N_2067,N_2084);
or U3384 (N_3384,N_2557,N_2002);
nand U3385 (N_3385,N_2413,N_2382);
and U3386 (N_3386,N_2638,N_2271);
and U3387 (N_3387,N_2445,N_2155);
or U3388 (N_3388,N_2685,N_2017);
nor U3389 (N_3389,N_2856,N_2254);
nor U3390 (N_3390,N_2088,N_2258);
nand U3391 (N_3391,N_2288,N_2951);
or U3392 (N_3392,N_2667,N_2417);
nor U3393 (N_3393,N_2707,N_2866);
nor U3394 (N_3394,N_2120,N_2599);
or U3395 (N_3395,N_2464,N_2255);
or U3396 (N_3396,N_2379,N_2606);
nor U3397 (N_3397,N_2115,N_2077);
and U3398 (N_3398,N_2927,N_2931);
nor U3399 (N_3399,N_2768,N_2492);
and U3400 (N_3400,N_2450,N_2625);
nand U3401 (N_3401,N_2955,N_2974);
xor U3402 (N_3402,N_2527,N_2317);
and U3403 (N_3403,N_2669,N_2263);
nor U3404 (N_3404,N_2150,N_2130);
or U3405 (N_3405,N_2870,N_2144);
or U3406 (N_3406,N_2484,N_2718);
nor U3407 (N_3407,N_2021,N_2001);
and U3408 (N_3408,N_2071,N_2780);
and U3409 (N_3409,N_2306,N_2121);
nand U3410 (N_3410,N_2323,N_2025);
and U3411 (N_3411,N_2999,N_2687);
nand U3412 (N_3412,N_2580,N_2248);
and U3413 (N_3413,N_2882,N_2568);
xnor U3414 (N_3414,N_2275,N_2053);
or U3415 (N_3415,N_2529,N_2648);
nor U3416 (N_3416,N_2466,N_2943);
and U3417 (N_3417,N_2978,N_2656);
and U3418 (N_3418,N_2188,N_2816);
xor U3419 (N_3419,N_2104,N_2630);
xnor U3420 (N_3420,N_2092,N_2348);
and U3421 (N_3421,N_2033,N_2374);
nor U3422 (N_3422,N_2431,N_2256);
or U3423 (N_3423,N_2632,N_2602);
xnor U3424 (N_3424,N_2966,N_2244);
and U3425 (N_3425,N_2321,N_2960);
xor U3426 (N_3426,N_2496,N_2098);
xnor U3427 (N_3427,N_2462,N_2359);
nand U3428 (N_3428,N_2222,N_2203);
nor U3429 (N_3429,N_2692,N_2933);
nand U3430 (N_3430,N_2597,N_2108);
or U3431 (N_3431,N_2157,N_2826);
or U3432 (N_3432,N_2968,N_2497);
nor U3433 (N_3433,N_2037,N_2789);
nand U3434 (N_3434,N_2897,N_2353);
and U3435 (N_3435,N_2904,N_2811);
nand U3436 (N_3436,N_2429,N_2948);
nor U3437 (N_3437,N_2828,N_2435);
nor U3438 (N_3438,N_2598,N_2128);
nor U3439 (N_3439,N_2600,N_2143);
and U3440 (N_3440,N_2862,N_2970);
xor U3441 (N_3441,N_2686,N_2444);
and U3442 (N_3442,N_2161,N_2174);
and U3443 (N_3443,N_2884,N_2900);
nor U3444 (N_3444,N_2044,N_2486);
or U3445 (N_3445,N_2014,N_2532);
and U3446 (N_3446,N_2178,N_2459);
nor U3447 (N_3447,N_2370,N_2788);
nor U3448 (N_3448,N_2515,N_2125);
xnor U3449 (N_3449,N_2668,N_2113);
nor U3450 (N_3450,N_2881,N_2919);
and U3451 (N_3451,N_2947,N_2183);
xor U3452 (N_3452,N_2825,N_2402);
or U3453 (N_3453,N_2742,N_2074);
or U3454 (N_3454,N_2783,N_2794);
and U3455 (N_3455,N_2777,N_2503);
or U3456 (N_3456,N_2863,N_2342);
nand U3457 (N_3457,N_2643,N_2314);
nor U3458 (N_3458,N_2845,N_2003);
and U3459 (N_3459,N_2251,N_2127);
and U3460 (N_3460,N_2858,N_2366);
and U3461 (N_3461,N_2886,N_2068);
nand U3462 (N_3462,N_2172,N_2443);
or U3463 (N_3463,N_2280,N_2564);
and U3464 (N_3464,N_2888,N_2554);
nand U3465 (N_3465,N_2019,N_2201);
xor U3466 (N_3466,N_2398,N_2159);
nand U3467 (N_3467,N_2051,N_2397);
nand U3468 (N_3468,N_2312,N_2041);
nand U3469 (N_3469,N_2555,N_2060);
or U3470 (N_3470,N_2593,N_2934);
nor U3471 (N_3471,N_2701,N_2876);
xor U3472 (N_3472,N_2706,N_2124);
nand U3473 (N_3473,N_2151,N_2324);
nor U3474 (N_3474,N_2293,N_2894);
nor U3475 (N_3475,N_2371,N_2196);
nand U3476 (N_3476,N_2838,N_2354);
and U3477 (N_3477,N_2416,N_2213);
xnor U3478 (N_3478,N_2550,N_2272);
xnor U3479 (N_3479,N_2790,N_2168);
nor U3480 (N_3480,N_2167,N_2840);
nor U3481 (N_3481,N_2942,N_2626);
or U3482 (N_3482,N_2605,N_2986);
nor U3483 (N_3483,N_2241,N_2814);
and U3484 (N_3484,N_2447,N_2693);
and U3485 (N_3485,N_2541,N_2849);
or U3486 (N_3486,N_2962,N_2540);
or U3487 (N_3487,N_2050,N_2424);
nor U3488 (N_3488,N_2500,N_2289);
xor U3489 (N_3489,N_2979,N_2299);
or U3490 (N_3490,N_2896,N_2913);
nor U3491 (N_3491,N_2571,N_2949);
nor U3492 (N_3492,N_2871,N_2531);
or U3493 (N_3493,N_2291,N_2513);
nand U3494 (N_3494,N_2283,N_2136);
or U3495 (N_3495,N_2928,N_2270);
nor U3496 (N_3496,N_2005,N_2233);
xnor U3497 (N_3497,N_2616,N_2344);
nand U3498 (N_3498,N_2745,N_2646);
xor U3499 (N_3499,N_2548,N_2153);
nand U3500 (N_3500,N_2403,N_2223);
xor U3501 (N_3501,N_2729,N_2296);
and U3502 (N_3502,N_2730,N_2392);
xnor U3503 (N_3503,N_2796,N_2250);
nor U3504 (N_3504,N_2550,N_2267);
nor U3505 (N_3505,N_2773,N_2930);
and U3506 (N_3506,N_2727,N_2020);
nand U3507 (N_3507,N_2454,N_2989);
xor U3508 (N_3508,N_2821,N_2473);
and U3509 (N_3509,N_2568,N_2765);
or U3510 (N_3510,N_2251,N_2991);
nand U3511 (N_3511,N_2690,N_2645);
nor U3512 (N_3512,N_2222,N_2032);
nor U3513 (N_3513,N_2214,N_2868);
or U3514 (N_3514,N_2594,N_2624);
or U3515 (N_3515,N_2146,N_2044);
nor U3516 (N_3516,N_2841,N_2378);
and U3517 (N_3517,N_2497,N_2763);
and U3518 (N_3518,N_2516,N_2374);
xnor U3519 (N_3519,N_2458,N_2601);
nor U3520 (N_3520,N_2889,N_2313);
or U3521 (N_3521,N_2789,N_2672);
xnor U3522 (N_3522,N_2094,N_2691);
or U3523 (N_3523,N_2022,N_2713);
nand U3524 (N_3524,N_2784,N_2692);
xnor U3525 (N_3525,N_2763,N_2275);
xor U3526 (N_3526,N_2639,N_2669);
or U3527 (N_3527,N_2810,N_2353);
nor U3528 (N_3528,N_2274,N_2774);
or U3529 (N_3529,N_2179,N_2598);
xor U3530 (N_3530,N_2164,N_2854);
xnor U3531 (N_3531,N_2281,N_2239);
nand U3532 (N_3532,N_2525,N_2828);
and U3533 (N_3533,N_2730,N_2414);
and U3534 (N_3534,N_2471,N_2271);
xnor U3535 (N_3535,N_2787,N_2688);
or U3536 (N_3536,N_2647,N_2896);
nor U3537 (N_3537,N_2482,N_2082);
nand U3538 (N_3538,N_2601,N_2616);
nand U3539 (N_3539,N_2649,N_2689);
and U3540 (N_3540,N_2189,N_2649);
nor U3541 (N_3541,N_2059,N_2743);
nor U3542 (N_3542,N_2388,N_2077);
nor U3543 (N_3543,N_2289,N_2322);
nand U3544 (N_3544,N_2950,N_2606);
nand U3545 (N_3545,N_2885,N_2384);
or U3546 (N_3546,N_2615,N_2353);
xor U3547 (N_3547,N_2772,N_2091);
or U3548 (N_3548,N_2573,N_2039);
nand U3549 (N_3549,N_2671,N_2406);
and U3550 (N_3550,N_2314,N_2494);
nand U3551 (N_3551,N_2168,N_2922);
and U3552 (N_3552,N_2002,N_2372);
nand U3553 (N_3553,N_2580,N_2962);
or U3554 (N_3554,N_2902,N_2878);
or U3555 (N_3555,N_2341,N_2268);
xor U3556 (N_3556,N_2936,N_2397);
and U3557 (N_3557,N_2276,N_2063);
nand U3558 (N_3558,N_2225,N_2790);
nand U3559 (N_3559,N_2596,N_2196);
nand U3560 (N_3560,N_2439,N_2456);
or U3561 (N_3561,N_2592,N_2262);
nand U3562 (N_3562,N_2251,N_2805);
nand U3563 (N_3563,N_2092,N_2416);
or U3564 (N_3564,N_2434,N_2752);
and U3565 (N_3565,N_2402,N_2662);
xnor U3566 (N_3566,N_2223,N_2130);
nor U3567 (N_3567,N_2307,N_2946);
nor U3568 (N_3568,N_2324,N_2762);
nand U3569 (N_3569,N_2601,N_2968);
xor U3570 (N_3570,N_2960,N_2630);
or U3571 (N_3571,N_2503,N_2368);
and U3572 (N_3572,N_2996,N_2859);
or U3573 (N_3573,N_2050,N_2959);
xnor U3574 (N_3574,N_2295,N_2652);
or U3575 (N_3575,N_2834,N_2523);
nand U3576 (N_3576,N_2651,N_2551);
nor U3577 (N_3577,N_2187,N_2418);
xnor U3578 (N_3578,N_2587,N_2064);
nor U3579 (N_3579,N_2544,N_2000);
xor U3580 (N_3580,N_2593,N_2024);
nand U3581 (N_3581,N_2796,N_2534);
xor U3582 (N_3582,N_2694,N_2640);
nand U3583 (N_3583,N_2349,N_2381);
nor U3584 (N_3584,N_2783,N_2921);
xnor U3585 (N_3585,N_2056,N_2709);
or U3586 (N_3586,N_2335,N_2023);
nand U3587 (N_3587,N_2335,N_2696);
or U3588 (N_3588,N_2325,N_2781);
xnor U3589 (N_3589,N_2980,N_2345);
xor U3590 (N_3590,N_2843,N_2219);
nor U3591 (N_3591,N_2093,N_2389);
and U3592 (N_3592,N_2548,N_2946);
xor U3593 (N_3593,N_2093,N_2201);
nand U3594 (N_3594,N_2016,N_2811);
xor U3595 (N_3595,N_2246,N_2336);
nand U3596 (N_3596,N_2687,N_2866);
nand U3597 (N_3597,N_2123,N_2027);
or U3598 (N_3598,N_2620,N_2547);
and U3599 (N_3599,N_2910,N_2790);
and U3600 (N_3600,N_2680,N_2619);
nand U3601 (N_3601,N_2421,N_2922);
nand U3602 (N_3602,N_2296,N_2662);
xor U3603 (N_3603,N_2617,N_2698);
nand U3604 (N_3604,N_2269,N_2203);
xor U3605 (N_3605,N_2360,N_2829);
xor U3606 (N_3606,N_2821,N_2111);
xnor U3607 (N_3607,N_2933,N_2965);
and U3608 (N_3608,N_2786,N_2131);
nor U3609 (N_3609,N_2833,N_2153);
and U3610 (N_3610,N_2971,N_2892);
nor U3611 (N_3611,N_2410,N_2758);
nand U3612 (N_3612,N_2511,N_2398);
xor U3613 (N_3613,N_2563,N_2722);
nor U3614 (N_3614,N_2619,N_2050);
xor U3615 (N_3615,N_2038,N_2223);
xor U3616 (N_3616,N_2074,N_2680);
nor U3617 (N_3617,N_2297,N_2105);
nand U3618 (N_3618,N_2256,N_2791);
and U3619 (N_3619,N_2204,N_2121);
or U3620 (N_3620,N_2061,N_2263);
nor U3621 (N_3621,N_2609,N_2017);
nor U3622 (N_3622,N_2565,N_2793);
xnor U3623 (N_3623,N_2121,N_2447);
nand U3624 (N_3624,N_2307,N_2609);
and U3625 (N_3625,N_2844,N_2205);
nor U3626 (N_3626,N_2317,N_2819);
nand U3627 (N_3627,N_2549,N_2944);
or U3628 (N_3628,N_2260,N_2759);
xor U3629 (N_3629,N_2419,N_2055);
xnor U3630 (N_3630,N_2996,N_2928);
nand U3631 (N_3631,N_2673,N_2958);
or U3632 (N_3632,N_2193,N_2375);
or U3633 (N_3633,N_2019,N_2503);
or U3634 (N_3634,N_2866,N_2136);
or U3635 (N_3635,N_2091,N_2828);
xnor U3636 (N_3636,N_2404,N_2318);
nor U3637 (N_3637,N_2862,N_2724);
and U3638 (N_3638,N_2224,N_2086);
and U3639 (N_3639,N_2389,N_2749);
xnor U3640 (N_3640,N_2981,N_2871);
nand U3641 (N_3641,N_2642,N_2522);
and U3642 (N_3642,N_2609,N_2793);
nor U3643 (N_3643,N_2029,N_2141);
or U3644 (N_3644,N_2932,N_2978);
or U3645 (N_3645,N_2263,N_2080);
and U3646 (N_3646,N_2377,N_2128);
nor U3647 (N_3647,N_2358,N_2927);
xor U3648 (N_3648,N_2236,N_2610);
nand U3649 (N_3649,N_2191,N_2528);
xnor U3650 (N_3650,N_2354,N_2446);
and U3651 (N_3651,N_2017,N_2778);
or U3652 (N_3652,N_2614,N_2550);
and U3653 (N_3653,N_2122,N_2109);
or U3654 (N_3654,N_2180,N_2585);
xnor U3655 (N_3655,N_2706,N_2460);
and U3656 (N_3656,N_2628,N_2697);
xor U3657 (N_3657,N_2122,N_2390);
and U3658 (N_3658,N_2354,N_2219);
nor U3659 (N_3659,N_2534,N_2484);
nand U3660 (N_3660,N_2843,N_2468);
nand U3661 (N_3661,N_2533,N_2911);
or U3662 (N_3662,N_2436,N_2493);
nor U3663 (N_3663,N_2484,N_2750);
or U3664 (N_3664,N_2761,N_2518);
nand U3665 (N_3665,N_2823,N_2314);
nand U3666 (N_3666,N_2887,N_2989);
and U3667 (N_3667,N_2571,N_2736);
nand U3668 (N_3668,N_2661,N_2733);
nor U3669 (N_3669,N_2311,N_2598);
or U3670 (N_3670,N_2160,N_2295);
nor U3671 (N_3671,N_2796,N_2967);
xor U3672 (N_3672,N_2826,N_2635);
nor U3673 (N_3673,N_2061,N_2700);
nor U3674 (N_3674,N_2126,N_2022);
or U3675 (N_3675,N_2980,N_2549);
nand U3676 (N_3676,N_2759,N_2243);
or U3677 (N_3677,N_2042,N_2941);
nand U3678 (N_3678,N_2605,N_2495);
xor U3679 (N_3679,N_2545,N_2919);
nand U3680 (N_3680,N_2937,N_2067);
nand U3681 (N_3681,N_2224,N_2545);
and U3682 (N_3682,N_2683,N_2354);
xnor U3683 (N_3683,N_2516,N_2074);
nor U3684 (N_3684,N_2558,N_2652);
and U3685 (N_3685,N_2081,N_2722);
nor U3686 (N_3686,N_2576,N_2001);
and U3687 (N_3687,N_2094,N_2842);
or U3688 (N_3688,N_2985,N_2151);
nor U3689 (N_3689,N_2216,N_2061);
nor U3690 (N_3690,N_2747,N_2113);
nand U3691 (N_3691,N_2967,N_2171);
or U3692 (N_3692,N_2676,N_2695);
or U3693 (N_3693,N_2508,N_2055);
and U3694 (N_3694,N_2155,N_2572);
and U3695 (N_3695,N_2133,N_2584);
xor U3696 (N_3696,N_2210,N_2309);
nor U3697 (N_3697,N_2573,N_2266);
nor U3698 (N_3698,N_2075,N_2545);
nand U3699 (N_3699,N_2453,N_2123);
and U3700 (N_3700,N_2547,N_2888);
nand U3701 (N_3701,N_2936,N_2207);
and U3702 (N_3702,N_2499,N_2654);
nand U3703 (N_3703,N_2572,N_2203);
nor U3704 (N_3704,N_2452,N_2897);
xor U3705 (N_3705,N_2907,N_2601);
and U3706 (N_3706,N_2690,N_2360);
and U3707 (N_3707,N_2798,N_2598);
xnor U3708 (N_3708,N_2794,N_2491);
nor U3709 (N_3709,N_2494,N_2745);
nand U3710 (N_3710,N_2504,N_2558);
xor U3711 (N_3711,N_2211,N_2396);
nand U3712 (N_3712,N_2066,N_2327);
or U3713 (N_3713,N_2698,N_2907);
nor U3714 (N_3714,N_2574,N_2896);
xor U3715 (N_3715,N_2335,N_2694);
xor U3716 (N_3716,N_2306,N_2296);
and U3717 (N_3717,N_2897,N_2815);
xor U3718 (N_3718,N_2937,N_2181);
or U3719 (N_3719,N_2224,N_2833);
xnor U3720 (N_3720,N_2187,N_2772);
xor U3721 (N_3721,N_2832,N_2034);
and U3722 (N_3722,N_2690,N_2196);
or U3723 (N_3723,N_2640,N_2525);
nand U3724 (N_3724,N_2546,N_2439);
or U3725 (N_3725,N_2293,N_2313);
or U3726 (N_3726,N_2869,N_2235);
and U3727 (N_3727,N_2697,N_2476);
or U3728 (N_3728,N_2951,N_2064);
or U3729 (N_3729,N_2903,N_2730);
nor U3730 (N_3730,N_2659,N_2602);
nand U3731 (N_3731,N_2946,N_2630);
nor U3732 (N_3732,N_2570,N_2612);
nor U3733 (N_3733,N_2910,N_2986);
xor U3734 (N_3734,N_2655,N_2149);
xnor U3735 (N_3735,N_2834,N_2169);
nor U3736 (N_3736,N_2858,N_2427);
and U3737 (N_3737,N_2394,N_2836);
nor U3738 (N_3738,N_2833,N_2857);
nand U3739 (N_3739,N_2190,N_2912);
and U3740 (N_3740,N_2740,N_2637);
and U3741 (N_3741,N_2732,N_2851);
and U3742 (N_3742,N_2485,N_2754);
or U3743 (N_3743,N_2753,N_2624);
nand U3744 (N_3744,N_2505,N_2080);
or U3745 (N_3745,N_2894,N_2840);
or U3746 (N_3746,N_2576,N_2070);
or U3747 (N_3747,N_2465,N_2799);
nor U3748 (N_3748,N_2215,N_2621);
or U3749 (N_3749,N_2019,N_2584);
and U3750 (N_3750,N_2875,N_2830);
or U3751 (N_3751,N_2902,N_2643);
nor U3752 (N_3752,N_2970,N_2802);
xnor U3753 (N_3753,N_2852,N_2418);
and U3754 (N_3754,N_2959,N_2133);
nand U3755 (N_3755,N_2451,N_2317);
nand U3756 (N_3756,N_2070,N_2737);
nand U3757 (N_3757,N_2103,N_2355);
and U3758 (N_3758,N_2485,N_2035);
nand U3759 (N_3759,N_2725,N_2116);
nand U3760 (N_3760,N_2828,N_2568);
xnor U3761 (N_3761,N_2617,N_2044);
and U3762 (N_3762,N_2547,N_2436);
or U3763 (N_3763,N_2978,N_2104);
or U3764 (N_3764,N_2304,N_2086);
and U3765 (N_3765,N_2332,N_2542);
or U3766 (N_3766,N_2929,N_2350);
nor U3767 (N_3767,N_2481,N_2292);
and U3768 (N_3768,N_2468,N_2039);
nor U3769 (N_3769,N_2818,N_2862);
nor U3770 (N_3770,N_2280,N_2850);
nand U3771 (N_3771,N_2553,N_2152);
nand U3772 (N_3772,N_2013,N_2463);
xor U3773 (N_3773,N_2440,N_2941);
xnor U3774 (N_3774,N_2102,N_2035);
and U3775 (N_3775,N_2171,N_2687);
and U3776 (N_3776,N_2996,N_2322);
or U3777 (N_3777,N_2726,N_2635);
nor U3778 (N_3778,N_2515,N_2406);
or U3779 (N_3779,N_2637,N_2921);
nand U3780 (N_3780,N_2468,N_2363);
xor U3781 (N_3781,N_2478,N_2226);
nand U3782 (N_3782,N_2150,N_2868);
and U3783 (N_3783,N_2156,N_2961);
nand U3784 (N_3784,N_2796,N_2618);
nand U3785 (N_3785,N_2700,N_2638);
nand U3786 (N_3786,N_2975,N_2538);
nand U3787 (N_3787,N_2641,N_2383);
nor U3788 (N_3788,N_2497,N_2122);
or U3789 (N_3789,N_2946,N_2747);
and U3790 (N_3790,N_2610,N_2728);
nand U3791 (N_3791,N_2292,N_2228);
or U3792 (N_3792,N_2872,N_2142);
nand U3793 (N_3793,N_2211,N_2198);
xor U3794 (N_3794,N_2787,N_2207);
and U3795 (N_3795,N_2128,N_2745);
nand U3796 (N_3796,N_2412,N_2762);
and U3797 (N_3797,N_2282,N_2900);
xor U3798 (N_3798,N_2927,N_2489);
nand U3799 (N_3799,N_2962,N_2827);
nor U3800 (N_3800,N_2808,N_2606);
and U3801 (N_3801,N_2956,N_2422);
nor U3802 (N_3802,N_2515,N_2041);
nor U3803 (N_3803,N_2993,N_2926);
xnor U3804 (N_3804,N_2729,N_2365);
and U3805 (N_3805,N_2924,N_2960);
xnor U3806 (N_3806,N_2701,N_2065);
xnor U3807 (N_3807,N_2910,N_2191);
nor U3808 (N_3808,N_2676,N_2267);
nor U3809 (N_3809,N_2126,N_2972);
xor U3810 (N_3810,N_2735,N_2936);
xor U3811 (N_3811,N_2204,N_2001);
or U3812 (N_3812,N_2167,N_2879);
or U3813 (N_3813,N_2491,N_2735);
nor U3814 (N_3814,N_2450,N_2894);
or U3815 (N_3815,N_2368,N_2151);
nand U3816 (N_3816,N_2576,N_2629);
nor U3817 (N_3817,N_2052,N_2482);
nor U3818 (N_3818,N_2822,N_2983);
nand U3819 (N_3819,N_2469,N_2099);
or U3820 (N_3820,N_2495,N_2757);
nor U3821 (N_3821,N_2072,N_2056);
and U3822 (N_3822,N_2691,N_2906);
or U3823 (N_3823,N_2445,N_2808);
xnor U3824 (N_3824,N_2707,N_2509);
and U3825 (N_3825,N_2212,N_2354);
nand U3826 (N_3826,N_2386,N_2633);
nand U3827 (N_3827,N_2472,N_2733);
and U3828 (N_3828,N_2453,N_2810);
and U3829 (N_3829,N_2142,N_2875);
and U3830 (N_3830,N_2499,N_2357);
or U3831 (N_3831,N_2864,N_2160);
and U3832 (N_3832,N_2300,N_2541);
nor U3833 (N_3833,N_2977,N_2633);
or U3834 (N_3834,N_2608,N_2008);
xor U3835 (N_3835,N_2172,N_2440);
xnor U3836 (N_3836,N_2540,N_2577);
and U3837 (N_3837,N_2197,N_2703);
nand U3838 (N_3838,N_2692,N_2833);
nand U3839 (N_3839,N_2263,N_2463);
or U3840 (N_3840,N_2552,N_2349);
or U3841 (N_3841,N_2982,N_2386);
xor U3842 (N_3842,N_2685,N_2275);
or U3843 (N_3843,N_2310,N_2397);
or U3844 (N_3844,N_2187,N_2150);
nor U3845 (N_3845,N_2687,N_2903);
nand U3846 (N_3846,N_2820,N_2785);
xor U3847 (N_3847,N_2313,N_2670);
nand U3848 (N_3848,N_2758,N_2740);
or U3849 (N_3849,N_2589,N_2923);
or U3850 (N_3850,N_2834,N_2373);
nor U3851 (N_3851,N_2136,N_2295);
and U3852 (N_3852,N_2206,N_2564);
or U3853 (N_3853,N_2013,N_2945);
xor U3854 (N_3854,N_2579,N_2680);
xnor U3855 (N_3855,N_2141,N_2636);
xnor U3856 (N_3856,N_2601,N_2292);
xnor U3857 (N_3857,N_2482,N_2857);
or U3858 (N_3858,N_2854,N_2759);
and U3859 (N_3859,N_2865,N_2204);
and U3860 (N_3860,N_2824,N_2308);
or U3861 (N_3861,N_2968,N_2033);
and U3862 (N_3862,N_2111,N_2370);
nand U3863 (N_3863,N_2631,N_2146);
or U3864 (N_3864,N_2253,N_2032);
or U3865 (N_3865,N_2506,N_2750);
nor U3866 (N_3866,N_2149,N_2517);
nand U3867 (N_3867,N_2831,N_2400);
nand U3868 (N_3868,N_2376,N_2772);
or U3869 (N_3869,N_2392,N_2610);
xor U3870 (N_3870,N_2358,N_2420);
nor U3871 (N_3871,N_2579,N_2735);
and U3872 (N_3872,N_2513,N_2861);
nor U3873 (N_3873,N_2656,N_2140);
or U3874 (N_3874,N_2626,N_2726);
or U3875 (N_3875,N_2884,N_2172);
xor U3876 (N_3876,N_2844,N_2360);
nand U3877 (N_3877,N_2962,N_2533);
or U3878 (N_3878,N_2315,N_2983);
or U3879 (N_3879,N_2940,N_2650);
or U3880 (N_3880,N_2613,N_2264);
nand U3881 (N_3881,N_2713,N_2172);
nor U3882 (N_3882,N_2384,N_2803);
nand U3883 (N_3883,N_2303,N_2374);
xnor U3884 (N_3884,N_2339,N_2166);
nor U3885 (N_3885,N_2377,N_2708);
or U3886 (N_3886,N_2284,N_2007);
xnor U3887 (N_3887,N_2330,N_2996);
or U3888 (N_3888,N_2991,N_2564);
nor U3889 (N_3889,N_2213,N_2655);
nor U3890 (N_3890,N_2618,N_2050);
or U3891 (N_3891,N_2693,N_2073);
xnor U3892 (N_3892,N_2411,N_2324);
xor U3893 (N_3893,N_2024,N_2764);
nor U3894 (N_3894,N_2058,N_2007);
nand U3895 (N_3895,N_2290,N_2379);
xor U3896 (N_3896,N_2832,N_2791);
xnor U3897 (N_3897,N_2066,N_2592);
nand U3898 (N_3898,N_2675,N_2152);
nor U3899 (N_3899,N_2871,N_2582);
nor U3900 (N_3900,N_2458,N_2966);
xor U3901 (N_3901,N_2838,N_2314);
nor U3902 (N_3902,N_2626,N_2751);
xnor U3903 (N_3903,N_2807,N_2687);
nand U3904 (N_3904,N_2906,N_2055);
and U3905 (N_3905,N_2278,N_2888);
xor U3906 (N_3906,N_2674,N_2383);
nor U3907 (N_3907,N_2783,N_2914);
nand U3908 (N_3908,N_2075,N_2038);
xor U3909 (N_3909,N_2955,N_2657);
xor U3910 (N_3910,N_2924,N_2012);
nor U3911 (N_3911,N_2047,N_2472);
nor U3912 (N_3912,N_2326,N_2783);
or U3913 (N_3913,N_2881,N_2233);
nand U3914 (N_3914,N_2652,N_2473);
and U3915 (N_3915,N_2445,N_2631);
or U3916 (N_3916,N_2489,N_2841);
or U3917 (N_3917,N_2052,N_2035);
nand U3918 (N_3918,N_2974,N_2378);
xor U3919 (N_3919,N_2236,N_2840);
or U3920 (N_3920,N_2914,N_2848);
xor U3921 (N_3921,N_2696,N_2076);
xnor U3922 (N_3922,N_2606,N_2071);
and U3923 (N_3923,N_2413,N_2901);
and U3924 (N_3924,N_2480,N_2019);
or U3925 (N_3925,N_2552,N_2081);
xnor U3926 (N_3926,N_2789,N_2111);
nand U3927 (N_3927,N_2399,N_2191);
or U3928 (N_3928,N_2208,N_2447);
and U3929 (N_3929,N_2082,N_2013);
and U3930 (N_3930,N_2007,N_2911);
xor U3931 (N_3931,N_2898,N_2220);
or U3932 (N_3932,N_2589,N_2252);
nand U3933 (N_3933,N_2098,N_2191);
or U3934 (N_3934,N_2138,N_2363);
or U3935 (N_3935,N_2334,N_2613);
or U3936 (N_3936,N_2916,N_2896);
xnor U3937 (N_3937,N_2117,N_2421);
or U3938 (N_3938,N_2722,N_2429);
nor U3939 (N_3939,N_2438,N_2663);
nand U3940 (N_3940,N_2100,N_2002);
nor U3941 (N_3941,N_2194,N_2554);
and U3942 (N_3942,N_2031,N_2304);
or U3943 (N_3943,N_2456,N_2873);
xnor U3944 (N_3944,N_2525,N_2836);
and U3945 (N_3945,N_2776,N_2042);
and U3946 (N_3946,N_2290,N_2775);
or U3947 (N_3947,N_2808,N_2478);
nor U3948 (N_3948,N_2540,N_2746);
xor U3949 (N_3949,N_2660,N_2017);
nand U3950 (N_3950,N_2028,N_2343);
and U3951 (N_3951,N_2763,N_2737);
and U3952 (N_3952,N_2088,N_2156);
or U3953 (N_3953,N_2557,N_2515);
nor U3954 (N_3954,N_2112,N_2412);
nand U3955 (N_3955,N_2194,N_2394);
nand U3956 (N_3956,N_2768,N_2006);
nor U3957 (N_3957,N_2177,N_2754);
nor U3958 (N_3958,N_2280,N_2960);
nor U3959 (N_3959,N_2482,N_2727);
xnor U3960 (N_3960,N_2405,N_2778);
xnor U3961 (N_3961,N_2608,N_2606);
xor U3962 (N_3962,N_2118,N_2028);
and U3963 (N_3963,N_2639,N_2513);
and U3964 (N_3964,N_2512,N_2672);
and U3965 (N_3965,N_2672,N_2781);
xor U3966 (N_3966,N_2750,N_2676);
xnor U3967 (N_3967,N_2597,N_2775);
nor U3968 (N_3968,N_2765,N_2759);
nor U3969 (N_3969,N_2377,N_2988);
or U3970 (N_3970,N_2126,N_2553);
xor U3971 (N_3971,N_2828,N_2204);
nand U3972 (N_3972,N_2605,N_2752);
or U3973 (N_3973,N_2958,N_2126);
xnor U3974 (N_3974,N_2740,N_2987);
xnor U3975 (N_3975,N_2572,N_2613);
nand U3976 (N_3976,N_2462,N_2347);
nor U3977 (N_3977,N_2851,N_2864);
and U3978 (N_3978,N_2815,N_2899);
and U3979 (N_3979,N_2349,N_2674);
and U3980 (N_3980,N_2830,N_2527);
nand U3981 (N_3981,N_2638,N_2589);
or U3982 (N_3982,N_2849,N_2108);
nand U3983 (N_3983,N_2483,N_2384);
or U3984 (N_3984,N_2467,N_2769);
xnor U3985 (N_3985,N_2204,N_2984);
xnor U3986 (N_3986,N_2421,N_2740);
xor U3987 (N_3987,N_2255,N_2739);
nor U3988 (N_3988,N_2994,N_2795);
xnor U3989 (N_3989,N_2177,N_2111);
or U3990 (N_3990,N_2410,N_2664);
xnor U3991 (N_3991,N_2040,N_2479);
and U3992 (N_3992,N_2574,N_2793);
nand U3993 (N_3993,N_2481,N_2384);
xor U3994 (N_3994,N_2498,N_2608);
and U3995 (N_3995,N_2867,N_2473);
and U3996 (N_3996,N_2059,N_2262);
and U3997 (N_3997,N_2929,N_2195);
nor U3998 (N_3998,N_2609,N_2315);
xor U3999 (N_3999,N_2209,N_2620);
nor U4000 (N_4000,N_3449,N_3018);
and U4001 (N_4001,N_3225,N_3993);
nor U4002 (N_4002,N_3618,N_3755);
and U4003 (N_4003,N_3948,N_3072);
xnor U4004 (N_4004,N_3375,N_3360);
xnor U4005 (N_4005,N_3278,N_3482);
nor U4006 (N_4006,N_3536,N_3147);
or U4007 (N_4007,N_3457,N_3281);
xnor U4008 (N_4008,N_3001,N_3363);
and U4009 (N_4009,N_3677,N_3878);
nor U4010 (N_4010,N_3953,N_3188);
and U4011 (N_4011,N_3686,N_3208);
xnor U4012 (N_4012,N_3101,N_3595);
or U4013 (N_4013,N_3582,N_3268);
nor U4014 (N_4014,N_3048,N_3136);
or U4015 (N_4015,N_3809,N_3507);
nor U4016 (N_4016,N_3213,N_3461);
nand U4017 (N_4017,N_3666,N_3726);
and U4018 (N_4018,N_3555,N_3608);
or U4019 (N_4019,N_3116,N_3504);
and U4020 (N_4020,N_3756,N_3763);
and U4021 (N_4021,N_3553,N_3391);
xor U4022 (N_4022,N_3509,N_3167);
and U4023 (N_4023,N_3826,N_3499);
and U4024 (N_4024,N_3532,N_3324);
xnor U4025 (N_4025,N_3660,N_3151);
nand U4026 (N_4026,N_3880,N_3096);
nor U4027 (N_4027,N_3684,N_3827);
nand U4028 (N_4028,N_3725,N_3359);
xor U4029 (N_4029,N_3970,N_3649);
nor U4030 (N_4030,N_3002,N_3577);
or U4031 (N_4031,N_3633,N_3697);
or U4032 (N_4032,N_3111,N_3205);
nor U4033 (N_4033,N_3495,N_3087);
and U4034 (N_4034,N_3169,N_3513);
xnor U4035 (N_4035,N_3635,N_3333);
nand U4036 (N_4036,N_3179,N_3837);
xnor U4037 (N_4037,N_3852,N_3855);
or U4038 (N_4038,N_3378,N_3645);
or U4039 (N_4039,N_3164,N_3185);
nand U4040 (N_4040,N_3551,N_3719);
nor U4041 (N_4041,N_3986,N_3815);
or U4042 (N_4042,N_3007,N_3424);
or U4043 (N_4043,N_3812,N_3266);
nor U4044 (N_4044,N_3610,N_3501);
nand U4045 (N_4045,N_3288,N_3983);
nor U4046 (N_4046,N_3958,N_3240);
xnor U4047 (N_4047,N_3506,N_3434);
or U4048 (N_4048,N_3286,N_3637);
or U4049 (N_4049,N_3956,N_3678);
xnor U4050 (N_4050,N_3881,N_3814);
or U4051 (N_4051,N_3023,N_3183);
xor U4052 (N_4052,N_3886,N_3828);
nand U4053 (N_4053,N_3954,N_3508);
and U4054 (N_4054,N_3031,N_3237);
nor U4055 (N_4055,N_3063,N_3847);
nor U4056 (N_4056,N_3831,N_3419);
nor U4057 (N_4057,N_3665,N_3123);
and U4058 (N_4058,N_3766,N_3634);
nand U4059 (N_4059,N_3918,N_3472);
or U4060 (N_4060,N_3068,N_3861);
or U4061 (N_4061,N_3190,N_3671);
and U4062 (N_4062,N_3284,N_3129);
nand U4063 (N_4063,N_3366,N_3061);
and U4064 (N_4064,N_3305,N_3247);
nand U4065 (N_4065,N_3309,N_3200);
xnor U4066 (N_4066,N_3965,N_3552);
nor U4067 (N_4067,N_3612,N_3028);
or U4068 (N_4068,N_3720,N_3590);
or U4069 (N_4069,N_3168,N_3897);
xor U4070 (N_4070,N_3148,N_3008);
or U4071 (N_4071,N_3891,N_3418);
xor U4072 (N_4072,N_3584,N_3734);
and U4073 (N_4073,N_3773,N_3193);
or U4074 (N_4074,N_3805,N_3331);
or U4075 (N_4075,N_3030,N_3664);
nand U4076 (N_4076,N_3176,N_3276);
nand U4077 (N_4077,N_3414,N_3682);
and U4078 (N_4078,N_3849,N_3848);
nand U4079 (N_4079,N_3264,N_3989);
and U4080 (N_4080,N_3067,N_3544);
nand U4081 (N_4081,N_3926,N_3298);
nand U4082 (N_4082,N_3561,N_3212);
or U4083 (N_4083,N_3013,N_3239);
xor U4084 (N_4084,N_3131,N_3026);
or U4085 (N_4085,N_3191,N_3708);
or U4086 (N_4086,N_3351,N_3250);
xor U4087 (N_4087,N_3079,N_3566);
nor U4088 (N_4088,N_3349,N_3877);
or U4089 (N_4089,N_3559,N_3905);
nand U4090 (N_4090,N_3711,N_3214);
nor U4091 (N_4091,N_3187,N_3384);
nor U4092 (N_4092,N_3489,N_3715);
and U4093 (N_4093,N_3174,N_3889);
nand U4094 (N_4094,N_3246,N_3476);
or U4095 (N_4095,N_3856,N_3862);
or U4096 (N_4096,N_3231,N_3177);
and U4097 (N_4097,N_3775,N_3710);
or U4098 (N_4098,N_3613,N_3153);
xnor U4099 (N_4099,N_3585,N_3735);
and U4100 (N_4100,N_3510,N_3640);
xnor U4101 (N_4101,N_3998,N_3873);
or U4102 (N_4102,N_3092,N_3841);
and U4103 (N_4103,N_3386,N_3497);
or U4104 (N_4104,N_3539,N_3235);
nor U4105 (N_4105,N_3394,N_3767);
or U4106 (N_4106,N_3738,N_3269);
nor U4107 (N_4107,N_3807,N_3337);
nand U4108 (N_4108,N_3620,N_3399);
xnor U4109 (N_4109,N_3749,N_3978);
xnor U4110 (N_4110,N_3003,N_3598);
and U4111 (N_4111,N_3854,N_3924);
or U4112 (N_4112,N_3084,N_3282);
nand U4113 (N_4113,N_3919,N_3724);
nand U4114 (N_4114,N_3939,N_3404);
or U4115 (N_4115,N_3059,N_3492);
nor U4116 (N_4116,N_3835,N_3938);
and U4117 (N_4117,N_3128,N_3731);
nand U4118 (N_4118,N_3690,N_3243);
nand U4119 (N_4119,N_3959,N_3599);
or U4120 (N_4120,N_3464,N_3152);
or U4121 (N_4121,N_3156,N_3011);
nand U4122 (N_4122,N_3853,N_3283);
nor U4123 (N_4123,N_3903,N_3244);
nand U4124 (N_4124,N_3935,N_3279);
nand U4125 (N_4125,N_3687,N_3103);
or U4126 (N_4126,N_3445,N_3803);
nand U4127 (N_4127,N_3933,N_3688);
or U4128 (N_4128,N_3535,N_3676);
nor U4129 (N_4129,N_3143,N_3727);
nor U4130 (N_4130,N_3981,N_3382);
nand U4131 (N_4131,N_3657,N_3440);
or U4132 (N_4132,N_3014,N_3203);
xnor U4133 (N_4133,N_3393,N_3703);
or U4134 (N_4134,N_3189,N_3651);
nor U4135 (N_4135,N_3516,N_3329);
and U4136 (N_4136,N_3844,N_3761);
nand U4137 (N_4137,N_3088,N_3549);
or U4138 (N_4138,N_3005,N_3994);
nor U4139 (N_4139,N_3291,N_3969);
xor U4140 (N_4140,N_3515,N_3452);
and U4141 (N_4141,N_3723,N_3916);
xor U4142 (N_4142,N_3209,N_3065);
or U4143 (N_4143,N_3460,N_3806);
and U4144 (N_4144,N_3811,N_3325);
nand U4145 (N_4145,N_3709,N_3304);
or U4146 (N_4146,N_3021,N_3721);
xnor U4147 (N_4147,N_3732,N_3217);
or U4148 (N_4148,N_3172,N_3348);
nor U4149 (N_4149,N_3303,N_3484);
or U4150 (N_4150,N_3318,N_3275);
nor U4151 (N_4151,N_3801,N_3915);
xor U4152 (N_4152,N_3797,N_3619);
xnor U4153 (N_4153,N_3597,N_3563);
xnor U4154 (N_4154,N_3421,N_3180);
xnor U4155 (N_4155,N_3019,N_3788);
nor U4156 (N_4156,N_3227,N_3796);
or U4157 (N_4157,N_3483,N_3471);
xor U4158 (N_4158,N_3262,N_3230);
xor U4159 (N_4159,N_3256,N_3140);
nor U4160 (N_4160,N_3373,N_3458);
nand U4161 (N_4161,N_3740,N_3494);
nor U4162 (N_4162,N_3794,N_3863);
xnor U4163 (N_4163,N_3338,N_3042);
nor U4164 (N_4164,N_3022,N_3545);
nand U4165 (N_4165,N_3611,N_3417);
or U4166 (N_4166,N_3737,N_3987);
or U4167 (N_4167,N_3783,N_3475);
nor U4168 (N_4168,N_3443,N_3255);
nor U4169 (N_4169,N_3564,N_3865);
nand U4170 (N_4170,N_3602,N_3940);
and U4171 (N_4171,N_3000,N_3631);
nor U4172 (N_4172,N_3742,N_3319);
xor U4173 (N_4173,N_3137,N_3377);
and U4174 (N_4174,N_3571,N_3728);
nor U4175 (N_4175,N_3789,N_3527);
and U4176 (N_4176,N_3330,N_3317);
nand U4177 (N_4177,N_3706,N_3656);
xor U4178 (N_4178,N_3301,N_3274);
nor U4179 (N_4179,N_3525,N_3692);
xnor U4180 (N_4180,N_3043,N_3114);
nand U4181 (N_4181,N_3748,N_3961);
nor U4182 (N_4182,N_3600,N_3874);
nor U4183 (N_4183,N_3952,N_3674);
or U4184 (N_4184,N_3922,N_3623);
xor U4185 (N_4185,N_3782,N_3477);
xor U4186 (N_4186,N_3966,N_3569);
xor U4187 (N_4187,N_3913,N_3923);
and U4188 (N_4188,N_3592,N_3292);
nor U4189 (N_4189,N_3699,N_3531);
xnor U4190 (N_4190,N_3523,N_3052);
nand U4191 (N_4191,N_3413,N_3166);
nor U4192 (N_4192,N_3354,N_3347);
xnor U4193 (N_4193,N_3265,N_3362);
or U4194 (N_4194,N_3219,N_3273);
or U4195 (N_4195,N_3197,N_3371);
nor U4196 (N_4196,N_3960,N_3696);
nor U4197 (N_4197,N_3066,N_3198);
xnor U4198 (N_4198,N_3132,N_3465);
nand U4199 (N_4199,N_3745,N_3270);
nand U4200 (N_4200,N_3834,N_3315);
nor U4201 (N_4201,N_3560,N_3636);
nor U4202 (N_4202,N_3558,N_3984);
xnor U4203 (N_4203,N_3943,N_3823);
and U4204 (N_4204,N_3448,N_3601);
nand U4205 (N_4205,N_3893,N_3397);
nand U4206 (N_4206,N_3327,N_3917);
and U4207 (N_4207,N_3647,N_3290);
xor U4208 (N_4208,N_3016,N_3914);
xnor U4209 (N_4209,N_3988,N_3175);
nand U4210 (N_4210,N_3937,N_3374);
nand U4211 (N_4211,N_3340,N_3381);
xor U4212 (N_4212,N_3196,N_3124);
and U4213 (N_4213,N_3125,N_3009);
and U4214 (N_4214,N_3260,N_3346);
nand U4215 (N_4215,N_3390,N_3236);
or U4216 (N_4216,N_3154,N_3353);
xnor U4217 (N_4217,N_3689,N_3867);
or U4218 (N_4218,N_3530,N_3102);
and U4219 (N_4219,N_3972,N_3357);
xnor U4220 (N_4220,N_3369,N_3929);
nor U4221 (N_4221,N_3479,N_3157);
and U4222 (N_4222,N_3053,N_3573);
xor U4223 (N_4223,N_3641,N_3866);
nand U4224 (N_4224,N_3964,N_3054);
nor U4225 (N_4225,N_3857,N_3076);
nor U4226 (N_4226,N_3947,N_3097);
or U4227 (N_4227,N_3086,N_3046);
nand U4228 (N_4228,N_3004,N_3928);
and U4229 (N_4229,N_3603,N_3580);
xnor U4230 (N_4230,N_3376,N_3522);
nor U4231 (N_4231,N_3769,N_3010);
and U4232 (N_4232,N_3765,N_3130);
nor U4233 (N_4233,N_3968,N_3077);
nand U4234 (N_4234,N_3594,N_3252);
nand U4235 (N_4235,N_3135,N_3578);
xor U4236 (N_4236,N_3163,N_3540);
nor U4237 (N_4237,N_3277,N_3342);
and U4238 (N_4238,N_3764,N_3034);
nor U4239 (N_4239,N_3436,N_3776);
nand U4240 (N_4240,N_3328,N_3502);
and U4241 (N_4241,N_3218,N_3165);
xor U4242 (N_4242,N_3757,N_3033);
nand U4243 (N_4243,N_3512,N_3316);
or U4244 (N_4244,N_3672,N_3659);
or U4245 (N_4245,N_3426,N_3473);
nor U4246 (N_4246,N_3155,N_3879);
xnor U4247 (N_4247,N_3120,N_3416);
xor U4248 (N_4248,N_3543,N_3907);
nand U4249 (N_4249,N_3693,N_3967);
and U4250 (N_4250,N_3184,N_3830);
and U4251 (N_4251,N_3463,N_3320);
nor U4252 (N_4252,N_3423,N_3712);
xnor U4253 (N_4253,N_3480,N_3661);
and U4254 (N_4254,N_3518,N_3220);
or U4255 (N_4255,N_3145,N_3127);
xor U4256 (N_4256,N_3704,N_3554);
or U4257 (N_4257,N_3985,N_3109);
or U4258 (N_4258,N_3846,N_3110);
nand U4259 (N_4259,N_3900,N_3596);
nor U4260 (N_4260,N_3833,N_3800);
xnor U4261 (N_4261,N_3071,N_3224);
and U4262 (N_4262,N_3950,N_3395);
or U4263 (N_4263,N_3838,N_3931);
nand U4264 (N_4264,N_3609,N_3272);
or U4265 (N_4265,N_3628,N_3468);
or U4266 (N_4266,N_3093,N_3367);
and U4267 (N_4267,N_3781,N_3158);
or U4268 (N_4268,N_3836,N_3379);
or U4269 (N_4269,N_3138,N_3344);
and U4270 (N_4270,N_3242,N_3817);
and U4271 (N_4271,N_3117,N_3029);
and U4272 (N_4272,N_3840,N_3717);
nand U4273 (N_4273,N_3149,N_3082);
xnor U4274 (N_4274,N_3352,N_3104);
nor U4275 (N_4275,N_3069,N_3562);
and U4276 (N_4276,N_3521,N_3420);
and U4277 (N_4277,N_3999,N_3181);
nor U4278 (N_4278,N_3744,N_3520);
and U4279 (N_4279,N_3868,N_3332);
or U4280 (N_4280,N_3245,N_3435);
and U4281 (N_4281,N_3334,N_3979);
nand U4282 (N_4282,N_3652,N_3750);
and U4283 (N_4283,N_3108,N_3977);
or U4284 (N_4284,N_3364,N_3779);
xor U4285 (N_4285,N_3056,N_3162);
or U4286 (N_4286,N_3695,N_3996);
nand U4287 (N_4287,N_3630,N_3410);
and U4288 (N_4288,N_3642,N_3751);
nand U4289 (N_4289,N_3997,N_3784);
nor U4290 (N_4290,N_3995,N_3466);
and U4291 (N_4291,N_3459,N_3538);
or U4292 (N_4292,N_3533,N_3112);
nand U4293 (N_4293,N_3300,N_3675);
xor U4294 (N_4294,N_3517,N_3622);
nor U4295 (N_4295,N_3505,N_3772);
or U4296 (N_4296,N_3429,N_3064);
nand U4297 (N_4297,N_3115,N_3790);
nand U4298 (N_4298,N_3638,N_3451);
and U4299 (N_4299,N_3040,N_3875);
nand U4300 (N_4300,N_3289,N_3850);
xor U4301 (N_4301,N_3644,N_3605);
or U4302 (N_4302,N_3144,N_3793);
and U4303 (N_4303,N_3439,N_3258);
and U4304 (N_4304,N_3643,N_3892);
nor U4305 (N_4305,N_3579,N_3430);
xor U4306 (N_4306,N_3894,N_3896);
or U4307 (N_4307,N_3139,N_3428);
and U4308 (N_4308,N_3588,N_3107);
or U4309 (N_4309,N_3752,N_3713);
nand U4310 (N_4310,N_3941,N_3982);
xnor U4311 (N_4311,N_3804,N_3780);
or U4312 (N_4312,N_3085,N_3587);
nand U4313 (N_4313,N_3350,N_3027);
xor U4314 (N_4314,N_3624,N_3910);
or U4315 (N_4315,N_3037,N_3795);
or U4316 (N_4316,N_3195,N_3670);
nor U4317 (N_4317,N_3658,N_3094);
and U4318 (N_4318,N_3625,N_3774);
nor U4319 (N_4319,N_3567,N_3146);
or U4320 (N_4320,N_3238,N_3669);
xor U4321 (N_4321,N_3741,N_3514);
nand U4322 (N_4322,N_3629,N_3639);
xor U4323 (N_4323,N_3528,N_3341);
nor U4324 (N_4324,N_3314,N_3075);
or U4325 (N_4325,N_3906,N_3911);
nand U4326 (N_4326,N_3422,N_3487);
nand U4327 (N_4327,N_3142,N_3621);
and U4328 (N_4328,N_3050,N_3663);
nor U4329 (N_4329,N_3100,N_3498);
xor U4330 (N_4330,N_3204,N_3051);
nand U4331 (N_4331,N_3589,N_3824);
nand U4332 (N_4332,N_3653,N_3486);
and U4333 (N_4333,N_3730,N_3470);
nand U4334 (N_4334,N_3973,N_3308);
and U4335 (N_4335,N_3488,N_3206);
or U4336 (N_4336,N_3326,N_3842);
nand U4337 (N_4337,N_3186,N_3261);
nor U4338 (N_4338,N_3716,N_3447);
nand U4339 (N_4339,N_3060,N_3141);
nor U4340 (N_4340,N_3032,N_3267);
xnor U4341 (N_4341,N_3234,N_3170);
xor U4342 (N_4342,N_3006,N_3872);
or U4343 (N_4343,N_3312,N_3078);
nand U4344 (N_4344,N_3839,N_3883);
and U4345 (N_4345,N_3223,N_3951);
nand U4346 (N_4346,N_3591,N_3182);
nand U4347 (N_4347,N_3388,N_3746);
or U4348 (N_4348,N_3932,N_3548);
nand U4349 (N_4349,N_3934,N_3581);
and U4350 (N_4350,N_3936,N_3882);
and U4351 (N_4351,N_3887,N_3792);
xnor U4352 (N_4352,N_3478,N_3098);
or U4353 (N_4353,N_3679,N_3869);
or U4354 (N_4354,N_3408,N_3524);
and U4355 (N_4355,N_3895,N_3285);
and U4356 (N_4356,N_3454,N_3899);
nor U4357 (N_4357,N_3074,N_3049);
and U4358 (N_4358,N_3925,N_3683);
xor U4359 (N_4359,N_3949,N_3758);
and U4360 (N_4360,N_3024,N_3118);
nand U4361 (N_4361,N_3534,N_3387);
xnor U4362 (N_4362,N_3963,N_3450);
and U4363 (N_4363,N_3930,N_3407);
nor U4364 (N_4364,N_3446,N_3992);
nor U4365 (N_4365,N_3015,N_3161);
nor U4366 (N_4366,N_3888,N_3550);
nand U4367 (N_4367,N_3062,N_3257);
and U4368 (N_4368,N_3248,N_3870);
or U4369 (N_4369,N_3485,N_3370);
or U4370 (N_4370,N_3226,N_3760);
or U4371 (N_4371,N_3798,N_3411);
and U4372 (N_4372,N_3680,N_3974);
nand U4373 (N_4373,N_3753,N_3747);
or U4374 (N_4374,N_3980,N_3705);
nand U4375 (N_4375,N_3576,N_3668);
nand U4376 (N_4376,N_3405,N_3770);
nor U4377 (N_4377,N_3380,N_3614);
or U4378 (N_4378,N_3392,N_3593);
and U4379 (N_4379,N_3462,N_3134);
nor U4380 (N_4380,N_3017,N_3080);
xor U4381 (N_4381,N_3047,N_3927);
and U4382 (N_4382,N_3481,N_3859);
nor U4383 (N_4383,N_3299,N_3171);
xor U4384 (N_4384,N_3133,N_3990);
nor U4385 (N_4385,N_3099,N_3648);
nand U4386 (N_4386,N_3339,N_3908);
or U4387 (N_4387,N_3718,N_3864);
xnor U4388 (N_4388,N_3105,N_3297);
xor U4389 (N_4389,N_3280,N_3194);
nand U4390 (N_4390,N_3920,N_3570);
and U4391 (N_4391,N_3012,N_3401);
and U4392 (N_4392,N_3041,N_3444);
xor U4393 (N_4393,N_3402,N_3490);
nand U4394 (N_4394,N_3736,N_3777);
and U4395 (N_4395,N_3909,N_3768);
and U4396 (N_4396,N_3091,N_3307);
or U4397 (N_4397,N_3372,N_3714);
and U4398 (N_4398,N_3229,N_3832);
xnor U4399 (N_4399,N_3568,N_3912);
or U4400 (N_4400,N_3627,N_3201);
or U4401 (N_4401,N_3890,N_3519);
and U4402 (N_4402,N_3150,N_3456);
nor U4403 (N_4403,N_3754,N_3119);
and U4404 (N_4404,N_3962,N_3415);
or U4405 (N_4405,N_3398,N_3762);
xnor U4406 (N_4406,N_3662,N_3921);
or U4407 (N_4407,N_3944,N_3356);
nor U4408 (N_4408,N_3607,N_3057);
and U4409 (N_4409,N_3843,N_3574);
and U4410 (N_4410,N_3361,N_3547);
xor U4411 (N_4411,N_3851,N_3210);
nor U4412 (N_4412,N_3400,N_3739);
xor U4413 (N_4413,N_3902,N_3722);
nand U4414 (N_4414,N_3083,N_3323);
xor U4415 (N_4415,N_3586,N_3432);
xnor U4416 (N_4416,N_3343,N_3442);
or U4417 (N_4417,N_3025,N_3496);
nand U4418 (N_4418,N_3813,N_3433);
and U4419 (N_4419,N_3691,N_3820);
or U4420 (N_4420,N_3787,N_3565);
nand U4421 (N_4421,N_3822,N_3336);
nor U4422 (N_4422,N_3606,N_3971);
or U4423 (N_4423,N_3073,N_3778);
nand U4424 (N_4424,N_3829,N_3310);
and U4425 (N_4425,N_3583,N_3816);
nor U4426 (N_4426,N_3694,N_3821);
and U4427 (N_4427,N_3808,N_3860);
xor U4428 (N_4428,N_3403,N_3311);
and U4429 (N_4429,N_3178,N_3385);
or U4430 (N_4430,N_3358,N_3654);
or U4431 (N_4431,N_3617,N_3898);
or U4432 (N_4432,N_3743,N_3626);
nor U4433 (N_4433,N_3904,N_3655);
nor U4434 (N_4434,N_3491,N_3058);
nand U4435 (N_4435,N_3529,N_3089);
or U4436 (N_4436,N_3556,N_3216);
nor U4437 (N_4437,N_3251,N_3818);
nor U4438 (N_4438,N_3975,N_3106);
nor U4439 (N_4439,N_3160,N_3045);
nand U4440 (N_4440,N_3035,N_3572);
and U4441 (N_4441,N_3557,N_3500);
nor U4442 (N_4442,N_3322,N_3537);
and U4443 (N_4443,N_3295,N_3791);
and U4444 (N_4444,N_3942,N_3474);
nand U4445 (N_4445,N_3700,N_3302);
nor U4446 (N_4446,N_3546,N_3173);
or U4447 (N_4447,N_3615,N_3876);
nand U4448 (N_4448,N_3228,N_3702);
or U4449 (N_4449,N_3389,N_3044);
nor U4450 (N_4450,N_3259,N_3222);
xor U4451 (N_4451,N_3232,N_3355);
xnor U4452 (N_4452,N_3604,N_3810);
nor U4453 (N_4453,N_3503,N_3294);
xor U4454 (N_4454,N_3122,N_3396);
xnor U4455 (N_4455,N_3365,N_3511);
and U4456 (N_4456,N_3667,N_3287);
nor U4457 (N_4457,N_3293,N_3254);
xnor U4458 (N_4458,N_3211,N_3453);
or U4459 (N_4459,N_3159,N_3202);
or U4460 (N_4460,N_3427,N_3090);
xor U4461 (N_4461,N_3406,N_3241);
and U4462 (N_4462,N_3575,N_3192);
and U4463 (N_4463,N_3802,N_3825);
or U4464 (N_4464,N_3976,N_3038);
or U4465 (N_4465,N_3707,N_3786);
nand U4466 (N_4466,N_3681,N_3345);
and U4467 (N_4467,N_3249,N_3113);
nor U4468 (N_4468,N_3271,N_3526);
or U4469 (N_4469,N_3207,N_3055);
nand U4470 (N_4470,N_3759,N_3785);
nand U4471 (N_4471,N_3884,N_3199);
xor U4472 (N_4472,N_3437,N_3215);
or U4473 (N_4473,N_3799,N_3221);
nor U4474 (N_4474,N_3039,N_3673);
nand U4475 (N_4475,N_3685,N_3126);
and U4476 (N_4476,N_3335,N_3296);
xnor U4477 (N_4477,N_3650,N_3493);
nand U4478 (N_4478,N_3646,N_3036);
and U4479 (N_4479,N_3306,N_3858);
nor U4480 (N_4480,N_3438,N_3431);
and U4481 (N_4481,N_3467,N_3819);
or U4482 (N_4482,N_3729,N_3542);
nor U4483 (N_4483,N_3901,N_3733);
xor U4484 (N_4484,N_3945,N_3946);
nand U4485 (N_4485,N_3409,N_3313);
nor U4486 (N_4486,N_3469,N_3233);
and U4487 (N_4487,N_3412,N_3701);
and U4488 (N_4488,N_3425,N_3441);
nand U4489 (N_4489,N_3698,N_3871);
nand U4490 (N_4490,N_3263,N_3632);
nand U4491 (N_4491,N_3455,N_3991);
nand U4492 (N_4492,N_3081,N_3383);
xnor U4493 (N_4493,N_3885,N_3095);
or U4494 (N_4494,N_3955,N_3616);
xor U4495 (N_4495,N_3541,N_3253);
and U4496 (N_4496,N_3845,N_3020);
nand U4497 (N_4497,N_3957,N_3070);
nor U4498 (N_4498,N_3771,N_3321);
xor U4499 (N_4499,N_3121,N_3368);
or U4500 (N_4500,N_3866,N_3501);
and U4501 (N_4501,N_3635,N_3585);
and U4502 (N_4502,N_3351,N_3520);
nand U4503 (N_4503,N_3433,N_3585);
nand U4504 (N_4504,N_3994,N_3021);
nand U4505 (N_4505,N_3715,N_3717);
or U4506 (N_4506,N_3089,N_3332);
nor U4507 (N_4507,N_3263,N_3380);
nand U4508 (N_4508,N_3092,N_3363);
or U4509 (N_4509,N_3714,N_3592);
nor U4510 (N_4510,N_3299,N_3687);
nor U4511 (N_4511,N_3953,N_3307);
and U4512 (N_4512,N_3773,N_3432);
nand U4513 (N_4513,N_3310,N_3080);
nor U4514 (N_4514,N_3321,N_3316);
or U4515 (N_4515,N_3101,N_3934);
or U4516 (N_4516,N_3811,N_3592);
nand U4517 (N_4517,N_3417,N_3268);
and U4518 (N_4518,N_3671,N_3540);
or U4519 (N_4519,N_3818,N_3520);
nor U4520 (N_4520,N_3659,N_3671);
nor U4521 (N_4521,N_3702,N_3477);
or U4522 (N_4522,N_3263,N_3576);
or U4523 (N_4523,N_3363,N_3483);
nand U4524 (N_4524,N_3979,N_3657);
and U4525 (N_4525,N_3512,N_3171);
or U4526 (N_4526,N_3635,N_3639);
xor U4527 (N_4527,N_3143,N_3921);
and U4528 (N_4528,N_3636,N_3816);
nand U4529 (N_4529,N_3287,N_3560);
and U4530 (N_4530,N_3533,N_3810);
and U4531 (N_4531,N_3478,N_3758);
and U4532 (N_4532,N_3789,N_3408);
xnor U4533 (N_4533,N_3715,N_3628);
and U4534 (N_4534,N_3197,N_3999);
xnor U4535 (N_4535,N_3846,N_3708);
nand U4536 (N_4536,N_3255,N_3412);
xor U4537 (N_4537,N_3661,N_3617);
nand U4538 (N_4538,N_3700,N_3828);
nand U4539 (N_4539,N_3648,N_3162);
or U4540 (N_4540,N_3534,N_3672);
xor U4541 (N_4541,N_3309,N_3323);
or U4542 (N_4542,N_3067,N_3988);
nand U4543 (N_4543,N_3562,N_3216);
or U4544 (N_4544,N_3342,N_3453);
nor U4545 (N_4545,N_3022,N_3151);
nor U4546 (N_4546,N_3585,N_3217);
xnor U4547 (N_4547,N_3547,N_3014);
nor U4548 (N_4548,N_3796,N_3581);
xor U4549 (N_4549,N_3849,N_3560);
nand U4550 (N_4550,N_3344,N_3204);
nor U4551 (N_4551,N_3006,N_3709);
nand U4552 (N_4552,N_3944,N_3238);
and U4553 (N_4553,N_3959,N_3703);
or U4554 (N_4554,N_3745,N_3198);
or U4555 (N_4555,N_3985,N_3369);
nand U4556 (N_4556,N_3357,N_3710);
nand U4557 (N_4557,N_3364,N_3763);
nand U4558 (N_4558,N_3566,N_3365);
nand U4559 (N_4559,N_3841,N_3733);
nor U4560 (N_4560,N_3230,N_3579);
nand U4561 (N_4561,N_3173,N_3926);
nand U4562 (N_4562,N_3732,N_3086);
xnor U4563 (N_4563,N_3771,N_3386);
or U4564 (N_4564,N_3621,N_3593);
xor U4565 (N_4565,N_3325,N_3789);
or U4566 (N_4566,N_3273,N_3926);
xnor U4567 (N_4567,N_3884,N_3652);
xnor U4568 (N_4568,N_3106,N_3356);
and U4569 (N_4569,N_3837,N_3825);
or U4570 (N_4570,N_3606,N_3328);
nand U4571 (N_4571,N_3635,N_3813);
xor U4572 (N_4572,N_3110,N_3709);
and U4573 (N_4573,N_3960,N_3726);
nor U4574 (N_4574,N_3008,N_3618);
and U4575 (N_4575,N_3113,N_3819);
nand U4576 (N_4576,N_3933,N_3859);
xor U4577 (N_4577,N_3437,N_3426);
xnor U4578 (N_4578,N_3325,N_3594);
or U4579 (N_4579,N_3825,N_3352);
or U4580 (N_4580,N_3825,N_3592);
xor U4581 (N_4581,N_3227,N_3113);
and U4582 (N_4582,N_3778,N_3821);
or U4583 (N_4583,N_3549,N_3628);
nor U4584 (N_4584,N_3595,N_3041);
xor U4585 (N_4585,N_3193,N_3765);
or U4586 (N_4586,N_3962,N_3849);
and U4587 (N_4587,N_3974,N_3872);
or U4588 (N_4588,N_3232,N_3059);
nand U4589 (N_4589,N_3917,N_3071);
nor U4590 (N_4590,N_3022,N_3179);
nor U4591 (N_4591,N_3867,N_3271);
xnor U4592 (N_4592,N_3718,N_3741);
xor U4593 (N_4593,N_3198,N_3310);
nor U4594 (N_4594,N_3111,N_3737);
and U4595 (N_4595,N_3251,N_3052);
nor U4596 (N_4596,N_3344,N_3820);
or U4597 (N_4597,N_3327,N_3158);
and U4598 (N_4598,N_3916,N_3779);
nand U4599 (N_4599,N_3722,N_3262);
or U4600 (N_4600,N_3617,N_3293);
or U4601 (N_4601,N_3434,N_3855);
and U4602 (N_4602,N_3742,N_3871);
nand U4603 (N_4603,N_3892,N_3389);
or U4604 (N_4604,N_3434,N_3123);
or U4605 (N_4605,N_3475,N_3580);
and U4606 (N_4606,N_3943,N_3054);
nand U4607 (N_4607,N_3589,N_3706);
nor U4608 (N_4608,N_3437,N_3229);
nor U4609 (N_4609,N_3884,N_3047);
nor U4610 (N_4610,N_3046,N_3344);
and U4611 (N_4611,N_3583,N_3725);
nand U4612 (N_4612,N_3124,N_3611);
nor U4613 (N_4613,N_3815,N_3720);
and U4614 (N_4614,N_3780,N_3859);
nand U4615 (N_4615,N_3432,N_3212);
nand U4616 (N_4616,N_3644,N_3476);
and U4617 (N_4617,N_3498,N_3564);
nand U4618 (N_4618,N_3092,N_3020);
nor U4619 (N_4619,N_3709,N_3536);
nor U4620 (N_4620,N_3868,N_3018);
nor U4621 (N_4621,N_3575,N_3228);
nor U4622 (N_4622,N_3428,N_3062);
xor U4623 (N_4623,N_3297,N_3729);
and U4624 (N_4624,N_3878,N_3200);
or U4625 (N_4625,N_3000,N_3202);
or U4626 (N_4626,N_3280,N_3283);
nor U4627 (N_4627,N_3675,N_3575);
nor U4628 (N_4628,N_3147,N_3533);
and U4629 (N_4629,N_3378,N_3865);
xor U4630 (N_4630,N_3635,N_3897);
xor U4631 (N_4631,N_3079,N_3594);
or U4632 (N_4632,N_3555,N_3716);
nor U4633 (N_4633,N_3412,N_3244);
nor U4634 (N_4634,N_3212,N_3166);
nand U4635 (N_4635,N_3930,N_3225);
or U4636 (N_4636,N_3184,N_3360);
or U4637 (N_4637,N_3824,N_3552);
nand U4638 (N_4638,N_3764,N_3576);
xnor U4639 (N_4639,N_3561,N_3443);
and U4640 (N_4640,N_3722,N_3808);
nor U4641 (N_4641,N_3541,N_3958);
xor U4642 (N_4642,N_3063,N_3563);
nor U4643 (N_4643,N_3771,N_3478);
nand U4644 (N_4644,N_3873,N_3235);
and U4645 (N_4645,N_3816,N_3024);
xnor U4646 (N_4646,N_3918,N_3200);
or U4647 (N_4647,N_3498,N_3133);
or U4648 (N_4648,N_3202,N_3899);
xnor U4649 (N_4649,N_3499,N_3870);
nor U4650 (N_4650,N_3630,N_3323);
and U4651 (N_4651,N_3304,N_3485);
and U4652 (N_4652,N_3480,N_3884);
and U4653 (N_4653,N_3972,N_3284);
xnor U4654 (N_4654,N_3376,N_3476);
xnor U4655 (N_4655,N_3231,N_3280);
xnor U4656 (N_4656,N_3849,N_3528);
xor U4657 (N_4657,N_3734,N_3853);
xor U4658 (N_4658,N_3336,N_3710);
nand U4659 (N_4659,N_3597,N_3566);
nand U4660 (N_4660,N_3956,N_3769);
nand U4661 (N_4661,N_3532,N_3591);
xor U4662 (N_4662,N_3315,N_3274);
or U4663 (N_4663,N_3945,N_3504);
nor U4664 (N_4664,N_3023,N_3051);
nand U4665 (N_4665,N_3138,N_3756);
and U4666 (N_4666,N_3228,N_3370);
and U4667 (N_4667,N_3377,N_3538);
nand U4668 (N_4668,N_3919,N_3058);
nand U4669 (N_4669,N_3785,N_3901);
or U4670 (N_4670,N_3772,N_3821);
xnor U4671 (N_4671,N_3040,N_3933);
or U4672 (N_4672,N_3381,N_3995);
or U4673 (N_4673,N_3059,N_3656);
nand U4674 (N_4674,N_3353,N_3947);
and U4675 (N_4675,N_3347,N_3653);
nor U4676 (N_4676,N_3182,N_3779);
nor U4677 (N_4677,N_3510,N_3278);
nor U4678 (N_4678,N_3605,N_3897);
nand U4679 (N_4679,N_3804,N_3923);
nand U4680 (N_4680,N_3123,N_3944);
nand U4681 (N_4681,N_3415,N_3565);
or U4682 (N_4682,N_3953,N_3331);
nor U4683 (N_4683,N_3921,N_3640);
nand U4684 (N_4684,N_3311,N_3600);
nand U4685 (N_4685,N_3085,N_3755);
and U4686 (N_4686,N_3608,N_3986);
xnor U4687 (N_4687,N_3924,N_3895);
nor U4688 (N_4688,N_3647,N_3630);
or U4689 (N_4689,N_3922,N_3919);
and U4690 (N_4690,N_3097,N_3746);
nand U4691 (N_4691,N_3497,N_3221);
or U4692 (N_4692,N_3265,N_3731);
and U4693 (N_4693,N_3517,N_3774);
xor U4694 (N_4694,N_3108,N_3853);
nand U4695 (N_4695,N_3557,N_3258);
and U4696 (N_4696,N_3552,N_3475);
xor U4697 (N_4697,N_3298,N_3101);
nand U4698 (N_4698,N_3047,N_3166);
and U4699 (N_4699,N_3210,N_3456);
nor U4700 (N_4700,N_3550,N_3820);
xnor U4701 (N_4701,N_3457,N_3367);
or U4702 (N_4702,N_3548,N_3442);
and U4703 (N_4703,N_3742,N_3327);
or U4704 (N_4704,N_3988,N_3386);
nor U4705 (N_4705,N_3187,N_3588);
and U4706 (N_4706,N_3614,N_3581);
and U4707 (N_4707,N_3437,N_3519);
xor U4708 (N_4708,N_3290,N_3249);
or U4709 (N_4709,N_3780,N_3638);
nand U4710 (N_4710,N_3493,N_3527);
xor U4711 (N_4711,N_3533,N_3305);
xnor U4712 (N_4712,N_3175,N_3753);
nor U4713 (N_4713,N_3833,N_3404);
or U4714 (N_4714,N_3160,N_3379);
or U4715 (N_4715,N_3418,N_3421);
and U4716 (N_4716,N_3232,N_3172);
or U4717 (N_4717,N_3709,N_3452);
nand U4718 (N_4718,N_3621,N_3614);
xnor U4719 (N_4719,N_3318,N_3256);
or U4720 (N_4720,N_3198,N_3813);
or U4721 (N_4721,N_3582,N_3524);
or U4722 (N_4722,N_3240,N_3851);
nor U4723 (N_4723,N_3201,N_3933);
xnor U4724 (N_4724,N_3842,N_3235);
nor U4725 (N_4725,N_3875,N_3013);
nand U4726 (N_4726,N_3883,N_3756);
nor U4727 (N_4727,N_3488,N_3708);
nand U4728 (N_4728,N_3332,N_3740);
or U4729 (N_4729,N_3059,N_3010);
xor U4730 (N_4730,N_3644,N_3278);
and U4731 (N_4731,N_3580,N_3793);
xnor U4732 (N_4732,N_3524,N_3748);
or U4733 (N_4733,N_3651,N_3778);
nor U4734 (N_4734,N_3266,N_3045);
nor U4735 (N_4735,N_3552,N_3746);
nand U4736 (N_4736,N_3878,N_3165);
or U4737 (N_4737,N_3983,N_3381);
xor U4738 (N_4738,N_3227,N_3373);
xor U4739 (N_4739,N_3910,N_3781);
or U4740 (N_4740,N_3651,N_3586);
nand U4741 (N_4741,N_3238,N_3319);
or U4742 (N_4742,N_3198,N_3444);
nor U4743 (N_4743,N_3625,N_3893);
or U4744 (N_4744,N_3622,N_3998);
nor U4745 (N_4745,N_3702,N_3845);
and U4746 (N_4746,N_3851,N_3133);
or U4747 (N_4747,N_3060,N_3198);
nand U4748 (N_4748,N_3685,N_3902);
nand U4749 (N_4749,N_3502,N_3106);
or U4750 (N_4750,N_3124,N_3110);
nor U4751 (N_4751,N_3580,N_3440);
nor U4752 (N_4752,N_3457,N_3825);
nor U4753 (N_4753,N_3563,N_3421);
nor U4754 (N_4754,N_3919,N_3796);
nand U4755 (N_4755,N_3021,N_3174);
or U4756 (N_4756,N_3331,N_3292);
nand U4757 (N_4757,N_3981,N_3834);
nand U4758 (N_4758,N_3795,N_3504);
nor U4759 (N_4759,N_3263,N_3804);
or U4760 (N_4760,N_3475,N_3258);
and U4761 (N_4761,N_3348,N_3819);
nand U4762 (N_4762,N_3877,N_3087);
and U4763 (N_4763,N_3291,N_3159);
and U4764 (N_4764,N_3660,N_3432);
xnor U4765 (N_4765,N_3762,N_3710);
or U4766 (N_4766,N_3131,N_3499);
nand U4767 (N_4767,N_3131,N_3976);
or U4768 (N_4768,N_3303,N_3642);
nor U4769 (N_4769,N_3420,N_3996);
and U4770 (N_4770,N_3045,N_3945);
xnor U4771 (N_4771,N_3225,N_3037);
and U4772 (N_4772,N_3883,N_3367);
and U4773 (N_4773,N_3385,N_3068);
xnor U4774 (N_4774,N_3771,N_3876);
nand U4775 (N_4775,N_3940,N_3142);
xor U4776 (N_4776,N_3537,N_3814);
nor U4777 (N_4777,N_3309,N_3317);
and U4778 (N_4778,N_3865,N_3311);
xnor U4779 (N_4779,N_3009,N_3091);
nand U4780 (N_4780,N_3340,N_3136);
and U4781 (N_4781,N_3470,N_3885);
nor U4782 (N_4782,N_3197,N_3200);
nand U4783 (N_4783,N_3435,N_3686);
or U4784 (N_4784,N_3412,N_3754);
nand U4785 (N_4785,N_3527,N_3627);
or U4786 (N_4786,N_3201,N_3365);
nor U4787 (N_4787,N_3175,N_3324);
nand U4788 (N_4788,N_3613,N_3282);
xor U4789 (N_4789,N_3790,N_3957);
xor U4790 (N_4790,N_3416,N_3186);
or U4791 (N_4791,N_3320,N_3365);
or U4792 (N_4792,N_3093,N_3285);
nand U4793 (N_4793,N_3739,N_3257);
and U4794 (N_4794,N_3112,N_3669);
or U4795 (N_4795,N_3754,N_3880);
or U4796 (N_4796,N_3504,N_3977);
nor U4797 (N_4797,N_3559,N_3451);
or U4798 (N_4798,N_3702,N_3137);
nand U4799 (N_4799,N_3219,N_3323);
and U4800 (N_4800,N_3782,N_3903);
nand U4801 (N_4801,N_3298,N_3151);
or U4802 (N_4802,N_3519,N_3939);
nand U4803 (N_4803,N_3363,N_3946);
nor U4804 (N_4804,N_3585,N_3041);
xor U4805 (N_4805,N_3300,N_3309);
and U4806 (N_4806,N_3814,N_3740);
xnor U4807 (N_4807,N_3281,N_3441);
xnor U4808 (N_4808,N_3299,N_3573);
nor U4809 (N_4809,N_3374,N_3654);
nand U4810 (N_4810,N_3206,N_3389);
and U4811 (N_4811,N_3174,N_3198);
xnor U4812 (N_4812,N_3402,N_3400);
or U4813 (N_4813,N_3450,N_3430);
or U4814 (N_4814,N_3019,N_3654);
and U4815 (N_4815,N_3214,N_3821);
nor U4816 (N_4816,N_3896,N_3757);
nor U4817 (N_4817,N_3310,N_3966);
and U4818 (N_4818,N_3130,N_3308);
nor U4819 (N_4819,N_3642,N_3162);
xnor U4820 (N_4820,N_3823,N_3571);
or U4821 (N_4821,N_3504,N_3350);
and U4822 (N_4822,N_3805,N_3131);
or U4823 (N_4823,N_3799,N_3192);
or U4824 (N_4824,N_3765,N_3150);
nor U4825 (N_4825,N_3389,N_3222);
and U4826 (N_4826,N_3445,N_3179);
and U4827 (N_4827,N_3625,N_3340);
and U4828 (N_4828,N_3280,N_3344);
nand U4829 (N_4829,N_3928,N_3283);
nor U4830 (N_4830,N_3052,N_3491);
nand U4831 (N_4831,N_3537,N_3556);
nand U4832 (N_4832,N_3414,N_3464);
nand U4833 (N_4833,N_3598,N_3617);
nand U4834 (N_4834,N_3780,N_3070);
xnor U4835 (N_4835,N_3042,N_3395);
nor U4836 (N_4836,N_3817,N_3227);
or U4837 (N_4837,N_3819,N_3674);
and U4838 (N_4838,N_3772,N_3874);
or U4839 (N_4839,N_3974,N_3141);
nand U4840 (N_4840,N_3755,N_3429);
nand U4841 (N_4841,N_3037,N_3657);
or U4842 (N_4842,N_3187,N_3912);
or U4843 (N_4843,N_3282,N_3296);
nand U4844 (N_4844,N_3202,N_3200);
nor U4845 (N_4845,N_3474,N_3652);
or U4846 (N_4846,N_3802,N_3641);
xor U4847 (N_4847,N_3229,N_3212);
or U4848 (N_4848,N_3790,N_3395);
or U4849 (N_4849,N_3286,N_3806);
nand U4850 (N_4850,N_3028,N_3153);
xnor U4851 (N_4851,N_3099,N_3137);
or U4852 (N_4852,N_3718,N_3790);
xor U4853 (N_4853,N_3238,N_3492);
or U4854 (N_4854,N_3818,N_3914);
and U4855 (N_4855,N_3517,N_3358);
nand U4856 (N_4856,N_3681,N_3093);
xor U4857 (N_4857,N_3660,N_3597);
nor U4858 (N_4858,N_3189,N_3495);
or U4859 (N_4859,N_3919,N_3390);
and U4860 (N_4860,N_3730,N_3458);
nand U4861 (N_4861,N_3673,N_3259);
nor U4862 (N_4862,N_3552,N_3698);
and U4863 (N_4863,N_3362,N_3445);
and U4864 (N_4864,N_3367,N_3319);
nor U4865 (N_4865,N_3904,N_3338);
and U4866 (N_4866,N_3393,N_3578);
nor U4867 (N_4867,N_3943,N_3016);
or U4868 (N_4868,N_3340,N_3837);
or U4869 (N_4869,N_3266,N_3472);
and U4870 (N_4870,N_3440,N_3894);
nand U4871 (N_4871,N_3534,N_3295);
nor U4872 (N_4872,N_3109,N_3326);
xnor U4873 (N_4873,N_3748,N_3409);
and U4874 (N_4874,N_3782,N_3617);
nand U4875 (N_4875,N_3100,N_3840);
and U4876 (N_4876,N_3160,N_3872);
and U4877 (N_4877,N_3006,N_3968);
nand U4878 (N_4878,N_3505,N_3682);
or U4879 (N_4879,N_3841,N_3144);
xnor U4880 (N_4880,N_3971,N_3740);
or U4881 (N_4881,N_3653,N_3176);
and U4882 (N_4882,N_3515,N_3375);
xnor U4883 (N_4883,N_3536,N_3661);
nand U4884 (N_4884,N_3273,N_3081);
nor U4885 (N_4885,N_3820,N_3618);
nor U4886 (N_4886,N_3606,N_3676);
and U4887 (N_4887,N_3151,N_3471);
nor U4888 (N_4888,N_3901,N_3051);
nor U4889 (N_4889,N_3776,N_3574);
nor U4890 (N_4890,N_3286,N_3480);
nor U4891 (N_4891,N_3992,N_3813);
or U4892 (N_4892,N_3110,N_3241);
nand U4893 (N_4893,N_3858,N_3466);
or U4894 (N_4894,N_3803,N_3887);
nor U4895 (N_4895,N_3309,N_3515);
nand U4896 (N_4896,N_3399,N_3132);
nor U4897 (N_4897,N_3723,N_3730);
and U4898 (N_4898,N_3632,N_3888);
nor U4899 (N_4899,N_3783,N_3645);
nor U4900 (N_4900,N_3869,N_3306);
nand U4901 (N_4901,N_3959,N_3414);
nand U4902 (N_4902,N_3314,N_3087);
and U4903 (N_4903,N_3690,N_3128);
and U4904 (N_4904,N_3964,N_3983);
nand U4905 (N_4905,N_3335,N_3378);
xor U4906 (N_4906,N_3500,N_3492);
nor U4907 (N_4907,N_3768,N_3941);
nand U4908 (N_4908,N_3589,N_3556);
or U4909 (N_4909,N_3156,N_3104);
nor U4910 (N_4910,N_3760,N_3040);
and U4911 (N_4911,N_3767,N_3617);
xnor U4912 (N_4912,N_3301,N_3837);
nor U4913 (N_4913,N_3019,N_3094);
nand U4914 (N_4914,N_3187,N_3281);
or U4915 (N_4915,N_3108,N_3911);
nor U4916 (N_4916,N_3247,N_3780);
nor U4917 (N_4917,N_3172,N_3952);
nor U4918 (N_4918,N_3537,N_3237);
xnor U4919 (N_4919,N_3019,N_3877);
xor U4920 (N_4920,N_3161,N_3396);
nand U4921 (N_4921,N_3280,N_3368);
xnor U4922 (N_4922,N_3855,N_3507);
xnor U4923 (N_4923,N_3359,N_3447);
and U4924 (N_4924,N_3319,N_3031);
xor U4925 (N_4925,N_3177,N_3976);
or U4926 (N_4926,N_3599,N_3062);
nand U4927 (N_4927,N_3948,N_3760);
nand U4928 (N_4928,N_3664,N_3244);
nor U4929 (N_4929,N_3939,N_3211);
nand U4930 (N_4930,N_3942,N_3259);
or U4931 (N_4931,N_3237,N_3616);
xnor U4932 (N_4932,N_3668,N_3902);
and U4933 (N_4933,N_3062,N_3767);
or U4934 (N_4934,N_3414,N_3234);
and U4935 (N_4935,N_3532,N_3076);
nor U4936 (N_4936,N_3995,N_3490);
xor U4937 (N_4937,N_3815,N_3923);
nor U4938 (N_4938,N_3018,N_3174);
xor U4939 (N_4939,N_3510,N_3592);
nor U4940 (N_4940,N_3552,N_3386);
or U4941 (N_4941,N_3598,N_3300);
nand U4942 (N_4942,N_3728,N_3113);
or U4943 (N_4943,N_3930,N_3935);
xor U4944 (N_4944,N_3341,N_3110);
and U4945 (N_4945,N_3167,N_3388);
xnor U4946 (N_4946,N_3982,N_3803);
nand U4947 (N_4947,N_3211,N_3402);
and U4948 (N_4948,N_3183,N_3978);
nor U4949 (N_4949,N_3964,N_3579);
nand U4950 (N_4950,N_3609,N_3995);
nor U4951 (N_4951,N_3831,N_3168);
or U4952 (N_4952,N_3145,N_3642);
nor U4953 (N_4953,N_3870,N_3413);
nor U4954 (N_4954,N_3014,N_3726);
xnor U4955 (N_4955,N_3739,N_3653);
or U4956 (N_4956,N_3163,N_3475);
nand U4957 (N_4957,N_3218,N_3321);
nor U4958 (N_4958,N_3086,N_3325);
nor U4959 (N_4959,N_3625,N_3313);
nand U4960 (N_4960,N_3873,N_3784);
nor U4961 (N_4961,N_3000,N_3325);
nor U4962 (N_4962,N_3943,N_3100);
nand U4963 (N_4963,N_3832,N_3670);
and U4964 (N_4964,N_3357,N_3247);
and U4965 (N_4965,N_3138,N_3671);
and U4966 (N_4966,N_3213,N_3446);
or U4967 (N_4967,N_3640,N_3332);
and U4968 (N_4968,N_3232,N_3425);
nor U4969 (N_4969,N_3673,N_3230);
xnor U4970 (N_4970,N_3204,N_3488);
and U4971 (N_4971,N_3064,N_3375);
nand U4972 (N_4972,N_3623,N_3187);
xor U4973 (N_4973,N_3386,N_3378);
or U4974 (N_4974,N_3208,N_3868);
or U4975 (N_4975,N_3692,N_3026);
nor U4976 (N_4976,N_3091,N_3892);
nand U4977 (N_4977,N_3448,N_3836);
and U4978 (N_4978,N_3939,N_3244);
xor U4979 (N_4979,N_3880,N_3862);
and U4980 (N_4980,N_3787,N_3090);
xnor U4981 (N_4981,N_3737,N_3786);
nor U4982 (N_4982,N_3420,N_3877);
or U4983 (N_4983,N_3198,N_3464);
and U4984 (N_4984,N_3541,N_3424);
nand U4985 (N_4985,N_3109,N_3278);
nor U4986 (N_4986,N_3989,N_3132);
xor U4987 (N_4987,N_3468,N_3940);
nor U4988 (N_4988,N_3419,N_3727);
nor U4989 (N_4989,N_3605,N_3336);
nor U4990 (N_4990,N_3676,N_3414);
nor U4991 (N_4991,N_3320,N_3098);
nor U4992 (N_4992,N_3866,N_3414);
nor U4993 (N_4993,N_3339,N_3137);
nor U4994 (N_4994,N_3660,N_3030);
xnor U4995 (N_4995,N_3593,N_3151);
nor U4996 (N_4996,N_3920,N_3697);
and U4997 (N_4997,N_3750,N_3722);
or U4998 (N_4998,N_3746,N_3792);
nor U4999 (N_4999,N_3386,N_3135);
xnor UO_0 (O_0,N_4509,N_4818);
xor UO_1 (O_1,N_4079,N_4354);
xnor UO_2 (O_2,N_4291,N_4199);
nor UO_3 (O_3,N_4853,N_4062);
xnor UO_4 (O_4,N_4102,N_4901);
nor UO_5 (O_5,N_4266,N_4182);
nand UO_6 (O_6,N_4369,N_4116);
nand UO_7 (O_7,N_4977,N_4074);
nand UO_8 (O_8,N_4540,N_4181);
or UO_9 (O_9,N_4944,N_4472);
xnor UO_10 (O_10,N_4248,N_4159);
nand UO_11 (O_11,N_4920,N_4841);
or UO_12 (O_12,N_4714,N_4255);
xor UO_13 (O_13,N_4355,N_4249);
and UO_14 (O_14,N_4748,N_4707);
or UO_15 (O_15,N_4769,N_4389);
and UO_16 (O_16,N_4857,N_4398);
and UO_17 (O_17,N_4084,N_4782);
or UO_18 (O_18,N_4980,N_4987);
nand UO_19 (O_19,N_4912,N_4361);
nor UO_20 (O_20,N_4597,N_4542);
nor UO_21 (O_21,N_4646,N_4424);
nand UO_22 (O_22,N_4059,N_4170);
or UO_23 (O_23,N_4712,N_4340);
and UO_24 (O_24,N_4497,N_4185);
xnor UO_25 (O_25,N_4594,N_4531);
nand UO_26 (O_26,N_4871,N_4191);
nor UO_27 (O_27,N_4907,N_4690);
nor UO_28 (O_28,N_4023,N_4022);
and UO_29 (O_29,N_4534,N_4789);
or UO_30 (O_30,N_4142,N_4358);
or UO_31 (O_31,N_4109,N_4587);
nor UO_32 (O_32,N_4458,N_4283);
nor UO_33 (O_33,N_4858,N_4034);
xor UO_34 (O_34,N_4824,N_4021);
xnor UO_35 (O_35,N_4563,N_4918);
or UO_36 (O_36,N_4590,N_4156);
and UO_37 (O_37,N_4125,N_4719);
and UO_38 (O_38,N_4866,N_4219);
nor UO_39 (O_39,N_4019,N_4722);
nor UO_40 (O_40,N_4588,N_4864);
or UO_41 (O_41,N_4049,N_4263);
xnor UO_42 (O_42,N_4585,N_4682);
or UO_43 (O_43,N_4392,N_4859);
xnor UO_44 (O_44,N_4038,N_4881);
xnor UO_45 (O_45,N_4295,N_4578);
xor UO_46 (O_46,N_4231,N_4478);
xnor UO_47 (O_47,N_4727,N_4952);
and UO_48 (O_48,N_4670,N_4121);
and UO_49 (O_49,N_4312,N_4289);
and UO_50 (O_50,N_4026,N_4851);
and UO_51 (O_51,N_4042,N_4272);
nor UO_52 (O_52,N_4891,N_4463);
or UO_53 (O_53,N_4758,N_4954);
nor UO_54 (O_54,N_4568,N_4604);
xnor UO_55 (O_55,N_4147,N_4308);
nand UO_56 (O_56,N_4047,N_4090);
xnor UO_57 (O_57,N_4802,N_4091);
or UO_58 (O_58,N_4650,N_4676);
or UO_59 (O_59,N_4574,N_4486);
or UO_60 (O_60,N_4469,N_4518);
and UO_61 (O_61,N_4564,N_4737);
xor UO_62 (O_62,N_4488,N_4167);
and UO_63 (O_63,N_4257,N_4838);
nand UO_64 (O_64,N_4002,N_4755);
or UO_65 (O_65,N_4601,N_4775);
nand UO_66 (O_66,N_4797,N_4559);
or UO_67 (O_67,N_4863,N_4467);
xnor UO_68 (O_68,N_4697,N_4400);
or UO_69 (O_69,N_4583,N_4897);
nor UO_70 (O_70,N_4967,N_4784);
nor UO_71 (O_71,N_4211,N_4732);
or UO_72 (O_72,N_4834,N_4452);
xnor UO_73 (O_73,N_4081,N_4527);
or UO_74 (O_74,N_4155,N_4430);
or UO_75 (O_75,N_4652,N_4082);
or UO_76 (O_76,N_4875,N_4058);
nand UO_77 (O_77,N_4311,N_4238);
nand UO_78 (O_78,N_4489,N_4404);
and UO_79 (O_79,N_4649,N_4305);
nor UO_80 (O_80,N_4036,N_4947);
nand UO_81 (O_81,N_4966,N_4625);
xnor UO_82 (O_82,N_4150,N_4425);
xor UO_83 (O_83,N_4158,N_4414);
nor UO_84 (O_84,N_4213,N_4339);
nor UO_85 (O_85,N_4696,N_4270);
nor UO_86 (O_86,N_4229,N_4504);
or UO_87 (O_87,N_4956,N_4938);
nor UO_88 (O_88,N_4247,N_4940);
xor UO_89 (O_89,N_4485,N_4888);
nor UO_90 (O_90,N_4762,N_4456);
or UO_91 (O_91,N_4661,N_4372);
or UO_92 (O_92,N_4974,N_4324);
nand UO_93 (O_93,N_4576,N_4029);
xnor UO_94 (O_94,N_4613,N_4362);
nand UO_95 (O_95,N_4055,N_4950);
or UO_96 (O_96,N_4936,N_4939);
xor UO_97 (O_97,N_4522,N_4922);
nand UO_98 (O_98,N_4256,N_4344);
or UO_99 (O_99,N_4970,N_4284);
nor UO_100 (O_100,N_4179,N_4865);
nand UO_101 (O_101,N_4525,N_4387);
nand UO_102 (O_102,N_4268,N_4910);
and UO_103 (O_103,N_4551,N_4862);
or UO_104 (O_104,N_4635,N_4243);
and UO_105 (O_105,N_4433,N_4288);
or UO_106 (O_106,N_4890,N_4196);
xnor UO_107 (O_107,N_4946,N_4629);
xor UO_108 (O_108,N_4589,N_4602);
nor UO_109 (O_109,N_4795,N_4868);
nor UO_110 (O_110,N_4796,N_4064);
and UO_111 (O_111,N_4989,N_4407);
nand UO_112 (O_112,N_4253,N_4069);
xor UO_113 (O_113,N_4276,N_4207);
xnor UO_114 (O_114,N_4929,N_4086);
or UO_115 (O_115,N_4931,N_4020);
nand UO_116 (O_116,N_4442,N_4087);
or UO_117 (O_117,N_4450,N_4097);
nand UO_118 (O_118,N_4208,N_4605);
nand UO_119 (O_119,N_4935,N_4490);
nand UO_120 (O_120,N_4837,N_4892);
nor UO_121 (O_121,N_4790,N_4018);
nor UO_122 (O_122,N_4473,N_4379);
nand UO_123 (O_123,N_4814,N_4454);
nor UO_124 (O_124,N_4043,N_4048);
nor UO_125 (O_125,N_4607,N_4012);
nand UO_126 (O_126,N_4135,N_4927);
xor UO_127 (O_127,N_4730,N_4318);
or UO_128 (O_128,N_4129,N_4298);
xnor UO_129 (O_129,N_4076,N_4752);
or UO_130 (O_130,N_4330,N_4130);
xnor UO_131 (O_131,N_4511,N_4742);
nand UO_132 (O_132,N_4582,N_4500);
and UO_133 (O_133,N_4981,N_4721);
xor UO_134 (O_134,N_4827,N_4329);
nor UO_135 (O_135,N_4679,N_4390);
nand UO_136 (O_136,N_4612,N_4005);
and UO_137 (O_137,N_4325,N_4152);
xor UO_138 (O_138,N_4346,N_4523);
nand UO_139 (O_139,N_4193,N_4338);
or UO_140 (O_140,N_4861,N_4111);
nor UO_141 (O_141,N_4112,N_4376);
nor UO_142 (O_142,N_4971,N_4239);
nor UO_143 (O_143,N_4725,N_4225);
xor UO_144 (O_144,N_4184,N_4320);
xnor UO_145 (O_145,N_4519,N_4555);
nand UO_146 (O_146,N_4495,N_4009);
xor UO_147 (O_147,N_4416,N_4406);
nand UO_148 (O_148,N_4530,N_4529);
nand UO_149 (O_149,N_4774,N_4403);
xnor UO_150 (O_150,N_4835,N_4878);
xnor UO_151 (O_151,N_4615,N_4764);
or UO_152 (O_152,N_4139,N_4687);
xor UO_153 (O_153,N_4746,N_4089);
nand UO_154 (O_154,N_4672,N_4429);
nand UO_155 (O_155,N_4842,N_4335);
nor UO_156 (O_156,N_4397,N_4261);
and UO_157 (O_157,N_4506,N_4412);
nand UO_158 (O_158,N_4505,N_4264);
nor UO_159 (O_159,N_4538,N_4848);
nor UO_160 (O_160,N_4304,N_4805);
and UO_161 (O_161,N_4877,N_4095);
nand UO_162 (O_162,N_4075,N_4846);
nor UO_163 (O_163,N_4080,N_4516);
nand UO_164 (O_164,N_4294,N_4117);
nand UO_165 (O_165,N_4665,N_4259);
nand UO_166 (O_166,N_4777,N_4826);
nand UO_167 (O_167,N_4809,N_4356);
and UO_168 (O_168,N_4819,N_4290);
and UO_169 (O_169,N_4203,N_4926);
nand UO_170 (O_170,N_4694,N_4017);
and UO_171 (O_171,N_4114,N_4278);
or UO_172 (O_172,N_4209,N_4180);
nor UO_173 (O_173,N_4514,N_4681);
nor UO_174 (O_174,N_4894,N_4919);
or UO_175 (O_175,N_4385,N_4183);
nor UO_176 (O_176,N_4526,N_4711);
nand UO_177 (O_177,N_4065,N_4508);
nand UO_178 (O_178,N_4380,N_4071);
xor UO_179 (O_179,N_4874,N_4146);
or UO_180 (O_180,N_4566,N_4083);
and UO_181 (O_181,N_4422,N_4098);
nand UO_182 (O_182,N_4680,N_4134);
and UO_183 (O_183,N_4991,N_4833);
or UO_184 (O_184,N_4177,N_4492);
xnor UO_185 (O_185,N_4993,N_4787);
and UO_186 (O_186,N_4749,N_4695);
and UO_187 (O_187,N_4924,N_4448);
or UO_188 (O_188,N_4713,N_4241);
nand UO_189 (O_189,N_4963,N_4767);
xnor UO_190 (O_190,N_4381,N_4364);
and UO_191 (O_191,N_4623,N_4337);
and UO_192 (O_192,N_4378,N_4148);
nor UO_193 (O_193,N_4197,N_4475);
or UO_194 (O_194,N_4157,N_4621);
xnor UO_195 (O_195,N_4024,N_4326);
nor UO_196 (O_196,N_4192,N_4353);
xnor UO_197 (O_197,N_4915,N_4303);
nand UO_198 (O_198,N_4393,N_4011);
or UO_199 (O_199,N_4194,N_4474);
or UO_200 (O_200,N_4128,N_4648);
nor UO_201 (O_201,N_4739,N_4908);
nand UO_202 (O_202,N_4960,N_4446);
or UO_203 (O_203,N_4759,N_4836);
or UO_204 (O_204,N_4973,N_4724);
or UO_205 (O_205,N_4662,N_4427);
and UO_206 (O_206,N_4360,N_4396);
xnor UO_207 (O_207,N_4245,N_4060);
xnor UO_208 (O_208,N_4198,N_4321);
nor UO_209 (O_209,N_4479,N_4934);
nor UO_210 (O_210,N_4549,N_4914);
xor UO_211 (O_211,N_4778,N_4124);
xnor UO_212 (O_212,N_4840,N_4046);
nor UO_213 (O_213,N_4483,N_4898);
or UO_214 (O_214,N_4120,N_4743);
or UO_215 (O_215,N_4258,N_4013);
and UO_216 (O_216,N_4410,N_4375);
and UO_217 (O_217,N_4791,N_4738);
nor UO_218 (O_218,N_4131,N_4078);
and UO_219 (O_219,N_4773,N_4668);
and UO_220 (O_220,N_4384,N_4882);
nand UO_221 (O_221,N_4119,N_4010);
or UO_222 (O_222,N_4688,N_4154);
or UO_223 (O_223,N_4230,N_4319);
and UO_224 (O_224,N_4162,N_4825);
nand UO_225 (O_225,N_4413,N_4684);
nor UO_226 (O_226,N_4336,N_4100);
nor UO_227 (O_227,N_4443,N_4235);
or UO_228 (O_228,N_4766,N_4671);
or UO_229 (O_229,N_4507,N_4447);
or UO_230 (O_230,N_4584,N_4189);
and UO_231 (O_231,N_4561,N_4365);
nor UO_232 (O_232,N_4223,N_4332);
or UO_233 (O_233,N_4251,N_4792);
and UO_234 (O_234,N_4832,N_4656);
xnor UO_235 (O_235,N_4172,N_4357);
or UO_236 (O_236,N_4122,N_4761);
nand UO_237 (O_237,N_4616,N_4622);
nor UO_238 (O_238,N_4873,N_4953);
or UO_239 (O_239,N_4515,N_4770);
and UO_240 (O_240,N_4099,N_4173);
and UO_241 (O_241,N_4242,N_4132);
xor UO_242 (O_242,N_4554,N_4799);
nand UO_243 (O_243,N_4883,N_4710);
or UO_244 (O_244,N_4813,N_4893);
nor UO_245 (O_245,N_4817,N_4677);
and UO_246 (O_246,N_4718,N_4260);
nor UO_247 (O_247,N_4341,N_4418);
nand UO_248 (O_248,N_4227,N_4528);
nor UO_249 (O_249,N_4708,N_4373);
or UO_250 (O_250,N_4405,N_4314);
and UO_251 (O_251,N_4066,N_4978);
and UO_252 (O_252,N_4955,N_4088);
and UO_253 (O_253,N_4118,N_4945);
and UO_254 (O_254,N_4942,N_4692);
nand UO_255 (O_255,N_4094,N_4550);
or UO_256 (O_256,N_4502,N_4905);
nand UO_257 (O_257,N_4481,N_4498);
xor UO_258 (O_258,N_4783,N_4439);
nand UO_259 (O_259,N_4803,N_4277);
xnor UO_260 (O_260,N_4962,N_4581);
xor UO_261 (O_261,N_4562,N_4215);
and UO_262 (O_262,N_4577,N_4323);
xnor UO_263 (O_263,N_4937,N_4210);
nand UO_264 (O_264,N_4889,N_4176);
nor UO_265 (O_265,N_4281,N_4145);
and UO_266 (O_266,N_4644,N_4096);
xnor UO_267 (O_267,N_4843,N_4660);
and UO_268 (O_268,N_4190,N_4847);
or UO_269 (O_269,N_4169,N_4441);
nand UO_270 (O_270,N_4110,N_4123);
and UO_271 (O_271,N_4471,N_4560);
nor UO_272 (O_272,N_4630,N_4726);
nand UO_273 (O_273,N_4880,N_4343);
nand UO_274 (O_274,N_4830,N_4027);
or UO_275 (O_275,N_4524,N_4916);
nand UO_276 (O_276,N_4212,N_4965);
nor UO_277 (O_277,N_4431,N_4438);
or UO_278 (O_278,N_4164,N_4460);
or UO_279 (O_279,N_4226,N_4627);
or UO_280 (O_280,N_4595,N_4923);
nor UO_281 (O_281,N_4301,N_4421);
nor UO_282 (O_282,N_4733,N_4811);
or UO_283 (O_283,N_4611,N_4558);
xor UO_284 (O_284,N_4028,N_4051);
xor UO_285 (O_285,N_4828,N_4178);
and UO_286 (O_286,N_4659,N_4720);
or UO_287 (O_287,N_4423,N_4045);
and UO_288 (O_288,N_4331,N_4572);
nor UO_289 (O_289,N_4855,N_4293);
nor UO_290 (O_290,N_4651,N_4411);
nor UO_291 (O_291,N_4599,N_4909);
nor UO_292 (O_292,N_4204,N_4108);
and UO_293 (O_293,N_4772,N_4370);
xnor UO_294 (O_294,N_4533,N_4415);
nand UO_295 (O_295,N_4280,N_4911);
or UO_296 (O_296,N_4317,N_4921);
or UO_297 (O_297,N_4580,N_4221);
nand UO_298 (O_298,N_4140,N_4068);
xor UO_299 (O_299,N_4653,N_4419);
nand UO_300 (O_300,N_4141,N_4698);
nor UO_301 (O_301,N_4151,N_4477);
or UO_302 (O_302,N_4408,N_4961);
and UO_303 (O_303,N_4975,N_4821);
and UO_304 (O_304,N_4643,N_4262);
and UO_305 (O_305,N_4070,N_4753);
and UO_306 (O_306,N_4969,N_4067);
nor UO_307 (O_307,N_4449,N_4768);
and UO_308 (O_308,N_4972,N_4933);
xor UO_309 (O_309,N_4008,N_4501);
nand UO_310 (O_310,N_4063,N_4876);
and UO_311 (O_311,N_4457,N_4349);
nor UO_312 (O_312,N_4445,N_4806);
or UO_313 (O_313,N_4482,N_4996);
nor UO_314 (O_314,N_4334,N_4654);
or UO_315 (O_315,N_4313,N_4628);
nand UO_316 (O_316,N_4994,N_4417);
or UO_317 (O_317,N_4535,N_4976);
and UO_318 (O_318,N_4854,N_4663);
and UO_319 (O_319,N_4872,N_4327);
xnor UO_320 (O_320,N_4499,N_4267);
nand UO_321 (O_321,N_4741,N_4030);
nand UO_322 (O_322,N_4902,N_4685);
and UO_323 (O_323,N_4025,N_4216);
nand UO_324 (O_324,N_4539,N_4236);
nor UO_325 (O_325,N_4547,N_4852);
nand UO_326 (O_326,N_4061,N_4982);
xnor UO_327 (O_327,N_4913,N_4949);
or UO_328 (O_328,N_4113,N_4553);
nor UO_329 (O_329,N_4943,N_4609);
nor UO_330 (O_330,N_4756,N_4282);
and UO_331 (O_331,N_4217,N_4517);
and UO_332 (O_332,N_4368,N_4274);
xnor UO_333 (O_333,N_4503,N_4342);
nand UO_334 (O_334,N_4636,N_4548);
xnor UO_335 (O_335,N_4484,N_4073);
xnor UO_336 (O_336,N_4958,N_4491);
and UO_337 (O_337,N_4153,N_4265);
or UO_338 (O_338,N_4983,N_4296);
nor UO_339 (O_339,N_4480,N_4299);
or UO_340 (O_340,N_4675,N_4691);
nand UO_341 (O_341,N_4461,N_4925);
and UO_342 (O_342,N_4808,N_4544);
nand UO_343 (O_343,N_4839,N_4006);
or UO_344 (O_344,N_4620,N_4310);
and UO_345 (O_345,N_4039,N_4686);
and UO_346 (O_346,N_4896,N_4033);
nand UO_347 (O_347,N_4168,N_4103);
xnor UO_348 (O_348,N_4143,N_4435);
or UO_349 (O_349,N_4437,N_4546);
or UO_350 (O_350,N_4205,N_4571);
xnor UO_351 (O_351,N_4736,N_4701);
xor UO_352 (O_352,N_4860,N_4237);
or UO_353 (O_353,N_4693,N_4683);
nor UO_354 (O_354,N_4885,N_4990);
nor UO_355 (O_355,N_4166,N_4812);
xor UO_356 (O_356,N_4287,N_4968);
or UO_357 (O_357,N_4420,N_4886);
or UO_358 (O_358,N_4041,N_4930);
nand UO_359 (O_359,N_4513,N_4136);
nor UO_360 (O_360,N_4664,N_4092);
and UO_361 (O_361,N_4444,N_4716);
and UO_362 (O_362,N_4850,N_4964);
and UO_363 (O_363,N_4815,N_4780);
and UO_364 (O_364,N_4402,N_4606);
and UO_365 (O_365,N_4271,N_4816);
xor UO_366 (O_366,N_4106,N_4723);
and UO_367 (O_367,N_4887,N_4798);
or UO_368 (O_368,N_4307,N_4333);
xnor UO_369 (O_369,N_4928,N_4126);
nand UO_370 (O_370,N_4161,N_4985);
nand UO_371 (O_371,N_4781,N_4906);
and UO_372 (O_372,N_4297,N_4844);
and UO_373 (O_373,N_4031,N_4222);
xor UO_374 (O_374,N_4638,N_4292);
nor UO_375 (O_375,N_4986,N_4984);
nand UO_376 (O_376,N_4521,N_4352);
or UO_377 (O_377,N_4144,N_4674);
nor UO_378 (O_378,N_4520,N_4639);
or UO_379 (O_379,N_4988,N_4037);
nand UO_380 (O_380,N_4077,N_4941);
or UO_381 (O_381,N_4593,N_4001);
nand UO_382 (O_382,N_4363,N_4220);
xnor UO_383 (O_383,N_4149,N_4598);
nand UO_384 (O_384,N_4246,N_4669);
or UO_385 (O_385,N_4667,N_4273);
and UO_386 (O_386,N_4705,N_4655);
xnor UO_387 (O_387,N_4371,N_4747);
nand UO_388 (O_388,N_4093,N_4040);
nor UO_389 (O_389,N_4462,N_4309);
nand UO_390 (O_390,N_4250,N_4476);
or UO_391 (O_391,N_4127,N_4496);
or UO_392 (O_392,N_4306,N_4382);
or UO_393 (O_393,N_4232,N_4493);
nor UO_394 (O_394,N_4374,N_4647);
xor UO_395 (O_395,N_4032,N_4948);
and UO_396 (O_396,N_4056,N_4793);
and UO_397 (O_397,N_4804,N_4884);
xor UO_398 (O_398,N_4849,N_4904);
nor UO_399 (O_399,N_4275,N_4600);
or UO_400 (O_400,N_4206,N_4658);
nand UO_401 (O_401,N_4269,N_4543);
xnor UO_402 (O_402,N_4586,N_4432);
xnor UO_403 (O_403,N_4800,N_4254);
and UO_404 (O_404,N_4101,N_4728);
or UO_405 (O_405,N_4997,N_4579);
or UO_406 (O_406,N_4453,N_4856);
xnor UO_407 (O_407,N_4637,N_4218);
nand UO_408 (O_408,N_4545,N_4731);
or UO_409 (O_409,N_4645,N_4409);
nand UO_410 (O_410,N_4391,N_4556);
or UO_411 (O_411,N_4359,N_4632);
nand UO_412 (O_412,N_4634,N_4750);
and UO_413 (O_413,N_4673,N_4072);
nand UO_414 (O_414,N_4322,N_4532);
nand UO_415 (O_415,N_4440,N_4642);
xor UO_416 (O_416,N_4744,N_4401);
and UO_417 (O_417,N_4703,N_4328);
xnor UO_418 (O_418,N_4633,N_4794);
xnor UO_419 (O_419,N_4917,N_4557);
nand UO_420 (O_420,N_4591,N_4428);
and UO_421 (O_421,N_4786,N_4494);
nand UO_422 (O_422,N_4807,N_4570);
nand UO_423 (O_423,N_4831,N_4366);
and UO_424 (O_424,N_4785,N_4512);
xor UO_425 (O_425,N_4107,N_4138);
nand UO_426 (O_426,N_4436,N_4776);
xor UO_427 (O_427,N_4171,N_4286);
nor UO_428 (O_428,N_4619,N_4302);
and UO_429 (O_429,N_4823,N_4788);
or UO_430 (O_430,N_4201,N_4715);
xnor UO_431 (O_431,N_4105,N_4959);
xor UO_432 (O_432,N_4300,N_4000);
nor UO_433 (O_433,N_4351,N_4455);
xor UO_434 (O_434,N_4765,N_4057);
nor UO_435 (O_435,N_4610,N_4678);
nor UO_436 (O_436,N_4007,N_4751);
and UO_437 (O_437,N_4240,N_4569);
nand UO_438 (O_438,N_4729,N_4536);
nand UO_439 (O_439,N_4552,N_4186);
or UO_440 (O_440,N_4754,N_4470);
and UO_441 (O_441,N_4187,N_4175);
and UO_442 (O_442,N_4200,N_4163);
or UO_443 (O_443,N_4016,N_4734);
and UO_444 (O_444,N_4757,N_4315);
nor UO_445 (O_445,N_4052,N_4347);
and UO_446 (O_446,N_4573,N_4992);
or UO_447 (O_447,N_4468,N_4195);
or UO_448 (O_448,N_4900,N_4626);
and UO_449 (O_449,N_4657,N_4388);
xnor UO_450 (O_450,N_4999,N_4487);
nand UO_451 (O_451,N_4345,N_4133);
xor UO_452 (O_452,N_4044,N_4234);
xnor UO_453 (O_453,N_4244,N_4004);
nor UO_454 (O_454,N_4867,N_4592);
and UO_455 (O_455,N_4214,N_4053);
xnor UO_456 (O_456,N_4386,N_4666);
or UO_457 (O_457,N_4704,N_4202);
or UO_458 (O_458,N_4640,N_4845);
and UO_459 (O_459,N_4596,N_4957);
or UO_460 (O_460,N_4541,N_4348);
xor UO_461 (O_461,N_4085,N_4434);
nand UO_462 (O_462,N_4137,N_4394);
nor UO_463 (O_463,N_4465,N_4735);
and UO_464 (O_464,N_4165,N_4224);
and UO_465 (O_465,N_4820,N_4350);
xor UO_466 (O_466,N_4608,N_4932);
nor UO_467 (O_467,N_4631,N_4709);
xnor UO_468 (O_468,N_4451,N_4115);
nor UO_469 (O_469,N_4869,N_4464);
xor UO_470 (O_470,N_4763,N_4895);
nor UO_471 (O_471,N_4706,N_4979);
nor UO_472 (O_472,N_4537,N_4383);
or UO_473 (O_473,N_4810,N_4998);
and UO_474 (O_474,N_4879,N_4003);
nor UO_475 (O_475,N_4565,N_4014);
nand UO_476 (O_476,N_4617,N_4035);
nand UO_477 (O_477,N_4285,N_4104);
xnor UO_478 (O_478,N_4575,N_4951);
nand UO_479 (O_479,N_4618,N_4822);
nor UO_480 (O_480,N_4903,N_4801);
xor UO_481 (O_481,N_4740,N_4466);
xnor UO_482 (O_482,N_4717,N_4567);
and UO_483 (O_483,N_4829,N_4614);
or UO_484 (O_484,N_4760,N_4779);
nand UO_485 (O_485,N_4641,N_4160);
nand UO_486 (O_486,N_4995,N_4699);
and UO_487 (O_487,N_4870,N_4426);
xnor UO_488 (O_488,N_4054,N_4603);
or UO_489 (O_489,N_4367,N_4233);
or UO_490 (O_490,N_4279,N_4745);
and UO_491 (O_491,N_4510,N_4689);
nor UO_492 (O_492,N_4188,N_4252);
nand UO_493 (O_493,N_4174,N_4316);
nand UO_494 (O_494,N_4624,N_4771);
and UO_495 (O_495,N_4700,N_4377);
nand UO_496 (O_496,N_4899,N_4459);
or UO_497 (O_497,N_4050,N_4702);
nand UO_498 (O_498,N_4395,N_4399);
or UO_499 (O_499,N_4015,N_4228);
nand UO_500 (O_500,N_4839,N_4937);
nand UO_501 (O_501,N_4574,N_4061);
nand UO_502 (O_502,N_4015,N_4458);
and UO_503 (O_503,N_4760,N_4682);
or UO_504 (O_504,N_4370,N_4460);
nor UO_505 (O_505,N_4552,N_4364);
nor UO_506 (O_506,N_4863,N_4214);
xor UO_507 (O_507,N_4048,N_4693);
or UO_508 (O_508,N_4474,N_4130);
nor UO_509 (O_509,N_4461,N_4147);
nand UO_510 (O_510,N_4741,N_4919);
nor UO_511 (O_511,N_4090,N_4204);
xnor UO_512 (O_512,N_4863,N_4424);
xnor UO_513 (O_513,N_4156,N_4023);
and UO_514 (O_514,N_4586,N_4457);
nand UO_515 (O_515,N_4217,N_4388);
or UO_516 (O_516,N_4819,N_4641);
and UO_517 (O_517,N_4543,N_4541);
nand UO_518 (O_518,N_4165,N_4914);
xnor UO_519 (O_519,N_4377,N_4728);
nand UO_520 (O_520,N_4692,N_4097);
and UO_521 (O_521,N_4094,N_4139);
or UO_522 (O_522,N_4902,N_4621);
nor UO_523 (O_523,N_4841,N_4170);
or UO_524 (O_524,N_4697,N_4822);
xor UO_525 (O_525,N_4287,N_4066);
nor UO_526 (O_526,N_4942,N_4707);
xnor UO_527 (O_527,N_4615,N_4047);
and UO_528 (O_528,N_4874,N_4698);
and UO_529 (O_529,N_4910,N_4112);
or UO_530 (O_530,N_4477,N_4643);
and UO_531 (O_531,N_4682,N_4319);
nand UO_532 (O_532,N_4990,N_4222);
xor UO_533 (O_533,N_4464,N_4391);
xnor UO_534 (O_534,N_4485,N_4994);
nand UO_535 (O_535,N_4208,N_4096);
or UO_536 (O_536,N_4450,N_4636);
xor UO_537 (O_537,N_4439,N_4451);
nor UO_538 (O_538,N_4897,N_4205);
or UO_539 (O_539,N_4836,N_4890);
xor UO_540 (O_540,N_4422,N_4943);
and UO_541 (O_541,N_4010,N_4240);
or UO_542 (O_542,N_4117,N_4807);
xor UO_543 (O_543,N_4795,N_4266);
nor UO_544 (O_544,N_4467,N_4106);
or UO_545 (O_545,N_4037,N_4064);
nand UO_546 (O_546,N_4491,N_4647);
and UO_547 (O_547,N_4339,N_4120);
nand UO_548 (O_548,N_4265,N_4832);
nor UO_549 (O_549,N_4264,N_4414);
nor UO_550 (O_550,N_4455,N_4144);
or UO_551 (O_551,N_4159,N_4552);
and UO_552 (O_552,N_4568,N_4325);
and UO_553 (O_553,N_4695,N_4265);
xor UO_554 (O_554,N_4831,N_4313);
xor UO_555 (O_555,N_4346,N_4195);
nor UO_556 (O_556,N_4979,N_4146);
or UO_557 (O_557,N_4837,N_4828);
or UO_558 (O_558,N_4299,N_4495);
nand UO_559 (O_559,N_4810,N_4136);
nor UO_560 (O_560,N_4249,N_4014);
and UO_561 (O_561,N_4797,N_4316);
and UO_562 (O_562,N_4450,N_4599);
nand UO_563 (O_563,N_4872,N_4685);
xnor UO_564 (O_564,N_4049,N_4050);
and UO_565 (O_565,N_4566,N_4921);
or UO_566 (O_566,N_4255,N_4975);
and UO_567 (O_567,N_4235,N_4264);
xor UO_568 (O_568,N_4751,N_4738);
nand UO_569 (O_569,N_4966,N_4350);
or UO_570 (O_570,N_4355,N_4292);
nor UO_571 (O_571,N_4695,N_4288);
xor UO_572 (O_572,N_4089,N_4815);
xor UO_573 (O_573,N_4175,N_4643);
xnor UO_574 (O_574,N_4806,N_4753);
nand UO_575 (O_575,N_4315,N_4038);
nor UO_576 (O_576,N_4763,N_4695);
nor UO_577 (O_577,N_4194,N_4013);
nand UO_578 (O_578,N_4527,N_4385);
nor UO_579 (O_579,N_4259,N_4318);
nand UO_580 (O_580,N_4812,N_4875);
nor UO_581 (O_581,N_4679,N_4755);
nor UO_582 (O_582,N_4120,N_4725);
xnor UO_583 (O_583,N_4228,N_4466);
nand UO_584 (O_584,N_4680,N_4811);
or UO_585 (O_585,N_4974,N_4793);
nand UO_586 (O_586,N_4271,N_4009);
and UO_587 (O_587,N_4689,N_4550);
nor UO_588 (O_588,N_4466,N_4542);
or UO_589 (O_589,N_4836,N_4102);
and UO_590 (O_590,N_4393,N_4394);
nor UO_591 (O_591,N_4003,N_4390);
xnor UO_592 (O_592,N_4253,N_4408);
nor UO_593 (O_593,N_4270,N_4411);
xnor UO_594 (O_594,N_4484,N_4884);
nor UO_595 (O_595,N_4296,N_4047);
nor UO_596 (O_596,N_4555,N_4742);
or UO_597 (O_597,N_4916,N_4274);
nand UO_598 (O_598,N_4657,N_4727);
xor UO_599 (O_599,N_4304,N_4146);
nand UO_600 (O_600,N_4211,N_4455);
and UO_601 (O_601,N_4319,N_4168);
nor UO_602 (O_602,N_4385,N_4422);
xnor UO_603 (O_603,N_4891,N_4987);
or UO_604 (O_604,N_4736,N_4226);
xnor UO_605 (O_605,N_4540,N_4897);
xor UO_606 (O_606,N_4991,N_4453);
xnor UO_607 (O_607,N_4870,N_4146);
nand UO_608 (O_608,N_4631,N_4511);
nor UO_609 (O_609,N_4820,N_4270);
nand UO_610 (O_610,N_4523,N_4972);
and UO_611 (O_611,N_4858,N_4685);
xor UO_612 (O_612,N_4483,N_4853);
nand UO_613 (O_613,N_4469,N_4903);
nand UO_614 (O_614,N_4088,N_4617);
nor UO_615 (O_615,N_4794,N_4758);
xnor UO_616 (O_616,N_4633,N_4718);
or UO_617 (O_617,N_4744,N_4317);
or UO_618 (O_618,N_4233,N_4190);
nand UO_619 (O_619,N_4203,N_4293);
xor UO_620 (O_620,N_4902,N_4865);
and UO_621 (O_621,N_4853,N_4600);
xor UO_622 (O_622,N_4937,N_4555);
and UO_623 (O_623,N_4695,N_4594);
nor UO_624 (O_624,N_4167,N_4618);
nand UO_625 (O_625,N_4155,N_4739);
and UO_626 (O_626,N_4042,N_4978);
nand UO_627 (O_627,N_4591,N_4411);
and UO_628 (O_628,N_4035,N_4535);
and UO_629 (O_629,N_4309,N_4094);
and UO_630 (O_630,N_4694,N_4637);
and UO_631 (O_631,N_4258,N_4311);
nor UO_632 (O_632,N_4117,N_4057);
xor UO_633 (O_633,N_4869,N_4315);
nor UO_634 (O_634,N_4274,N_4171);
and UO_635 (O_635,N_4339,N_4929);
xnor UO_636 (O_636,N_4889,N_4646);
or UO_637 (O_637,N_4173,N_4683);
nor UO_638 (O_638,N_4029,N_4077);
and UO_639 (O_639,N_4332,N_4772);
nor UO_640 (O_640,N_4885,N_4884);
or UO_641 (O_641,N_4920,N_4258);
xor UO_642 (O_642,N_4609,N_4448);
or UO_643 (O_643,N_4282,N_4019);
and UO_644 (O_644,N_4965,N_4411);
and UO_645 (O_645,N_4025,N_4620);
xor UO_646 (O_646,N_4046,N_4468);
nand UO_647 (O_647,N_4896,N_4805);
nand UO_648 (O_648,N_4324,N_4337);
nand UO_649 (O_649,N_4886,N_4288);
or UO_650 (O_650,N_4764,N_4646);
and UO_651 (O_651,N_4594,N_4730);
and UO_652 (O_652,N_4823,N_4352);
xnor UO_653 (O_653,N_4973,N_4692);
xor UO_654 (O_654,N_4356,N_4270);
and UO_655 (O_655,N_4525,N_4856);
nor UO_656 (O_656,N_4365,N_4230);
or UO_657 (O_657,N_4426,N_4013);
nand UO_658 (O_658,N_4203,N_4630);
nor UO_659 (O_659,N_4215,N_4685);
xnor UO_660 (O_660,N_4783,N_4080);
or UO_661 (O_661,N_4001,N_4660);
nor UO_662 (O_662,N_4888,N_4900);
or UO_663 (O_663,N_4066,N_4210);
and UO_664 (O_664,N_4169,N_4924);
nor UO_665 (O_665,N_4325,N_4916);
or UO_666 (O_666,N_4266,N_4543);
nand UO_667 (O_667,N_4976,N_4451);
and UO_668 (O_668,N_4925,N_4144);
nand UO_669 (O_669,N_4286,N_4437);
and UO_670 (O_670,N_4062,N_4227);
and UO_671 (O_671,N_4219,N_4252);
nor UO_672 (O_672,N_4440,N_4053);
nand UO_673 (O_673,N_4222,N_4464);
nand UO_674 (O_674,N_4527,N_4052);
xnor UO_675 (O_675,N_4893,N_4514);
xor UO_676 (O_676,N_4815,N_4247);
nor UO_677 (O_677,N_4166,N_4536);
and UO_678 (O_678,N_4610,N_4454);
xor UO_679 (O_679,N_4648,N_4853);
and UO_680 (O_680,N_4612,N_4658);
or UO_681 (O_681,N_4505,N_4664);
and UO_682 (O_682,N_4828,N_4985);
nand UO_683 (O_683,N_4968,N_4244);
xor UO_684 (O_684,N_4439,N_4797);
nor UO_685 (O_685,N_4609,N_4488);
nand UO_686 (O_686,N_4861,N_4041);
nand UO_687 (O_687,N_4420,N_4487);
nor UO_688 (O_688,N_4722,N_4159);
nor UO_689 (O_689,N_4621,N_4517);
nand UO_690 (O_690,N_4521,N_4653);
nand UO_691 (O_691,N_4800,N_4154);
and UO_692 (O_692,N_4581,N_4813);
xor UO_693 (O_693,N_4405,N_4260);
nand UO_694 (O_694,N_4925,N_4850);
xor UO_695 (O_695,N_4609,N_4007);
nand UO_696 (O_696,N_4428,N_4665);
nor UO_697 (O_697,N_4289,N_4175);
or UO_698 (O_698,N_4878,N_4544);
or UO_699 (O_699,N_4088,N_4157);
or UO_700 (O_700,N_4344,N_4022);
and UO_701 (O_701,N_4145,N_4595);
or UO_702 (O_702,N_4664,N_4943);
and UO_703 (O_703,N_4499,N_4582);
or UO_704 (O_704,N_4441,N_4584);
nor UO_705 (O_705,N_4309,N_4410);
xor UO_706 (O_706,N_4534,N_4059);
nor UO_707 (O_707,N_4817,N_4479);
xor UO_708 (O_708,N_4820,N_4661);
nor UO_709 (O_709,N_4749,N_4794);
nand UO_710 (O_710,N_4421,N_4626);
nor UO_711 (O_711,N_4385,N_4734);
xor UO_712 (O_712,N_4228,N_4742);
and UO_713 (O_713,N_4357,N_4805);
nor UO_714 (O_714,N_4068,N_4411);
nor UO_715 (O_715,N_4670,N_4875);
nor UO_716 (O_716,N_4589,N_4318);
and UO_717 (O_717,N_4334,N_4637);
or UO_718 (O_718,N_4763,N_4437);
nor UO_719 (O_719,N_4825,N_4747);
xor UO_720 (O_720,N_4838,N_4873);
xnor UO_721 (O_721,N_4445,N_4694);
nor UO_722 (O_722,N_4575,N_4314);
nor UO_723 (O_723,N_4660,N_4556);
or UO_724 (O_724,N_4305,N_4820);
and UO_725 (O_725,N_4920,N_4701);
xor UO_726 (O_726,N_4170,N_4194);
or UO_727 (O_727,N_4189,N_4435);
xor UO_728 (O_728,N_4956,N_4311);
or UO_729 (O_729,N_4620,N_4315);
or UO_730 (O_730,N_4354,N_4242);
nand UO_731 (O_731,N_4025,N_4872);
xnor UO_732 (O_732,N_4984,N_4566);
nand UO_733 (O_733,N_4007,N_4075);
nand UO_734 (O_734,N_4741,N_4519);
nor UO_735 (O_735,N_4918,N_4617);
nand UO_736 (O_736,N_4292,N_4018);
nand UO_737 (O_737,N_4777,N_4214);
xor UO_738 (O_738,N_4122,N_4063);
or UO_739 (O_739,N_4957,N_4435);
nand UO_740 (O_740,N_4896,N_4938);
nand UO_741 (O_741,N_4701,N_4988);
nand UO_742 (O_742,N_4346,N_4481);
and UO_743 (O_743,N_4670,N_4202);
or UO_744 (O_744,N_4802,N_4324);
xnor UO_745 (O_745,N_4905,N_4130);
or UO_746 (O_746,N_4477,N_4923);
and UO_747 (O_747,N_4407,N_4191);
nand UO_748 (O_748,N_4702,N_4081);
or UO_749 (O_749,N_4403,N_4694);
nand UO_750 (O_750,N_4890,N_4007);
and UO_751 (O_751,N_4538,N_4526);
nor UO_752 (O_752,N_4860,N_4107);
and UO_753 (O_753,N_4439,N_4747);
or UO_754 (O_754,N_4858,N_4010);
nand UO_755 (O_755,N_4095,N_4586);
xnor UO_756 (O_756,N_4212,N_4439);
nand UO_757 (O_757,N_4916,N_4509);
or UO_758 (O_758,N_4569,N_4992);
xor UO_759 (O_759,N_4798,N_4727);
xnor UO_760 (O_760,N_4258,N_4753);
xor UO_761 (O_761,N_4688,N_4225);
nand UO_762 (O_762,N_4884,N_4685);
and UO_763 (O_763,N_4949,N_4766);
and UO_764 (O_764,N_4811,N_4220);
xor UO_765 (O_765,N_4382,N_4622);
xnor UO_766 (O_766,N_4336,N_4728);
nor UO_767 (O_767,N_4568,N_4413);
nand UO_768 (O_768,N_4511,N_4365);
or UO_769 (O_769,N_4994,N_4189);
nor UO_770 (O_770,N_4393,N_4988);
and UO_771 (O_771,N_4178,N_4459);
or UO_772 (O_772,N_4175,N_4591);
and UO_773 (O_773,N_4778,N_4221);
xnor UO_774 (O_774,N_4882,N_4412);
xor UO_775 (O_775,N_4175,N_4297);
xnor UO_776 (O_776,N_4360,N_4009);
nand UO_777 (O_777,N_4405,N_4095);
nand UO_778 (O_778,N_4755,N_4144);
or UO_779 (O_779,N_4773,N_4809);
nor UO_780 (O_780,N_4744,N_4594);
xnor UO_781 (O_781,N_4101,N_4396);
nand UO_782 (O_782,N_4543,N_4521);
nor UO_783 (O_783,N_4935,N_4569);
or UO_784 (O_784,N_4340,N_4175);
or UO_785 (O_785,N_4210,N_4223);
or UO_786 (O_786,N_4905,N_4271);
or UO_787 (O_787,N_4354,N_4784);
nor UO_788 (O_788,N_4166,N_4159);
or UO_789 (O_789,N_4096,N_4962);
or UO_790 (O_790,N_4806,N_4772);
or UO_791 (O_791,N_4787,N_4020);
or UO_792 (O_792,N_4983,N_4793);
or UO_793 (O_793,N_4437,N_4670);
or UO_794 (O_794,N_4467,N_4331);
or UO_795 (O_795,N_4218,N_4877);
xor UO_796 (O_796,N_4067,N_4149);
xor UO_797 (O_797,N_4612,N_4968);
and UO_798 (O_798,N_4661,N_4011);
nor UO_799 (O_799,N_4826,N_4183);
nor UO_800 (O_800,N_4570,N_4806);
or UO_801 (O_801,N_4319,N_4156);
nand UO_802 (O_802,N_4045,N_4317);
xnor UO_803 (O_803,N_4113,N_4444);
or UO_804 (O_804,N_4291,N_4791);
and UO_805 (O_805,N_4621,N_4016);
and UO_806 (O_806,N_4011,N_4571);
nand UO_807 (O_807,N_4743,N_4133);
nand UO_808 (O_808,N_4916,N_4849);
nand UO_809 (O_809,N_4243,N_4674);
nand UO_810 (O_810,N_4840,N_4001);
nand UO_811 (O_811,N_4628,N_4009);
nand UO_812 (O_812,N_4959,N_4468);
xor UO_813 (O_813,N_4996,N_4940);
nand UO_814 (O_814,N_4377,N_4513);
and UO_815 (O_815,N_4502,N_4599);
and UO_816 (O_816,N_4559,N_4576);
or UO_817 (O_817,N_4805,N_4122);
nand UO_818 (O_818,N_4001,N_4889);
or UO_819 (O_819,N_4529,N_4409);
and UO_820 (O_820,N_4493,N_4956);
and UO_821 (O_821,N_4687,N_4338);
xor UO_822 (O_822,N_4796,N_4503);
and UO_823 (O_823,N_4331,N_4426);
nor UO_824 (O_824,N_4346,N_4855);
nand UO_825 (O_825,N_4117,N_4088);
and UO_826 (O_826,N_4262,N_4620);
or UO_827 (O_827,N_4942,N_4631);
and UO_828 (O_828,N_4952,N_4672);
nor UO_829 (O_829,N_4120,N_4062);
or UO_830 (O_830,N_4183,N_4294);
and UO_831 (O_831,N_4941,N_4175);
nor UO_832 (O_832,N_4328,N_4723);
nor UO_833 (O_833,N_4229,N_4254);
and UO_834 (O_834,N_4952,N_4008);
or UO_835 (O_835,N_4333,N_4259);
or UO_836 (O_836,N_4174,N_4278);
nor UO_837 (O_837,N_4896,N_4510);
xor UO_838 (O_838,N_4894,N_4595);
nor UO_839 (O_839,N_4381,N_4723);
or UO_840 (O_840,N_4068,N_4291);
or UO_841 (O_841,N_4645,N_4630);
nand UO_842 (O_842,N_4312,N_4404);
or UO_843 (O_843,N_4972,N_4715);
nand UO_844 (O_844,N_4161,N_4077);
nand UO_845 (O_845,N_4479,N_4597);
nand UO_846 (O_846,N_4192,N_4992);
nor UO_847 (O_847,N_4719,N_4959);
and UO_848 (O_848,N_4588,N_4203);
and UO_849 (O_849,N_4552,N_4573);
nand UO_850 (O_850,N_4994,N_4010);
and UO_851 (O_851,N_4385,N_4691);
and UO_852 (O_852,N_4123,N_4043);
and UO_853 (O_853,N_4812,N_4117);
or UO_854 (O_854,N_4182,N_4106);
or UO_855 (O_855,N_4672,N_4961);
nor UO_856 (O_856,N_4047,N_4956);
and UO_857 (O_857,N_4445,N_4134);
nor UO_858 (O_858,N_4363,N_4794);
nor UO_859 (O_859,N_4969,N_4692);
xnor UO_860 (O_860,N_4842,N_4278);
xnor UO_861 (O_861,N_4554,N_4035);
xnor UO_862 (O_862,N_4848,N_4086);
nand UO_863 (O_863,N_4559,N_4712);
and UO_864 (O_864,N_4399,N_4362);
nor UO_865 (O_865,N_4943,N_4619);
or UO_866 (O_866,N_4248,N_4130);
nand UO_867 (O_867,N_4252,N_4955);
or UO_868 (O_868,N_4145,N_4671);
xor UO_869 (O_869,N_4269,N_4895);
or UO_870 (O_870,N_4767,N_4991);
nor UO_871 (O_871,N_4722,N_4221);
nor UO_872 (O_872,N_4504,N_4621);
or UO_873 (O_873,N_4632,N_4314);
or UO_874 (O_874,N_4037,N_4659);
or UO_875 (O_875,N_4968,N_4870);
nor UO_876 (O_876,N_4011,N_4480);
xor UO_877 (O_877,N_4387,N_4340);
or UO_878 (O_878,N_4109,N_4358);
nor UO_879 (O_879,N_4518,N_4999);
or UO_880 (O_880,N_4352,N_4810);
nand UO_881 (O_881,N_4210,N_4362);
and UO_882 (O_882,N_4198,N_4589);
nand UO_883 (O_883,N_4250,N_4433);
nand UO_884 (O_884,N_4346,N_4242);
nand UO_885 (O_885,N_4994,N_4208);
nor UO_886 (O_886,N_4036,N_4584);
and UO_887 (O_887,N_4903,N_4132);
xor UO_888 (O_888,N_4151,N_4285);
nand UO_889 (O_889,N_4886,N_4297);
nand UO_890 (O_890,N_4501,N_4292);
or UO_891 (O_891,N_4639,N_4055);
xor UO_892 (O_892,N_4853,N_4363);
xnor UO_893 (O_893,N_4790,N_4875);
and UO_894 (O_894,N_4151,N_4798);
nand UO_895 (O_895,N_4312,N_4810);
xnor UO_896 (O_896,N_4370,N_4784);
and UO_897 (O_897,N_4225,N_4311);
nor UO_898 (O_898,N_4240,N_4093);
or UO_899 (O_899,N_4324,N_4012);
or UO_900 (O_900,N_4956,N_4737);
xnor UO_901 (O_901,N_4314,N_4615);
nand UO_902 (O_902,N_4122,N_4574);
xnor UO_903 (O_903,N_4910,N_4452);
and UO_904 (O_904,N_4776,N_4891);
and UO_905 (O_905,N_4439,N_4088);
nor UO_906 (O_906,N_4952,N_4053);
xnor UO_907 (O_907,N_4474,N_4122);
nand UO_908 (O_908,N_4921,N_4026);
nand UO_909 (O_909,N_4372,N_4724);
nor UO_910 (O_910,N_4343,N_4440);
nand UO_911 (O_911,N_4140,N_4839);
or UO_912 (O_912,N_4840,N_4218);
nand UO_913 (O_913,N_4031,N_4497);
nor UO_914 (O_914,N_4458,N_4926);
nand UO_915 (O_915,N_4755,N_4689);
nand UO_916 (O_916,N_4595,N_4723);
nand UO_917 (O_917,N_4231,N_4503);
nor UO_918 (O_918,N_4345,N_4454);
and UO_919 (O_919,N_4124,N_4485);
nor UO_920 (O_920,N_4354,N_4992);
nand UO_921 (O_921,N_4191,N_4244);
nor UO_922 (O_922,N_4864,N_4911);
and UO_923 (O_923,N_4568,N_4138);
and UO_924 (O_924,N_4465,N_4968);
nand UO_925 (O_925,N_4055,N_4923);
or UO_926 (O_926,N_4062,N_4189);
nand UO_927 (O_927,N_4162,N_4771);
xor UO_928 (O_928,N_4845,N_4739);
nand UO_929 (O_929,N_4619,N_4525);
or UO_930 (O_930,N_4425,N_4116);
and UO_931 (O_931,N_4381,N_4207);
or UO_932 (O_932,N_4395,N_4988);
xor UO_933 (O_933,N_4718,N_4459);
xnor UO_934 (O_934,N_4518,N_4793);
xnor UO_935 (O_935,N_4077,N_4584);
and UO_936 (O_936,N_4926,N_4394);
nand UO_937 (O_937,N_4951,N_4449);
and UO_938 (O_938,N_4864,N_4647);
xor UO_939 (O_939,N_4962,N_4347);
xor UO_940 (O_940,N_4889,N_4143);
xnor UO_941 (O_941,N_4804,N_4028);
or UO_942 (O_942,N_4402,N_4330);
nor UO_943 (O_943,N_4608,N_4903);
nand UO_944 (O_944,N_4802,N_4511);
nand UO_945 (O_945,N_4248,N_4400);
nor UO_946 (O_946,N_4390,N_4543);
nor UO_947 (O_947,N_4072,N_4024);
nor UO_948 (O_948,N_4546,N_4927);
and UO_949 (O_949,N_4460,N_4169);
nor UO_950 (O_950,N_4827,N_4060);
nor UO_951 (O_951,N_4749,N_4461);
nor UO_952 (O_952,N_4589,N_4309);
or UO_953 (O_953,N_4007,N_4006);
nand UO_954 (O_954,N_4022,N_4252);
nor UO_955 (O_955,N_4381,N_4354);
and UO_956 (O_956,N_4182,N_4651);
nand UO_957 (O_957,N_4140,N_4353);
nor UO_958 (O_958,N_4905,N_4114);
xnor UO_959 (O_959,N_4664,N_4054);
xor UO_960 (O_960,N_4421,N_4228);
and UO_961 (O_961,N_4813,N_4132);
and UO_962 (O_962,N_4202,N_4756);
nand UO_963 (O_963,N_4080,N_4318);
xnor UO_964 (O_964,N_4812,N_4931);
xnor UO_965 (O_965,N_4345,N_4906);
xnor UO_966 (O_966,N_4110,N_4031);
nor UO_967 (O_967,N_4266,N_4322);
nor UO_968 (O_968,N_4098,N_4685);
and UO_969 (O_969,N_4907,N_4439);
or UO_970 (O_970,N_4680,N_4922);
xnor UO_971 (O_971,N_4384,N_4020);
nor UO_972 (O_972,N_4388,N_4316);
xor UO_973 (O_973,N_4934,N_4077);
and UO_974 (O_974,N_4291,N_4576);
and UO_975 (O_975,N_4788,N_4917);
nand UO_976 (O_976,N_4718,N_4047);
or UO_977 (O_977,N_4798,N_4455);
nand UO_978 (O_978,N_4169,N_4031);
nor UO_979 (O_979,N_4096,N_4031);
nand UO_980 (O_980,N_4585,N_4627);
or UO_981 (O_981,N_4001,N_4842);
nor UO_982 (O_982,N_4365,N_4044);
or UO_983 (O_983,N_4535,N_4944);
or UO_984 (O_984,N_4960,N_4747);
nor UO_985 (O_985,N_4275,N_4475);
nor UO_986 (O_986,N_4675,N_4972);
nor UO_987 (O_987,N_4905,N_4430);
nand UO_988 (O_988,N_4230,N_4172);
and UO_989 (O_989,N_4799,N_4540);
nor UO_990 (O_990,N_4874,N_4048);
or UO_991 (O_991,N_4960,N_4284);
nor UO_992 (O_992,N_4924,N_4418);
nand UO_993 (O_993,N_4716,N_4895);
xnor UO_994 (O_994,N_4213,N_4254);
xnor UO_995 (O_995,N_4940,N_4991);
xnor UO_996 (O_996,N_4516,N_4111);
nand UO_997 (O_997,N_4006,N_4491);
nand UO_998 (O_998,N_4344,N_4169);
nor UO_999 (O_999,N_4429,N_4421);
endmodule