module basic_750_5000_1000_50_levels_5xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
nand U0 (N_0,In_109,In_377);
nand U1 (N_1,In_134,In_528);
xor U2 (N_2,In_499,In_725);
nand U3 (N_3,In_687,In_391);
and U4 (N_4,In_630,In_339);
nor U5 (N_5,In_380,In_596);
xnor U6 (N_6,In_437,In_254);
nand U7 (N_7,In_588,In_705);
nor U8 (N_8,In_697,In_464);
nand U9 (N_9,In_652,In_500);
nor U10 (N_10,In_592,In_653);
nor U11 (N_11,In_442,In_407);
nor U12 (N_12,In_600,In_123);
and U13 (N_13,In_477,In_89);
nand U14 (N_14,In_34,In_505);
and U15 (N_15,In_272,In_122);
xnor U16 (N_16,In_397,In_96);
and U17 (N_17,In_712,In_703);
nand U18 (N_18,In_269,In_153);
nor U19 (N_19,In_516,In_206);
nand U20 (N_20,In_243,In_502);
nor U21 (N_21,In_620,In_44);
nand U22 (N_22,In_237,In_195);
nand U23 (N_23,In_574,In_527);
or U24 (N_24,In_404,In_340);
or U25 (N_25,In_250,In_587);
nand U26 (N_26,In_7,In_576);
xnor U27 (N_27,In_646,In_410);
xor U28 (N_28,In_10,In_655);
xnor U29 (N_29,In_119,In_113);
xor U30 (N_30,In_227,In_615);
nand U31 (N_31,In_275,In_204);
nand U32 (N_32,In_638,In_190);
or U33 (N_33,In_737,In_333);
or U34 (N_34,In_2,In_367);
or U35 (N_35,In_445,In_682);
nor U36 (N_36,In_656,In_173);
or U37 (N_37,In_523,In_738);
and U38 (N_38,In_559,In_337);
nand U39 (N_39,In_110,In_688);
nand U40 (N_40,In_28,In_520);
and U41 (N_41,In_14,In_362);
nor U42 (N_42,In_98,In_709);
or U43 (N_43,In_542,In_411);
and U44 (N_44,In_130,In_599);
and U45 (N_45,In_632,In_621);
and U46 (N_46,In_364,In_617);
or U47 (N_47,In_475,In_316);
nand U48 (N_48,In_570,In_235);
or U49 (N_49,In_580,In_627);
nand U50 (N_50,In_461,In_234);
nor U51 (N_51,In_504,In_37);
nand U52 (N_52,In_481,In_13);
and U53 (N_53,In_558,In_251);
nor U54 (N_54,In_555,In_536);
or U55 (N_55,In_701,In_112);
nor U56 (N_56,In_565,In_101);
nand U57 (N_57,In_661,In_641);
or U58 (N_58,In_405,In_288);
and U59 (N_59,In_749,In_708);
nor U60 (N_60,In_539,In_663);
nand U61 (N_61,In_566,In_293);
and U62 (N_62,In_350,In_32);
and U63 (N_63,In_295,In_205);
and U64 (N_64,In_665,In_106);
or U65 (N_65,In_616,In_549);
or U66 (N_66,In_42,In_317);
nor U67 (N_67,In_121,In_718);
or U68 (N_68,In_595,In_302);
nor U69 (N_69,In_38,In_69);
or U70 (N_70,In_714,In_309);
and U71 (N_71,In_660,In_470);
or U72 (N_72,In_294,In_374);
or U73 (N_73,In_526,In_468);
or U74 (N_74,In_540,In_624);
xor U75 (N_75,In_79,In_139);
nor U76 (N_76,In_508,In_512);
xor U77 (N_77,In_572,In_614);
and U78 (N_78,In_132,In_56);
nor U79 (N_79,In_399,In_51);
xnor U80 (N_80,In_165,In_544);
or U81 (N_81,In_233,In_246);
and U82 (N_82,In_240,In_267);
nor U83 (N_83,In_290,In_433);
and U84 (N_84,In_222,In_23);
nand U85 (N_85,In_747,In_730);
and U86 (N_86,In_264,In_715);
or U87 (N_87,In_328,In_462);
nor U88 (N_88,In_637,In_142);
nand U89 (N_89,In_353,In_678);
or U90 (N_90,In_488,In_211);
or U91 (N_91,In_623,In_131);
and U92 (N_92,In_16,In_382);
xor U93 (N_93,In_514,In_739);
nor U94 (N_94,In_63,In_591);
nor U95 (N_95,In_440,In_58);
and U96 (N_96,In_219,In_619);
or U97 (N_97,In_363,In_390);
xnor U98 (N_98,In_720,In_188);
and U99 (N_99,In_732,In_152);
nand U100 (N_100,In_327,In_117);
or U101 (N_101,In_118,N_45);
and U102 (N_102,In_585,N_94);
or U103 (N_103,In_681,In_444);
or U104 (N_104,In_114,In_429);
and U105 (N_105,N_92,In_179);
or U106 (N_106,N_9,In_210);
and U107 (N_107,In_17,In_169);
nand U108 (N_108,In_304,N_46);
or U109 (N_109,In_493,In_693);
nor U110 (N_110,In_248,In_313);
xnor U111 (N_111,In_149,In_184);
or U112 (N_112,In_628,In_704);
nor U113 (N_113,In_307,In_263);
nor U114 (N_114,In_668,In_322);
nand U115 (N_115,N_53,In_719);
or U116 (N_116,In_355,In_177);
and U117 (N_117,In_11,In_1);
nand U118 (N_118,In_498,In_633);
and U119 (N_119,In_352,In_335);
nand U120 (N_120,In_722,In_430);
nor U121 (N_121,In_291,In_529);
or U122 (N_122,N_81,In_373);
xnor U123 (N_123,In_40,In_519);
or U124 (N_124,In_608,In_650);
nor U125 (N_125,In_170,In_606);
nand U126 (N_126,In_76,In_143);
or U127 (N_127,In_438,In_490);
and U128 (N_128,In_278,In_224);
nand U129 (N_129,N_90,In_479);
and U130 (N_130,In_103,N_22);
and U131 (N_131,In_135,In_568);
or U132 (N_132,N_48,N_2);
xnor U133 (N_133,In_65,In_324);
and U134 (N_134,In_408,In_181);
and U135 (N_135,In_187,In_601);
nor U136 (N_136,In_217,In_318);
nand U137 (N_137,In_748,In_5);
and U138 (N_138,In_631,In_483);
nor U139 (N_139,In_239,In_501);
xnor U140 (N_140,N_30,In_120);
nor U141 (N_141,In_597,In_236);
nand U142 (N_142,In_182,In_77);
nor U143 (N_143,In_582,In_292);
or U144 (N_144,N_44,N_17);
and U145 (N_145,In_244,In_742);
nor U146 (N_146,In_30,In_50);
or U147 (N_147,N_31,In_667);
xor U148 (N_148,In_225,In_90);
and U149 (N_149,In_396,In_629);
and U150 (N_150,N_24,In_107);
or U151 (N_151,In_141,In_562);
or U152 (N_152,In_154,In_604);
nor U153 (N_153,In_435,In_389);
nor U154 (N_154,In_651,In_716);
xnor U155 (N_155,In_265,In_700);
or U156 (N_156,In_645,In_453);
nor U157 (N_157,In_329,In_456);
nand U158 (N_158,In_70,In_221);
nor U159 (N_159,In_392,In_127);
and U160 (N_160,In_670,In_586);
and U161 (N_161,N_41,In_743);
or U162 (N_162,In_622,In_679);
nor U163 (N_163,In_745,In_330);
xnor U164 (N_164,In_603,In_241);
or U165 (N_165,In_354,In_35);
and U166 (N_166,In_43,In_68);
or U167 (N_167,N_49,In_415);
or U168 (N_168,In_276,In_201);
nand U169 (N_169,In_18,N_36);
nand U170 (N_170,N_27,In_87);
and U171 (N_171,In_451,In_115);
nand U172 (N_172,In_398,In_185);
nand U173 (N_173,In_268,In_496);
xnor U174 (N_174,In_360,In_326);
nand U175 (N_175,In_286,In_345);
nand U176 (N_176,N_26,In_534);
nor U177 (N_177,In_465,In_375);
nand U178 (N_178,N_85,In_431);
nand U179 (N_179,N_18,In_197);
nand U180 (N_180,In_625,In_53);
or U181 (N_181,N_80,In_62);
or U182 (N_182,In_680,N_93);
xor U183 (N_183,In_140,In_494);
xnor U184 (N_184,In_721,In_247);
nor U185 (N_185,In_563,In_575);
nand U186 (N_186,In_192,In_281);
xor U187 (N_187,In_521,In_129);
nor U188 (N_188,In_454,In_282);
and U189 (N_189,In_24,In_649);
nor U190 (N_190,In_138,In_448);
nand U191 (N_191,In_232,In_66);
nor U192 (N_192,In_33,In_172);
nand U193 (N_193,In_683,In_436);
and U194 (N_194,In_507,In_164);
nand U195 (N_195,In_561,In_194);
nor U196 (N_196,N_8,In_497);
and U197 (N_197,In_666,N_95);
nor U198 (N_198,In_299,In_711);
and U199 (N_199,In_532,In_581);
nand U200 (N_200,N_120,In_171);
nand U201 (N_201,In_452,In_57);
xnor U202 (N_202,In_341,In_515);
nand U203 (N_203,In_160,N_114);
nand U204 (N_204,In_612,In_102);
nand U205 (N_205,N_178,In_82);
nor U206 (N_206,In_212,N_57);
nor U207 (N_207,In_86,In_664);
nor U208 (N_208,In_551,N_82);
nand U209 (N_209,In_696,N_160);
or U210 (N_210,N_21,In_108);
and U211 (N_211,In_301,In_15);
xor U212 (N_212,N_38,In_594);
nand U213 (N_213,In_554,In_19);
and U214 (N_214,In_417,N_163);
or U215 (N_215,In_157,In_458);
and U216 (N_216,In_538,In_6);
nand U217 (N_217,In_424,N_16);
and U218 (N_218,N_137,In_460);
and U219 (N_219,In_491,In_459);
nand U220 (N_220,In_256,In_611);
and U221 (N_221,In_208,N_153);
or U222 (N_222,In_480,In_657);
or U223 (N_223,In_635,In_48);
nor U224 (N_224,N_116,In_351);
or U225 (N_225,In_297,N_154);
and U226 (N_226,In_686,In_510);
nand U227 (N_227,N_145,N_139);
or U228 (N_228,In_713,In_416);
and U229 (N_229,In_55,In_150);
or U230 (N_230,In_73,In_163);
nor U231 (N_231,In_613,In_673);
or U232 (N_232,N_127,In_511);
nor U233 (N_233,In_216,N_76);
xnor U234 (N_234,In_746,N_193);
nor U235 (N_235,In_209,In_81);
or U236 (N_236,In_403,In_677);
nor U237 (N_237,In_226,In_280);
xnor U238 (N_238,In_409,N_158);
xnor U239 (N_239,In_27,In_506);
xnor U240 (N_240,In_387,N_58);
and U241 (N_241,In_258,In_671);
nor U242 (N_242,In_552,In_257);
nor U243 (N_243,In_503,In_723);
nand U244 (N_244,In_394,N_88);
and U245 (N_245,In_530,N_188);
and U246 (N_246,In_545,N_155);
and U247 (N_247,In_8,In_71);
or U248 (N_248,In_471,N_75);
xnor U249 (N_249,In_648,In_384);
or U250 (N_250,In_395,N_89);
xor U251 (N_251,In_36,In_144);
nand U252 (N_252,In_126,In_361);
or U253 (N_253,In_20,In_128);
nand U254 (N_254,In_383,In_553);
or U255 (N_255,In_724,In_550);
and U256 (N_256,N_199,In_402);
xnor U257 (N_257,N_118,N_28);
and U258 (N_258,In_266,In_344);
nor U259 (N_259,In_378,In_474);
nand U260 (N_260,N_37,In_67);
or U261 (N_261,In_357,In_425);
and U262 (N_262,In_684,N_171);
nand U263 (N_263,In_298,N_87);
or U264 (N_264,In_734,In_690);
nand U265 (N_265,In_533,In_610);
and U266 (N_266,N_190,In_427);
nand U267 (N_267,N_142,N_91);
and U268 (N_268,In_426,In_111);
or U269 (N_269,In_428,In_578);
and U270 (N_270,In_406,In_289);
xnor U271 (N_271,In_412,In_450);
nor U272 (N_272,In_717,In_158);
nand U273 (N_273,N_164,In_423);
and U274 (N_274,In_741,In_543);
or U275 (N_275,In_370,In_249);
or U276 (N_276,In_524,N_112);
nor U277 (N_277,In_31,N_3);
or U278 (N_278,N_108,N_42);
xor U279 (N_279,In_99,In_733);
or U280 (N_280,In_385,In_420);
xor U281 (N_281,In_567,In_0);
or U282 (N_282,N_12,In_509);
and U283 (N_283,In_283,In_12);
nand U284 (N_284,N_198,In_434);
nor U285 (N_285,N_197,In_605);
nor U286 (N_286,In_230,In_287);
and U287 (N_287,N_79,In_388);
or U288 (N_288,In_541,N_123);
or U289 (N_289,In_707,In_432);
nor U290 (N_290,In_369,In_180);
nor U291 (N_291,In_311,In_3);
or U292 (N_292,In_694,N_68);
or U293 (N_293,In_348,In_535);
and U294 (N_294,In_215,In_174);
nor U295 (N_295,In_92,In_640);
and U296 (N_296,In_61,In_736);
nand U297 (N_297,In_303,In_368);
and U298 (N_298,N_146,In_331);
and U299 (N_299,In_695,In_482);
and U300 (N_300,In_356,In_238);
and U301 (N_301,In_325,N_13);
xor U302 (N_302,In_161,N_32);
nand U303 (N_303,In_47,N_221);
nand U304 (N_304,N_299,In_259);
nand U305 (N_305,N_39,N_202);
or U306 (N_306,N_74,N_61);
nand U307 (N_307,N_291,In_472);
nand U308 (N_308,N_35,N_292);
or U309 (N_309,In_176,In_607);
and U310 (N_310,In_556,N_7);
and U311 (N_311,N_288,N_135);
nand U312 (N_312,N_66,In_358);
or U313 (N_313,In_484,In_308);
nor U314 (N_314,N_238,N_64);
or U315 (N_315,N_111,N_281);
nor U316 (N_316,In_252,N_141);
nand U317 (N_317,In_22,In_421);
nor U318 (N_318,In_151,N_138);
or U319 (N_319,N_173,N_234);
nand U320 (N_320,In_347,N_147);
and U321 (N_321,In_159,In_45);
nand U322 (N_322,N_150,N_296);
nand U323 (N_323,N_266,N_132);
or U324 (N_324,In_49,In_148);
or U325 (N_325,N_268,In_386);
xnor U326 (N_326,N_279,In_473);
and U327 (N_327,N_59,N_203);
or U328 (N_328,N_119,N_200);
xnor U329 (N_329,In_518,N_216);
nand U330 (N_330,In_546,In_75);
and U331 (N_331,N_206,N_233);
nand U332 (N_332,N_252,In_343);
and U333 (N_333,In_39,N_51);
nor U334 (N_334,In_727,N_129);
nand U335 (N_335,In_467,N_162);
nor U336 (N_336,In_124,N_34);
xor U337 (N_337,N_263,In_193);
nor U338 (N_338,In_366,In_320);
and U339 (N_339,In_279,In_306);
and U340 (N_340,N_23,N_255);
nand U341 (N_341,N_294,In_379);
nor U342 (N_342,N_124,In_441);
and U343 (N_343,In_489,N_174);
nor U344 (N_344,In_218,In_569);
xor U345 (N_345,In_202,N_33);
xnor U346 (N_346,In_26,In_220);
nand U347 (N_347,In_207,N_151);
nor U348 (N_348,In_175,In_199);
xor U349 (N_349,In_228,In_531);
and U350 (N_350,In_332,In_372);
or U351 (N_351,In_583,In_547);
nor U352 (N_352,N_283,In_60);
xor U353 (N_353,In_495,N_77);
nand U354 (N_354,N_157,N_47);
and U355 (N_355,N_180,In_659);
and U356 (N_356,In_94,In_273);
and U357 (N_357,In_242,N_69);
xor U358 (N_358,In_699,N_5);
nand U359 (N_359,N_84,In_145);
nand U360 (N_360,N_217,N_259);
nand U361 (N_361,N_205,In_579);
nor U362 (N_362,N_253,In_413);
and U363 (N_363,In_274,N_176);
nor U364 (N_364,In_557,In_323);
xnor U365 (N_365,N_215,N_103);
nor U366 (N_366,In_261,In_72);
xnor U367 (N_367,N_71,In_46);
xor U368 (N_368,In_731,In_305);
and U369 (N_369,In_702,N_228);
and U370 (N_370,In_137,In_478);
and U371 (N_371,In_271,N_54);
nor U372 (N_372,In_676,In_643);
nand U373 (N_373,N_168,In_85);
and U374 (N_374,N_240,N_78);
xor U375 (N_375,N_227,In_310);
and U376 (N_376,N_265,N_65);
nand U377 (N_377,N_148,N_184);
or U378 (N_378,N_297,In_729);
xor U379 (N_379,In_706,N_128);
nor U380 (N_380,In_548,N_167);
nor U381 (N_381,N_237,In_400);
nand U382 (N_382,In_83,N_140);
xnor U383 (N_383,In_74,N_133);
xor U384 (N_384,N_243,N_271);
nor U385 (N_385,N_86,N_286);
nor U386 (N_386,In_589,N_246);
nand U387 (N_387,N_115,N_159);
nor U388 (N_388,N_14,N_100);
and U389 (N_389,In_213,N_70);
and U390 (N_390,In_639,In_674);
and U391 (N_391,In_381,In_537);
nand U392 (N_392,N_214,In_21);
nand U393 (N_393,In_487,In_376);
nor U394 (N_394,In_486,In_334);
xor U395 (N_395,N_289,In_439);
or U396 (N_396,In_446,N_67);
nor U397 (N_397,N_149,N_275);
nand U398 (N_398,N_290,In_573);
nand U399 (N_399,In_618,N_165);
or U400 (N_400,N_101,N_192);
xor U401 (N_401,In_231,In_609);
or U402 (N_402,N_381,N_363);
and U403 (N_403,N_396,In_214);
nand U404 (N_404,In_178,In_476);
and U405 (N_405,N_229,N_63);
and U406 (N_406,N_326,In_196);
and U407 (N_407,In_186,In_95);
nand U408 (N_408,N_357,In_560);
nor U409 (N_409,N_332,N_122);
nor U410 (N_410,In_443,N_183);
and U411 (N_411,N_371,N_179);
and U412 (N_412,In_200,N_322);
or U413 (N_413,In_321,N_372);
nor U414 (N_414,In_270,In_744);
xnor U415 (N_415,N_52,N_56);
nor U416 (N_416,N_218,N_274);
nand U417 (N_417,N_280,N_97);
xnor U418 (N_418,N_273,N_232);
nand U419 (N_419,In_669,In_245);
or U420 (N_420,N_143,In_593);
nand U421 (N_421,N_373,N_96);
nor U422 (N_422,N_316,N_60);
or U423 (N_423,N_204,In_590);
or U424 (N_424,N_113,N_210);
xnor U425 (N_425,In_191,N_231);
xor U426 (N_426,N_376,N_305);
nand U427 (N_427,N_327,N_29);
nor U428 (N_428,In_168,N_117);
xnor U429 (N_429,In_223,In_685);
or U430 (N_430,N_15,In_300);
nand U431 (N_431,N_394,N_339);
or U432 (N_432,In_675,N_258);
or U433 (N_433,In_419,In_156);
nand U434 (N_434,In_296,N_248);
nand U435 (N_435,N_107,N_393);
and U436 (N_436,N_312,N_20);
nand U437 (N_437,In_203,N_99);
and U438 (N_438,N_211,N_110);
or U439 (N_439,In_162,N_359);
xor U440 (N_440,N_222,In_91);
nor U441 (N_441,In_492,N_11);
xnor U442 (N_442,In_662,N_313);
xnor U443 (N_443,N_249,N_19);
nand U444 (N_444,In_52,N_336);
nand U445 (N_445,N_340,N_317);
or U446 (N_446,N_350,N_385);
and U447 (N_447,N_43,N_194);
or U448 (N_448,In_602,In_93);
xor U449 (N_449,N_378,N_310);
nand U450 (N_450,N_364,N_309);
nand U451 (N_451,In_455,In_584);
or U452 (N_452,N_379,N_349);
and U453 (N_453,N_342,N_177);
or U454 (N_454,In_253,N_374);
xnor U455 (N_455,In_285,In_525);
nor U456 (N_456,N_302,In_100);
or U457 (N_457,In_658,In_105);
xnor U458 (N_458,In_571,N_308);
nand U459 (N_459,N_241,N_382);
or U460 (N_460,In_691,N_195);
or U461 (N_461,N_182,N_347);
or U462 (N_462,N_370,N_351);
nand U463 (N_463,N_10,N_315);
nand U464 (N_464,N_161,In_59);
or U465 (N_465,N_172,N_366);
xor U466 (N_466,N_247,In_469);
or U467 (N_467,N_144,N_166);
and U468 (N_468,In_342,N_334);
and U469 (N_469,N_300,N_276);
nor U470 (N_470,In_167,N_337);
nand U471 (N_471,In_726,In_9);
or U472 (N_472,N_272,In_183);
or U473 (N_473,N_367,N_83);
nand U474 (N_474,In_255,N_354);
nand U475 (N_475,In_577,N_387);
or U476 (N_476,In_393,In_229);
and U477 (N_477,N_348,N_356);
and U478 (N_478,N_377,N_345);
nor U479 (N_479,N_239,N_224);
nor U480 (N_480,In_41,N_225);
and U481 (N_481,N_126,N_353);
or U482 (N_482,In_314,N_220);
nor U483 (N_483,In_349,N_295);
xnor U484 (N_484,N_72,N_196);
nand U485 (N_485,N_304,N_170);
nor U486 (N_486,In_485,In_315);
nor U487 (N_487,N_257,N_329);
xor U488 (N_488,N_397,N_355);
xor U489 (N_489,N_213,N_344);
nor U490 (N_490,N_298,N_331);
nor U491 (N_491,N_311,N_321);
or U492 (N_492,N_391,In_365);
and U493 (N_493,In_78,N_175);
or U494 (N_494,In_338,N_125);
xor U495 (N_495,In_564,In_319);
nor U496 (N_496,N_104,N_169);
or U497 (N_497,N_181,N_267);
nand U498 (N_498,N_223,In_104);
or U499 (N_499,In_634,N_365);
nand U500 (N_500,N_136,In_654);
or U501 (N_501,N_346,N_201);
and U502 (N_502,N_380,N_398);
or U503 (N_503,In_155,N_453);
nand U504 (N_504,N_325,N_486);
or U505 (N_505,In_64,N_368);
nor U506 (N_506,In_277,N_264);
or U507 (N_507,N_493,In_84);
or U508 (N_508,In_25,N_460);
nand U509 (N_509,N_287,N_335);
nand U510 (N_510,N_341,N_260);
xnor U511 (N_511,N_423,N_496);
nor U512 (N_512,N_375,N_405);
or U513 (N_513,N_474,N_278);
or U514 (N_514,In_136,N_109);
nand U515 (N_515,N_293,N_388);
or U516 (N_516,N_441,N_130);
xnor U517 (N_517,In_125,N_207);
nand U518 (N_518,N_481,N_465);
nor U519 (N_519,N_408,In_262);
nor U520 (N_520,N_434,N_450);
and U521 (N_521,N_429,N_383);
nand U522 (N_522,N_358,N_50);
and U523 (N_523,N_417,N_156);
nand U524 (N_524,N_438,N_361);
nand U525 (N_525,N_414,N_484);
nand U526 (N_526,N_328,N_256);
and U527 (N_527,N_473,N_134);
or U528 (N_528,N_462,In_147);
nor U529 (N_529,N_319,N_468);
or U530 (N_530,N_424,N_457);
or U531 (N_531,N_235,In_54);
or U532 (N_532,N_422,N_419);
nor U533 (N_533,In_598,N_485);
xnor U534 (N_534,N_284,N_320);
and U535 (N_535,N_4,In_146);
nand U536 (N_536,N_40,N_245);
nand U537 (N_537,N_446,N_212);
xnor U538 (N_538,N_230,N_73);
or U539 (N_539,In_449,N_187);
nand U540 (N_540,N_282,N_421);
or U541 (N_541,N_492,In_710);
nor U542 (N_542,In_80,N_458);
and U543 (N_543,In_692,N_412);
or U544 (N_544,N_55,N_389);
and U545 (N_545,N_413,In_198);
nand U546 (N_546,N_226,N_490);
and U547 (N_547,N_303,N_435);
xnor U548 (N_548,N_415,N_437);
or U549 (N_549,N_470,N_219);
nor U550 (N_550,N_6,N_121);
nand U551 (N_551,N_244,N_467);
or U552 (N_552,N_324,N_440);
and U553 (N_553,N_476,In_689);
nand U554 (N_554,N_25,N_452);
nor U555 (N_555,N_208,N_487);
nand U556 (N_556,N_480,N_475);
nand U557 (N_557,N_323,N_403);
nand U558 (N_558,In_735,N_426);
nand U559 (N_559,N_461,N_343);
and U560 (N_560,N_269,In_422);
nor U561 (N_561,In_728,In_457);
xnor U562 (N_562,N_436,N_352);
or U563 (N_563,In_133,N_410);
xor U564 (N_564,N_0,N_445);
and U565 (N_565,N_499,N_406);
xnor U566 (N_566,N_392,In_418);
and U567 (N_567,N_463,N_464);
nor U568 (N_568,N_98,N_186);
nor U569 (N_569,In_672,N_236);
or U570 (N_570,N_442,In_740);
and U571 (N_571,N_444,In_447);
nor U572 (N_572,N_400,In_513);
or U573 (N_573,N_449,N_131);
nand U574 (N_574,N_477,N_430);
and U575 (N_575,In_284,In_401);
xor U576 (N_576,N_451,N_285);
and U577 (N_577,N_185,N_395);
nand U578 (N_578,N_209,N_251);
and U579 (N_579,N_407,In_414);
or U580 (N_580,N_416,N_433);
and U581 (N_581,In_97,N_455);
nand U582 (N_582,N_447,N_270);
xor U583 (N_583,N_152,In_642);
and U584 (N_584,In_336,N_254);
or U585 (N_585,N_262,N_472);
or U586 (N_586,N_191,In_626);
xnor U587 (N_587,N_401,In_260);
and U588 (N_588,N_390,N_469);
or U589 (N_589,N_431,N_498);
and U590 (N_590,N_250,N_411);
and U591 (N_591,N_491,N_307);
nor U592 (N_592,N_314,N_338);
nand U593 (N_593,N_386,N_242);
xor U594 (N_594,N_102,N_360);
nand U595 (N_595,N_456,In_698);
and U596 (N_596,N_277,N_494);
and U597 (N_597,N_301,In_4);
xor U598 (N_598,N_427,In_636);
and U599 (N_599,N_428,N_443);
nor U600 (N_600,N_524,N_525);
nand U601 (N_601,N_550,N_483);
xnor U602 (N_602,N_548,N_553);
and U603 (N_603,N_333,N_589);
nand U604 (N_604,N_564,In_463);
nor U605 (N_605,N_512,N_591);
nor U606 (N_606,In_312,N_561);
and U607 (N_607,N_478,N_479);
and U608 (N_608,N_544,N_516);
and U609 (N_609,N_513,N_1);
nand U610 (N_610,N_559,N_570);
and U611 (N_611,N_552,N_555);
or U612 (N_612,N_261,N_523);
and U613 (N_613,N_409,N_585);
or U614 (N_614,N_576,N_106);
nor U615 (N_615,N_511,N_558);
or U616 (N_616,N_466,N_532);
or U617 (N_617,N_563,N_569);
or U618 (N_618,N_540,N_535);
nor U619 (N_619,In_517,N_542);
nor U620 (N_620,N_592,In_371);
or U621 (N_621,In_644,N_584);
xnor U622 (N_622,N_536,N_556);
nand U623 (N_623,N_598,N_515);
or U624 (N_624,N_547,N_574);
nor U625 (N_625,N_541,N_509);
or U626 (N_626,N_579,In_166);
or U627 (N_627,In_359,N_578);
or U628 (N_628,N_521,N_565);
nor U629 (N_629,N_554,In_466);
and U630 (N_630,N_562,N_384);
nand U631 (N_631,N_573,N_420);
and U632 (N_632,N_588,N_567);
nand U633 (N_633,N_551,N_514);
nand U634 (N_634,N_418,N_549);
or U635 (N_635,N_526,N_575);
and U636 (N_636,N_505,N_543);
and U637 (N_637,N_501,N_580);
nor U638 (N_638,N_594,N_318);
and U639 (N_639,N_507,N_432);
nor U640 (N_640,N_529,N_572);
and U641 (N_641,N_362,N_510);
and U642 (N_642,N_582,N_503);
or U643 (N_643,N_399,N_571);
and U644 (N_644,N_528,N_587);
nor U645 (N_645,N_189,N_577);
nor U646 (N_646,N_522,In_88);
nand U647 (N_647,N_402,N_497);
or U648 (N_648,N_404,N_471);
xor U649 (N_649,N_519,N_527);
and U650 (N_650,N_500,N_506);
nand U651 (N_651,N_596,N_586);
and U652 (N_652,In_29,N_581);
nor U653 (N_653,N_504,N_545);
nor U654 (N_654,N_425,N_531);
nor U655 (N_655,N_537,N_520);
nor U656 (N_656,N_508,N_369);
and U657 (N_657,N_534,N_330);
nor U658 (N_658,N_533,N_595);
and U659 (N_659,N_439,N_590);
and U660 (N_660,N_306,N_518);
and U661 (N_661,N_454,N_482);
or U662 (N_662,In_346,N_546);
or U663 (N_663,N_489,N_538);
xor U664 (N_664,In_189,N_495);
nor U665 (N_665,N_517,N_448);
or U666 (N_666,N_488,In_116);
or U667 (N_667,In_522,N_599);
nand U668 (N_668,In_647,N_502);
and U669 (N_669,N_566,N_459);
and U670 (N_670,N_597,N_530);
or U671 (N_671,N_568,N_62);
and U672 (N_672,N_583,N_105);
xnor U673 (N_673,N_560,N_539);
nand U674 (N_674,N_557,N_593);
nand U675 (N_675,N_537,N_583);
xor U676 (N_676,N_594,N_579);
nor U677 (N_677,N_540,N_572);
nand U678 (N_678,N_532,N_330);
nand U679 (N_679,N_432,N_556);
or U680 (N_680,N_598,N_595);
and U681 (N_681,In_647,N_545);
and U682 (N_682,N_577,N_525);
and U683 (N_683,N_570,In_312);
or U684 (N_684,N_509,N_540);
and U685 (N_685,N_333,N_538);
nand U686 (N_686,N_471,N_533);
nand U687 (N_687,N_591,N_532);
xor U688 (N_688,In_371,N_409);
nand U689 (N_689,N_540,N_553);
nor U690 (N_690,N_369,N_512);
xnor U691 (N_691,N_560,N_579);
or U692 (N_692,N_526,N_536);
nand U693 (N_693,In_371,N_594);
nor U694 (N_694,N_514,N_566);
nor U695 (N_695,N_544,N_521);
or U696 (N_696,N_599,N_479);
xnor U697 (N_697,N_569,N_525);
xnor U698 (N_698,N_106,N_581);
nor U699 (N_699,N_594,N_597);
or U700 (N_700,N_651,N_688);
and U701 (N_701,N_690,N_658);
nor U702 (N_702,N_653,N_610);
and U703 (N_703,N_633,N_616);
nand U704 (N_704,N_642,N_606);
nor U705 (N_705,N_686,N_601);
and U706 (N_706,N_655,N_685);
xnor U707 (N_707,N_695,N_649);
nor U708 (N_708,N_613,N_634);
or U709 (N_709,N_692,N_630);
nand U710 (N_710,N_632,N_609);
nor U711 (N_711,N_624,N_672);
and U712 (N_712,N_693,N_665);
nor U713 (N_713,N_683,N_619);
and U714 (N_714,N_660,N_622);
or U715 (N_715,N_694,N_643);
nor U716 (N_716,N_679,N_618);
or U717 (N_717,N_627,N_620);
nand U718 (N_718,N_607,N_659);
nor U719 (N_719,N_696,N_639);
nor U720 (N_720,N_645,N_675);
nor U721 (N_721,N_623,N_628);
nor U722 (N_722,N_625,N_641);
nor U723 (N_723,N_611,N_677);
or U724 (N_724,N_614,N_650);
nand U725 (N_725,N_603,N_662);
nand U726 (N_726,N_637,N_698);
or U727 (N_727,N_654,N_663);
nor U728 (N_728,N_644,N_681);
and U729 (N_729,N_669,N_647);
nand U730 (N_730,N_699,N_668);
nor U731 (N_731,N_676,N_682);
nor U732 (N_732,N_612,N_648);
or U733 (N_733,N_657,N_600);
or U734 (N_734,N_661,N_678);
nand U735 (N_735,N_697,N_671);
and U736 (N_736,N_640,N_656);
nand U737 (N_737,N_689,N_635);
nand U738 (N_738,N_626,N_673);
nor U739 (N_739,N_615,N_666);
nor U740 (N_740,N_664,N_617);
nand U741 (N_741,N_608,N_680);
and U742 (N_742,N_605,N_638);
nor U743 (N_743,N_629,N_602);
and U744 (N_744,N_636,N_674);
or U745 (N_745,N_667,N_691);
nand U746 (N_746,N_604,N_687);
or U747 (N_747,N_646,N_652);
nand U748 (N_748,N_670,N_631);
or U749 (N_749,N_621,N_684);
and U750 (N_750,N_669,N_624);
nor U751 (N_751,N_683,N_691);
or U752 (N_752,N_697,N_695);
and U753 (N_753,N_680,N_658);
xnor U754 (N_754,N_647,N_682);
and U755 (N_755,N_678,N_673);
nand U756 (N_756,N_607,N_674);
and U757 (N_757,N_624,N_645);
nand U758 (N_758,N_695,N_604);
or U759 (N_759,N_616,N_638);
and U760 (N_760,N_662,N_665);
nand U761 (N_761,N_631,N_662);
xnor U762 (N_762,N_677,N_696);
nand U763 (N_763,N_682,N_691);
nor U764 (N_764,N_698,N_628);
nor U765 (N_765,N_667,N_675);
nand U766 (N_766,N_685,N_635);
or U767 (N_767,N_648,N_674);
nor U768 (N_768,N_684,N_642);
nor U769 (N_769,N_664,N_627);
nor U770 (N_770,N_698,N_612);
nand U771 (N_771,N_639,N_629);
or U772 (N_772,N_603,N_634);
nor U773 (N_773,N_683,N_672);
or U774 (N_774,N_694,N_601);
xnor U775 (N_775,N_664,N_686);
nor U776 (N_776,N_686,N_690);
and U777 (N_777,N_638,N_606);
nor U778 (N_778,N_617,N_609);
and U779 (N_779,N_691,N_673);
or U780 (N_780,N_628,N_608);
or U781 (N_781,N_660,N_668);
nor U782 (N_782,N_672,N_679);
and U783 (N_783,N_667,N_611);
nor U784 (N_784,N_645,N_642);
and U785 (N_785,N_633,N_648);
or U786 (N_786,N_642,N_643);
xnor U787 (N_787,N_634,N_665);
nand U788 (N_788,N_647,N_632);
or U789 (N_789,N_604,N_655);
and U790 (N_790,N_688,N_637);
nand U791 (N_791,N_667,N_681);
and U792 (N_792,N_649,N_638);
nand U793 (N_793,N_657,N_647);
and U794 (N_794,N_644,N_626);
and U795 (N_795,N_681,N_664);
nor U796 (N_796,N_612,N_633);
and U797 (N_797,N_699,N_633);
nor U798 (N_798,N_649,N_675);
or U799 (N_799,N_657,N_698);
xor U800 (N_800,N_727,N_740);
and U801 (N_801,N_795,N_700);
or U802 (N_802,N_746,N_707);
or U803 (N_803,N_733,N_799);
and U804 (N_804,N_713,N_774);
nand U805 (N_805,N_716,N_770);
nor U806 (N_806,N_750,N_798);
or U807 (N_807,N_715,N_741);
nor U808 (N_808,N_734,N_737);
and U809 (N_809,N_759,N_724);
nor U810 (N_810,N_708,N_714);
nor U811 (N_811,N_794,N_767);
nor U812 (N_812,N_756,N_703);
xnor U813 (N_813,N_764,N_753);
and U814 (N_814,N_717,N_728);
nand U815 (N_815,N_791,N_785);
nor U816 (N_816,N_783,N_796);
nand U817 (N_817,N_712,N_787);
or U818 (N_818,N_718,N_769);
and U819 (N_819,N_705,N_771);
nor U820 (N_820,N_710,N_789);
or U821 (N_821,N_719,N_722);
or U822 (N_822,N_720,N_736);
and U823 (N_823,N_721,N_779);
nor U824 (N_824,N_765,N_731);
or U825 (N_825,N_784,N_739);
or U826 (N_826,N_777,N_723);
and U827 (N_827,N_763,N_711);
nor U828 (N_828,N_773,N_778);
nand U829 (N_829,N_751,N_793);
or U830 (N_830,N_761,N_757);
and U831 (N_831,N_755,N_729);
xnor U832 (N_832,N_726,N_792);
xor U833 (N_833,N_776,N_744);
nand U834 (N_834,N_768,N_758);
nor U835 (N_835,N_775,N_742);
and U836 (N_836,N_760,N_747);
nor U837 (N_837,N_749,N_797);
nand U838 (N_838,N_743,N_754);
xor U839 (N_839,N_732,N_762);
and U840 (N_840,N_772,N_766);
nand U841 (N_841,N_738,N_780);
and U842 (N_842,N_745,N_752);
nor U843 (N_843,N_701,N_704);
or U844 (N_844,N_782,N_730);
nand U845 (N_845,N_709,N_735);
nand U846 (N_846,N_702,N_781);
or U847 (N_847,N_748,N_790);
or U848 (N_848,N_788,N_706);
nor U849 (N_849,N_786,N_725);
and U850 (N_850,N_789,N_709);
and U851 (N_851,N_711,N_719);
and U852 (N_852,N_728,N_745);
nor U853 (N_853,N_736,N_761);
nand U854 (N_854,N_792,N_786);
and U855 (N_855,N_764,N_703);
nand U856 (N_856,N_759,N_799);
nand U857 (N_857,N_722,N_711);
nand U858 (N_858,N_787,N_754);
nor U859 (N_859,N_782,N_742);
nand U860 (N_860,N_777,N_749);
nand U861 (N_861,N_706,N_796);
nor U862 (N_862,N_797,N_708);
or U863 (N_863,N_757,N_729);
and U864 (N_864,N_753,N_788);
nand U865 (N_865,N_754,N_759);
or U866 (N_866,N_765,N_738);
nor U867 (N_867,N_715,N_712);
or U868 (N_868,N_784,N_790);
and U869 (N_869,N_793,N_795);
and U870 (N_870,N_773,N_724);
or U871 (N_871,N_719,N_763);
nor U872 (N_872,N_763,N_757);
nand U873 (N_873,N_711,N_764);
nor U874 (N_874,N_700,N_777);
nor U875 (N_875,N_709,N_780);
and U876 (N_876,N_713,N_726);
and U877 (N_877,N_738,N_775);
or U878 (N_878,N_780,N_790);
or U879 (N_879,N_735,N_738);
nor U880 (N_880,N_710,N_768);
xor U881 (N_881,N_774,N_795);
xnor U882 (N_882,N_780,N_775);
and U883 (N_883,N_706,N_782);
nor U884 (N_884,N_771,N_764);
nor U885 (N_885,N_767,N_746);
or U886 (N_886,N_768,N_763);
and U887 (N_887,N_716,N_760);
and U888 (N_888,N_749,N_778);
and U889 (N_889,N_717,N_725);
nor U890 (N_890,N_775,N_710);
or U891 (N_891,N_719,N_750);
and U892 (N_892,N_742,N_723);
or U893 (N_893,N_709,N_746);
or U894 (N_894,N_765,N_727);
or U895 (N_895,N_766,N_794);
xnor U896 (N_896,N_764,N_704);
nor U897 (N_897,N_768,N_747);
nor U898 (N_898,N_769,N_786);
xor U899 (N_899,N_711,N_741);
or U900 (N_900,N_891,N_870);
and U901 (N_901,N_863,N_816);
xnor U902 (N_902,N_871,N_876);
and U903 (N_903,N_803,N_864);
and U904 (N_904,N_835,N_878);
nand U905 (N_905,N_853,N_860);
and U906 (N_906,N_857,N_859);
and U907 (N_907,N_837,N_800);
nand U908 (N_908,N_895,N_873);
nand U909 (N_909,N_802,N_889);
or U910 (N_910,N_882,N_825);
and U911 (N_911,N_804,N_810);
and U912 (N_912,N_832,N_849);
or U913 (N_913,N_828,N_894);
nor U914 (N_914,N_899,N_809);
nor U915 (N_915,N_884,N_807);
nand U916 (N_916,N_893,N_839);
nor U917 (N_917,N_836,N_898);
nand U918 (N_918,N_842,N_866);
nor U919 (N_919,N_879,N_813);
or U920 (N_920,N_872,N_818);
nor U921 (N_921,N_874,N_847);
and U922 (N_922,N_829,N_856);
nor U923 (N_923,N_848,N_812);
nor U924 (N_924,N_814,N_883);
nand U925 (N_925,N_888,N_892);
nand U926 (N_926,N_890,N_877);
and U927 (N_927,N_861,N_840);
nor U928 (N_928,N_831,N_801);
and U929 (N_929,N_886,N_881);
xnor U930 (N_930,N_820,N_819);
nand U931 (N_931,N_885,N_806);
or U932 (N_932,N_811,N_815);
and U933 (N_933,N_869,N_822);
nand U934 (N_934,N_851,N_875);
nand U935 (N_935,N_808,N_843);
and U936 (N_936,N_834,N_817);
nor U937 (N_937,N_846,N_887);
and U938 (N_938,N_826,N_824);
and U939 (N_939,N_827,N_850);
nor U940 (N_940,N_880,N_897);
or U941 (N_941,N_821,N_855);
and U942 (N_942,N_896,N_867);
or U943 (N_943,N_858,N_854);
nand U944 (N_944,N_865,N_844);
xor U945 (N_945,N_838,N_845);
xor U946 (N_946,N_868,N_852);
or U947 (N_947,N_823,N_862);
nand U948 (N_948,N_841,N_805);
nand U949 (N_949,N_833,N_830);
or U950 (N_950,N_804,N_873);
or U951 (N_951,N_809,N_812);
nor U952 (N_952,N_878,N_854);
nand U953 (N_953,N_839,N_834);
nand U954 (N_954,N_825,N_893);
and U955 (N_955,N_890,N_824);
or U956 (N_956,N_896,N_884);
or U957 (N_957,N_880,N_840);
nor U958 (N_958,N_837,N_895);
nand U959 (N_959,N_850,N_890);
nand U960 (N_960,N_813,N_872);
xnor U961 (N_961,N_847,N_867);
nor U962 (N_962,N_833,N_843);
nor U963 (N_963,N_849,N_810);
nor U964 (N_964,N_823,N_819);
nor U965 (N_965,N_883,N_868);
nand U966 (N_966,N_800,N_892);
or U967 (N_967,N_837,N_858);
nand U968 (N_968,N_846,N_849);
nand U969 (N_969,N_823,N_811);
or U970 (N_970,N_853,N_893);
and U971 (N_971,N_845,N_868);
nand U972 (N_972,N_885,N_861);
or U973 (N_973,N_878,N_852);
or U974 (N_974,N_833,N_876);
or U975 (N_975,N_869,N_818);
or U976 (N_976,N_836,N_839);
xor U977 (N_977,N_871,N_801);
xnor U978 (N_978,N_867,N_899);
or U979 (N_979,N_834,N_898);
or U980 (N_980,N_872,N_829);
nor U981 (N_981,N_887,N_837);
nor U982 (N_982,N_836,N_873);
xor U983 (N_983,N_841,N_821);
or U984 (N_984,N_842,N_861);
nor U985 (N_985,N_866,N_807);
or U986 (N_986,N_803,N_821);
nand U987 (N_987,N_802,N_883);
nand U988 (N_988,N_822,N_876);
and U989 (N_989,N_893,N_828);
or U990 (N_990,N_812,N_837);
and U991 (N_991,N_800,N_883);
nand U992 (N_992,N_854,N_859);
or U993 (N_993,N_899,N_817);
or U994 (N_994,N_809,N_877);
nor U995 (N_995,N_892,N_837);
and U996 (N_996,N_871,N_872);
nor U997 (N_997,N_893,N_845);
nand U998 (N_998,N_800,N_857);
or U999 (N_999,N_856,N_841);
xnor U1000 (N_1000,N_977,N_986);
xor U1001 (N_1001,N_960,N_990);
or U1002 (N_1002,N_930,N_934);
and U1003 (N_1003,N_979,N_944);
nand U1004 (N_1004,N_955,N_950);
nor U1005 (N_1005,N_971,N_903);
nand U1006 (N_1006,N_943,N_993);
and U1007 (N_1007,N_921,N_953);
nor U1008 (N_1008,N_969,N_909);
nand U1009 (N_1009,N_965,N_905);
or U1010 (N_1010,N_954,N_985);
nor U1011 (N_1011,N_920,N_913);
or U1012 (N_1012,N_992,N_927);
and U1013 (N_1013,N_972,N_932);
nand U1014 (N_1014,N_975,N_962);
nand U1015 (N_1015,N_918,N_973);
or U1016 (N_1016,N_931,N_904);
and U1017 (N_1017,N_906,N_947);
or U1018 (N_1018,N_945,N_938);
and U1019 (N_1019,N_958,N_933);
xor U1020 (N_1020,N_901,N_937);
and U1021 (N_1021,N_956,N_939);
and U1022 (N_1022,N_961,N_968);
and U1023 (N_1023,N_967,N_998);
nor U1024 (N_1024,N_959,N_995);
xnor U1025 (N_1025,N_970,N_974);
nand U1026 (N_1026,N_942,N_989);
or U1027 (N_1027,N_987,N_925);
and U1028 (N_1028,N_949,N_908);
and U1029 (N_1029,N_928,N_902);
and U1030 (N_1030,N_923,N_984);
xor U1031 (N_1031,N_917,N_935);
or U1032 (N_1032,N_994,N_952);
and U1033 (N_1033,N_900,N_951);
nor U1034 (N_1034,N_991,N_978);
nand U1035 (N_1035,N_999,N_924);
and U1036 (N_1036,N_996,N_983);
or U1037 (N_1037,N_976,N_919);
nor U1038 (N_1038,N_914,N_915);
nor U1039 (N_1039,N_916,N_910);
or U1040 (N_1040,N_980,N_911);
nand U1041 (N_1041,N_982,N_926);
or U1042 (N_1042,N_957,N_936);
nand U1043 (N_1043,N_988,N_912);
and U1044 (N_1044,N_966,N_964);
xor U1045 (N_1045,N_963,N_948);
xnor U1046 (N_1046,N_997,N_941);
and U1047 (N_1047,N_981,N_907);
or U1048 (N_1048,N_929,N_946);
or U1049 (N_1049,N_940,N_922);
and U1050 (N_1050,N_936,N_959);
or U1051 (N_1051,N_906,N_920);
or U1052 (N_1052,N_964,N_995);
and U1053 (N_1053,N_973,N_901);
nor U1054 (N_1054,N_980,N_934);
xor U1055 (N_1055,N_984,N_930);
and U1056 (N_1056,N_945,N_964);
and U1057 (N_1057,N_929,N_921);
and U1058 (N_1058,N_993,N_936);
or U1059 (N_1059,N_984,N_974);
nor U1060 (N_1060,N_962,N_945);
nor U1061 (N_1061,N_964,N_901);
nand U1062 (N_1062,N_910,N_911);
nand U1063 (N_1063,N_932,N_975);
xnor U1064 (N_1064,N_904,N_943);
nand U1065 (N_1065,N_962,N_980);
nor U1066 (N_1066,N_919,N_957);
or U1067 (N_1067,N_980,N_957);
nand U1068 (N_1068,N_912,N_950);
or U1069 (N_1069,N_927,N_991);
nand U1070 (N_1070,N_988,N_907);
and U1071 (N_1071,N_971,N_926);
nand U1072 (N_1072,N_950,N_966);
xor U1073 (N_1073,N_996,N_916);
and U1074 (N_1074,N_961,N_959);
nor U1075 (N_1075,N_905,N_917);
nand U1076 (N_1076,N_944,N_999);
nand U1077 (N_1077,N_962,N_956);
nor U1078 (N_1078,N_981,N_989);
nor U1079 (N_1079,N_921,N_900);
nand U1080 (N_1080,N_957,N_902);
nor U1081 (N_1081,N_913,N_995);
xnor U1082 (N_1082,N_958,N_999);
and U1083 (N_1083,N_910,N_941);
or U1084 (N_1084,N_975,N_922);
xor U1085 (N_1085,N_995,N_991);
nand U1086 (N_1086,N_904,N_920);
nand U1087 (N_1087,N_985,N_968);
nand U1088 (N_1088,N_951,N_996);
nor U1089 (N_1089,N_951,N_912);
or U1090 (N_1090,N_923,N_903);
nor U1091 (N_1091,N_944,N_940);
or U1092 (N_1092,N_957,N_948);
or U1093 (N_1093,N_962,N_951);
nor U1094 (N_1094,N_975,N_926);
or U1095 (N_1095,N_978,N_948);
nand U1096 (N_1096,N_933,N_914);
and U1097 (N_1097,N_934,N_990);
or U1098 (N_1098,N_917,N_953);
nand U1099 (N_1099,N_983,N_967);
nand U1100 (N_1100,N_1033,N_1093);
or U1101 (N_1101,N_1006,N_1084);
or U1102 (N_1102,N_1041,N_1040);
nand U1103 (N_1103,N_1024,N_1014);
nor U1104 (N_1104,N_1028,N_1065);
or U1105 (N_1105,N_1052,N_1050);
or U1106 (N_1106,N_1005,N_1077);
and U1107 (N_1107,N_1001,N_1009);
nand U1108 (N_1108,N_1059,N_1020);
and U1109 (N_1109,N_1025,N_1067);
and U1110 (N_1110,N_1056,N_1079);
nor U1111 (N_1111,N_1000,N_1090);
nand U1112 (N_1112,N_1029,N_1013);
nand U1113 (N_1113,N_1082,N_1073);
xor U1114 (N_1114,N_1034,N_1046);
or U1115 (N_1115,N_1002,N_1018);
and U1116 (N_1116,N_1030,N_1016);
nor U1117 (N_1117,N_1088,N_1089);
nor U1118 (N_1118,N_1064,N_1061);
nor U1119 (N_1119,N_1031,N_1091);
and U1120 (N_1120,N_1078,N_1095);
nand U1121 (N_1121,N_1045,N_1021);
nor U1122 (N_1122,N_1081,N_1060);
nor U1123 (N_1123,N_1037,N_1043);
and U1124 (N_1124,N_1074,N_1069);
or U1125 (N_1125,N_1097,N_1012);
nor U1126 (N_1126,N_1083,N_1054);
or U1127 (N_1127,N_1008,N_1026);
nand U1128 (N_1128,N_1098,N_1068);
nor U1129 (N_1129,N_1072,N_1076);
and U1130 (N_1130,N_1055,N_1011);
xor U1131 (N_1131,N_1007,N_1051);
and U1132 (N_1132,N_1071,N_1003);
or U1133 (N_1133,N_1062,N_1010);
and U1134 (N_1134,N_1048,N_1038);
and U1135 (N_1135,N_1053,N_1015);
or U1136 (N_1136,N_1085,N_1080);
nand U1137 (N_1137,N_1044,N_1087);
or U1138 (N_1138,N_1017,N_1032);
or U1139 (N_1139,N_1070,N_1049);
and U1140 (N_1140,N_1066,N_1099);
nand U1141 (N_1141,N_1022,N_1035);
and U1142 (N_1142,N_1042,N_1004);
xor U1143 (N_1143,N_1036,N_1096);
xnor U1144 (N_1144,N_1092,N_1058);
nand U1145 (N_1145,N_1023,N_1086);
and U1146 (N_1146,N_1094,N_1075);
xor U1147 (N_1147,N_1027,N_1019);
or U1148 (N_1148,N_1039,N_1063);
nand U1149 (N_1149,N_1057,N_1047);
and U1150 (N_1150,N_1094,N_1061);
nand U1151 (N_1151,N_1009,N_1008);
nand U1152 (N_1152,N_1027,N_1097);
or U1153 (N_1153,N_1098,N_1053);
nand U1154 (N_1154,N_1003,N_1094);
xnor U1155 (N_1155,N_1044,N_1002);
nor U1156 (N_1156,N_1007,N_1088);
or U1157 (N_1157,N_1067,N_1030);
nand U1158 (N_1158,N_1093,N_1099);
or U1159 (N_1159,N_1051,N_1095);
or U1160 (N_1160,N_1023,N_1008);
and U1161 (N_1161,N_1015,N_1051);
nand U1162 (N_1162,N_1097,N_1083);
nand U1163 (N_1163,N_1062,N_1089);
and U1164 (N_1164,N_1088,N_1010);
nand U1165 (N_1165,N_1026,N_1000);
nor U1166 (N_1166,N_1004,N_1098);
nor U1167 (N_1167,N_1056,N_1039);
nor U1168 (N_1168,N_1021,N_1097);
nor U1169 (N_1169,N_1042,N_1051);
nand U1170 (N_1170,N_1023,N_1069);
nand U1171 (N_1171,N_1059,N_1040);
and U1172 (N_1172,N_1017,N_1009);
nand U1173 (N_1173,N_1075,N_1078);
or U1174 (N_1174,N_1027,N_1021);
nor U1175 (N_1175,N_1000,N_1086);
nand U1176 (N_1176,N_1038,N_1053);
and U1177 (N_1177,N_1048,N_1077);
or U1178 (N_1178,N_1012,N_1083);
and U1179 (N_1179,N_1069,N_1040);
nand U1180 (N_1180,N_1043,N_1026);
or U1181 (N_1181,N_1005,N_1003);
and U1182 (N_1182,N_1056,N_1010);
or U1183 (N_1183,N_1042,N_1095);
xnor U1184 (N_1184,N_1000,N_1041);
nor U1185 (N_1185,N_1015,N_1005);
and U1186 (N_1186,N_1009,N_1012);
and U1187 (N_1187,N_1009,N_1061);
xnor U1188 (N_1188,N_1047,N_1024);
xnor U1189 (N_1189,N_1096,N_1024);
or U1190 (N_1190,N_1095,N_1067);
and U1191 (N_1191,N_1021,N_1007);
nand U1192 (N_1192,N_1052,N_1084);
nand U1193 (N_1193,N_1064,N_1025);
and U1194 (N_1194,N_1003,N_1096);
nand U1195 (N_1195,N_1087,N_1011);
nand U1196 (N_1196,N_1059,N_1083);
nand U1197 (N_1197,N_1060,N_1088);
nor U1198 (N_1198,N_1019,N_1046);
nor U1199 (N_1199,N_1035,N_1011);
and U1200 (N_1200,N_1140,N_1149);
nor U1201 (N_1201,N_1133,N_1130);
nor U1202 (N_1202,N_1181,N_1173);
nand U1203 (N_1203,N_1192,N_1103);
xnor U1204 (N_1204,N_1137,N_1144);
nand U1205 (N_1205,N_1152,N_1110);
nor U1206 (N_1206,N_1113,N_1172);
or U1207 (N_1207,N_1163,N_1179);
xor U1208 (N_1208,N_1124,N_1125);
nand U1209 (N_1209,N_1114,N_1115);
or U1210 (N_1210,N_1197,N_1128);
nor U1211 (N_1211,N_1117,N_1198);
and U1212 (N_1212,N_1101,N_1146);
and U1213 (N_1213,N_1112,N_1199);
or U1214 (N_1214,N_1184,N_1142);
nor U1215 (N_1215,N_1136,N_1161);
and U1216 (N_1216,N_1190,N_1127);
and U1217 (N_1217,N_1119,N_1196);
nor U1218 (N_1218,N_1121,N_1174);
nand U1219 (N_1219,N_1194,N_1132);
nand U1220 (N_1220,N_1153,N_1164);
nand U1221 (N_1221,N_1175,N_1151);
or U1222 (N_1222,N_1176,N_1170);
nand U1223 (N_1223,N_1191,N_1131);
xor U1224 (N_1224,N_1193,N_1143);
nor U1225 (N_1225,N_1189,N_1150);
xnor U1226 (N_1226,N_1129,N_1148);
or U1227 (N_1227,N_1182,N_1177);
nand U1228 (N_1228,N_1102,N_1158);
nand U1229 (N_1229,N_1116,N_1118);
nand U1230 (N_1230,N_1168,N_1155);
and U1231 (N_1231,N_1109,N_1123);
nand U1232 (N_1232,N_1162,N_1145);
nor U1233 (N_1233,N_1167,N_1139);
and U1234 (N_1234,N_1165,N_1147);
or U1235 (N_1235,N_1156,N_1135);
or U1236 (N_1236,N_1188,N_1141);
and U1237 (N_1237,N_1154,N_1178);
nand U1238 (N_1238,N_1108,N_1120);
xnor U1239 (N_1239,N_1186,N_1157);
nor U1240 (N_1240,N_1195,N_1169);
nand U1241 (N_1241,N_1166,N_1160);
nand U1242 (N_1242,N_1185,N_1100);
nor U1243 (N_1243,N_1107,N_1187);
and U1244 (N_1244,N_1159,N_1106);
or U1245 (N_1245,N_1122,N_1104);
nand U1246 (N_1246,N_1111,N_1134);
xnor U1247 (N_1247,N_1183,N_1138);
and U1248 (N_1248,N_1105,N_1180);
and U1249 (N_1249,N_1171,N_1126);
nand U1250 (N_1250,N_1109,N_1190);
and U1251 (N_1251,N_1123,N_1164);
nor U1252 (N_1252,N_1112,N_1142);
nand U1253 (N_1253,N_1160,N_1111);
and U1254 (N_1254,N_1129,N_1186);
or U1255 (N_1255,N_1169,N_1188);
nor U1256 (N_1256,N_1100,N_1195);
and U1257 (N_1257,N_1129,N_1175);
nor U1258 (N_1258,N_1115,N_1165);
and U1259 (N_1259,N_1109,N_1162);
nand U1260 (N_1260,N_1178,N_1116);
nor U1261 (N_1261,N_1193,N_1186);
or U1262 (N_1262,N_1128,N_1184);
nand U1263 (N_1263,N_1142,N_1179);
or U1264 (N_1264,N_1139,N_1180);
and U1265 (N_1265,N_1119,N_1101);
nand U1266 (N_1266,N_1161,N_1164);
xnor U1267 (N_1267,N_1176,N_1123);
nand U1268 (N_1268,N_1102,N_1134);
and U1269 (N_1269,N_1136,N_1107);
nor U1270 (N_1270,N_1185,N_1198);
nand U1271 (N_1271,N_1190,N_1178);
nor U1272 (N_1272,N_1180,N_1182);
nand U1273 (N_1273,N_1100,N_1122);
nor U1274 (N_1274,N_1152,N_1131);
xnor U1275 (N_1275,N_1185,N_1174);
nand U1276 (N_1276,N_1176,N_1180);
and U1277 (N_1277,N_1166,N_1150);
or U1278 (N_1278,N_1135,N_1120);
nand U1279 (N_1279,N_1160,N_1165);
nor U1280 (N_1280,N_1139,N_1122);
and U1281 (N_1281,N_1183,N_1127);
or U1282 (N_1282,N_1110,N_1119);
or U1283 (N_1283,N_1157,N_1143);
nor U1284 (N_1284,N_1122,N_1172);
or U1285 (N_1285,N_1146,N_1153);
or U1286 (N_1286,N_1169,N_1135);
and U1287 (N_1287,N_1157,N_1118);
nor U1288 (N_1288,N_1153,N_1133);
and U1289 (N_1289,N_1180,N_1173);
nand U1290 (N_1290,N_1183,N_1120);
nand U1291 (N_1291,N_1126,N_1117);
nand U1292 (N_1292,N_1187,N_1199);
or U1293 (N_1293,N_1173,N_1101);
or U1294 (N_1294,N_1199,N_1134);
nand U1295 (N_1295,N_1171,N_1124);
or U1296 (N_1296,N_1171,N_1182);
xnor U1297 (N_1297,N_1168,N_1144);
xor U1298 (N_1298,N_1148,N_1178);
xnor U1299 (N_1299,N_1107,N_1188);
nand U1300 (N_1300,N_1204,N_1234);
or U1301 (N_1301,N_1295,N_1296);
nor U1302 (N_1302,N_1228,N_1220);
or U1303 (N_1303,N_1294,N_1217);
or U1304 (N_1304,N_1230,N_1209);
nand U1305 (N_1305,N_1264,N_1221);
nand U1306 (N_1306,N_1243,N_1258);
or U1307 (N_1307,N_1298,N_1200);
and U1308 (N_1308,N_1259,N_1244);
nor U1309 (N_1309,N_1267,N_1212);
xor U1310 (N_1310,N_1246,N_1208);
nor U1311 (N_1311,N_1292,N_1253);
nor U1312 (N_1312,N_1242,N_1250);
or U1313 (N_1313,N_1260,N_1222);
nor U1314 (N_1314,N_1238,N_1269);
nor U1315 (N_1315,N_1203,N_1299);
nor U1316 (N_1316,N_1290,N_1249);
nor U1317 (N_1317,N_1287,N_1241);
nor U1318 (N_1318,N_1233,N_1285);
nor U1319 (N_1319,N_1207,N_1236);
xor U1320 (N_1320,N_1276,N_1237);
or U1321 (N_1321,N_1291,N_1279);
xnor U1322 (N_1322,N_1274,N_1235);
nand U1323 (N_1323,N_1213,N_1286);
nand U1324 (N_1324,N_1265,N_1293);
nor U1325 (N_1325,N_1229,N_1262);
nand U1326 (N_1326,N_1211,N_1263);
xnor U1327 (N_1327,N_1210,N_1215);
or U1328 (N_1328,N_1257,N_1232);
and U1329 (N_1329,N_1281,N_1270);
or U1330 (N_1330,N_1261,N_1283);
xor U1331 (N_1331,N_1218,N_1214);
nand U1332 (N_1332,N_1272,N_1273);
and U1333 (N_1333,N_1248,N_1288);
and U1334 (N_1334,N_1206,N_1266);
and U1335 (N_1335,N_1202,N_1239);
and U1336 (N_1336,N_1240,N_1251);
or U1337 (N_1337,N_1224,N_1201);
nand U1338 (N_1338,N_1275,N_1245);
and U1339 (N_1339,N_1254,N_1231);
nor U1340 (N_1340,N_1268,N_1223);
nand U1341 (N_1341,N_1226,N_1297);
or U1342 (N_1342,N_1205,N_1271);
or U1343 (N_1343,N_1280,N_1278);
xnor U1344 (N_1344,N_1252,N_1247);
nor U1345 (N_1345,N_1225,N_1219);
and U1346 (N_1346,N_1227,N_1284);
or U1347 (N_1347,N_1255,N_1282);
nor U1348 (N_1348,N_1256,N_1216);
or U1349 (N_1349,N_1289,N_1277);
nor U1350 (N_1350,N_1239,N_1263);
nor U1351 (N_1351,N_1267,N_1243);
or U1352 (N_1352,N_1269,N_1256);
and U1353 (N_1353,N_1236,N_1251);
nor U1354 (N_1354,N_1240,N_1233);
nand U1355 (N_1355,N_1248,N_1269);
nand U1356 (N_1356,N_1299,N_1260);
or U1357 (N_1357,N_1234,N_1225);
nand U1358 (N_1358,N_1282,N_1253);
or U1359 (N_1359,N_1262,N_1286);
nor U1360 (N_1360,N_1239,N_1208);
nand U1361 (N_1361,N_1227,N_1285);
nor U1362 (N_1362,N_1283,N_1210);
nand U1363 (N_1363,N_1236,N_1204);
or U1364 (N_1364,N_1237,N_1233);
nor U1365 (N_1365,N_1242,N_1252);
or U1366 (N_1366,N_1236,N_1278);
nor U1367 (N_1367,N_1233,N_1298);
nand U1368 (N_1368,N_1288,N_1246);
nand U1369 (N_1369,N_1284,N_1205);
and U1370 (N_1370,N_1235,N_1248);
xnor U1371 (N_1371,N_1202,N_1284);
nor U1372 (N_1372,N_1200,N_1217);
nor U1373 (N_1373,N_1220,N_1299);
or U1374 (N_1374,N_1221,N_1275);
or U1375 (N_1375,N_1237,N_1272);
xnor U1376 (N_1376,N_1282,N_1265);
nor U1377 (N_1377,N_1216,N_1244);
or U1378 (N_1378,N_1227,N_1298);
or U1379 (N_1379,N_1288,N_1233);
xor U1380 (N_1380,N_1278,N_1210);
and U1381 (N_1381,N_1238,N_1256);
nor U1382 (N_1382,N_1218,N_1281);
or U1383 (N_1383,N_1224,N_1267);
nor U1384 (N_1384,N_1257,N_1204);
or U1385 (N_1385,N_1299,N_1269);
nor U1386 (N_1386,N_1226,N_1279);
and U1387 (N_1387,N_1215,N_1286);
nand U1388 (N_1388,N_1221,N_1278);
or U1389 (N_1389,N_1245,N_1203);
or U1390 (N_1390,N_1200,N_1213);
and U1391 (N_1391,N_1231,N_1245);
or U1392 (N_1392,N_1257,N_1230);
nor U1393 (N_1393,N_1268,N_1235);
or U1394 (N_1394,N_1276,N_1282);
and U1395 (N_1395,N_1243,N_1285);
and U1396 (N_1396,N_1259,N_1215);
or U1397 (N_1397,N_1264,N_1203);
and U1398 (N_1398,N_1294,N_1261);
xnor U1399 (N_1399,N_1255,N_1297);
nor U1400 (N_1400,N_1303,N_1305);
and U1401 (N_1401,N_1345,N_1340);
or U1402 (N_1402,N_1395,N_1320);
xor U1403 (N_1403,N_1306,N_1365);
or U1404 (N_1404,N_1338,N_1339);
and U1405 (N_1405,N_1335,N_1309);
and U1406 (N_1406,N_1385,N_1356);
or U1407 (N_1407,N_1396,N_1324);
xor U1408 (N_1408,N_1322,N_1318);
or U1409 (N_1409,N_1379,N_1382);
nor U1410 (N_1410,N_1376,N_1307);
nor U1411 (N_1411,N_1333,N_1310);
and U1412 (N_1412,N_1378,N_1397);
xnor U1413 (N_1413,N_1311,N_1360);
nor U1414 (N_1414,N_1358,N_1313);
xnor U1415 (N_1415,N_1330,N_1363);
nand U1416 (N_1416,N_1399,N_1304);
nor U1417 (N_1417,N_1380,N_1369);
and U1418 (N_1418,N_1326,N_1347);
and U1419 (N_1419,N_1386,N_1321);
nor U1420 (N_1420,N_1353,N_1364);
xor U1421 (N_1421,N_1349,N_1375);
nor U1422 (N_1422,N_1336,N_1348);
and U1423 (N_1423,N_1370,N_1312);
and U1424 (N_1424,N_1323,N_1381);
or U1425 (N_1425,N_1373,N_1372);
nand U1426 (N_1426,N_1317,N_1394);
nor U1427 (N_1427,N_1361,N_1398);
and U1428 (N_1428,N_1301,N_1355);
and U1429 (N_1429,N_1341,N_1362);
nor U1430 (N_1430,N_1390,N_1328);
and U1431 (N_1431,N_1319,N_1388);
and U1432 (N_1432,N_1314,N_1302);
and U1433 (N_1433,N_1392,N_1357);
nand U1434 (N_1434,N_1393,N_1366);
or U1435 (N_1435,N_1300,N_1354);
and U1436 (N_1436,N_1344,N_1337);
nand U1437 (N_1437,N_1377,N_1351);
or U1438 (N_1438,N_1383,N_1331);
xnor U1439 (N_1439,N_1391,N_1352);
or U1440 (N_1440,N_1316,N_1315);
nor U1441 (N_1441,N_1387,N_1325);
nor U1442 (N_1442,N_1329,N_1374);
or U1443 (N_1443,N_1342,N_1346);
and U1444 (N_1444,N_1367,N_1343);
or U1445 (N_1445,N_1334,N_1384);
nor U1446 (N_1446,N_1389,N_1371);
xor U1447 (N_1447,N_1359,N_1368);
or U1448 (N_1448,N_1350,N_1332);
or U1449 (N_1449,N_1308,N_1327);
nand U1450 (N_1450,N_1326,N_1316);
nor U1451 (N_1451,N_1342,N_1399);
nand U1452 (N_1452,N_1369,N_1316);
and U1453 (N_1453,N_1346,N_1367);
and U1454 (N_1454,N_1387,N_1301);
and U1455 (N_1455,N_1381,N_1383);
nor U1456 (N_1456,N_1312,N_1372);
nand U1457 (N_1457,N_1360,N_1316);
and U1458 (N_1458,N_1397,N_1337);
or U1459 (N_1459,N_1317,N_1302);
nand U1460 (N_1460,N_1327,N_1363);
and U1461 (N_1461,N_1325,N_1373);
and U1462 (N_1462,N_1328,N_1375);
and U1463 (N_1463,N_1367,N_1340);
nor U1464 (N_1464,N_1375,N_1335);
nor U1465 (N_1465,N_1363,N_1377);
nor U1466 (N_1466,N_1315,N_1387);
or U1467 (N_1467,N_1362,N_1305);
nand U1468 (N_1468,N_1387,N_1310);
xnor U1469 (N_1469,N_1303,N_1388);
nand U1470 (N_1470,N_1309,N_1332);
nor U1471 (N_1471,N_1334,N_1346);
or U1472 (N_1472,N_1348,N_1358);
nand U1473 (N_1473,N_1379,N_1363);
nor U1474 (N_1474,N_1378,N_1382);
or U1475 (N_1475,N_1343,N_1306);
nand U1476 (N_1476,N_1371,N_1308);
and U1477 (N_1477,N_1373,N_1385);
nor U1478 (N_1478,N_1308,N_1391);
and U1479 (N_1479,N_1340,N_1336);
nor U1480 (N_1480,N_1395,N_1357);
nand U1481 (N_1481,N_1353,N_1312);
and U1482 (N_1482,N_1392,N_1371);
nand U1483 (N_1483,N_1320,N_1304);
nor U1484 (N_1484,N_1347,N_1316);
nand U1485 (N_1485,N_1314,N_1386);
nand U1486 (N_1486,N_1349,N_1359);
or U1487 (N_1487,N_1365,N_1385);
and U1488 (N_1488,N_1392,N_1368);
nand U1489 (N_1489,N_1317,N_1320);
xor U1490 (N_1490,N_1318,N_1399);
xor U1491 (N_1491,N_1387,N_1360);
or U1492 (N_1492,N_1317,N_1342);
or U1493 (N_1493,N_1328,N_1371);
or U1494 (N_1494,N_1361,N_1346);
or U1495 (N_1495,N_1356,N_1302);
and U1496 (N_1496,N_1341,N_1330);
xnor U1497 (N_1497,N_1334,N_1375);
xor U1498 (N_1498,N_1339,N_1332);
and U1499 (N_1499,N_1324,N_1356);
nor U1500 (N_1500,N_1445,N_1472);
xor U1501 (N_1501,N_1442,N_1454);
nand U1502 (N_1502,N_1433,N_1466);
nor U1503 (N_1503,N_1400,N_1447);
and U1504 (N_1504,N_1456,N_1494);
nor U1505 (N_1505,N_1499,N_1403);
nand U1506 (N_1506,N_1423,N_1458);
nand U1507 (N_1507,N_1414,N_1431);
or U1508 (N_1508,N_1459,N_1469);
or U1509 (N_1509,N_1452,N_1430);
nor U1510 (N_1510,N_1405,N_1420);
and U1511 (N_1511,N_1421,N_1488);
and U1512 (N_1512,N_1481,N_1475);
nor U1513 (N_1513,N_1467,N_1464);
nand U1514 (N_1514,N_1453,N_1461);
nor U1515 (N_1515,N_1498,N_1478);
or U1516 (N_1516,N_1432,N_1471);
nor U1517 (N_1517,N_1495,N_1409);
and U1518 (N_1518,N_1415,N_1428);
or U1519 (N_1519,N_1476,N_1455);
and U1520 (N_1520,N_1473,N_1407);
and U1521 (N_1521,N_1439,N_1406);
nand U1522 (N_1522,N_1402,N_1465);
or U1523 (N_1523,N_1484,N_1427);
nor U1524 (N_1524,N_1480,N_1411);
nor U1525 (N_1525,N_1436,N_1487);
and U1526 (N_1526,N_1491,N_1468);
or U1527 (N_1527,N_1470,N_1441);
nor U1528 (N_1528,N_1404,N_1422);
nand U1529 (N_1529,N_1443,N_1460);
nor U1530 (N_1530,N_1492,N_1457);
nand U1531 (N_1531,N_1462,N_1418);
or U1532 (N_1532,N_1429,N_1419);
or U1533 (N_1533,N_1477,N_1449);
or U1534 (N_1534,N_1485,N_1438);
nor U1535 (N_1535,N_1401,N_1451);
or U1536 (N_1536,N_1408,N_1493);
or U1537 (N_1537,N_1448,N_1463);
xor U1538 (N_1538,N_1489,N_1416);
and U1539 (N_1539,N_1486,N_1450);
nand U1540 (N_1540,N_1435,N_1434);
nand U1541 (N_1541,N_1446,N_1417);
nand U1542 (N_1542,N_1425,N_1424);
nor U1543 (N_1543,N_1496,N_1426);
xnor U1544 (N_1544,N_1482,N_1474);
or U1545 (N_1545,N_1483,N_1490);
nand U1546 (N_1546,N_1440,N_1497);
and U1547 (N_1547,N_1444,N_1413);
or U1548 (N_1548,N_1412,N_1410);
nor U1549 (N_1549,N_1479,N_1437);
and U1550 (N_1550,N_1476,N_1440);
and U1551 (N_1551,N_1489,N_1475);
or U1552 (N_1552,N_1416,N_1490);
or U1553 (N_1553,N_1400,N_1461);
or U1554 (N_1554,N_1419,N_1422);
nand U1555 (N_1555,N_1410,N_1435);
or U1556 (N_1556,N_1470,N_1435);
nand U1557 (N_1557,N_1460,N_1411);
and U1558 (N_1558,N_1444,N_1423);
xnor U1559 (N_1559,N_1491,N_1423);
nand U1560 (N_1560,N_1478,N_1404);
or U1561 (N_1561,N_1432,N_1451);
nand U1562 (N_1562,N_1495,N_1403);
and U1563 (N_1563,N_1479,N_1450);
nand U1564 (N_1564,N_1440,N_1486);
and U1565 (N_1565,N_1430,N_1418);
or U1566 (N_1566,N_1413,N_1455);
nand U1567 (N_1567,N_1426,N_1413);
and U1568 (N_1568,N_1492,N_1498);
or U1569 (N_1569,N_1408,N_1449);
xor U1570 (N_1570,N_1431,N_1426);
nor U1571 (N_1571,N_1461,N_1407);
and U1572 (N_1572,N_1478,N_1431);
or U1573 (N_1573,N_1453,N_1415);
nor U1574 (N_1574,N_1401,N_1404);
and U1575 (N_1575,N_1450,N_1485);
nand U1576 (N_1576,N_1446,N_1473);
nor U1577 (N_1577,N_1419,N_1490);
and U1578 (N_1578,N_1417,N_1494);
and U1579 (N_1579,N_1457,N_1454);
nand U1580 (N_1580,N_1413,N_1433);
xor U1581 (N_1581,N_1404,N_1442);
nand U1582 (N_1582,N_1434,N_1462);
nor U1583 (N_1583,N_1498,N_1411);
and U1584 (N_1584,N_1462,N_1455);
or U1585 (N_1585,N_1482,N_1468);
nand U1586 (N_1586,N_1404,N_1403);
nand U1587 (N_1587,N_1404,N_1426);
and U1588 (N_1588,N_1457,N_1436);
nor U1589 (N_1589,N_1432,N_1427);
or U1590 (N_1590,N_1427,N_1438);
nor U1591 (N_1591,N_1433,N_1476);
nor U1592 (N_1592,N_1412,N_1411);
and U1593 (N_1593,N_1410,N_1466);
nand U1594 (N_1594,N_1409,N_1491);
nand U1595 (N_1595,N_1482,N_1436);
and U1596 (N_1596,N_1440,N_1451);
xor U1597 (N_1597,N_1436,N_1470);
or U1598 (N_1598,N_1460,N_1495);
nor U1599 (N_1599,N_1449,N_1446);
and U1600 (N_1600,N_1522,N_1511);
nor U1601 (N_1601,N_1583,N_1517);
xnor U1602 (N_1602,N_1528,N_1533);
or U1603 (N_1603,N_1568,N_1516);
xnor U1604 (N_1604,N_1526,N_1508);
nand U1605 (N_1605,N_1546,N_1536);
and U1606 (N_1606,N_1589,N_1585);
nand U1607 (N_1607,N_1509,N_1532);
nor U1608 (N_1608,N_1544,N_1574);
or U1609 (N_1609,N_1524,N_1579);
nand U1610 (N_1610,N_1538,N_1539);
xor U1611 (N_1611,N_1588,N_1519);
nor U1612 (N_1612,N_1529,N_1534);
or U1613 (N_1613,N_1512,N_1561);
nor U1614 (N_1614,N_1558,N_1557);
nor U1615 (N_1615,N_1530,N_1543);
nand U1616 (N_1616,N_1555,N_1513);
nor U1617 (N_1617,N_1523,N_1590);
nand U1618 (N_1618,N_1518,N_1571);
or U1619 (N_1619,N_1586,N_1535);
nand U1620 (N_1620,N_1515,N_1505);
xor U1621 (N_1621,N_1506,N_1559);
nand U1622 (N_1622,N_1567,N_1576);
and U1623 (N_1623,N_1594,N_1537);
and U1624 (N_1624,N_1562,N_1560);
nand U1625 (N_1625,N_1570,N_1502);
nand U1626 (N_1626,N_1595,N_1596);
nand U1627 (N_1627,N_1507,N_1552);
and U1628 (N_1628,N_1593,N_1565);
nor U1629 (N_1629,N_1521,N_1587);
and U1630 (N_1630,N_1592,N_1582);
and U1631 (N_1631,N_1551,N_1577);
nand U1632 (N_1632,N_1564,N_1563);
xnor U1633 (N_1633,N_1547,N_1578);
and U1634 (N_1634,N_1599,N_1520);
or U1635 (N_1635,N_1591,N_1554);
nand U1636 (N_1636,N_1572,N_1514);
and U1637 (N_1637,N_1504,N_1549);
and U1638 (N_1638,N_1525,N_1501);
and U1639 (N_1639,N_1597,N_1598);
or U1640 (N_1640,N_1541,N_1542);
nand U1641 (N_1641,N_1581,N_1556);
nand U1642 (N_1642,N_1573,N_1566);
nand U1643 (N_1643,N_1527,N_1531);
nor U1644 (N_1644,N_1510,N_1580);
xnor U1645 (N_1645,N_1503,N_1550);
nand U1646 (N_1646,N_1553,N_1569);
nand U1647 (N_1647,N_1540,N_1575);
nand U1648 (N_1648,N_1545,N_1584);
and U1649 (N_1649,N_1500,N_1548);
nand U1650 (N_1650,N_1509,N_1573);
or U1651 (N_1651,N_1573,N_1594);
nor U1652 (N_1652,N_1588,N_1554);
nand U1653 (N_1653,N_1506,N_1540);
nand U1654 (N_1654,N_1502,N_1508);
nand U1655 (N_1655,N_1573,N_1532);
nor U1656 (N_1656,N_1589,N_1583);
xnor U1657 (N_1657,N_1540,N_1532);
and U1658 (N_1658,N_1531,N_1514);
nor U1659 (N_1659,N_1516,N_1505);
or U1660 (N_1660,N_1530,N_1539);
xnor U1661 (N_1661,N_1558,N_1522);
xor U1662 (N_1662,N_1569,N_1523);
or U1663 (N_1663,N_1572,N_1535);
nand U1664 (N_1664,N_1589,N_1588);
nand U1665 (N_1665,N_1539,N_1529);
or U1666 (N_1666,N_1538,N_1549);
nor U1667 (N_1667,N_1540,N_1514);
nand U1668 (N_1668,N_1569,N_1520);
xnor U1669 (N_1669,N_1514,N_1544);
nor U1670 (N_1670,N_1559,N_1574);
nor U1671 (N_1671,N_1554,N_1515);
or U1672 (N_1672,N_1535,N_1580);
nor U1673 (N_1673,N_1555,N_1520);
xor U1674 (N_1674,N_1555,N_1536);
nand U1675 (N_1675,N_1516,N_1515);
nor U1676 (N_1676,N_1510,N_1574);
xor U1677 (N_1677,N_1536,N_1598);
or U1678 (N_1678,N_1573,N_1503);
or U1679 (N_1679,N_1554,N_1548);
nand U1680 (N_1680,N_1533,N_1523);
nand U1681 (N_1681,N_1559,N_1564);
or U1682 (N_1682,N_1526,N_1505);
nor U1683 (N_1683,N_1531,N_1583);
nand U1684 (N_1684,N_1507,N_1575);
nor U1685 (N_1685,N_1565,N_1552);
nand U1686 (N_1686,N_1598,N_1504);
and U1687 (N_1687,N_1596,N_1571);
or U1688 (N_1688,N_1525,N_1527);
nor U1689 (N_1689,N_1514,N_1529);
and U1690 (N_1690,N_1543,N_1500);
and U1691 (N_1691,N_1508,N_1566);
nand U1692 (N_1692,N_1543,N_1580);
and U1693 (N_1693,N_1504,N_1559);
nor U1694 (N_1694,N_1534,N_1547);
nand U1695 (N_1695,N_1589,N_1503);
and U1696 (N_1696,N_1549,N_1546);
nand U1697 (N_1697,N_1584,N_1511);
nor U1698 (N_1698,N_1574,N_1598);
and U1699 (N_1699,N_1534,N_1526);
nor U1700 (N_1700,N_1685,N_1613);
nor U1701 (N_1701,N_1621,N_1698);
nor U1702 (N_1702,N_1649,N_1681);
nand U1703 (N_1703,N_1630,N_1673);
and U1704 (N_1704,N_1665,N_1674);
nand U1705 (N_1705,N_1610,N_1671);
nand U1706 (N_1706,N_1695,N_1643);
nand U1707 (N_1707,N_1645,N_1684);
xnor U1708 (N_1708,N_1687,N_1658);
xor U1709 (N_1709,N_1686,N_1691);
and U1710 (N_1710,N_1656,N_1666);
nor U1711 (N_1711,N_1668,N_1638);
nand U1712 (N_1712,N_1600,N_1694);
nor U1713 (N_1713,N_1629,N_1678);
nand U1714 (N_1714,N_1647,N_1611);
nor U1715 (N_1715,N_1637,N_1651);
and U1716 (N_1716,N_1607,N_1601);
and U1717 (N_1717,N_1667,N_1628);
nor U1718 (N_1718,N_1605,N_1603);
nor U1719 (N_1719,N_1644,N_1642);
nor U1720 (N_1720,N_1670,N_1617);
or U1721 (N_1721,N_1615,N_1689);
or U1722 (N_1722,N_1683,N_1639);
nand U1723 (N_1723,N_1672,N_1640);
nand U1724 (N_1724,N_1624,N_1663);
and U1725 (N_1725,N_1606,N_1682);
or U1726 (N_1726,N_1692,N_1627);
or U1727 (N_1727,N_1619,N_1677);
nand U1728 (N_1728,N_1661,N_1676);
and U1729 (N_1729,N_1608,N_1679);
or U1730 (N_1730,N_1657,N_1622);
or U1731 (N_1731,N_1626,N_1618);
nor U1732 (N_1732,N_1669,N_1646);
or U1733 (N_1733,N_1634,N_1648);
or U1734 (N_1734,N_1697,N_1633);
xor U1735 (N_1735,N_1660,N_1655);
or U1736 (N_1736,N_1632,N_1620);
nand U1737 (N_1737,N_1641,N_1635);
nand U1738 (N_1738,N_1631,N_1699);
or U1739 (N_1739,N_1664,N_1659);
and U1740 (N_1740,N_1604,N_1636);
nand U1741 (N_1741,N_1625,N_1609);
or U1742 (N_1742,N_1650,N_1616);
or U1743 (N_1743,N_1696,N_1623);
or U1744 (N_1744,N_1693,N_1675);
nor U1745 (N_1745,N_1654,N_1602);
nor U1746 (N_1746,N_1652,N_1614);
or U1747 (N_1747,N_1688,N_1680);
or U1748 (N_1748,N_1690,N_1653);
nand U1749 (N_1749,N_1662,N_1612);
nand U1750 (N_1750,N_1687,N_1604);
and U1751 (N_1751,N_1626,N_1657);
nand U1752 (N_1752,N_1605,N_1628);
nand U1753 (N_1753,N_1615,N_1681);
nor U1754 (N_1754,N_1621,N_1636);
or U1755 (N_1755,N_1612,N_1693);
nand U1756 (N_1756,N_1609,N_1608);
nor U1757 (N_1757,N_1671,N_1602);
and U1758 (N_1758,N_1616,N_1692);
or U1759 (N_1759,N_1622,N_1692);
or U1760 (N_1760,N_1663,N_1661);
nor U1761 (N_1761,N_1694,N_1679);
nor U1762 (N_1762,N_1612,N_1641);
nand U1763 (N_1763,N_1643,N_1662);
nor U1764 (N_1764,N_1652,N_1648);
nor U1765 (N_1765,N_1600,N_1645);
nor U1766 (N_1766,N_1694,N_1620);
nand U1767 (N_1767,N_1691,N_1632);
nor U1768 (N_1768,N_1667,N_1648);
nand U1769 (N_1769,N_1617,N_1627);
or U1770 (N_1770,N_1662,N_1608);
or U1771 (N_1771,N_1661,N_1623);
and U1772 (N_1772,N_1611,N_1683);
nor U1773 (N_1773,N_1622,N_1689);
and U1774 (N_1774,N_1696,N_1612);
nor U1775 (N_1775,N_1615,N_1619);
xor U1776 (N_1776,N_1675,N_1618);
nor U1777 (N_1777,N_1651,N_1662);
and U1778 (N_1778,N_1682,N_1632);
nor U1779 (N_1779,N_1601,N_1684);
nor U1780 (N_1780,N_1614,N_1643);
nand U1781 (N_1781,N_1641,N_1658);
and U1782 (N_1782,N_1675,N_1676);
nand U1783 (N_1783,N_1668,N_1680);
nor U1784 (N_1784,N_1618,N_1695);
nand U1785 (N_1785,N_1690,N_1615);
nor U1786 (N_1786,N_1629,N_1660);
nor U1787 (N_1787,N_1698,N_1617);
nor U1788 (N_1788,N_1634,N_1652);
or U1789 (N_1789,N_1610,N_1655);
and U1790 (N_1790,N_1686,N_1653);
or U1791 (N_1791,N_1622,N_1635);
and U1792 (N_1792,N_1649,N_1642);
nand U1793 (N_1793,N_1638,N_1699);
and U1794 (N_1794,N_1656,N_1694);
nor U1795 (N_1795,N_1674,N_1697);
nor U1796 (N_1796,N_1628,N_1646);
nor U1797 (N_1797,N_1662,N_1648);
and U1798 (N_1798,N_1690,N_1699);
or U1799 (N_1799,N_1657,N_1691);
or U1800 (N_1800,N_1747,N_1741);
and U1801 (N_1801,N_1750,N_1787);
or U1802 (N_1802,N_1772,N_1767);
or U1803 (N_1803,N_1717,N_1716);
and U1804 (N_1804,N_1773,N_1784);
nand U1805 (N_1805,N_1779,N_1730);
or U1806 (N_1806,N_1749,N_1791);
nand U1807 (N_1807,N_1701,N_1780);
nor U1808 (N_1808,N_1756,N_1706);
nor U1809 (N_1809,N_1704,N_1740);
nor U1810 (N_1810,N_1721,N_1743);
nor U1811 (N_1811,N_1789,N_1792);
nand U1812 (N_1812,N_1724,N_1778);
nand U1813 (N_1813,N_1713,N_1742);
or U1814 (N_1814,N_1769,N_1723);
nand U1815 (N_1815,N_1746,N_1783);
nand U1816 (N_1816,N_1763,N_1735);
nand U1817 (N_1817,N_1745,N_1702);
xor U1818 (N_1818,N_1736,N_1764);
xor U1819 (N_1819,N_1754,N_1733);
and U1820 (N_1820,N_1744,N_1725);
or U1821 (N_1821,N_1705,N_1719);
and U1822 (N_1822,N_1765,N_1775);
xnor U1823 (N_1823,N_1727,N_1795);
nand U1824 (N_1824,N_1752,N_1739);
nor U1825 (N_1825,N_1766,N_1734);
nor U1826 (N_1826,N_1759,N_1790);
or U1827 (N_1827,N_1753,N_1796);
xor U1828 (N_1828,N_1711,N_1710);
nand U1829 (N_1829,N_1720,N_1728);
nand U1830 (N_1830,N_1709,N_1722);
nor U1831 (N_1831,N_1751,N_1760);
nor U1832 (N_1832,N_1755,N_1726);
nand U1833 (N_1833,N_1799,N_1707);
nor U1834 (N_1834,N_1715,N_1708);
nand U1835 (N_1835,N_1718,N_1798);
and U1836 (N_1836,N_1700,N_1737);
nor U1837 (N_1837,N_1774,N_1794);
or U1838 (N_1838,N_1786,N_1703);
and U1839 (N_1839,N_1757,N_1785);
and U1840 (N_1840,N_1781,N_1793);
and U1841 (N_1841,N_1776,N_1748);
and U1842 (N_1842,N_1762,N_1714);
xnor U1843 (N_1843,N_1777,N_1782);
and U1844 (N_1844,N_1729,N_1761);
nor U1845 (N_1845,N_1797,N_1758);
and U1846 (N_1846,N_1768,N_1731);
or U1847 (N_1847,N_1788,N_1770);
or U1848 (N_1848,N_1712,N_1738);
nor U1849 (N_1849,N_1771,N_1732);
nor U1850 (N_1850,N_1720,N_1795);
or U1851 (N_1851,N_1728,N_1788);
nand U1852 (N_1852,N_1700,N_1708);
xor U1853 (N_1853,N_1759,N_1776);
nand U1854 (N_1854,N_1752,N_1717);
nand U1855 (N_1855,N_1710,N_1755);
and U1856 (N_1856,N_1725,N_1783);
nand U1857 (N_1857,N_1752,N_1713);
nor U1858 (N_1858,N_1728,N_1738);
and U1859 (N_1859,N_1769,N_1726);
and U1860 (N_1860,N_1726,N_1735);
and U1861 (N_1861,N_1779,N_1721);
nor U1862 (N_1862,N_1708,N_1725);
xor U1863 (N_1863,N_1790,N_1770);
and U1864 (N_1864,N_1755,N_1761);
nand U1865 (N_1865,N_1747,N_1779);
xnor U1866 (N_1866,N_1772,N_1797);
nand U1867 (N_1867,N_1719,N_1798);
or U1868 (N_1868,N_1735,N_1715);
and U1869 (N_1869,N_1718,N_1727);
or U1870 (N_1870,N_1774,N_1736);
nand U1871 (N_1871,N_1786,N_1741);
nand U1872 (N_1872,N_1779,N_1725);
nand U1873 (N_1873,N_1759,N_1707);
or U1874 (N_1874,N_1710,N_1701);
nand U1875 (N_1875,N_1730,N_1758);
and U1876 (N_1876,N_1782,N_1748);
or U1877 (N_1877,N_1797,N_1749);
nand U1878 (N_1878,N_1736,N_1702);
and U1879 (N_1879,N_1772,N_1721);
and U1880 (N_1880,N_1762,N_1742);
nor U1881 (N_1881,N_1792,N_1740);
or U1882 (N_1882,N_1714,N_1702);
nand U1883 (N_1883,N_1751,N_1701);
nor U1884 (N_1884,N_1734,N_1788);
and U1885 (N_1885,N_1735,N_1729);
nor U1886 (N_1886,N_1721,N_1791);
or U1887 (N_1887,N_1762,N_1759);
nor U1888 (N_1888,N_1785,N_1702);
or U1889 (N_1889,N_1778,N_1734);
or U1890 (N_1890,N_1771,N_1708);
xor U1891 (N_1891,N_1770,N_1727);
nor U1892 (N_1892,N_1710,N_1796);
or U1893 (N_1893,N_1759,N_1721);
nor U1894 (N_1894,N_1701,N_1772);
and U1895 (N_1895,N_1710,N_1779);
and U1896 (N_1896,N_1744,N_1787);
or U1897 (N_1897,N_1793,N_1719);
nor U1898 (N_1898,N_1787,N_1742);
or U1899 (N_1899,N_1789,N_1729);
and U1900 (N_1900,N_1864,N_1891);
and U1901 (N_1901,N_1841,N_1815);
xor U1902 (N_1902,N_1896,N_1825);
and U1903 (N_1903,N_1876,N_1883);
and U1904 (N_1904,N_1853,N_1888);
or U1905 (N_1905,N_1873,N_1817);
and U1906 (N_1906,N_1868,N_1816);
nand U1907 (N_1907,N_1863,N_1851);
nor U1908 (N_1908,N_1848,N_1861);
nor U1909 (N_1909,N_1886,N_1893);
and U1910 (N_1910,N_1824,N_1871);
or U1911 (N_1911,N_1807,N_1874);
and U1912 (N_1912,N_1801,N_1885);
and U1913 (N_1913,N_1829,N_1828);
nor U1914 (N_1914,N_1823,N_1830);
nor U1915 (N_1915,N_1882,N_1890);
and U1916 (N_1916,N_1831,N_1838);
xnor U1917 (N_1917,N_1810,N_1865);
nor U1918 (N_1918,N_1809,N_1870);
nor U1919 (N_1919,N_1854,N_1814);
nand U1920 (N_1920,N_1820,N_1872);
nor U1921 (N_1921,N_1899,N_1835);
xor U1922 (N_1922,N_1827,N_1840);
nand U1923 (N_1923,N_1826,N_1812);
xor U1924 (N_1924,N_1808,N_1858);
nand U1925 (N_1925,N_1822,N_1866);
xor U1926 (N_1926,N_1894,N_1862);
nand U1927 (N_1927,N_1877,N_1869);
nor U1928 (N_1928,N_1802,N_1897);
and U1929 (N_1929,N_1843,N_1800);
and U1930 (N_1930,N_1833,N_1879);
nor U1931 (N_1931,N_1860,N_1855);
and U1932 (N_1932,N_1819,N_1880);
and U1933 (N_1933,N_1806,N_1867);
xor U1934 (N_1934,N_1805,N_1878);
nand U1935 (N_1935,N_1836,N_1832);
or U1936 (N_1936,N_1846,N_1887);
and U1937 (N_1937,N_1884,N_1839);
nor U1938 (N_1938,N_1842,N_1892);
nor U1939 (N_1939,N_1845,N_1821);
nand U1940 (N_1940,N_1813,N_1811);
nor U1941 (N_1941,N_1847,N_1837);
and U1942 (N_1942,N_1818,N_1895);
and U1943 (N_1943,N_1881,N_1889);
or U1944 (N_1944,N_1844,N_1898);
nand U1945 (N_1945,N_1834,N_1850);
nor U1946 (N_1946,N_1859,N_1804);
nand U1947 (N_1947,N_1849,N_1857);
or U1948 (N_1948,N_1875,N_1856);
nor U1949 (N_1949,N_1852,N_1803);
nor U1950 (N_1950,N_1816,N_1867);
nor U1951 (N_1951,N_1892,N_1836);
nand U1952 (N_1952,N_1813,N_1805);
nand U1953 (N_1953,N_1827,N_1810);
or U1954 (N_1954,N_1872,N_1895);
nor U1955 (N_1955,N_1844,N_1896);
nand U1956 (N_1956,N_1856,N_1872);
or U1957 (N_1957,N_1878,N_1825);
nand U1958 (N_1958,N_1884,N_1877);
nand U1959 (N_1959,N_1866,N_1869);
xnor U1960 (N_1960,N_1838,N_1885);
nor U1961 (N_1961,N_1803,N_1882);
or U1962 (N_1962,N_1812,N_1811);
or U1963 (N_1963,N_1854,N_1855);
and U1964 (N_1964,N_1845,N_1875);
and U1965 (N_1965,N_1868,N_1885);
and U1966 (N_1966,N_1806,N_1815);
nor U1967 (N_1967,N_1885,N_1822);
or U1968 (N_1968,N_1894,N_1806);
or U1969 (N_1969,N_1823,N_1875);
xnor U1970 (N_1970,N_1893,N_1871);
or U1971 (N_1971,N_1885,N_1882);
nor U1972 (N_1972,N_1890,N_1822);
and U1973 (N_1973,N_1885,N_1876);
or U1974 (N_1974,N_1896,N_1879);
nand U1975 (N_1975,N_1884,N_1831);
or U1976 (N_1976,N_1814,N_1874);
nor U1977 (N_1977,N_1808,N_1832);
and U1978 (N_1978,N_1865,N_1829);
nor U1979 (N_1979,N_1874,N_1884);
and U1980 (N_1980,N_1823,N_1857);
nand U1981 (N_1981,N_1891,N_1815);
and U1982 (N_1982,N_1878,N_1873);
nand U1983 (N_1983,N_1886,N_1891);
nor U1984 (N_1984,N_1863,N_1825);
and U1985 (N_1985,N_1814,N_1895);
and U1986 (N_1986,N_1815,N_1865);
nor U1987 (N_1987,N_1835,N_1831);
nor U1988 (N_1988,N_1886,N_1816);
or U1989 (N_1989,N_1860,N_1865);
xnor U1990 (N_1990,N_1851,N_1839);
nand U1991 (N_1991,N_1888,N_1847);
and U1992 (N_1992,N_1882,N_1872);
and U1993 (N_1993,N_1864,N_1882);
and U1994 (N_1994,N_1840,N_1821);
xnor U1995 (N_1995,N_1872,N_1809);
or U1996 (N_1996,N_1836,N_1809);
and U1997 (N_1997,N_1823,N_1888);
or U1998 (N_1998,N_1874,N_1817);
nor U1999 (N_1999,N_1841,N_1874);
nor U2000 (N_2000,N_1985,N_1909);
nand U2001 (N_2001,N_1927,N_1983);
nand U2002 (N_2002,N_1905,N_1931);
nor U2003 (N_2003,N_1957,N_1944);
or U2004 (N_2004,N_1951,N_1968);
and U2005 (N_2005,N_1966,N_1961);
or U2006 (N_2006,N_1936,N_1942);
nand U2007 (N_2007,N_1929,N_1992);
xor U2008 (N_2008,N_1945,N_1902);
nand U2009 (N_2009,N_1903,N_1984);
nand U2010 (N_2010,N_1915,N_1962);
nand U2011 (N_2011,N_1978,N_1963);
nor U2012 (N_2012,N_1959,N_1946);
nor U2013 (N_2013,N_1965,N_1986);
nor U2014 (N_2014,N_1921,N_1954);
or U2015 (N_2015,N_1914,N_1926);
nand U2016 (N_2016,N_1906,N_1976);
nor U2017 (N_2017,N_1960,N_1923);
or U2018 (N_2018,N_1933,N_1989);
and U2019 (N_2019,N_1930,N_1973);
and U2020 (N_2020,N_1991,N_1917);
or U2021 (N_2021,N_1972,N_1990);
nand U2022 (N_2022,N_1941,N_1964);
nor U2023 (N_2023,N_1928,N_1943);
nand U2024 (N_2024,N_1974,N_1908);
and U2025 (N_2025,N_1918,N_1956);
and U2026 (N_2026,N_1994,N_1900);
nor U2027 (N_2027,N_1958,N_1949);
nand U2028 (N_2028,N_1910,N_1907);
nor U2029 (N_2029,N_1969,N_1981);
and U2030 (N_2030,N_1938,N_1916);
and U2031 (N_2031,N_1996,N_1947);
and U2032 (N_2032,N_1901,N_1987);
and U2033 (N_2033,N_1979,N_1932);
or U2034 (N_2034,N_1919,N_1924);
nor U2035 (N_2035,N_1935,N_1970);
nor U2036 (N_2036,N_1940,N_1995);
nor U2037 (N_2037,N_1937,N_1939);
and U2038 (N_2038,N_1955,N_1971);
xor U2039 (N_2039,N_1982,N_1950);
nor U2040 (N_2040,N_1975,N_1922);
nand U2041 (N_2041,N_1913,N_1952);
nand U2042 (N_2042,N_1920,N_1993);
and U2043 (N_2043,N_1999,N_1977);
xor U2044 (N_2044,N_1948,N_1934);
nand U2045 (N_2045,N_1911,N_1980);
xnor U2046 (N_2046,N_1967,N_1988);
nor U2047 (N_2047,N_1912,N_1925);
and U2048 (N_2048,N_1997,N_1998);
or U2049 (N_2049,N_1904,N_1953);
and U2050 (N_2050,N_1928,N_1965);
or U2051 (N_2051,N_1911,N_1907);
and U2052 (N_2052,N_1943,N_1929);
nand U2053 (N_2053,N_1933,N_1994);
or U2054 (N_2054,N_1918,N_1993);
and U2055 (N_2055,N_1914,N_1935);
nand U2056 (N_2056,N_1989,N_1920);
or U2057 (N_2057,N_1992,N_1921);
nor U2058 (N_2058,N_1939,N_1997);
and U2059 (N_2059,N_1979,N_1957);
or U2060 (N_2060,N_1968,N_1956);
nand U2061 (N_2061,N_1999,N_1974);
or U2062 (N_2062,N_1934,N_1938);
and U2063 (N_2063,N_1977,N_1946);
or U2064 (N_2064,N_1967,N_1924);
or U2065 (N_2065,N_1996,N_1927);
or U2066 (N_2066,N_1900,N_1923);
nand U2067 (N_2067,N_1928,N_1932);
nand U2068 (N_2068,N_1962,N_1901);
nand U2069 (N_2069,N_1909,N_1967);
or U2070 (N_2070,N_1922,N_1956);
or U2071 (N_2071,N_1929,N_1981);
and U2072 (N_2072,N_1978,N_1942);
or U2073 (N_2073,N_1922,N_1977);
nor U2074 (N_2074,N_1977,N_1931);
or U2075 (N_2075,N_1913,N_1941);
nor U2076 (N_2076,N_1924,N_1911);
nor U2077 (N_2077,N_1925,N_1911);
and U2078 (N_2078,N_1926,N_1972);
xor U2079 (N_2079,N_1956,N_1966);
and U2080 (N_2080,N_1908,N_1999);
and U2081 (N_2081,N_1942,N_1996);
or U2082 (N_2082,N_1917,N_1985);
nor U2083 (N_2083,N_1993,N_1934);
nor U2084 (N_2084,N_1959,N_1932);
and U2085 (N_2085,N_1913,N_1962);
nand U2086 (N_2086,N_1920,N_1928);
nor U2087 (N_2087,N_1932,N_1939);
or U2088 (N_2088,N_1923,N_1998);
nor U2089 (N_2089,N_1907,N_1992);
nand U2090 (N_2090,N_1998,N_1965);
nand U2091 (N_2091,N_1913,N_1944);
nor U2092 (N_2092,N_1997,N_1993);
or U2093 (N_2093,N_1957,N_1946);
nor U2094 (N_2094,N_1942,N_1955);
nor U2095 (N_2095,N_1955,N_1973);
nor U2096 (N_2096,N_1931,N_1993);
or U2097 (N_2097,N_1987,N_1912);
and U2098 (N_2098,N_1918,N_1922);
or U2099 (N_2099,N_1995,N_1921);
xnor U2100 (N_2100,N_2026,N_2073);
and U2101 (N_2101,N_2066,N_2083);
nand U2102 (N_2102,N_2002,N_2050);
or U2103 (N_2103,N_2053,N_2078);
nand U2104 (N_2104,N_2087,N_2051);
nand U2105 (N_2105,N_2059,N_2012);
xnor U2106 (N_2106,N_2027,N_2034);
nor U2107 (N_2107,N_2075,N_2038);
nor U2108 (N_2108,N_2028,N_2046);
nor U2109 (N_2109,N_2084,N_2030);
nand U2110 (N_2110,N_2019,N_2041);
and U2111 (N_2111,N_2022,N_2095);
or U2112 (N_2112,N_2011,N_2061);
xnor U2113 (N_2113,N_2070,N_2089);
and U2114 (N_2114,N_2094,N_2099);
xnor U2115 (N_2115,N_2097,N_2093);
nand U2116 (N_2116,N_2092,N_2009);
and U2117 (N_2117,N_2015,N_2003);
xor U2118 (N_2118,N_2045,N_2031);
or U2119 (N_2119,N_2001,N_2074);
nand U2120 (N_2120,N_2090,N_2021);
nor U2121 (N_2121,N_2004,N_2007);
and U2122 (N_2122,N_2048,N_2005);
or U2123 (N_2123,N_2056,N_2096);
and U2124 (N_2124,N_2077,N_2072);
nor U2125 (N_2125,N_2008,N_2064);
nand U2126 (N_2126,N_2037,N_2071);
xor U2127 (N_2127,N_2054,N_2040);
nand U2128 (N_2128,N_2055,N_2020);
and U2129 (N_2129,N_2068,N_2085);
xnor U2130 (N_2130,N_2088,N_2010);
or U2131 (N_2131,N_2076,N_2082);
xnor U2132 (N_2132,N_2063,N_2052);
nor U2133 (N_2133,N_2067,N_2032);
and U2134 (N_2134,N_2025,N_2043);
nand U2135 (N_2135,N_2016,N_2014);
or U2136 (N_2136,N_2017,N_2086);
or U2137 (N_2137,N_2080,N_2091);
xnor U2138 (N_2138,N_2039,N_2018);
and U2139 (N_2139,N_2029,N_2098);
nand U2140 (N_2140,N_2065,N_2081);
nand U2141 (N_2141,N_2013,N_2079);
and U2142 (N_2142,N_2033,N_2024);
nor U2143 (N_2143,N_2006,N_2044);
nor U2144 (N_2144,N_2000,N_2023);
nand U2145 (N_2145,N_2042,N_2047);
and U2146 (N_2146,N_2035,N_2058);
nand U2147 (N_2147,N_2049,N_2069);
or U2148 (N_2148,N_2036,N_2060);
nand U2149 (N_2149,N_2057,N_2062);
or U2150 (N_2150,N_2057,N_2000);
nor U2151 (N_2151,N_2092,N_2098);
and U2152 (N_2152,N_2082,N_2070);
or U2153 (N_2153,N_2033,N_2099);
nor U2154 (N_2154,N_2091,N_2025);
or U2155 (N_2155,N_2038,N_2047);
or U2156 (N_2156,N_2067,N_2058);
and U2157 (N_2157,N_2021,N_2078);
xnor U2158 (N_2158,N_2094,N_2011);
or U2159 (N_2159,N_2061,N_2067);
and U2160 (N_2160,N_2023,N_2001);
nand U2161 (N_2161,N_2050,N_2027);
and U2162 (N_2162,N_2011,N_2023);
and U2163 (N_2163,N_2003,N_2075);
xor U2164 (N_2164,N_2087,N_2073);
or U2165 (N_2165,N_2011,N_2008);
nand U2166 (N_2166,N_2020,N_2031);
nand U2167 (N_2167,N_2040,N_2059);
xor U2168 (N_2168,N_2005,N_2088);
nor U2169 (N_2169,N_2001,N_2066);
and U2170 (N_2170,N_2018,N_2067);
and U2171 (N_2171,N_2088,N_2076);
nor U2172 (N_2172,N_2034,N_2086);
or U2173 (N_2173,N_2075,N_2092);
nor U2174 (N_2174,N_2047,N_2089);
and U2175 (N_2175,N_2067,N_2013);
or U2176 (N_2176,N_2068,N_2018);
and U2177 (N_2177,N_2030,N_2016);
or U2178 (N_2178,N_2045,N_2063);
and U2179 (N_2179,N_2043,N_2007);
or U2180 (N_2180,N_2049,N_2064);
nand U2181 (N_2181,N_2025,N_2047);
nand U2182 (N_2182,N_2059,N_2053);
nor U2183 (N_2183,N_2096,N_2050);
or U2184 (N_2184,N_2057,N_2006);
and U2185 (N_2185,N_2066,N_2005);
nand U2186 (N_2186,N_2054,N_2052);
xnor U2187 (N_2187,N_2092,N_2010);
nor U2188 (N_2188,N_2077,N_2043);
nand U2189 (N_2189,N_2064,N_2021);
xnor U2190 (N_2190,N_2003,N_2035);
or U2191 (N_2191,N_2005,N_2016);
and U2192 (N_2192,N_2047,N_2032);
or U2193 (N_2193,N_2084,N_2027);
nor U2194 (N_2194,N_2009,N_2005);
nand U2195 (N_2195,N_2028,N_2012);
xnor U2196 (N_2196,N_2004,N_2039);
nor U2197 (N_2197,N_2058,N_2052);
or U2198 (N_2198,N_2045,N_2042);
or U2199 (N_2199,N_2010,N_2069);
nor U2200 (N_2200,N_2150,N_2142);
nor U2201 (N_2201,N_2190,N_2168);
xnor U2202 (N_2202,N_2107,N_2122);
and U2203 (N_2203,N_2117,N_2129);
nor U2204 (N_2204,N_2188,N_2134);
or U2205 (N_2205,N_2171,N_2103);
nor U2206 (N_2206,N_2140,N_2136);
and U2207 (N_2207,N_2153,N_2132);
nand U2208 (N_2208,N_2176,N_2172);
nand U2209 (N_2209,N_2151,N_2119);
or U2210 (N_2210,N_2154,N_2111);
nor U2211 (N_2211,N_2169,N_2127);
nand U2212 (N_2212,N_2177,N_2161);
nor U2213 (N_2213,N_2141,N_2197);
nand U2214 (N_2214,N_2100,N_2184);
and U2215 (N_2215,N_2126,N_2106);
or U2216 (N_2216,N_2158,N_2191);
xor U2217 (N_2217,N_2109,N_2178);
nor U2218 (N_2218,N_2113,N_2164);
or U2219 (N_2219,N_2114,N_2124);
and U2220 (N_2220,N_2123,N_2128);
and U2221 (N_2221,N_2199,N_2170);
nor U2222 (N_2222,N_2102,N_2160);
nor U2223 (N_2223,N_2193,N_2147);
xor U2224 (N_2224,N_2104,N_2125);
or U2225 (N_2225,N_2156,N_2115);
or U2226 (N_2226,N_2121,N_2137);
nor U2227 (N_2227,N_2131,N_2120);
or U2228 (N_2228,N_2159,N_2166);
and U2229 (N_2229,N_2135,N_2157);
and U2230 (N_2230,N_2105,N_2133);
nand U2231 (N_2231,N_2144,N_2138);
nor U2232 (N_2232,N_2101,N_2116);
nor U2233 (N_2233,N_2118,N_2139);
or U2234 (N_2234,N_2185,N_2186);
nand U2235 (N_2235,N_2162,N_2174);
or U2236 (N_2236,N_2146,N_2145);
xnor U2237 (N_2237,N_2181,N_2112);
nor U2238 (N_2238,N_2110,N_2148);
nand U2239 (N_2239,N_2152,N_2163);
nand U2240 (N_2240,N_2167,N_2175);
or U2241 (N_2241,N_2194,N_2182);
or U2242 (N_2242,N_2130,N_2155);
and U2243 (N_2243,N_2165,N_2192);
or U2244 (N_2244,N_2189,N_2183);
nand U2245 (N_2245,N_2143,N_2180);
nand U2246 (N_2246,N_2195,N_2196);
nand U2247 (N_2247,N_2187,N_2108);
nand U2248 (N_2248,N_2149,N_2179);
and U2249 (N_2249,N_2173,N_2198);
nand U2250 (N_2250,N_2154,N_2195);
or U2251 (N_2251,N_2184,N_2134);
and U2252 (N_2252,N_2172,N_2108);
nand U2253 (N_2253,N_2176,N_2160);
xnor U2254 (N_2254,N_2158,N_2182);
or U2255 (N_2255,N_2102,N_2124);
nand U2256 (N_2256,N_2132,N_2100);
nor U2257 (N_2257,N_2182,N_2174);
and U2258 (N_2258,N_2153,N_2184);
nor U2259 (N_2259,N_2185,N_2127);
and U2260 (N_2260,N_2142,N_2137);
nor U2261 (N_2261,N_2116,N_2161);
and U2262 (N_2262,N_2130,N_2197);
nor U2263 (N_2263,N_2177,N_2106);
or U2264 (N_2264,N_2126,N_2121);
nand U2265 (N_2265,N_2160,N_2128);
nor U2266 (N_2266,N_2136,N_2179);
or U2267 (N_2267,N_2186,N_2195);
nor U2268 (N_2268,N_2129,N_2126);
or U2269 (N_2269,N_2117,N_2101);
and U2270 (N_2270,N_2192,N_2173);
or U2271 (N_2271,N_2159,N_2101);
and U2272 (N_2272,N_2154,N_2196);
and U2273 (N_2273,N_2146,N_2134);
nor U2274 (N_2274,N_2185,N_2190);
nand U2275 (N_2275,N_2178,N_2148);
xnor U2276 (N_2276,N_2181,N_2191);
nor U2277 (N_2277,N_2189,N_2101);
and U2278 (N_2278,N_2117,N_2149);
nand U2279 (N_2279,N_2120,N_2145);
and U2280 (N_2280,N_2178,N_2163);
xnor U2281 (N_2281,N_2104,N_2134);
or U2282 (N_2282,N_2181,N_2193);
nand U2283 (N_2283,N_2107,N_2128);
nor U2284 (N_2284,N_2186,N_2157);
nand U2285 (N_2285,N_2169,N_2190);
or U2286 (N_2286,N_2110,N_2154);
or U2287 (N_2287,N_2146,N_2155);
and U2288 (N_2288,N_2116,N_2168);
or U2289 (N_2289,N_2111,N_2138);
nand U2290 (N_2290,N_2108,N_2105);
xnor U2291 (N_2291,N_2150,N_2159);
xor U2292 (N_2292,N_2142,N_2140);
xnor U2293 (N_2293,N_2103,N_2175);
and U2294 (N_2294,N_2156,N_2157);
nor U2295 (N_2295,N_2141,N_2158);
and U2296 (N_2296,N_2136,N_2195);
and U2297 (N_2297,N_2139,N_2177);
nor U2298 (N_2298,N_2170,N_2139);
nor U2299 (N_2299,N_2112,N_2145);
xor U2300 (N_2300,N_2218,N_2252);
xor U2301 (N_2301,N_2287,N_2299);
and U2302 (N_2302,N_2204,N_2225);
or U2303 (N_2303,N_2297,N_2228);
xnor U2304 (N_2304,N_2217,N_2211);
and U2305 (N_2305,N_2270,N_2273);
nand U2306 (N_2306,N_2293,N_2236);
nand U2307 (N_2307,N_2229,N_2213);
nor U2308 (N_2308,N_2223,N_2242);
nor U2309 (N_2309,N_2208,N_2251);
and U2310 (N_2310,N_2230,N_2209);
nor U2311 (N_2311,N_2274,N_2216);
or U2312 (N_2312,N_2222,N_2240);
or U2313 (N_2313,N_2214,N_2210);
or U2314 (N_2314,N_2263,N_2291);
or U2315 (N_2315,N_2212,N_2245);
nor U2316 (N_2316,N_2239,N_2250);
xnor U2317 (N_2317,N_2255,N_2265);
and U2318 (N_2318,N_2244,N_2221);
and U2319 (N_2319,N_2281,N_2290);
xor U2320 (N_2320,N_2206,N_2298);
nor U2321 (N_2321,N_2205,N_2271);
nand U2322 (N_2322,N_2266,N_2215);
and U2323 (N_2323,N_2233,N_2267);
xor U2324 (N_2324,N_2203,N_2226);
nand U2325 (N_2325,N_2269,N_2220);
nor U2326 (N_2326,N_2289,N_2256);
nor U2327 (N_2327,N_2232,N_2277);
or U2328 (N_2328,N_2237,N_2257);
or U2329 (N_2329,N_2285,N_2243);
nor U2330 (N_2330,N_2207,N_2235);
or U2331 (N_2331,N_2279,N_2241);
nand U2332 (N_2332,N_2238,N_2201);
or U2333 (N_2333,N_2248,N_2261);
nor U2334 (N_2334,N_2296,N_2260);
or U2335 (N_2335,N_2200,N_2259);
and U2336 (N_2336,N_2288,N_2282);
nor U2337 (N_2337,N_2264,N_2219);
nor U2338 (N_2338,N_2275,N_2224);
or U2339 (N_2339,N_2284,N_2227);
and U2340 (N_2340,N_2268,N_2286);
or U2341 (N_2341,N_2249,N_2292);
or U2342 (N_2342,N_2262,N_2231);
or U2343 (N_2343,N_2294,N_2280);
nand U2344 (N_2344,N_2202,N_2253);
xnor U2345 (N_2345,N_2272,N_2258);
and U2346 (N_2346,N_2234,N_2246);
and U2347 (N_2347,N_2278,N_2295);
nand U2348 (N_2348,N_2247,N_2254);
nor U2349 (N_2349,N_2276,N_2283);
nand U2350 (N_2350,N_2243,N_2281);
xor U2351 (N_2351,N_2219,N_2212);
and U2352 (N_2352,N_2292,N_2240);
xnor U2353 (N_2353,N_2215,N_2201);
nor U2354 (N_2354,N_2295,N_2233);
or U2355 (N_2355,N_2251,N_2253);
nand U2356 (N_2356,N_2276,N_2252);
xnor U2357 (N_2357,N_2260,N_2235);
nor U2358 (N_2358,N_2230,N_2215);
nor U2359 (N_2359,N_2240,N_2284);
xnor U2360 (N_2360,N_2231,N_2287);
or U2361 (N_2361,N_2239,N_2277);
and U2362 (N_2362,N_2269,N_2274);
and U2363 (N_2363,N_2287,N_2255);
nand U2364 (N_2364,N_2246,N_2228);
and U2365 (N_2365,N_2260,N_2263);
and U2366 (N_2366,N_2250,N_2236);
nand U2367 (N_2367,N_2287,N_2274);
xnor U2368 (N_2368,N_2204,N_2251);
or U2369 (N_2369,N_2210,N_2215);
xnor U2370 (N_2370,N_2282,N_2287);
xnor U2371 (N_2371,N_2212,N_2258);
and U2372 (N_2372,N_2262,N_2267);
nor U2373 (N_2373,N_2287,N_2271);
and U2374 (N_2374,N_2255,N_2211);
and U2375 (N_2375,N_2249,N_2293);
and U2376 (N_2376,N_2299,N_2239);
xnor U2377 (N_2377,N_2280,N_2246);
nor U2378 (N_2378,N_2214,N_2279);
nand U2379 (N_2379,N_2286,N_2257);
or U2380 (N_2380,N_2266,N_2289);
xor U2381 (N_2381,N_2295,N_2287);
or U2382 (N_2382,N_2280,N_2253);
and U2383 (N_2383,N_2235,N_2231);
xnor U2384 (N_2384,N_2297,N_2278);
xnor U2385 (N_2385,N_2288,N_2220);
nor U2386 (N_2386,N_2211,N_2249);
nor U2387 (N_2387,N_2273,N_2298);
xor U2388 (N_2388,N_2254,N_2218);
xnor U2389 (N_2389,N_2257,N_2269);
nand U2390 (N_2390,N_2219,N_2284);
nor U2391 (N_2391,N_2223,N_2277);
or U2392 (N_2392,N_2232,N_2203);
nor U2393 (N_2393,N_2206,N_2227);
nand U2394 (N_2394,N_2229,N_2205);
nor U2395 (N_2395,N_2280,N_2240);
nand U2396 (N_2396,N_2249,N_2286);
nand U2397 (N_2397,N_2220,N_2236);
nand U2398 (N_2398,N_2241,N_2272);
nand U2399 (N_2399,N_2233,N_2269);
xnor U2400 (N_2400,N_2311,N_2353);
and U2401 (N_2401,N_2306,N_2315);
nor U2402 (N_2402,N_2337,N_2318);
or U2403 (N_2403,N_2313,N_2372);
nor U2404 (N_2404,N_2363,N_2362);
or U2405 (N_2405,N_2346,N_2393);
or U2406 (N_2406,N_2375,N_2371);
and U2407 (N_2407,N_2364,N_2342);
or U2408 (N_2408,N_2369,N_2314);
and U2409 (N_2409,N_2316,N_2339);
or U2410 (N_2410,N_2386,N_2330);
and U2411 (N_2411,N_2394,N_2321);
xor U2412 (N_2412,N_2352,N_2381);
or U2413 (N_2413,N_2359,N_2309);
nand U2414 (N_2414,N_2335,N_2378);
or U2415 (N_2415,N_2301,N_2308);
nor U2416 (N_2416,N_2323,N_2326);
and U2417 (N_2417,N_2354,N_2327);
and U2418 (N_2418,N_2347,N_2340);
nand U2419 (N_2419,N_2374,N_2317);
and U2420 (N_2420,N_2390,N_2380);
nor U2421 (N_2421,N_2396,N_2331);
nor U2422 (N_2422,N_2350,N_2357);
xor U2423 (N_2423,N_2303,N_2341);
nor U2424 (N_2424,N_2360,N_2398);
and U2425 (N_2425,N_2361,N_2302);
and U2426 (N_2426,N_2348,N_2377);
nor U2427 (N_2427,N_2376,N_2395);
nor U2428 (N_2428,N_2387,N_2344);
or U2429 (N_2429,N_2355,N_2343);
nand U2430 (N_2430,N_2373,N_2368);
or U2431 (N_2431,N_2379,N_2392);
and U2432 (N_2432,N_2324,N_2367);
nor U2433 (N_2433,N_2336,N_2389);
nor U2434 (N_2434,N_2334,N_2319);
nor U2435 (N_2435,N_2333,N_2349);
or U2436 (N_2436,N_2307,N_2310);
nor U2437 (N_2437,N_2312,N_2384);
and U2438 (N_2438,N_2351,N_2325);
nor U2439 (N_2439,N_2399,N_2305);
nand U2440 (N_2440,N_2397,N_2329);
nor U2441 (N_2441,N_2332,N_2322);
and U2442 (N_2442,N_2356,N_2385);
nand U2443 (N_2443,N_2366,N_2370);
nand U2444 (N_2444,N_2304,N_2358);
and U2445 (N_2445,N_2338,N_2391);
nor U2446 (N_2446,N_2300,N_2328);
nand U2447 (N_2447,N_2365,N_2345);
or U2448 (N_2448,N_2383,N_2382);
nand U2449 (N_2449,N_2388,N_2320);
nor U2450 (N_2450,N_2309,N_2327);
and U2451 (N_2451,N_2361,N_2328);
nor U2452 (N_2452,N_2312,N_2355);
and U2453 (N_2453,N_2323,N_2355);
nor U2454 (N_2454,N_2374,N_2322);
nor U2455 (N_2455,N_2348,N_2383);
or U2456 (N_2456,N_2390,N_2394);
and U2457 (N_2457,N_2381,N_2384);
xnor U2458 (N_2458,N_2305,N_2358);
nor U2459 (N_2459,N_2344,N_2349);
and U2460 (N_2460,N_2361,N_2332);
nand U2461 (N_2461,N_2354,N_2373);
nand U2462 (N_2462,N_2304,N_2398);
xor U2463 (N_2463,N_2329,N_2344);
xnor U2464 (N_2464,N_2322,N_2367);
or U2465 (N_2465,N_2338,N_2379);
nand U2466 (N_2466,N_2373,N_2341);
or U2467 (N_2467,N_2365,N_2342);
or U2468 (N_2468,N_2341,N_2344);
nor U2469 (N_2469,N_2383,N_2324);
xnor U2470 (N_2470,N_2316,N_2327);
or U2471 (N_2471,N_2354,N_2300);
xnor U2472 (N_2472,N_2331,N_2314);
and U2473 (N_2473,N_2369,N_2311);
nor U2474 (N_2474,N_2308,N_2360);
and U2475 (N_2475,N_2341,N_2356);
and U2476 (N_2476,N_2346,N_2313);
or U2477 (N_2477,N_2316,N_2379);
xor U2478 (N_2478,N_2399,N_2361);
nand U2479 (N_2479,N_2339,N_2345);
or U2480 (N_2480,N_2399,N_2390);
and U2481 (N_2481,N_2341,N_2332);
and U2482 (N_2482,N_2327,N_2311);
nor U2483 (N_2483,N_2301,N_2370);
and U2484 (N_2484,N_2382,N_2364);
xor U2485 (N_2485,N_2353,N_2358);
and U2486 (N_2486,N_2344,N_2358);
xnor U2487 (N_2487,N_2330,N_2308);
and U2488 (N_2488,N_2378,N_2360);
nor U2489 (N_2489,N_2315,N_2366);
xnor U2490 (N_2490,N_2394,N_2358);
nor U2491 (N_2491,N_2300,N_2375);
and U2492 (N_2492,N_2388,N_2337);
nor U2493 (N_2493,N_2341,N_2367);
or U2494 (N_2494,N_2370,N_2328);
nand U2495 (N_2495,N_2367,N_2318);
nor U2496 (N_2496,N_2392,N_2388);
and U2497 (N_2497,N_2347,N_2398);
or U2498 (N_2498,N_2385,N_2306);
xor U2499 (N_2499,N_2306,N_2393);
or U2500 (N_2500,N_2483,N_2470);
and U2501 (N_2501,N_2477,N_2462);
or U2502 (N_2502,N_2487,N_2455);
or U2503 (N_2503,N_2410,N_2405);
nor U2504 (N_2504,N_2402,N_2423);
and U2505 (N_2505,N_2441,N_2425);
nand U2506 (N_2506,N_2436,N_2432);
nand U2507 (N_2507,N_2475,N_2468);
nor U2508 (N_2508,N_2480,N_2452);
nor U2509 (N_2509,N_2478,N_2454);
nor U2510 (N_2510,N_2444,N_2493);
nor U2511 (N_2511,N_2416,N_2456);
and U2512 (N_2512,N_2431,N_2448);
or U2513 (N_2513,N_2471,N_2479);
xor U2514 (N_2514,N_2496,N_2427);
and U2515 (N_2515,N_2429,N_2474);
nor U2516 (N_2516,N_2495,N_2400);
or U2517 (N_2517,N_2457,N_2435);
and U2518 (N_2518,N_2445,N_2430);
or U2519 (N_2519,N_2491,N_2409);
or U2520 (N_2520,N_2428,N_2460);
nand U2521 (N_2521,N_2499,N_2473);
nand U2522 (N_2522,N_2414,N_2418);
nand U2523 (N_2523,N_2465,N_2467);
or U2524 (N_2524,N_2492,N_2469);
nand U2525 (N_2525,N_2415,N_2459);
or U2526 (N_2526,N_2407,N_2489);
or U2527 (N_2527,N_2424,N_2494);
and U2528 (N_2528,N_2437,N_2417);
or U2529 (N_2529,N_2472,N_2488);
xor U2530 (N_2530,N_2498,N_2421);
nor U2531 (N_2531,N_2446,N_2408);
nor U2532 (N_2532,N_2497,N_2453);
nor U2533 (N_2533,N_2484,N_2451);
nand U2534 (N_2534,N_2434,N_2485);
nand U2535 (N_2535,N_2438,N_2412);
nor U2536 (N_2536,N_2420,N_2422);
or U2537 (N_2537,N_2450,N_2481);
or U2538 (N_2538,N_2406,N_2426);
nor U2539 (N_2539,N_2433,N_2449);
and U2540 (N_2540,N_2419,N_2442);
xor U2541 (N_2541,N_2458,N_2476);
or U2542 (N_2542,N_2404,N_2466);
or U2543 (N_2543,N_2440,N_2461);
or U2544 (N_2544,N_2443,N_2439);
xnor U2545 (N_2545,N_2403,N_2490);
nor U2546 (N_2546,N_2447,N_2413);
and U2547 (N_2547,N_2482,N_2401);
or U2548 (N_2548,N_2463,N_2411);
and U2549 (N_2549,N_2486,N_2464);
nor U2550 (N_2550,N_2426,N_2405);
nor U2551 (N_2551,N_2404,N_2483);
and U2552 (N_2552,N_2448,N_2413);
xnor U2553 (N_2553,N_2468,N_2496);
nand U2554 (N_2554,N_2432,N_2464);
and U2555 (N_2555,N_2407,N_2481);
xor U2556 (N_2556,N_2486,N_2409);
nand U2557 (N_2557,N_2469,N_2459);
nor U2558 (N_2558,N_2401,N_2486);
xnor U2559 (N_2559,N_2416,N_2491);
nor U2560 (N_2560,N_2452,N_2402);
and U2561 (N_2561,N_2464,N_2435);
and U2562 (N_2562,N_2480,N_2461);
nor U2563 (N_2563,N_2436,N_2498);
and U2564 (N_2564,N_2419,N_2434);
and U2565 (N_2565,N_2482,N_2407);
and U2566 (N_2566,N_2404,N_2432);
nor U2567 (N_2567,N_2438,N_2450);
nor U2568 (N_2568,N_2401,N_2439);
nor U2569 (N_2569,N_2402,N_2443);
nor U2570 (N_2570,N_2496,N_2480);
nor U2571 (N_2571,N_2440,N_2441);
or U2572 (N_2572,N_2452,N_2403);
xor U2573 (N_2573,N_2496,N_2484);
and U2574 (N_2574,N_2429,N_2485);
nand U2575 (N_2575,N_2477,N_2459);
or U2576 (N_2576,N_2498,N_2490);
nand U2577 (N_2577,N_2495,N_2477);
xor U2578 (N_2578,N_2486,N_2405);
or U2579 (N_2579,N_2410,N_2494);
nor U2580 (N_2580,N_2450,N_2443);
or U2581 (N_2581,N_2492,N_2477);
and U2582 (N_2582,N_2438,N_2483);
or U2583 (N_2583,N_2490,N_2439);
xnor U2584 (N_2584,N_2471,N_2401);
nand U2585 (N_2585,N_2457,N_2497);
xnor U2586 (N_2586,N_2451,N_2470);
and U2587 (N_2587,N_2448,N_2471);
nor U2588 (N_2588,N_2477,N_2483);
or U2589 (N_2589,N_2446,N_2424);
or U2590 (N_2590,N_2485,N_2470);
nor U2591 (N_2591,N_2483,N_2445);
nand U2592 (N_2592,N_2483,N_2451);
nor U2593 (N_2593,N_2457,N_2411);
and U2594 (N_2594,N_2456,N_2497);
or U2595 (N_2595,N_2416,N_2407);
nand U2596 (N_2596,N_2468,N_2470);
nor U2597 (N_2597,N_2451,N_2430);
or U2598 (N_2598,N_2497,N_2428);
nand U2599 (N_2599,N_2432,N_2461);
nand U2600 (N_2600,N_2517,N_2589);
nand U2601 (N_2601,N_2522,N_2573);
xor U2602 (N_2602,N_2510,N_2567);
nand U2603 (N_2603,N_2588,N_2546);
and U2604 (N_2604,N_2590,N_2514);
or U2605 (N_2605,N_2592,N_2504);
nor U2606 (N_2606,N_2506,N_2585);
or U2607 (N_2607,N_2547,N_2525);
xnor U2608 (N_2608,N_2551,N_2536);
or U2609 (N_2609,N_2501,N_2596);
and U2610 (N_2610,N_2503,N_2576);
or U2611 (N_2611,N_2584,N_2594);
nor U2612 (N_2612,N_2561,N_2532);
nand U2613 (N_2613,N_2597,N_2515);
or U2614 (N_2614,N_2570,N_2558);
and U2615 (N_2615,N_2580,N_2559);
nand U2616 (N_2616,N_2507,N_2513);
and U2617 (N_2617,N_2562,N_2538);
nor U2618 (N_2618,N_2595,N_2524);
nor U2619 (N_2619,N_2540,N_2557);
nor U2620 (N_2620,N_2518,N_2581);
or U2621 (N_2621,N_2577,N_2578);
or U2622 (N_2622,N_2565,N_2575);
or U2623 (N_2623,N_2568,N_2550);
xor U2624 (N_2624,N_2502,N_2539);
nand U2625 (N_2625,N_2548,N_2587);
nand U2626 (N_2626,N_2512,N_2523);
or U2627 (N_2627,N_2544,N_2519);
nand U2628 (N_2628,N_2531,N_2505);
nand U2629 (N_2629,N_2591,N_2560);
nor U2630 (N_2630,N_2572,N_2508);
or U2631 (N_2631,N_2579,N_2528);
nand U2632 (N_2632,N_2500,N_2556);
nand U2633 (N_2633,N_2541,N_2526);
xnor U2634 (N_2634,N_2527,N_2574);
or U2635 (N_2635,N_2516,N_2593);
xnor U2636 (N_2636,N_2564,N_2509);
nand U2637 (N_2637,N_2599,N_2566);
and U2638 (N_2638,N_2521,N_2582);
or U2639 (N_2639,N_2542,N_2569);
nor U2640 (N_2640,N_2529,N_2586);
nand U2641 (N_2641,N_2553,N_2535);
nand U2642 (N_2642,N_2598,N_2537);
and U2643 (N_2643,N_2534,N_2571);
nand U2644 (N_2644,N_2583,N_2552);
nand U2645 (N_2645,N_2511,N_2555);
nand U2646 (N_2646,N_2549,N_2533);
and U2647 (N_2647,N_2543,N_2520);
nand U2648 (N_2648,N_2554,N_2545);
xor U2649 (N_2649,N_2563,N_2530);
and U2650 (N_2650,N_2567,N_2566);
and U2651 (N_2651,N_2548,N_2516);
or U2652 (N_2652,N_2544,N_2521);
and U2653 (N_2653,N_2562,N_2539);
and U2654 (N_2654,N_2568,N_2556);
xnor U2655 (N_2655,N_2528,N_2537);
and U2656 (N_2656,N_2594,N_2525);
nor U2657 (N_2657,N_2599,N_2547);
and U2658 (N_2658,N_2580,N_2592);
nand U2659 (N_2659,N_2511,N_2529);
nand U2660 (N_2660,N_2552,N_2511);
nand U2661 (N_2661,N_2574,N_2518);
and U2662 (N_2662,N_2503,N_2554);
nand U2663 (N_2663,N_2532,N_2511);
and U2664 (N_2664,N_2555,N_2589);
and U2665 (N_2665,N_2545,N_2580);
nand U2666 (N_2666,N_2541,N_2503);
nand U2667 (N_2667,N_2541,N_2561);
or U2668 (N_2668,N_2505,N_2558);
xor U2669 (N_2669,N_2591,N_2548);
or U2670 (N_2670,N_2582,N_2590);
nor U2671 (N_2671,N_2591,N_2538);
nor U2672 (N_2672,N_2556,N_2508);
nor U2673 (N_2673,N_2593,N_2524);
or U2674 (N_2674,N_2564,N_2533);
xnor U2675 (N_2675,N_2520,N_2576);
xnor U2676 (N_2676,N_2540,N_2550);
or U2677 (N_2677,N_2595,N_2523);
xnor U2678 (N_2678,N_2523,N_2575);
nand U2679 (N_2679,N_2593,N_2563);
nor U2680 (N_2680,N_2571,N_2514);
nand U2681 (N_2681,N_2526,N_2506);
and U2682 (N_2682,N_2524,N_2597);
nand U2683 (N_2683,N_2562,N_2516);
xnor U2684 (N_2684,N_2535,N_2529);
nor U2685 (N_2685,N_2541,N_2537);
nor U2686 (N_2686,N_2594,N_2521);
and U2687 (N_2687,N_2550,N_2582);
nand U2688 (N_2688,N_2570,N_2588);
and U2689 (N_2689,N_2583,N_2522);
nand U2690 (N_2690,N_2597,N_2533);
and U2691 (N_2691,N_2584,N_2579);
and U2692 (N_2692,N_2597,N_2510);
nor U2693 (N_2693,N_2585,N_2533);
nand U2694 (N_2694,N_2504,N_2563);
or U2695 (N_2695,N_2597,N_2520);
or U2696 (N_2696,N_2585,N_2574);
xnor U2697 (N_2697,N_2520,N_2593);
or U2698 (N_2698,N_2583,N_2591);
and U2699 (N_2699,N_2576,N_2570);
or U2700 (N_2700,N_2692,N_2680);
nor U2701 (N_2701,N_2638,N_2688);
nor U2702 (N_2702,N_2661,N_2689);
nand U2703 (N_2703,N_2629,N_2686);
or U2704 (N_2704,N_2662,N_2615);
and U2705 (N_2705,N_2669,N_2697);
and U2706 (N_2706,N_2600,N_2636);
nand U2707 (N_2707,N_2652,N_2687);
or U2708 (N_2708,N_2622,N_2676);
or U2709 (N_2709,N_2668,N_2657);
nor U2710 (N_2710,N_2602,N_2639);
xor U2711 (N_2711,N_2646,N_2637);
and U2712 (N_2712,N_2691,N_2653);
and U2713 (N_2713,N_2665,N_2619);
and U2714 (N_2714,N_2633,N_2612);
nand U2715 (N_2715,N_2614,N_2630);
nor U2716 (N_2716,N_2677,N_2666);
xnor U2717 (N_2717,N_2675,N_2651);
or U2718 (N_2718,N_2682,N_2672);
and U2719 (N_2719,N_2611,N_2603);
or U2720 (N_2720,N_2696,N_2607);
nor U2721 (N_2721,N_2644,N_2634);
nand U2722 (N_2722,N_2690,N_2640);
nand U2723 (N_2723,N_2608,N_2667);
and U2724 (N_2724,N_2670,N_2658);
or U2725 (N_2725,N_2685,N_2601);
and U2726 (N_2726,N_2660,N_2698);
or U2727 (N_2727,N_2699,N_2635);
or U2728 (N_2728,N_2681,N_2616);
and U2729 (N_2729,N_2613,N_2626);
or U2730 (N_2730,N_2604,N_2674);
xnor U2731 (N_2731,N_2673,N_2645);
or U2732 (N_2732,N_2632,N_2695);
nor U2733 (N_2733,N_2648,N_2606);
or U2734 (N_2734,N_2617,N_2694);
or U2735 (N_2735,N_2628,N_2643);
and U2736 (N_2736,N_2610,N_2631);
nor U2737 (N_2737,N_2693,N_2655);
nand U2738 (N_2738,N_2642,N_2627);
and U2739 (N_2739,N_2659,N_2683);
nand U2740 (N_2740,N_2641,N_2679);
xor U2741 (N_2741,N_2649,N_2671);
nor U2742 (N_2742,N_2647,N_2618);
xor U2743 (N_2743,N_2605,N_2620);
nor U2744 (N_2744,N_2624,N_2656);
nor U2745 (N_2745,N_2684,N_2678);
nand U2746 (N_2746,N_2664,N_2625);
or U2747 (N_2747,N_2663,N_2609);
xnor U2748 (N_2748,N_2654,N_2650);
nor U2749 (N_2749,N_2621,N_2623);
or U2750 (N_2750,N_2671,N_2647);
nand U2751 (N_2751,N_2679,N_2651);
xor U2752 (N_2752,N_2691,N_2616);
xnor U2753 (N_2753,N_2650,N_2632);
or U2754 (N_2754,N_2681,N_2684);
and U2755 (N_2755,N_2672,N_2636);
or U2756 (N_2756,N_2620,N_2669);
nand U2757 (N_2757,N_2667,N_2687);
or U2758 (N_2758,N_2662,N_2650);
nor U2759 (N_2759,N_2609,N_2683);
nor U2760 (N_2760,N_2601,N_2631);
nor U2761 (N_2761,N_2645,N_2658);
and U2762 (N_2762,N_2620,N_2630);
nor U2763 (N_2763,N_2670,N_2611);
nor U2764 (N_2764,N_2650,N_2607);
nor U2765 (N_2765,N_2632,N_2610);
or U2766 (N_2766,N_2692,N_2688);
xnor U2767 (N_2767,N_2693,N_2611);
nor U2768 (N_2768,N_2691,N_2636);
or U2769 (N_2769,N_2617,N_2616);
nand U2770 (N_2770,N_2676,N_2609);
nand U2771 (N_2771,N_2630,N_2628);
and U2772 (N_2772,N_2622,N_2672);
nor U2773 (N_2773,N_2686,N_2676);
xor U2774 (N_2774,N_2608,N_2675);
nand U2775 (N_2775,N_2681,N_2656);
nand U2776 (N_2776,N_2670,N_2609);
nand U2777 (N_2777,N_2609,N_2632);
and U2778 (N_2778,N_2604,N_2668);
nand U2779 (N_2779,N_2639,N_2688);
and U2780 (N_2780,N_2628,N_2610);
nor U2781 (N_2781,N_2609,N_2615);
or U2782 (N_2782,N_2674,N_2648);
or U2783 (N_2783,N_2603,N_2634);
nand U2784 (N_2784,N_2668,N_2664);
or U2785 (N_2785,N_2602,N_2685);
and U2786 (N_2786,N_2626,N_2635);
nand U2787 (N_2787,N_2680,N_2616);
or U2788 (N_2788,N_2613,N_2631);
nor U2789 (N_2789,N_2634,N_2668);
xnor U2790 (N_2790,N_2620,N_2681);
nor U2791 (N_2791,N_2651,N_2673);
or U2792 (N_2792,N_2656,N_2631);
or U2793 (N_2793,N_2644,N_2609);
xnor U2794 (N_2794,N_2671,N_2609);
or U2795 (N_2795,N_2643,N_2691);
nor U2796 (N_2796,N_2618,N_2652);
or U2797 (N_2797,N_2650,N_2613);
nand U2798 (N_2798,N_2672,N_2658);
and U2799 (N_2799,N_2658,N_2695);
and U2800 (N_2800,N_2726,N_2718);
and U2801 (N_2801,N_2759,N_2731);
or U2802 (N_2802,N_2764,N_2749);
nand U2803 (N_2803,N_2748,N_2730);
nor U2804 (N_2804,N_2723,N_2716);
nand U2805 (N_2805,N_2753,N_2713);
nand U2806 (N_2806,N_2735,N_2776);
nand U2807 (N_2807,N_2798,N_2783);
nand U2808 (N_2808,N_2724,N_2741);
and U2809 (N_2809,N_2797,N_2743);
or U2810 (N_2810,N_2717,N_2772);
nor U2811 (N_2811,N_2789,N_2763);
and U2812 (N_2812,N_2701,N_2769);
xor U2813 (N_2813,N_2762,N_2719);
nor U2814 (N_2814,N_2768,N_2733);
nor U2815 (N_2815,N_2779,N_2746);
and U2816 (N_2816,N_2761,N_2740);
nand U2817 (N_2817,N_2765,N_2705);
and U2818 (N_2818,N_2736,N_2738);
and U2819 (N_2819,N_2714,N_2706);
and U2820 (N_2820,N_2785,N_2770);
and U2821 (N_2821,N_2775,N_2737);
or U2822 (N_2822,N_2794,N_2744);
or U2823 (N_2823,N_2773,N_2781);
or U2824 (N_2824,N_2766,N_2792);
or U2825 (N_2825,N_2727,N_2782);
and U2826 (N_2826,N_2777,N_2728);
or U2827 (N_2827,N_2725,N_2703);
or U2828 (N_2828,N_2742,N_2734);
nor U2829 (N_2829,N_2739,N_2732);
nor U2830 (N_2830,N_2700,N_2786);
or U2831 (N_2831,N_2708,N_2787);
or U2832 (N_2832,N_2788,N_2704);
nor U2833 (N_2833,N_2754,N_2720);
and U2834 (N_2834,N_2760,N_2757);
or U2835 (N_2835,N_2793,N_2702);
xnor U2836 (N_2836,N_2767,N_2750);
and U2837 (N_2837,N_2774,N_2722);
or U2838 (N_2838,N_2747,N_2752);
nor U2839 (N_2839,N_2709,N_2721);
nand U2840 (N_2840,N_2715,N_2780);
nand U2841 (N_2841,N_2707,N_2751);
and U2842 (N_2842,N_2771,N_2799);
xor U2843 (N_2843,N_2791,N_2790);
and U2844 (N_2844,N_2755,N_2756);
nand U2845 (N_2845,N_2745,N_2710);
nor U2846 (N_2846,N_2795,N_2729);
nor U2847 (N_2847,N_2712,N_2778);
and U2848 (N_2848,N_2711,N_2796);
or U2849 (N_2849,N_2758,N_2784);
nand U2850 (N_2850,N_2748,N_2757);
nand U2851 (N_2851,N_2709,N_2799);
nor U2852 (N_2852,N_2739,N_2799);
nor U2853 (N_2853,N_2767,N_2718);
nand U2854 (N_2854,N_2728,N_2776);
or U2855 (N_2855,N_2725,N_2748);
nand U2856 (N_2856,N_2791,N_2710);
nand U2857 (N_2857,N_2778,N_2761);
and U2858 (N_2858,N_2740,N_2791);
nand U2859 (N_2859,N_2760,N_2750);
and U2860 (N_2860,N_2739,N_2786);
nand U2861 (N_2861,N_2741,N_2715);
and U2862 (N_2862,N_2745,N_2714);
and U2863 (N_2863,N_2754,N_2765);
nand U2864 (N_2864,N_2793,N_2781);
or U2865 (N_2865,N_2707,N_2744);
or U2866 (N_2866,N_2712,N_2748);
and U2867 (N_2867,N_2736,N_2768);
and U2868 (N_2868,N_2762,N_2768);
or U2869 (N_2869,N_2752,N_2712);
nand U2870 (N_2870,N_2750,N_2765);
nor U2871 (N_2871,N_2747,N_2734);
xnor U2872 (N_2872,N_2707,N_2724);
nor U2873 (N_2873,N_2720,N_2703);
nand U2874 (N_2874,N_2758,N_2744);
xnor U2875 (N_2875,N_2702,N_2790);
and U2876 (N_2876,N_2720,N_2765);
and U2877 (N_2877,N_2735,N_2792);
nor U2878 (N_2878,N_2792,N_2759);
nand U2879 (N_2879,N_2744,N_2733);
nor U2880 (N_2880,N_2775,N_2711);
and U2881 (N_2881,N_2725,N_2712);
nor U2882 (N_2882,N_2775,N_2713);
nor U2883 (N_2883,N_2721,N_2751);
and U2884 (N_2884,N_2715,N_2712);
nor U2885 (N_2885,N_2719,N_2766);
nand U2886 (N_2886,N_2767,N_2733);
or U2887 (N_2887,N_2748,N_2722);
nor U2888 (N_2888,N_2736,N_2794);
or U2889 (N_2889,N_2714,N_2774);
nand U2890 (N_2890,N_2797,N_2737);
xnor U2891 (N_2891,N_2730,N_2709);
and U2892 (N_2892,N_2703,N_2748);
nand U2893 (N_2893,N_2758,N_2757);
xor U2894 (N_2894,N_2712,N_2714);
or U2895 (N_2895,N_2744,N_2741);
nand U2896 (N_2896,N_2739,N_2781);
nor U2897 (N_2897,N_2771,N_2723);
or U2898 (N_2898,N_2794,N_2707);
nor U2899 (N_2899,N_2739,N_2740);
or U2900 (N_2900,N_2898,N_2879);
and U2901 (N_2901,N_2802,N_2818);
or U2902 (N_2902,N_2854,N_2841);
nor U2903 (N_2903,N_2856,N_2847);
xnor U2904 (N_2904,N_2892,N_2870);
nor U2905 (N_2905,N_2803,N_2827);
or U2906 (N_2906,N_2899,N_2881);
nand U2907 (N_2907,N_2839,N_2840);
nand U2908 (N_2908,N_2884,N_2885);
or U2909 (N_2909,N_2897,N_2846);
and U2910 (N_2910,N_2886,N_2814);
or U2911 (N_2911,N_2833,N_2804);
nand U2912 (N_2912,N_2861,N_2820);
nor U2913 (N_2913,N_2844,N_2865);
nand U2914 (N_2914,N_2888,N_2864);
nor U2915 (N_2915,N_2894,N_2807);
xor U2916 (N_2916,N_2806,N_2890);
or U2917 (N_2917,N_2821,N_2862);
nand U2918 (N_2918,N_2809,N_2877);
nand U2919 (N_2919,N_2817,N_2883);
nor U2920 (N_2920,N_2811,N_2875);
xor U2921 (N_2921,N_2868,N_2843);
nand U2922 (N_2922,N_2826,N_2829);
or U2923 (N_2923,N_2822,N_2855);
or U2924 (N_2924,N_2812,N_2832);
xor U2925 (N_2925,N_2849,N_2834);
and U2926 (N_2926,N_2824,N_2842);
nor U2927 (N_2927,N_2845,N_2863);
nand U2928 (N_2928,N_2823,N_2873);
xor U2929 (N_2929,N_2895,N_2808);
and U2930 (N_2930,N_2866,N_2860);
nor U2931 (N_2931,N_2859,N_2880);
or U2932 (N_2932,N_2831,N_2852);
and U2933 (N_2933,N_2867,N_2825);
or U2934 (N_2934,N_2850,N_2857);
nor U2935 (N_2935,N_2816,N_2835);
nand U2936 (N_2936,N_2837,N_2819);
nor U2937 (N_2937,N_2872,N_2813);
or U2938 (N_2938,N_2889,N_2893);
or U2939 (N_2939,N_2896,N_2874);
or U2940 (N_2940,N_2891,N_2887);
or U2941 (N_2941,N_2815,N_2869);
nor U2942 (N_2942,N_2838,N_2828);
or U2943 (N_2943,N_2810,N_2878);
nor U2944 (N_2944,N_2882,N_2853);
nor U2945 (N_2945,N_2858,N_2830);
or U2946 (N_2946,N_2800,N_2871);
xor U2947 (N_2947,N_2805,N_2876);
nor U2948 (N_2948,N_2851,N_2836);
nor U2949 (N_2949,N_2848,N_2801);
nor U2950 (N_2950,N_2830,N_2878);
and U2951 (N_2951,N_2869,N_2898);
nand U2952 (N_2952,N_2868,N_2842);
or U2953 (N_2953,N_2812,N_2828);
and U2954 (N_2954,N_2809,N_2803);
nor U2955 (N_2955,N_2801,N_2879);
nor U2956 (N_2956,N_2867,N_2804);
nor U2957 (N_2957,N_2892,N_2896);
nand U2958 (N_2958,N_2838,N_2845);
and U2959 (N_2959,N_2878,N_2867);
and U2960 (N_2960,N_2883,N_2899);
and U2961 (N_2961,N_2814,N_2893);
nor U2962 (N_2962,N_2846,N_2872);
nand U2963 (N_2963,N_2850,N_2887);
nand U2964 (N_2964,N_2823,N_2805);
xor U2965 (N_2965,N_2894,N_2806);
nor U2966 (N_2966,N_2871,N_2883);
nand U2967 (N_2967,N_2829,N_2836);
nand U2968 (N_2968,N_2883,N_2874);
nand U2969 (N_2969,N_2895,N_2873);
xor U2970 (N_2970,N_2875,N_2821);
nand U2971 (N_2971,N_2849,N_2875);
nand U2972 (N_2972,N_2827,N_2822);
nand U2973 (N_2973,N_2855,N_2802);
nand U2974 (N_2974,N_2831,N_2884);
and U2975 (N_2975,N_2881,N_2818);
and U2976 (N_2976,N_2841,N_2808);
nand U2977 (N_2977,N_2842,N_2874);
or U2978 (N_2978,N_2836,N_2840);
nand U2979 (N_2979,N_2860,N_2881);
nand U2980 (N_2980,N_2834,N_2813);
or U2981 (N_2981,N_2857,N_2848);
nor U2982 (N_2982,N_2841,N_2863);
or U2983 (N_2983,N_2855,N_2885);
nand U2984 (N_2984,N_2872,N_2898);
nor U2985 (N_2985,N_2833,N_2810);
nand U2986 (N_2986,N_2810,N_2863);
and U2987 (N_2987,N_2865,N_2810);
nor U2988 (N_2988,N_2842,N_2801);
and U2989 (N_2989,N_2886,N_2864);
nor U2990 (N_2990,N_2828,N_2830);
nor U2991 (N_2991,N_2849,N_2856);
nor U2992 (N_2992,N_2827,N_2865);
and U2993 (N_2993,N_2873,N_2801);
and U2994 (N_2994,N_2847,N_2823);
nor U2995 (N_2995,N_2828,N_2808);
and U2996 (N_2996,N_2836,N_2872);
or U2997 (N_2997,N_2881,N_2842);
nor U2998 (N_2998,N_2845,N_2886);
and U2999 (N_2999,N_2891,N_2840);
and U3000 (N_3000,N_2921,N_2989);
nor U3001 (N_3001,N_2996,N_2935);
and U3002 (N_3002,N_2953,N_2978);
nor U3003 (N_3003,N_2991,N_2909);
or U3004 (N_3004,N_2971,N_2941);
xor U3005 (N_3005,N_2961,N_2904);
and U3006 (N_3006,N_2992,N_2988);
nor U3007 (N_3007,N_2962,N_2929);
nor U3008 (N_3008,N_2920,N_2965);
nand U3009 (N_3009,N_2932,N_2934);
or U3010 (N_3010,N_2925,N_2979);
nand U3011 (N_3011,N_2942,N_2915);
or U3012 (N_3012,N_2956,N_2918);
nor U3013 (N_3013,N_2970,N_2923);
nand U3014 (N_3014,N_2931,N_2903);
and U3015 (N_3015,N_2940,N_2933);
nor U3016 (N_3016,N_2913,N_2998);
or U3017 (N_3017,N_2946,N_2950);
or U3018 (N_3018,N_2901,N_2930);
xor U3019 (N_3019,N_2972,N_2982);
nand U3020 (N_3020,N_2995,N_2900);
and U3021 (N_3021,N_2977,N_2924);
nand U3022 (N_3022,N_2919,N_2976);
nand U3023 (N_3023,N_2905,N_2960);
nor U3024 (N_3024,N_2926,N_2983);
nor U3025 (N_3025,N_2994,N_2959);
nor U3026 (N_3026,N_2912,N_2943);
xor U3027 (N_3027,N_2947,N_2927);
nand U3028 (N_3028,N_2999,N_2922);
or U3029 (N_3029,N_2916,N_2975);
xor U3030 (N_3030,N_2908,N_2911);
nor U3031 (N_3031,N_2907,N_2986);
nor U3032 (N_3032,N_2997,N_2984);
or U3033 (N_3033,N_2910,N_2968);
nand U3034 (N_3034,N_2928,N_2949);
xor U3035 (N_3035,N_2945,N_2954);
or U3036 (N_3036,N_2987,N_2993);
xor U3037 (N_3037,N_2936,N_2974);
and U3038 (N_3038,N_2948,N_2955);
nand U3039 (N_3039,N_2938,N_2952);
or U3040 (N_3040,N_2906,N_2964);
nand U3041 (N_3041,N_2902,N_2969);
nor U3042 (N_3042,N_2963,N_2951);
nor U3043 (N_3043,N_2939,N_2973);
and U3044 (N_3044,N_2990,N_2981);
and U3045 (N_3045,N_2985,N_2958);
xor U3046 (N_3046,N_2937,N_2957);
nor U3047 (N_3047,N_2914,N_2917);
nand U3048 (N_3048,N_2967,N_2944);
and U3049 (N_3049,N_2980,N_2966);
and U3050 (N_3050,N_2933,N_2971);
or U3051 (N_3051,N_2984,N_2979);
nor U3052 (N_3052,N_2990,N_2991);
or U3053 (N_3053,N_2914,N_2925);
xnor U3054 (N_3054,N_2961,N_2976);
nor U3055 (N_3055,N_2968,N_2947);
and U3056 (N_3056,N_2983,N_2957);
nor U3057 (N_3057,N_2923,N_2917);
and U3058 (N_3058,N_2999,N_2978);
or U3059 (N_3059,N_2903,N_2942);
nand U3060 (N_3060,N_2915,N_2945);
nor U3061 (N_3061,N_2993,N_2958);
or U3062 (N_3062,N_2991,N_2949);
nand U3063 (N_3063,N_2971,N_2906);
and U3064 (N_3064,N_2932,N_2938);
or U3065 (N_3065,N_2987,N_2963);
xnor U3066 (N_3066,N_2913,N_2908);
nor U3067 (N_3067,N_2904,N_2985);
nor U3068 (N_3068,N_2912,N_2980);
nand U3069 (N_3069,N_2963,N_2907);
or U3070 (N_3070,N_2980,N_2913);
nor U3071 (N_3071,N_2939,N_2959);
xor U3072 (N_3072,N_2967,N_2974);
nand U3073 (N_3073,N_2957,N_2932);
and U3074 (N_3074,N_2908,N_2981);
nand U3075 (N_3075,N_2944,N_2991);
and U3076 (N_3076,N_2982,N_2961);
xnor U3077 (N_3077,N_2912,N_2902);
or U3078 (N_3078,N_2928,N_2963);
nand U3079 (N_3079,N_2946,N_2991);
and U3080 (N_3080,N_2964,N_2957);
nor U3081 (N_3081,N_2944,N_2975);
and U3082 (N_3082,N_2906,N_2930);
nor U3083 (N_3083,N_2948,N_2912);
nor U3084 (N_3084,N_2959,N_2912);
or U3085 (N_3085,N_2964,N_2937);
or U3086 (N_3086,N_2927,N_2958);
nor U3087 (N_3087,N_2990,N_2960);
and U3088 (N_3088,N_2934,N_2971);
or U3089 (N_3089,N_2948,N_2936);
or U3090 (N_3090,N_2986,N_2983);
nand U3091 (N_3091,N_2953,N_2946);
or U3092 (N_3092,N_2938,N_2999);
nor U3093 (N_3093,N_2930,N_2940);
nor U3094 (N_3094,N_2910,N_2936);
and U3095 (N_3095,N_2928,N_2960);
or U3096 (N_3096,N_2970,N_2998);
and U3097 (N_3097,N_2912,N_2952);
nor U3098 (N_3098,N_2953,N_2908);
nor U3099 (N_3099,N_2941,N_2957);
nor U3100 (N_3100,N_3068,N_3073);
or U3101 (N_3101,N_3015,N_3026);
nand U3102 (N_3102,N_3057,N_3076);
xor U3103 (N_3103,N_3046,N_3006);
nand U3104 (N_3104,N_3091,N_3053);
nand U3105 (N_3105,N_3047,N_3041);
and U3106 (N_3106,N_3023,N_3094);
nor U3107 (N_3107,N_3084,N_3097);
nor U3108 (N_3108,N_3028,N_3067);
nor U3109 (N_3109,N_3051,N_3010);
xor U3110 (N_3110,N_3048,N_3052);
xor U3111 (N_3111,N_3004,N_3071);
nor U3112 (N_3112,N_3016,N_3056);
and U3113 (N_3113,N_3039,N_3065);
or U3114 (N_3114,N_3096,N_3003);
nand U3115 (N_3115,N_3055,N_3092);
and U3116 (N_3116,N_3095,N_3070);
nand U3117 (N_3117,N_3043,N_3019);
nand U3118 (N_3118,N_3090,N_3099);
nand U3119 (N_3119,N_3042,N_3049);
nor U3120 (N_3120,N_3066,N_3088);
nor U3121 (N_3121,N_3080,N_3093);
nand U3122 (N_3122,N_3029,N_3007);
or U3123 (N_3123,N_3038,N_3098);
nor U3124 (N_3124,N_3075,N_3025);
and U3125 (N_3125,N_3074,N_3013);
nand U3126 (N_3126,N_3058,N_3000);
or U3127 (N_3127,N_3044,N_3086);
nor U3128 (N_3128,N_3005,N_3030);
nand U3129 (N_3129,N_3087,N_3037);
xor U3130 (N_3130,N_3020,N_3033);
nor U3131 (N_3131,N_3014,N_3083);
or U3132 (N_3132,N_3061,N_3011);
and U3133 (N_3133,N_3021,N_3009);
nor U3134 (N_3134,N_3017,N_3034);
or U3135 (N_3135,N_3018,N_3060);
nand U3136 (N_3136,N_3024,N_3085);
nor U3137 (N_3137,N_3077,N_3082);
xnor U3138 (N_3138,N_3063,N_3012);
nor U3139 (N_3139,N_3054,N_3072);
nand U3140 (N_3140,N_3078,N_3064);
xor U3141 (N_3141,N_3069,N_3050);
nand U3142 (N_3142,N_3062,N_3081);
and U3143 (N_3143,N_3036,N_3040);
xor U3144 (N_3144,N_3035,N_3027);
nor U3145 (N_3145,N_3089,N_3008);
and U3146 (N_3146,N_3002,N_3022);
nor U3147 (N_3147,N_3031,N_3001);
and U3148 (N_3148,N_3032,N_3079);
nand U3149 (N_3149,N_3059,N_3045);
and U3150 (N_3150,N_3016,N_3037);
nor U3151 (N_3151,N_3070,N_3085);
or U3152 (N_3152,N_3064,N_3047);
or U3153 (N_3153,N_3071,N_3092);
or U3154 (N_3154,N_3092,N_3060);
nor U3155 (N_3155,N_3037,N_3067);
nand U3156 (N_3156,N_3086,N_3072);
or U3157 (N_3157,N_3023,N_3046);
and U3158 (N_3158,N_3094,N_3036);
and U3159 (N_3159,N_3027,N_3088);
xnor U3160 (N_3160,N_3064,N_3057);
xor U3161 (N_3161,N_3061,N_3077);
nand U3162 (N_3162,N_3049,N_3017);
nand U3163 (N_3163,N_3000,N_3095);
nor U3164 (N_3164,N_3030,N_3014);
nor U3165 (N_3165,N_3092,N_3080);
xnor U3166 (N_3166,N_3027,N_3009);
and U3167 (N_3167,N_3060,N_3078);
and U3168 (N_3168,N_3030,N_3001);
nor U3169 (N_3169,N_3015,N_3043);
xor U3170 (N_3170,N_3085,N_3087);
xor U3171 (N_3171,N_3072,N_3010);
nand U3172 (N_3172,N_3027,N_3048);
nand U3173 (N_3173,N_3022,N_3065);
or U3174 (N_3174,N_3036,N_3071);
xor U3175 (N_3175,N_3069,N_3088);
nor U3176 (N_3176,N_3027,N_3014);
nor U3177 (N_3177,N_3088,N_3034);
nand U3178 (N_3178,N_3087,N_3090);
nor U3179 (N_3179,N_3049,N_3078);
nand U3180 (N_3180,N_3097,N_3057);
and U3181 (N_3181,N_3032,N_3003);
or U3182 (N_3182,N_3072,N_3065);
and U3183 (N_3183,N_3092,N_3097);
and U3184 (N_3184,N_3028,N_3037);
nor U3185 (N_3185,N_3061,N_3099);
and U3186 (N_3186,N_3015,N_3093);
nand U3187 (N_3187,N_3093,N_3017);
and U3188 (N_3188,N_3089,N_3018);
nor U3189 (N_3189,N_3053,N_3082);
nand U3190 (N_3190,N_3059,N_3024);
and U3191 (N_3191,N_3033,N_3028);
or U3192 (N_3192,N_3098,N_3010);
xor U3193 (N_3193,N_3071,N_3079);
or U3194 (N_3194,N_3011,N_3010);
or U3195 (N_3195,N_3023,N_3031);
or U3196 (N_3196,N_3027,N_3068);
and U3197 (N_3197,N_3018,N_3086);
xnor U3198 (N_3198,N_3074,N_3069);
or U3199 (N_3199,N_3003,N_3045);
nor U3200 (N_3200,N_3186,N_3197);
nand U3201 (N_3201,N_3188,N_3125);
nor U3202 (N_3202,N_3102,N_3142);
and U3203 (N_3203,N_3109,N_3179);
xor U3204 (N_3204,N_3135,N_3131);
nor U3205 (N_3205,N_3191,N_3111);
nor U3206 (N_3206,N_3140,N_3136);
nand U3207 (N_3207,N_3161,N_3120);
nand U3208 (N_3208,N_3139,N_3192);
nor U3209 (N_3209,N_3119,N_3194);
and U3210 (N_3210,N_3173,N_3137);
xnor U3211 (N_3211,N_3129,N_3134);
nor U3212 (N_3212,N_3115,N_3175);
or U3213 (N_3213,N_3101,N_3132);
and U3214 (N_3214,N_3177,N_3189);
nor U3215 (N_3215,N_3126,N_3155);
nor U3216 (N_3216,N_3127,N_3116);
nor U3217 (N_3217,N_3150,N_3146);
nand U3218 (N_3218,N_3199,N_3167);
nand U3219 (N_3219,N_3145,N_3178);
or U3220 (N_3220,N_3107,N_3196);
and U3221 (N_3221,N_3187,N_3163);
nand U3222 (N_3222,N_3166,N_3157);
nor U3223 (N_3223,N_3180,N_3112);
and U3224 (N_3224,N_3130,N_3143);
and U3225 (N_3225,N_3160,N_3118);
xnor U3226 (N_3226,N_3162,N_3195);
xor U3227 (N_3227,N_3172,N_3152);
and U3228 (N_3228,N_3122,N_3181);
or U3229 (N_3229,N_3151,N_3138);
or U3230 (N_3230,N_3105,N_3158);
nand U3231 (N_3231,N_3148,N_3176);
nor U3232 (N_3232,N_3170,N_3121);
or U3233 (N_3233,N_3114,N_3153);
nor U3234 (N_3234,N_3156,N_3154);
or U3235 (N_3235,N_3183,N_3124);
or U3236 (N_3236,N_3182,N_3128);
and U3237 (N_3237,N_3104,N_3193);
xnor U3238 (N_3238,N_3108,N_3110);
or U3239 (N_3239,N_3185,N_3165);
xnor U3240 (N_3240,N_3106,N_3149);
nand U3241 (N_3241,N_3198,N_3159);
and U3242 (N_3242,N_3169,N_3184);
or U3243 (N_3243,N_3171,N_3144);
or U3244 (N_3244,N_3141,N_3147);
nor U3245 (N_3245,N_3174,N_3190);
and U3246 (N_3246,N_3103,N_3164);
and U3247 (N_3247,N_3117,N_3123);
or U3248 (N_3248,N_3133,N_3100);
nor U3249 (N_3249,N_3168,N_3113);
or U3250 (N_3250,N_3127,N_3113);
nor U3251 (N_3251,N_3126,N_3182);
or U3252 (N_3252,N_3185,N_3105);
or U3253 (N_3253,N_3129,N_3157);
and U3254 (N_3254,N_3113,N_3133);
or U3255 (N_3255,N_3163,N_3191);
or U3256 (N_3256,N_3168,N_3126);
nand U3257 (N_3257,N_3127,N_3111);
and U3258 (N_3258,N_3165,N_3135);
and U3259 (N_3259,N_3198,N_3121);
or U3260 (N_3260,N_3192,N_3100);
and U3261 (N_3261,N_3156,N_3186);
nand U3262 (N_3262,N_3103,N_3180);
nor U3263 (N_3263,N_3125,N_3149);
xor U3264 (N_3264,N_3187,N_3189);
nor U3265 (N_3265,N_3106,N_3184);
or U3266 (N_3266,N_3189,N_3199);
and U3267 (N_3267,N_3183,N_3153);
nand U3268 (N_3268,N_3188,N_3149);
nor U3269 (N_3269,N_3163,N_3166);
xor U3270 (N_3270,N_3166,N_3126);
nor U3271 (N_3271,N_3185,N_3127);
nand U3272 (N_3272,N_3122,N_3148);
and U3273 (N_3273,N_3162,N_3145);
nand U3274 (N_3274,N_3182,N_3157);
nand U3275 (N_3275,N_3127,N_3135);
or U3276 (N_3276,N_3107,N_3163);
nor U3277 (N_3277,N_3157,N_3122);
nor U3278 (N_3278,N_3121,N_3153);
nand U3279 (N_3279,N_3107,N_3177);
or U3280 (N_3280,N_3165,N_3169);
and U3281 (N_3281,N_3171,N_3199);
or U3282 (N_3282,N_3159,N_3110);
nor U3283 (N_3283,N_3177,N_3198);
or U3284 (N_3284,N_3163,N_3129);
xnor U3285 (N_3285,N_3154,N_3115);
nand U3286 (N_3286,N_3126,N_3174);
xnor U3287 (N_3287,N_3144,N_3101);
and U3288 (N_3288,N_3154,N_3147);
or U3289 (N_3289,N_3109,N_3102);
nand U3290 (N_3290,N_3174,N_3163);
xor U3291 (N_3291,N_3137,N_3109);
and U3292 (N_3292,N_3197,N_3176);
and U3293 (N_3293,N_3153,N_3135);
and U3294 (N_3294,N_3172,N_3137);
or U3295 (N_3295,N_3155,N_3148);
nor U3296 (N_3296,N_3131,N_3100);
and U3297 (N_3297,N_3113,N_3181);
nor U3298 (N_3298,N_3144,N_3174);
or U3299 (N_3299,N_3126,N_3133);
nor U3300 (N_3300,N_3263,N_3248);
nor U3301 (N_3301,N_3206,N_3275);
nand U3302 (N_3302,N_3294,N_3246);
or U3303 (N_3303,N_3220,N_3219);
or U3304 (N_3304,N_3288,N_3241);
nand U3305 (N_3305,N_3266,N_3287);
nand U3306 (N_3306,N_3222,N_3298);
nor U3307 (N_3307,N_3283,N_3236);
and U3308 (N_3308,N_3281,N_3284);
nand U3309 (N_3309,N_3285,N_3289);
nor U3310 (N_3310,N_3271,N_3218);
and U3311 (N_3311,N_3226,N_3257);
or U3312 (N_3312,N_3253,N_3221);
nor U3313 (N_3313,N_3274,N_3244);
xor U3314 (N_3314,N_3227,N_3205);
nand U3315 (N_3315,N_3209,N_3292);
nor U3316 (N_3316,N_3265,N_3297);
or U3317 (N_3317,N_3213,N_3237);
xor U3318 (N_3318,N_3242,N_3223);
nor U3319 (N_3319,N_3217,N_3295);
nand U3320 (N_3320,N_3207,N_3239);
and U3321 (N_3321,N_3280,N_3278);
or U3322 (N_3322,N_3291,N_3234);
nand U3323 (N_3323,N_3210,N_3270);
nor U3324 (N_3324,N_3240,N_3211);
or U3325 (N_3325,N_3228,N_3250);
and U3326 (N_3326,N_3215,N_3268);
or U3327 (N_3327,N_3261,N_3224);
or U3328 (N_3328,N_3277,N_3200);
or U3329 (N_3329,N_3296,N_3290);
nand U3330 (N_3330,N_3230,N_3243);
nand U3331 (N_3331,N_3229,N_3212);
xor U3332 (N_3332,N_3255,N_3225);
or U3333 (N_3333,N_3272,N_3276);
xnor U3334 (N_3334,N_3249,N_3201);
xnor U3335 (N_3335,N_3231,N_3203);
nor U3336 (N_3336,N_3299,N_3258);
nand U3337 (N_3337,N_3235,N_3204);
nor U3338 (N_3338,N_3286,N_3202);
nor U3339 (N_3339,N_3293,N_3214);
or U3340 (N_3340,N_3282,N_3262);
nor U3341 (N_3341,N_3232,N_3208);
nand U3342 (N_3342,N_3245,N_3267);
and U3343 (N_3343,N_3216,N_3252);
nand U3344 (N_3344,N_3233,N_3238);
or U3345 (N_3345,N_3269,N_3279);
nor U3346 (N_3346,N_3259,N_3256);
nand U3347 (N_3347,N_3247,N_3251);
and U3348 (N_3348,N_3264,N_3260);
nor U3349 (N_3349,N_3254,N_3273);
nand U3350 (N_3350,N_3217,N_3229);
xnor U3351 (N_3351,N_3235,N_3260);
nand U3352 (N_3352,N_3261,N_3272);
and U3353 (N_3353,N_3221,N_3284);
and U3354 (N_3354,N_3286,N_3271);
nor U3355 (N_3355,N_3248,N_3219);
nand U3356 (N_3356,N_3258,N_3293);
and U3357 (N_3357,N_3263,N_3252);
xnor U3358 (N_3358,N_3240,N_3239);
and U3359 (N_3359,N_3211,N_3212);
or U3360 (N_3360,N_3270,N_3243);
or U3361 (N_3361,N_3255,N_3200);
nand U3362 (N_3362,N_3271,N_3212);
xnor U3363 (N_3363,N_3206,N_3223);
or U3364 (N_3364,N_3278,N_3235);
and U3365 (N_3365,N_3287,N_3275);
and U3366 (N_3366,N_3250,N_3220);
or U3367 (N_3367,N_3274,N_3262);
nand U3368 (N_3368,N_3209,N_3275);
and U3369 (N_3369,N_3257,N_3270);
and U3370 (N_3370,N_3245,N_3251);
or U3371 (N_3371,N_3210,N_3282);
or U3372 (N_3372,N_3269,N_3266);
nand U3373 (N_3373,N_3245,N_3299);
nor U3374 (N_3374,N_3213,N_3210);
or U3375 (N_3375,N_3290,N_3253);
nor U3376 (N_3376,N_3285,N_3245);
nor U3377 (N_3377,N_3218,N_3259);
nand U3378 (N_3378,N_3211,N_3200);
nor U3379 (N_3379,N_3237,N_3289);
and U3380 (N_3380,N_3220,N_3272);
nand U3381 (N_3381,N_3257,N_3205);
nor U3382 (N_3382,N_3238,N_3247);
nor U3383 (N_3383,N_3256,N_3204);
and U3384 (N_3384,N_3230,N_3292);
and U3385 (N_3385,N_3257,N_3227);
and U3386 (N_3386,N_3203,N_3238);
or U3387 (N_3387,N_3248,N_3242);
or U3388 (N_3388,N_3210,N_3249);
nor U3389 (N_3389,N_3284,N_3217);
and U3390 (N_3390,N_3202,N_3276);
xor U3391 (N_3391,N_3299,N_3213);
and U3392 (N_3392,N_3272,N_3279);
and U3393 (N_3393,N_3205,N_3221);
and U3394 (N_3394,N_3239,N_3216);
xnor U3395 (N_3395,N_3232,N_3229);
and U3396 (N_3396,N_3237,N_3211);
nor U3397 (N_3397,N_3292,N_3278);
and U3398 (N_3398,N_3269,N_3250);
nand U3399 (N_3399,N_3222,N_3283);
and U3400 (N_3400,N_3387,N_3388);
or U3401 (N_3401,N_3382,N_3342);
nor U3402 (N_3402,N_3384,N_3395);
nand U3403 (N_3403,N_3392,N_3319);
or U3404 (N_3404,N_3343,N_3310);
xnor U3405 (N_3405,N_3352,N_3341);
and U3406 (N_3406,N_3348,N_3327);
nand U3407 (N_3407,N_3316,N_3377);
nor U3408 (N_3408,N_3338,N_3366);
or U3409 (N_3409,N_3361,N_3360);
nor U3410 (N_3410,N_3340,N_3325);
nand U3411 (N_3411,N_3302,N_3336);
nand U3412 (N_3412,N_3380,N_3337);
xnor U3413 (N_3413,N_3381,N_3356);
nand U3414 (N_3414,N_3371,N_3318);
or U3415 (N_3415,N_3303,N_3376);
nor U3416 (N_3416,N_3332,N_3367);
nand U3417 (N_3417,N_3312,N_3359);
nand U3418 (N_3418,N_3347,N_3315);
nor U3419 (N_3419,N_3368,N_3331);
and U3420 (N_3420,N_3357,N_3301);
xor U3421 (N_3421,N_3358,N_3345);
nor U3422 (N_3422,N_3349,N_3326);
nor U3423 (N_3423,N_3363,N_3393);
nor U3424 (N_3424,N_3394,N_3346);
nor U3425 (N_3425,N_3353,N_3314);
or U3426 (N_3426,N_3375,N_3391);
and U3427 (N_3427,N_3379,N_3320);
or U3428 (N_3428,N_3397,N_3365);
and U3429 (N_3429,N_3323,N_3350);
or U3430 (N_3430,N_3396,N_3311);
nor U3431 (N_3431,N_3399,N_3383);
nor U3432 (N_3432,N_3306,N_3344);
nor U3433 (N_3433,N_3378,N_3369);
nand U3434 (N_3434,N_3304,N_3390);
or U3435 (N_3435,N_3333,N_3385);
and U3436 (N_3436,N_3322,N_3307);
nor U3437 (N_3437,N_3374,N_3389);
xor U3438 (N_3438,N_3370,N_3305);
nand U3439 (N_3439,N_3300,N_3354);
nor U3440 (N_3440,N_3351,N_3324);
nand U3441 (N_3441,N_3328,N_3355);
nand U3442 (N_3442,N_3339,N_3398);
and U3443 (N_3443,N_3317,N_3335);
or U3444 (N_3444,N_3364,N_3309);
nand U3445 (N_3445,N_3321,N_3308);
and U3446 (N_3446,N_3334,N_3386);
nand U3447 (N_3447,N_3313,N_3362);
nor U3448 (N_3448,N_3329,N_3372);
or U3449 (N_3449,N_3373,N_3330);
or U3450 (N_3450,N_3349,N_3330);
xor U3451 (N_3451,N_3335,N_3336);
xnor U3452 (N_3452,N_3358,N_3366);
and U3453 (N_3453,N_3369,N_3368);
xnor U3454 (N_3454,N_3319,N_3378);
or U3455 (N_3455,N_3313,N_3375);
nand U3456 (N_3456,N_3330,N_3370);
nand U3457 (N_3457,N_3375,N_3363);
and U3458 (N_3458,N_3303,N_3365);
nand U3459 (N_3459,N_3338,N_3319);
nand U3460 (N_3460,N_3371,N_3389);
nand U3461 (N_3461,N_3360,N_3392);
or U3462 (N_3462,N_3327,N_3375);
or U3463 (N_3463,N_3337,N_3324);
nand U3464 (N_3464,N_3312,N_3345);
and U3465 (N_3465,N_3399,N_3321);
and U3466 (N_3466,N_3323,N_3302);
or U3467 (N_3467,N_3330,N_3332);
nand U3468 (N_3468,N_3323,N_3336);
nand U3469 (N_3469,N_3393,N_3374);
and U3470 (N_3470,N_3341,N_3317);
nor U3471 (N_3471,N_3317,N_3325);
and U3472 (N_3472,N_3375,N_3371);
or U3473 (N_3473,N_3363,N_3311);
and U3474 (N_3474,N_3308,N_3384);
or U3475 (N_3475,N_3399,N_3360);
nor U3476 (N_3476,N_3334,N_3346);
nor U3477 (N_3477,N_3364,N_3344);
and U3478 (N_3478,N_3373,N_3386);
nor U3479 (N_3479,N_3385,N_3314);
and U3480 (N_3480,N_3307,N_3386);
nand U3481 (N_3481,N_3301,N_3315);
nand U3482 (N_3482,N_3391,N_3370);
nor U3483 (N_3483,N_3368,N_3315);
nor U3484 (N_3484,N_3302,N_3327);
or U3485 (N_3485,N_3301,N_3362);
nand U3486 (N_3486,N_3374,N_3334);
or U3487 (N_3487,N_3381,N_3317);
nand U3488 (N_3488,N_3340,N_3386);
or U3489 (N_3489,N_3312,N_3379);
or U3490 (N_3490,N_3352,N_3350);
nor U3491 (N_3491,N_3328,N_3314);
or U3492 (N_3492,N_3371,N_3316);
or U3493 (N_3493,N_3320,N_3310);
nand U3494 (N_3494,N_3337,N_3391);
and U3495 (N_3495,N_3313,N_3374);
xor U3496 (N_3496,N_3367,N_3375);
nand U3497 (N_3497,N_3317,N_3399);
nor U3498 (N_3498,N_3350,N_3322);
or U3499 (N_3499,N_3391,N_3344);
or U3500 (N_3500,N_3400,N_3445);
nand U3501 (N_3501,N_3497,N_3441);
and U3502 (N_3502,N_3472,N_3428);
nor U3503 (N_3503,N_3415,N_3463);
and U3504 (N_3504,N_3466,N_3443);
nor U3505 (N_3505,N_3495,N_3419);
and U3506 (N_3506,N_3496,N_3455);
nand U3507 (N_3507,N_3491,N_3407);
nor U3508 (N_3508,N_3431,N_3411);
nand U3509 (N_3509,N_3406,N_3462);
nand U3510 (N_3510,N_3489,N_3486);
xnor U3511 (N_3511,N_3460,N_3482);
and U3512 (N_3512,N_3464,N_3468);
nand U3513 (N_3513,N_3401,N_3457);
or U3514 (N_3514,N_3454,N_3417);
or U3515 (N_3515,N_3448,N_3418);
and U3516 (N_3516,N_3442,N_3447);
and U3517 (N_3517,N_3453,N_3424);
and U3518 (N_3518,N_3476,N_3426);
xor U3519 (N_3519,N_3429,N_3446);
nor U3520 (N_3520,N_3433,N_3402);
xor U3521 (N_3521,N_3469,N_3475);
nand U3522 (N_3522,N_3409,N_3492);
and U3523 (N_3523,N_3473,N_3410);
xor U3524 (N_3524,N_3434,N_3456);
and U3525 (N_3525,N_3499,N_3459);
and U3526 (N_3526,N_3437,N_3405);
and U3527 (N_3527,N_3450,N_3404);
nand U3528 (N_3528,N_3449,N_3471);
or U3529 (N_3529,N_3440,N_3465);
nor U3530 (N_3530,N_3412,N_3451);
and U3531 (N_3531,N_3481,N_3485);
nor U3532 (N_3532,N_3444,N_3474);
or U3533 (N_3533,N_3427,N_3480);
and U3534 (N_3534,N_3467,N_3435);
nand U3535 (N_3535,N_3436,N_3477);
xor U3536 (N_3536,N_3425,N_3461);
and U3537 (N_3537,N_3421,N_3416);
or U3538 (N_3538,N_3408,N_3430);
or U3539 (N_3539,N_3438,N_3423);
nand U3540 (N_3540,N_3414,N_3432);
nor U3541 (N_3541,N_3494,N_3420);
nor U3542 (N_3542,N_3479,N_3493);
or U3543 (N_3543,N_3403,N_3413);
nand U3544 (N_3544,N_3484,N_3478);
or U3545 (N_3545,N_3487,N_3458);
nand U3546 (N_3546,N_3452,N_3470);
nand U3547 (N_3547,N_3490,N_3422);
nand U3548 (N_3548,N_3439,N_3498);
and U3549 (N_3549,N_3488,N_3483);
xor U3550 (N_3550,N_3415,N_3499);
or U3551 (N_3551,N_3473,N_3471);
or U3552 (N_3552,N_3416,N_3429);
and U3553 (N_3553,N_3497,N_3419);
or U3554 (N_3554,N_3481,N_3498);
nor U3555 (N_3555,N_3439,N_3479);
xnor U3556 (N_3556,N_3459,N_3482);
nor U3557 (N_3557,N_3481,N_3457);
and U3558 (N_3558,N_3428,N_3474);
xor U3559 (N_3559,N_3439,N_3445);
nand U3560 (N_3560,N_3492,N_3486);
nand U3561 (N_3561,N_3498,N_3455);
or U3562 (N_3562,N_3423,N_3497);
or U3563 (N_3563,N_3499,N_3414);
nor U3564 (N_3564,N_3405,N_3409);
nor U3565 (N_3565,N_3400,N_3458);
nand U3566 (N_3566,N_3444,N_3407);
or U3567 (N_3567,N_3455,N_3430);
nand U3568 (N_3568,N_3489,N_3408);
and U3569 (N_3569,N_3493,N_3422);
and U3570 (N_3570,N_3492,N_3484);
nand U3571 (N_3571,N_3471,N_3479);
and U3572 (N_3572,N_3443,N_3464);
nand U3573 (N_3573,N_3456,N_3428);
nand U3574 (N_3574,N_3452,N_3463);
nand U3575 (N_3575,N_3499,N_3433);
nor U3576 (N_3576,N_3400,N_3433);
and U3577 (N_3577,N_3421,N_3424);
or U3578 (N_3578,N_3495,N_3467);
and U3579 (N_3579,N_3472,N_3466);
nand U3580 (N_3580,N_3487,N_3462);
or U3581 (N_3581,N_3410,N_3408);
nand U3582 (N_3582,N_3450,N_3493);
or U3583 (N_3583,N_3464,N_3414);
xnor U3584 (N_3584,N_3437,N_3481);
nor U3585 (N_3585,N_3496,N_3408);
nor U3586 (N_3586,N_3410,N_3470);
nand U3587 (N_3587,N_3425,N_3434);
nand U3588 (N_3588,N_3444,N_3440);
nand U3589 (N_3589,N_3487,N_3402);
or U3590 (N_3590,N_3426,N_3497);
xor U3591 (N_3591,N_3478,N_3498);
and U3592 (N_3592,N_3432,N_3491);
nor U3593 (N_3593,N_3451,N_3485);
nor U3594 (N_3594,N_3435,N_3489);
or U3595 (N_3595,N_3472,N_3483);
nor U3596 (N_3596,N_3477,N_3478);
or U3597 (N_3597,N_3422,N_3407);
nand U3598 (N_3598,N_3476,N_3480);
or U3599 (N_3599,N_3445,N_3431);
nand U3600 (N_3600,N_3594,N_3505);
or U3601 (N_3601,N_3579,N_3597);
nand U3602 (N_3602,N_3502,N_3578);
nor U3603 (N_3603,N_3559,N_3537);
and U3604 (N_3604,N_3573,N_3501);
and U3605 (N_3605,N_3533,N_3527);
nand U3606 (N_3606,N_3581,N_3596);
nand U3607 (N_3607,N_3561,N_3550);
and U3608 (N_3608,N_3562,N_3558);
xnor U3609 (N_3609,N_3515,N_3521);
nand U3610 (N_3610,N_3507,N_3514);
or U3611 (N_3611,N_3593,N_3590);
or U3612 (N_3612,N_3531,N_3524);
xnor U3613 (N_3613,N_3511,N_3570);
or U3614 (N_3614,N_3568,N_3555);
nor U3615 (N_3615,N_3523,N_3571);
and U3616 (N_3616,N_3532,N_3545);
nor U3617 (N_3617,N_3565,N_3574);
nor U3618 (N_3618,N_3512,N_3504);
nor U3619 (N_3619,N_3569,N_3583);
or U3620 (N_3620,N_3575,N_3572);
nand U3621 (N_3621,N_3547,N_3584);
nand U3622 (N_3622,N_3548,N_3522);
xnor U3623 (N_3623,N_3539,N_3503);
or U3624 (N_3624,N_3566,N_3589);
and U3625 (N_3625,N_3557,N_3599);
and U3626 (N_3626,N_3517,N_3543);
nor U3627 (N_3627,N_3595,N_3509);
and U3628 (N_3628,N_3567,N_3506);
nor U3629 (N_3629,N_3549,N_3551);
or U3630 (N_3630,N_3554,N_3534);
or U3631 (N_3631,N_3544,N_3510);
or U3632 (N_3632,N_3564,N_3528);
nor U3633 (N_3633,N_3582,N_3529);
nand U3634 (N_3634,N_3513,N_3538);
nor U3635 (N_3635,N_3576,N_3592);
and U3636 (N_3636,N_3546,N_3560);
and U3637 (N_3637,N_3535,N_3552);
nand U3638 (N_3638,N_3525,N_3541);
or U3639 (N_3639,N_3530,N_3508);
and U3640 (N_3640,N_3542,N_3588);
xnor U3641 (N_3641,N_3536,N_3520);
or U3642 (N_3642,N_3585,N_3563);
and U3643 (N_3643,N_3516,N_3598);
nor U3644 (N_3644,N_3577,N_3519);
nor U3645 (N_3645,N_3518,N_3553);
nor U3646 (N_3646,N_3591,N_3556);
nor U3647 (N_3647,N_3540,N_3586);
nand U3648 (N_3648,N_3526,N_3500);
and U3649 (N_3649,N_3587,N_3580);
nand U3650 (N_3650,N_3565,N_3560);
and U3651 (N_3651,N_3516,N_3570);
nand U3652 (N_3652,N_3590,N_3554);
nand U3653 (N_3653,N_3510,N_3547);
and U3654 (N_3654,N_3561,N_3582);
or U3655 (N_3655,N_3560,N_3513);
and U3656 (N_3656,N_3526,N_3543);
nor U3657 (N_3657,N_3522,N_3502);
and U3658 (N_3658,N_3533,N_3524);
or U3659 (N_3659,N_3545,N_3562);
nor U3660 (N_3660,N_3599,N_3550);
nor U3661 (N_3661,N_3580,N_3568);
nand U3662 (N_3662,N_3555,N_3535);
or U3663 (N_3663,N_3544,N_3571);
and U3664 (N_3664,N_3556,N_3553);
nor U3665 (N_3665,N_3598,N_3553);
xor U3666 (N_3666,N_3502,N_3535);
nand U3667 (N_3667,N_3538,N_3574);
nor U3668 (N_3668,N_3562,N_3503);
or U3669 (N_3669,N_3519,N_3563);
xnor U3670 (N_3670,N_3505,N_3571);
nor U3671 (N_3671,N_3523,N_3592);
and U3672 (N_3672,N_3549,N_3534);
and U3673 (N_3673,N_3539,N_3574);
nand U3674 (N_3674,N_3528,N_3504);
and U3675 (N_3675,N_3554,N_3535);
nor U3676 (N_3676,N_3555,N_3530);
nor U3677 (N_3677,N_3556,N_3596);
xor U3678 (N_3678,N_3507,N_3524);
nor U3679 (N_3679,N_3593,N_3586);
xor U3680 (N_3680,N_3541,N_3592);
nor U3681 (N_3681,N_3552,N_3512);
and U3682 (N_3682,N_3548,N_3520);
and U3683 (N_3683,N_3556,N_3546);
or U3684 (N_3684,N_3548,N_3583);
nor U3685 (N_3685,N_3543,N_3587);
nor U3686 (N_3686,N_3578,N_3575);
nor U3687 (N_3687,N_3573,N_3555);
and U3688 (N_3688,N_3531,N_3578);
nand U3689 (N_3689,N_3576,N_3577);
or U3690 (N_3690,N_3583,N_3586);
nor U3691 (N_3691,N_3575,N_3508);
nand U3692 (N_3692,N_3575,N_3558);
nor U3693 (N_3693,N_3591,N_3521);
or U3694 (N_3694,N_3578,N_3538);
nor U3695 (N_3695,N_3561,N_3503);
xor U3696 (N_3696,N_3569,N_3519);
nor U3697 (N_3697,N_3579,N_3530);
nand U3698 (N_3698,N_3517,N_3520);
nor U3699 (N_3699,N_3594,N_3543);
nor U3700 (N_3700,N_3674,N_3608);
nor U3701 (N_3701,N_3678,N_3684);
nor U3702 (N_3702,N_3676,N_3600);
and U3703 (N_3703,N_3644,N_3647);
nor U3704 (N_3704,N_3628,N_3603);
and U3705 (N_3705,N_3623,N_3605);
or U3706 (N_3706,N_3669,N_3653);
nand U3707 (N_3707,N_3680,N_3624);
or U3708 (N_3708,N_3643,N_3677);
and U3709 (N_3709,N_3689,N_3612);
or U3710 (N_3710,N_3662,N_3640);
nor U3711 (N_3711,N_3655,N_3637);
and U3712 (N_3712,N_3666,N_3616);
and U3713 (N_3713,N_3607,N_3671);
and U3714 (N_3714,N_3692,N_3694);
nand U3715 (N_3715,N_3675,N_3697);
nand U3716 (N_3716,N_3696,N_3615);
and U3717 (N_3717,N_3688,N_3681);
and U3718 (N_3718,N_3652,N_3633);
nor U3719 (N_3719,N_3611,N_3650);
nor U3720 (N_3720,N_3610,N_3642);
and U3721 (N_3721,N_3619,N_3632);
nand U3722 (N_3722,N_3654,N_3651);
and U3723 (N_3723,N_3686,N_3679);
and U3724 (N_3724,N_3609,N_3687);
or U3725 (N_3725,N_3645,N_3602);
or U3726 (N_3726,N_3672,N_3614);
and U3727 (N_3727,N_3639,N_3690);
and U3728 (N_3728,N_3630,N_3636);
and U3729 (N_3729,N_3661,N_3604);
nand U3730 (N_3730,N_3665,N_3646);
xor U3731 (N_3731,N_3685,N_3691);
or U3732 (N_3732,N_3668,N_3613);
xnor U3733 (N_3733,N_3626,N_3618);
nor U3734 (N_3734,N_3648,N_3670);
nand U3735 (N_3735,N_3658,N_3683);
and U3736 (N_3736,N_3638,N_3693);
and U3737 (N_3737,N_3629,N_3627);
or U3738 (N_3738,N_3635,N_3660);
or U3739 (N_3739,N_3601,N_3606);
nand U3740 (N_3740,N_3634,N_3663);
xnor U3741 (N_3741,N_3673,N_3649);
nand U3742 (N_3742,N_3617,N_3620);
nor U3743 (N_3743,N_3631,N_3625);
or U3744 (N_3744,N_3656,N_3641);
or U3745 (N_3745,N_3659,N_3657);
nor U3746 (N_3746,N_3695,N_3698);
or U3747 (N_3747,N_3664,N_3622);
or U3748 (N_3748,N_3682,N_3621);
and U3749 (N_3749,N_3699,N_3667);
nand U3750 (N_3750,N_3657,N_3647);
and U3751 (N_3751,N_3632,N_3686);
nor U3752 (N_3752,N_3681,N_3685);
nand U3753 (N_3753,N_3638,N_3625);
and U3754 (N_3754,N_3626,N_3644);
nand U3755 (N_3755,N_3662,N_3612);
and U3756 (N_3756,N_3605,N_3644);
nand U3757 (N_3757,N_3624,N_3688);
or U3758 (N_3758,N_3661,N_3633);
or U3759 (N_3759,N_3698,N_3683);
and U3760 (N_3760,N_3674,N_3691);
xnor U3761 (N_3761,N_3665,N_3638);
and U3762 (N_3762,N_3663,N_3694);
and U3763 (N_3763,N_3603,N_3685);
and U3764 (N_3764,N_3692,N_3607);
and U3765 (N_3765,N_3680,N_3633);
xor U3766 (N_3766,N_3673,N_3650);
and U3767 (N_3767,N_3626,N_3684);
nand U3768 (N_3768,N_3650,N_3613);
nand U3769 (N_3769,N_3684,N_3681);
nor U3770 (N_3770,N_3666,N_3659);
nand U3771 (N_3771,N_3646,N_3699);
and U3772 (N_3772,N_3621,N_3604);
and U3773 (N_3773,N_3623,N_3608);
nor U3774 (N_3774,N_3648,N_3664);
nor U3775 (N_3775,N_3650,N_3680);
or U3776 (N_3776,N_3690,N_3695);
or U3777 (N_3777,N_3675,N_3672);
nand U3778 (N_3778,N_3665,N_3676);
nor U3779 (N_3779,N_3652,N_3635);
or U3780 (N_3780,N_3620,N_3630);
nand U3781 (N_3781,N_3633,N_3618);
xnor U3782 (N_3782,N_3672,N_3616);
nand U3783 (N_3783,N_3681,N_3601);
nor U3784 (N_3784,N_3688,N_3692);
or U3785 (N_3785,N_3686,N_3657);
nor U3786 (N_3786,N_3635,N_3686);
and U3787 (N_3787,N_3644,N_3697);
xnor U3788 (N_3788,N_3696,N_3657);
or U3789 (N_3789,N_3672,N_3607);
xor U3790 (N_3790,N_3655,N_3617);
nor U3791 (N_3791,N_3665,N_3642);
or U3792 (N_3792,N_3613,N_3624);
xor U3793 (N_3793,N_3656,N_3690);
and U3794 (N_3794,N_3680,N_3679);
nor U3795 (N_3795,N_3636,N_3607);
and U3796 (N_3796,N_3655,N_3682);
nor U3797 (N_3797,N_3601,N_3683);
or U3798 (N_3798,N_3676,N_3686);
nor U3799 (N_3799,N_3609,N_3606);
nand U3800 (N_3800,N_3798,N_3754);
nand U3801 (N_3801,N_3713,N_3740);
or U3802 (N_3802,N_3718,N_3717);
and U3803 (N_3803,N_3728,N_3712);
nor U3804 (N_3804,N_3719,N_3720);
nand U3805 (N_3805,N_3741,N_3775);
nor U3806 (N_3806,N_3770,N_3766);
and U3807 (N_3807,N_3753,N_3746);
and U3808 (N_3808,N_3776,N_3771);
or U3809 (N_3809,N_3793,N_3796);
nor U3810 (N_3810,N_3777,N_3739);
nor U3811 (N_3811,N_3706,N_3714);
or U3812 (N_3812,N_3769,N_3723);
and U3813 (N_3813,N_3725,N_3787);
nand U3814 (N_3814,N_3780,N_3797);
xnor U3815 (N_3815,N_3778,N_3722);
and U3816 (N_3816,N_3760,N_3734);
nor U3817 (N_3817,N_3784,N_3715);
or U3818 (N_3818,N_3711,N_3773);
nand U3819 (N_3819,N_3705,N_3721);
nor U3820 (N_3820,N_3745,N_3789);
or U3821 (N_3821,N_3765,N_3786);
or U3822 (N_3822,N_3772,N_3733);
nor U3823 (N_3823,N_3737,N_3757);
xor U3824 (N_3824,N_3779,N_3788);
or U3825 (N_3825,N_3792,N_3747);
nor U3826 (N_3826,N_3729,N_3716);
and U3827 (N_3827,N_3752,N_3761);
and U3828 (N_3828,N_3700,N_3742);
and U3829 (N_3829,N_3799,N_3781);
xnor U3830 (N_3830,N_3744,N_3709);
and U3831 (N_3831,N_3710,N_3762);
and U3832 (N_3832,N_3732,N_3791);
nand U3833 (N_3833,N_3748,N_3701);
nor U3834 (N_3834,N_3703,N_3727);
and U3835 (N_3835,N_3708,N_3795);
xor U3836 (N_3836,N_3743,N_3749);
nand U3837 (N_3837,N_3738,N_3751);
nand U3838 (N_3838,N_3768,N_3782);
nor U3839 (N_3839,N_3767,N_3736);
xor U3840 (N_3840,N_3763,N_3774);
or U3841 (N_3841,N_3794,N_3724);
nor U3842 (N_3842,N_3730,N_3758);
nand U3843 (N_3843,N_3759,N_3750);
nand U3844 (N_3844,N_3764,N_3704);
nor U3845 (N_3845,N_3726,N_3756);
xor U3846 (N_3846,N_3707,N_3783);
or U3847 (N_3847,N_3731,N_3785);
nor U3848 (N_3848,N_3755,N_3790);
or U3849 (N_3849,N_3702,N_3735);
and U3850 (N_3850,N_3753,N_3709);
nand U3851 (N_3851,N_3728,N_3729);
and U3852 (N_3852,N_3765,N_3762);
and U3853 (N_3853,N_3776,N_3725);
and U3854 (N_3854,N_3731,N_3776);
xor U3855 (N_3855,N_3716,N_3750);
nor U3856 (N_3856,N_3704,N_3781);
and U3857 (N_3857,N_3751,N_3701);
nand U3858 (N_3858,N_3728,N_3723);
and U3859 (N_3859,N_3705,N_3731);
and U3860 (N_3860,N_3745,N_3700);
nor U3861 (N_3861,N_3756,N_3787);
and U3862 (N_3862,N_3760,N_3736);
xnor U3863 (N_3863,N_3781,N_3770);
and U3864 (N_3864,N_3758,N_3753);
or U3865 (N_3865,N_3755,N_3738);
xor U3866 (N_3866,N_3765,N_3737);
or U3867 (N_3867,N_3742,N_3728);
nor U3868 (N_3868,N_3727,N_3775);
nand U3869 (N_3869,N_3717,N_3743);
nor U3870 (N_3870,N_3734,N_3711);
nor U3871 (N_3871,N_3700,N_3720);
or U3872 (N_3872,N_3754,N_3728);
nand U3873 (N_3873,N_3718,N_3709);
nand U3874 (N_3874,N_3763,N_3728);
xnor U3875 (N_3875,N_3730,N_3741);
xor U3876 (N_3876,N_3770,N_3785);
nand U3877 (N_3877,N_3724,N_3722);
nand U3878 (N_3878,N_3780,N_3772);
and U3879 (N_3879,N_3709,N_3785);
and U3880 (N_3880,N_3783,N_3701);
xnor U3881 (N_3881,N_3705,N_3708);
nand U3882 (N_3882,N_3778,N_3725);
and U3883 (N_3883,N_3765,N_3752);
nor U3884 (N_3884,N_3728,N_3778);
xnor U3885 (N_3885,N_3780,N_3738);
and U3886 (N_3886,N_3702,N_3767);
nand U3887 (N_3887,N_3700,N_3771);
and U3888 (N_3888,N_3706,N_3795);
nor U3889 (N_3889,N_3733,N_3740);
and U3890 (N_3890,N_3710,N_3794);
and U3891 (N_3891,N_3781,N_3765);
or U3892 (N_3892,N_3710,N_3751);
or U3893 (N_3893,N_3736,N_3701);
and U3894 (N_3894,N_3763,N_3735);
or U3895 (N_3895,N_3718,N_3784);
xnor U3896 (N_3896,N_3796,N_3769);
and U3897 (N_3897,N_3750,N_3729);
or U3898 (N_3898,N_3777,N_3737);
nor U3899 (N_3899,N_3786,N_3735);
and U3900 (N_3900,N_3805,N_3879);
xnor U3901 (N_3901,N_3896,N_3889);
nand U3902 (N_3902,N_3855,N_3899);
nor U3903 (N_3903,N_3863,N_3822);
or U3904 (N_3904,N_3867,N_3825);
nor U3905 (N_3905,N_3824,N_3866);
xnor U3906 (N_3906,N_3830,N_3852);
or U3907 (N_3907,N_3850,N_3878);
nand U3908 (N_3908,N_3884,N_3885);
or U3909 (N_3909,N_3864,N_3833);
nand U3910 (N_3910,N_3897,N_3860);
nand U3911 (N_3911,N_3875,N_3894);
nand U3912 (N_3912,N_3826,N_3876);
nand U3913 (N_3913,N_3810,N_3893);
nand U3914 (N_3914,N_3883,N_3851);
nor U3915 (N_3915,N_3848,N_3816);
or U3916 (N_3916,N_3853,N_3869);
nand U3917 (N_3917,N_3871,N_3831);
nand U3918 (N_3918,N_3837,N_3812);
nor U3919 (N_3919,N_3817,N_3820);
nor U3920 (N_3920,N_3807,N_3815);
xnor U3921 (N_3921,N_3841,N_3880);
nand U3922 (N_3922,N_3877,N_3814);
xnor U3923 (N_3923,N_3874,N_3865);
xor U3924 (N_3924,N_3846,N_3828);
or U3925 (N_3925,N_3827,N_3888);
and U3926 (N_3926,N_3829,N_3802);
and U3927 (N_3927,N_3887,N_3823);
or U3928 (N_3928,N_3806,N_3845);
and U3929 (N_3929,N_3834,N_3859);
nor U3930 (N_3930,N_3857,N_3838);
or U3931 (N_3931,N_3882,N_3804);
and U3932 (N_3932,N_3842,N_3836);
and U3933 (N_3933,N_3800,N_3818);
xor U3934 (N_3934,N_3868,N_3821);
or U3935 (N_3935,N_3861,N_3843);
xnor U3936 (N_3936,N_3811,N_3849);
or U3937 (N_3937,N_3844,N_3891);
and U3938 (N_3938,N_3892,N_3839);
and U3939 (N_3939,N_3832,N_3856);
nand U3940 (N_3940,N_3840,N_3858);
or U3941 (N_3941,N_3809,N_3847);
and U3942 (N_3942,N_3895,N_3813);
and U3943 (N_3943,N_3801,N_3808);
and U3944 (N_3944,N_3870,N_3890);
xor U3945 (N_3945,N_3835,N_3854);
nand U3946 (N_3946,N_3886,N_3803);
nor U3947 (N_3947,N_3881,N_3898);
and U3948 (N_3948,N_3872,N_3873);
xor U3949 (N_3949,N_3862,N_3819);
nand U3950 (N_3950,N_3850,N_3831);
and U3951 (N_3951,N_3847,N_3832);
or U3952 (N_3952,N_3852,N_3814);
nand U3953 (N_3953,N_3802,N_3847);
or U3954 (N_3954,N_3887,N_3849);
nand U3955 (N_3955,N_3848,N_3842);
and U3956 (N_3956,N_3852,N_3847);
or U3957 (N_3957,N_3898,N_3888);
nand U3958 (N_3958,N_3880,N_3839);
and U3959 (N_3959,N_3887,N_3877);
or U3960 (N_3960,N_3858,N_3892);
or U3961 (N_3961,N_3886,N_3804);
or U3962 (N_3962,N_3886,N_3893);
and U3963 (N_3963,N_3824,N_3851);
or U3964 (N_3964,N_3867,N_3871);
and U3965 (N_3965,N_3896,N_3862);
or U3966 (N_3966,N_3896,N_3820);
nor U3967 (N_3967,N_3895,N_3825);
nor U3968 (N_3968,N_3844,N_3805);
and U3969 (N_3969,N_3891,N_3818);
or U3970 (N_3970,N_3865,N_3884);
xnor U3971 (N_3971,N_3856,N_3808);
nor U3972 (N_3972,N_3862,N_3820);
or U3973 (N_3973,N_3808,N_3814);
nand U3974 (N_3974,N_3824,N_3821);
and U3975 (N_3975,N_3857,N_3888);
nor U3976 (N_3976,N_3851,N_3842);
nor U3977 (N_3977,N_3889,N_3858);
or U3978 (N_3978,N_3849,N_3854);
and U3979 (N_3979,N_3827,N_3854);
nand U3980 (N_3980,N_3871,N_3862);
or U3981 (N_3981,N_3869,N_3833);
nor U3982 (N_3982,N_3872,N_3847);
xnor U3983 (N_3983,N_3899,N_3821);
nor U3984 (N_3984,N_3886,N_3878);
and U3985 (N_3985,N_3877,N_3846);
nor U3986 (N_3986,N_3858,N_3835);
or U3987 (N_3987,N_3863,N_3821);
nor U3988 (N_3988,N_3854,N_3855);
and U3989 (N_3989,N_3886,N_3826);
and U3990 (N_3990,N_3841,N_3869);
nor U3991 (N_3991,N_3827,N_3825);
or U3992 (N_3992,N_3836,N_3858);
or U3993 (N_3993,N_3899,N_3850);
and U3994 (N_3994,N_3891,N_3849);
nand U3995 (N_3995,N_3828,N_3800);
nand U3996 (N_3996,N_3862,N_3838);
xor U3997 (N_3997,N_3845,N_3886);
nand U3998 (N_3998,N_3846,N_3870);
and U3999 (N_3999,N_3862,N_3803);
or U4000 (N_4000,N_3970,N_3913);
xor U4001 (N_4001,N_3926,N_3936);
nand U4002 (N_4002,N_3946,N_3920);
and U4003 (N_4003,N_3923,N_3968);
nand U4004 (N_4004,N_3972,N_3939);
nor U4005 (N_4005,N_3982,N_3911);
nand U4006 (N_4006,N_3960,N_3967);
nand U4007 (N_4007,N_3918,N_3990);
nor U4008 (N_4008,N_3979,N_3941);
or U4009 (N_4009,N_3925,N_3949);
or U4010 (N_4010,N_3916,N_3955);
and U4011 (N_4011,N_3977,N_3954);
and U4012 (N_4012,N_3997,N_3910);
nand U4013 (N_4013,N_3952,N_3956);
nor U4014 (N_4014,N_3933,N_3993);
nor U4015 (N_4015,N_3947,N_3986);
nand U4016 (N_4016,N_3905,N_3928);
or U4017 (N_4017,N_3973,N_3943);
or U4018 (N_4018,N_3981,N_3938);
or U4019 (N_4019,N_3976,N_3924);
or U4020 (N_4020,N_3994,N_3931);
nand U4021 (N_4021,N_3909,N_3922);
and U4022 (N_4022,N_3950,N_3987);
and U4023 (N_4023,N_3998,N_3921);
nand U4024 (N_4024,N_3945,N_3991);
and U4025 (N_4025,N_3958,N_3961);
or U4026 (N_4026,N_3989,N_3908);
and U4027 (N_4027,N_3959,N_3996);
nand U4028 (N_4028,N_3957,N_3900);
nand U4029 (N_4029,N_3965,N_3901);
or U4030 (N_4030,N_3906,N_3940);
nand U4031 (N_4031,N_3992,N_3902);
nand U4032 (N_4032,N_3944,N_3914);
nor U4033 (N_4033,N_3903,N_3912);
and U4034 (N_4034,N_3974,N_3937);
xor U4035 (N_4035,N_3975,N_3953);
nand U4036 (N_4036,N_3969,N_3932);
nor U4037 (N_4037,N_3915,N_3999);
xor U4038 (N_4038,N_3907,N_3995);
nor U4039 (N_4039,N_3927,N_3978);
nor U4040 (N_4040,N_3951,N_3948);
nand U4041 (N_4041,N_3930,N_3980);
nor U4042 (N_4042,N_3963,N_3904);
or U4043 (N_4043,N_3971,N_3934);
or U4044 (N_4044,N_3942,N_3985);
and U4045 (N_4045,N_3935,N_3919);
nor U4046 (N_4046,N_3966,N_3983);
nor U4047 (N_4047,N_3962,N_3964);
nand U4048 (N_4048,N_3929,N_3984);
nor U4049 (N_4049,N_3988,N_3917);
or U4050 (N_4050,N_3989,N_3934);
or U4051 (N_4051,N_3921,N_3941);
nor U4052 (N_4052,N_3981,N_3958);
and U4053 (N_4053,N_3973,N_3912);
nand U4054 (N_4054,N_3968,N_3998);
or U4055 (N_4055,N_3979,N_3973);
xor U4056 (N_4056,N_3926,N_3997);
nand U4057 (N_4057,N_3980,N_3920);
and U4058 (N_4058,N_3918,N_3987);
xor U4059 (N_4059,N_3913,N_3900);
nand U4060 (N_4060,N_3949,N_3968);
and U4061 (N_4061,N_3993,N_3984);
or U4062 (N_4062,N_3951,N_3989);
nand U4063 (N_4063,N_3982,N_3975);
or U4064 (N_4064,N_3919,N_3903);
nor U4065 (N_4065,N_3975,N_3915);
or U4066 (N_4066,N_3976,N_3939);
or U4067 (N_4067,N_3934,N_3906);
or U4068 (N_4068,N_3998,N_3924);
nor U4069 (N_4069,N_3963,N_3906);
or U4070 (N_4070,N_3934,N_3956);
nor U4071 (N_4071,N_3955,N_3993);
nand U4072 (N_4072,N_3945,N_3946);
or U4073 (N_4073,N_3912,N_3965);
and U4074 (N_4074,N_3981,N_3925);
nor U4075 (N_4075,N_3968,N_3913);
and U4076 (N_4076,N_3914,N_3995);
or U4077 (N_4077,N_3921,N_3908);
or U4078 (N_4078,N_3958,N_3985);
nor U4079 (N_4079,N_3950,N_3951);
nand U4080 (N_4080,N_3952,N_3992);
nand U4081 (N_4081,N_3968,N_3957);
nand U4082 (N_4082,N_3979,N_3962);
and U4083 (N_4083,N_3914,N_3939);
or U4084 (N_4084,N_3936,N_3972);
nor U4085 (N_4085,N_3965,N_3968);
and U4086 (N_4086,N_3995,N_3943);
nor U4087 (N_4087,N_3939,N_3989);
or U4088 (N_4088,N_3964,N_3912);
nand U4089 (N_4089,N_3905,N_3926);
nor U4090 (N_4090,N_3906,N_3976);
nand U4091 (N_4091,N_3967,N_3989);
nor U4092 (N_4092,N_3929,N_3939);
and U4093 (N_4093,N_3965,N_3946);
and U4094 (N_4094,N_3992,N_3921);
nor U4095 (N_4095,N_3940,N_3911);
and U4096 (N_4096,N_3916,N_3960);
nor U4097 (N_4097,N_3973,N_3902);
or U4098 (N_4098,N_3986,N_3998);
nor U4099 (N_4099,N_3976,N_3940);
nand U4100 (N_4100,N_4041,N_4055);
nand U4101 (N_4101,N_4054,N_4016);
nor U4102 (N_4102,N_4057,N_4064);
or U4103 (N_4103,N_4089,N_4094);
and U4104 (N_4104,N_4021,N_4097);
nor U4105 (N_4105,N_4080,N_4072);
and U4106 (N_4106,N_4098,N_4027);
nor U4107 (N_4107,N_4035,N_4062);
or U4108 (N_4108,N_4044,N_4034);
and U4109 (N_4109,N_4022,N_4050);
nor U4110 (N_4110,N_4066,N_4086);
or U4111 (N_4111,N_4006,N_4085);
xor U4112 (N_4112,N_4067,N_4031);
and U4113 (N_4113,N_4005,N_4040);
xor U4114 (N_4114,N_4036,N_4018);
xor U4115 (N_4115,N_4008,N_4015);
nand U4116 (N_4116,N_4019,N_4090);
or U4117 (N_4117,N_4047,N_4082);
or U4118 (N_4118,N_4013,N_4003);
and U4119 (N_4119,N_4049,N_4012);
and U4120 (N_4120,N_4033,N_4079);
and U4121 (N_4121,N_4026,N_4032);
or U4122 (N_4122,N_4092,N_4060);
nor U4123 (N_4123,N_4096,N_4077);
nand U4124 (N_4124,N_4071,N_4048);
and U4125 (N_4125,N_4068,N_4083);
nand U4126 (N_4126,N_4070,N_4078);
or U4127 (N_4127,N_4023,N_4051);
and U4128 (N_4128,N_4028,N_4029);
nor U4129 (N_4129,N_4061,N_4088);
nand U4130 (N_4130,N_4017,N_4099);
or U4131 (N_4131,N_4001,N_4075);
and U4132 (N_4132,N_4074,N_4073);
nand U4133 (N_4133,N_4069,N_4065);
nor U4134 (N_4134,N_4076,N_4039);
and U4135 (N_4135,N_4087,N_4058);
nor U4136 (N_4136,N_4063,N_4002);
nand U4137 (N_4137,N_4024,N_4020);
and U4138 (N_4138,N_4081,N_4000);
nor U4139 (N_4139,N_4037,N_4038);
or U4140 (N_4140,N_4010,N_4011);
nor U4141 (N_4141,N_4042,N_4091);
nor U4142 (N_4142,N_4052,N_4004);
xnor U4143 (N_4143,N_4056,N_4093);
or U4144 (N_4144,N_4007,N_4045);
and U4145 (N_4145,N_4084,N_4030);
nand U4146 (N_4146,N_4009,N_4059);
or U4147 (N_4147,N_4053,N_4043);
and U4148 (N_4148,N_4014,N_4025);
nand U4149 (N_4149,N_4095,N_4046);
or U4150 (N_4150,N_4081,N_4077);
nor U4151 (N_4151,N_4060,N_4041);
or U4152 (N_4152,N_4054,N_4076);
xor U4153 (N_4153,N_4020,N_4045);
or U4154 (N_4154,N_4038,N_4035);
or U4155 (N_4155,N_4099,N_4012);
and U4156 (N_4156,N_4014,N_4033);
or U4157 (N_4157,N_4022,N_4085);
nand U4158 (N_4158,N_4006,N_4081);
or U4159 (N_4159,N_4079,N_4000);
nor U4160 (N_4160,N_4072,N_4012);
nor U4161 (N_4161,N_4002,N_4062);
xnor U4162 (N_4162,N_4093,N_4084);
and U4163 (N_4163,N_4023,N_4063);
nor U4164 (N_4164,N_4057,N_4051);
nand U4165 (N_4165,N_4089,N_4007);
nor U4166 (N_4166,N_4013,N_4040);
nand U4167 (N_4167,N_4029,N_4032);
and U4168 (N_4168,N_4083,N_4097);
or U4169 (N_4169,N_4019,N_4067);
and U4170 (N_4170,N_4041,N_4012);
xnor U4171 (N_4171,N_4079,N_4019);
nor U4172 (N_4172,N_4045,N_4046);
nor U4173 (N_4173,N_4028,N_4084);
and U4174 (N_4174,N_4014,N_4080);
nor U4175 (N_4175,N_4061,N_4085);
and U4176 (N_4176,N_4039,N_4075);
or U4177 (N_4177,N_4015,N_4052);
and U4178 (N_4178,N_4050,N_4077);
and U4179 (N_4179,N_4047,N_4000);
nand U4180 (N_4180,N_4054,N_4028);
nand U4181 (N_4181,N_4033,N_4045);
and U4182 (N_4182,N_4058,N_4005);
and U4183 (N_4183,N_4056,N_4060);
xnor U4184 (N_4184,N_4046,N_4022);
or U4185 (N_4185,N_4097,N_4074);
nand U4186 (N_4186,N_4000,N_4063);
or U4187 (N_4187,N_4085,N_4089);
or U4188 (N_4188,N_4001,N_4094);
nand U4189 (N_4189,N_4025,N_4068);
nor U4190 (N_4190,N_4065,N_4059);
and U4191 (N_4191,N_4003,N_4033);
and U4192 (N_4192,N_4019,N_4059);
and U4193 (N_4193,N_4059,N_4097);
nor U4194 (N_4194,N_4077,N_4015);
or U4195 (N_4195,N_4075,N_4018);
xnor U4196 (N_4196,N_4043,N_4061);
nand U4197 (N_4197,N_4011,N_4076);
nor U4198 (N_4198,N_4047,N_4085);
nor U4199 (N_4199,N_4085,N_4003);
or U4200 (N_4200,N_4158,N_4130);
and U4201 (N_4201,N_4175,N_4177);
and U4202 (N_4202,N_4117,N_4111);
and U4203 (N_4203,N_4144,N_4169);
nor U4204 (N_4204,N_4120,N_4142);
nor U4205 (N_4205,N_4171,N_4195);
and U4206 (N_4206,N_4164,N_4129);
nor U4207 (N_4207,N_4104,N_4118);
nor U4208 (N_4208,N_4178,N_4149);
or U4209 (N_4209,N_4137,N_4191);
or U4210 (N_4210,N_4115,N_4190);
nor U4211 (N_4211,N_4152,N_4173);
xor U4212 (N_4212,N_4102,N_4124);
or U4213 (N_4213,N_4127,N_4131);
nand U4214 (N_4214,N_4194,N_4189);
xnor U4215 (N_4215,N_4160,N_4167);
and U4216 (N_4216,N_4133,N_4122);
nor U4217 (N_4217,N_4192,N_4110);
xnor U4218 (N_4218,N_4125,N_4163);
xor U4219 (N_4219,N_4151,N_4150);
nor U4220 (N_4220,N_4198,N_4119);
nand U4221 (N_4221,N_4196,N_4146);
nor U4222 (N_4222,N_4145,N_4165);
nand U4223 (N_4223,N_4139,N_4181);
nand U4224 (N_4224,N_4186,N_4116);
nor U4225 (N_4225,N_4193,N_4199);
nand U4226 (N_4226,N_4101,N_4157);
nand U4227 (N_4227,N_4174,N_4162);
and U4228 (N_4228,N_4123,N_4170);
xnor U4229 (N_4229,N_4148,N_4182);
or U4230 (N_4230,N_4183,N_4113);
xnor U4231 (N_4231,N_4141,N_4184);
and U4232 (N_4232,N_4105,N_4179);
or U4233 (N_4233,N_4126,N_4135);
nand U4234 (N_4234,N_4103,N_4168);
nand U4235 (N_4235,N_4100,N_4140);
nor U4236 (N_4236,N_4109,N_4188);
and U4237 (N_4237,N_4153,N_4176);
nand U4238 (N_4238,N_4187,N_4128);
xnor U4239 (N_4239,N_4143,N_4108);
nand U4240 (N_4240,N_4166,N_4136);
and U4241 (N_4241,N_4156,N_4154);
or U4242 (N_4242,N_4114,N_4106);
and U4243 (N_4243,N_4107,N_4172);
or U4244 (N_4244,N_4147,N_4159);
nand U4245 (N_4245,N_4112,N_4134);
xor U4246 (N_4246,N_4180,N_4132);
or U4247 (N_4247,N_4155,N_4138);
nand U4248 (N_4248,N_4197,N_4161);
and U4249 (N_4249,N_4185,N_4121);
and U4250 (N_4250,N_4115,N_4159);
nor U4251 (N_4251,N_4177,N_4194);
and U4252 (N_4252,N_4156,N_4181);
and U4253 (N_4253,N_4177,N_4156);
or U4254 (N_4254,N_4169,N_4123);
or U4255 (N_4255,N_4199,N_4168);
nand U4256 (N_4256,N_4109,N_4141);
and U4257 (N_4257,N_4131,N_4196);
or U4258 (N_4258,N_4167,N_4163);
nor U4259 (N_4259,N_4196,N_4134);
nor U4260 (N_4260,N_4117,N_4179);
nor U4261 (N_4261,N_4142,N_4109);
and U4262 (N_4262,N_4170,N_4111);
and U4263 (N_4263,N_4118,N_4168);
or U4264 (N_4264,N_4118,N_4141);
nand U4265 (N_4265,N_4143,N_4149);
and U4266 (N_4266,N_4183,N_4187);
nand U4267 (N_4267,N_4171,N_4156);
nand U4268 (N_4268,N_4125,N_4100);
or U4269 (N_4269,N_4127,N_4198);
nor U4270 (N_4270,N_4162,N_4141);
nor U4271 (N_4271,N_4136,N_4151);
xnor U4272 (N_4272,N_4146,N_4139);
nor U4273 (N_4273,N_4170,N_4191);
xor U4274 (N_4274,N_4105,N_4108);
nor U4275 (N_4275,N_4194,N_4186);
xor U4276 (N_4276,N_4131,N_4152);
or U4277 (N_4277,N_4184,N_4183);
and U4278 (N_4278,N_4182,N_4194);
or U4279 (N_4279,N_4133,N_4151);
nand U4280 (N_4280,N_4198,N_4195);
nand U4281 (N_4281,N_4173,N_4143);
nor U4282 (N_4282,N_4113,N_4124);
nand U4283 (N_4283,N_4158,N_4172);
xnor U4284 (N_4284,N_4174,N_4140);
nor U4285 (N_4285,N_4196,N_4124);
nor U4286 (N_4286,N_4114,N_4107);
or U4287 (N_4287,N_4193,N_4120);
and U4288 (N_4288,N_4144,N_4116);
and U4289 (N_4289,N_4134,N_4114);
nand U4290 (N_4290,N_4103,N_4162);
nand U4291 (N_4291,N_4138,N_4113);
or U4292 (N_4292,N_4109,N_4158);
xor U4293 (N_4293,N_4125,N_4155);
or U4294 (N_4294,N_4135,N_4166);
nand U4295 (N_4295,N_4193,N_4191);
and U4296 (N_4296,N_4148,N_4116);
nor U4297 (N_4297,N_4119,N_4159);
or U4298 (N_4298,N_4193,N_4123);
and U4299 (N_4299,N_4135,N_4119);
or U4300 (N_4300,N_4281,N_4232);
or U4301 (N_4301,N_4205,N_4210);
nor U4302 (N_4302,N_4294,N_4217);
or U4303 (N_4303,N_4216,N_4278);
nand U4304 (N_4304,N_4248,N_4207);
xor U4305 (N_4305,N_4263,N_4231);
nor U4306 (N_4306,N_4246,N_4271);
nor U4307 (N_4307,N_4285,N_4242);
nand U4308 (N_4308,N_4243,N_4274);
nor U4309 (N_4309,N_4229,N_4250);
xnor U4310 (N_4310,N_4286,N_4213);
nor U4311 (N_4311,N_4225,N_4245);
nor U4312 (N_4312,N_4208,N_4262);
or U4313 (N_4313,N_4260,N_4235);
and U4314 (N_4314,N_4266,N_4237);
nor U4315 (N_4315,N_4206,N_4254);
nand U4316 (N_4316,N_4288,N_4273);
and U4317 (N_4317,N_4203,N_4283);
or U4318 (N_4318,N_4298,N_4277);
nand U4319 (N_4319,N_4290,N_4226);
nand U4320 (N_4320,N_4299,N_4253);
xor U4321 (N_4321,N_4264,N_4219);
or U4322 (N_4322,N_4238,N_4292);
xnor U4323 (N_4323,N_4230,N_4222);
or U4324 (N_4324,N_4202,N_4236);
nand U4325 (N_4325,N_4227,N_4247);
nand U4326 (N_4326,N_4295,N_4221);
or U4327 (N_4327,N_4267,N_4244);
xnor U4328 (N_4328,N_4265,N_4270);
nor U4329 (N_4329,N_4215,N_4223);
nor U4330 (N_4330,N_4293,N_4269);
and U4331 (N_4331,N_4249,N_4284);
and U4332 (N_4332,N_4239,N_4276);
nor U4333 (N_4333,N_4296,N_4287);
nor U4334 (N_4334,N_4224,N_4291);
or U4335 (N_4335,N_4214,N_4272);
and U4336 (N_4336,N_4220,N_4252);
xor U4337 (N_4337,N_4261,N_4200);
nand U4338 (N_4338,N_4218,N_4204);
nand U4339 (N_4339,N_4257,N_4233);
nand U4340 (N_4340,N_4275,N_4279);
nor U4341 (N_4341,N_4209,N_4251);
nor U4342 (N_4342,N_4259,N_4268);
nor U4343 (N_4343,N_4256,N_4212);
and U4344 (N_4344,N_4211,N_4240);
nor U4345 (N_4345,N_4280,N_4282);
nor U4346 (N_4346,N_4258,N_4297);
nand U4347 (N_4347,N_4201,N_4234);
nor U4348 (N_4348,N_4289,N_4228);
or U4349 (N_4349,N_4255,N_4241);
nor U4350 (N_4350,N_4299,N_4280);
and U4351 (N_4351,N_4290,N_4223);
xor U4352 (N_4352,N_4252,N_4228);
nand U4353 (N_4353,N_4219,N_4225);
or U4354 (N_4354,N_4275,N_4291);
or U4355 (N_4355,N_4243,N_4204);
nand U4356 (N_4356,N_4205,N_4283);
nand U4357 (N_4357,N_4220,N_4281);
and U4358 (N_4358,N_4273,N_4264);
or U4359 (N_4359,N_4213,N_4237);
xnor U4360 (N_4360,N_4255,N_4257);
nand U4361 (N_4361,N_4235,N_4248);
xor U4362 (N_4362,N_4288,N_4238);
or U4363 (N_4363,N_4257,N_4256);
nor U4364 (N_4364,N_4231,N_4274);
and U4365 (N_4365,N_4243,N_4238);
nor U4366 (N_4366,N_4266,N_4230);
nor U4367 (N_4367,N_4218,N_4293);
or U4368 (N_4368,N_4281,N_4245);
or U4369 (N_4369,N_4290,N_4285);
or U4370 (N_4370,N_4257,N_4251);
or U4371 (N_4371,N_4222,N_4204);
xnor U4372 (N_4372,N_4257,N_4203);
and U4373 (N_4373,N_4294,N_4256);
nor U4374 (N_4374,N_4283,N_4287);
and U4375 (N_4375,N_4244,N_4200);
and U4376 (N_4376,N_4296,N_4215);
nand U4377 (N_4377,N_4201,N_4207);
or U4378 (N_4378,N_4255,N_4277);
or U4379 (N_4379,N_4216,N_4200);
nor U4380 (N_4380,N_4214,N_4271);
or U4381 (N_4381,N_4212,N_4261);
and U4382 (N_4382,N_4253,N_4279);
or U4383 (N_4383,N_4215,N_4269);
nand U4384 (N_4384,N_4261,N_4283);
and U4385 (N_4385,N_4239,N_4292);
nor U4386 (N_4386,N_4247,N_4285);
or U4387 (N_4387,N_4256,N_4230);
nor U4388 (N_4388,N_4251,N_4235);
and U4389 (N_4389,N_4212,N_4280);
nor U4390 (N_4390,N_4223,N_4252);
nor U4391 (N_4391,N_4278,N_4292);
and U4392 (N_4392,N_4267,N_4255);
nand U4393 (N_4393,N_4295,N_4250);
and U4394 (N_4394,N_4229,N_4225);
and U4395 (N_4395,N_4289,N_4275);
nor U4396 (N_4396,N_4228,N_4259);
or U4397 (N_4397,N_4248,N_4218);
xnor U4398 (N_4398,N_4225,N_4221);
or U4399 (N_4399,N_4270,N_4212);
or U4400 (N_4400,N_4302,N_4370);
or U4401 (N_4401,N_4396,N_4352);
nand U4402 (N_4402,N_4308,N_4349);
nand U4403 (N_4403,N_4377,N_4399);
and U4404 (N_4404,N_4318,N_4342);
nand U4405 (N_4405,N_4378,N_4311);
or U4406 (N_4406,N_4363,N_4393);
nand U4407 (N_4407,N_4330,N_4392);
nor U4408 (N_4408,N_4367,N_4382);
nor U4409 (N_4409,N_4358,N_4300);
or U4410 (N_4410,N_4316,N_4375);
nor U4411 (N_4411,N_4306,N_4356);
nand U4412 (N_4412,N_4337,N_4334);
nand U4413 (N_4413,N_4322,N_4313);
xnor U4414 (N_4414,N_4338,N_4387);
nand U4415 (N_4415,N_4343,N_4353);
or U4416 (N_4416,N_4325,N_4365);
or U4417 (N_4417,N_4321,N_4351);
nor U4418 (N_4418,N_4340,N_4398);
nor U4419 (N_4419,N_4303,N_4357);
nor U4420 (N_4420,N_4383,N_4355);
or U4421 (N_4421,N_4344,N_4320);
or U4422 (N_4422,N_4366,N_4362);
nand U4423 (N_4423,N_4345,N_4326);
nand U4424 (N_4424,N_4372,N_4339);
xor U4425 (N_4425,N_4374,N_4359);
nor U4426 (N_4426,N_4335,N_4336);
nor U4427 (N_4427,N_4394,N_4389);
nor U4428 (N_4428,N_4368,N_4397);
nand U4429 (N_4429,N_4310,N_4323);
nand U4430 (N_4430,N_4341,N_4348);
nand U4431 (N_4431,N_4379,N_4369);
nand U4432 (N_4432,N_4312,N_4385);
xor U4433 (N_4433,N_4384,N_4346);
nand U4434 (N_4434,N_4301,N_4328);
or U4435 (N_4435,N_4381,N_4373);
nor U4436 (N_4436,N_4317,N_4329);
and U4437 (N_4437,N_4371,N_4376);
and U4438 (N_4438,N_4314,N_4327);
and U4439 (N_4439,N_4350,N_4307);
nand U4440 (N_4440,N_4380,N_4324);
or U4441 (N_4441,N_4309,N_4315);
or U4442 (N_4442,N_4391,N_4354);
nor U4443 (N_4443,N_4386,N_4390);
and U4444 (N_4444,N_4304,N_4305);
nand U4445 (N_4445,N_4395,N_4331);
nand U4446 (N_4446,N_4347,N_4332);
and U4447 (N_4447,N_4388,N_4319);
nor U4448 (N_4448,N_4361,N_4360);
and U4449 (N_4449,N_4364,N_4333);
nand U4450 (N_4450,N_4369,N_4371);
xnor U4451 (N_4451,N_4312,N_4378);
nor U4452 (N_4452,N_4360,N_4345);
or U4453 (N_4453,N_4312,N_4393);
nand U4454 (N_4454,N_4382,N_4363);
and U4455 (N_4455,N_4397,N_4356);
nor U4456 (N_4456,N_4313,N_4332);
or U4457 (N_4457,N_4396,N_4367);
nor U4458 (N_4458,N_4383,N_4393);
or U4459 (N_4459,N_4337,N_4392);
nand U4460 (N_4460,N_4374,N_4300);
and U4461 (N_4461,N_4324,N_4333);
or U4462 (N_4462,N_4334,N_4311);
nand U4463 (N_4463,N_4350,N_4328);
and U4464 (N_4464,N_4396,N_4344);
nor U4465 (N_4465,N_4382,N_4312);
and U4466 (N_4466,N_4355,N_4313);
nor U4467 (N_4467,N_4381,N_4365);
and U4468 (N_4468,N_4383,N_4308);
nor U4469 (N_4469,N_4368,N_4388);
and U4470 (N_4470,N_4376,N_4362);
nor U4471 (N_4471,N_4362,N_4348);
nor U4472 (N_4472,N_4385,N_4314);
and U4473 (N_4473,N_4333,N_4341);
and U4474 (N_4474,N_4380,N_4309);
and U4475 (N_4475,N_4305,N_4354);
or U4476 (N_4476,N_4393,N_4345);
nor U4477 (N_4477,N_4308,N_4351);
or U4478 (N_4478,N_4318,N_4378);
nor U4479 (N_4479,N_4340,N_4362);
or U4480 (N_4480,N_4378,N_4383);
nor U4481 (N_4481,N_4312,N_4362);
nand U4482 (N_4482,N_4302,N_4313);
and U4483 (N_4483,N_4348,N_4331);
nor U4484 (N_4484,N_4353,N_4325);
xor U4485 (N_4485,N_4327,N_4339);
and U4486 (N_4486,N_4345,N_4371);
nand U4487 (N_4487,N_4309,N_4322);
nand U4488 (N_4488,N_4361,N_4316);
xnor U4489 (N_4489,N_4307,N_4363);
and U4490 (N_4490,N_4316,N_4394);
or U4491 (N_4491,N_4314,N_4336);
xor U4492 (N_4492,N_4391,N_4363);
nor U4493 (N_4493,N_4339,N_4337);
nand U4494 (N_4494,N_4393,N_4361);
or U4495 (N_4495,N_4366,N_4301);
and U4496 (N_4496,N_4334,N_4389);
nand U4497 (N_4497,N_4311,N_4377);
nor U4498 (N_4498,N_4313,N_4361);
nor U4499 (N_4499,N_4388,N_4393);
nor U4500 (N_4500,N_4458,N_4428);
nor U4501 (N_4501,N_4433,N_4463);
and U4502 (N_4502,N_4462,N_4464);
or U4503 (N_4503,N_4480,N_4418);
nor U4504 (N_4504,N_4496,N_4429);
xor U4505 (N_4505,N_4423,N_4424);
or U4506 (N_4506,N_4425,N_4414);
or U4507 (N_4507,N_4448,N_4498);
nor U4508 (N_4508,N_4432,N_4446);
nand U4509 (N_4509,N_4475,N_4419);
nor U4510 (N_4510,N_4474,N_4416);
nand U4511 (N_4511,N_4461,N_4465);
and U4512 (N_4512,N_4412,N_4497);
and U4513 (N_4513,N_4487,N_4452);
nand U4514 (N_4514,N_4499,N_4420);
xnor U4515 (N_4515,N_4473,N_4410);
and U4516 (N_4516,N_4489,N_4482);
and U4517 (N_4517,N_4495,N_4454);
nor U4518 (N_4518,N_4401,N_4456);
nor U4519 (N_4519,N_4453,N_4457);
nor U4520 (N_4520,N_4427,N_4434);
nand U4521 (N_4521,N_4493,N_4404);
nand U4522 (N_4522,N_4491,N_4478);
nor U4523 (N_4523,N_4466,N_4402);
and U4524 (N_4524,N_4445,N_4407);
or U4525 (N_4525,N_4488,N_4447);
nor U4526 (N_4526,N_4486,N_4439);
nand U4527 (N_4527,N_4421,N_4413);
or U4528 (N_4528,N_4469,N_4455);
or U4529 (N_4529,N_4409,N_4411);
nor U4530 (N_4530,N_4405,N_4449);
nor U4531 (N_4531,N_4426,N_4435);
and U4532 (N_4532,N_4481,N_4467);
or U4533 (N_4533,N_4451,N_4494);
or U4534 (N_4534,N_4470,N_4479);
and U4535 (N_4535,N_4415,N_4492);
nor U4536 (N_4536,N_4437,N_4408);
nand U4537 (N_4537,N_4406,N_4490);
nor U4538 (N_4538,N_4441,N_4417);
or U4539 (N_4539,N_4476,N_4442);
and U4540 (N_4540,N_4477,N_4440);
or U4541 (N_4541,N_4403,N_4471);
nand U4542 (N_4542,N_4443,N_4400);
nand U4543 (N_4543,N_4460,N_4436);
nand U4544 (N_4544,N_4444,N_4484);
nor U4545 (N_4545,N_4468,N_4422);
nand U4546 (N_4546,N_4485,N_4430);
nand U4547 (N_4547,N_4450,N_4459);
or U4548 (N_4548,N_4438,N_4472);
xor U4549 (N_4549,N_4483,N_4431);
xor U4550 (N_4550,N_4473,N_4456);
nor U4551 (N_4551,N_4420,N_4411);
and U4552 (N_4552,N_4407,N_4498);
and U4553 (N_4553,N_4418,N_4499);
nor U4554 (N_4554,N_4444,N_4439);
nor U4555 (N_4555,N_4470,N_4497);
nor U4556 (N_4556,N_4432,N_4491);
or U4557 (N_4557,N_4460,N_4403);
or U4558 (N_4558,N_4401,N_4413);
nand U4559 (N_4559,N_4454,N_4447);
nor U4560 (N_4560,N_4487,N_4438);
and U4561 (N_4561,N_4429,N_4420);
nor U4562 (N_4562,N_4484,N_4457);
or U4563 (N_4563,N_4431,N_4489);
or U4564 (N_4564,N_4419,N_4466);
nand U4565 (N_4565,N_4453,N_4498);
nor U4566 (N_4566,N_4496,N_4465);
nand U4567 (N_4567,N_4416,N_4408);
nor U4568 (N_4568,N_4495,N_4465);
and U4569 (N_4569,N_4453,N_4423);
nand U4570 (N_4570,N_4461,N_4452);
and U4571 (N_4571,N_4464,N_4460);
nor U4572 (N_4572,N_4483,N_4485);
nand U4573 (N_4573,N_4411,N_4488);
nand U4574 (N_4574,N_4485,N_4494);
and U4575 (N_4575,N_4487,N_4475);
nand U4576 (N_4576,N_4485,N_4416);
and U4577 (N_4577,N_4463,N_4470);
and U4578 (N_4578,N_4414,N_4469);
nor U4579 (N_4579,N_4458,N_4423);
and U4580 (N_4580,N_4428,N_4491);
xnor U4581 (N_4581,N_4450,N_4427);
nor U4582 (N_4582,N_4468,N_4482);
and U4583 (N_4583,N_4445,N_4484);
or U4584 (N_4584,N_4488,N_4492);
and U4585 (N_4585,N_4483,N_4441);
or U4586 (N_4586,N_4439,N_4494);
and U4587 (N_4587,N_4434,N_4485);
or U4588 (N_4588,N_4449,N_4409);
nor U4589 (N_4589,N_4440,N_4409);
or U4590 (N_4590,N_4497,N_4479);
nand U4591 (N_4591,N_4416,N_4429);
nand U4592 (N_4592,N_4403,N_4483);
and U4593 (N_4593,N_4421,N_4400);
nand U4594 (N_4594,N_4402,N_4451);
nor U4595 (N_4595,N_4431,N_4424);
or U4596 (N_4596,N_4470,N_4408);
nor U4597 (N_4597,N_4413,N_4430);
nand U4598 (N_4598,N_4473,N_4479);
nor U4599 (N_4599,N_4478,N_4418);
nor U4600 (N_4600,N_4568,N_4540);
nand U4601 (N_4601,N_4579,N_4560);
or U4602 (N_4602,N_4526,N_4510);
or U4603 (N_4603,N_4533,N_4553);
nand U4604 (N_4604,N_4524,N_4506);
nand U4605 (N_4605,N_4539,N_4507);
or U4606 (N_4606,N_4552,N_4523);
nand U4607 (N_4607,N_4555,N_4550);
nand U4608 (N_4608,N_4554,N_4512);
and U4609 (N_4609,N_4536,N_4580);
nand U4610 (N_4610,N_4573,N_4578);
nand U4611 (N_4611,N_4530,N_4570);
nand U4612 (N_4612,N_4503,N_4547);
nand U4613 (N_4613,N_4516,N_4504);
nor U4614 (N_4614,N_4527,N_4549);
nand U4615 (N_4615,N_4586,N_4567);
xnor U4616 (N_4616,N_4592,N_4569);
or U4617 (N_4617,N_4520,N_4597);
and U4618 (N_4618,N_4528,N_4521);
or U4619 (N_4619,N_4517,N_4563);
or U4620 (N_4620,N_4591,N_4543);
or U4621 (N_4621,N_4593,N_4588);
nand U4622 (N_4622,N_4585,N_4508);
nor U4623 (N_4623,N_4582,N_4529);
nor U4624 (N_4624,N_4546,N_4574);
nand U4625 (N_4625,N_4500,N_4515);
or U4626 (N_4626,N_4566,N_4590);
and U4627 (N_4627,N_4589,N_4557);
or U4628 (N_4628,N_4561,N_4575);
and U4629 (N_4629,N_4502,N_4596);
and U4630 (N_4630,N_4511,N_4537);
xnor U4631 (N_4631,N_4513,N_4584);
and U4632 (N_4632,N_4562,N_4598);
or U4633 (N_4633,N_4559,N_4501);
and U4634 (N_4634,N_4522,N_4525);
xor U4635 (N_4635,N_4583,N_4594);
xnor U4636 (N_4636,N_4571,N_4534);
xor U4637 (N_4637,N_4531,N_4587);
nor U4638 (N_4638,N_4572,N_4542);
nand U4639 (N_4639,N_4551,N_4505);
nand U4640 (N_4640,N_4576,N_4518);
or U4641 (N_4641,N_4541,N_4581);
nor U4642 (N_4642,N_4532,N_4577);
or U4643 (N_4643,N_4564,N_4544);
or U4644 (N_4644,N_4558,N_4509);
nand U4645 (N_4645,N_4595,N_4556);
nand U4646 (N_4646,N_4519,N_4545);
or U4647 (N_4647,N_4535,N_4599);
and U4648 (N_4648,N_4548,N_4538);
nand U4649 (N_4649,N_4514,N_4565);
and U4650 (N_4650,N_4584,N_4508);
and U4651 (N_4651,N_4548,N_4591);
xnor U4652 (N_4652,N_4548,N_4514);
or U4653 (N_4653,N_4546,N_4580);
nor U4654 (N_4654,N_4506,N_4589);
nand U4655 (N_4655,N_4500,N_4569);
nor U4656 (N_4656,N_4582,N_4575);
or U4657 (N_4657,N_4519,N_4553);
and U4658 (N_4658,N_4502,N_4514);
or U4659 (N_4659,N_4551,N_4548);
or U4660 (N_4660,N_4508,N_4533);
nand U4661 (N_4661,N_4519,N_4582);
and U4662 (N_4662,N_4584,N_4543);
and U4663 (N_4663,N_4559,N_4554);
nand U4664 (N_4664,N_4544,N_4521);
xnor U4665 (N_4665,N_4544,N_4535);
or U4666 (N_4666,N_4547,N_4528);
nand U4667 (N_4667,N_4546,N_4549);
nand U4668 (N_4668,N_4591,N_4534);
nand U4669 (N_4669,N_4541,N_4538);
or U4670 (N_4670,N_4542,N_4573);
and U4671 (N_4671,N_4526,N_4565);
and U4672 (N_4672,N_4505,N_4516);
and U4673 (N_4673,N_4537,N_4563);
and U4674 (N_4674,N_4505,N_4537);
and U4675 (N_4675,N_4539,N_4530);
nand U4676 (N_4676,N_4530,N_4508);
or U4677 (N_4677,N_4542,N_4553);
and U4678 (N_4678,N_4508,N_4532);
nor U4679 (N_4679,N_4535,N_4598);
nor U4680 (N_4680,N_4575,N_4542);
nand U4681 (N_4681,N_4551,N_4588);
or U4682 (N_4682,N_4526,N_4504);
and U4683 (N_4683,N_4550,N_4501);
xnor U4684 (N_4684,N_4530,N_4517);
or U4685 (N_4685,N_4532,N_4555);
nor U4686 (N_4686,N_4553,N_4592);
nor U4687 (N_4687,N_4579,N_4512);
and U4688 (N_4688,N_4516,N_4599);
nor U4689 (N_4689,N_4528,N_4597);
nand U4690 (N_4690,N_4556,N_4501);
nand U4691 (N_4691,N_4565,N_4502);
and U4692 (N_4692,N_4556,N_4517);
nand U4693 (N_4693,N_4565,N_4577);
xor U4694 (N_4694,N_4581,N_4510);
nor U4695 (N_4695,N_4500,N_4589);
nor U4696 (N_4696,N_4534,N_4507);
nor U4697 (N_4697,N_4561,N_4506);
nand U4698 (N_4698,N_4560,N_4547);
or U4699 (N_4699,N_4514,N_4576);
nor U4700 (N_4700,N_4625,N_4646);
or U4701 (N_4701,N_4654,N_4614);
or U4702 (N_4702,N_4679,N_4692);
or U4703 (N_4703,N_4662,N_4612);
or U4704 (N_4704,N_4673,N_4642);
nand U4705 (N_4705,N_4630,N_4652);
xnor U4706 (N_4706,N_4670,N_4622);
nor U4707 (N_4707,N_4695,N_4620);
nand U4708 (N_4708,N_4660,N_4666);
and U4709 (N_4709,N_4623,N_4686);
or U4710 (N_4710,N_4619,N_4636);
nand U4711 (N_4711,N_4665,N_4610);
and U4712 (N_4712,N_4635,N_4604);
and U4713 (N_4713,N_4653,N_4637);
and U4714 (N_4714,N_4603,N_4668);
and U4715 (N_4715,N_4606,N_4659);
and U4716 (N_4716,N_4697,N_4651);
xnor U4717 (N_4717,N_4617,N_4641);
nor U4718 (N_4718,N_4634,N_4616);
nor U4719 (N_4719,N_4672,N_4627);
or U4720 (N_4720,N_4631,N_4685);
nor U4721 (N_4721,N_4655,N_4680);
or U4722 (N_4722,N_4676,N_4601);
and U4723 (N_4723,N_4691,N_4687);
and U4724 (N_4724,N_4664,N_4600);
or U4725 (N_4725,N_4693,N_4657);
nand U4726 (N_4726,N_4645,N_4694);
xor U4727 (N_4727,N_4633,N_4639);
nor U4728 (N_4728,N_4650,N_4643);
nor U4729 (N_4729,N_4667,N_4632);
and U4730 (N_4730,N_4688,N_4611);
nor U4731 (N_4731,N_4621,N_4648);
or U4732 (N_4732,N_4698,N_4644);
or U4733 (N_4733,N_4690,N_4684);
xnor U4734 (N_4734,N_4629,N_4689);
or U4735 (N_4735,N_4609,N_4607);
nand U4736 (N_4736,N_4675,N_4656);
or U4737 (N_4737,N_4658,N_4661);
nand U4738 (N_4738,N_4640,N_4663);
nor U4739 (N_4739,N_4618,N_4638);
nor U4740 (N_4740,N_4696,N_4628);
and U4741 (N_4741,N_4649,N_4602);
xnor U4742 (N_4742,N_4626,N_4681);
xnor U4743 (N_4743,N_4674,N_4671);
and U4744 (N_4744,N_4624,N_4647);
nand U4745 (N_4745,N_4605,N_4677);
nor U4746 (N_4746,N_4615,N_4682);
and U4747 (N_4747,N_4669,N_4699);
or U4748 (N_4748,N_4683,N_4678);
nor U4749 (N_4749,N_4613,N_4608);
nand U4750 (N_4750,N_4627,N_4666);
or U4751 (N_4751,N_4690,N_4652);
xnor U4752 (N_4752,N_4673,N_4694);
or U4753 (N_4753,N_4608,N_4636);
nand U4754 (N_4754,N_4647,N_4614);
and U4755 (N_4755,N_4667,N_4648);
nand U4756 (N_4756,N_4682,N_4695);
nand U4757 (N_4757,N_4676,N_4651);
nand U4758 (N_4758,N_4696,N_4618);
or U4759 (N_4759,N_4626,N_4683);
and U4760 (N_4760,N_4689,N_4658);
xnor U4761 (N_4761,N_4677,N_4657);
and U4762 (N_4762,N_4621,N_4622);
and U4763 (N_4763,N_4695,N_4654);
nor U4764 (N_4764,N_4636,N_4690);
or U4765 (N_4765,N_4671,N_4649);
and U4766 (N_4766,N_4604,N_4660);
xor U4767 (N_4767,N_4602,N_4660);
and U4768 (N_4768,N_4602,N_4646);
nand U4769 (N_4769,N_4661,N_4684);
or U4770 (N_4770,N_4699,N_4611);
nand U4771 (N_4771,N_4618,N_4649);
or U4772 (N_4772,N_4654,N_4682);
and U4773 (N_4773,N_4690,N_4635);
or U4774 (N_4774,N_4661,N_4649);
nor U4775 (N_4775,N_4610,N_4629);
or U4776 (N_4776,N_4674,N_4691);
or U4777 (N_4777,N_4662,N_4680);
and U4778 (N_4778,N_4610,N_4642);
or U4779 (N_4779,N_4691,N_4616);
nand U4780 (N_4780,N_4632,N_4692);
nor U4781 (N_4781,N_4601,N_4649);
or U4782 (N_4782,N_4632,N_4690);
xnor U4783 (N_4783,N_4693,N_4604);
and U4784 (N_4784,N_4692,N_4652);
and U4785 (N_4785,N_4662,N_4655);
or U4786 (N_4786,N_4606,N_4660);
nand U4787 (N_4787,N_4647,N_4679);
nand U4788 (N_4788,N_4690,N_4691);
nor U4789 (N_4789,N_4623,N_4642);
or U4790 (N_4790,N_4651,N_4625);
xnor U4791 (N_4791,N_4600,N_4668);
nor U4792 (N_4792,N_4609,N_4629);
nand U4793 (N_4793,N_4633,N_4678);
nand U4794 (N_4794,N_4663,N_4603);
and U4795 (N_4795,N_4650,N_4660);
nor U4796 (N_4796,N_4606,N_4680);
nand U4797 (N_4797,N_4675,N_4613);
and U4798 (N_4798,N_4629,N_4695);
nand U4799 (N_4799,N_4638,N_4680);
and U4800 (N_4800,N_4784,N_4745);
nor U4801 (N_4801,N_4777,N_4761);
and U4802 (N_4802,N_4778,N_4791);
and U4803 (N_4803,N_4722,N_4783);
and U4804 (N_4804,N_4727,N_4743);
nor U4805 (N_4805,N_4782,N_4730);
or U4806 (N_4806,N_4780,N_4793);
nand U4807 (N_4807,N_4751,N_4706);
or U4808 (N_4808,N_4746,N_4701);
or U4809 (N_4809,N_4715,N_4726);
nand U4810 (N_4810,N_4779,N_4764);
or U4811 (N_4811,N_4772,N_4705);
nor U4812 (N_4812,N_4771,N_4799);
or U4813 (N_4813,N_4704,N_4750);
nand U4814 (N_4814,N_4718,N_4728);
xor U4815 (N_4815,N_4717,N_4759);
nor U4816 (N_4816,N_4725,N_4736);
xor U4817 (N_4817,N_4747,N_4742);
or U4818 (N_4818,N_4765,N_4732);
xor U4819 (N_4819,N_4798,N_4740);
nor U4820 (N_4820,N_4720,N_4775);
nor U4821 (N_4821,N_4794,N_4738);
nor U4822 (N_4822,N_4785,N_4723);
nor U4823 (N_4823,N_4707,N_4741);
nor U4824 (N_4824,N_4716,N_4762);
and U4825 (N_4825,N_4756,N_4795);
nor U4826 (N_4826,N_4797,N_4787);
xnor U4827 (N_4827,N_4790,N_4709);
nor U4828 (N_4828,N_4792,N_4776);
nor U4829 (N_4829,N_4739,N_4703);
nand U4830 (N_4830,N_4769,N_4760);
nor U4831 (N_4831,N_4748,N_4773);
xnor U4832 (N_4832,N_4767,N_4753);
and U4833 (N_4833,N_4700,N_4724);
nand U4834 (N_4834,N_4766,N_4763);
and U4835 (N_4835,N_4734,N_4749);
nand U4836 (N_4836,N_4755,N_4713);
nor U4837 (N_4837,N_4786,N_4719);
and U4838 (N_4838,N_4737,N_4770);
nand U4839 (N_4839,N_4744,N_4774);
and U4840 (N_4840,N_4735,N_4733);
nor U4841 (N_4841,N_4714,N_4712);
nor U4842 (N_4842,N_4752,N_4729);
or U4843 (N_4843,N_4781,N_4757);
nand U4844 (N_4844,N_4710,N_4721);
xor U4845 (N_4845,N_4731,N_4711);
and U4846 (N_4846,N_4796,N_4789);
and U4847 (N_4847,N_4708,N_4702);
nand U4848 (N_4848,N_4758,N_4788);
xnor U4849 (N_4849,N_4768,N_4754);
or U4850 (N_4850,N_4775,N_4755);
or U4851 (N_4851,N_4743,N_4752);
or U4852 (N_4852,N_4765,N_4724);
or U4853 (N_4853,N_4776,N_4783);
and U4854 (N_4854,N_4783,N_4754);
or U4855 (N_4855,N_4707,N_4702);
and U4856 (N_4856,N_4729,N_4784);
nand U4857 (N_4857,N_4720,N_4733);
nor U4858 (N_4858,N_4746,N_4742);
nor U4859 (N_4859,N_4737,N_4728);
and U4860 (N_4860,N_4773,N_4751);
nand U4861 (N_4861,N_4778,N_4788);
or U4862 (N_4862,N_4785,N_4713);
and U4863 (N_4863,N_4729,N_4739);
nor U4864 (N_4864,N_4741,N_4736);
nor U4865 (N_4865,N_4723,N_4782);
or U4866 (N_4866,N_4741,N_4770);
nor U4867 (N_4867,N_4785,N_4756);
nor U4868 (N_4868,N_4721,N_4749);
or U4869 (N_4869,N_4768,N_4777);
or U4870 (N_4870,N_4706,N_4737);
and U4871 (N_4871,N_4702,N_4760);
nor U4872 (N_4872,N_4760,N_4713);
and U4873 (N_4873,N_4787,N_4753);
nand U4874 (N_4874,N_4794,N_4760);
nand U4875 (N_4875,N_4759,N_4730);
nor U4876 (N_4876,N_4721,N_4747);
nand U4877 (N_4877,N_4778,N_4777);
or U4878 (N_4878,N_4788,N_4747);
nand U4879 (N_4879,N_4755,N_4728);
or U4880 (N_4880,N_4709,N_4732);
nor U4881 (N_4881,N_4718,N_4780);
and U4882 (N_4882,N_4786,N_4778);
or U4883 (N_4883,N_4719,N_4712);
or U4884 (N_4884,N_4741,N_4718);
nor U4885 (N_4885,N_4737,N_4791);
and U4886 (N_4886,N_4720,N_4746);
xor U4887 (N_4887,N_4763,N_4721);
nor U4888 (N_4888,N_4725,N_4750);
xnor U4889 (N_4889,N_4750,N_4740);
nor U4890 (N_4890,N_4778,N_4717);
nor U4891 (N_4891,N_4745,N_4702);
or U4892 (N_4892,N_4753,N_4760);
nand U4893 (N_4893,N_4714,N_4735);
or U4894 (N_4894,N_4760,N_4700);
xor U4895 (N_4895,N_4775,N_4759);
or U4896 (N_4896,N_4722,N_4719);
and U4897 (N_4897,N_4799,N_4703);
nand U4898 (N_4898,N_4785,N_4738);
nand U4899 (N_4899,N_4793,N_4773);
xnor U4900 (N_4900,N_4885,N_4888);
or U4901 (N_4901,N_4878,N_4828);
or U4902 (N_4902,N_4887,N_4882);
nand U4903 (N_4903,N_4879,N_4807);
nor U4904 (N_4904,N_4865,N_4831);
or U4905 (N_4905,N_4850,N_4810);
and U4906 (N_4906,N_4894,N_4812);
xnor U4907 (N_4907,N_4881,N_4847);
or U4908 (N_4908,N_4895,N_4832);
or U4909 (N_4909,N_4835,N_4857);
nand U4910 (N_4910,N_4809,N_4815);
nor U4911 (N_4911,N_4822,N_4801);
nand U4912 (N_4912,N_4833,N_4821);
and U4913 (N_4913,N_4873,N_4808);
and U4914 (N_4914,N_4839,N_4870);
nor U4915 (N_4915,N_4859,N_4884);
xor U4916 (N_4916,N_4880,N_4892);
nor U4917 (N_4917,N_4830,N_4875);
nor U4918 (N_4918,N_4846,N_4891);
nor U4919 (N_4919,N_4841,N_4871);
nand U4920 (N_4920,N_4826,N_4823);
or U4921 (N_4921,N_4843,N_4813);
xnor U4922 (N_4922,N_4817,N_4877);
xor U4923 (N_4923,N_4844,N_4800);
nor U4924 (N_4924,N_4890,N_4852);
xnor U4925 (N_4925,N_4849,N_4806);
nand U4926 (N_4926,N_4818,N_4853);
xor U4927 (N_4927,N_4834,N_4862);
or U4928 (N_4928,N_4819,N_4855);
nor U4929 (N_4929,N_4898,N_4886);
nand U4930 (N_4930,N_4840,N_4836);
xnor U4931 (N_4931,N_4854,N_4876);
and U4932 (N_4932,N_4861,N_4805);
and U4933 (N_4933,N_4883,N_4803);
or U4934 (N_4934,N_4868,N_4896);
or U4935 (N_4935,N_4837,N_4811);
nand U4936 (N_4936,N_4820,N_4872);
nor U4937 (N_4937,N_4864,N_4889);
nor U4938 (N_4938,N_4851,N_4863);
nand U4939 (N_4939,N_4856,N_4838);
nand U4940 (N_4940,N_4814,N_4860);
nand U4941 (N_4941,N_4842,N_4897);
nand U4942 (N_4942,N_4804,N_4858);
or U4943 (N_4943,N_4825,N_4829);
nand U4944 (N_4944,N_4824,N_4816);
nand U4945 (N_4945,N_4802,N_4874);
and U4946 (N_4946,N_4893,N_4866);
nand U4947 (N_4947,N_4869,N_4848);
xor U4948 (N_4948,N_4899,N_4867);
nor U4949 (N_4949,N_4827,N_4845);
and U4950 (N_4950,N_4876,N_4812);
nand U4951 (N_4951,N_4839,N_4814);
nor U4952 (N_4952,N_4866,N_4824);
or U4953 (N_4953,N_4802,N_4842);
nor U4954 (N_4954,N_4808,N_4828);
nand U4955 (N_4955,N_4856,N_4821);
xnor U4956 (N_4956,N_4874,N_4862);
or U4957 (N_4957,N_4884,N_4804);
xor U4958 (N_4958,N_4879,N_4877);
nand U4959 (N_4959,N_4830,N_4883);
and U4960 (N_4960,N_4836,N_4825);
and U4961 (N_4961,N_4806,N_4891);
xnor U4962 (N_4962,N_4851,N_4891);
nor U4963 (N_4963,N_4874,N_4857);
nand U4964 (N_4964,N_4804,N_4829);
nand U4965 (N_4965,N_4835,N_4855);
and U4966 (N_4966,N_4853,N_4805);
nor U4967 (N_4967,N_4828,N_4849);
nor U4968 (N_4968,N_4848,N_4889);
nor U4969 (N_4969,N_4811,N_4868);
nor U4970 (N_4970,N_4814,N_4869);
and U4971 (N_4971,N_4831,N_4866);
nor U4972 (N_4972,N_4809,N_4843);
nand U4973 (N_4973,N_4894,N_4820);
xnor U4974 (N_4974,N_4876,N_4877);
and U4975 (N_4975,N_4893,N_4809);
or U4976 (N_4976,N_4833,N_4831);
and U4977 (N_4977,N_4840,N_4897);
and U4978 (N_4978,N_4809,N_4811);
nand U4979 (N_4979,N_4832,N_4868);
nor U4980 (N_4980,N_4816,N_4806);
xor U4981 (N_4981,N_4826,N_4800);
nor U4982 (N_4982,N_4824,N_4807);
nand U4983 (N_4983,N_4837,N_4872);
or U4984 (N_4984,N_4876,N_4862);
nand U4985 (N_4985,N_4879,N_4804);
nor U4986 (N_4986,N_4887,N_4864);
and U4987 (N_4987,N_4893,N_4894);
nor U4988 (N_4988,N_4830,N_4874);
and U4989 (N_4989,N_4898,N_4832);
nand U4990 (N_4990,N_4885,N_4899);
nor U4991 (N_4991,N_4875,N_4857);
or U4992 (N_4992,N_4829,N_4897);
or U4993 (N_4993,N_4823,N_4803);
nor U4994 (N_4994,N_4802,N_4844);
nand U4995 (N_4995,N_4895,N_4898);
or U4996 (N_4996,N_4817,N_4822);
or U4997 (N_4997,N_4853,N_4897);
nand U4998 (N_4998,N_4813,N_4824);
or U4999 (N_4999,N_4891,N_4803);
nor UO_0 (O_0,N_4922,N_4903);
and UO_1 (O_1,N_4982,N_4983);
and UO_2 (O_2,N_4936,N_4999);
or UO_3 (O_3,N_4941,N_4976);
nand UO_4 (O_4,N_4991,N_4997);
nand UO_5 (O_5,N_4933,N_4904);
or UO_6 (O_6,N_4913,N_4908);
or UO_7 (O_7,N_4958,N_4961);
or UO_8 (O_8,N_4964,N_4907);
nor UO_9 (O_9,N_4930,N_4931);
and UO_10 (O_10,N_4902,N_4998);
and UO_11 (O_11,N_4969,N_4995);
xnor UO_12 (O_12,N_4950,N_4945);
or UO_13 (O_13,N_4948,N_4915);
or UO_14 (O_14,N_4914,N_4975);
and UO_15 (O_15,N_4919,N_4910);
nor UO_16 (O_16,N_4909,N_4938);
xor UO_17 (O_17,N_4926,N_4956);
nor UO_18 (O_18,N_4934,N_4925);
nand UO_19 (O_19,N_4921,N_4900);
or UO_20 (O_20,N_4905,N_4949);
nand UO_21 (O_21,N_4953,N_4987);
or UO_22 (O_22,N_4920,N_4960);
and UO_23 (O_23,N_4993,N_4990);
or UO_24 (O_24,N_4988,N_4935);
or UO_25 (O_25,N_4992,N_4974);
nor UO_26 (O_26,N_4937,N_4981);
and UO_27 (O_27,N_4955,N_4972);
or UO_28 (O_28,N_4965,N_4927);
and UO_29 (O_29,N_4951,N_4917);
nand UO_30 (O_30,N_4906,N_4978);
or UO_31 (O_31,N_4943,N_4912);
and UO_32 (O_32,N_4962,N_4947);
nor UO_33 (O_33,N_4973,N_4959);
or UO_34 (O_34,N_4980,N_4952);
xor UO_35 (O_35,N_4911,N_4923);
nor UO_36 (O_36,N_4967,N_4929);
nor UO_37 (O_37,N_4940,N_4994);
xnor UO_38 (O_38,N_4963,N_4977);
and UO_39 (O_39,N_4942,N_4954);
or UO_40 (O_40,N_4939,N_4944);
or UO_41 (O_41,N_4989,N_4985);
and UO_42 (O_42,N_4984,N_4971);
nor UO_43 (O_43,N_4996,N_4957);
nand UO_44 (O_44,N_4901,N_4916);
nand UO_45 (O_45,N_4932,N_4968);
or UO_46 (O_46,N_4924,N_4979);
or UO_47 (O_47,N_4966,N_4946);
nor UO_48 (O_48,N_4928,N_4986);
or UO_49 (O_49,N_4970,N_4918);
nand UO_50 (O_50,N_4940,N_4914);
or UO_51 (O_51,N_4912,N_4994);
nand UO_52 (O_52,N_4924,N_4963);
and UO_53 (O_53,N_4914,N_4915);
nand UO_54 (O_54,N_4951,N_4989);
nand UO_55 (O_55,N_4970,N_4905);
nand UO_56 (O_56,N_4993,N_4999);
nand UO_57 (O_57,N_4976,N_4971);
nand UO_58 (O_58,N_4987,N_4914);
and UO_59 (O_59,N_4973,N_4970);
or UO_60 (O_60,N_4962,N_4914);
and UO_61 (O_61,N_4949,N_4984);
nand UO_62 (O_62,N_4904,N_4994);
xnor UO_63 (O_63,N_4985,N_4916);
nor UO_64 (O_64,N_4987,N_4988);
or UO_65 (O_65,N_4986,N_4930);
nor UO_66 (O_66,N_4912,N_4920);
nand UO_67 (O_67,N_4933,N_4934);
and UO_68 (O_68,N_4900,N_4935);
nor UO_69 (O_69,N_4950,N_4955);
or UO_70 (O_70,N_4959,N_4903);
or UO_71 (O_71,N_4919,N_4970);
and UO_72 (O_72,N_4949,N_4947);
xor UO_73 (O_73,N_4969,N_4963);
nand UO_74 (O_74,N_4945,N_4911);
or UO_75 (O_75,N_4996,N_4978);
nor UO_76 (O_76,N_4968,N_4915);
and UO_77 (O_77,N_4957,N_4910);
and UO_78 (O_78,N_4919,N_4964);
or UO_79 (O_79,N_4996,N_4920);
or UO_80 (O_80,N_4993,N_4909);
nand UO_81 (O_81,N_4984,N_4911);
or UO_82 (O_82,N_4962,N_4907);
nor UO_83 (O_83,N_4991,N_4988);
and UO_84 (O_84,N_4967,N_4997);
or UO_85 (O_85,N_4941,N_4986);
or UO_86 (O_86,N_4956,N_4985);
or UO_87 (O_87,N_4973,N_4960);
nand UO_88 (O_88,N_4927,N_4970);
and UO_89 (O_89,N_4908,N_4960);
nand UO_90 (O_90,N_4954,N_4993);
and UO_91 (O_91,N_4912,N_4988);
and UO_92 (O_92,N_4911,N_4952);
and UO_93 (O_93,N_4905,N_4965);
xor UO_94 (O_94,N_4935,N_4964);
xor UO_95 (O_95,N_4985,N_4991);
nand UO_96 (O_96,N_4921,N_4909);
and UO_97 (O_97,N_4936,N_4938);
or UO_98 (O_98,N_4983,N_4987);
and UO_99 (O_99,N_4943,N_4979);
nor UO_100 (O_100,N_4979,N_4988);
or UO_101 (O_101,N_4909,N_4968);
nor UO_102 (O_102,N_4976,N_4909);
nand UO_103 (O_103,N_4909,N_4900);
and UO_104 (O_104,N_4986,N_4923);
or UO_105 (O_105,N_4991,N_4941);
nand UO_106 (O_106,N_4993,N_4930);
nand UO_107 (O_107,N_4922,N_4954);
and UO_108 (O_108,N_4965,N_4997);
or UO_109 (O_109,N_4991,N_4922);
or UO_110 (O_110,N_4969,N_4983);
or UO_111 (O_111,N_4945,N_4993);
or UO_112 (O_112,N_4977,N_4986);
nand UO_113 (O_113,N_4941,N_4932);
or UO_114 (O_114,N_4973,N_4922);
and UO_115 (O_115,N_4959,N_4915);
nand UO_116 (O_116,N_4987,N_4931);
and UO_117 (O_117,N_4956,N_4935);
or UO_118 (O_118,N_4945,N_4909);
nor UO_119 (O_119,N_4920,N_4913);
xor UO_120 (O_120,N_4997,N_4944);
nand UO_121 (O_121,N_4941,N_4965);
nand UO_122 (O_122,N_4984,N_4951);
or UO_123 (O_123,N_4919,N_4974);
or UO_124 (O_124,N_4950,N_4918);
nand UO_125 (O_125,N_4999,N_4976);
or UO_126 (O_126,N_4904,N_4963);
nor UO_127 (O_127,N_4953,N_4979);
nand UO_128 (O_128,N_4956,N_4907);
nand UO_129 (O_129,N_4907,N_4998);
and UO_130 (O_130,N_4929,N_4984);
nor UO_131 (O_131,N_4950,N_4989);
or UO_132 (O_132,N_4925,N_4955);
and UO_133 (O_133,N_4973,N_4952);
and UO_134 (O_134,N_4922,N_4999);
nor UO_135 (O_135,N_4908,N_4995);
nand UO_136 (O_136,N_4962,N_4943);
xnor UO_137 (O_137,N_4972,N_4940);
xnor UO_138 (O_138,N_4956,N_4927);
nand UO_139 (O_139,N_4936,N_4967);
and UO_140 (O_140,N_4914,N_4964);
or UO_141 (O_141,N_4960,N_4918);
nand UO_142 (O_142,N_4938,N_4960);
nor UO_143 (O_143,N_4941,N_4908);
nand UO_144 (O_144,N_4940,N_4999);
nor UO_145 (O_145,N_4976,N_4924);
and UO_146 (O_146,N_4995,N_4902);
or UO_147 (O_147,N_4928,N_4938);
or UO_148 (O_148,N_4950,N_4906);
xor UO_149 (O_149,N_4935,N_4999);
and UO_150 (O_150,N_4997,N_4906);
nand UO_151 (O_151,N_4962,N_4963);
xnor UO_152 (O_152,N_4944,N_4936);
xnor UO_153 (O_153,N_4972,N_4997);
nor UO_154 (O_154,N_4916,N_4984);
and UO_155 (O_155,N_4982,N_4978);
xor UO_156 (O_156,N_4919,N_4984);
and UO_157 (O_157,N_4958,N_4943);
nor UO_158 (O_158,N_4966,N_4925);
nor UO_159 (O_159,N_4924,N_4943);
nor UO_160 (O_160,N_4924,N_4982);
nor UO_161 (O_161,N_4956,N_4994);
nand UO_162 (O_162,N_4925,N_4974);
and UO_163 (O_163,N_4960,N_4959);
and UO_164 (O_164,N_4925,N_4950);
xor UO_165 (O_165,N_4987,N_4977);
or UO_166 (O_166,N_4925,N_4926);
xor UO_167 (O_167,N_4977,N_4992);
and UO_168 (O_168,N_4987,N_4946);
or UO_169 (O_169,N_4972,N_4979);
nor UO_170 (O_170,N_4918,N_4917);
or UO_171 (O_171,N_4984,N_4975);
nand UO_172 (O_172,N_4970,N_4986);
or UO_173 (O_173,N_4929,N_4987);
xor UO_174 (O_174,N_4954,N_4926);
nor UO_175 (O_175,N_4931,N_4948);
and UO_176 (O_176,N_4928,N_4903);
nand UO_177 (O_177,N_4946,N_4918);
or UO_178 (O_178,N_4947,N_4981);
nor UO_179 (O_179,N_4917,N_4940);
nor UO_180 (O_180,N_4934,N_4949);
nor UO_181 (O_181,N_4996,N_4992);
and UO_182 (O_182,N_4945,N_4973);
or UO_183 (O_183,N_4926,N_4915);
or UO_184 (O_184,N_4961,N_4975);
or UO_185 (O_185,N_4946,N_4906);
xor UO_186 (O_186,N_4942,N_4969);
or UO_187 (O_187,N_4940,N_4931);
nor UO_188 (O_188,N_4920,N_4901);
nand UO_189 (O_189,N_4966,N_4928);
or UO_190 (O_190,N_4935,N_4967);
xor UO_191 (O_191,N_4940,N_4977);
or UO_192 (O_192,N_4908,N_4970);
nand UO_193 (O_193,N_4900,N_4933);
and UO_194 (O_194,N_4909,N_4998);
or UO_195 (O_195,N_4948,N_4921);
nor UO_196 (O_196,N_4927,N_4996);
or UO_197 (O_197,N_4908,N_4950);
and UO_198 (O_198,N_4918,N_4997);
or UO_199 (O_199,N_4934,N_4937);
nand UO_200 (O_200,N_4994,N_4982);
and UO_201 (O_201,N_4953,N_4965);
nand UO_202 (O_202,N_4997,N_4971);
nand UO_203 (O_203,N_4919,N_4936);
nand UO_204 (O_204,N_4955,N_4993);
or UO_205 (O_205,N_4954,N_4997);
nor UO_206 (O_206,N_4999,N_4925);
or UO_207 (O_207,N_4999,N_4961);
and UO_208 (O_208,N_4926,N_4982);
nand UO_209 (O_209,N_4980,N_4911);
nor UO_210 (O_210,N_4901,N_4988);
and UO_211 (O_211,N_4948,N_4963);
and UO_212 (O_212,N_4948,N_4994);
nor UO_213 (O_213,N_4935,N_4978);
and UO_214 (O_214,N_4924,N_4904);
nand UO_215 (O_215,N_4900,N_4964);
or UO_216 (O_216,N_4956,N_4991);
nor UO_217 (O_217,N_4977,N_4954);
xnor UO_218 (O_218,N_4922,N_4998);
nand UO_219 (O_219,N_4931,N_4965);
or UO_220 (O_220,N_4915,N_4925);
nand UO_221 (O_221,N_4968,N_4989);
nand UO_222 (O_222,N_4911,N_4946);
nor UO_223 (O_223,N_4940,N_4969);
nand UO_224 (O_224,N_4988,N_4969);
nor UO_225 (O_225,N_4916,N_4944);
and UO_226 (O_226,N_4902,N_4997);
and UO_227 (O_227,N_4923,N_4975);
and UO_228 (O_228,N_4971,N_4978);
or UO_229 (O_229,N_4907,N_4918);
and UO_230 (O_230,N_4972,N_4948);
nand UO_231 (O_231,N_4995,N_4906);
nor UO_232 (O_232,N_4907,N_4999);
or UO_233 (O_233,N_4960,N_4905);
or UO_234 (O_234,N_4943,N_4959);
nand UO_235 (O_235,N_4967,N_4999);
and UO_236 (O_236,N_4953,N_4958);
or UO_237 (O_237,N_4966,N_4972);
nand UO_238 (O_238,N_4928,N_4958);
or UO_239 (O_239,N_4953,N_4925);
nand UO_240 (O_240,N_4971,N_4948);
nand UO_241 (O_241,N_4924,N_4966);
and UO_242 (O_242,N_4973,N_4932);
nand UO_243 (O_243,N_4981,N_4900);
or UO_244 (O_244,N_4939,N_4966);
or UO_245 (O_245,N_4913,N_4924);
and UO_246 (O_246,N_4930,N_4904);
nand UO_247 (O_247,N_4985,N_4967);
nor UO_248 (O_248,N_4974,N_4987);
and UO_249 (O_249,N_4952,N_4948);
xnor UO_250 (O_250,N_4900,N_4913);
nor UO_251 (O_251,N_4918,N_4948);
nand UO_252 (O_252,N_4995,N_4949);
xnor UO_253 (O_253,N_4937,N_4910);
or UO_254 (O_254,N_4983,N_4923);
nand UO_255 (O_255,N_4985,N_4926);
and UO_256 (O_256,N_4989,N_4992);
nand UO_257 (O_257,N_4976,N_4932);
nor UO_258 (O_258,N_4984,N_4930);
xor UO_259 (O_259,N_4909,N_4980);
and UO_260 (O_260,N_4997,N_4934);
nor UO_261 (O_261,N_4978,N_4979);
xor UO_262 (O_262,N_4923,N_4933);
nand UO_263 (O_263,N_4920,N_4925);
xnor UO_264 (O_264,N_4961,N_4982);
nor UO_265 (O_265,N_4917,N_4946);
or UO_266 (O_266,N_4968,N_4908);
and UO_267 (O_267,N_4962,N_4979);
or UO_268 (O_268,N_4961,N_4969);
or UO_269 (O_269,N_4950,N_4994);
xor UO_270 (O_270,N_4927,N_4964);
nand UO_271 (O_271,N_4990,N_4973);
xnor UO_272 (O_272,N_4995,N_4914);
or UO_273 (O_273,N_4923,N_4954);
and UO_274 (O_274,N_4926,N_4928);
and UO_275 (O_275,N_4949,N_4933);
nor UO_276 (O_276,N_4941,N_4979);
nor UO_277 (O_277,N_4941,N_4906);
nand UO_278 (O_278,N_4911,N_4914);
or UO_279 (O_279,N_4960,N_4946);
nand UO_280 (O_280,N_4943,N_4913);
nand UO_281 (O_281,N_4999,N_4991);
or UO_282 (O_282,N_4904,N_4968);
nor UO_283 (O_283,N_4981,N_4923);
nor UO_284 (O_284,N_4921,N_4957);
nor UO_285 (O_285,N_4943,N_4921);
nor UO_286 (O_286,N_4932,N_4912);
nand UO_287 (O_287,N_4917,N_4938);
nor UO_288 (O_288,N_4997,N_4905);
nor UO_289 (O_289,N_4922,N_4918);
and UO_290 (O_290,N_4931,N_4978);
nor UO_291 (O_291,N_4938,N_4958);
nand UO_292 (O_292,N_4993,N_4924);
or UO_293 (O_293,N_4907,N_4944);
xor UO_294 (O_294,N_4958,N_4917);
nor UO_295 (O_295,N_4916,N_4935);
nor UO_296 (O_296,N_4967,N_4990);
or UO_297 (O_297,N_4954,N_4919);
or UO_298 (O_298,N_4966,N_4933);
and UO_299 (O_299,N_4930,N_4910);
nor UO_300 (O_300,N_4996,N_4919);
or UO_301 (O_301,N_4931,N_4910);
nor UO_302 (O_302,N_4901,N_4925);
or UO_303 (O_303,N_4933,N_4992);
and UO_304 (O_304,N_4961,N_4947);
xnor UO_305 (O_305,N_4958,N_4972);
and UO_306 (O_306,N_4923,N_4939);
nand UO_307 (O_307,N_4945,N_4959);
and UO_308 (O_308,N_4990,N_4953);
nand UO_309 (O_309,N_4989,N_4969);
and UO_310 (O_310,N_4924,N_4970);
nor UO_311 (O_311,N_4953,N_4975);
xor UO_312 (O_312,N_4946,N_4980);
nand UO_313 (O_313,N_4995,N_4970);
or UO_314 (O_314,N_4917,N_4998);
nand UO_315 (O_315,N_4982,N_4997);
and UO_316 (O_316,N_4952,N_4939);
nand UO_317 (O_317,N_4921,N_4961);
or UO_318 (O_318,N_4916,N_4905);
nor UO_319 (O_319,N_4991,N_4911);
nor UO_320 (O_320,N_4910,N_4909);
or UO_321 (O_321,N_4927,N_4953);
nor UO_322 (O_322,N_4952,N_4979);
nor UO_323 (O_323,N_4959,N_4907);
or UO_324 (O_324,N_4996,N_4910);
nand UO_325 (O_325,N_4982,N_4988);
or UO_326 (O_326,N_4960,N_4978);
nor UO_327 (O_327,N_4998,N_4974);
xor UO_328 (O_328,N_4981,N_4975);
and UO_329 (O_329,N_4991,N_4937);
or UO_330 (O_330,N_4960,N_4900);
nand UO_331 (O_331,N_4976,N_4949);
nor UO_332 (O_332,N_4994,N_4990);
and UO_333 (O_333,N_4989,N_4929);
and UO_334 (O_334,N_4998,N_4936);
xor UO_335 (O_335,N_4963,N_4968);
and UO_336 (O_336,N_4979,N_4955);
nand UO_337 (O_337,N_4960,N_4997);
nor UO_338 (O_338,N_4966,N_4951);
or UO_339 (O_339,N_4976,N_4987);
and UO_340 (O_340,N_4902,N_4947);
and UO_341 (O_341,N_4935,N_4992);
nand UO_342 (O_342,N_4996,N_4986);
nand UO_343 (O_343,N_4974,N_4970);
or UO_344 (O_344,N_4941,N_4936);
xor UO_345 (O_345,N_4903,N_4930);
nand UO_346 (O_346,N_4944,N_4983);
nor UO_347 (O_347,N_4947,N_4988);
or UO_348 (O_348,N_4955,N_4942);
and UO_349 (O_349,N_4928,N_4904);
nand UO_350 (O_350,N_4906,N_4999);
nor UO_351 (O_351,N_4958,N_4949);
nand UO_352 (O_352,N_4921,N_4962);
or UO_353 (O_353,N_4985,N_4976);
and UO_354 (O_354,N_4949,N_4982);
xnor UO_355 (O_355,N_4973,N_4992);
or UO_356 (O_356,N_4996,N_4909);
nor UO_357 (O_357,N_4944,N_4925);
nand UO_358 (O_358,N_4987,N_4944);
nand UO_359 (O_359,N_4939,N_4929);
and UO_360 (O_360,N_4916,N_4957);
nand UO_361 (O_361,N_4995,N_4979);
and UO_362 (O_362,N_4920,N_4964);
nor UO_363 (O_363,N_4965,N_4968);
or UO_364 (O_364,N_4903,N_4984);
or UO_365 (O_365,N_4923,N_4908);
nand UO_366 (O_366,N_4983,N_4918);
and UO_367 (O_367,N_4944,N_4982);
nor UO_368 (O_368,N_4909,N_4953);
and UO_369 (O_369,N_4997,N_4935);
nand UO_370 (O_370,N_4926,N_4962);
nand UO_371 (O_371,N_4956,N_4905);
nand UO_372 (O_372,N_4935,N_4926);
nand UO_373 (O_373,N_4905,N_4980);
nor UO_374 (O_374,N_4950,N_4984);
and UO_375 (O_375,N_4907,N_4951);
and UO_376 (O_376,N_4993,N_4958);
nand UO_377 (O_377,N_4996,N_4907);
and UO_378 (O_378,N_4904,N_4927);
and UO_379 (O_379,N_4948,N_4903);
nand UO_380 (O_380,N_4946,N_4995);
nand UO_381 (O_381,N_4997,N_4920);
nand UO_382 (O_382,N_4930,N_4942);
or UO_383 (O_383,N_4943,N_4902);
nand UO_384 (O_384,N_4996,N_4940);
nand UO_385 (O_385,N_4999,N_4903);
nand UO_386 (O_386,N_4900,N_4932);
or UO_387 (O_387,N_4901,N_4973);
and UO_388 (O_388,N_4952,N_4907);
and UO_389 (O_389,N_4945,N_4989);
nor UO_390 (O_390,N_4905,N_4906);
nand UO_391 (O_391,N_4976,N_4950);
nor UO_392 (O_392,N_4912,N_4973);
or UO_393 (O_393,N_4930,N_4972);
or UO_394 (O_394,N_4986,N_4935);
xnor UO_395 (O_395,N_4970,N_4916);
nor UO_396 (O_396,N_4931,N_4990);
or UO_397 (O_397,N_4988,N_4938);
or UO_398 (O_398,N_4912,N_4917);
and UO_399 (O_399,N_4991,N_4907);
xnor UO_400 (O_400,N_4991,N_4949);
or UO_401 (O_401,N_4903,N_4997);
and UO_402 (O_402,N_4934,N_4901);
xor UO_403 (O_403,N_4989,N_4900);
and UO_404 (O_404,N_4960,N_4993);
and UO_405 (O_405,N_4960,N_4924);
or UO_406 (O_406,N_4962,N_4938);
nor UO_407 (O_407,N_4926,N_4940);
nand UO_408 (O_408,N_4996,N_4922);
nor UO_409 (O_409,N_4969,N_4973);
nor UO_410 (O_410,N_4931,N_4949);
nor UO_411 (O_411,N_4920,N_4963);
nand UO_412 (O_412,N_4925,N_4954);
or UO_413 (O_413,N_4903,N_4937);
and UO_414 (O_414,N_4973,N_4944);
nor UO_415 (O_415,N_4918,N_4998);
or UO_416 (O_416,N_4974,N_4939);
or UO_417 (O_417,N_4914,N_4959);
xor UO_418 (O_418,N_4915,N_4987);
or UO_419 (O_419,N_4927,N_4999);
nor UO_420 (O_420,N_4913,N_4994);
xnor UO_421 (O_421,N_4933,N_4901);
nor UO_422 (O_422,N_4967,N_4937);
and UO_423 (O_423,N_4915,N_4916);
or UO_424 (O_424,N_4962,N_4900);
xnor UO_425 (O_425,N_4915,N_4979);
or UO_426 (O_426,N_4938,N_4934);
nor UO_427 (O_427,N_4983,N_4962);
nor UO_428 (O_428,N_4987,N_4955);
nand UO_429 (O_429,N_4904,N_4960);
nand UO_430 (O_430,N_4942,N_4941);
or UO_431 (O_431,N_4940,N_4961);
xnor UO_432 (O_432,N_4976,N_4960);
or UO_433 (O_433,N_4910,N_4904);
or UO_434 (O_434,N_4983,N_4953);
nor UO_435 (O_435,N_4964,N_4929);
nand UO_436 (O_436,N_4945,N_4952);
or UO_437 (O_437,N_4952,N_4988);
nand UO_438 (O_438,N_4950,N_4940);
nand UO_439 (O_439,N_4920,N_4903);
nand UO_440 (O_440,N_4939,N_4945);
nand UO_441 (O_441,N_4998,N_4954);
nor UO_442 (O_442,N_4956,N_4987);
and UO_443 (O_443,N_4947,N_4984);
and UO_444 (O_444,N_4985,N_4908);
nand UO_445 (O_445,N_4981,N_4956);
nand UO_446 (O_446,N_4934,N_4962);
nand UO_447 (O_447,N_4976,N_4969);
nand UO_448 (O_448,N_4958,N_4988);
nand UO_449 (O_449,N_4906,N_4960);
nor UO_450 (O_450,N_4974,N_4969);
xnor UO_451 (O_451,N_4963,N_4955);
xor UO_452 (O_452,N_4994,N_4970);
and UO_453 (O_453,N_4928,N_4976);
xor UO_454 (O_454,N_4992,N_4944);
nor UO_455 (O_455,N_4934,N_4900);
nand UO_456 (O_456,N_4904,N_4983);
nor UO_457 (O_457,N_4971,N_4938);
nor UO_458 (O_458,N_4981,N_4974);
xnor UO_459 (O_459,N_4932,N_4959);
or UO_460 (O_460,N_4924,N_4948);
or UO_461 (O_461,N_4988,N_4955);
and UO_462 (O_462,N_4917,N_4984);
and UO_463 (O_463,N_4967,N_4998);
nor UO_464 (O_464,N_4923,N_4966);
and UO_465 (O_465,N_4959,N_4970);
and UO_466 (O_466,N_4927,N_4974);
xnor UO_467 (O_467,N_4921,N_4904);
nor UO_468 (O_468,N_4905,N_4915);
nand UO_469 (O_469,N_4913,N_4988);
or UO_470 (O_470,N_4980,N_4977);
nor UO_471 (O_471,N_4929,N_4934);
nor UO_472 (O_472,N_4902,N_4930);
or UO_473 (O_473,N_4994,N_4992);
or UO_474 (O_474,N_4904,N_4991);
nor UO_475 (O_475,N_4972,N_4968);
nor UO_476 (O_476,N_4901,N_4991);
nor UO_477 (O_477,N_4963,N_4957);
or UO_478 (O_478,N_4993,N_4947);
and UO_479 (O_479,N_4987,N_4923);
nor UO_480 (O_480,N_4971,N_4906);
nor UO_481 (O_481,N_4940,N_4942);
nor UO_482 (O_482,N_4959,N_4954);
nand UO_483 (O_483,N_4975,N_4957);
xnor UO_484 (O_484,N_4935,N_4976);
and UO_485 (O_485,N_4909,N_4960);
or UO_486 (O_486,N_4971,N_4943);
nand UO_487 (O_487,N_4974,N_4993);
and UO_488 (O_488,N_4956,N_4973);
xnor UO_489 (O_489,N_4927,N_4957);
and UO_490 (O_490,N_4963,N_4951);
nor UO_491 (O_491,N_4978,N_4987);
nor UO_492 (O_492,N_4992,N_4958);
and UO_493 (O_493,N_4985,N_4909);
nor UO_494 (O_494,N_4928,N_4991);
nor UO_495 (O_495,N_4996,N_4912);
nand UO_496 (O_496,N_4921,N_4947);
and UO_497 (O_497,N_4901,N_4902);
nand UO_498 (O_498,N_4966,N_4911);
nand UO_499 (O_499,N_4952,N_4937);
or UO_500 (O_500,N_4987,N_4919);
and UO_501 (O_501,N_4925,N_4971);
or UO_502 (O_502,N_4995,N_4985);
or UO_503 (O_503,N_4996,N_4928);
and UO_504 (O_504,N_4946,N_4976);
or UO_505 (O_505,N_4945,N_4978);
and UO_506 (O_506,N_4916,N_4934);
nor UO_507 (O_507,N_4922,N_4900);
or UO_508 (O_508,N_4971,N_4904);
and UO_509 (O_509,N_4934,N_4975);
nor UO_510 (O_510,N_4952,N_4924);
xnor UO_511 (O_511,N_4937,N_4912);
or UO_512 (O_512,N_4911,N_4998);
nor UO_513 (O_513,N_4903,N_4991);
nor UO_514 (O_514,N_4933,N_4925);
nor UO_515 (O_515,N_4951,N_4990);
and UO_516 (O_516,N_4964,N_4911);
nand UO_517 (O_517,N_4988,N_4964);
nand UO_518 (O_518,N_4964,N_4946);
and UO_519 (O_519,N_4950,N_4968);
nand UO_520 (O_520,N_4989,N_4906);
nand UO_521 (O_521,N_4923,N_4979);
xor UO_522 (O_522,N_4953,N_4928);
and UO_523 (O_523,N_4970,N_4964);
and UO_524 (O_524,N_4975,N_4937);
or UO_525 (O_525,N_4921,N_4940);
xor UO_526 (O_526,N_4992,N_4914);
or UO_527 (O_527,N_4969,N_4992);
xor UO_528 (O_528,N_4991,N_4940);
nand UO_529 (O_529,N_4940,N_4993);
nor UO_530 (O_530,N_4937,N_4962);
and UO_531 (O_531,N_4916,N_4973);
and UO_532 (O_532,N_4994,N_4934);
and UO_533 (O_533,N_4942,N_4987);
or UO_534 (O_534,N_4954,N_4953);
nand UO_535 (O_535,N_4926,N_4973);
or UO_536 (O_536,N_4998,N_4931);
or UO_537 (O_537,N_4968,N_4962);
and UO_538 (O_538,N_4971,N_4982);
or UO_539 (O_539,N_4960,N_4977);
xor UO_540 (O_540,N_4939,N_4912);
xor UO_541 (O_541,N_4950,N_4900);
or UO_542 (O_542,N_4979,N_4910);
xnor UO_543 (O_543,N_4949,N_4996);
nor UO_544 (O_544,N_4996,N_4959);
or UO_545 (O_545,N_4911,N_4956);
nand UO_546 (O_546,N_4982,N_4904);
nor UO_547 (O_547,N_4936,N_4971);
and UO_548 (O_548,N_4934,N_4932);
nor UO_549 (O_549,N_4931,N_4967);
and UO_550 (O_550,N_4952,N_4943);
and UO_551 (O_551,N_4969,N_4953);
xor UO_552 (O_552,N_4905,N_4918);
and UO_553 (O_553,N_4993,N_4976);
or UO_554 (O_554,N_4912,N_4979);
or UO_555 (O_555,N_4986,N_4968);
xnor UO_556 (O_556,N_4948,N_4932);
nor UO_557 (O_557,N_4951,N_4920);
nor UO_558 (O_558,N_4985,N_4975);
or UO_559 (O_559,N_4956,N_4939);
nor UO_560 (O_560,N_4992,N_4981);
xnor UO_561 (O_561,N_4901,N_4962);
nand UO_562 (O_562,N_4941,N_4964);
and UO_563 (O_563,N_4964,N_4939);
and UO_564 (O_564,N_4976,N_4981);
or UO_565 (O_565,N_4908,N_4965);
nand UO_566 (O_566,N_4965,N_4904);
or UO_567 (O_567,N_4978,N_4956);
xor UO_568 (O_568,N_4986,N_4912);
or UO_569 (O_569,N_4903,N_4966);
nor UO_570 (O_570,N_4956,N_4963);
nor UO_571 (O_571,N_4916,N_4945);
nor UO_572 (O_572,N_4921,N_4923);
nor UO_573 (O_573,N_4980,N_4917);
xnor UO_574 (O_574,N_4944,N_4922);
or UO_575 (O_575,N_4966,N_4973);
nand UO_576 (O_576,N_4998,N_4972);
and UO_577 (O_577,N_4978,N_4976);
and UO_578 (O_578,N_4955,N_4976);
nor UO_579 (O_579,N_4986,N_4978);
nand UO_580 (O_580,N_4938,N_4998);
and UO_581 (O_581,N_4976,N_4980);
and UO_582 (O_582,N_4928,N_4930);
or UO_583 (O_583,N_4949,N_4948);
and UO_584 (O_584,N_4990,N_4988);
nand UO_585 (O_585,N_4942,N_4933);
nor UO_586 (O_586,N_4999,N_4941);
and UO_587 (O_587,N_4901,N_4911);
nor UO_588 (O_588,N_4907,N_4916);
or UO_589 (O_589,N_4914,N_4967);
or UO_590 (O_590,N_4977,N_4969);
nand UO_591 (O_591,N_4983,N_4912);
nand UO_592 (O_592,N_4944,N_4905);
nand UO_593 (O_593,N_4937,N_4918);
or UO_594 (O_594,N_4974,N_4932);
or UO_595 (O_595,N_4922,N_4912);
and UO_596 (O_596,N_4937,N_4913);
and UO_597 (O_597,N_4948,N_4913);
xor UO_598 (O_598,N_4923,N_4909);
nor UO_599 (O_599,N_4964,N_4985);
nor UO_600 (O_600,N_4941,N_4905);
nor UO_601 (O_601,N_4904,N_4993);
nand UO_602 (O_602,N_4946,N_4956);
xnor UO_603 (O_603,N_4986,N_4937);
nand UO_604 (O_604,N_4950,N_4957);
nor UO_605 (O_605,N_4971,N_4918);
nor UO_606 (O_606,N_4983,N_4999);
and UO_607 (O_607,N_4909,N_4925);
nand UO_608 (O_608,N_4984,N_4908);
and UO_609 (O_609,N_4948,N_4985);
nand UO_610 (O_610,N_4932,N_4906);
xnor UO_611 (O_611,N_4959,N_4984);
nor UO_612 (O_612,N_4901,N_4903);
or UO_613 (O_613,N_4959,N_4909);
nor UO_614 (O_614,N_4915,N_4902);
and UO_615 (O_615,N_4997,N_4978);
and UO_616 (O_616,N_4933,N_4920);
nand UO_617 (O_617,N_4941,N_4920);
nand UO_618 (O_618,N_4960,N_4922);
xor UO_619 (O_619,N_4956,N_4920);
or UO_620 (O_620,N_4935,N_4991);
and UO_621 (O_621,N_4948,N_4916);
and UO_622 (O_622,N_4900,N_4993);
nor UO_623 (O_623,N_4995,N_4950);
nor UO_624 (O_624,N_4950,N_4985);
nor UO_625 (O_625,N_4994,N_4993);
and UO_626 (O_626,N_4963,N_4919);
and UO_627 (O_627,N_4954,N_4931);
or UO_628 (O_628,N_4998,N_4977);
xor UO_629 (O_629,N_4981,N_4941);
xnor UO_630 (O_630,N_4993,N_4922);
nand UO_631 (O_631,N_4996,N_4952);
and UO_632 (O_632,N_4949,N_4961);
xor UO_633 (O_633,N_4942,N_4964);
and UO_634 (O_634,N_4904,N_4986);
nor UO_635 (O_635,N_4916,N_4969);
xor UO_636 (O_636,N_4908,N_4951);
or UO_637 (O_637,N_4986,N_4967);
and UO_638 (O_638,N_4976,N_4966);
and UO_639 (O_639,N_4997,N_4936);
and UO_640 (O_640,N_4980,N_4945);
or UO_641 (O_641,N_4958,N_4935);
and UO_642 (O_642,N_4929,N_4941);
nor UO_643 (O_643,N_4964,N_4959);
or UO_644 (O_644,N_4942,N_4919);
nor UO_645 (O_645,N_4971,N_4910);
nor UO_646 (O_646,N_4946,N_4970);
and UO_647 (O_647,N_4913,N_4976);
xnor UO_648 (O_648,N_4920,N_4977);
nand UO_649 (O_649,N_4976,N_4919);
nand UO_650 (O_650,N_4977,N_4922);
nand UO_651 (O_651,N_4911,N_4947);
nor UO_652 (O_652,N_4966,N_4908);
nand UO_653 (O_653,N_4964,N_4967);
or UO_654 (O_654,N_4998,N_4997);
or UO_655 (O_655,N_4957,N_4937);
and UO_656 (O_656,N_4990,N_4950);
nand UO_657 (O_657,N_4918,N_4947);
nor UO_658 (O_658,N_4911,N_4961);
nand UO_659 (O_659,N_4953,N_4939);
nor UO_660 (O_660,N_4972,N_4937);
or UO_661 (O_661,N_4982,N_4907);
xnor UO_662 (O_662,N_4933,N_4999);
xnor UO_663 (O_663,N_4953,N_4915);
nor UO_664 (O_664,N_4964,N_4923);
and UO_665 (O_665,N_4970,N_4921);
nand UO_666 (O_666,N_4980,N_4983);
nor UO_667 (O_667,N_4991,N_4947);
nor UO_668 (O_668,N_4991,N_4954);
nor UO_669 (O_669,N_4908,N_4914);
and UO_670 (O_670,N_4918,N_4916);
nand UO_671 (O_671,N_4990,N_4995);
nand UO_672 (O_672,N_4946,N_4934);
and UO_673 (O_673,N_4944,N_4920);
and UO_674 (O_674,N_4954,N_4929);
or UO_675 (O_675,N_4960,N_4949);
nand UO_676 (O_676,N_4910,N_4984);
and UO_677 (O_677,N_4958,N_4914);
nand UO_678 (O_678,N_4949,N_4929);
nand UO_679 (O_679,N_4990,N_4935);
or UO_680 (O_680,N_4930,N_4960);
xor UO_681 (O_681,N_4968,N_4942);
nor UO_682 (O_682,N_4922,N_4941);
or UO_683 (O_683,N_4953,N_4945);
nand UO_684 (O_684,N_4988,N_4921);
xnor UO_685 (O_685,N_4932,N_4926);
nor UO_686 (O_686,N_4967,N_4924);
nand UO_687 (O_687,N_4928,N_4912);
nand UO_688 (O_688,N_4900,N_4982);
nor UO_689 (O_689,N_4948,N_4979);
or UO_690 (O_690,N_4988,N_4911);
nand UO_691 (O_691,N_4993,N_4963);
nor UO_692 (O_692,N_4965,N_4917);
nor UO_693 (O_693,N_4980,N_4924);
nor UO_694 (O_694,N_4917,N_4925);
and UO_695 (O_695,N_4915,N_4969);
and UO_696 (O_696,N_4999,N_4985);
nor UO_697 (O_697,N_4967,N_4955);
nor UO_698 (O_698,N_4954,N_4967);
xor UO_699 (O_699,N_4962,N_4977);
nand UO_700 (O_700,N_4937,N_4998);
nor UO_701 (O_701,N_4983,N_4973);
or UO_702 (O_702,N_4913,N_4958);
nand UO_703 (O_703,N_4993,N_4933);
nand UO_704 (O_704,N_4984,N_4926);
nand UO_705 (O_705,N_4980,N_4942);
and UO_706 (O_706,N_4948,N_4942);
nand UO_707 (O_707,N_4943,N_4946);
nor UO_708 (O_708,N_4958,N_4965);
nor UO_709 (O_709,N_4969,N_4993);
nor UO_710 (O_710,N_4945,N_4965);
nor UO_711 (O_711,N_4935,N_4929);
xor UO_712 (O_712,N_4975,N_4972);
nor UO_713 (O_713,N_4959,N_4967);
and UO_714 (O_714,N_4959,N_4908);
nand UO_715 (O_715,N_4968,N_4941);
nand UO_716 (O_716,N_4993,N_4973);
xnor UO_717 (O_717,N_4951,N_4910);
nand UO_718 (O_718,N_4987,N_4925);
or UO_719 (O_719,N_4961,N_4965);
nor UO_720 (O_720,N_4931,N_4988);
nor UO_721 (O_721,N_4937,N_4932);
nand UO_722 (O_722,N_4917,N_4927);
nor UO_723 (O_723,N_4938,N_4990);
or UO_724 (O_724,N_4916,N_4910);
nand UO_725 (O_725,N_4940,N_4904);
xnor UO_726 (O_726,N_4931,N_4915);
nor UO_727 (O_727,N_4910,N_4997);
nand UO_728 (O_728,N_4925,N_4900);
and UO_729 (O_729,N_4927,N_4906);
nand UO_730 (O_730,N_4934,N_4970);
nor UO_731 (O_731,N_4937,N_4907);
nor UO_732 (O_732,N_4938,N_4902);
and UO_733 (O_733,N_4982,N_4918);
nand UO_734 (O_734,N_4999,N_4958);
nand UO_735 (O_735,N_4991,N_4951);
or UO_736 (O_736,N_4941,N_4997);
nand UO_737 (O_737,N_4989,N_4948);
xor UO_738 (O_738,N_4909,N_4978);
and UO_739 (O_739,N_4913,N_4930);
xnor UO_740 (O_740,N_4950,N_4956);
nand UO_741 (O_741,N_4904,N_4975);
or UO_742 (O_742,N_4959,N_4927);
nand UO_743 (O_743,N_4993,N_4939);
and UO_744 (O_744,N_4954,N_4928);
nand UO_745 (O_745,N_4908,N_4915);
nand UO_746 (O_746,N_4937,N_4948);
nand UO_747 (O_747,N_4905,N_4919);
or UO_748 (O_748,N_4916,N_4980);
nand UO_749 (O_749,N_4927,N_4986);
nand UO_750 (O_750,N_4994,N_4915);
nor UO_751 (O_751,N_4966,N_4961);
nor UO_752 (O_752,N_4983,N_4949);
xor UO_753 (O_753,N_4982,N_4956);
nor UO_754 (O_754,N_4939,N_4975);
nor UO_755 (O_755,N_4976,N_4923);
or UO_756 (O_756,N_4998,N_4975);
or UO_757 (O_757,N_4957,N_4989);
or UO_758 (O_758,N_4957,N_4959);
nand UO_759 (O_759,N_4973,N_4991);
xor UO_760 (O_760,N_4901,N_4908);
nand UO_761 (O_761,N_4984,N_4945);
nand UO_762 (O_762,N_4952,N_4961);
nand UO_763 (O_763,N_4943,N_4968);
nand UO_764 (O_764,N_4960,N_4948);
or UO_765 (O_765,N_4975,N_4968);
and UO_766 (O_766,N_4993,N_4970);
or UO_767 (O_767,N_4997,N_4990);
xnor UO_768 (O_768,N_4976,N_4973);
nand UO_769 (O_769,N_4948,N_4976);
nand UO_770 (O_770,N_4917,N_4952);
nor UO_771 (O_771,N_4912,N_4985);
nand UO_772 (O_772,N_4916,N_4921);
nand UO_773 (O_773,N_4949,N_4972);
nand UO_774 (O_774,N_4915,N_4974);
and UO_775 (O_775,N_4977,N_4955);
and UO_776 (O_776,N_4982,N_4970);
and UO_777 (O_777,N_4933,N_4954);
or UO_778 (O_778,N_4963,N_4997);
nand UO_779 (O_779,N_4968,N_4959);
nor UO_780 (O_780,N_4927,N_4947);
or UO_781 (O_781,N_4965,N_4977);
and UO_782 (O_782,N_4944,N_4994);
and UO_783 (O_783,N_4954,N_4979);
nand UO_784 (O_784,N_4910,N_4958);
nor UO_785 (O_785,N_4968,N_4960);
and UO_786 (O_786,N_4965,N_4939);
nand UO_787 (O_787,N_4980,N_4912);
nor UO_788 (O_788,N_4930,N_4947);
nor UO_789 (O_789,N_4934,N_4978);
nand UO_790 (O_790,N_4938,N_4972);
nand UO_791 (O_791,N_4952,N_4926);
xnor UO_792 (O_792,N_4918,N_4910);
or UO_793 (O_793,N_4952,N_4940);
or UO_794 (O_794,N_4984,N_4964);
nor UO_795 (O_795,N_4937,N_4974);
nor UO_796 (O_796,N_4977,N_4918);
and UO_797 (O_797,N_4986,N_4966);
nand UO_798 (O_798,N_4923,N_4937);
and UO_799 (O_799,N_4921,N_4907);
nor UO_800 (O_800,N_4914,N_4923);
nor UO_801 (O_801,N_4960,N_4929);
and UO_802 (O_802,N_4925,N_4949);
nor UO_803 (O_803,N_4952,N_4983);
xor UO_804 (O_804,N_4962,N_4952);
or UO_805 (O_805,N_4944,N_4962);
or UO_806 (O_806,N_4934,N_4903);
nand UO_807 (O_807,N_4935,N_4947);
or UO_808 (O_808,N_4963,N_4985);
or UO_809 (O_809,N_4930,N_4961);
or UO_810 (O_810,N_4902,N_4925);
nor UO_811 (O_811,N_4910,N_4969);
and UO_812 (O_812,N_4925,N_4960);
and UO_813 (O_813,N_4956,N_4922);
nor UO_814 (O_814,N_4972,N_4918);
nor UO_815 (O_815,N_4959,N_4918);
nand UO_816 (O_816,N_4953,N_4940);
nor UO_817 (O_817,N_4970,N_4983);
and UO_818 (O_818,N_4917,N_4972);
or UO_819 (O_819,N_4990,N_4930);
and UO_820 (O_820,N_4996,N_4926);
nor UO_821 (O_821,N_4950,N_4928);
and UO_822 (O_822,N_4971,N_4940);
and UO_823 (O_823,N_4954,N_4963);
or UO_824 (O_824,N_4994,N_4946);
or UO_825 (O_825,N_4930,N_4963);
nand UO_826 (O_826,N_4961,N_4935);
and UO_827 (O_827,N_4918,N_4929);
or UO_828 (O_828,N_4972,N_4902);
and UO_829 (O_829,N_4990,N_4958);
nor UO_830 (O_830,N_4972,N_4912);
or UO_831 (O_831,N_4935,N_4981);
nand UO_832 (O_832,N_4931,N_4912);
xor UO_833 (O_833,N_4967,N_4994);
nor UO_834 (O_834,N_4936,N_4993);
or UO_835 (O_835,N_4925,N_4924);
xor UO_836 (O_836,N_4934,N_4910);
or UO_837 (O_837,N_4974,N_4908);
nor UO_838 (O_838,N_4956,N_4993);
and UO_839 (O_839,N_4950,N_4923);
nor UO_840 (O_840,N_4927,N_4934);
or UO_841 (O_841,N_4931,N_4986);
nand UO_842 (O_842,N_4926,N_4927);
nor UO_843 (O_843,N_4983,N_4957);
xor UO_844 (O_844,N_4900,N_4924);
nor UO_845 (O_845,N_4926,N_4976);
nor UO_846 (O_846,N_4927,N_4951);
xor UO_847 (O_847,N_4971,N_4903);
nor UO_848 (O_848,N_4979,N_4994);
nor UO_849 (O_849,N_4919,N_4944);
nor UO_850 (O_850,N_4994,N_4921);
or UO_851 (O_851,N_4981,N_4985);
or UO_852 (O_852,N_4964,N_4973);
xnor UO_853 (O_853,N_4916,N_4979);
xor UO_854 (O_854,N_4976,N_4945);
nand UO_855 (O_855,N_4946,N_4908);
nor UO_856 (O_856,N_4925,N_4906);
or UO_857 (O_857,N_4969,N_4929);
xnor UO_858 (O_858,N_4946,N_4942);
nand UO_859 (O_859,N_4980,N_4991);
xor UO_860 (O_860,N_4933,N_4939);
and UO_861 (O_861,N_4975,N_4941);
nor UO_862 (O_862,N_4904,N_4969);
nor UO_863 (O_863,N_4923,N_4945);
nand UO_864 (O_864,N_4984,N_4979);
nand UO_865 (O_865,N_4949,N_4968);
and UO_866 (O_866,N_4914,N_4996);
and UO_867 (O_867,N_4908,N_4936);
or UO_868 (O_868,N_4931,N_4905);
nor UO_869 (O_869,N_4941,N_4917);
nand UO_870 (O_870,N_4927,N_4913);
nand UO_871 (O_871,N_4988,N_4932);
and UO_872 (O_872,N_4938,N_4943);
nand UO_873 (O_873,N_4939,N_4960);
nor UO_874 (O_874,N_4940,N_4948);
nand UO_875 (O_875,N_4998,N_4919);
nand UO_876 (O_876,N_4942,N_4906);
or UO_877 (O_877,N_4972,N_4923);
or UO_878 (O_878,N_4989,N_4958);
and UO_879 (O_879,N_4953,N_4977);
nor UO_880 (O_880,N_4990,N_4929);
nor UO_881 (O_881,N_4952,N_4987);
xnor UO_882 (O_882,N_4914,N_4989);
nand UO_883 (O_883,N_4961,N_4979);
xnor UO_884 (O_884,N_4977,N_4973);
or UO_885 (O_885,N_4993,N_4991);
or UO_886 (O_886,N_4967,N_4946);
or UO_887 (O_887,N_4944,N_4901);
or UO_888 (O_888,N_4975,N_4900);
or UO_889 (O_889,N_4915,N_4947);
or UO_890 (O_890,N_4920,N_4949);
xor UO_891 (O_891,N_4954,N_4957);
or UO_892 (O_892,N_4992,N_4922);
or UO_893 (O_893,N_4967,N_4995);
and UO_894 (O_894,N_4984,N_4992);
xor UO_895 (O_895,N_4917,N_4908);
xnor UO_896 (O_896,N_4967,N_4965);
nand UO_897 (O_897,N_4962,N_4915);
and UO_898 (O_898,N_4954,N_4940);
nor UO_899 (O_899,N_4967,N_4930);
nor UO_900 (O_900,N_4980,N_4963);
or UO_901 (O_901,N_4966,N_4921);
nand UO_902 (O_902,N_4951,N_4964);
nor UO_903 (O_903,N_4953,N_4995);
xor UO_904 (O_904,N_4947,N_4983);
or UO_905 (O_905,N_4989,N_4984);
nor UO_906 (O_906,N_4938,N_4935);
or UO_907 (O_907,N_4958,N_4930);
and UO_908 (O_908,N_4930,N_4997);
and UO_909 (O_909,N_4990,N_4952);
nand UO_910 (O_910,N_4960,N_4990);
nor UO_911 (O_911,N_4982,N_4967);
nand UO_912 (O_912,N_4983,N_4979);
or UO_913 (O_913,N_4990,N_4902);
nand UO_914 (O_914,N_4990,N_4981);
and UO_915 (O_915,N_4927,N_4990);
or UO_916 (O_916,N_4978,N_4905);
and UO_917 (O_917,N_4969,N_4925);
and UO_918 (O_918,N_4948,N_4973);
nor UO_919 (O_919,N_4943,N_4992);
nand UO_920 (O_920,N_4936,N_4984);
nand UO_921 (O_921,N_4964,N_4934);
or UO_922 (O_922,N_4947,N_4939);
nor UO_923 (O_923,N_4971,N_4965);
nor UO_924 (O_924,N_4955,N_4931);
or UO_925 (O_925,N_4922,N_4963);
and UO_926 (O_926,N_4907,N_4932);
nor UO_927 (O_927,N_4989,N_4976);
nand UO_928 (O_928,N_4907,N_4928);
or UO_929 (O_929,N_4906,N_4980);
nand UO_930 (O_930,N_4935,N_4950);
nand UO_931 (O_931,N_4962,N_4956);
and UO_932 (O_932,N_4979,N_4991);
or UO_933 (O_933,N_4955,N_4954);
xor UO_934 (O_934,N_4907,N_4989);
nor UO_935 (O_935,N_4936,N_4915);
and UO_936 (O_936,N_4975,N_4922);
nand UO_937 (O_937,N_4973,N_4961);
and UO_938 (O_938,N_4937,N_4919);
xnor UO_939 (O_939,N_4906,N_4953);
nand UO_940 (O_940,N_4949,N_4903);
xor UO_941 (O_941,N_4962,N_4996);
or UO_942 (O_942,N_4929,N_4919);
and UO_943 (O_943,N_4908,N_4916);
or UO_944 (O_944,N_4917,N_4920);
xnor UO_945 (O_945,N_4950,N_4907);
and UO_946 (O_946,N_4940,N_4933);
and UO_947 (O_947,N_4950,N_4922);
nand UO_948 (O_948,N_4929,N_4985);
nor UO_949 (O_949,N_4955,N_4927);
or UO_950 (O_950,N_4933,N_4955);
or UO_951 (O_951,N_4928,N_4908);
and UO_952 (O_952,N_4981,N_4918);
nand UO_953 (O_953,N_4944,N_4937);
and UO_954 (O_954,N_4913,N_4960);
and UO_955 (O_955,N_4968,N_4974);
and UO_956 (O_956,N_4909,N_4957);
nor UO_957 (O_957,N_4994,N_4963);
nand UO_958 (O_958,N_4962,N_4964);
or UO_959 (O_959,N_4962,N_4939);
or UO_960 (O_960,N_4954,N_4987);
nor UO_961 (O_961,N_4967,N_4927);
nand UO_962 (O_962,N_4948,N_4922);
nor UO_963 (O_963,N_4988,N_4981);
xnor UO_964 (O_964,N_4952,N_4981);
and UO_965 (O_965,N_4901,N_4919);
nand UO_966 (O_966,N_4941,N_4938);
xnor UO_967 (O_967,N_4968,N_4957);
or UO_968 (O_968,N_4905,N_4908);
nand UO_969 (O_969,N_4919,N_4952);
xnor UO_970 (O_970,N_4994,N_4983);
nand UO_971 (O_971,N_4905,N_4929);
nor UO_972 (O_972,N_4925,N_4918);
xnor UO_973 (O_973,N_4909,N_4943);
nor UO_974 (O_974,N_4943,N_4933);
and UO_975 (O_975,N_4970,N_4996);
or UO_976 (O_976,N_4904,N_4985);
nand UO_977 (O_977,N_4937,N_4961);
or UO_978 (O_978,N_4920,N_4979);
or UO_979 (O_979,N_4907,N_4980);
nor UO_980 (O_980,N_4967,N_4960);
or UO_981 (O_981,N_4962,N_4932);
nand UO_982 (O_982,N_4907,N_4973);
or UO_983 (O_983,N_4988,N_4906);
and UO_984 (O_984,N_4964,N_4925);
and UO_985 (O_985,N_4949,N_4910);
nand UO_986 (O_986,N_4928,N_4960);
or UO_987 (O_987,N_4911,N_4916);
nor UO_988 (O_988,N_4985,N_4993);
nor UO_989 (O_989,N_4975,N_4988);
nor UO_990 (O_990,N_4942,N_4934);
nand UO_991 (O_991,N_4967,N_4941);
nor UO_992 (O_992,N_4954,N_4956);
and UO_993 (O_993,N_4952,N_4992);
nand UO_994 (O_994,N_4963,N_4983);
nor UO_995 (O_995,N_4911,N_4977);
xnor UO_996 (O_996,N_4921,N_4928);
nand UO_997 (O_997,N_4921,N_4927);
or UO_998 (O_998,N_4926,N_4955);
nand UO_999 (O_999,N_4953,N_4918);
endmodule