module basic_2500_25000_3000_4_levels_10xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18791,N_18792,N_18793,N_18795,N_18796,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19348,N_19350,N_19351,N_19352,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19409,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19456,N_19458,N_19459,N_19460,N_19461,N_19462,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19570,N_19571,N_19572,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19612,N_19613,N_19614,N_19615,N_19616,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19765,N_19766,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19878,N_19879,N_19880,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19990,N_19991,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20255,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20638,N_20639,N_20640,N_20641,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20704,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20837,N_20838,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20939,N_20940,N_20941,N_20942,N_20943,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20968,N_20969,N_20970,N_20971,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22073,N_22075,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22243,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22266,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22884,N_22886,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23151,N_23152,N_23153,N_23154,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23163,N_23164,N_23165,N_23166,N_23167,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23386,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23397,N_23398,N_23399,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23451,N_23452,N_23453,N_23454,N_23455,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23524,N_23525,N_23526,N_23529,N_23530,N_23531,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23663,N_23664,N_23665,N_23666,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24189,N_24190,N_24191,N_24192,N_24193,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24227,N_24228,N_24229,N_24231,N_24232,N_24233,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24450,N_24451,N_24452,N_24453,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24526,N_24527,N_24528,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24595,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24830,N_24831,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
nor U0 (N_0,In_2167,In_1629);
nand U1 (N_1,In_277,In_1633);
or U2 (N_2,In_529,In_553);
nor U3 (N_3,In_542,In_1434);
or U4 (N_4,In_2078,In_1285);
nor U5 (N_5,In_49,In_488);
nand U6 (N_6,In_1335,In_84);
xor U7 (N_7,In_308,In_1523);
or U8 (N_8,In_1910,In_1982);
or U9 (N_9,In_325,In_2129);
nand U10 (N_10,In_297,In_501);
or U11 (N_11,In_2401,In_919);
xor U12 (N_12,In_988,In_1121);
xor U13 (N_13,In_285,In_1256);
nor U14 (N_14,In_2337,In_268);
nor U15 (N_15,In_579,In_1677);
nor U16 (N_16,In_2189,In_651);
nor U17 (N_17,In_143,In_1004);
or U18 (N_18,In_1291,In_332);
nand U19 (N_19,In_1811,In_54);
or U20 (N_20,In_1708,In_1003);
or U21 (N_21,In_2320,In_2289);
and U22 (N_22,In_371,In_18);
nor U23 (N_23,In_1372,In_992);
xor U24 (N_24,In_2229,In_1337);
xnor U25 (N_25,In_2066,In_2334);
and U26 (N_26,In_2427,In_342);
nor U27 (N_27,In_2236,In_1338);
nand U28 (N_28,In_1565,In_892);
or U29 (N_29,In_961,In_215);
xor U30 (N_30,In_203,In_964);
nor U31 (N_31,In_1240,In_2291);
nand U32 (N_32,In_1119,In_2110);
nand U33 (N_33,In_2330,In_1018);
and U34 (N_34,In_798,In_2365);
nor U35 (N_35,In_1689,In_7);
or U36 (N_36,In_2484,In_1414);
or U37 (N_37,In_686,In_408);
nand U38 (N_38,In_594,In_814);
or U39 (N_39,In_2234,In_2059);
nand U40 (N_40,In_2125,In_924);
nor U41 (N_41,In_345,In_1459);
and U42 (N_42,In_1660,In_106);
nand U43 (N_43,In_2079,In_618);
or U44 (N_44,In_1485,In_741);
and U45 (N_45,In_469,In_2016);
or U46 (N_46,In_978,In_44);
or U47 (N_47,In_101,In_2475);
nand U48 (N_48,In_1248,In_2428);
or U49 (N_49,In_104,In_1635);
xor U50 (N_50,In_989,In_1996);
or U51 (N_51,In_2028,In_1552);
nor U52 (N_52,In_74,In_53);
xor U53 (N_53,In_2213,In_1581);
xor U54 (N_54,In_1894,In_1957);
nor U55 (N_55,In_421,In_1024);
or U56 (N_56,In_167,In_1508);
or U57 (N_57,In_1012,In_827);
and U58 (N_58,In_129,In_2457);
or U59 (N_59,In_2172,In_1199);
nor U60 (N_60,In_677,In_1695);
nor U61 (N_61,In_1649,In_2317);
or U62 (N_62,In_2239,In_1593);
xor U63 (N_63,In_657,In_326);
nand U64 (N_64,In_1662,In_728);
nand U65 (N_65,In_874,In_1317);
and U66 (N_66,In_770,In_492);
nand U67 (N_67,In_1318,In_619);
and U68 (N_68,In_1916,In_2178);
and U69 (N_69,In_1229,In_710);
nand U70 (N_70,In_1504,In_2177);
xor U71 (N_71,In_2212,In_957);
nor U72 (N_72,In_1682,In_890);
and U73 (N_73,In_687,In_969);
or U74 (N_74,In_1930,In_2131);
nor U75 (N_75,In_1223,In_1102);
xnor U76 (N_76,In_1895,In_720);
and U77 (N_77,In_170,In_506);
nand U78 (N_78,In_438,In_1439);
or U79 (N_79,In_2262,In_2254);
xnor U80 (N_80,In_416,In_394);
nor U81 (N_81,In_1650,In_1652);
xor U82 (N_82,In_29,In_478);
and U83 (N_83,In_2490,In_1070);
nand U84 (N_84,In_1819,In_854);
or U85 (N_85,In_1539,In_468);
nand U86 (N_86,In_2116,In_1106);
nand U87 (N_87,In_731,In_1701);
xnor U88 (N_88,In_580,In_562);
xnor U89 (N_89,In_2366,In_1661);
nand U90 (N_90,In_1261,In_1901);
nor U91 (N_91,In_25,In_43);
nand U92 (N_92,In_2030,In_664);
nor U93 (N_93,In_665,In_1554);
and U94 (N_94,In_1158,In_2286);
and U95 (N_95,In_292,In_337);
nor U96 (N_96,In_2064,In_2048);
nand U97 (N_97,In_935,In_1688);
nand U98 (N_98,In_1623,In_191);
xnor U99 (N_99,In_1950,In_251);
or U100 (N_100,In_682,In_1495);
nand U101 (N_101,In_1812,In_637);
or U102 (N_102,In_2150,In_2235);
nand U103 (N_103,In_2308,In_1553);
and U104 (N_104,In_109,In_1050);
and U105 (N_105,In_1540,In_2082);
nand U106 (N_106,In_913,In_1309);
xnor U107 (N_107,In_2447,In_1207);
nand U108 (N_108,In_206,In_1191);
or U109 (N_109,In_333,In_2070);
xnor U110 (N_110,In_1541,In_2029);
nor U111 (N_111,In_70,In_863);
or U112 (N_112,In_1983,In_1155);
xnor U113 (N_113,In_749,In_1000);
and U114 (N_114,In_458,In_1469);
nor U115 (N_115,In_914,In_771);
and U116 (N_116,In_2441,In_1943);
or U117 (N_117,In_275,In_1900);
xnor U118 (N_118,In_2203,In_1296);
and U119 (N_119,In_320,In_633);
and U120 (N_120,In_1783,In_64);
nand U121 (N_121,In_0,In_1888);
nor U122 (N_122,In_952,In_1039);
xnor U123 (N_123,In_1374,In_1858);
and U124 (N_124,In_1678,In_1952);
nor U125 (N_125,In_1923,In_1690);
xor U126 (N_126,In_647,In_703);
xnor U127 (N_127,In_62,In_641);
xnor U128 (N_128,In_2223,In_330);
nor U129 (N_129,In_689,In_464);
xor U130 (N_130,In_733,In_395);
nor U131 (N_131,In_716,In_1966);
and U132 (N_132,In_397,In_1700);
and U133 (N_133,In_2329,In_1714);
nand U134 (N_134,In_213,In_1879);
nor U135 (N_135,In_323,In_1319);
xnor U136 (N_136,In_183,In_1630);
and U137 (N_137,In_462,In_410);
nand U138 (N_138,In_773,In_937);
nor U139 (N_139,In_2080,In_1043);
nor U140 (N_140,In_2423,In_1839);
nor U141 (N_141,In_2180,In_552);
nand U142 (N_142,In_893,In_42);
nand U143 (N_143,In_1235,In_1809);
nand U144 (N_144,In_487,In_1236);
nand U145 (N_145,In_2268,In_1073);
nor U146 (N_146,In_1233,In_1842);
xor U147 (N_147,In_1594,In_1878);
or U148 (N_148,In_2250,In_1245);
nand U149 (N_149,In_2220,In_2311);
nor U150 (N_150,In_356,In_638);
xnor U151 (N_151,In_1868,In_1692);
and U152 (N_152,In_910,In_931);
nand U153 (N_153,In_1873,In_2073);
and U154 (N_154,In_1150,In_1186);
xnor U155 (N_155,In_1090,In_1549);
or U156 (N_156,In_1383,In_1333);
or U157 (N_157,In_1611,In_1767);
and U158 (N_158,In_1215,In_746);
and U159 (N_159,In_790,In_176);
or U160 (N_160,In_936,In_584);
xor U161 (N_161,In_963,In_1848);
nor U162 (N_162,In_2335,In_1250);
or U163 (N_163,In_1672,In_2394);
or U164 (N_164,In_2202,In_1417);
or U165 (N_165,In_2256,In_169);
xnor U166 (N_166,In_1258,In_1411);
nand U167 (N_167,In_12,In_1620);
xor U168 (N_168,In_1307,In_2276);
or U169 (N_169,In_670,In_1449);
and U170 (N_170,In_1711,In_157);
nand U171 (N_171,In_1359,In_219);
nand U172 (N_172,In_1356,In_1008);
nand U173 (N_173,In_712,In_627);
nor U174 (N_174,In_968,In_1889);
nor U175 (N_175,In_1755,In_2032);
xnor U176 (N_176,In_1136,In_583);
xor U177 (N_177,In_2010,In_1213);
xnor U178 (N_178,In_2410,In_862);
and U179 (N_179,In_923,In_872);
nor U180 (N_180,In_22,In_2340);
or U181 (N_181,In_2356,In_1077);
nor U182 (N_182,In_119,In_1212);
or U183 (N_183,In_445,In_2305);
nor U184 (N_184,In_2299,In_130);
xnor U185 (N_185,In_2181,In_611);
xnor U186 (N_186,In_1935,In_2314);
nand U187 (N_187,In_1597,In_2104);
nor U188 (N_188,In_14,In_2168);
xnor U189 (N_189,In_287,In_582);
xnor U190 (N_190,In_1796,In_1156);
nand U191 (N_191,In_2369,In_1748);
xnor U192 (N_192,In_1360,In_73);
and U193 (N_193,In_303,In_1817);
nand U194 (N_194,In_1573,In_1159);
xor U195 (N_195,In_2053,In_126);
or U196 (N_196,In_1621,In_1052);
and U197 (N_197,In_227,In_412);
nand U198 (N_198,In_449,In_1152);
xnor U199 (N_199,In_1896,In_1036);
nor U200 (N_200,In_2316,In_1071);
xor U201 (N_201,In_1316,In_207);
nand U202 (N_202,In_768,In_948);
and U203 (N_203,In_391,In_1745);
xnor U204 (N_204,In_1232,In_1415);
and U205 (N_205,In_2009,In_1886);
nand U206 (N_206,In_97,In_2143);
and U207 (N_207,In_1577,In_1699);
or U208 (N_208,In_294,In_1228);
and U209 (N_209,In_2021,In_2406);
xnor U210 (N_210,In_2197,In_1007);
nor U211 (N_211,In_1367,In_2140);
or U212 (N_212,In_1441,In_1277);
or U213 (N_213,In_1385,In_1428);
xnor U214 (N_214,In_1149,In_2085);
xor U215 (N_215,In_1416,In_933);
nand U216 (N_216,In_274,In_1917);
or U217 (N_217,In_451,In_699);
and U218 (N_218,In_1967,In_1078);
and U219 (N_219,In_244,In_692);
nand U220 (N_220,In_2222,In_2007);
xnor U221 (N_221,In_1275,In_1642);
nor U222 (N_222,In_444,In_1295);
xnor U223 (N_223,In_452,In_1663);
or U224 (N_224,In_1366,In_1311);
xnor U225 (N_225,In_2122,In_1913);
and U226 (N_226,In_1736,In_1404);
or U227 (N_227,In_672,In_884);
and U228 (N_228,In_837,In_1499);
xor U229 (N_229,In_1516,In_2405);
nor U230 (N_230,In_1457,In_1548);
nor U231 (N_231,In_1522,In_598);
or U232 (N_232,In_1587,In_3);
nor U233 (N_233,In_2040,In_900);
xor U234 (N_234,In_929,In_727);
nor U235 (N_235,In_1310,In_1022);
nand U236 (N_236,In_1481,In_860);
nand U237 (N_237,In_1501,In_1697);
or U238 (N_238,In_319,In_2138);
nor U239 (N_239,In_431,In_1502);
or U240 (N_240,In_508,In_818);
xor U241 (N_241,In_1954,In_678);
nor U242 (N_242,In_1009,In_1231);
and U243 (N_243,In_1624,In_98);
or U244 (N_244,In_1182,In_132);
and U245 (N_245,In_31,In_1473);
nor U246 (N_246,In_858,In_2169);
nor U247 (N_247,In_1118,In_171);
nor U248 (N_248,In_2350,In_1470);
xor U249 (N_249,In_376,In_1626);
nand U250 (N_250,In_1949,In_573);
or U251 (N_251,In_543,In_402);
nor U252 (N_252,In_1120,In_1846);
nand U253 (N_253,In_168,In_1547);
and U254 (N_254,In_2240,In_1062);
xor U255 (N_255,In_2469,In_2407);
and U256 (N_256,In_1162,In_1486);
nand U257 (N_257,In_2483,In_2446);
nor U258 (N_258,In_269,In_1780);
and U259 (N_259,In_2024,In_28);
and U260 (N_260,In_321,In_1902);
or U261 (N_261,In_1599,In_526);
nand U262 (N_262,In_2493,In_512);
and U263 (N_263,In_2257,In_1413);
or U264 (N_264,In_732,In_1487);
or U265 (N_265,In_569,In_1055);
nor U266 (N_266,In_2105,In_1422);
nand U267 (N_267,In_2165,In_1694);
or U268 (N_268,In_585,In_446);
nand U269 (N_269,In_908,In_898);
xnor U270 (N_270,In_1369,In_1904);
and U271 (N_271,In_2309,In_32);
nand U272 (N_272,In_1320,In_2345);
nor U273 (N_273,In_1881,In_640);
and U274 (N_274,In_2155,In_1133);
xnor U275 (N_275,In_1453,In_570);
xor U276 (N_276,In_1801,In_1451);
and U277 (N_277,In_71,In_63);
and U278 (N_278,In_907,In_2249);
nor U279 (N_279,In_674,In_1669);
nand U280 (N_280,In_242,In_440);
xor U281 (N_281,In_750,In_883);
and U282 (N_282,In_1167,In_473);
or U283 (N_283,In_561,In_1860);
nor U284 (N_284,In_614,In_2280);
xnor U285 (N_285,In_804,In_987);
or U286 (N_286,In_347,In_803);
nor U287 (N_287,In_226,In_1631);
xnor U288 (N_288,In_2126,In_554);
and U289 (N_289,In_99,In_1201);
xor U290 (N_290,In_1365,In_2057);
and U291 (N_291,In_655,In_1237);
nand U292 (N_292,In_1342,In_648);
or U293 (N_293,In_430,In_2343);
nor U294 (N_294,In_288,In_1665);
nand U295 (N_295,In_2243,In_1177);
nand U296 (N_296,In_1196,In_2230);
xnor U297 (N_297,In_539,In_271);
nor U298 (N_298,In_2419,In_1825);
nor U299 (N_299,In_2045,In_146);
or U300 (N_300,In_1853,In_1550);
and U301 (N_301,In_125,In_1183);
and U302 (N_302,In_825,In_660);
xnor U303 (N_303,In_234,In_1426);
and U304 (N_304,In_489,In_374);
xor U305 (N_305,In_255,In_1076);
nand U306 (N_306,In_179,In_1300);
xnor U307 (N_307,In_1371,In_1659);
and U308 (N_308,In_2355,In_1019);
nor U309 (N_309,In_1668,In_1172);
or U310 (N_310,In_658,In_1980);
xor U311 (N_311,In_1444,In_160);
xnor U312 (N_312,In_401,In_1572);
or U313 (N_313,In_2036,In_517);
nor U314 (N_314,In_328,In_329);
xnor U315 (N_315,In_2395,In_950);
xor U316 (N_316,In_1072,In_474);
nor U317 (N_317,In_607,In_511);
nand U318 (N_318,In_1443,In_695);
xor U319 (N_319,In_2420,In_1568);
and U320 (N_320,In_849,In_797);
xnor U321 (N_321,In_2098,In_1313);
xnor U322 (N_322,In_237,In_2393);
nor U323 (N_323,In_2107,In_1253);
nand U324 (N_324,In_1604,In_1438);
nand U325 (N_325,In_2184,In_566);
nor U326 (N_326,In_2491,In_1476);
and U327 (N_327,In_1037,In_1925);
nor U328 (N_328,In_2092,In_2101);
or U329 (N_329,In_1016,In_405);
or U330 (N_330,In_1618,In_2325);
and U331 (N_331,In_1589,In_1776);
or U332 (N_332,In_127,In_1869);
or U333 (N_333,In_1951,In_902);
or U334 (N_334,In_235,In_1376);
nor U335 (N_335,In_1091,In_1086);
xor U336 (N_336,In_1208,In_1727);
nor U337 (N_337,In_1029,In_264);
and U338 (N_338,In_1892,In_1322);
or U339 (N_339,In_339,In_2488);
and U340 (N_340,In_1056,In_1065);
nand U341 (N_341,In_1084,In_1085);
xor U342 (N_342,In_954,In_1254);
nor U343 (N_343,In_1176,In_1974);
xnor U344 (N_344,In_1559,In_810);
and U345 (N_345,In_2193,In_472);
xor U346 (N_346,In_1068,In_1989);
nand U347 (N_347,In_9,In_681);
nor U348 (N_348,In_1837,In_1990);
nand U349 (N_349,In_525,In_909);
nand U350 (N_350,In_1829,In_1586);
or U351 (N_351,In_1128,In_33);
nand U352 (N_352,In_358,In_2231);
and U353 (N_353,In_1020,In_2108);
xor U354 (N_354,In_789,In_1195);
and U355 (N_355,In_2304,In_1127);
nor U356 (N_356,In_2409,In_365);
nand U357 (N_357,In_1484,In_2121);
nand U358 (N_358,In_1619,In_1002);
or U359 (N_359,In_335,In_375);
xnor U360 (N_360,In_1259,In_299);
xor U361 (N_361,In_153,In_2112);
nand U362 (N_362,In_772,In_1440);
nand U363 (N_363,In_1800,In_576);
nand U364 (N_364,In_505,In_2035);
or U365 (N_365,In_1081,In_1864);
xor U366 (N_366,In_2091,In_1973);
and U367 (N_367,In_996,In_2421);
nand U368 (N_368,In_1703,In_1542);
and U369 (N_369,In_2402,In_916);
or U370 (N_370,In_1643,In_174);
and U371 (N_371,In_1349,In_194);
nand U372 (N_372,In_1724,In_2429);
xnor U373 (N_373,In_1806,In_532);
nor U374 (N_374,In_926,In_531);
nor U375 (N_375,In_1646,In_558);
or U376 (N_376,In_2044,In_875);
xor U377 (N_377,In_217,In_248);
nor U378 (N_378,In_2001,In_2000);
xnor U379 (N_379,In_1206,In_1716);
and U380 (N_380,In_305,In_1557);
and U381 (N_381,In_229,In_2451);
xnor U382 (N_382,In_1493,In_806);
and U383 (N_383,In_938,In_1912);
or U384 (N_384,In_1725,In_2210);
nor U385 (N_385,In_1644,In_231);
and U386 (N_386,In_813,In_466);
and U387 (N_387,In_2414,In_1681);
xnor U388 (N_388,In_1092,In_463);
or U389 (N_389,In_1911,In_190);
nor U390 (N_390,In_581,In_108);
nor U391 (N_391,In_840,In_578);
xnor U392 (N_392,In_2282,In_1992);
nand U393 (N_393,In_2283,In_448);
nor U394 (N_394,In_362,In_260);
and U395 (N_395,In_37,In_384);
xor U396 (N_396,In_2200,In_943);
nand U397 (N_397,In_1521,In_117);
nand U398 (N_398,In_1976,In_548);
or U399 (N_399,In_621,In_1962);
nor U400 (N_400,In_1622,In_1737);
or U401 (N_401,In_2374,In_1421);
or U402 (N_402,In_1221,In_10);
nor U403 (N_403,In_663,In_821);
or U404 (N_404,In_1392,In_414);
nor U405 (N_405,In_626,In_145);
nor U406 (N_406,In_2123,In_724);
and U407 (N_407,In_1777,In_2430);
and U408 (N_408,In_2068,In_36);
or U409 (N_409,In_2496,In_2326);
or U410 (N_410,In_1270,In_705);
and U411 (N_411,In_2300,In_2417);
xnor U412 (N_412,In_2312,In_546);
nor U413 (N_413,In_1373,In_1814);
xor U414 (N_414,In_2096,In_1382);
or U415 (N_415,In_1153,In_1676);
or U416 (N_416,In_182,In_1774);
and U417 (N_417,In_2400,In_23);
or U418 (N_418,In_2004,In_162);
xor U419 (N_419,In_1192,In_2359);
nor U420 (N_420,In_541,In_291);
nand U421 (N_421,In_265,In_538);
nand U422 (N_422,In_859,In_1197);
nor U423 (N_423,In_740,In_2338);
xor U424 (N_424,In_1592,In_2095);
xor U425 (N_425,In_639,In_1107);
and U426 (N_426,In_1760,In_461);
and U427 (N_427,In_1798,In_459);
or U428 (N_428,In_1882,In_2411);
or U429 (N_429,In_4,In_2087);
nand U430 (N_430,In_2333,In_1097);
and U431 (N_431,In_864,In_1137);
xnor U432 (N_432,In_141,In_2198);
nand U433 (N_433,In_60,In_1855);
nor U434 (N_434,In_2377,In_1362);
nor U435 (N_435,In_1719,In_2495);
nor U436 (N_436,In_513,In_953);
nand U437 (N_437,In_1707,In_2379);
nor U438 (N_438,In_1844,In_1200);
xor U439 (N_439,In_1564,In_767);
or U440 (N_440,In_2327,In_1132);
and U441 (N_441,In_1123,In_249);
xor U442 (N_442,In_1509,In_1909);
nand U443 (N_443,In_2255,In_795);
nor U444 (N_444,In_497,In_382);
xor U445 (N_445,In_544,In_564);
nor U446 (N_446,In_1517,In_1040);
nor U447 (N_447,In_1303,In_1608);
and U448 (N_448,In_201,In_1721);
and U449 (N_449,In_694,In_1276);
nor U450 (N_450,In_1792,In_165);
xnor U451 (N_451,In_1265,In_1804);
nor U452 (N_452,In_1247,In_1391);
nor U453 (N_453,In_338,In_1095);
nand U454 (N_454,In_111,In_296);
and U455 (N_455,In_372,In_877);
nor U456 (N_456,In_481,In_87);
nor U457 (N_457,In_197,In_199);
and U458 (N_458,In_152,In_1647);
and U459 (N_459,In_59,In_1885);
xnor U460 (N_460,In_2347,In_2093);
xnor U461 (N_461,In_2214,In_587);
nor U462 (N_462,In_1046,In_2237);
xnor U463 (N_463,In_2245,In_343);
and U464 (N_464,In_2382,In_1591);
or U465 (N_465,In_366,In_1430);
xor U466 (N_466,In_2415,In_1185);
xnor U467 (N_467,In_1188,In_711);
nor U468 (N_468,In_1160,In_1808);
or U469 (N_469,In_1728,In_2301);
nand U470 (N_470,In_2246,In_995);
nand U471 (N_471,In_1234,In_2216);
nand U472 (N_472,In_1928,In_1856);
nor U473 (N_473,In_1429,In_1435);
and U474 (N_474,In_494,In_1972);
and U475 (N_475,In_522,In_1306);
or U476 (N_476,In_1344,In_450);
and U477 (N_477,In_1474,In_439);
nor U478 (N_478,In_150,In_1741);
nand U479 (N_479,In_475,In_982);
nor U480 (N_480,In_1111,In_1532);
and U481 (N_481,In_1433,In_1929);
and U482 (N_482,In_1015,In_1174);
nand U483 (N_483,In_142,In_1375);
or U484 (N_484,In_1044,In_2310);
xnor U485 (N_485,In_1991,In_605);
xor U486 (N_486,In_528,In_1788);
and U487 (N_487,In_156,In_1899);
nor U488 (N_488,In_945,In_1080);
or U489 (N_489,In_94,In_51);
nor U490 (N_490,In_1216,In_427);
xor U491 (N_491,In_828,In_419);
and U492 (N_492,In_1791,In_379);
or U493 (N_493,In_2319,In_1328);
xor U494 (N_494,In_1987,In_1238);
nor U495 (N_495,In_509,In_1556);
xor U496 (N_496,In_1513,In_91);
and U497 (N_497,In_1988,In_1299);
xnor U498 (N_498,In_1288,In_2206);
and U499 (N_499,In_399,In_742);
nor U500 (N_500,In_1761,In_1883);
nor U501 (N_501,In_2290,In_355);
nand U502 (N_502,In_600,In_747);
nand U503 (N_503,In_1857,In_189);
nand U504 (N_504,In_2362,In_1875);
xnor U505 (N_505,In_113,In_1833);
and U506 (N_506,In_897,In_1771);
or U507 (N_507,In_1872,In_787);
nor U508 (N_508,In_224,In_2367);
nor U509 (N_509,In_2058,In_2132);
or U510 (N_510,In_1500,In_1570);
or U511 (N_511,In_2031,In_307);
or U512 (N_512,In_2477,In_1965);
and U513 (N_513,In_649,In_76);
nand U514 (N_514,In_426,In_1750);
xnor U515 (N_515,In_949,In_2281);
xnor U516 (N_516,In_2348,In_911);
nor U517 (N_517,In_1514,In_2373);
nor U518 (N_518,In_2144,In_1740);
nand U519 (N_519,In_904,In_30);
and U520 (N_520,In_373,In_2005);
or U521 (N_521,In_809,In_1454);
and U522 (N_522,In_934,In_1865);
or U523 (N_523,In_2323,In_1613);
nor U524 (N_524,In_1460,In_245);
and U525 (N_525,In_2357,In_2011);
or U526 (N_526,In_369,In_1402);
and U527 (N_527,In_1031,In_1718);
nand U528 (N_528,In_1887,In_122);
nand U529 (N_529,In_1468,In_388);
xor U530 (N_530,In_1610,In_2462);
xor U531 (N_531,In_889,In_40);
and U532 (N_532,In_2391,In_2055);
and U533 (N_533,In_1066,In_2090);
or U534 (N_534,In_972,In_2196);
nor U535 (N_535,In_1790,In_315);
nor U536 (N_536,In_1753,In_2445);
and U537 (N_537,In_290,In_1087);
or U538 (N_538,In_403,In_1498);
xnor U539 (N_539,In_181,In_880);
nand U540 (N_540,In_6,In_2071);
nand U541 (N_541,In_1038,In_601);
xnor U542 (N_542,In_2434,In_1945);
nand U543 (N_543,In_1446,In_1948);
nor U544 (N_544,In_232,In_688);
xnor U545 (N_545,In_2302,In_1103);
or U546 (N_546,In_443,In_1380);
or U547 (N_547,In_1585,In_1011);
and U548 (N_548,In_841,In_1851);
xnor U549 (N_549,In_560,In_2099);
xnor U550 (N_550,In_1332,In_1561);
or U551 (N_551,In_1387,In_348);
nand U552 (N_552,In_1870,In_2185);
nor U553 (N_553,In_918,In_134);
xnor U554 (N_554,In_927,In_2042);
or U555 (N_555,In_92,In_2145);
nand U556 (N_556,In_1045,In_799);
or U557 (N_557,In_653,In_976);
nand U558 (N_558,In_236,In_2052);
nor U559 (N_559,In_613,In_2135);
nor U560 (N_560,In_673,In_721);
nor U561 (N_561,In_811,In_1089);
or U562 (N_562,In_20,In_1742);
nand U563 (N_563,In_959,In_1480);
or U564 (N_564,In_2443,In_832);
nor U565 (N_565,In_2069,In_2474);
nor U566 (N_566,In_1189,In_1243);
xnor U567 (N_567,In_381,In_1271);
xnor U568 (N_568,In_941,In_851);
xor U569 (N_569,In_1117,In_370);
or U570 (N_570,In_634,In_2067);
or U571 (N_571,In_490,In_434);
nand U572 (N_572,In_1769,In_2346);
and U573 (N_573,In_2043,In_302);
nand U574 (N_574,In_2298,In_344);
xor U575 (N_575,In_739,In_2472);
nor U576 (N_576,In_1920,In_2267);
and U577 (N_577,In_1601,In_1255);
or U578 (N_578,In_460,In_1351);
nand U579 (N_579,In_1114,In_606);
nor U580 (N_580,In_1632,In_383);
nand U581 (N_581,In_932,In_572);
nor U582 (N_582,In_1048,In_1698);
and U583 (N_583,In_1401,In_1298);
xnor U584 (N_584,In_1903,In_424);
nor U585 (N_585,In_885,In_764);
or U586 (N_586,In_1357,In_792);
nor U587 (N_587,In_1267,In_1057);
xnor U588 (N_588,In_1358,In_1558);
nor U589 (N_589,In_2455,In_1927);
or U590 (N_590,In_1739,In_1831);
or U591 (N_591,In_1035,In_1503);
or U592 (N_592,In_823,In_2361);
and U593 (N_593,In_2228,In_856);
xnor U594 (N_594,In_2065,In_2106);
or U595 (N_595,In_75,In_718);
nor U596 (N_596,In_2127,In_878);
xor U597 (N_597,In_2269,In_1705);
nand U598 (N_598,In_1361,In_1757);
or U599 (N_599,In_1571,In_1448);
nor U600 (N_600,In_368,In_985);
nor U601 (N_601,In_2397,In_2015);
nand U602 (N_602,In_971,In_791);
or U603 (N_603,In_2061,In_1775);
or U604 (N_604,In_602,In_1813);
nor U605 (N_605,In_624,In_1098);
nand U606 (N_606,In_1252,In_1069);
xnor U607 (N_607,In_273,In_906);
nand U608 (N_608,In_2479,In_1759);
xor U609 (N_609,In_46,In_436);
and U610 (N_610,In_2375,In_2440);
xor U611 (N_611,In_100,In_378);
or U612 (N_612,In_195,In_510);
or U613 (N_613,In_967,In_1406);
and U614 (N_614,In_829,In_1063);
nand U615 (N_615,In_423,In_1214);
xor U616 (N_616,In_1292,In_2439);
nor U617 (N_617,In_364,In_816);
nor U618 (N_618,In_1388,In_1985);
and U619 (N_619,In_1734,In_1524);
and U620 (N_620,In_2060,In_387);
nand U621 (N_621,In_1386,In_409);
or U622 (N_622,In_1679,In_1193);
or U623 (N_623,In_1249,In_2014);
or U624 (N_624,In_2436,In_680);
nand U625 (N_625,In_1125,In_1674);
or U626 (N_626,In_2103,In_1684);
or U627 (N_627,In_455,In_599);
or U628 (N_628,In_1545,In_1505);
xnor U629 (N_629,In_1653,In_719);
nor U630 (N_630,In_1496,In_2251);
and U631 (N_631,In_124,In_482);
nor U632 (N_632,In_2195,In_1704);
xor U633 (N_633,In_1764,In_1067);
nand U634 (N_634,In_1266,In_930);
xor U635 (N_635,In_1350,In_1984);
nor U636 (N_636,In_1732,In_2404);
xor U637 (N_637,In_784,In_392);
or U638 (N_638,In_1262,In_1331);
nand U639 (N_639,In_857,In_1058);
and U640 (N_640,In_295,In_515);
or U641 (N_641,In_565,In_1109);
and U642 (N_642,In_1510,In_1315);
and U643 (N_643,In_899,In_2008);
or U644 (N_644,In_230,In_1768);
nor U645 (N_645,In_2431,In_214);
or U646 (N_646,In_1931,In_453);
or U647 (N_647,In_1937,In_121);
and U648 (N_648,In_1148,In_1340);
nor U649 (N_649,In_2279,In_1787);
or U650 (N_650,In_2154,In_1364);
and U651 (N_651,In_351,In_1467);
nor U652 (N_652,In_1284,In_1347);
or U653 (N_653,In_1906,In_1600);
xnor U654 (N_654,In_1582,In_622);
or U655 (N_655,In_432,In_1260);
nand U656 (N_656,In_1343,In_1013);
nand U657 (N_657,In_2452,In_2063);
and U658 (N_658,In_272,In_1239);
nor U659 (N_659,In_1054,In_1617);
nand U660 (N_660,In_2118,In_1115);
nor U661 (N_661,In_1922,In_175);
nand U662 (N_662,In_270,In_223);
nand U663 (N_663,In_2023,In_2435);
nor U664 (N_664,In_845,In_407);
nor U665 (N_665,In_545,In_667);
nand U666 (N_666,In_751,In_2056);
or U667 (N_667,In_1507,In_1534);
and U668 (N_668,In_1849,In_683);
xor U669 (N_669,In_311,In_1293);
or U670 (N_670,In_390,In_123);
nor U671 (N_671,In_527,In_1006);
xor U672 (N_672,In_1970,In_1169);
xnor U673 (N_673,In_433,In_1224);
nor U674 (N_674,In_386,In_334);
nor U675 (N_675,In_775,In_1489);
or U676 (N_676,In_955,In_357);
nor U677 (N_677,In_2238,In_1921);
xnor U678 (N_678,In_1477,In_2466);
or U679 (N_679,In_2442,In_429);
xnor U680 (N_680,In_1978,In_1938);
and U681 (N_681,In_1497,In_1168);
xnor U682 (N_682,In_905,In_2219);
nand U683 (N_683,In_340,In_1575);
nand U684 (N_684,In_148,In_2470);
and U685 (N_685,In_228,In_973);
or U686 (N_686,In_193,In_47);
nor U687 (N_687,In_523,In_1794);
nand U688 (N_688,In_212,In_783);
nor U689 (N_689,In_2342,In_630);
and U690 (N_690,In_2114,In_1543);
xor U691 (N_691,In_1636,In_1838);
nand U692 (N_692,In_354,In_1204);
xor U693 (N_693,In_970,In_822);
nand U694 (N_694,In_625,In_2038);
or U695 (N_695,In_1656,In_1605);
xnor U696 (N_696,In_58,In_2387);
nor U697 (N_697,In_882,In_617);
nor U698 (N_698,In_1947,In_812);
nor U699 (N_699,In_676,In_2482);
and U700 (N_700,In_1290,In_2297);
nand U701 (N_701,In_891,In_1027);
and U702 (N_702,In_442,In_2344);
and U703 (N_703,In_2295,In_1466);
or U704 (N_704,In_652,In_1395);
xor U705 (N_705,In_1670,In_1820);
nand U706 (N_706,In_2364,In_1816);
nor U707 (N_707,In_1614,In_656);
nand U708 (N_708,In_1423,In_240);
nand U709 (N_709,In_2385,In_1230);
or U710 (N_710,In_2471,In_428);
xnor U711 (N_711,In_1032,In_1094);
xor U712 (N_712,In_13,In_1126);
nor U713 (N_713,In_502,In_389);
or U714 (N_714,In_815,In_164);
xor U715 (N_715,In_1108,In_77);
and U716 (N_716,In_1730,In_253);
xor U717 (N_717,In_1850,In_2456);
or U718 (N_718,In_282,In_894);
nand U719 (N_719,In_2187,In_210);
or U720 (N_720,In_1696,In_616);
or U721 (N_721,In_805,In_831);
or U722 (N_722,In_922,In_1348);
xnor U723 (N_723,In_353,In_888);
or U724 (N_724,In_2292,In_276);
and U725 (N_725,In_2476,In_2152);
xor U726 (N_726,In_2183,In_1100);
nor U727 (N_727,In_1995,In_93);
and U728 (N_728,In_855,In_131);
xor U729 (N_729,In_2148,In_1683);
and U730 (N_730,In_1835,In_309);
xor U731 (N_731,In_2339,In_1841);
and U732 (N_732,In_250,In_1602);
and U733 (N_733,In_2275,In_67);
or U734 (N_734,In_1834,In_817);
or U735 (N_735,In_868,In_1763);
or U736 (N_736,In_491,In_519);
nand U737 (N_737,In_499,In_278);
xor U738 (N_738,In_1297,In_781);
and U739 (N_739,In_713,In_1124);
nand U740 (N_740,In_1823,In_1143);
nand U741 (N_741,In_796,In_836);
nor U742 (N_742,In_1799,In_735);
nand U743 (N_743,In_650,In_1393);
xor U744 (N_744,In_1723,In_283);
and U745 (N_745,In_1781,In_2368);
xnor U746 (N_746,In_2336,In_1641);
nand U747 (N_747,In_1165,In_159);
nand U748 (N_748,In_1263,In_1596);
and U749 (N_749,In_1979,In_1612);
or U750 (N_750,In_761,In_1110);
xnor U751 (N_751,In_2448,In_2006);
and U752 (N_752,In_755,In_2084);
xor U753 (N_753,In_847,In_1112);
or U754 (N_754,In_597,In_2158);
nor U755 (N_755,In_1005,In_1566);
xnor U756 (N_756,In_2389,In_846);
and U757 (N_757,In_1179,In_1934);
xor U758 (N_758,In_361,In_1093);
or U759 (N_759,In_56,In_1282);
or U760 (N_760,In_848,In_259);
or U761 (N_761,In_1797,In_774);
nand U762 (N_762,In_1960,In_838);
xnor U763 (N_763,In_1525,In_1907);
or U764 (N_764,In_1409,In_842);
xnor U765 (N_765,In_2136,In_1981);
or U766 (N_766,In_377,In_1722);
xnor U767 (N_767,In_1268,In_2039);
or U768 (N_768,In_2225,In_715);
nand U769 (N_769,In_80,In_135);
nor U770 (N_770,In_95,In_479);
nand U771 (N_771,In_1251,In_1749);
xor U772 (N_772,In_1533,In_2438);
nor U773 (N_773,In_2188,In_246);
xor U774 (N_774,In_794,In_1744);
xor U775 (N_775,In_568,In_400);
and U776 (N_776,In_1437,In_138);
nor U777 (N_777,In_714,In_644);
or U778 (N_778,In_1609,In_21);
xor U779 (N_779,In_866,In_708);
and U780 (N_780,In_1475,In_1494);
and U781 (N_781,In_1866,In_586);
nand U782 (N_782,In_2226,In_700);
nor U783 (N_783,In_2272,In_779);
nand U784 (N_784,In_2321,In_2050);
xor U785 (N_785,In_612,In_754);
and U786 (N_786,In_984,In_2481);
and U787 (N_787,In_2190,In_1023);
nand U788 (N_788,In_2156,In_951);
nor U789 (N_789,In_2422,In_879);
or U790 (N_790,In_90,In_1419);
xnor U791 (N_791,In_1847,In_2318);
xnor U792 (N_792,In_1770,In_668);
nor U793 (N_793,In_238,In_1175);
xor U794 (N_794,In_2485,In_2072);
nor U795 (N_795,In_2161,In_2497);
nand U796 (N_796,In_2285,In_2117);
xor U797 (N_797,In_636,In_939);
nor U798 (N_798,In_209,In_1327);
and U799 (N_799,In_420,In_1257);
xnor U800 (N_800,In_516,In_331);
and U801 (N_801,In_1264,In_1088);
nand U802 (N_802,In_722,In_629);
or U803 (N_803,In_1479,In_2332);
xor U804 (N_804,In_966,In_34);
nor U805 (N_805,In_1836,In_915);
or U806 (N_806,In_2041,In_981);
nor U807 (N_807,In_486,In_1975);
nor U808 (N_808,In_1187,In_1772);
nor U809 (N_809,In_1803,In_136);
nand U810 (N_810,In_2075,In_802);
nand U811 (N_811,In_697,In_1940);
nor U812 (N_812,In_974,In_1702);
nand U813 (N_813,In_2062,In_2351);
and U814 (N_814,In_406,In_350);
nor U815 (N_815,In_1166,In_1639);
and U816 (N_816,In_2,In_745);
and U817 (N_817,In_1051,In_2227);
and U818 (N_818,In_1890,In_2371);
or U819 (N_819,In_593,In_808);
nor U820 (N_820,In_262,In_1607);
xor U821 (N_821,In_1616,In_643);
or U822 (N_822,In_1272,In_202);
or U823 (N_823,In_48,In_1170);
and U824 (N_824,In_314,In_2054);
and U825 (N_825,In_1955,In_1933);
nor U826 (N_826,In_172,In_780);
xnor U827 (N_827,In_2151,In_577);
xnor U828 (N_828,In_1033,In_2175);
xor U829 (N_829,In_17,In_595);
or U830 (N_830,In_15,In_457);
nor U831 (N_831,In_1047,In_1651);
and U832 (N_832,In_1648,In_317);
xnor U833 (N_833,In_327,In_1025);
or U834 (N_834,In_999,In_1447);
nor U835 (N_835,In_39,In_2027);
and U836 (N_836,In_2322,In_1717);
xor U837 (N_837,In_2412,In_896);
nand U838 (N_838,In_575,In_1139);
and U839 (N_839,In_1969,In_1560);
or U840 (N_840,In_876,In_2384);
nand U841 (N_841,In_1325,In_1511);
and U842 (N_842,In_865,In_441);
nor U843 (N_843,In_1464,In_1142);
or U844 (N_844,In_279,In_559);
nor U845 (N_845,In_2437,In_16);
or U846 (N_846,In_873,In_693);
nand U847 (N_847,In_782,In_1205);
nand U848 (N_848,In_977,In_1334);
and U849 (N_849,In_1286,In_1598);
nor U850 (N_850,In_2247,In_1352);
and U851 (N_851,In_867,In_2164);
xor U852 (N_852,In_2208,In_1898);
nand U853 (N_853,In_1779,In_940);
or U854 (N_854,In_2233,In_196);
and U855 (N_855,In_2489,In_1105);
nor U856 (N_856,In_318,In_1871);
and U857 (N_857,In_363,In_2221);
nand U858 (N_858,In_881,In_590);
nor U859 (N_859,In_1304,In_2363);
or U860 (N_860,In_1314,In_1782);
or U861 (N_861,In_642,In_2086);
xor U862 (N_862,In_704,In_997);
nand U863 (N_863,In_1171,In_556);
xnor U864 (N_864,In_843,In_1424);
nand U865 (N_865,In_233,In_180);
or U866 (N_866,In_833,In_2460);
or U867 (N_867,In_1488,In_1762);
nor U868 (N_868,In_2047,In_140);
xnor U869 (N_869,In_2204,In_435);
nand U870 (N_870,In_1953,In_1964);
nor U871 (N_871,In_417,In_2303);
and U872 (N_872,In_820,In_2386);
and U873 (N_873,In_1673,In_1420);
nand U874 (N_874,In_447,In_2137);
or U875 (N_875,In_1151,In_2157);
xor U876 (N_876,In_2287,In_2341);
xnor U877 (N_877,In_498,In_2294);
nand U878 (N_878,In_2025,In_1184);
and U879 (N_879,In_1640,In_1400);
nor U880 (N_880,In_86,In_2002);
and U881 (N_881,In_1458,In_1789);
xor U882 (N_882,In_1843,In_1324);
and U883 (N_883,In_313,In_85);
and U884 (N_884,In_1551,In_646);
nand U885 (N_885,In_962,In_990);
or U886 (N_886,In_1807,In_1378);
nand U887 (N_887,In_322,In_41);
nand U888 (N_888,In_1720,In_550);
nand U889 (N_889,In_483,In_2147);
or U890 (N_890,In_684,In_2100);
and U891 (N_891,In_535,In_2113);
nand U892 (N_892,In_1956,In_2487);
nor U893 (N_893,In_38,In_819);
nand U894 (N_894,In_1060,In_1959);
xnor U895 (N_895,In_1246,In_1203);
and U896 (N_896,In_946,In_102);
and U897 (N_897,In_1283,In_110);
or U898 (N_898,In_1691,In_2083);
and U899 (N_899,In_669,In_425);
nor U900 (N_900,In_1010,In_1977);
or U901 (N_901,In_107,In_1667);
xor U902 (N_902,In_1999,In_198);
or U903 (N_903,In_221,In_1218);
xor U904 (N_904,In_1219,In_1138);
or U905 (N_905,In_592,In_1064);
and U906 (N_906,In_1932,In_2454);
xnor U907 (N_907,In_520,In_1519);
nand U908 (N_908,In_1758,In_1028);
xnor U909 (N_909,In_1997,In_2315);
nand U910 (N_910,In_958,In_2173);
nand U911 (N_911,In_861,In_81);
nand U912 (N_912,In_45,In_2174);
or U913 (N_913,In_729,In_1014);
nor U914 (N_914,In_826,In_631);
xnor U915 (N_915,In_1731,In_66);
xnor U916 (N_916,In_533,In_1963);
xnor U917 (N_917,In_1874,In_2259);
nor U918 (N_918,In_1,In_1733);
nand U919 (N_919,In_1030,In_2179);
nor U920 (N_920,In_1805,In_105);
nand U921 (N_921,In_184,In_2232);
xnor U922 (N_922,In_2244,In_2383);
and U923 (N_923,In_204,In_2022);
xnor U924 (N_924,In_993,In_524);
nor U925 (N_925,In_1830,In_547);
xnor U926 (N_926,In_393,In_218);
nand U927 (N_927,In_2018,In_470);
nand U928 (N_928,In_886,In_68);
xnor U929 (N_929,In_1942,In_2217);
xor U930 (N_930,In_2120,In_752);
and U931 (N_931,In_2020,In_920);
and U932 (N_932,In_112,In_776);
and U933 (N_933,In_2358,In_1919);
xnor U934 (N_934,In_1765,In_2324);
and U935 (N_935,In_1530,In_1821);
xor U936 (N_936,In_1729,In_2124);
nand U937 (N_937,In_2307,In_2046);
xnor U938 (N_938,In_1747,In_1785);
and U939 (N_939,In_551,In_2293);
xnor U940 (N_940,In_1828,In_1113);
and U941 (N_941,In_2372,In_557);
nand U942 (N_942,In_2453,In_1287);
xnor U943 (N_943,In_1135,In_690);
nand U944 (N_944,In_5,In_1946);
nand U945 (N_945,In_1655,In_1515);
or U946 (N_946,In_1795,In_2378);
nand U947 (N_947,In_980,In_1897);
nand U948 (N_948,In_177,In_293);
nor U949 (N_949,In_1824,In_903);
nand U950 (N_950,In_55,In_2088);
or U951 (N_951,In_2199,In_1583);
or U952 (N_952,In_871,In_2433);
nand U953 (N_953,In_1810,In_975);
or U954 (N_954,In_1880,In_1017);
nor U955 (N_955,In_1021,In_1274);
or U956 (N_956,In_1778,In_1305);
nand U957 (N_957,In_2499,In_50);
or U958 (N_958,In_78,In_415);
nor U959 (N_959,In_2186,In_2026);
or U960 (N_960,In_2313,In_61);
and U961 (N_961,In_500,In_2170);
nand U962 (N_962,In_589,In_166);
nand U963 (N_963,In_844,In_1625);
nor U964 (N_964,In_2130,In_155);
or U965 (N_965,In_385,In_2077);
nand U966 (N_966,In_114,In_1506);
and U967 (N_967,In_1280,In_2037);
nor U968 (N_968,In_1083,In_1178);
nor U969 (N_969,In_1527,In_163);
nand U970 (N_970,In_1994,In_1961);
and U971 (N_971,In_763,In_281);
nand U972 (N_972,In_2215,In_52);
nor U973 (N_973,In_2146,In_1308);
and U974 (N_974,In_1936,In_2376);
or U975 (N_975,In_2013,In_252);
or U976 (N_976,In_1059,In_1329);
xor U977 (N_977,In_1323,In_1450);
nor U978 (N_978,In_887,In_2353);
nand U979 (N_979,In_284,In_800);
or U980 (N_980,In_1198,In_901);
xor U981 (N_981,In_192,In_1241);
and U982 (N_982,In_912,In_2494);
or U983 (N_983,In_1958,In_161);
and U984 (N_984,In_1405,In_1355);
or U985 (N_985,In_1859,In_2192);
nand U986 (N_986,In_1226,In_726);
or U987 (N_987,In_2258,In_239);
nand U988 (N_988,In_2252,In_1715);
nand U989 (N_989,In_2413,In_1726);
nor U990 (N_990,In_154,In_1891);
and U991 (N_991,In_1034,In_404);
nor U992 (N_992,In_1321,In_222);
xnor U993 (N_993,In_1227,In_1535);
and U994 (N_994,In_496,In_2166);
and U995 (N_995,In_991,In_2260);
and U996 (N_996,In_2424,In_2133);
xnor U997 (N_997,In_26,In_1968);
and U998 (N_998,In_380,In_2241);
nand U999 (N_999,In_2182,In_1463);
or U1000 (N_1000,In_1104,In_917);
nor U1001 (N_1001,In_286,In_2296);
nand U1002 (N_1002,In_1471,In_2458);
xor U1003 (N_1003,In_2094,In_2408);
nor U1004 (N_1004,In_1242,In_1377);
nand U1005 (N_1005,In_495,In_2160);
xor U1006 (N_1006,In_316,In_1173);
nor U1007 (N_1007,In_1082,In_2418);
and U1008 (N_1008,In_852,In_1445);
xor U1009 (N_1009,In_2306,In_1854);
or U1010 (N_1010,In_608,In_2207);
nand U1011 (N_1011,In_2218,In_173);
and U1012 (N_1012,In_762,In_1294);
nand U1013 (N_1013,In_1330,In_476);
nor U1014 (N_1014,In_11,In_1042);
nor U1015 (N_1015,In_1157,In_83);
and U1016 (N_1016,In_247,In_2468);
xnor U1017 (N_1017,In_1590,In_225);
xnor U1018 (N_1018,In_8,In_118);
or U1019 (N_1019,In_563,In_2162);
or U1020 (N_1020,In_1281,In_1408);
or U1021 (N_1021,In_352,In_1465);
nand U1022 (N_1022,In_1784,In_1312);
or U1023 (N_1023,In_2486,In_1738);
or U1024 (N_1024,In_2163,In_1410);
nand U1025 (N_1025,In_701,In_1706);
and U1026 (N_1026,In_757,In_1379);
nand U1027 (N_1027,In_835,In_1893);
nand U1028 (N_1028,In_1544,In_1822);
xnor U1029 (N_1029,In_2492,In_422);
nand U1030 (N_1030,In_986,In_133);
or U1031 (N_1031,In_1595,In_2134);
nand U1032 (N_1032,In_1049,In_514);
nand U1033 (N_1033,In_610,In_691);
xnor U1034 (N_1034,In_137,In_1101);
or U1035 (N_1035,In_1026,In_744);
nor U1036 (N_1036,In_1862,In_1826);
nor U1037 (N_1037,In_824,In_753);
nand U1038 (N_1038,In_834,In_2019);
or U1039 (N_1039,In_1278,In_2352);
or U1040 (N_1040,In_88,In_571);
xor U1041 (N_1041,In_1161,In_1129);
nand U1042 (N_1042,In_679,In_2049);
nor U1043 (N_1043,In_2102,In_2416);
xor U1044 (N_1044,In_298,In_1217);
nor U1045 (N_1045,In_1353,In_1210);
and U1046 (N_1046,In_398,In_696);
or U1047 (N_1047,In_1412,In_1455);
nor U1048 (N_1048,In_870,In_2109);
or U1049 (N_1049,In_1418,In_2467);
and U1050 (N_1050,In_654,In_1852);
or U1051 (N_1051,In_1462,In_1134);
and U1052 (N_1052,In_2270,In_759);
or U1053 (N_1053,In_2284,In_2277);
nor U1054 (N_1054,In_1075,In_1074);
or U1055 (N_1055,In_1710,In_604);
and U1056 (N_1056,In_503,In_2432);
and U1057 (N_1057,In_2271,In_349);
nor U1058 (N_1058,In_2153,In_1302);
or U1059 (N_1059,In_1537,In_2425);
nand U1060 (N_1060,In_555,In_2380);
or U1061 (N_1061,In_267,In_2331);
nor U1062 (N_1062,In_1390,In_1914);
or U1063 (N_1063,In_1584,In_1154);
nand U1064 (N_1064,In_256,In_1202);
or U1065 (N_1065,In_778,In_2263);
xor U1066 (N_1066,In_632,In_839);
and U1067 (N_1067,In_2265,In_2224);
nor U1068 (N_1068,In_2426,In_675);
and U1069 (N_1069,In_1399,In_2349);
nor U1070 (N_1070,In_310,In_702);
nor U1071 (N_1071,In_1491,In_1472);
nor U1072 (N_1072,In_1645,In_942);
or U1073 (N_1073,In_540,In_336);
nor U1074 (N_1074,In_116,In_756);
and U1075 (N_1075,In_2354,In_2399);
nor U1076 (N_1076,In_1538,In_2176);
nor U1077 (N_1077,In_72,In_2076);
nand U1078 (N_1078,In_1756,In_2390);
nand U1079 (N_1079,In_1180,In_2017);
nand U1080 (N_1080,In_2074,In_465);
or U1081 (N_1081,In_418,In_2205);
or U1082 (N_1082,In_1713,In_128);
or U1083 (N_1083,In_1941,In_709);
nand U1084 (N_1084,In_1482,In_1637);
nand U1085 (N_1085,In_574,In_1666);
nor U1086 (N_1086,In_1918,In_707);
nor U1087 (N_1087,In_2209,In_1579);
or U1088 (N_1088,In_1709,In_1536);
or U1089 (N_1089,In_1746,In_2274);
or U1090 (N_1090,In_1766,In_1396);
nand U1091 (N_1091,In_1394,In_777);
and U1092 (N_1092,In_1490,In_1867);
and U1093 (N_1093,In_27,In_1752);
and U1094 (N_1094,In_567,In_1815);
or U1095 (N_1095,In_1876,In_1555);
nor U1096 (N_1096,In_1628,In_1671);
xnor U1097 (N_1097,In_1147,In_471);
and U1098 (N_1098,In_216,In_1658);
xnor U1099 (N_1099,In_623,In_2398);
nor U1100 (N_1100,In_1531,In_960);
nor U1101 (N_1101,In_480,In_115);
and U1102 (N_1102,In_367,In_304);
or U1103 (N_1103,In_24,In_220);
xor U1104 (N_1104,In_2381,In_628);
nor U1105 (N_1105,In_1432,In_1578);
xor U1106 (N_1106,In_1427,In_1863);
nand U1107 (N_1107,In_1574,In_147);
or U1108 (N_1108,In_1567,In_254);
nor U1109 (N_1109,In_1877,In_944);
and U1110 (N_1110,In_983,In_1526);
xor U1111 (N_1111,In_925,In_1520);
or U1112 (N_1112,In_1397,In_1743);
or U1113 (N_1113,In_1053,In_35);
nor U1114 (N_1114,In_850,In_725);
nor U1115 (N_1115,In_1576,In_1915);
or U1116 (N_1116,In_2261,In_765);
and U1117 (N_1117,In_786,In_2211);
nand U1118 (N_1118,In_484,In_1685);
and U1119 (N_1119,In_79,In_853);
nor U1120 (N_1120,In_2097,In_596);
nor U1121 (N_1121,In_96,In_2119);
and U1122 (N_1122,In_186,In_1735);
nor U1123 (N_1123,In_2360,In_2012);
nor U1124 (N_1124,In_258,In_2248);
and U1125 (N_1125,In_2403,In_2149);
nand U1126 (N_1126,In_1346,In_1225);
nand U1127 (N_1127,In_2370,In_738);
nand U1128 (N_1128,In_1924,In_1827);
nand U1129 (N_1129,In_346,In_1712);
or U1130 (N_1130,In_2266,In_736);
xnor U1131 (N_1131,In_301,In_1456);
nand U1132 (N_1132,In_306,In_1562);
nand U1133 (N_1133,In_241,In_534);
xnor U1134 (N_1134,In_801,In_1194);
nand U1135 (N_1135,In_1793,In_243);
and U1136 (N_1136,In_1301,In_1289);
and U1137 (N_1137,In_671,In_1483);
xnor U1138 (N_1138,In_766,In_2388);
and U1139 (N_1139,In_1339,In_1627);
or U1140 (N_1140,In_549,In_1546);
xor U1141 (N_1141,In_139,In_89);
and U1142 (N_1142,In_65,In_706);
nor U1143 (N_1143,In_1381,In_2480);
or U1144 (N_1144,In_1211,In_717);
nor U1145 (N_1145,In_396,In_2473);
xnor U1146 (N_1146,In_1664,In_261);
xor U1147 (N_1147,In_2463,In_666);
or U1148 (N_1148,In_211,In_324);
nor U1149 (N_1149,In_1818,In_456);
nand U1150 (N_1150,In_1657,In_2201);
or U1151 (N_1151,In_1122,In_609);
or U1152 (N_1152,In_1634,In_1140);
nand U1153 (N_1153,In_807,In_645);
nand U1154 (N_1154,In_185,In_1425);
and U1155 (N_1155,In_2034,In_979);
nand U1156 (N_1156,In_1363,In_1181);
and U1157 (N_1157,In_869,In_1096);
nand U1158 (N_1158,In_1686,In_620);
xor U1159 (N_1159,In_1861,In_1190);
and U1160 (N_1160,In_19,In_965);
xnor U1161 (N_1161,In_769,In_359);
xor U1162 (N_1162,In_2392,In_2171);
nand U1163 (N_1163,In_521,In_1273);
and U1164 (N_1164,In_200,In_748);
nor U1165 (N_1165,In_2033,In_1905);
nor U1166 (N_1166,In_289,In_1244);
and U1167 (N_1167,In_2459,In_1431);
xor U1168 (N_1168,In_69,In_1832);
or U1169 (N_1169,In_300,In_1222);
or U1170 (N_1170,In_698,In_437);
xnor U1171 (N_1171,In_1370,In_2444);
nor U1172 (N_1172,In_2264,In_454);
nor U1173 (N_1173,In_1986,In_103);
and U1174 (N_1174,In_2139,In_2089);
xor U1175 (N_1175,In_956,In_1130);
nand U1176 (N_1176,In_591,In_2328);
xnor U1177 (N_1177,In_1693,In_1407);
xor U1178 (N_1178,In_1141,In_1269);
nand U1179 (N_1179,In_2465,In_1588);
xnor U1180 (N_1180,In_921,In_1163);
xnor U1181 (N_1181,In_1389,In_187);
nor U1182 (N_1182,In_57,In_2128);
nand U1183 (N_1183,In_208,In_158);
or U1184 (N_1184,In_1680,In_1326);
xnor U1185 (N_1185,In_1131,In_659);
or U1186 (N_1186,In_2141,In_537);
nor U1187 (N_1187,In_1452,In_785);
and U1188 (N_1188,In_1041,In_144);
xnor U1189 (N_1189,In_928,In_1687);
nor U1190 (N_1190,In_1754,In_2278);
nand U1191 (N_1191,In_205,In_1802);
and U1192 (N_1192,In_1638,In_280);
xnor U1193 (N_1193,In_178,In_830);
nor U1194 (N_1194,In_188,In_1993);
nor U1195 (N_1195,In_507,In_2288);
nor U1196 (N_1196,In_1518,In_1209);
nand U1197 (N_1197,In_2081,In_149);
nor U1198 (N_1198,In_2478,In_2464);
nand U1199 (N_1199,In_1345,In_467);
or U1200 (N_1200,In_1436,In_661);
or U1201 (N_1201,In_1998,In_1569);
nor U1202 (N_1202,In_2142,In_1442);
and U1203 (N_1203,In_760,In_312);
nor U1204 (N_1204,In_2159,In_662);
xnor U1205 (N_1205,In_1146,In_2253);
or U1206 (N_1206,In_477,In_2273);
or U1207 (N_1207,In_2396,In_1336);
xor U1208 (N_1208,In_493,In_1845);
or U1209 (N_1209,In_758,In_1971);
or U1210 (N_1210,In_1944,In_1061);
xor U1211 (N_1211,In_263,In_82);
nor U1212 (N_1212,In_266,In_120);
and U1213 (N_1213,In_413,In_1615);
xnor U1214 (N_1214,In_1145,In_257);
nor U1215 (N_1215,In_1939,In_2194);
or U1216 (N_1216,In_1840,In_1354);
and U1217 (N_1217,In_793,In_737);
nor U1218 (N_1218,In_485,In_1675);
nor U1219 (N_1219,In_1079,In_530);
and U1220 (N_1220,In_1654,In_2449);
nor U1221 (N_1221,In_723,In_994);
xor U1222 (N_1222,In_1398,In_1492);
nor U1223 (N_1223,In_1773,In_1341);
and U1224 (N_1224,In_615,In_2191);
and U1225 (N_1225,In_1001,In_1478);
or U1226 (N_1226,In_1164,In_2003);
or U1227 (N_1227,In_2450,In_1884);
or U1228 (N_1228,In_1528,In_998);
nand U1229 (N_1229,In_1144,In_2051);
and U1230 (N_1230,In_730,In_2115);
nand U1231 (N_1231,In_588,In_635);
or U1232 (N_1232,In_518,In_1116);
xnor U1233 (N_1233,In_1384,In_1908);
and U1234 (N_1234,In_2242,In_895);
and U1235 (N_1235,In_685,In_2111);
and U1236 (N_1236,In_947,In_1751);
or U1237 (N_1237,In_1786,In_2461);
nand U1238 (N_1238,In_1368,In_1563);
nor U1239 (N_1239,In_536,In_341);
xor U1240 (N_1240,In_1529,In_1279);
or U1241 (N_1241,In_1099,In_504);
xnor U1242 (N_1242,In_1926,In_411);
or U1243 (N_1243,In_734,In_1403);
nand U1244 (N_1244,In_1580,In_151);
and U1245 (N_1245,In_788,In_1512);
and U1246 (N_1246,In_1461,In_603);
xor U1247 (N_1247,In_1603,In_1220);
xnor U1248 (N_1248,In_2498,In_360);
xor U1249 (N_1249,In_1606,In_743);
nor U1250 (N_1250,In_1874,In_252);
and U1251 (N_1251,In_423,In_1619);
nand U1252 (N_1252,In_1097,In_958);
and U1253 (N_1253,In_1122,In_2316);
nor U1254 (N_1254,In_993,In_142);
xor U1255 (N_1255,In_1171,In_1845);
nor U1256 (N_1256,In_1982,In_1036);
or U1257 (N_1257,In_277,In_409);
xor U1258 (N_1258,In_2116,In_691);
nor U1259 (N_1259,In_235,In_25);
nand U1260 (N_1260,In_644,In_1623);
and U1261 (N_1261,In_1017,In_218);
nor U1262 (N_1262,In_2304,In_231);
or U1263 (N_1263,In_2145,In_219);
xnor U1264 (N_1264,In_189,In_2236);
nor U1265 (N_1265,In_668,In_1803);
nand U1266 (N_1266,In_661,In_1433);
or U1267 (N_1267,In_1478,In_1715);
nand U1268 (N_1268,In_1476,In_2056);
and U1269 (N_1269,In_635,In_2307);
and U1270 (N_1270,In_1562,In_1247);
nand U1271 (N_1271,In_1535,In_1339);
and U1272 (N_1272,In_290,In_152);
xnor U1273 (N_1273,In_2358,In_1859);
xor U1274 (N_1274,In_2254,In_263);
xor U1275 (N_1275,In_640,In_1124);
nand U1276 (N_1276,In_2286,In_2437);
nor U1277 (N_1277,In_341,In_976);
xor U1278 (N_1278,In_829,In_1459);
xor U1279 (N_1279,In_1453,In_96);
xnor U1280 (N_1280,In_1686,In_1880);
or U1281 (N_1281,In_2352,In_1899);
xor U1282 (N_1282,In_755,In_2224);
xnor U1283 (N_1283,In_697,In_1974);
and U1284 (N_1284,In_2025,In_1852);
or U1285 (N_1285,In_1222,In_1829);
nand U1286 (N_1286,In_1033,In_1975);
nand U1287 (N_1287,In_933,In_1083);
nand U1288 (N_1288,In_462,In_2109);
and U1289 (N_1289,In_1115,In_2034);
nand U1290 (N_1290,In_1465,In_1201);
or U1291 (N_1291,In_70,In_981);
or U1292 (N_1292,In_354,In_979);
and U1293 (N_1293,In_799,In_949);
or U1294 (N_1294,In_922,In_970);
and U1295 (N_1295,In_1674,In_122);
and U1296 (N_1296,In_1762,In_5);
and U1297 (N_1297,In_645,In_2497);
nand U1298 (N_1298,In_810,In_2360);
and U1299 (N_1299,In_2338,In_673);
or U1300 (N_1300,In_299,In_2060);
nand U1301 (N_1301,In_854,In_1461);
nor U1302 (N_1302,In_1127,In_506);
xnor U1303 (N_1303,In_27,In_2341);
and U1304 (N_1304,In_1576,In_780);
nand U1305 (N_1305,In_2099,In_595);
or U1306 (N_1306,In_0,In_624);
xor U1307 (N_1307,In_843,In_382);
nand U1308 (N_1308,In_1444,In_1886);
or U1309 (N_1309,In_763,In_895);
xnor U1310 (N_1310,In_57,In_1375);
xor U1311 (N_1311,In_840,In_2458);
nor U1312 (N_1312,In_324,In_1636);
nor U1313 (N_1313,In_1071,In_893);
and U1314 (N_1314,In_699,In_217);
nor U1315 (N_1315,In_2001,In_602);
nand U1316 (N_1316,In_172,In_1600);
nor U1317 (N_1317,In_1209,In_2121);
nand U1318 (N_1318,In_92,In_2043);
xor U1319 (N_1319,In_2256,In_668);
or U1320 (N_1320,In_99,In_981);
xor U1321 (N_1321,In_2497,In_2016);
nand U1322 (N_1322,In_1201,In_1545);
and U1323 (N_1323,In_731,In_1019);
nand U1324 (N_1324,In_2478,In_366);
nand U1325 (N_1325,In_1747,In_240);
nand U1326 (N_1326,In_1971,In_1681);
or U1327 (N_1327,In_2062,In_1109);
nand U1328 (N_1328,In_320,In_363);
nor U1329 (N_1329,In_788,In_1845);
and U1330 (N_1330,In_87,In_689);
or U1331 (N_1331,In_1420,In_665);
or U1332 (N_1332,In_1744,In_1215);
nor U1333 (N_1333,In_889,In_262);
xnor U1334 (N_1334,In_397,In_2488);
or U1335 (N_1335,In_129,In_1075);
or U1336 (N_1336,In_1237,In_1286);
nor U1337 (N_1337,In_1783,In_1046);
nand U1338 (N_1338,In_317,In_1567);
nor U1339 (N_1339,In_152,In_1721);
nor U1340 (N_1340,In_1802,In_177);
xnor U1341 (N_1341,In_195,In_854);
xnor U1342 (N_1342,In_906,In_2301);
nand U1343 (N_1343,In_472,In_974);
xnor U1344 (N_1344,In_1684,In_2018);
or U1345 (N_1345,In_116,In_1892);
and U1346 (N_1346,In_1667,In_2413);
or U1347 (N_1347,In_633,In_1520);
xor U1348 (N_1348,In_2167,In_968);
xor U1349 (N_1349,In_148,In_200);
nor U1350 (N_1350,In_1852,In_1114);
and U1351 (N_1351,In_1217,In_344);
nand U1352 (N_1352,In_2147,In_1657);
and U1353 (N_1353,In_51,In_2043);
nand U1354 (N_1354,In_497,In_121);
nor U1355 (N_1355,In_554,In_2206);
and U1356 (N_1356,In_1545,In_810);
xnor U1357 (N_1357,In_2374,In_2041);
or U1358 (N_1358,In_1054,In_2292);
or U1359 (N_1359,In_1200,In_986);
nor U1360 (N_1360,In_1330,In_1020);
and U1361 (N_1361,In_1459,In_2215);
nand U1362 (N_1362,In_474,In_182);
or U1363 (N_1363,In_2197,In_2497);
and U1364 (N_1364,In_64,In_2464);
xor U1365 (N_1365,In_762,In_178);
nand U1366 (N_1366,In_1436,In_2208);
nor U1367 (N_1367,In_2239,In_545);
nor U1368 (N_1368,In_1915,In_1253);
nand U1369 (N_1369,In_1304,In_1327);
or U1370 (N_1370,In_2185,In_1029);
nor U1371 (N_1371,In_1809,In_302);
nor U1372 (N_1372,In_2309,In_177);
xor U1373 (N_1373,In_1779,In_670);
nand U1374 (N_1374,In_168,In_124);
xor U1375 (N_1375,In_2111,In_75);
or U1376 (N_1376,In_1680,In_2044);
nand U1377 (N_1377,In_2168,In_255);
or U1378 (N_1378,In_2039,In_1414);
and U1379 (N_1379,In_1417,In_1688);
or U1380 (N_1380,In_1611,In_804);
xor U1381 (N_1381,In_1768,In_637);
nor U1382 (N_1382,In_1542,In_1852);
nor U1383 (N_1383,In_1935,In_120);
and U1384 (N_1384,In_2295,In_1024);
nor U1385 (N_1385,In_2124,In_166);
nand U1386 (N_1386,In_1462,In_541);
nor U1387 (N_1387,In_1190,In_2044);
nor U1388 (N_1388,In_2246,In_136);
xnor U1389 (N_1389,In_2237,In_1156);
or U1390 (N_1390,In_1297,In_502);
or U1391 (N_1391,In_2262,In_2116);
or U1392 (N_1392,In_2190,In_741);
and U1393 (N_1393,In_1606,In_765);
nand U1394 (N_1394,In_1363,In_418);
nor U1395 (N_1395,In_1358,In_617);
nand U1396 (N_1396,In_959,In_842);
nor U1397 (N_1397,In_2396,In_1977);
nand U1398 (N_1398,In_230,In_2205);
nor U1399 (N_1399,In_2157,In_2442);
and U1400 (N_1400,In_1142,In_1290);
nor U1401 (N_1401,In_952,In_627);
nor U1402 (N_1402,In_1608,In_1880);
xnor U1403 (N_1403,In_873,In_754);
or U1404 (N_1404,In_2439,In_1697);
nor U1405 (N_1405,In_2180,In_2198);
xnor U1406 (N_1406,In_723,In_2091);
nand U1407 (N_1407,In_1036,In_1489);
nor U1408 (N_1408,In_198,In_532);
and U1409 (N_1409,In_838,In_264);
nor U1410 (N_1410,In_1338,In_46);
xnor U1411 (N_1411,In_1192,In_2237);
xnor U1412 (N_1412,In_2407,In_717);
or U1413 (N_1413,In_1103,In_1031);
or U1414 (N_1414,In_1077,In_2171);
nor U1415 (N_1415,In_1252,In_1388);
nand U1416 (N_1416,In_1382,In_1186);
nor U1417 (N_1417,In_1779,In_1088);
xnor U1418 (N_1418,In_1337,In_1098);
or U1419 (N_1419,In_1477,In_628);
xor U1420 (N_1420,In_1759,In_1868);
xnor U1421 (N_1421,In_447,In_1218);
or U1422 (N_1422,In_115,In_1955);
or U1423 (N_1423,In_1551,In_1434);
nand U1424 (N_1424,In_621,In_805);
and U1425 (N_1425,In_991,In_652);
nand U1426 (N_1426,In_655,In_1685);
and U1427 (N_1427,In_2377,In_1232);
nand U1428 (N_1428,In_595,In_2218);
and U1429 (N_1429,In_2331,In_406);
nor U1430 (N_1430,In_1389,In_2309);
and U1431 (N_1431,In_1835,In_1552);
or U1432 (N_1432,In_523,In_634);
and U1433 (N_1433,In_613,In_789);
nand U1434 (N_1434,In_1029,In_20);
and U1435 (N_1435,In_2411,In_385);
nor U1436 (N_1436,In_1718,In_2255);
nand U1437 (N_1437,In_1424,In_1970);
nand U1438 (N_1438,In_2345,In_2044);
nor U1439 (N_1439,In_2118,In_1416);
nor U1440 (N_1440,In_336,In_1234);
nand U1441 (N_1441,In_1774,In_1570);
xnor U1442 (N_1442,In_548,In_1875);
and U1443 (N_1443,In_1107,In_1054);
and U1444 (N_1444,In_1468,In_195);
or U1445 (N_1445,In_1633,In_1298);
or U1446 (N_1446,In_418,In_2291);
xnor U1447 (N_1447,In_97,In_2481);
nor U1448 (N_1448,In_830,In_1363);
nor U1449 (N_1449,In_1905,In_1779);
nand U1450 (N_1450,In_529,In_528);
xnor U1451 (N_1451,In_1944,In_618);
nand U1452 (N_1452,In_689,In_845);
nand U1453 (N_1453,In_2434,In_118);
or U1454 (N_1454,In_2311,In_1138);
xor U1455 (N_1455,In_247,In_2311);
and U1456 (N_1456,In_16,In_1709);
nor U1457 (N_1457,In_2330,In_237);
and U1458 (N_1458,In_2327,In_976);
xor U1459 (N_1459,In_2239,In_1442);
nor U1460 (N_1460,In_2181,In_2454);
or U1461 (N_1461,In_66,In_1542);
xnor U1462 (N_1462,In_390,In_255);
or U1463 (N_1463,In_2331,In_236);
nor U1464 (N_1464,In_609,In_1851);
and U1465 (N_1465,In_2093,In_1266);
nor U1466 (N_1466,In_2386,In_2069);
or U1467 (N_1467,In_2325,In_1169);
and U1468 (N_1468,In_2100,In_591);
xnor U1469 (N_1469,In_1640,In_687);
nand U1470 (N_1470,In_1432,In_1385);
and U1471 (N_1471,In_1820,In_490);
and U1472 (N_1472,In_2025,In_1441);
and U1473 (N_1473,In_325,In_2135);
nand U1474 (N_1474,In_1578,In_341);
xnor U1475 (N_1475,In_1353,In_2460);
or U1476 (N_1476,In_1841,In_800);
xnor U1477 (N_1477,In_2339,In_1016);
or U1478 (N_1478,In_1251,In_1532);
or U1479 (N_1479,In_2434,In_473);
nor U1480 (N_1480,In_1689,In_1791);
or U1481 (N_1481,In_1299,In_1804);
nor U1482 (N_1482,In_922,In_689);
and U1483 (N_1483,In_784,In_1063);
or U1484 (N_1484,In_1370,In_2445);
nand U1485 (N_1485,In_169,In_1748);
nor U1486 (N_1486,In_2000,In_237);
nor U1487 (N_1487,In_17,In_2430);
nor U1488 (N_1488,In_629,In_962);
or U1489 (N_1489,In_6,In_620);
nand U1490 (N_1490,In_825,In_1202);
nor U1491 (N_1491,In_1817,In_841);
and U1492 (N_1492,In_1610,In_1415);
or U1493 (N_1493,In_166,In_2232);
nand U1494 (N_1494,In_141,In_1834);
nor U1495 (N_1495,In_1476,In_29);
xor U1496 (N_1496,In_660,In_2449);
and U1497 (N_1497,In_686,In_1838);
and U1498 (N_1498,In_369,In_258);
nand U1499 (N_1499,In_249,In_1070);
nand U1500 (N_1500,In_1282,In_1437);
and U1501 (N_1501,In_2125,In_1818);
or U1502 (N_1502,In_741,In_189);
xnor U1503 (N_1503,In_1606,In_489);
nand U1504 (N_1504,In_2186,In_439);
or U1505 (N_1505,In_2477,In_237);
nor U1506 (N_1506,In_1387,In_2462);
nor U1507 (N_1507,In_1546,In_1875);
and U1508 (N_1508,In_2306,In_700);
or U1509 (N_1509,In_1411,In_1722);
and U1510 (N_1510,In_1445,In_2001);
nand U1511 (N_1511,In_1146,In_953);
or U1512 (N_1512,In_392,In_25);
or U1513 (N_1513,In_463,In_446);
nor U1514 (N_1514,In_22,In_1273);
xor U1515 (N_1515,In_2421,In_1418);
xnor U1516 (N_1516,In_1853,In_1131);
or U1517 (N_1517,In_1546,In_538);
nor U1518 (N_1518,In_244,In_355);
nand U1519 (N_1519,In_2027,In_440);
xnor U1520 (N_1520,In_945,In_1603);
and U1521 (N_1521,In_1628,In_1528);
nor U1522 (N_1522,In_1559,In_2176);
xnor U1523 (N_1523,In_2484,In_2387);
and U1524 (N_1524,In_2150,In_2259);
xor U1525 (N_1525,In_14,In_104);
and U1526 (N_1526,In_948,In_824);
nand U1527 (N_1527,In_1857,In_2245);
nand U1528 (N_1528,In_1404,In_1495);
nand U1529 (N_1529,In_640,In_1088);
nor U1530 (N_1530,In_1306,In_1687);
nand U1531 (N_1531,In_347,In_1617);
xor U1532 (N_1532,In_769,In_241);
or U1533 (N_1533,In_1884,In_112);
nor U1534 (N_1534,In_1290,In_26);
nor U1535 (N_1535,In_1586,In_78);
nor U1536 (N_1536,In_1249,In_516);
nand U1537 (N_1537,In_2324,In_1464);
and U1538 (N_1538,In_1035,In_1821);
nand U1539 (N_1539,In_130,In_1581);
or U1540 (N_1540,In_1268,In_727);
or U1541 (N_1541,In_1446,In_648);
nor U1542 (N_1542,In_434,In_2374);
and U1543 (N_1543,In_1547,In_2395);
xor U1544 (N_1544,In_822,In_2388);
xnor U1545 (N_1545,In_338,In_1851);
nor U1546 (N_1546,In_25,In_1128);
nor U1547 (N_1547,In_179,In_1147);
nand U1548 (N_1548,In_1714,In_2100);
xnor U1549 (N_1549,In_2075,In_2335);
and U1550 (N_1550,In_545,In_945);
xnor U1551 (N_1551,In_1666,In_1174);
or U1552 (N_1552,In_1043,In_1805);
and U1553 (N_1553,In_556,In_2329);
xnor U1554 (N_1554,In_2283,In_1927);
nor U1555 (N_1555,In_556,In_100);
xnor U1556 (N_1556,In_1061,In_103);
and U1557 (N_1557,In_849,In_1763);
xor U1558 (N_1558,In_479,In_850);
and U1559 (N_1559,In_1222,In_591);
nand U1560 (N_1560,In_327,In_2128);
nor U1561 (N_1561,In_1925,In_398);
nand U1562 (N_1562,In_2459,In_954);
xor U1563 (N_1563,In_2313,In_2115);
or U1564 (N_1564,In_2315,In_937);
xor U1565 (N_1565,In_2028,In_550);
and U1566 (N_1566,In_1855,In_2382);
or U1567 (N_1567,In_1779,In_324);
and U1568 (N_1568,In_1653,In_2028);
and U1569 (N_1569,In_1968,In_1157);
xnor U1570 (N_1570,In_2298,In_1309);
nor U1571 (N_1571,In_2488,In_2074);
and U1572 (N_1572,In_324,In_896);
nor U1573 (N_1573,In_1913,In_2228);
xor U1574 (N_1574,In_1230,In_711);
xnor U1575 (N_1575,In_737,In_2070);
xnor U1576 (N_1576,In_1237,In_303);
nor U1577 (N_1577,In_877,In_656);
xor U1578 (N_1578,In_780,In_244);
nor U1579 (N_1579,In_230,In_2483);
nand U1580 (N_1580,In_97,In_765);
or U1581 (N_1581,In_1233,In_1873);
nand U1582 (N_1582,In_1532,In_2148);
nand U1583 (N_1583,In_204,In_2404);
and U1584 (N_1584,In_112,In_2443);
xnor U1585 (N_1585,In_1179,In_2209);
or U1586 (N_1586,In_426,In_2215);
xnor U1587 (N_1587,In_683,In_1492);
or U1588 (N_1588,In_2153,In_1638);
nand U1589 (N_1589,In_1289,In_2297);
xor U1590 (N_1590,In_1863,In_635);
or U1591 (N_1591,In_2086,In_354);
or U1592 (N_1592,In_1115,In_2027);
and U1593 (N_1593,In_1555,In_434);
and U1594 (N_1594,In_1658,In_979);
and U1595 (N_1595,In_269,In_931);
and U1596 (N_1596,In_822,In_352);
nor U1597 (N_1597,In_499,In_2471);
nand U1598 (N_1598,In_749,In_2279);
xnor U1599 (N_1599,In_1985,In_1028);
or U1600 (N_1600,In_1596,In_2084);
and U1601 (N_1601,In_1019,In_2141);
nand U1602 (N_1602,In_2355,In_2229);
nand U1603 (N_1603,In_543,In_1529);
and U1604 (N_1604,In_1978,In_1849);
nor U1605 (N_1605,In_378,In_192);
or U1606 (N_1606,In_2209,In_758);
or U1607 (N_1607,In_383,In_1961);
nor U1608 (N_1608,In_185,In_1464);
nor U1609 (N_1609,In_350,In_137);
or U1610 (N_1610,In_1782,In_1692);
nor U1611 (N_1611,In_762,In_192);
xnor U1612 (N_1612,In_658,In_111);
nand U1613 (N_1613,In_2433,In_75);
or U1614 (N_1614,In_1367,In_745);
xor U1615 (N_1615,In_1747,In_2329);
or U1616 (N_1616,In_2094,In_422);
or U1617 (N_1617,In_808,In_1022);
or U1618 (N_1618,In_2234,In_180);
nand U1619 (N_1619,In_2438,In_2132);
and U1620 (N_1620,In_710,In_1922);
nor U1621 (N_1621,In_927,In_2340);
nor U1622 (N_1622,In_1684,In_722);
nand U1623 (N_1623,In_1499,In_2076);
and U1624 (N_1624,In_1689,In_2140);
nor U1625 (N_1625,In_221,In_2349);
or U1626 (N_1626,In_333,In_353);
nand U1627 (N_1627,In_2171,In_501);
and U1628 (N_1628,In_408,In_1078);
and U1629 (N_1629,In_167,In_2482);
or U1630 (N_1630,In_171,In_1993);
and U1631 (N_1631,In_2251,In_1242);
xnor U1632 (N_1632,In_1441,In_1502);
xor U1633 (N_1633,In_1020,In_924);
xor U1634 (N_1634,In_2039,In_398);
nor U1635 (N_1635,In_1815,In_1457);
xor U1636 (N_1636,In_122,In_1288);
xnor U1637 (N_1637,In_2039,In_1782);
xnor U1638 (N_1638,In_2226,In_491);
nor U1639 (N_1639,In_936,In_2045);
xor U1640 (N_1640,In_2254,In_2494);
and U1641 (N_1641,In_1158,In_550);
nor U1642 (N_1642,In_77,In_2195);
nor U1643 (N_1643,In_2356,In_1258);
and U1644 (N_1644,In_238,In_1944);
xnor U1645 (N_1645,In_1739,In_419);
and U1646 (N_1646,In_2387,In_1159);
xor U1647 (N_1647,In_2299,In_932);
nor U1648 (N_1648,In_2494,In_1189);
xor U1649 (N_1649,In_622,In_94);
and U1650 (N_1650,In_33,In_34);
and U1651 (N_1651,In_762,In_2079);
or U1652 (N_1652,In_505,In_1523);
and U1653 (N_1653,In_915,In_2056);
xor U1654 (N_1654,In_1082,In_2469);
nor U1655 (N_1655,In_114,In_944);
or U1656 (N_1656,In_536,In_405);
nor U1657 (N_1657,In_837,In_1393);
or U1658 (N_1658,In_949,In_1118);
nor U1659 (N_1659,In_1646,In_2302);
nand U1660 (N_1660,In_1242,In_1597);
xor U1661 (N_1661,In_961,In_1325);
or U1662 (N_1662,In_589,In_2158);
and U1663 (N_1663,In_1119,In_84);
xor U1664 (N_1664,In_324,In_1344);
or U1665 (N_1665,In_401,In_147);
nor U1666 (N_1666,In_605,In_1804);
nor U1667 (N_1667,In_910,In_387);
or U1668 (N_1668,In_1756,In_49);
or U1669 (N_1669,In_566,In_2464);
nor U1670 (N_1670,In_635,In_974);
nand U1671 (N_1671,In_1048,In_1977);
or U1672 (N_1672,In_1981,In_2337);
nand U1673 (N_1673,In_637,In_1519);
xor U1674 (N_1674,In_2038,In_1244);
xor U1675 (N_1675,In_919,In_911);
xnor U1676 (N_1676,In_683,In_1792);
xor U1677 (N_1677,In_324,In_1842);
nand U1678 (N_1678,In_776,In_2392);
or U1679 (N_1679,In_779,In_430);
nor U1680 (N_1680,In_547,In_561);
nand U1681 (N_1681,In_2226,In_2424);
xor U1682 (N_1682,In_228,In_1321);
and U1683 (N_1683,In_1584,In_948);
nor U1684 (N_1684,In_1301,In_13);
and U1685 (N_1685,In_1066,In_1596);
nand U1686 (N_1686,In_303,In_1529);
nor U1687 (N_1687,In_731,In_1565);
or U1688 (N_1688,In_223,In_611);
nor U1689 (N_1689,In_408,In_1725);
and U1690 (N_1690,In_445,In_1200);
nand U1691 (N_1691,In_458,In_1256);
nor U1692 (N_1692,In_2308,In_884);
or U1693 (N_1693,In_799,In_1035);
xnor U1694 (N_1694,In_1798,In_1553);
nand U1695 (N_1695,In_2228,In_1226);
and U1696 (N_1696,In_924,In_1406);
or U1697 (N_1697,In_7,In_1044);
xor U1698 (N_1698,In_932,In_1316);
nor U1699 (N_1699,In_113,In_263);
or U1700 (N_1700,In_1752,In_529);
and U1701 (N_1701,In_1239,In_283);
nand U1702 (N_1702,In_767,In_1526);
or U1703 (N_1703,In_467,In_2432);
nor U1704 (N_1704,In_67,In_1463);
nor U1705 (N_1705,In_1082,In_2005);
nand U1706 (N_1706,In_1152,In_2443);
nand U1707 (N_1707,In_768,In_1680);
nand U1708 (N_1708,In_604,In_2058);
and U1709 (N_1709,In_61,In_1776);
nor U1710 (N_1710,In_1797,In_676);
or U1711 (N_1711,In_917,In_322);
nor U1712 (N_1712,In_781,In_2398);
nand U1713 (N_1713,In_310,In_754);
xor U1714 (N_1714,In_1164,In_1576);
nor U1715 (N_1715,In_150,In_1403);
or U1716 (N_1716,In_920,In_236);
or U1717 (N_1717,In_617,In_288);
nand U1718 (N_1718,In_1833,In_492);
xnor U1719 (N_1719,In_409,In_2397);
xor U1720 (N_1720,In_686,In_1133);
and U1721 (N_1721,In_1359,In_1882);
and U1722 (N_1722,In_639,In_301);
xnor U1723 (N_1723,In_2345,In_983);
nor U1724 (N_1724,In_437,In_597);
nor U1725 (N_1725,In_1312,In_203);
nand U1726 (N_1726,In_1191,In_1715);
and U1727 (N_1727,In_1111,In_2);
xor U1728 (N_1728,In_1593,In_617);
and U1729 (N_1729,In_313,In_789);
nand U1730 (N_1730,In_1797,In_2141);
nand U1731 (N_1731,In_1880,In_1649);
xnor U1732 (N_1732,In_1849,In_1738);
nand U1733 (N_1733,In_2177,In_1842);
or U1734 (N_1734,In_2126,In_2429);
or U1735 (N_1735,In_1646,In_774);
xnor U1736 (N_1736,In_1464,In_605);
nor U1737 (N_1737,In_1090,In_2408);
nand U1738 (N_1738,In_2164,In_1151);
nand U1739 (N_1739,In_242,In_636);
and U1740 (N_1740,In_243,In_792);
nand U1741 (N_1741,In_2373,In_258);
nor U1742 (N_1742,In_316,In_1967);
nand U1743 (N_1743,In_1433,In_1906);
xor U1744 (N_1744,In_453,In_1472);
nor U1745 (N_1745,In_1823,In_2286);
and U1746 (N_1746,In_1091,In_533);
xor U1747 (N_1747,In_817,In_298);
nand U1748 (N_1748,In_2095,In_1829);
or U1749 (N_1749,In_797,In_343);
or U1750 (N_1750,In_330,In_1569);
or U1751 (N_1751,In_1240,In_1172);
nor U1752 (N_1752,In_1402,In_754);
nand U1753 (N_1753,In_1882,In_1082);
nand U1754 (N_1754,In_1748,In_364);
and U1755 (N_1755,In_669,In_1625);
and U1756 (N_1756,In_1768,In_1016);
nand U1757 (N_1757,In_1665,In_106);
xnor U1758 (N_1758,In_2451,In_1198);
or U1759 (N_1759,In_2302,In_1352);
and U1760 (N_1760,In_2201,In_490);
nor U1761 (N_1761,In_2332,In_72);
nor U1762 (N_1762,In_1576,In_1432);
or U1763 (N_1763,In_1598,In_596);
xnor U1764 (N_1764,In_1868,In_1649);
nand U1765 (N_1765,In_271,In_2009);
or U1766 (N_1766,In_125,In_634);
nand U1767 (N_1767,In_1656,In_1553);
or U1768 (N_1768,In_1186,In_443);
xnor U1769 (N_1769,In_672,In_1946);
nand U1770 (N_1770,In_345,In_858);
nor U1771 (N_1771,In_463,In_2057);
xnor U1772 (N_1772,In_789,In_1577);
nor U1773 (N_1773,In_888,In_1485);
nand U1774 (N_1774,In_1996,In_2332);
nor U1775 (N_1775,In_1245,In_719);
nand U1776 (N_1776,In_1385,In_2162);
xor U1777 (N_1777,In_843,In_1964);
xnor U1778 (N_1778,In_1867,In_2448);
and U1779 (N_1779,In_1628,In_1401);
xor U1780 (N_1780,In_1339,In_147);
xor U1781 (N_1781,In_1030,In_2250);
nor U1782 (N_1782,In_2420,In_876);
or U1783 (N_1783,In_1584,In_945);
or U1784 (N_1784,In_391,In_2277);
xnor U1785 (N_1785,In_1468,In_2435);
and U1786 (N_1786,In_1297,In_1537);
or U1787 (N_1787,In_1352,In_237);
xnor U1788 (N_1788,In_454,In_823);
nor U1789 (N_1789,In_1702,In_1317);
nor U1790 (N_1790,In_22,In_1134);
or U1791 (N_1791,In_1975,In_799);
and U1792 (N_1792,In_1891,In_2315);
nand U1793 (N_1793,In_1421,In_2095);
and U1794 (N_1794,In_1765,In_679);
xor U1795 (N_1795,In_288,In_1304);
nor U1796 (N_1796,In_1124,In_468);
nor U1797 (N_1797,In_1378,In_125);
xor U1798 (N_1798,In_1532,In_2023);
or U1799 (N_1799,In_1157,In_1329);
and U1800 (N_1800,In_1782,In_146);
nand U1801 (N_1801,In_617,In_46);
or U1802 (N_1802,In_1664,In_1700);
nand U1803 (N_1803,In_694,In_1208);
or U1804 (N_1804,In_1233,In_2248);
or U1805 (N_1805,In_456,In_2044);
and U1806 (N_1806,In_815,In_963);
or U1807 (N_1807,In_1432,In_1783);
nand U1808 (N_1808,In_2139,In_750);
or U1809 (N_1809,In_645,In_1356);
xnor U1810 (N_1810,In_247,In_1884);
xnor U1811 (N_1811,In_1711,In_1950);
and U1812 (N_1812,In_2459,In_1174);
xor U1813 (N_1813,In_162,In_1274);
and U1814 (N_1814,In_2404,In_1508);
and U1815 (N_1815,In_1613,In_758);
xnor U1816 (N_1816,In_1007,In_2391);
nor U1817 (N_1817,In_2422,In_1527);
nor U1818 (N_1818,In_2361,In_1109);
nor U1819 (N_1819,In_615,In_2426);
nor U1820 (N_1820,In_1575,In_2120);
or U1821 (N_1821,In_795,In_1041);
xor U1822 (N_1822,In_572,In_501);
nor U1823 (N_1823,In_326,In_359);
nor U1824 (N_1824,In_2381,In_718);
nor U1825 (N_1825,In_1802,In_624);
nor U1826 (N_1826,In_1235,In_1164);
nand U1827 (N_1827,In_1828,In_1639);
nor U1828 (N_1828,In_563,In_2265);
or U1829 (N_1829,In_521,In_1408);
xor U1830 (N_1830,In_1402,In_1474);
xnor U1831 (N_1831,In_644,In_1021);
and U1832 (N_1832,In_168,In_1950);
nand U1833 (N_1833,In_1572,In_1077);
or U1834 (N_1834,In_844,In_1802);
xnor U1835 (N_1835,In_2204,In_2172);
xor U1836 (N_1836,In_2080,In_559);
nand U1837 (N_1837,In_51,In_724);
and U1838 (N_1838,In_640,In_1142);
and U1839 (N_1839,In_965,In_462);
nand U1840 (N_1840,In_425,In_634);
nor U1841 (N_1841,In_2081,In_1956);
nand U1842 (N_1842,In_982,In_790);
and U1843 (N_1843,In_1754,In_2202);
nand U1844 (N_1844,In_324,In_1724);
nand U1845 (N_1845,In_121,In_1501);
nand U1846 (N_1846,In_2029,In_961);
xor U1847 (N_1847,In_818,In_772);
and U1848 (N_1848,In_1295,In_642);
nor U1849 (N_1849,In_2481,In_1494);
nand U1850 (N_1850,In_825,In_520);
or U1851 (N_1851,In_578,In_1823);
or U1852 (N_1852,In_235,In_970);
nand U1853 (N_1853,In_1066,In_1808);
nor U1854 (N_1854,In_2335,In_1743);
and U1855 (N_1855,In_1901,In_506);
xor U1856 (N_1856,In_2227,In_2100);
xor U1857 (N_1857,In_27,In_1747);
nand U1858 (N_1858,In_2249,In_326);
xnor U1859 (N_1859,In_1689,In_451);
and U1860 (N_1860,In_2279,In_118);
nand U1861 (N_1861,In_1196,In_1484);
nor U1862 (N_1862,In_267,In_1381);
and U1863 (N_1863,In_249,In_1297);
and U1864 (N_1864,In_697,In_716);
and U1865 (N_1865,In_1572,In_1627);
or U1866 (N_1866,In_1982,In_1072);
or U1867 (N_1867,In_510,In_363);
xor U1868 (N_1868,In_651,In_738);
or U1869 (N_1869,In_2139,In_1980);
or U1870 (N_1870,In_731,In_996);
xnor U1871 (N_1871,In_2303,In_1354);
xor U1872 (N_1872,In_2479,In_474);
or U1873 (N_1873,In_975,In_2333);
nor U1874 (N_1874,In_1682,In_1369);
nand U1875 (N_1875,In_127,In_614);
or U1876 (N_1876,In_1644,In_849);
nor U1877 (N_1877,In_334,In_2467);
nand U1878 (N_1878,In_948,In_786);
or U1879 (N_1879,In_2045,In_2292);
nor U1880 (N_1880,In_549,In_1784);
xor U1881 (N_1881,In_77,In_85);
nor U1882 (N_1882,In_1281,In_1997);
and U1883 (N_1883,In_790,In_1720);
nand U1884 (N_1884,In_1247,In_28);
nand U1885 (N_1885,In_2229,In_493);
and U1886 (N_1886,In_176,In_49);
or U1887 (N_1887,In_941,In_1557);
and U1888 (N_1888,In_139,In_546);
or U1889 (N_1889,In_1316,In_1740);
and U1890 (N_1890,In_1709,In_1657);
xor U1891 (N_1891,In_1172,In_895);
xor U1892 (N_1892,In_583,In_2354);
nor U1893 (N_1893,In_1960,In_1402);
xnor U1894 (N_1894,In_1688,In_1012);
xnor U1895 (N_1895,In_1097,In_1322);
nor U1896 (N_1896,In_1960,In_1070);
or U1897 (N_1897,In_2424,In_1479);
or U1898 (N_1898,In_2081,In_1563);
nand U1899 (N_1899,In_942,In_2427);
xor U1900 (N_1900,In_1676,In_285);
nor U1901 (N_1901,In_1216,In_193);
or U1902 (N_1902,In_2281,In_610);
nor U1903 (N_1903,In_1468,In_77);
or U1904 (N_1904,In_1899,In_1169);
or U1905 (N_1905,In_1969,In_1179);
xor U1906 (N_1906,In_120,In_925);
nor U1907 (N_1907,In_1383,In_666);
nor U1908 (N_1908,In_474,In_346);
xnor U1909 (N_1909,In_2471,In_1016);
and U1910 (N_1910,In_2327,In_2193);
nor U1911 (N_1911,In_1171,In_2145);
or U1912 (N_1912,In_2210,In_143);
nor U1913 (N_1913,In_105,In_1362);
nand U1914 (N_1914,In_244,In_1449);
or U1915 (N_1915,In_1576,In_953);
nor U1916 (N_1916,In_2341,In_833);
nor U1917 (N_1917,In_2356,In_1233);
and U1918 (N_1918,In_778,In_2258);
nor U1919 (N_1919,In_52,In_2356);
nand U1920 (N_1920,In_2435,In_2087);
nor U1921 (N_1921,In_1137,In_2302);
nand U1922 (N_1922,In_638,In_1701);
nand U1923 (N_1923,In_816,In_1388);
and U1924 (N_1924,In_1216,In_1005);
and U1925 (N_1925,In_870,In_1828);
nor U1926 (N_1926,In_1019,In_311);
nand U1927 (N_1927,In_488,In_1588);
nand U1928 (N_1928,In_2147,In_2429);
nand U1929 (N_1929,In_474,In_1840);
or U1930 (N_1930,In_1805,In_2210);
nor U1931 (N_1931,In_2134,In_557);
or U1932 (N_1932,In_818,In_417);
xnor U1933 (N_1933,In_1942,In_1084);
or U1934 (N_1934,In_155,In_2339);
nand U1935 (N_1935,In_522,In_2454);
and U1936 (N_1936,In_49,In_2425);
nor U1937 (N_1937,In_1030,In_2009);
or U1938 (N_1938,In_617,In_1439);
and U1939 (N_1939,In_2362,In_1524);
and U1940 (N_1940,In_2250,In_258);
xor U1941 (N_1941,In_1395,In_1104);
nand U1942 (N_1942,In_248,In_1351);
nor U1943 (N_1943,In_1794,In_1123);
xor U1944 (N_1944,In_629,In_266);
nand U1945 (N_1945,In_958,In_1616);
nand U1946 (N_1946,In_657,In_2081);
nor U1947 (N_1947,In_1520,In_2275);
xor U1948 (N_1948,In_2285,In_2400);
nand U1949 (N_1949,In_2453,In_2367);
xnor U1950 (N_1950,In_1364,In_145);
and U1951 (N_1951,In_2314,In_1775);
and U1952 (N_1952,In_892,In_1976);
xor U1953 (N_1953,In_1449,In_756);
xnor U1954 (N_1954,In_67,In_2215);
nor U1955 (N_1955,In_32,In_105);
nor U1956 (N_1956,In_939,In_2171);
and U1957 (N_1957,In_248,In_2078);
xor U1958 (N_1958,In_885,In_1674);
nor U1959 (N_1959,In_20,In_1952);
and U1960 (N_1960,In_1263,In_1210);
xnor U1961 (N_1961,In_1882,In_2377);
xor U1962 (N_1962,In_530,In_1457);
or U1963 (N_1963,In_379,In_1883);
xor U1964 (N_1964,In_2462,In_324);
and U1965 (N_1965,In_1180,In_1647);
nor U1966 (N_1966,In_1331,In_2410);
nor U1967 (N_1967,In_483,In_1455);
nand U1968 (N_1968,In_1352,In_2133);
and U1969 (N_1969,In_67,In_879);
and U1970 (N_1970,In_1818,In_691);
xnor U1971 (N_1971,In_2381,In_1226);
and U1972 (N_1972,In_1610,In_31);
or U1973 (N_1973,In_1660,In_237);
nor U1974 (N_1974,In_234,In_285);
nand U1975 (N_1975,In_2199,In_41);
xor U1976 (N_1976,In_1318,In_257);
or U1977 (N_1977,In_550,In_1807);
and U1978 (N_1978,In_517,In_2203);
nor U1979 (N_1979,In_969,In_2320);
or U1980 (N_1980,In_1845,In_1187);
nor U1981 (N_1981,In_2179,In_1988);
nor U1982 (N_1982,In_634,In_2408);
nand U1983 (N_1983,In_932,In_1004);
nand U1984 (N_1984,In_1420,In_51);
or U1985 (N_1985,In_411,In_1301);
and U1986 (N_1986,In_725,In_357);
nand U1987 (N_1987,In_914,In_897);
nand U1988 (N_1988,In_1414,In_817);
nand U1989 (N_1989,In_1989,In_2130);
or U1990 (N_1990,In_1341,In_306);
or U1991 (N_1991,In_1055,In_2039);
xor U1992 (N_1992,In_104,In_1656);
nor U1993 (N_1993,In_1086,In_328);
xor U1994 (N_1994,In_454,In_1685);
nand U1995 (N_1995,In_446,In_1302);
nand U1996 (N_1996,In_1723,In_2320);
nand U1997 (N_1997,In_1498,In_1804);
or U1998 (N_1998,In_202,In_1722);
and U1999 (N_1999,In_1060,In_1015);
and U2000 (N_2000,In_1054,In_1513);
or U2001 (N_2001,In_1821,In_362);
xor U2002 (N_2002,In_307,In_1583);
xnor U2003 (N_2003,In_1261,In_592);
nand U2004 (N_2004,In_1879,In_640);
nor U2005 (N_2005,In_380,In_1189);
xor U2006 (N_2006,In_2146,In_440);
xor U2007 (N_2007,In_2088,In_1453);
or U2008 (N_2008,In_803,In_2476);
nand U2009 (N_2009,In_960,In_1218);
nor U2010 (N_2010,In_1205,In_1653);
nand U2011 (N_2011,In_1672,In_1577);
xnor U2012 (N_2012,In_1077,In_1419);
and U2013 (N_2013,In_931,In_2021);
nand U2014 (N_2014,In_99,In_746);
and U2015 (N_2015,In_2111,In_1560);
xor U2016 (N_2016,In_391,In_2487);
xnor U2017 (N_2017,In_967,In_317);
xnor U2018 (N_2018,In_1746,In_909);
xor U2019 (N_2019,In_1787,In_66);
nand U2020 (N_2020,In_869,In_1899);
xor U2021 (N_2021,In_2436,In_747);
or U2022 (N_2022,In_960,In_2415);
nor U2023 (N_2023,In_2334,In_1671);
and U2024 (N_2024,In_2221,In_1601);
or U2025 (N_2025,In_2226,In_2068);
xor U2026 (N_2026,In_607,In_1544);
nor U2027 (N_2027,In_2307,In_776);
xnor U2028 (N_2028,In_1014,In_2008);
and U2029 (N_2029,In_1734,In_508);
and U2030 (N_2030,In_1379,In_865);
nor U2031 (N_2031,In_1874,In_162);
and U2032 (N_2032,In_2112,In_799);
or U2033 (N_2033,In_426,In_1648);
nand U2034 (N_2034,In_1390,In_1460);
nand U2035 (N_2035,In_1131,In_1860);
xor U2036 (N_2036,In_1592,In_1853);
and U2037 (N_2037,In_562,In_1288);
nand U2038 (N_2038,In_1277,In_1836);
or U2039 (N_2039,In_1340,In_1237);
and U2040 (N_2040,In_1573,In_1581);
xor U2041 (N_2041,In_2044,In_1794);
and U2042 (N_2042,In_37,In_2210);
xor U2043 (N_2043,In_528,In_1563);
nand U2044 (N_2044,In_48,In_1954);
or U2045 (N_2045,In_2250,In_645);
nor U2046 (N_2046,In_742,In_893);
or U2047 (N_2047,In_222,In_920);
and U2048 (N_2048,In_1854,In_35);
xor U2049 (N_2049,In_2182,In_378);
nand U2050 (N_2050,In_645,In_500);
or U2051 (N_2051,In_1475,In_416);
and U2052 (N_2052,In_249,In_1514);
nand U2053 (N_2053,In_708,In_308);
and U2054 (N_2054,In_396,In_1644);
or U2055 (N_2055,In_1395,In_646);
and U2056 (N_2056,In_1131,In_291);
nor U2057 (N_2057,In_65,In_338);
nor U2058 (N_2058,In_1431,In_699);
nand U2059 (N_2059,In_2254,In_1627);
nand U2060 (N_2060,In_1543,In_1356);
and U2061 (N_2061,In_899,In_707);
or U2062 (N_2062,In_104,In_288);
or U2063 (N_2063,In_412,In_867);
nand U2064 (N_2064,In_117,In_2195);
nand U2065 (N_2065,In_1950,In_78);
nand U2066 (N_2066,In_600,In_1683);
or U2067 (N_2067,In_1733,In_2326);
nand U2068 (N_2068,In_1391,In_201);
nor U2069 (N_2069,In_1898,In_56);
and U2070 (N_2070,In_1225,In_1003);
and U2071 (N_2071,In_2363,In_2164);
and U2072 (N_2072,In_647,In_1978);
or U2073 (N_2073,In_2008,In_1419);
and U2074 (N_2074,In_1415,In_1597);
and U2075 (N_2075,In_2072,In_1705);
and U2076 (N_2076,In_1898,In_2179);
and U2077 (N_2077,In_2264,In_1592);
and U2078 (N_2078,In_1614,In_385);
nand U2079 (N_2079,In_2360,In_1821);
and U2080 (N_2080,In_1690,In_999);
and U2081 (N_2081,In_173,In_1785);
nor U2082 (N_2082,In_551,In_329);
nor U2083 (N_2083,In_1893,In_130);
nor U2084 (N_2084,In_1816,In_457);
nand U2085 (N_2085,In_240,In_1451);
or U2086 (N_2086,In_2007,In_133);
nor U2087 (N_2087,In_2373,In_306);
xor U2088 (N_2088,In_1976,In_1170);
nand U2089 (N_2089,In_780,In_1328);
and U2090 (N_2090,In_1286,In_585);
xnor U2091 (N_2091,In_288,In_351);
xnor U2092 (N_2092,In_1173,In_1791);
or U2093 (N_2093,In_1969,In_2018);
nor U2094 (N_2094,In_114,In_1852);
and U2095 (N_2095,In_1419,In_1675);
and U2096 (N_2096,In_85,In_1816);
nor U2097 (N_2097,In_781,In_1183);
xnor U2098 (N_2098,In_627,In_1108);
and U2099 (N_2099,In_295,In_746);
and U2100 (N_2100,In_836,In_2147);
xor U2101 (N_2101,In_1134,In_2350);
nand U2102 (N_2102,In_1951,In_1298);
and U2103 (N_2103,In_1198,In_2218);
xnor U2104 (N_2104,In_2004,In_2413);
nand U2105 (N_2105,In_1728,In_940);
nor U2106 (N_2106,In_2032,In_325);
nor U2107 (N_2107,In_141,In_1894);
nor U2108 (N_2108,In_1010,In_563);
nand U2109 (N_2109,In_1919,In_1836);
xor U2110 (N_2110,In_1195,In_339);
nand U2111 (N_2111,In_1190,In_99);
nand U2112 (N_2112,In_1883,In_2276);
xnor U2113 (N_2113,In_1192,In_593);
or U2114 (N_2114,In_1523,In_677);
xor U2115 (N_2115,In_1894,In_1389);
nor U2116 (N_2116,In_303,In_2285);
or U2117 (N_2117,In_1886,In_721);
or U2118 (N_2118,In_1058,In_756);
and U2119 (N_2119,In_1759,In_635);
and U2120 (N_2120,In_2467,In_1293);
nand U2121 (N_2121,In_2245,In_2353);
and U2122 (N_2122,In_2191,In_2373);
or U2123 (N_2123,In_656,In_439);
nand U2124 (N_2124,In_1490,In_885);
xnor U2125 (N_2125,In_1955,In_2010);
xor U2126 (N_2126,In_1508,In_1901);
or U2127 (N_2127,In_2353,In_1459);
or U2128 (N_2128,In_394,In_1799);
or U2129 (N_2129,In_1225,In_1285);
and U2130 (N_2130,In_2364,In_711);
xnor U2131 (N_2131,In_1138,In_779);
nor U2132 (N_2132,In_582,In_589);
and U2133 (N_2133,In_1409,In_1774);
and U2134 (N_2134,In_1374,In_183);
nor U2135 (N_2135,In_1358,In_1737);
nand U2136 (N_2136,In_2330,In_633);
nand U2137 (N_2137,In_2309,In_1603);
nand U2138 (N_2138,In_2100,In_229);
and U2139 (N_2139,In_65,In_2412);
and U2140 (N_2140,In_575,In_969);
nor U2141 (N_2141,In_1420,In_963);
nor U2142 (N_2142,In_2083,In_1421);
nor U2143 (N_2143,In_582,In_381);
nand U2144 (N_2144,In_2304,In_1746);
xor U2145 (N_2145,In_788,In_1973);
nand U2146 (N_2146,In_807,In_2191);
and U2147 (N_2147,In_828,In_1339);
xnor U2148 (N_2148,In_2479,In_1229);
or U2149 (N_2149,In_93,In_1657);
nand U2150 (N_2150,In_469,In_764);
nor U2151 (N_2151,In_1182,In_760);
xor U2152 (N_2152,In_953,In_2247);
xnor U2153 (N_2153,In_1451,In_838);
xor U2154 (N_2154,In_509,In_547);
nand U2155 (N_2155,In_1953,In_2348);
and U2156 (N_2156,In_1078,In_757);
xor U2157 (N_2157,In_1320,In_2136);
xnor U2158 (N_2158,In_383,In_692);
nand U2159 (N_2159,In_258,In_756);
and U2160 (N_2160,In_432,In_561);
or U2161 (N_2161,In_1246,In_715);
nor U2162 (N_2162,In_1902,In_1343);
xor U2163 (N_2163,In_1837,In_288);
nand U2164 (N_2164,In_640,In_707);
nand U2165 (N_2165,In_2028,In_1841);
nand U2166 (N_2166,In_158,In_2201);
xnor U2167 (N_2167,In_445,In_1003);
nor U2168 (N_2168,In_883,In_990);
nor U2169 (N_2169,In_2118,In_644);
and U2170 (N_2170,In_1593,In_748);
or U2171 (N_2171,In_714,In_1944);
and U2172 (N_2172,In_1609,In_962);
or U2173 (N_2173,In_1042,In_200);
nor U2174 (N_2174,In_2352,In_2354);
nor U2175 (N_2175,In_1491,In_376);
or U2176 (N_2176,In_239,In_318);
and U2177 (N_2177,In_44,In_1698);
xor U2178 (N_2178,In_1614,In_1295);
or U2179 (N_2179,In_1156,In_1299);
nor U2180 (N_2180,In_2236,In_1911);
nor U2181 (N_2181,In_1403,In_2324);
nand U2182 (N_2182,In_2221,In_701);
xor U2183 (N_2183,In_1565,In_1815);
nor U2184 (N_2184,In_864,In_1328);
xnor U2185 (N_2185,In_2413,In_44);
nor U2186 (N_2186,In_1067,In_385);
xnor U2187 (N_2187,In_259,In_703);
nor U2188 (N_2188,In_1804,In_1511);
nand U2189 (N_2189,In_2060,In_1520);
or U2190 (N_2190,In_1736,In_1809);
xnor U2191 (N_2191,In_2105,In_1569);
xnor U2192 (N_2192,In_407,In_184);
xnor U2193 (N_2193,In_1300,In_591);
or U2194 (N_2194,In_757,In_1600);
xor U2195 (N_2195,In_1850,In_824);
or U2196 (N_2196,In_1042,In_1524);
or U2197 (N_2197,In_1090,In_795);
and U2198 (N_2198,In_841,In_25);
nor U2199 (N_2199,In_230,In_2224);
and U2200 (N_2200,In_223,In_1979);
nor U2201 (N_2201,In_2493,In_173);
nor U2202 (N_2202,In_641,In_1367);
nor U2203 (N_2203,In_2486,In_2255);
nand U2204 (N_2204,In_377,In_1798);
nor U2205 (N_2205,In_936,In_2014);
and U2206 (N_2206,In_1991,In_314);
xor U2207 (N_2207,In_181,In_1750);
and U2208 (N_2208,In_501,In_336);
xor U2209 (N_2209,In_1293,In_853);
nand U2210 (N_2210,In_185,In_845);
and U2211 (N_2211,In_490,In_1811);
and U2212 (N_2212,In_1159,In_1324);
nand U2213 (N_2213,In_1871,In_205);
and U2214 (N_2214,In_2311,In_1751);
nor U2215 (N_2215,In_2348,In_865);
nor U2216 (N_2216,In_974,In_298);
and U2217 (N_2217,In_1069,In_789);
and U2218 (N_2218,In_1407,In_812);
or U2219 (N_2219,In_1604,In_1679);
nor U2220 (N_2220,In_2385,In_766);
or U2221 (N_2221,In_2375,In_855);
or U2222 (N_2222,In_1692,In_1740);
nor U2223 (N_2223,In_2343,In_1485);
nand U2224 (N_2224,In_2204,In_1073);
nor U2225 (N_2225,In_939,In_49);
nand U2226 (N_2226,In_1461,In_996);
and U2227 (N_2227,In_544,In_1058);
and U2228 (N_2228,In_714,In_431);
nor U2229 (N_2229,In_119,In_189);
and U2230 (N_2230,In_835,In_1776);
nor U2231 (N_2231,In_1259,In_2209);
xor U2232 (N_2232,In_551,In_1709);
nor U2233 (N_2233,In_809,In_2024);
nand U2234 (N_2234,In_784,In_244);
and U2235 (N_2235,In_789,In_1501);
nor U2236 (N_2236,In_2398,In_88);
nor U2237 (N_2237,In_1436,In_1005);
nand U2238 (N_2238,In_1527,In_1666);
or U2239 (N_2239,In_1844,In_2415);
or U2240 (N_2240,In_1912,In_2083);
and U2241 (N_2241,In_1372,In_79);
or U2242 (N_2242,In_2405,In_2223);
and U2243 (N_2243,In_2028,In_1549);
and U2244 (N_2244,In_1857,In_2180);
xnor U2245 (N_2245,In_1535,In_1938);
xor U2246 (N_2246,In_1550,In_439);
nand U2247 (N_2247,In_938,In_2148);
nor U2248 (N_2248,In_2434,In_758);
xnor U2249 (N_2249,In_500,In_1220);
or U2250 (N_2250,In_739,In_1740);
xnor U2251 (N_2251,In_1383,In_1166);
nor U2252 (N_2252,In_392,In_1698);
or U2253 (N_2253,In_150,In_1002);
or U2254 (N_2254,In_2427,In_698);
xor U2255 (N_2255,In_1305,In_2249);
or U2256 (N_2256,In_1443,In_33);
and U2257 (N_2257,In_2246,In_1365);
xnor U2258 (N_2258,In_387,In_175);
or U2259 (N_2259,In_831,In_1510);
and U2260 (N_2260,In_1104,In_761);
and U2261 (N_2261,In_645,In_808);
xor U2262 (N_2262,In_538,In_150);
or U2263 (N_2263,In_559,In_1634);
xnor U2264 (N_2264,In_1616,In_1953);
nand U2265 (N_2265,In_1267,In_1217);
nand U2266 (N_2266,In_488,In_1798);
nor U2267 (N_2267,In_494,In_130);
nand U2268 (N_2268,In_2388,In_1009);
and U2269 (N_2269,In_1432,In_168);
and U2270 (N_2270,In_2301,In_1892);
nand U2271 (N_2271,In_133,In_1683);
nor U2272 (N_2272,In_2156,In_1796);
nor U2273 (N_2273,In_1185,In_1610);
xor U2274 (N_2274,In_1151,In_2378);
nand U2275 (N_2275,In_1185,In_295);
or U2276 (N_2276,In_715,In_2264);
nand U2277 (N_2277,In_1607,In_2078);
nand U2278 (N_2278,In_2135,In_230);
xor U2279 (N_2279,In_159,In_537);
nor U2280 (N_2280,In_1811,In_518);
nor U2281 (N_2281,In_280,In_2444);
nor U2282 (N_2282,In_30,In_328);
or U2283 (N_2283,In_701,In_125);
nor U2284 (N_2284,In_396,In_7);
xor U2285 (N_2285,In_128,In_916);
nor U2286 (N_2286,In_987,In_998);
or U2287 (N_2287,In_2167,In_840);
xor U2288 (N_2288,In_686,In_1938);
nand U2289 (N_2289,In_529,In_408);
nand U2290 (N_2290,In_1102,In_368);
xor U2291 (N_2291,In_1037,In_2469);
nand U2292 (N_2292,In_1002,In_428);
xor U2293 (N_2293,In_141,In_307);
nor U2294 (N_2294,In_1312,In_503);
nor U2295 (N_2295,In_2141,In_2259);
nor U2296 (N_2296,In_1553,In_427);
or U2297 (N_2297,In_2279,In_1832);
or U2298 (N_2298,In_2213,In_2002);
xnor U2299 (N_2299,In_1065,In_1847);
and U2300 (N_2300,In_1717,In_1481);
or U2301 (N_2301,In_388,In_1336);
and U2302 (N_2302,In_1846,In_859);
xor U2303 (N_2303,In_797,In_683);
nor U2304 (N_2304,In_1131,In_2463);
nor U2305 (N_2305,In_1330,In_2456);
xnor U2306 (N_2306,In_953,In_545);
nor U2307 (N_2307,In_2379,In_190);
and U2308 (N_2308,In_840,In_495);
and U2309 (N_2309,In_1815,In_1432);
xor U2310 (N_2310,In_84,In_2364);
nor U2311 (N_2311,In_287,In_884);
nor U2312 (N_2312,In_1150,In_207);
and U2313 (N_2313,In_960,In_1460);
or U2314 (N_2314,In_1094,In_1060);
nor U2315 (N_2315,In_762,In_1259);
xor U2316 (N_2316,In_1189,In_694);
nand U2317 (N_2317,In_1236,In_2269);
or U2318 (N_2318,In_1710,In_718);
or U2319 (N_2319,In_896,In_1703);
nor U2320 (N_2320,In_475,In_76);
or U2321 (N_2321,In_28,In_843);
xnor U2322 (N_2322,In_1034,In_2319);
nor U2323 (N_2323,In_1080,In_1146);
xor U2324 (N_2324,In_917,In_937);
or U2325 (N_2325,In_1261,In_704);
or U2326 (N_2326,In_2087,In_1052);
xor U2327 (N_2327,In_809,In_187);
and U2328 (N_2328,In_283,In_1465);
nand U2329 (N_2329,In_1191,In_2031);
or U2330 (N_2330,In_2250,In_997);
nor U2331 (N_2331,In_1827,In_2033);
nand U2332 (N_2332,In_754,In_2356);
nand U2333 (N_2333,In_2129,In_1102);
xnor U2334 (N_2334,In_1858,In_582);
or U2335 (N_2335,In_976,In_839);
and U2336 (N_2336,In_349,In_1586);
nor U2337 (N_2337,In_326,In_2356);
nand U2338 (N_2338,In_783,In_1893);
xnor U2339 (N_2339,In_1933,In_1220);
or U2340 (N_2340,In_1271,In_1392);
xnor U2341 (N_2341,In_154,In_2021);
xor U2342 (N_2342,In_1341,In_1963);
and U2343 (N_2343,In_1984,In_464);
xnor U2344 (N_2344,In_1010,In_1238);
and U2345 (N_2345,In_1905,In_2235);
nand U2346 (N_2346,In_1192,In_1255);
nor U2347 (N_2347,In_2459,In_832);
or U2348 (N_2348,In_858,In_715);
or U2349 (N_2349,In_1533,In_1712);
nor U2350 (N_2350,In_1252,In_131);
nor U2351 (N_2351,In_1306,In_464);
and U2352 (N_2352,In_1629,In_219);
nor U2353 (N_2353,In_289,In_1738);
or U2354 (N_2354,In_1015,In_2441);
nand U2355 (N_2355,In_1544,In_2403);
and U2356 (N_2356,In_1549,In_1544);
or U2357 (N_2357,In_276,In_1915);
and U2358 (N_2358,In_1336,In_198);
nand U2359 (N_2359,In_2032,In_1225);
or U2360 (N_2360,In_1546,In_1745);
nand U2361 (N_2361,In_1587,In_250);
nor U2362 (N_2362,In_583,In_2391);
nand U2363 (N_2363,In_80,In_1298);
nor U2364 (N_2364,In_84,In_60);
xor U2365 (N_2365,In_925,In_1164);
nor U2366 (N_2366,In_670,In_1905);
xnor U2367 (N_2367,In_1899,In_1808);
or U2368 (N_2368,In_1124,In_2011);
or U2369 (N_2369,In_329,In_1749);
xor U2370 (N_2370,In_1673,In_443);
and U2371 (N_2371,In_9,In_634);
and U2372 (N_2372,In_197,In_933);
and U2373 (N_2373,In_737,In_444);
nor U2374 (N_2374,In_2035,In_1721);
nand U2375 (N_2375,In_1151,In_148);
or U2376 (N_2376,In_1431,In_784);
nor U2377 (N_2377,In_1635,In_1569);
and U2378 (N_2378,In_598,In_754);
or U2379 (N_2379,In_294,In_1570);
nor U2380 (N_2380,In_7,In_30);
nand U2381 (N_2381,In_2024,In_1263);
xnor U2382 (N_2382,In_340,In_1882);
nand U2383 (N_2383,In_2229,In_2196);
nor U2384 (N_2384,In_2167,In_869);
nor U2385 (N_2385,In_1082,In_402);
nor U2386 (N_2386,In_2199,In_1936);
nand U2387 (N_2387,In_2042,In_2399);
nor U2388 (N_2388,In_1857,In_112);
and U2389 (N_2389,In_1582,In_1767);
xor U2390 (N_2390,In_467,In_1049);
xor U2391 (N_2391,In_1187,In_1932);
and U2392 (N_2392,In_607,In_1177);
and U2393 (N_2393,In_98,In_1260);
nand U2394 (N_2394,In_419,In_1896);
or U2395 (N_2395,In_323,In_1118);
and U2396 (N_2396,In_1074,In_709);
and U2397 (N_2397,In_1443,In_2484);
and U2398 (N_2398,In_1486,In_2149);
nor U2399 (N_2399,In_1498,In_877);
nand U2400 (N_2400,In_1577,In_256);
and U2401 (N_2401,In_1134,In_2031);
or U2402 (N_2402,In_1346,In_835);
nand U2403 (N_2403,In_340,In_650);
or U2404 (N_2404,In_1496,In_2194);
or U2405 (N_2405,In_1757,In_1837);
or U2406 (N_2406,In_282,In_1300);
nor U2407 (N_2407,In_2257,In_1320);
or U2408 (N_2408,In_665,In_164);
or U2409 (N_2409,In_2130,In_610);
xor U2410 (N_2410,In_2294,In_775);
and U2411 (N_2411,In_1274,In_201);
nand U2412 (N_2412,In_1637,In_1184);
xor U2413 (N_2413,In_1833,In_714);
xor U2414 (N_2414,In_2005,In_2431);
and U2415 (N_2415,In_2437,In_1300);
xnor U2416 (N_2416,In_1262,In_1602);
or U2417 (N_2417,In_2277,In_1559);
nor U2418 (N_2418,In_862,In_523);
and U2419 (N_2419,In_720,In_2427);
nor U2420 (N_2420,In_655,In_1028);
nand U2421 (N_2421,In_1963,In_500);
nor U2422 (N_2422,In_759,In_184);
nor U2423 (N_2423,In_2426,In_357);
nand U2424 (N_2424,In_1346,In_1135);
and U2425 (N_2425,In_1135,In_1479);
xor U2426 (N_2426,In_693,In_1175);
and U2427 (N_2427,In_424,In_1596);
or U2428 (N_2428,In_1085,In_2245);
nand U2429 (N_2429,In_940,In_1937);
xnor U2430 (N_2430,In_1920,In_339);
xor U2431 (N_2431,In_176,In_174);
xor U2432 (N_2432,In_1351,In_1473);
nand U2433 (N_2433,In_316,In_834);
nor U2434 (N_2434,In_592,In_1168);
nand U2435 (N_2435,In_2438,In_939);
nand U2436 (N_2436,In_525,In_2011);
or U2437 (N_2437,In_2074,In_155);
or U2438 (N_2438,In_523,In_1202);
nor U2439 (N_2439,In_860,In_2341);
nor U2440 (N_2440,In_2153,In_212);
nor U2441 (N_2441,In_2185,In_956);
xor U2442 (N_2442,In_419,In_1207);
nand U2443 (N_2443,In_1648,In_2323);
or U2444 (N_2444,In_1437,In_1038);
and U2445 (N_2445,In_1543,In_2081);
nand U2446 (N_2446,In_1288,In_799);
xor U2447 (N_2447,In_589,In_566);
nor U2448 (N_2448,In_755,In_2219);
or U2449 (N_2449,In_1954,In_1338);
xnor U2450 (N_2450,In_1047,In_2232);
or U2451 (N_2451,In_1668,In_1713);
or U2452 (N_2452,In_852,In_753);
xor U2453 (N_2453,In_360,In_1594);
nand U2454 (N_2454,In_1494,In_998);
xnor U2455 (N_2455,In_2361,In_2047);
or U2456 (N_2456,In_2456,In_2339);
nand U2457 (N_2457,In_1569,In_1024);
nand U2458 (N_2458,In_685,In_2335);
or U2459 (N_2459,In_1732,In_1548);
xor U2460 (N_2460,In_1360,In_2003);
or U2461 (N_2461,In_1230,In_772);
and U2462 (N_2462,In_2392,In_1817);
nand U2463 (N_2463,In_2278,In_1548);
nor U2464 (N_2464,In_845,In_527);
nor U2465 (N_2465,In_2438,In_1736);
nor U2466 (N_2466,In_1898,In_909);
nand U2467 (N_2467,In_1078,In_813);
or U2468 (N_2468,In_168,In_300);
or U2469 (N_2469,In_2312,In_2467);
xnor U2470 (N_2470,In_390,In_988);
and U2471 (N_2471,In_2488,In_1667);
or U2472 (N_2472,In_97,In_1614);
nand U2473 (N_2473,In_736,In_1314);
nor U2474 (N_2474,In_54,In_469);
xnor U2475 (N_2475,In_1740,In_9);
nand U2476 (N_2476,In_1651,In_57);
nand U2477 (N_2477,In_368,In_605);
nand U2478 (N_2478,In_121,In_316);
xor U2479 (N_2479,In_1162,In_1479);
nand U2480 (N_2480,In_1224,In_401);
and U2481 (N_2481,In_1919,In_787);
or U2482 (N_2482,In_1448,In_1647);
xor U2483 (N_2483,In_276,In_915);
and U2484 (N_2484,In_1835,In_1127);
and U2485 (N_2485,In_400,In_2281);
or U2486 (N_2486,In_1035,In_1528);
or U2487 (N_2487,In_1552,In_630);
nand U2488 (N_2488,In_1468,In_602);
or U2489 (N_2489,In_1661,In_1504);
nor U2490 (N_2490,In_865,In_1351);
nor U2491 (N_2491,In_2174,In_1204);
or U2492 (N_2492,In_2391,In_1637);
or U2493 (N_2493,In_2278,In_1255);
and U2494 (N_2494,In_575,In_1905);
nor U2495 (N_2495,In_625,In_888);
nor U2496 (N_2496,In_165,In_744);
nand U2497 (N_2497,In_1981,In_966);
nor U2498 (N_2498,In_806,In_2294);
nor U2499 (N_2499,In_550,In_1615);
and U2500 (N_2500,In_2078,In_999);
nand U2501 (N_2501,In_1044,In_990);
and U2502 (N_2502,In_1525,In_2391);
nand U2503 (N_2503,In_889,In_1828);
xor U2504 (N_2504,In_1855,In_1371);
nor U2505 (N_2505,In_2278,In_2056);
and U2506 (N_2506,In_2244,In_1562);
and U2507 (N_2507,In_1200,In_272);
nand U2508 (N_2508,In_1580,In_602);
or U2509 (N_2509,In_1056,In_714);
nor U2510 (N_2510,In_2371,In_929);
xor U2511 (N_2511,In_1319,In_631);
and U2512 (N_2512,In_51,In_577);
and U2513 (N_2513,In_1300,In_654);
xor U2514 (N_2514,In_487,In_853);
xnor U2515 (N_2515,In_1919,In_1362);
and U2516 (N_2516,In_261,In_1361);
nor U2517 (N_2517,In_2223,In_396);
and U2518 (N_2518,In_1196,In_1676);
or U2519 (N_2519,In_810,In_2066);
and U2520 (N_2520,In_1321,In_1400);
xnor U2521 (N_2521,In_1232,In_609);
nand U2522 (N_2522,In_886,In_1658);
nand U2523 (N_2523,In_1180,In_1684);
nor U2524 (N_2524,In_510,In_262);
nor U2525 (N_2525,In_2057,In_379);
nor U2526 (N_2526,In_1313,In_1885);
or U2527 (N_2527,In_2369,In_1979);
nor U2528 (N_2528,In_1581,In_397);
and U2529 (N_2529,In_43,In_2173);
nand U2530 (N_2530,In_657,In_2310);
or U2531 (N_2531,In_1479,In_1898);
nor U2532 (N_2532,In_850,In_1387);
nor U2533 (N_2533,In_1953,In_1169);
nand U2534 (N_2534,In_1789,In_702);
nand U2535 (N_2535,In_296,In_1669);
xnor U2536 (N_2536,In_1680,In_2404);
or U2537 (N_2537,In_1718,In_210);
or U2538 (N_2538,In_698,In_1122);
or U2539 (N_2539,In_374,In_1635);
xnor U2540 (N_2540,In_449,In_1728);
or U2541 (N_2541,In_413,In_0);
nand U2542 (N_2542,In_725,In_801);
and U2543 (N_2543,In_2421,In_1559);
or U2544 (N_2544,In_165,In_1071);
xnor U2545 (N_2545,In_1435,In_1940);
nor U2546 (N_2546,In_324,In_255);
and U2547 (N_2547,In_348,In_405);
or U2548 (N_2548,In_1424,In_50);
or U2549 (N_2549,In_1461,In_192);
and U2550 (N_2550,In_442,In_129);
xnor U2551 (N_2551,In_1203,In_144);
or U2552 (N_2552,In_248,In_267);
nand U2553 (N_2553,In_416,In_1326);
nand U2554 (N_2554,In_195,In_1107);
nand U2555 (N_2555,In_1597,In_104);
nand U2556 (N_2556,In_772,In_483);
nor U2557 (N_2557,In_2251,In_879);
xor U2558 (N_2558,In_1377,In_695);
nand U2559 (N_2559,In_1219,In_521);
and U2560 (N_2560,In_397,In_2201);
or U2561 (N_2561,In_2275,In_147);
and U2562 (N_2562,In_2317,In_978);
or U2563 (N_2563,In_261,In_975);
or U2564 (N_2564,In_1981,In_1750);
nand U2565 (N_2565,In_35,In_1094);
nand U2566 (N_2566,In_664,In_947);
and U2567 (N_2567,In_2432,In_1405);
and U2568 (N_2568,In_1333,In_95);
or U2569 (N_2569,In_205,In_554);
nor U2570 (N_2570,In_618,In_753);
or U2571 (N_2571,In_2163,In_1355);
or U2572 (N_2572,In_2333,In_2346);
nand U2573 (N_2573,In_469,In_1285);
nand U2574 (N_2574,In_1235,In_955);
nor U2575 (N_2575,In_515,In_1400);
or U2576 (N_2576,In_792,In_812);
and U2577 (N_2577,In_2113,In_990);
and U2578 (N_2578,In_1255,In_310);
or U2579 (N_2579,In_238,In_654);
nor U2580 (N_2580,In_273,In_1137);
nor U2581 (N_2581,In_2003,In_515);
nor U2582 (N_2582,In_845,In_1747);
or U2583 (N_2583,In_1792,In_697);
nor U2584 (N_2584,In_227,In_713);
nand U2585 (N_2585,In_1693,In_384);
and U2586 (N_2586,In_2035,In_1865);
xor U2587 (N_2587,In_277,In_1029);
xnor U2588 (N_2588,In_687,In_1042);
or U2589 (N_2589,In_2146,In_2349);
nor U2590 (N_2590,In_603,In_817);
and U2591 (N_2591,In_184,In_1615);
or U2592 (N_2592,In_279,In_142);
or U2593 (N_2593,In_1109,In_228);
or U2594 (N_2594,In_1614,In_886);
nor U2595 (N_2595,In_1281,In_1118);
nor U2596 (N_2596,In_209,In_2260);
and U2597 (N_2597,In_674,In_1019);
and U2598 (N_2598,In_2250,In_260);
nand U2599 (N_2599,In_2253,In_86);
xor U2600 (N_2600,In_1975,In_396);
nand U2601 (N_2601,In_1163,In_2292);
nand U2602 (N_2602,In_615,In_666);
and U2603 (N_2603,In_2213,In_299);
or U2604 (N_2604,In_2097,In_2224);
or U2605 (N_2605,In_1369,In_2361);
and U2606 (N_2606,In_1668,In_2267);
or U2607 (N_2607,In_2066,In_1529);
or U2608 (N_2608,In_2325,In_321);
nand U2609 (N_2609,In_611,In_2327);
nor U2610 (N_2610,In_2268,In_54);
or U2611 (N_2611,In_1915,In_1771);
and U2612 (N_2612,In_1973,In_2325);
xnor U2613 (N_2613,In_173,In_33);
xnor U2614 (N_2614,In_2371,In_1948);
nand U2615 (N_2615,In_548,In_1561);
nor U2616 (N_2616,In_678,In_1849);
xor U2617 (N_2617,In_1971,In_818);
xnor U2618 (N_2618,In_555,In_1137);
or U2619 (N_2619,In_77,In_1598);
or U2620 (N_2620,In_1682,In_1061);
xnor U2621 (N_2621,In_10,In_2214);
nand U2622 (N_2622,In_140,In_835);
nand U2623 (N_2623,In_1971,In_371);
xor U2624 (N_2624,In_2487,In_798);
nand U2625 (N_2625,In_559,In_1700);
nor U2626 (N_2626,In_1585,In_500);
xnor U2627 (N_2627,In_1520,In_2469);
xor U2628 (N_2628,In_83,In_2029);
nand U2629 (N_2629,In_170,In_726);
nand U2630 (N_2630,In_1669,In_2446);
or U2631 (N_2631,In_1516,In_660);
nand U2632 (N_2632,In_1242,In_1866);
and U2633 (N_2633,In_2093,In_1533);
or U2634 (N_2634,In_1738,In_1755);
or U2635 (N_2635,In_762,In_106);
and U2636 (N_2636,In_439,In_50);
nor U2637 (N_2637,In_2135,In_536);
nor U2638 (N_2638,In_748,In_860);
xnor U2639 (N_2639,In_1501,In_2388);
or U2640 (N_2640,In_2078,In_862);
xor U2641 (N_2641,In_2026,In_364);
nand U2642 (N_2642,In_399,In_560);
xor U2643 (N_2643,In_12,In_2477);
xor U2644 (N_2644,In_1879,In_1463);
nand U2645 (N_2645,In_467,In_224);
and U2646 (N_2646,In_1144,In_1095);
or U2647 (N_2647,In_62,In_2317);
nor U2648 (N_2648,In_1733,In_1322);
nand U2649 (N_2649,In_2317,In_1821);
nand U2650 (N_2650,In_724,In_726);
nor U2651 (N_2651,In_2193,In_1139);
and U2652 (N_2652,In_1521,In_2299);
and U2653 (N_2653,In_2378,In_6);
nor U2654 (N_2654,In_1718,In_1505);
nor U2655 (N_2655,In_2050,In_2004);
nor U2656 (N_2656,In_1086,In_1684);
nor U2657 (N_2657,In_1970,In_2150);
or U2658 (N_2658,In_651,In_1808);
nand U2659 (N_2659,In_1002,In_1893);
and U2660 (N_2660,In_1040,In_896);
nand U2661 (N_2661,In_1378,In_301);
or U2662 (N_2662,In_392,In_776);
nor U2663 (N_2663,In_412,In_672);
or U2664 (N_2664,In_518,In_2483);
xor U2665 (N_2665,In_2424,In_234);
and U2666 (N_2666,In_257,In_2217);
or U2667 (N_2667,In_7,In_1372);
nor U2668 (N_2668,In_89,In_152);
nand U2669 (N_2669,In_1777,In_2475);
nor U2670 (N_2670,In_1199,In_279);
nand U2671 (N_2671,In_847,In_1276);
nor U2672 (N_2672,In_1271,In_655);
nand U2673 (N_2673,In_50,In_1686);
or U2674 (N_2674,In_2266,In_1632);
nor U2675 (N_2675,In_1713,In_521);
xor U2676 (N_2676,In_1671,In_1888);
xnor U2677 (N_2677,In_389,In_772);
xor U2678 (N_2678,In_2071,In_2413);
and U2679 (N_2679,In_1368,In_59);
nand U2680 (N_2680,In_1707,In_2498);
xor U2681 (N_2681,In_316,In_63);
xnor U2682 (N_2682,In_681,In_1234);
or U2683 (N_2683,In_1390,In_1755);
or U2684 (N_2684,In_1741,In_228);
xnor U2685 (N_2685,In_1719,In_1547);
nor U2686 (N_2686,In_1588,In_1070);
and U2687 (N_2687,In_2133,In_1035);
or U2688 (N_2688,In_2067,In_258);
xnor U2689 (N_2689,In_103,In_2361);
nor U2690 (N_2690,In_1272,In_2264);
nand U2691 (N_2691,In_2025,In_508);
and U2692 (N_2692,In_1660,In_1450);
nor U2693 (N_2693,In_636,In_1507);
xnor U2694 (N_2694,In_1656,In_1526);
xnor U2695 (N_2695,In_168,In_1356);
or U2696 (N_2696,In_1563,In_1693);
xnor U2697 (N_2697,In_1115,In_2012);
nand U2698 (N_2698,In_1460,In_670);
nand U2699 (N_2699,In_2327,In_1140);
or U2700 (N_2700,In_502,In_640);
nor U2701 (N_2701,In_620,In_987);
nand U2702 (N_2702,In_150,In_1847);
or U2703 (N_2703,In_1887,In_298);
nand U2704 (N_2704,In_951,In_1601);
or U2705 (N_2705,In_1799,In_117);
and U2706 (N_2706,In_2087,In_171);
or U2707 (N_2707,In_1118,In_1001);
xnor U2708 (N_2708,In_2182,In_2120);
nand U2709 (N_2709,In_2260,In_1296);
xor U2710 (N_2710,In_673,In_2307);
nand U2711 (N_2711,In_107,In_494);
or U2712 (N_2712,In_2290,In_2234);
or U2713 (N_2713,In_160,In_362);
or U2714 (N_2714,In_2034,In_250);
nor U2715 (N_2715,In_412,In_1008);
nand U2716 (N_2716,In_1771,In_1739);
nor U2717 (N_2717,In_683,In_1345);
nand U2718 (N_2718,In_2118,In_535);
xor U2719 (N_2719,In_36,In_1033);
or U2720 (N_2720,In_1003,In_325);
nand U2721 (N_2721,In_44,In_2097);
nand U2722 (N_2722,In_776,In_1483);
nand U2723 (N_2723,In_1942,In_551);
nor U2724 (N_2724,In_2085,In_1391);
xnor U2725 (N_2725,In_678,In_872);
xnor U2726 (N_2726,In_1648,In_1006);
nand U2727 (N_2727,In_1483,In_2040);
nor U2728 (N_2728,In_1167,In_615);
nand U2729 (N_2729,In_2053,In_1457);
nand U2730 (N_2730,In_218,In_2446);
and U2731 (N_2731,In_651,In_1730);
xnor U2732 (N_2732,In_2306,In_453);
nor U2733 (N_2733,In_2434,In_1063);
nor U2734 (N_2734,In_1631,In_1482);
nor U2735 (N_2735,In_748,In_1366);
or U2736 (N_2736,In_2246,In_28);
or U2737 (N_2737,In_681,In_592);
nor U2738 (N_2738,In_1971,In_5);
and U2739 (N_2739,In_312,In_2462);
or U2740 (N_2740,In_2223,In_196);
nand U2741 (N_2741,In_163,In_1303);
nand U2742 (N_2742,In_1092,In_13);
or U2743 (N_2743,In_177,In_1105);
and U2744 (N_2744,In_1337,In_324);
and U2745 (N_2745,In_2177,In_2031);
nor U2746 (N_2746,In_488,In_2256);
nor U2747 (N_2747,In_901,In_78);
and U2748 (N_2748,In_957,In_2006);
xor U2749 (N_2749,In_1293,In_1522);
xnor U2750 (N_2750,In_427,In_747);
nand U2751 (N_2751,In_24,In_1692);
and U2752 (N_2752,In_643,In_1189);
and U2753 (N_2753,In_34,In_932);
and U2754 (N_2754,In_19,In_1691);
nor U2755 (N_2755,In_904,In_273);
or U2756 (N_2756,In_978,In_202);
nor U2757 (N_2757,In_997,In_1380);
xnor U2758 (N_2758,In_537,In_1935);
or U2759 (N_2759,In_523,In_118);
nand U2760 (N_2760,In_2278,In_1737);
xnor U2761 (N_2761,In_2275,In_2443);
nand U2762 (N_2762,In_1185,In_917);
or U2763 (N_2763,In_2177,In_1759);
xnor U2764 (N_2764,In_1339,In_1888);
or U2765 (N_2765,In_568,In_1655);
nor U2766 (N_2766,In_1662,In_1251);
nand U2767 (N_2767,In_486,In_421);
xnor U2768 (N_2768,In_1144,In_221);
nand U2769 (N_2769,In_1479,In_2136);
nor U2770 (N_2770,In_1932,In_1854);
and U2771 (N_2771,In_1505,In_18);
nor U2772 (N_2772,In_2164,In_1942);
or U2773 (N_2773,In_1887,In_990);
and U2774 (N_2774,In_1449,In_966);
or U2775 (N_2775,In_560,In_1165);
and U2776 (N_2776,In_1083,In_589);
and U2777 (N_2777,In_2060,In_1294);
or U2778 (N_2778,In_222,In_1307);
nor U2779 (N_2779,In_2172,In_345);
nand U2780 (N_2780,In_2038,In_459);
nand U2781 (N_2781,In_1842,In_97);
nor U2782 (N_2782,In_2185,In_1254);
xnor U2783 (N_2783,In_252,In_1322);
and U2784 (N_2784,In_2291,In_746);
nor U2785 (N_2785,In_2411,In_686);
or U2786 (N_2786,In_982,In_856);
or U2787 (N_2787,In_67,In_2085);
xnor U2788 (N_2788,In_51,In_1344);
and U2789 (N_2789,In_591,In_849);
and U2790 (N_2790,In_1988,In_2306);
xnor U2791 (N_2791,In_1542,In_209);
nor U2792 (N_2792,In_1826,In_1786);
nand U2793 (N_2793,In_509,In_1781);
xnor U2794 (N_2794,In_934,In_2195);
nand U2795 (N_2795,In_571,In_1767);
or U2796 (N_2796,In_796,In_294);
or U2797 (N_2797,In_556,In_1642);
nand U2798 (N_2798,In_2367,In_1846);
and U2799 (N_2799,In_1955,In_778);
and U2800 (N_2800,In_1271,In_992);
nor U2801 (N_2801,In_2030,In_882);
nand U2802 (N_2802,In_986,In_1671);
nor U2803 (N_2803,In_1499,In_675);
or U2804 (N_2804,In_2141,In_1623);
and U2805 (N_2805,In_1624,In_468);
nand U2806 (N_2806,In_435,In_312);
nor U2807 (N_2807,In_2033,In_818);
nand U2808 (N_2808,In_2313,In_480);
and U2809 (N_2809,In_1989,In_1036);
and U2810 (N_2810,In_168,In_1695);
nand U2811 (N_2811,In_2236,In_2077);
xor U2812 (N_2812,In_821,In_61);
nand U2813 (N_2813,In_976,In_263);
nor U2814 (N_2814,In_318,In_1767);
or U2815 (N_2815,In_751,In_406);
nand U2816 (N_2816,In_1314,In_2158);
and U2817 (N_2817,In_1940,In_1168);
xor U2818 (N_2818,In_2460,In_252);
and U2819 (N_2819,In_451,In_224);
nand U2820 (N_2820,In_2320,In_1408);
xnor U2821 (N_2821,In_367,In_1135);
nor U2822 (N_2822,In_845,In_857);
or U2823 (N_2823,In_479,In_1447);
xnor U2824 (N_2824,In_1107,In_1226);
xnor U2825 (N_2825,In_1406,In_528);
or U2826 (N_2826,In_742,In_1786);
nor U2827 (N_2827,In_1614,In_570);
nand U2828 (N_2828,In_166,In_778);
nand U2829 (N_2829,In_1642,In_730);
and U2830 (N_2830,In_1625,In_1551);
or U2831 (N_2831,In_1648,In_367);
nand U2832 (N_2832,In_2301,In_658);
nor U2833 (N_2833,In_496,In_2251);
nor U2834 (N_2834,In_851,In_1355);
nor U2835 (N_2835,In_1827,In_1628);
nor U2836 (N_2836,In_598,In_2472);
nor U2837 (N_2837,In_1911,In_2068);
nor U2838 (N_2838,In_1116,In_378);
and U2839 (N_2839,In_1810,In_1865);
nor U2840 (N_2840,In_2314,In_1748);
or U2841 (N_2841,In_63,In_1766);
and U2842 (N_2842,In_563,In_1285);
or U2843 (N_2843,In_624,In_296);
or U2844 (N_2844,In_812,In_1285);
xor U2845 (N_2845,In_1108,In_963);
xnor U2846 (N_2846,In_789,In_574);
nand U2847 (N_2847,In_1693,In_1609);
nor U2848 (N_2848,In_1190,In_1943);
xor U2849 (N_2849,In_2387,In_1615);
xor U2850 (N_2850,In_1196,In_542);
and U2851 (N_2851,In_354,In_2180);
nand U2852 (N_2852,In_2465,In_1116);
xor U2853 (N_2853,In_500,In_2128);
nand U2854 (N_2854,In_2039,In_649);
nor U2855 (N_2855,In_825,In_431);
xnor U2856 (N_2856,In_813,In_279);
xor U2857 (N_2857,In_577,In_1735);
xnor U2858 (N_2858,In_222,In_1587);
or U2859 (N_2859,In_1117,In_1874);
xnor U2860 (N_2860,In_216,In_2219);
and U2861 (N_2861,In_145,In_1161);
nand U2862 (N_2862,In_934,In_2267);
nand U2863 (N_2863,In_1083,In_881);
and U2864 (N_2864,In_1529,In_1116);
or U2865 (N_2865,In_2347,In_709);
nand U2866 (N_2866,In_1010,In_588);
xnor U2867 (N_2867,In_2033,In_1544);
xor U2868 (N_2868,In_650,In_2);
xnor U2869 (N_2869,In_2304,In_669);
nor U2870 (N_2870,In_611,In_987);
and U2871 (N_2871,In_2417,In_1847);
nand U2872 (N_2872,In_2036,In_812);
nor U2873 (N_2873,In_2317,In_1128);
nand U2874 (N_2874,In_1151,In_1719);
nand U2875 (N_2875,In_1172,In_1490);
or U2876 (N_2876,In_1167,In_2412);
xor U2877 (N_2877,In_2115,In_1687);
or U2878 (N_2878,In_915,In_660);
nor U2879 (N_2879,In_1916,In_797);
and U2880 (N_2880,In_766,In_715);
and U2881 (N_2881,In_611,In_2234);
nand U2882 (N_2882,In_2257,In_2164);
and U2883 (N_2883,In_878,In_1373);
and U2884 (N_2884,In_2010,In_2310);
nor U2885 (N_2885,In_2422,In_821);
nor U2886 (N_2886,In_1313,In_2214);
nor U2887 (N_2887,In_2480,In_2035);
and U2888 (N_2888,In_836,In_725);
and U2889 (N_2889,In_279,In_391);
nand U2890 (N_2890,In_1681,In_2174);
nand U2891 (N_2891,In_964,In_1531);
and U2892 (N_2892,In_2189,In_805);
nand U2893 (N_2893,In_678,In_958);
and U2894 (N_2894,In_1622,In_1879);
nand U2895 (N_2895,In_2332,In_833);
or U2896 (N_2896,In_1069,In_1782);
and U2897 (N_2897,In_924,In_1);
nand U2898 (N_2898,In_1136,In_465);
nor U2899 (N_2899,In_1264,In_2182);
nor U2900 (N_2900,In_266,In_1418);
xnor U2901 (N_2901,In_2004,In_760);
or U2902 (N_2902,In_2100,In_35);
nand U2903 (N_2903,In_1301,In_2028);
or U2904 (N_2904,In_2402,In_1912);
nand U2905 (N_2905,In_881,In_2172);
or U2906 (N_2906,In_2438,In_2115);
xnor U2907 (N_2907,In_643,In_89);
and U2908 (N_2908,In_2213,In_1791);
and U2909 (N_2909,In_936,In_1787);
or U2910 (N_2910,In_2085,In_697);
or U2911 (N_2911,In_621,In_946);
nand U2912 (N_2912,In_2067,In_1782);
and U2913 (N_2913,In_133,In_761);
or U2914 (N_2914,In_48,In_1637);
nor U2915 (N_2915,In_2472,In_1697);
and U2916 (N_2916,In_1947,In_980);
nor U2917 (N_2917,In_152,In_725);
nand U2918 (N_2918,In_314,In_2467);
nor U2919 (N_2919,In_2466,In_330);
nand U2920 (N_2920,In_2141,In_1592);
nand U2921 (N_2921,In_322,In_119);
nand U2922 (N_2922,In_2185,In_2018);
xnor U2923 (N_2923,In_657,In_1928);
or U2924 (N_2924,In_2469,In_1923);
nor U2925 (N_2925,In_1826,In_494);
or U2926 (N_2926,In_1724,In_1665);
nand U2927 (N_2927,In_1046,In_1292);
nand U2928 (N_2928,In_1302,In_1185);
and U2929 (N_2929,In_2079,In_296);
or U2930 (N_2930,In_2129,In_767);
nand U2931 (N_2931,In_1581,In_910);
nor U2932 (N_2932,In_2074,In_1553);
nor U2933 (N_2933,In_450,In_2324);
or U2934 (N_2934,In_672,In_116);
and U2935 (N_2935,In_1760,In_841);
nor U2936 (N_2936,In_2226,In_1358);
xor U2937 (N_2937,In_1559,In_318);
or U2938 (N_2938,In_2284,In_2485);
xnor U2939 (N_2939,In_669,In_2398);
nor U2940 (N_2940,In_1256,In_1913);
or U2941 (N_2941,In_472,In_737);
nand U2942 (N_2942,In_4,In_2309);
and U2943 (N_2943,In_2448,In_372);
and U2944 (N_2944,In_2386,In_327);
and U2945 (N_2945,In_2471,In_1205);
xnor U2946 (N_2946,In_882,In_2115);
nand U2947 (N_2947,In_455,In_1277);
nor U2948 (N_2948,In_280,In_2306);
nor U2949 (N_2949,In_579,In_2385);
or U2950 (N_2950,In_305,In_1266);
nand U2951 (N_2951,In_291,In_2479);
nand U2952 (N_2952,In_2395,In_28);
nor U2953 (N_2953,In_1816,In_2177);
and U2954 (N_2954,In_81,In_660);
and U2955 (N_2955,In_2220,In_276);
nor U2956 (N_2956,In_2089,In_2318);
nor U2957 (N_2957,In_283,In_958);
and U2958 (N_2958,In_1449,In_693);
or U2959 (N_2959,In_1216,In_2128);
nand U2960 (N_2960,In_1100,In_753);
xor U2961 (N_2961,In_1066,In_1186);
nand U2962 (N_2962,In_1313,In_2094);
or U2963 (N_2963,In_1047,In_396);
nor U2964 (N_2964,In_2432,In_1640);
nor U2965 (N_2965,In_1949,In_2175);
nor U2966 (N_2966,In_1985,In_96);
nor U2967 (N_2967,In_1005,In_23);
nand U2968 (N_2968,In_914,In_2069);
nand U2969 (N_2969,In_2404,In_1841);
nand U2970 (N_2970,In_1271,In_435);
and U2971 (N_2971,In_2385,In_2452);
xnor U2972 (N_2972,In_1577,In_1025);
and U2973 (N_2973,In_480,In_2366);
nand U2974 (N_2974,In_1564,In_1019);
nand U2975 (N_2975,In_599,In_80);
or U2976 (N_2976,In_1156,In_637);
nand U2977 (N_2977,In_540,In_1089);
or U2978 (N_2978,In_1465,In_895);
nand U2979 (N_2979,In_2287,In_1576);
xnor U2980 (N_2980,In_805,In_390);
xnor U2981 (N_2981,In_1417,In_2111);
or U2982 (N_2982,In_1613,In_1838);
nand U2983 (N_2983,In_450,In_2343);
xnor U2984 (N_2984,In_1467,In_123);
or U2985 (N_2985,In_1703,In_1283);
and U2986 (N_2986,In_1133,In_1067);
xor U2987 (N_2987,In_1126,In_1925);
or U2988 (N_2988,In_236,In_2210);
or U2989 (N_2989,In_1301,In_2155);
xor U2990 (N_2990,In_2144,In_635);
and U2991 (N_2991,In_1984,In_800);
xor U2992 (N_2992,In_1556,In_2150);
or U2993 (N_2993,In_1932,In_1055);
nand U2994 (N_2994,In_33,In_1268);
or U2995 (N_2995,In_181,In_1932);
and U2996 (N_2996,In_1408,In_2200);
nand U2997 (N_2997,In_353,In_1965);
nand U2998 (N_2998,In_1928,In_1849);
and U2999 (N_2999,In_1926,In_655);
xnor U3000 (N_3000,In_34,In_688);
nand U3001 (N_3001,In_35,In_2079);
or U3002 (N_3002,In_265,In_2324);
nor U3003 (N_3003,In_1397,In_1295);
xor U3004 (N_3004,In_71,In_495);
nand U3005 (N_3005,In_1548,In_522);
nand U3006 (N_3006,In_1276,In_1440);
nor U3007 (N_3007,In_48,In_392);
or U3008 (N_3008,In_611,In_1021);
or U3009 (N_3009,In_470,In_2364);
xor U3010 (N_3010,In_2250,In_165);
nor U3011 (N_3011,In_1905,In_948);
nor U3012 (N_3012,In_2049,In_2261);
or U3013 (N_3013,In_2140,In_2428);
nand U3014 (N_3014,In_848,In_1261);
or U3015 (N_3015,In_1887,In_1435);
nor U3016 (N_3016,In_1222,In_1580);
xor U3017 (N_3017,In_1464,In_230);
nand U3018 (N_3018,In_2172,In_871);
or U3019 (N_3019,In_12,In_593);
nor U3020 (N_3020,In_1916,In_2211);
nand U3021 (N_3021,In_974,In_1924);
nand U3022 (N_3022,In_1006,In_967);
or U3023 (N_3023,In_754,In_2102);
nand U3024 (N_3024,In_1731,In_481);
or U3025 (N_3025,In_342,In_1696);
nor U3026 (N_3026,In_1258,In_688);
or U3027 (N_3027,In_1121,In_1850);
nand U3028 (N_3028,In_1574,In_1280);
nand U3029 (N_3029,In_1238,In_1132);
nand U3030 (N_3030,In_2140,In_2279);
nand U3031 (N_3031,In_1921,In_96);
xor U3032 (N_3032,In_2453,In_1841);
nor U3033 (N_3033,In_851,In_105);
nand U3034 (N_3034,In_666,In_737);
xnor U3035 (N_3035,In_461,In_984);
nor U3036 (N_3036,In_535,In_810);
nand U3037 (N_3037,In_1619,In_390);
nand U3038 (N_3038,In_170,In_237);
or U3039 (N_3039,In_1653,In_2043);
nor U3040 (N_3040,In_727,In_2030);
xor U3041 (N_3041,In_1780,In_59);
and U3042 (N_3042,In_777,In_1294);
nor U3043 (N_3043,In_349,In_633);
xnor U3044 (N_3044,In_2025,In_2078);
xor U3045 (N_3045,In_1896,In_1498);
or U3046 (N_3046,In_2383,In_223);
xor U3047 (N_3047,In_871,In_1043);
xor U3048 (N_3048,In_1971,In_2190);
nor U3049 (N_3049,In_743,In_1662);
and U3050 (N_3050,In_2032,In_2184);
and U3051 (N_3051,In_1117,In_1647);
nor U3052 (N_3052,In_130,In_902);
and U3053 (N_3053,In_41,In_1545);
and U3054 (N_3054,In_2437,In_1454);
nor U3055 (N_3055,In_165,In_2172);
nor U3056 (N_3056,In_1041,In_1925);
and U3057 (N_3057,In_1692,In_2423);
nand U3058 (N_3058,In_517,In_906);
and U3059 (N_3059,In_2264,In_1598);
xnor U3060 (N_3060,In_203,In_1064);
nor U3061 (N_3061,In_1028,In_1933);
xor U3062 (N_3062,In_376,In_2087);
nand U3063 (N_3063,In_1626,In_1084);
and U3064 (N_3064,In_2332,In_2067);
or U3065 (N_3065,In_1546,In_2155);
and U3066 (N_3066,In_1299,In_426);
nand U3067 (N_3067,In_1877,In_411);
and U3068 (N_3068,In_2068,In_500);
or U3069 (N_3069,In_1659,In_1687);
xnor U3070 (N_3070,In_2198,In_834);
nand U3071 (N_3071,In_73,In_15);
and U3072 (N_3072,In_352,In_813);
xnor U3073 (N_3073,In_1828,In_42);
and U3074 (N_3074,In_1309,In_2266);
or U3075 (N_3075,In_1566,In_2308);
or U3076 (N_3076,In_1338,In_2429);
nor U3077 (N_3077,In_2047,In_896);
nand U3078 (N_3078,In_2194,In_308);
nor U3079 (N_3079,In_2245,In_1835);
xnor U3080 (N_3080,In_2351,In_793);
or U3081 (N_3081,In_616,In_330);
and U3082 (N_3082,In_1694,In_549);
or U3083 (N_3083,In_1366,In_1949);
nor U3084 (N_3084,In_891,In_42);
xnor U3085 (N_3085,In_1514,In_99);
or U3086 (N_3086,In_1626,In_1682);
nand U3087 (N_3087,In_761,In_699);
or U3088 (N_3088,In_1094,In_2368);
or U3089 (N_3089,In_1010,In_1998);
or U3090 (N_3090,In_106,In_1803);
or U3091 (N_3091,In_1315,In_586);
xnor U3092 (N_3092,In_1431,In_1010);
nor U3093 (N_3093,In_1823,In_1056);
nand U3094 (N_3094,In_1946,In_2102);
or U3095 (N_3095,In_2329,In_1453);
nor U3096 (N_3096,In_2172,In_652);
and U3097 (N_3097,In_2028,In_957);
or U3098 (N_3098,In_69,In_1086);
or U3099 (N_3099,In_2182,In_1111);
xnor U3100 (N_3100,In_1222,In_440);
nand U3101 (N_3101,In_1352,In_1633);
nand U3102 (N_3102,In_726,In_1378);
or U3103 (N_3103,In_2479,In_1126);
nor U3104 (N_3104,In_321,In_564);
or U3105 (N_3105,In_1705,In_709);
xor U3106 (N_3106,In_2064,In_212);
nand U3107 (N_3107,In_1900,In_1152);
and U3108 (N_3108,In_827,In_1028);
nor U3109 (N_3109,In_2329,In_1475);
and U3110 (N_3110,In_528,In_1485);
nand U3111 (N_3111,In_1462,In_854);
or U3112 (N_3112,In_1728,In_2086);
or U3113 (N_3113,In_1606,In_1139);
and U3114 (N_3114,In_2152,In_2231);
nor U3115 (N_3115,In_1919,In_1514);
and U3116 (N_3116,In_438,In_2441);
or U3117 (N_3117,In_2180,In_1602);
and U3118 (N_3118,In_1830,In_2479);
nand U3119 (N_3119,In_658,In_977);
xnor U3120 (N_3120,In_1333,In_905);
or U3121 (N_3121,In_2360,In_1569);
nor U3122 (N_3122,In_859,In_1089);
xnor U3123 (N_3123,In_2395,In_1617);
xnor U3124 (N_3124,In_2081,In_813);
nand U3125 (N_3125,In_2066,In_1129);
and U3126 (N_3126,In_2080,In_1335);
xnor U3127 (N_3127,In_2485,In_1042);
or U3128 (N_3128,In_588,In_1015);
or U3129 (N_3129,In_1673,In_1761);
and U3130 (N_3130,In_1225,In_2239);
xor U3131 (N_3131,In_0,In_123);
xor U3132 (N_3132,In_2384,In_1623);
or U3133 (N_3133,In_1883,In_611);
nor U3134 (N_3134,In_1987,In_479);
and U3135 (N_3135,In_2318,In_920);
nor U3136 (N_3136,In_1627,In_699);
and U3137 (N_3137,In_1960,In_2012);
nor U3138 (N_3138,In_968,In_2293);
xnor U3139 (N_3139,In_1550,In_2000);
or U3140 (N_3140,In_51,In_140);
nand U3141 (N_3141,In_312,In_1835);
nand U3142 (N_3142,In_291,In_1278);
or U3143 (N_3143,In_1367,In_153);
and U3144 (N_3144,In_114,In_389);
and U3145 (N_3145,In_89,In_524);
xnor U3146 (N_3146,In_929,In_10);
nand U3147 (N_3147,In_782,In_1925);
or U3148 (N_3148,In_2190,In_1271);
nor U3149 (N_3149,In_1663,In_2357);
nand U3150 (N_3150,In_2422,In_1158);
xor U3151 (N_3151,In_1018,In_1368);
and U3152 (N_3152,In_266,In_740);
nand U3153 (N_3153,In_1727,In_2257);
nand U3154 (N_3154,In_155,In_304);
nand U3155 (N_3155,In_1616,In_1565);
or U3156 (N_3156,In_871,In_2076);
xor U3157 (N_3157,In_385,In_1162);
or U3158 (N_3158,In_1190,In_607);
or U3159 (N_3159,In_943,In_830);
xnor U3160 (N_3160,In_1872,In_2116);
and U3161 (N_3161,In_1481,In_2435);
nand U3162 (N_3162,In_1016,In_1484);
or U3163 (N_3163,In_1925,In_2402);
or U3164 (N_3164,In_823,In_961);
or U3165 (N_3165,In_1027,In_1110);
or U3166 (N_3166,In_1141,In_2261);
or U3167 (N_3167,In_442,In_740);
nand U3168 (N_3168,In_665,In_1390);
and U3169 (N_3169,In_1920,In_2145);
xor U3170 (N_3170,In_2117,In_1458);
nor U3171 (N_3171,In_2285,In_1594);
nand U3172 (N_3172,In_1247,In_2428);
and U3173 (N_3173,In_2092,In_1234);
nand U3174 (N_3174,In_1569,In_482);
xor U3175 (N_3175,In_2496,In_1763);
and U3176 (N_3176,In_1926,In_1440);
xor U3177 (N_3177,In_1949,In_989);
and U3178 (N_3178,In_2008,In_2434);
nand U3179 (N_3179,In_48,In_1033);
or U3180 (N_3180,In_1374,In_2259);
nor U3181 (N_3181,In_2494,In_1558);
or U3182 (N_3182,In_516,In_1050);
xor U3183 (N_3183,In_1533,In_595);
nand U3184 (N_3184,In_1020,In_863);
or U3185 (N_3185,In_880,In_490);
or U3186 (N_3186,In_585,In_1151);
nand U3187 (N_3187,In_651,In_104);
or U3188 (N_3188,In_900,In_1546);
nor U3189 (N_3189,In_724,In_120);
or U3190 (N_3190,In_684,In_248);
or U3191 (N_3191,In_1430,In_1267);
nor U3192 (N_3192,In_1678,In_1266);
or U3193 (N_3193,In_536,In_393);
and U3194 (N_3194,In_882,In_1108);
nand U3195 (N_3195,In_2199,In_2410);
nor U3196 (N_3196,In_504,In_26);
nand U3197 (N_3197,In_1842,In_711);
nand U3198 (N_3198,In_464,In_885);
nor U3199 (N_3199,In_128,In_1257);
and U3200 (N_3200,In_1860,In_1127);
nand U3201 (N_3201,In_558,In_2203);
nor U3202 (N_3202,In_1385,In_1106);
and U3203 (N_3203,In_530,In_2336);
or U3204 (N_3204,In_1776,In_1412);
and U3205 (N_3205,In_1056,In_826);
nand U3206 (N_3206,In_301,In_1538);
nor U3207 (N_3207,In_842,In_2363);
or U3208 (N_3208,In_724,In_440);
xnor U3209 (N_3209,In_1994,In_852);
nand U3210 (N_3210,In_1135,In_2082);
or U3211 (N_3211,In_869,In_554);
and U3212 (N_3212,In_407,In_2294);
or U3213 (N_3213,In_862,In_589);
and U3214 (N_3214,In_1673,In_1426);
or U3215 (N_3215,In_2415,In_1057);
nand U3216 (N_3216,In_2211,In_720);
nand U3217 (N_3217,In_178,In_2012);
nand U3218 (N_3218,In_590,In_1070);
or U3219 (N_3219,In_1359,In_501);
and U3220 (N_3220,In_2335,In_1629);
xnor U3221 (N_3221,In_2222,In_2168);
or U3222 (N_3222,In_1182,In_922);
nand U3223 (N_3223,In_456,In_1391);
nor U3224 (N_3224,In_1632,In_851);
or U3225 (N_3225,In_1239,In_2244);
nand U3226 (N_3226,In_1200,In_1426);
and U3227 (N_3227,In_831,In_1340);
nor U3228 (N_3228,In_2291,In_1611);
xor U3229 (N_3229,In_2340,In_1682);
nor U3230 (N_3230,In_731,In_480);
nor U3231 (N_3231,In_200,In_2085);
nor U3232 (N_3232,In_2102,In_1584);
nand U3233 (N_3233,In_2189,In_1645);
xor U3234 (N_3234,In_1985,In_2340);
xor U3235 (N_3235,In_1833,In_2004);
nand U3236 (N_3236,In_2053,In_2124);
or U3237 (N_3237,In_2213,In_2162);
nand U3238 (N_3238,In_1287,In_1030);
nand U3239 (N_3239,In_796,In_1559);
nand U3240 (N_3240,In_1654,In_2134);
nor U3241 (N_3241,In_1767,In_1195);
or U3242 (N_3242,In_1895,In_1281);
or U3243 (N_3243,In_663,In_393);
nand U3244 (N_3244,In_421,In_1636);
or U3245 (N_3245,In_660,In_59);
or U3246 (N_3246,In_2317,In_1970);
nand U3247 (N_3247,In_467,In_161);
xor U3248 (N_3248,In_1523,In_1638);
nand U3249 (N_3249,In_2119,In_953);
and U3250 (N_3250,In_893,In_854);
nor U3251 (N_3251,In_1007,In_1708);
and U3252 (N_3252,In_2329,In_363);
or U3253 (N_3253,In_2122,In_1779);
nor U3254 (N_3254,In_4,In_1479);
or U3255 (N_3255,In_2463,In_892);
nand U3256 (N_3256,In_955,In_2298);
nand U3257 (N_3257,In_177,In_1740);
and U3258 (N_3258,In_2094,In_278);
and U3259 (N_3259,In_954,In_1465);
nor U3260 (N_3260,In_131,In_1139);
nor U3261 (N_3261,In_1090,In_2383);
xnor U3262 (N_3262,In_656,In_1543);
nand U3263 (N_3263,In_1752,In_2306);
or U3264 (N_3264,In_1611,In_258);
xor U3265 (N_3265,In_922,In_1054);
nand U3266 (N_3266,In_562,In_678);
and U3267 (N_3267,In_1287,In_755);
xor U3268 (N_3268,In_548,In_490);
nor U3269 (N_3269,In_770,In_836);
xor U3270 (N_3270,In_312,In_563);
nand U3271 (N_3271,In_2372,In_487);
nor U3272 (N_3272,In_774,In_731);
nor U3273 (N_3273,In_2069,In_1230);
xor U3274 (N_3274,In_118,In_1009);
and U3275 (N_3275,In_343,In_355);
nor U3276 (N_3276,In_581,In_1802);
nand U3277 (N_3277,In_1688,In_1923);
or U3278 (N_3278,In_499,In_300);
nor U3279 (N_3279,In_556,In_2114);
or U3280 (N_3280,In_1911,In_577);
nand U3281 (N_3281,In_785,In_789);
nor U3282 (N_3282,In_597,In_1804);
xnor U3283 (N_3283,In_876,In_2069);
nand U3284 (N_3284,In_710,In_1666);
or U3285 (N_3285,In_2427,In_43);
and U3286 (N_3286,In_517,In_1549);
and U3287 (N_3287,In_2132,In_1896);
or U3288 (N_3288,In_2081,In_135);
or U3289 (N_3289,In_1387,In_600);
nand U3290 (N_3290,In_1715,In_1587);
xor U3291 (N_3291,In_784,In_2285);
xnor U3292 (N_3292,In_275,In_1935);
and U3293 (N_3293,In_1448,In_892);
xor U3294 (N_3294,In_1884,In_47);
xnor U3295 (N_3295,In_1016,In_2182);
or U3296 (N_3296,In_2403,In_528);
nor U3297 (N_3297,In_2482,In_384);
and U3298 (N_3298,In_1912,In_683);
xnor U3299 (N_3299,In_1615,In_1021);
or U3300 (N_3300,In_2490,In_527);
and U3301 (N_3301,In_755,In_1393);
nand U3302 (N_3302,In_2232,In_2295);
nor U3303 (N_3303,In_2495,In_1424);
or U3304 (N_3304,In_1274,In_1115);
nand U3305 (N_3305,In_2069,In_1536);
and U3306 (N_3306,In_2472,In_419);
xnor U3307 (N_3307,In_453,In_1718);
and U3308 (N_3308,In_1791,In_1081);
or U3309 (N_3309,In_2003,In_1713);
nand U3310 (N_3310,In_2304,In_921);
and U3311 (N_3311,In_690,In_1093);
nor U3312 (N_3312,In_1020,In_224);
or U3313 (N_3313,In_1871,In_1968);
nand U3314 (N_3314,In_1982,In_1267);
or U3315 (N_3315,In_135,In_1574);
nand U3316 (N_3316,In_1229,In_2370);
nand U3317 (N_3317,In_2082,In_1887);
and U3318 (N_3318,In_2026,In_1128);
xor U3319 (N_3319,In_1928,In_557);
or U3320 (N_3320,In_909,In_215);
nor U3321 (N_3321,In_2413,In_1980);
xor U3322 (N_3322,In_195,In_992);
and U3323 (N_3323,In_1058,In_2186);
nand U3324 (N_3324,In_581,In_2327);
nand U3325 (N_3325,In_1076,In_2472);
nor U3326 (N_3326,In_657,In_976);
xor U3327 (N_3327,In_579,In_991);
xor U3328 (N_3328,In_1784,In_709);
and U3329 (N_3329,In_2442,In_283);
nor U3330 (N_3330,In_1213,In_614);
and U3331 (N_3331,In_2029,In_1706);
nand U3332 (N_3332,In_15,In_2039);
or U3333 (N_3333,In_1712,In_35);
xor U3334 (N_3334,In_1178,In_732);
xor U3335 (N_3335,In_1181,In_702);
xor U3336 (N_3336,In_978,In_31);
nand U3337 (N_3337,In_473,In_572);
and U3338 (N_3338,In_38,In_1417);
and U3339 (N_3339,In_915,In_682);
or U3340 (N_3340,In_1126,In_298);
nand U3341 (N_3341,In_1850,In_238);
nor U3342 (N_3342,In_27,In_1789);
nor U3343 (N_3343,In_1033,In_1059);
xor U3344 (N_3344,In_2009,In_882);
nor U3345 (N_3345,In_1572,In_833);
and U3346 (N_3346,In_65,In_711);
nor U3347 (N_3347,In_537,In_1825);
xor U3348 (N_3348,In_1042,In_213);
or U3349 (N_3349,In_628,In_36);
xnor U3350 (N_3350,In_2369,In_2230);
nand U3351 (N_3351,In_1451,In_245);
xor U3352 (N_3352,In_606,In_1993);
nand U3353 (N_3353,In_1872,In_979);
xor U3354 (N_3354,In_811,In_216);
xor U3355 (N_3355,In_2378,In_131);
or U3356 (N_3356,In_412,In_1176);
nor U3357 (N_3357,In_235,In_381);
nor U3358 (N_3358,In_218,In_174);
xnor U3359 (N_3359,In_1694,In_1638);
or U3360 (N_3360,In_1753,In_2375);
xnor U3361 (N_3361,In_1317,In_2414);
or U3362 (N_3362,In_1983,In_577);
nor U3363 (N_3363,In_423,In_1764);
or U3364 (N_3364,In_222,In_1162);
and U3365 (N_3365,In_1170,In_438);
and U3366 (N_3366,In_2020,In_1761);
nor U3367 (N_3367,In_843,In_827);
nand U3368 (N_3368,In_58,In_1130);
and U3369 (N_3369,In_1317,In_1599);
nand U3370 (N_3370,In_947,In_2238);
xnor U3371 (N_3371,In_1406,In_2315);
or U3372 (N_3372,In_475,In_1998);
and U3373 (N_3373,In_2473,In_660);
nor U3374 (N_3374,In_2027,In_1925);
nor U3375 (N_3375,In_2495,In_2410);
or U3376 (N_3376,In_580,In_71);
or U3377 (N_3377,In_2064,In_1489);
or U3378 (N_3378,In_1959,In_1180);
nand U3379 (N_3379,In_726,In_1250);
xnor U3380 (N_3380,In_789,In_864);
and U3381 (N_3381,In_1225,In_1128);
or U3382 (N_3382,In_1989,In_227);
and U3383 (N_3383,In_2029,In_1627);
or U3384 (N_3384,In_1104,In_111);
nor U3385 (N_3385,In_2159,In_1584);
nor U3386 (N_3386,In_2435,In_1172);
nand U3387 (N_3387,In_198,In_29);
nor U3388 (N_3388,In_1300,In_368);
nor U3389 (N_3389,In_2093,In_1295);
and U3390 (N_3390,In_1098,In_1651);
xor U3391 (N_3391,In_1461,In_1707);
xnor U3392 (N_3392,In_1744,In_1988);
nand U3393 (N_3393,In_2371,In_1836);
xor U3394 (N_3394,In_373,In_274);
nor U3395 (N_3395,In_2378,In_1797);
nand U3396 (N_3396,In_1226,In_2043);
nand U3397 (N_3397,In_1776,In_1777);
and U3398 (N_3398,In_611,In_708);
nor U3399 (N_3399,In_1424,In_871);
nand U3400 (N_3400,In_325,In_715);
and U3401 (N_3401,In_1322,In_2037);
or U3402 (N_3402,In_551,In_2090);
nand U3403 (N_3403,In_1378,In_672);
nor U3404 (N_3404,In_2462,In_2391);
nand U3405 (N_3405,In_1904,In_1461);
or U3406 (N_3406,In_857,In_908);
xnor U3407 (N_3407,In_1818,In_2111);
nor U3408 (N_3408,In_252,In_120);
nor U3409 (N_3409,In_1999,In_446);
and U3410 (N_3410,In_191,In_2425);
nand U3411 (N_3411,In_321,In_146);
or U3412 (N_3412,In_1184,In_562);
xnor U3413 (N_3413,In_321,In_2006);
nor U3414 (N_3414,In_1053,In_443);
nor U3415 (N_3415,In_2306,In_1527);
nor U3416 (N_3416,In_1736,In_861);
xor U3417 (N_3417,In_1823,In_2336);
and U3418 (N_3418,In_1533,In_2229);
or U3419 (N_3419,In_1422,In_326);
nand U3420 (N_3420,In_1320,In_1218);
or U3421 (N_3421,In_375,In_2243);
nand U3422 (N_3422,In_1854,In_988);
or U3423 (N_3423,In_127,In_1886);
xnor U3424 (N_3424,In_1186,In_1819);
xnor U3425 (N_3425,In_1597,In_2429);
nor U3426 (N_3426,In_1381,In_1867);
and U3427 (N_3427,In_2350,In_2307);
xor U3428 (N_3428,In_2314,In_2131);
xnor U3429 (N_3429,In_1422,In_241);
xor U3430 (N_3430,In_1581,In_995);
nor U3431 (N_3431,In_1456,In_732);
nand U3432 (N_3432,In_35,In_1698);
nor U3433 (N_3433,In_2147,In_1264);
or U3434 (N_3434,In_1084,In_1541);
nand U3435 (N_3435,In_675,In_1915);
nor U3436 (N_3436,In_1385,In_250);
nand U3437 (N_3437,In_930,In_143);
or U3438 (N_3438,In_382,In_521);
xor U3439 (N_3439,In_2406,In_1456);
xor U3440 (N_3440,In_1515,In_1413);
xnor U3441 (N_3441,In_1821,In_59);
nand U3442 (N_3442,In_767,In_900);
nand U3443 (N_3443,In_2053,In_1702);
or U3444 (N_3444,In_1460,In_844);
or U3445 (N_3445,In_112,In_2154);
and U3446 (N_3446,In_1694,In_1212);
and U3447 (N_3447,In_1525,In_1710);
and U3448 (N_3448,In_471,In_1602);
nor U3449 (N_3449,In_670,In_1663);
xnor U3450 (N_3450,In_1948,In_287);
or U3451 (N_3451,In_2385,In_866);
nand U3452 (N_3452,In_2027,In_381);
nand U3453 (N_3453,In_1157,In_292);
or U3454 (N_3454,In_1786,In_341);
nand U3455 (N_3455,In_779,In_306);
nand U3456 (N_3456,In_2343,In_1532);
or U3457 (N_3457,In_135,In_2378);
xnor U3458 (N_3458,In_1354,In_519);
or U3459 (N_3459,In_1220,In_1619);
or U3460 (N_3460,In_2186,In_1201);
nor U3461 (N_3461,In_1134,In_2112);
and U3462 (N_3462,In_1980,In_953);
xor U3463 (N_3463,In_1205,In_312);
and U3464 (N_3464,In_732,In_1239);
or U3465 (N_3465,In_574,In_18);
or U3466 (N_3466,In_797,In_547);
nor U3467 (N_3467,In_235,In_798);
nor U3468 (N_3468,In_464,In_1093);
nor U3469 (N_3469,In_267,In_774);
nor U3470 (N_3470,In_33,In_679);
or U3471 (N_3471,In_1910,In_2256);
nand U3472 (N_3472,In_546,In_615);
xor U3473 (N_3473,In_1111,In_612);
or U3474 (N_3474,In_1483,In_2445);
nand U3475 (N_3475,In_138,In_2143);
or U3476 (N_3476,In_82,In_477);
and U3477 (N_3477,In_1036,In_1184);
and U3478 (N_3478,In_66,In_68);
and U3479 (N_3479,In_1083,In_2300);
and U3480 (N_3480,In_1653,In_2219);
xor U3481 (N_3481,In_1817,In_1239);
nor U3482 (N_3482,In_951,In_855);
xnor U3483 (N_3483,In_1568,In_1389);
or U3484 (N_3484,In_836,In_1348);
nor U3485 (N_3485,In_1248,In_1390);
and U3486 (N_3486,In_776,In_865);
nand U3487 (N_3487,In_2436,In_163);
nor U3488 (N_3488,In_1561,In_1298);
xnor U3489 (N_3489,In_696,In_1586);
and U3490 (N_3490,In_1767,In_2139);
nor U3491 (N_3491,In_1769,In_502);
and U3492 (N_3492,In_2051,In_720);
or U3493 (N_3493,In_1349,In_2096);
and U3494 (N_3494,In_1810,In_993);
xnor U3495 (N_3495,In_1087,In_1179);
xor U3496 (N_3496,In_1071,In_906);
or U3497 (N_3497,In_1922,In_2210);
nor U3498 (N_3498,In_28,In_1917);
or U3499 (N_3499,In_283,In_1552);
or U3500 (N_3500,In_1578,In_1255);
xor U3501 (N_3501,In_1965,In_570);
and U3502 (N_3502,In_1119,In_1303);
and U3503 (N_3503,In_2436,In_2117);
nand U3504 (N_3504,In_826,In_871);
nand U3505 (N_3505,In_1774,In_243);
nor U3506 (N_3506,In_515,In_93);
nor U3507 (N_3507,In_679,In_1317);
nand U3508 (N_3508,In_2358,In_43);
nand U3509 (N_3509,In_2059,In_55);
and U3510 (N_3510,In_313,In_1703);
nand U3511 (N_3511,In_2353,In_1322);
and U3512 (N_3512,In_392,In_1917);
xnor U3513 (N_3513,In_1857,In_1520);
or U3514 (N_3514,In_2381,In_1452);
and U3515 (N_3515,In_2385,In_388);
nand U3516 (N_3516,In_895,In_1786);
xor U3517 (N_3517,In_2331,In_2351);
or U3518 (N_3518,In_934,In_2199);
and U3519 (N_3519,In_2335,In_1354);
and U3520 (N_3520,In_1788,In_281);
nor U3521 (N_3521,In_1753,In_355);
and U3522 (N_3522,In_1668,In_1448);
or U3523 (N_3523,In_2079,In_562);
nand U3524 (N_3524,In_228,In_1599);
xor U3525 (N_3525,In_2384,In_694);
and U3526 (N_3526,In_149,In_1406);
or U3527 (N_3527,In_1951,In_862);
and U3528 (N_3528,In_383,In_1217);
or U3529 (N_3529,In_738,In_2036);
xor U3530 (N_3530,In_931,In_1443);
nor U3531 (N_3531,In_2304,In_1233);
and U3532 (N_3532,In_1064,In_605);
nand U3533 (N_3533,In_28,In_879);
nand U3534 (N_3534,In_1062,In_995);
nand U3535 (N_3535,In_1280,In_113);
or U3536 (N_3536,In_758,In_211);
xor U3537 (N_3537,In_33,In_2025);
and U3538 (N_3538,In_2417,In_1092);
xor U3539 (N_3539,In_273,In_9);
and U3540 (N_3540,In_2212,In_14);
or U3541 (N_3541,In_326,In_2481);
nor U3542 (N_3542,In_2210,In_206);
nor U3543 (N_3543,In_2343,In_1584);
nor U3544 (N_3544,In_2122,In_1086);
nand U3545 (N_3545,In_1019,In_232);
xor U3546 (N_3546,In_246,In_2112);
xor U3547 (N_3547,In_790,In_480);
and U3548 (N_3548,In_2077,In_777);
nor U3549 (N_3549,In_1367,In_1610);
nor U3550 (N_3550,In_2144,In_2117);
or U3551 (N_3551,In_1151,In_942);
nor U3552 (N_3552,In_1981,In_2321);
xor U3553 (N_3553,In_1239,In_850);
and U3554 (N_3554,In_734,In_80);
nand U3555 (N_3555,In_286,In_2153);
xor U3556 (N_3556,In_574,In_928);
nand U3557 (N_3557,In_1339,In_2139);
or U3558 (N_3558,In_2244,In_1865);
xor U3559 (N_3559,In_877,In_403);
or U3560 (N_3560,In_120,In_1476);
nand U3561 (N_3561,In_1615,In_196);
xnor U3562 (N_3562,In_56,In_485);
or U3563 (N_3563,In_1567,In_2156);
and U3564 (N_3564,In_100,In_1514);
nor U3565 (N_3565,In_819,In_880);
and U3566 (N_3566,In_15,In_848);
nor U3567 (N_3567,In_1844,In_1563);
or U3568 (N_3568,In_1877,In_2244);
and U3569 (N_3569,In_1722,In_2363);
nor U3570 (N_3570,In_2179,In_41);
and U3571 (N_3571,In_36,In_557);
or U3572 (N_3572,In_2001,In_1106);
nand U3573 (N_3573,In_1333,In_931);
or U3574 (N_3574,In_599,In_1356);
xor U3575 (N_3575,In_613,In_769);
nor U3576 (N_3576,In_2133,In_910);
and U3577 (N_3577,In_167,In_895);
and U3578 (N_3578,In_857,In_1725);
or U3579 (N_3579,In_2485,In_1721);
or U3580 (N_3580,In_1706,In_2011);
xnor U3581 (N_3581,In_681,In_1695);
nand U3582 (N_3582,In_86,In_1942);
and U3583 (N_3583,In_1540,In_236);
or U3584 (N_3584,In_1023,In_1818);
nor U3585 (N_3585,In_1671,In_404);
or U3586 (N_3586,In_862,In_2347);
or U3587 (N_3587,In_2003,In_1893);
nand U3588 (N_3588,In_1414,In_1093);
nor U3589 (N_3589,In_1285,In_2255);
nor U3590 (N_3590,In_1029,In_1286);
or U3591 (N_3591,In_484,In_1167);
nor U3592 (N_3592,In_1681,In_494);
or U3593 (N_3593,In_751,In_2111);
xor U3594 (N_3594,In_1970,In_1060);
and U3595 (N_3595,In_413,In_734);
xnor U3596 (N_3596,In_1610,In_2300);
nor U3597 (N_3597,In_2235,In_1503);
and U3598 (N_3598,In_697,In_1501);
nand U3599 (N_3599,In_1249,In_1574);
and U3600 (N_3600,In_60,In_739);
nor U3601 (N_3601,In_338,In_808);
nand U3602 (N_3602,In_1677,In_2387);
xnor U3603 (N_3603,In_398,In_2023);
nor U3604 (N_3604,In_1934,In_2467);
and U3605 (N_3605,In_955,In_1477);
nor U3606 (N_3606,In_2074,In_1277);
nand U3607 (N_3607,In_542,In_2446);
xor U3608 (N_3608,In_1818,In_108);
and U3609 (N_3609,In_394,In_1977);
or U3610 (N_3610,In_875,In_2221);
nand U3611 (N_3611,In_603,In_572);
nand U3612 (N_3612,In_1188,In_1539);
nand U3613 (N_3613,In_1778,In_1602);
or U3614 (N_3614,In_678,In_619);
or U3615 (N_3615,In_1265,In_789);
or U3616 (N_3616,In_1752,In_2471);
xor U3617 (N_3617,In_848,In_196);
and U3618 (N_3618,In_1982,In_2352);
nand U3619 (N_3619,In_2179,In_2377);
xor U3620 (N_3620,In_1551,In_2386);
or U3621 (N_3621,In_851,In_1100);
and U3622 (N_3622,In_2372,In_2015);
nor U3623 (N_3623,In_1481,In_1740);
and U3624 (N_3624,In_2077,In_656);
nor U3625 (N_3625,In_1797,In_2432);
nand U3626 (N_3626,In_1013,In_2497);
nand U3627 (N_3627,In_1536,In_2300);
and U3628 (N_3628,In_1130,In_2094);
nor U3629 (N_3629,In_2173,In_263);
and U3630 (N_3630,In_130,In_2380);
and U3631 (N_3631,In_788,In_514);
nor U3632 (N_3632,In_2032,In_1078);
xor U3633 (N_3633,In_1255,In_515);
xnor U3634 (N_3634,In_616,In_1764);
nand U3635 (N_3635,In_2311,In_234);
nand U3636 (N_3636,In_2228,In_159);
xor U3637 (N_3637,In_1767,In_1029);
nand U3638 (N_3638,In_1920,In_2322);
or U3639 (N_3639,In_2134,In_2484);
xor U3640 (N_3640,In_2068,In_1937);
and U3641 (N_3641,In_1117,In_1887);
or U3642 (N_3642,In_462,In_695);
nand U3643 (N_3643,In_2265,In_223);
or U3644 (N_3644,In_2453,In_794);
and U3645 (N_3645,In_110,In_1287);
and U3646 (N_3646,In_1208,In_1923);
and U3647 (N_3647,In_1609,In_2242);
and U3648 (N_3648,In_296,In_1212);
and U3649 (N_3649,In_1491,In_1202);
or U3650 (N_3650,In_613,In_1895);
nand U3651 (N_3651,In_1743,In_77);
and U3652 (N_3652,In_1186,In_913);
and U3653 (N_3653,In_1291,In_800);
nand U3654 (N_3654,In_495,In_1637);
and U3655 (N_3655,In_2337,In_2345);
and U3656 (N_3656,In_1394,In_747);
xor U3657 (N_3657,In_152,In_559);
nor U3658 (N_3658,In_1054,In_237);
xnor U3659 (N_3659,In_1307,In_1152);
xnor U3660 (N_3660,In_1084,In_1549);
or U3661 (N_3661,In_2318,In_237);
nand U3662 (N_3662,In_2041,In_669);
and U3663 (N_3663,In_2391,In_2224);
nand U3664 (N_3664,In_682,In_609);
and U3665 (N_3665,In_2343,In_2415);
nor U3666 (N_3666,In_1670,In_1311);
nor U3667 (N_3667,In_2298,In_2249);
nand U3668 (N_3668,In_2408,In_1654);
xnor U3669 (N_3669,In_1436,In_1659);
nor U3670 (N_3670,In_1966,In_966);
nand U3671 (N_3671,In_926,In_1160);
nor U3672 (N_3672,In_1683,In_1605);
nor U3673 (N_3673,In_1970,In_112);
and U3674 (N_3674,In_2136,In_1857);
or U3675 (N_3675,In_1938,In_1811);
xnor U3676 (N_3676,In_1027,In_1161);
and U3677 (N_3677,In_794,In_1182);
nand U3678 (N_3678,In_2430,In_869);
nor U3679 (N_3679,In_409,In_1962);
or U3680 (N_3680,In_2261,In_1423);
nand U3681 (N_3681,In_1514,In_816);
xor U3682 (N_3682,In_2111,In_1088);
nand U3683 (N_3683,In_1104,In_833);
xnor U3684 (N_3684,In_2334,In_1241);
or U3685 (N_3685,In_401,In_433);
nand U3686 (N_3686,In_1021,In_1556);
nor U3687 (N_3687,In_1919,In_1477);
and U3688 (N_3688,In_849,In_1874);
or U3689 (N_3689,In_1285,In_605);
or U3690 (N_3690,In_1281,In_991);
nand U3691 (N_3691,In_431,In_443);
nand U3692 (N_3692,In_1491,In_1997);
and U3693 (N_3693,In_1198,In_2122);
or U3694 (N_3694,In_1908,In_1626);
xnor U3695 (N_3695,In_1654,In_1323);
or U3696 (N_3696,In_1195,In_282);
and U3697 (N_3697,In_528,In_137);
and U3698 (N_3698,In_1952,In_504);
or U3699 (N_3699,In_473,In_513);
nor U3700 (N_3700,In_1615,In_1901);
and U3701 (N_3701,In_1798,In_2349);
xnor U3702 (N_3702,In_801,In_977);
xnor U3703 (N_3703,In_1574,In_1066);
nand U3704 (N_3704,In_1414,In_26);
xnor U3705 (N_3705,In_1376,In_1753);
and U3706 (N_3706,In_246,In_1759);
nor U3707 (N_3707,In_543,In_2144);
nand U3708 (N_3708,In_901,In_1977);
and U3709 (N_3709,In_646,In_1227);
and U3710 (N_3710,In_724,In_2278);
or U3711 (N_3711,In_824,In_680);
xor U3712 (N_3712,In_25,In_519);
and U3713 (N_3713,In_2008,In_127);
nand U3714 (N_3714,In_118,In_1974);
and U3715 (N_3715,In_1238,In_1450);
xor U3716 (N_3716,In_440,In_1452);
or U3717 (N_3717,In_103,In_2427);
xnor U3718 (N_3718,In_539,In_294);
and U3719 (N_3719,In_808,In_96);
xor U3720 (N_3720,In_962,In_2130);
or U3721 (N_3721,In_2124,In_1584);
nand U3722 (N_3722,In_644,In_2310);
nor U3723 (N_3723,In_2289,In_177);
nor U3724 (N_3724,In_1637,In_270);
xor U3725 (N_3725,In_2300,In_2077);
nor U3726 (N_3726,In_350,In_2221);
nor U3727 (N_3727,In_1958,In_744);
xnor U3728 (N_3728,In_2106,In_370);
or U3729 (N_3729,In_465,In_1239);
nand U3730 (N_3730,In_484,In_309);
xnor U3731 (N_3731,In_745,In_331);
nor U3732 (N_3732,In_1622,In_349);
and U3733 (N_3733,In_1518,In_1492);
xnor U3734 (N_3734,In_1678,In_2423);
nand U3735 (N_3735,In_1186,In_965);
or U3736 (N_3736,In_1630,In_2377);
nand U3737 (N_3737,In_1557,In_605);
nand U3738 (N_3738,In_1906,In_965);
nor U3739 (N_3739,In_2220,In_783);
or U3740 (N_3740,In_827,In_358);
or U3741 (N_3741,In_665,In_2137);
nor U3742 (N_3742,In_1280,In_679);
xnor U3743 (N_3743,In_2418,In_174);
nand U3744 (N_3744,In_2122,In_1593);
or U3745 (N_3745,In_1639,In_2432);
and U3746 (N_3746,In_1978,In_2243);
xor U3747 (N_3747,In_1772,In_78);
or U3748 (N_3748,In_76,In_611);
nor U3749 (N_3749,In_631,In_2302);
and U3750 (N_3750,In_1124,In_801);
xnor U3751 (N_3751,In_852,In_2470);
nand U3752 (N_3752,In_2427,In_1558);
or U3753 (N_3753,In_94,In_2069);
and U3754 (N_3754,In_791,In_1423);
xnor U3755 (N_3755,In_1676,In_1117);
nand U3756 (N_3756,In_1,In_452);
nor U3757 (N_3757,In_1833,In_2051);
xor U3758 (N_3758,In_2499,In_1218);
xor U3759 (N_3759,In_1063,In_532);
xor U3760 (N_3760,In_1080,In_2071);
nand U3761 (N_3761,In_2272,In_971);
and U3762 (N_3762,In_1316,In_1479);
nor U3763 (N_3763,In_1217,In_1370);
nand U3764 (N_3764,In_1493,In_1726);
nand U3765 (N_3765,In_635,In_146);
nor U3766 (N_3766,In_684,In_863);
nor U3767 (N_3767,In_836,In_1645);
nor U3768 (N_3768,In_2036,In_378);
xor U3769 (N_3769,In_68,In_2224);
xnor U3770 (N_3770,In_1446,In_2376);
nor U3771 (N_3771,In_1212,In_856);
nand U3772 (N_3772,In_600,In_2397);
nor U3773 (N_3773,In_853,In_1727);
nand U3774 (N_3774,In_1572,In_2192);
xor U3775 (N_3775,In_106,In_1769);
nand U3776 (N_3776,In_1010,In_1953);
or U3777 (N_3777,In_1976,In_1816);
and U3778 (N_3778,In_2380,In_1668);
nor U3779 (N_3779,In_1445,In_2409);
or U3780 (N_3780,In_1813,In_2488);
or U3781 (N_3781,In_996,In_1403);
nor U3782 (N_3782,In_2346,In_1052);
nor U3783 (N_3783,In_1364,In_1284);
xor U3784 (N_3784,In_526,In_1732);
and U3785 (N_3785,In_589,In_637);
and U3786 (N_3786,In_475,In_1019);
nor U3787 (N_3787,In_1183,In_1661);
nand U3788 (N_3788,In_533,In_1800);
nand U3789 (N_3789,In_1511,In_2018);
xor U3790 (N_3790,In_17,In_988);
and U3791 (N_3791,In_960,In_234);
xor U3792 (N_3792,In_2293,In_1071);
xnor U3793 (N_3793,In_1371,In_430);
and U3794 (N_3794,In_1639,In_1125);
nor U3795 (N_3795,In_2461,In_1439);
and U3796 (N_3796,In_1624,In_259);
nand U3797 (N_3797,In_657,In_1617);
xnor U3798 (N_3798,In_2470,In_2196);
nand U3799 (N_3799,In_1795,In_604);
nand U3800 (N_3800,In_1278,In_1237);
nor U3801 (N_3801,In_654,In_2435);
and U3802 (N_3802,In_1714,In_2152);
or U3803 (N_3803,In_1157,In_684);
nor U3804 (N_3804,In_1782,In_1165);
xor U3805 (N_3805,In_1842,In_1162);
or U3806 (N_3806,In_747,In_2188);
xor U3807 (N_3807,In_1947,In_967);
or U3808 (N_3808,In_523,In_2467);
and U3809 (N_3809,In_414,In_47);
nor U3810 (N_3810,In_1399,In_1076);
xnor U3811 (N_3811,In_2290,In_1222);
xor U3812 (N_3812,In_1190,In_1741);
xnor U3813 (N_3813,In_2239,In_1237);
nand U3814 (N_3814,In_1306,In_1);
nor U3815 (N_3815,In_1509,In_990);
or U3816 (N_3816,In_888,In_1416);
or U3817 (N_3817,In_349,In_853);
nor U3818 (N_3818,In_57,In_1005);
or U3819 (N_3819,In_1652,In_1774);
or U3820 (N_3820,In_503,In_964);
xnor U3821 (N_3821,In_423,In_361);
nand U3822 (N_3822,In_283,In_1722);
and U3823 (N_3823,In_329,In_87);
or U3824 (N_3824,In_1658,In_1727);
and U3825 (N_3825,In_348,In_2170);
nor U3826 (N_3826,In_1059,In_233);
and U3827 (N_3827,In_54,In_1508);
and U3828 (N_3828,In_2355,In_1853);
and U3829 (N_3829,In_2171,In_638);
nand U3830 (N_3830,In_639,In_1318);
and U3831 (N_3831,In_462,In_1105);
nor U3832 (N_3832,In_644,In_657);
xnor U3833 (N_3833,In_1839,In_1197);
and U3834 (N_3834,In_64,In_266);
nand U3835 (N_3835,In_77,In_2231);
nor U3836 (N_3836,In_1943,In_991);
or U3837 (N_3837,In_2326,In_1542);
nor U3838 (N_3838,In_2020,In_768);
and U3839 (N_3839,In_1140,In_1762);
nand U3840 (N_3840,In_606,In_139);
or U3841 (N_3841,In_416,In_1419);
and U3842 (N_3842,In_2289,In_2046);
xnor U3843 (N_3843,In_1740,In_279);
xor U3844 (N_3844,In_1741,In_585);
nor U3845 (N_3845,In_1492,In_746);
nor U3846 (N_3846,In_1670,In_169);
nor U3847 (N_3847,In_455,In_840);
nand U3848 (N_3848,In_2351,In_2266);
nand U3849 (N_3849,In_306,In_2261);
nand U3850 (N_3850,In_1114,In_1479);
xor U3851 (N_3851,In_106,In_158);
nand U3852 (N_3852,In_2262,In_799);
nand U3853 (N_3853,In_1303,In_58);
xor U3854 (N_3854,In_2111,In_1624);
or U3855 (N_3855,In_953,In_2136);
xnor U3856 (N_3856,In_1353,In_1801);
and U3857 (N_3857,In_766,In_1947);
nand U3858 (N_3858,In_123,In_1129);
xnor U3859 (N_3859,In_319,In_723);
or U3860 (N_3860,In_1881,In_1353);
and U3861 (N_3861,In_1754,In_245);
xnor U3862 (N_3862,In_443,In_871);
xor U3863 (N_3863,In_908,In_765);
nand U3864 (N_3864,In_742,In_1511);
nand U3865 (N_3865,In_1025,In_1729);
or U3866 (N_3866,In_1773,In_1985);
nor U3867 (N_3867,In_232,In_1240);
nor U3868 (N_3868,In_2246,In_269);
or U3869 (N_3869,In_76,In_212);
or U3870 (N_3870,In_949,In_163);
or U3871 (N_3871,In_901,In_798);
nor U3872 (N_3872,In_994,In_988);
nor U3873 (N_3873,In_2028,In_936);
nand U3874 (N_3874,In_2008,In_2133);
xor U3875 (N_3875,In_2132,In_593);
or U3876 (N_3876,In_1918,In_1409);
or U3877 (N_3877,In_1647,In_328);
and U3878 (N_3878,In_2026,In_314);
nand U3879 (N_3879,In_905,In_18);
nor U3880 (N_3880,In_236,In_766);
and U3881 (N_3881,In_1011,In_363);
xnor U3882 (N_3882,In_1596,In_87);
nor U3883 (N_3883,In_473,In_366);
xnor U3884 (N_3884,In_2194,In_825);
nor U3885 (N_3885,In_1267,In_1215);
or U3886 (N_3886,In_873,In_2201);
xnor U3887 (N_3887,In_41,In_1193);
and U3888 (N_3888,In_1285,In_2451);
and U3889 (N_3889,In_1616,In_760);
or U3890 (N_3890,In_30,In_1088);
xor U3891 (N_3891,In_591,In_610);
xnor U3892 (N_3892,In_102,In_2140);
nand U3893 (N_3893,In_2331,In_1882);
and U3894 (N_3894,In_7,In_76);
or U3895 (N_3895,In_481,In_1154);
nand U3896 (N_3896,In_1699,In_764);
or U3897 (N_3897,In_886,In_267);
nor U3898 (N_3898,In_599,In_1633);
xnor U3899 (N_3899,In_2203,In_1551);
xor U3900 (N_3900,In_946,In_2292);
and U3901 (N_3901,In_607,In_1756);
or U3902 (N_3902,In_1369,In_2418);
nand U3903 (N_3903,In_1821,In_293);
nand U3904 (N_3904,In_953,In_354);
and U3905 (N_3905,In_878,In_338);
nand U3906 (N_3906,In_939,In_68);
nor U3907 (N_3907,In_461,In_2456);
and U3908 (N_3908,In_424,In_1930);
xor U3909 (N_3909,In_2066,In_2293);
nand U3910 (N_3910,In_273,In_2187);
nor U3911 (N_3911,In_889,In_1522);
nor U3912 (N_3912,In_1441,In_1888);
and U3913 (N_3913,In_1402,In_661);
xor U3914 (N_3914,In_1705,In_1443);
and U3915 (N_3915,In_735,In_2262);
and U3916 (N_3916,In_1026,In_1702);
xor U3917 (N_3917,In_273,In_1086);
or U3918 (N_3918,In_820,In_166);
nor U3919 (N_3919,In_500,In_1246);
xnor U3920 (N_3920,In_516,In_456);
or U3921 (N_3921,In_1015,In_371);
nor U3922 (N_3922,In_429,In_41);
or U3923 (N_3923,In_789,In_2146);
nand U3924 (N_3924,In_270,In_2325);
xnor U3925 (N_3925,In_1189,In_415);
xnor U3926 (N_3926,In_115,In_2428);
nand U3927 (N_3927,In_1749,In_713);
or U3928 (N_3928,In_1762,In_1848);
nand U3929 (N_3929,In_1702,In_834);
or U3930 (N_3930,In_2292,In_1008);
or U3931 (N_3931,In_917,In_2137);
and U3932 (N_3932,In_2365,In_1646);
and U3933 (N_3933,In_1194,In_1795);
and U3934 (N_3934,In_1292,In_1496);
and U3935 (N_3935,In_1248,In_1710);
and U3936 (N_3936,In_2043,In_1336);
or U3937 (N_3937,In_648,In_1567);
nor U3938 (N_3938,In_606,In_1821);
or U3939 (N_3939,In_282,In_1430);
or U3940 (N_3940,In_1373,In_147);
or U3941 (N_3941,In_1194,In_1946);
and U3942 (N_3942,In_1318,In_1119);
and U3943 (N_3943,In_1527,In_1328);
nor U3944 (N_3944,In_749,In_1062);
or U3945 (N_3945,In_696,In_2300);
nand U3946 (N_3946,In_723,In_2231);
or U3947 (N_3947,In_1537,In_927);
xor U3948 (N_3948,In_605,In_2143);
and U3949 (N_3949,In_817,In_348);
nand U3950 (N_3950,In_2213,In_1752);
or U3951 (N_3951,In_1089,In_477);
xnor U3952 (N_3952,In_1804,In_329);
xnor U3953 (N_3953,In_110,In_650);
xor U3954 (N_3954,In_864,In_1006);
xor U3955 (N_3955,In_1725,In_2217);
xor U3956 (N_3956,In_1341,In_783);
nand U3957 (N_3957,In_46,In_1411);
nor U3958 (N_3958,In_600,In_378);
nor U3959 (N_3959,In_2460,In_954);
nand U3960 (N_3960,In_1385,In_1669);
xnor U3961 (N_3961,In_822,In_2472);
nand U3962 (N_3962,In_73,In_103);
or U3963 (N_3963,In_808,In_642);
or U3964 (N_3964,In_1768,In_442);
xor U3965 (N_3965,In_862,In_1038);
nor U3966 (N_3966,In_75,In_636);
or U3967 (N_3967,In_1451,In_1054);
or U3968 (N_3968,In_2004,In_118);
nor U3969 (N_3969,In_618,In_2120);
nand U3970 (N_3970,In_2434,In_1217);
nor U3971 (N_3971,In_244,In_2409);
nor U3972 (N_3972,In_1282,In_273);
nor U3973 (N_3973,In_316,In_1663);
and U3974 (N_3974,In_2046,In_1999);
and U3975 (N_3975,In_396,In_785);
nand U3976 (N_3976,In_1884,In_2223);
and U3977 (N_3977,In_1065,In_1479);
nor U3978 (N_3978,In_2158,In_788);
nor U3979 (N_3979,In_1956,In_2488);
xor U3980 (N_3980,In_1691,In_2115);
or U3981 (N_3981,In_1439,In_1646);
nand U3982 (N_3982,In_100,In_168);
and U3983 (N_3983,In_1119,In_1687);
or U3984 (N_3984,In_1101,In_1449);
or U3985 (N_3985,In_275,In_796);
xnor U3986 (N_3986,In_2383,In_2366);
xor U3987 (N_3987,In_558,In_2015);
xor U3988 (N_3988,In_1027,In_1767);
nor U3989 (N_3989,In_1140,In_1353);
and U3990 (N_3990,In_399,In_363);
and U3991 (N_3991,In_205,In_1129);
xor U3992 (N_3992,In_1738,In_1207);
or U3993 (N_3993,In_446,In_2004);
xnor U3994 (N_3994,In_1007,In_1025);
nor U3995 (N_3995,In_184,In_745);
xor U3996 (N_3996,In_649,In_1222);
or U3997 (N_3997,In_999,In_736);
xor U3998 (N_3998,In_572,In_605);
or U3999 (N_3999,In_379,In_2391);
xnor U4000 (N_4000,In_1128,In_1398);
nor U4001 (N_4001,In_1656,In_478);
xnor U4002 (N_4002,In_627,In_633);
nor U4003 (N_4003,In_534,In_1889);
nor U4004 (N_4004,In_862,In_1007);
xnor U4005 (N_4005,In_391,In_643);
xor U4006 (N_4006,In_99,In_415);
or U4007 (N_4007,In_223,In_436);
and U4008 (N_4008,In_2317,In_1504);
and U4009 (N_4009,In_1601,In_239);
nand U4010 (N_4010,In_2409,In_2172);
or U4011 (N_4011,In_313,In_179);
nor U4012 (N_4012,In_1044,In_2446);
xor U4013 (N_4013,In_660,In_1663);
and U4014 (N_4014,In_1570,In_207);
or U4015 (N_4015,In_688,In_2375);
xor U4016 (N_4016,In_646,In_374);
xor U4017 (N_4017,In_2073,In_1848);
xor U4018 (N_4018,In_698,In_600);
nor U4019 (N_4019,In_2185,In_1588);
and U4020 (N_4020,In_627,In_1739);
or U4021 (N_4021,In_1663,In_265);
or U4022 (N_4022,In_1487,In_1420);
nand U4023 (N_4023,In_2263,In_2394);
nand U4024 (N_4024,In_2468,In_2363);
and U4025 (N_4025,In_1107,In_2081);
or U4026 (N_4026,In_1097,In_246);
or U4027 (N_4027,In_931,In_948);
nor U4028 (N_4028,In_1936,In_1961);
xor U4029 (N_4029,In_495,In_2192);
or U4030 (N_4030,In_1141,In_512);
nor U4031 (N_4031,In_2234,In_2301);
nand U4032 (N_4032,In_241,In_1945);
nand U4033 (N_4033,In_1275,In_676);
nand U4034 (N_4034,In_252,In_2049);
nand U4035 (N_4035,In_2331,In_1908);
and U4036 (N_4036,In_1782,In_2263);
nor U4037 (N_4037,In_1657,In_2464);
nand U4038 (N_4038,In_1910,In_380);
nor U4039 (N_4039,In_2450,In_1777);
or U4040 (N_4040,In_411,In_1413);
or U4041 (N_4041,In_332,In_1925);
xnor U4042 (N_4042,In_1423,In_1125);
nand U4043 (N_4043,In_485,In_2045);
nand U4044 (N_4044,In_1748,In_1608);
or U4045 (N_4045,In_1139,In_1958);
and U4046 (N_4046,In_1919,In_1902);
and U4047 (N_4047,In_135,In_2171);
xnor U4048 (N_4048,In_610,In_1927);
xor U4049 (N_4049,In_1184,In_1920);
or U4050 (N_4050,In_501,In_1315);
nand U4051 (N_4051,In_1723,In_680);
and U4052 (N_4052,In_2136,In_1967);
nor U4053 (N_4053,In_1834,In_874);
or U4054 (N_4054,In_2324,In_740);
or U4055 (N_4055,In_341,In_188);
xnor U4056 (N_4056,In_961,In_954);
nor U4057 (N_4057,In_529,In_751);
nand U4058 (N_4058,In_1223,In_1025);
nand U4059 (N_4059,In_2302,In_1170);
nor U4060 (N_4060,In_1332,In_1707);
or U4061 (N_4061,In_377,In_610);
and U4062 (N_4062,In_1377,In_1788);
and U4063 (N_4063,In_2030,In_1786);
nor U4064 (N_4064,In_413,In_1920);
or U4065 (N_4065,In_871,In_181);
and U4066 (N_4066,In_953,In_1841);
and U4067 (N_4067,In_2378,In_1356);
xor U4068 (N_4068,In_2216,In_921);
or U4069 (N_4069,In_1048,In_1815);
nor U4070 (N_4070,In_857,In_1938);
and U4071 (N_4071,In_2017,In_1984);
or U4072 (N_4072,In_174,In_3);
xor U4073 (N_4073,In_2195,In_1177);
and U4074 (N_4074,In_360,In_1031);
and U4075 (N_4075,In_488,In_445);
and U4076 (N_4076,In_385,In_929);
nand U4077 (N_4077,In_1473,In_691);
nor U4078 (N_4078,In_1512,In_879);
nand U4079 (N_4079,In_879,In_903);
or U4080 (N_4080,In_1858,In_320);
and U4081 (N_4081,In_1127,In_2228);
nand U4082 (N_4082,In_1179,In_273);
xnor U4083 (N_4083,In_142,In_2351);
nand U4084 (N_4084,In_451,In_855);
and U4085 (N_4085,In_70,In_2289);
and U4086 (N_4086,In_1872,In_279);
nor U4087 (N_4087,In_1545,In_1011);
nor U4088 (N_4088,In_399,In_971);
nand U4089 (N_4089,In_179,In_737);
nand U4090 (N_4090,In_276,In_1071);
nand U4091 (N_4091,In_2289,In_1638);
xor U4092 (N_4092,In_702,In_2296);
nand U4093 (N_4093,In_1692,In_1952);
nor U4094 (N_4094,In_1015,In_1091);
xnor U4095 (N_4095,In_169,In_2004);
nand U4096 (N_4096,In_1193,In_1227);
xnor U4097 (N_4097,In_1316,In_750);
nor U4098 (N_4098,In_1203,In_1541);
xnor U4099 (N_4099,In_287,In_113);
and U4100 (N_4100,In_1532,In_1865);
nor U4101 (N_4101,In_1683,In_2495);
xnor U4102 (N_4102,In_2253,In_2203);
or U4103 (N_4103,In_2167,In_2247);
nor U4104 (N_4104,In_611,In_228);
nand U4105 (N_4105,In_1377,In_1613);
xor U4106 (N_4106,In_1795,In_1156);
and U4107 (N_4107,In_2466,In_1087);
nand U4108 (N_4108,In_1966,In_559);
xnor U4109 (N_4109,In_2155,In_1604);
nor U4110 (N_4110,In_8,In_1308);
or U4111 (N_4111,In_1852,In_2);
nand U4112 (N_4112,In_1576,In_554);
or U4113 (N_4113,In_1569,In_749);
and U4114 (N_4114,In_626,In_1422);
nand U4115 (N_4115,In_768,In_490);
or U4116 (N_4116,In_149,In_1635);
or U4117 (N_4117,In_914,In_821);
and U4118 (N_4118,In_2147,In_1211);
nand U4119 (N_4119,In_673,In_137);
and U4120 (N_4120,In_470,In_2261);
nor U4121 (N_4121,In_1338,In_174);
xnor U4122 (N_4122,In_1845,In_286);
nor U4123 (N_4123,In_977,In_12);
nor U4124 (N_4124,In_790,In_1083);
or U4125 (N_4125,In_2189,In_2011);
nand U4126 (N_4126,In_421,In_1026);
xnor U4127 (N_4127,In_310,In_579);
xnor U4128 (N_4128,In_341,In_1630);
nor U4129 (N_4129,In_1747,In_887);
xnor U4130 (N_4130,In_1898,In_455);
nor U4131 (N_4131,In_1074,In_774);
nor U4132 (N_4132,In_2362,In_821);
or U4133 (N_4133,In_1803,In_185);
nand U4134 (N_4134,In_1810,In_1819);
or U4135 (N_4135,In_1005,In_914);
or U4136 (N_4136,In_2047,In_2084);
and U4137 (N_4137,In_1574,In_597);
and U4138 (N_4138,In_1370,In_970);
or U4139 (N_4139,In_786,In_484);
xor U4140 (N_4140,In_2453,In_1837);
nor U4141 (N_4141,In_492,In_1187);
or U4142 (N_4142,In_302,In_1621);
nor U4143 (N_4143,In_1872,In_921);
nor U4144 (N_4144,In_821,In_1353);
nand U4145 (N_4145,In_1085,In_796);
and U4146 (N_4146,In_207,In_1034);
xnor U4147 (N_4147,In_1400,In_1531);
xor U4148 (N_4148,In_1507,In_1259);
nand U4149 (N_4149,In_1153,In_1393);
nor U4150 (N_4150,In_840,In_1141);
and U4151 (N_4151,In_1384,In_1409);
and U4152 (N_4152,In_1981,In_183);
nor U4153 (N_4153,In_405,In_1325);
or U4154 (N_4154,In_2092,In_1947);
nor U4155 (N_4155,In_84,In_760);
xor U4156 (N_4156,In_2261,In_2367);
nor U4157 (N_4157,In_1385,In_920);
nor U4158 (N_4158,In_1907,In_1910);
nand U4159 (N_4159,In_1011,In_628);
or U4160 (N_4160,In_71,In_1602);
or U4161 (N_4161,In_222,In_2434);
and U4162 (N_4162,In_2350,In_1165);
and U4163 (N_4163,In_1804,In_1113);
nand U4164 (N_4164,In_1667,In_1070);
or U4165 (N_4165,In_2273,In_2028);
nand U4166 (N_4166,In_493,In_1915);
nor U4167 (N_4167,In_367,In_2130);
and U4168 (N_4168,In_1538,In_101);
nand U4169 (N_4169,In_2005,In_1772);
or U4170 (N_4170,In_569,In_406);
or U4171 (N_4171,In_1146,In_498);
and U4172 (N_4172,In_2431,In_1376);
nor U4173 (N_4173,In_840,In_309);
or U4174 (N_4174,In_82,In_2070);
xnor U4175 (N_4175,In_2219,In_988);
nand U4176 (N_4176,In_673,In_608);
or U4177 (N_4177,In_1765,In_1672);
and U4178 (N_4178,In_1014,In_781);
nand U4179 (N_4179,In_1354,In_219);
nand U4180 (N_4180,In_2043,In_1715);
nor U4181 (N_4181,In_770,In_1005);
and U4182 (N_4182,In_1891,In_2029);
xnor U4183 (N_4183,In_59,In_1569);
nand U4184 (N_4184,In_385,In_1703);
and U4185 (N_4185,In_1098,In_2074);
and U4186 (N_4186,In_1203,In_1515);
nand U4187 (N_4187,In_2374,In_1678);
or U4188 (N_4188,In_2402,In_2132);
or U4189 (N_4189,In_1193,In_2014);
nand U4190 (N_4190,In_1833,In_2243);
nor U4191 (N_4191,In_542,In_88);
or U4192 (N_4192,In_955,In_445);
xnor U4193 (N_4193,In_710,In_2252);
xnor U4194 (N_4194,In_2122,In_1857);
nand U4195 (N_4195,In_306,In_680);
nor U4196 (N_4196,In_993,In_1334);
and U4197 (N_4197,In_2234,In_333);
or U4198 (N_4198,In_421,In_1300);
and U4199 (N_4199,In_977,In_1368);
nor U4200 (N_4200,In_1513,In_2416);
nand U4201 (N_4201,In_1261,In_962);
or U4202 (N_4202,In_452,In_1120);
or U4203 (N_4203,In_2484,In_2318);
nand U4204 (N_4204,In_937,In_1395);
or U4205 (N_4205,In_723,In_455);
xnor U4206 (N_4206,In_222,In_1125);
or U4207 (N_4207,In_2116,In_704);
nor U4208 (N_4208,In_744,In_1331);
nor U4209 (N_4209,In_2019,In_1407);
or U4210 (N_4210,In_1738,In_1079);
nor U4211 (N_4211,In_2232,In_1558);
xnor U4212 (N_4212,In_1102,In_1272);
and U4213 (N_4213,In_1628,In_2413);
or U4214 (N_4214,In_167,In_714);
and U4215 (N_4215,In_436,In_911);
or U4216 (N_4216,In_1354,In_660);
or U4217 (N_4217,In_2237,In_1983);
nor U4218 (N_4218,In_2205,In_1125);
and U4219 (N_4219,In_1524,In_1963);
xnor U4220 (N_4220,In_1274,In_1296);
and U4221 (N_4221,In_505,In_456);
nand U4222 (N_4222,In_950,In_2410);
nand U4223 (N_4223,In_652,In_1264);
and U4224 (N_4224,In_2034,In_773);
nand U4225 (N_4225,In_92,In_769);
and U4226 (N_4226,In_677,In_1095);
nor U4227 (N_4227,In_508,In_60);
nand U4228 (N_4228,In_234,In_1625);
or U4229 (N_4229,In_2424,In_2378);
and U4230 (N_4230,In_1686,In_1983);
xor U4231 (N_4231,In_2148,In_2393);
and U4232 (N_4232,In_357,In_2167);
xnor U4233 (N_4233,In_1672,In_1747);
or U4234 (N_4234,In_1069,In_496);
or U4235 (N_4235,In_239,In_1367);
and U4236 (N_4236,In_1075,In_913);
or U4237 (N_4237,In_1487,In_1528);
xnor U4238 (N_4238,In_2089,In_406);
nor U4239 (N_4239,In_55,In_19);
nor U4240 (N_4240,In_1385,In_1261);
nor U4241 (N_4241,In_2007,In_447);
nor U4242 (N_4242,In_15,In_802);
or U4243 (N_4243,In_2137,In_1559);
nor U4244 (N_4244,In_373,In_2152);
nand U4245 (N_4245,In_669,In_490);
and U4246 (N_4246,In_1447,In_1604);
or U4247 (N_4247,In_995,In_1717);
nor U4248 (N_4248,In_243,In_513);
xnor U4249 (N_4249,In_691,In_1460);
xor U4250 (N_4250,In_410,In_911);
and U4251 (N_4251,In_580,In_705);
nand U4252 (N_4252,In_779,In_984);
or U4253 (N_4253,In_685,In_453);
or U4254 (N_4254,In_137,In_2452);
and U4255 (N_4255,In_1744,In_2227);
nand U4256 (N_4256,In_524,In_1100);
nor U4257 (N_4257,In_2242,In_53);
nand U4258 (N_4258,In_930,In_2464);
nand U4259 (N_4259,In_1603,In_211);
nor U4260 (N_4260,In_968,In_2430);
xnor U4261 (N_4261,In_1579,In_1870);
or U4262 (N_4262,In_10,In_2286);
xnor U4263 (N_4263,In_245,In_1968);
xor U4264 (N_4264,In_1531,In_1384);
and U4265 (N_4265,In_1487,In_1729);
nor U4266 (N_4266,In_2441,In_63);
xor U4267 (N_4267,In_2436,In_2292);
nor U4268 (N_4268,In_165,In_174);
and U4269 (N_4269,In_1240,In_324);
xor U4270 (N_4270,In_2130,In_1225);
nor U4271 (N_4271,In_198,In_2373);
xnor U4272 (N_4272,In_781,In_2417);
xor U4273 (N_4273,In_883,In_1161);
nor U4274 (N_4274,In_740,In_542);
or U4275 (N_4275,In_2437,In_2214);
and U4276 (N_4276,In_1612,In_581);
nand U4277 (N_4277,In_1630,In_549);
or U4278 (N_4278,In_593,In_1277);
nor U4279 (N_4279,In_363,In_1601);
nor U4280 (N_4280,In_1739,In_1350);
and U4281 (N_4281,In_43,In_363);
nand U4282 (N_4282,In_614,In_1614);
or U4283 (N_4283,In_2128,In_198);
xnor U4284 (N_4284,In_1549,In_261);
or U4285 (N_4285,In_2023,In_2088);
xnor U4286 (N_4286,In_1170,In_1927);
nor U4287 (N_4287,In_2351,In_2079);
nor U4288 (N_4288,In_1208,In_2255);
xor U4289 (N_4289,In_605,In_2053);
and U4290 (N_4290,In_516,In_195);
or U4291 (N_4291,In_137,In_770);
or U4292 (N_4292,In_711,In_401);
and U4293 (N_4293,In_602,In_1624);
xnor U4294 (N_4294,In_78,In_2295);
and U4295 (N_4295,In_163,In_530);
and U4296 (N_4296,In_2337,In_1423);
or U4297 (N_4297,In_1205,In_1023);
nor U4298 (N_4298,In_1384,In_1243);
nor U4299 (N_4299,In_709,In_765);
nand U4300 (N_4300,In_1402,In_1725);
and U4301 (N_4301,In_892,In_459);
or U4302 (N_4302,In_585,In_671);
and U4303 (N_4303,In_138,In_1401);
or U4304 (N_4304,In_1963,In_1288);
nand U4305 (N_4305,In_2315,In_1055);
nand U4306 (N_4306,In_1296,In_1154);
nor U4307 (N_4307,In_217,In_878);
xor U4308 (N_4308,In_1430,In_2449);
xnor U4309 (N_4309,In_2056,In_654);
or U4310 (N_4310,In_2470,In_369);
and U4311 (N_4311,In_1344,In_1721);
xor U4312 (N_4312,In_1734,In_1768);
nand U4313 (N_4313,In_1307,In_2004);
nor U4314 (N_4314,In_1459,In_775);
and U4315 (N_4315,In_140,In_2316);
xnor U4316 (N_4316,In_2239,In_210);
nand U4317 (N_4317,In_1508,In_1121);
or U4318 (N_4318,In_645,In_2045);
or U4319 (N_4319,In_2222,In_541);
and U4320 (N_4320,In_329,In_1938);
xor U4321 (N_4321,In_1159,In_421);
and U4322 (N_4322,In_804,In_2012);
nor U4323 (N_4323,In_692,In_1033);
xnor U4324 (N_4324,In_1631,In_1272);
nand U4325 (N_4325,In_2190,In_1152);
xor U4326 (N_4326,In_1798,In_243);
nor U4327 (N_4327,In_2022,In_650);
nor U4328 (N_4328,In_681,In_695);
nor U4329 (N_4329,In_1200,In_2131);
nor U4330 (N_4330,In_1325,In_2122);
nor U4331 (N_4331,In_2444,In_1847);
nand U4332 (N_4332,In_83,In_2161);
nand U4333 (N_4333,In_1047,In_1816);
or U4334 (N_4334,In_1934,In_637);
or U4335 (N_4335,In_1508,In_1585);
xnor U4336 (N_4336,In_2231,In_818);
nand U4337 (N_4337,In_487,In_1091);
nor U4338 (N_4338,In_74,In_2157);
nand U4339 (N_4339,In_1185,In_1323);
nand U4340 (N_4340,In_1556,In_571);
nand U4341 (N_4341,In_927,In_1370);
xor U4342 (N_4342,In_1443,In_1924);
nor U4343 (N_4343,In_1528,In_1876);
or U4344 (N_4344,In_2050,In_574);
xnor U4345 (N_4345,In_1486,In_366);
nor U4346 (N_4346,In_1208,In_955);
xnor U4347 (N_4347,In_36,In_829);
xnor U4348 (N_4348,In_2446,In_249);
and U4349 (N_4349,In_2228,In_322);
or U4350 (N_4350,In_1172,In_1553);
xor U4351 (N_4351,In_706,In_1454);
and U4352 (N_4352,In_1633,In_1004);
or U4353 (N_4353,In_766,In_2272);
nor U4354 (N_4354,In_1930,In_973);
or U4355 (N_4355,In_1776,In_2096);
xnor U4356 (N_4356,In_890,In_537);
or U4357 (N_4357,In_1316,In_540);
nand U4358 (N_4358,In_60,In_2355);
nand U4359 (N_4359,In_657,In_703);
xor U4360 (N_4360,In_1914,In_1809);
or U4361 (N_4361,In_1184,In_1725);
nor U4362 (N_4362,In_1550,In_459);
nand U4363 (N_4363,In_1861,In_619);
xnor U4364 (N_4364,In_1714,In_259);
nor U4365 (N_4365,In_2022,In_203);
nand U4366 (N_4366,In_1245,In_640);
nor U4367 (N_4367,In_1716,In_2166);
nor U4368 (N_4368,In_570,In_903);
xor U4369 (N_4369,In_1944,In_795);
nor U4370 (N_4370,In_623,In_1554);
nor U4371 (N_4371,In_1443,In_252);
xnor U4372 (N_4372,In_1456,In_2193);
xor U4373 (N_4373,In_120,In_1703);
xnor U4374 (N_4374,In_625,In_1954);
nand U4375 (N_4375,In_1031,In_2158);
or U4376 (N_4376,In_256,In_2450);
and U4377 (N_4377,In_1800,In_2152);
nand U4378 (N_4378,In_1003,In_1);
or U4379 (N_4379,In_1627,In_1366);
nand U4380 (N_4380,In_567,In_631);
or U4381 (N_4381,In_301,In_1010);
or U4382 (N_4382,In_1212,In_166);
xnor U4383 (N_4383,In_2392,In_1663);
xor U4384 (N_4384,In_1529,In_1060);
xnor U4385 (N_4385,In_1700,In_493);
xor U4386 (N_4386,In_613,In_313);
nor U4387 (N_4387,In_692,In_2054);
and U4388 (N_4388,In_310,In_2238);
or U4389 (N_4389,In_33,In_1188);
xor U4390 (N_4390,In_417,In_2328);
nand U4391 (N_4391,In_450,In_1786);
xnor U4392 (N_4392,In_497,In_1280);
nor U4393 (N_4393,In_1613,In_1960);
nand U4394 (N_4394,In_1768,In_343);
xnor U4395 (N_4395,In_441,In_1331);
and U4396 (N_4396,In_1424,In_2270);
nor U4397 (N_4397,In_537,In_2394);
nand U4398 (N_4398,In_426,In_1546);
and U4399 (N_4399,In_2457,In_1203);
and U4400 (N_4400,In_1170,In_1661);
xnor U4401 (N_4401,In_568,In_949);
and U4402 (N_4402,In_2424,In_1974);
nand U4403 (N_4403,In_223,In_2235);
and U4404 (N_4404,In_166,In_357);
xnor U4405 (N_4405,In_1416,In_1404);
nor U4406 (N_4406,In_2388,In_932);
xnor U4407 (N_4407,In_1456,In_916);
nor U4408 (N_4408,In_1261,In_1415);
nand U4409 (N_4409,In_1778,In_742);
nor U4410 (N_4410,In_1027,In_699);
xor U4411 (N_4411,In_2354,In_301);
nand U4412 (N_4412,In_370,In_637);
nand U4413 (N_4413,In_1320,In_588);
and U4414 (N_4414,In_111,In_1792);
nand U4415 (N_4415,In_1289,In_1393);
or U4416 (N_4416,In_990,In_1928);
nand U4417 (N_4417,In_807,In_1797);
nand U4418 (N_4418,In_2419,In_1281);
nand U4419 (N_4419,In_1582,In_1448);
nor U4420 (N_4420,In_54,In_1475);
nor U4421 (N_4421,In_1064,In_965);
or U4422 (N_4422,In_783,In_411);
nand U4423 (N_4423,In_1860,In_488);
or U4424 (N_4424,In_1102,In_1836);
nor U4425 (N_4425,In_1828,In_1246);
nor U4426 (N_4426,In_904,In_2356);
xnor U4427 (N_4427,In_420,In_928);
and U4428 (N_4428,In_827,In_623);
nor U4429 (N_4429,In_1333,In_1220);
xnor U4430 (N_4430,In_718,In_1812);
xnor U4431 (N_4431,In_1455,In_830);
nor U4432 (N_4432,In_1378,In_1476);
nor U4433 (N_4433,In_385,In_660);
nand U4434 (N_4434,In_1567,In_378);
nand U4435 (N_4435,In_34,In_2046);
nand U4436 (N_4436,In_863,In_915);
nand U4437 (N_4437,In_520,In_744);
and U4438 (N_4438,In_1927,In_453);
nand U4439 (N_4439,In_424,In_909);
xnor U4440 (N_4440,In_1852,In_362);
nor U4441 (N_4441,In_671,In_251);
xor U4442 (N_4442,In_769,In_710);
or U4443 (N_4443,In_1981,In_431);
xor U4444 (N_4444,In_25,In_46);
xnor U4445 (N_4445,In_2106,In_1661);
nand U4446 (N_4446,In_607,In_470);
and U4447 (N_4447,In_1588,In_33);
or U4448 (N_4448,In_1924,In_495);
nor U4449 (N_4449,In_2412,In_61);
or U4450 (N_4450,In_980,In_927);
xnor U4451 (N_4451,In_2214,In_1749);
xor U4452 (N_4452,In_2257,In_506);
and U4453 (N_4453,In_1743,In_1277);
or U4454 (N_4454,In_720,In_301);
or U4455 (N_4455,In_1575,In_1831);
or U4456 (N_4456,In_671,In_187);
or U4457 (N_4457,In_1727,In_1642);
or U4458 (N_4458,In_1003,In_905);
nand U4459 (N_4459,In_2241,In_98);
nand U4460 (N_4460,In_850,In_1670);
xor U4461 (N_4461,In_197,In_2406);
or U4462 (N_4462,In_1349,In_1866);
xnor U4463 (N_4463,In_2180,In_2319);
nor U4464 (N_4464,In_2228,In_2411);
or U4465 (N_4465,In_2398,In_679);
and U4466 (N_4466,In_213,In_135);
and U4467 (N_4467,In_592,In_1125);
xnor U4468 (N_4468,In_892,In_642);
nor U4469 (N_4469,In_2326,In_2269);
or U4470 (N_4470,In_459,In_647);
or U4471 (N_4471,In_2401,In_396);
or U4472 (N_4472,In_1645,In_1952);
xnor U4473 (N_4473,In_2025,In_2423);
and U4474 (N_4474,In_1591,In_1610);
nor U4475 (N_4475,In_250,In_1411);
nor U4476 (N_4476,In_1480,In_2292);
and U4477 (N_4477,In_1771,In_1432);
or U4478 (N_4478,In_939,In_742);
and U4479 (N_4479,In_1795,In_18);
nor U4480 (N_4480,In_2006,In_1868);
nand U4481 (N_4481,In_1513,In_320);
xnor U4482 (N_4482,In_933,In_176);
and U4483 (N_4483,In_1390,In_822);
nand U4484 (N_4484,In_1275,In_817);
nand U4485 (N_4485,In_1931,In_1923);
and U4486 (N_4486,In_1538,In_71);
nor U4487 (N_4487,In_146,In_844);
nor U4488 (N_4488,In_269,In_860);
and U4489 (N_4489,In_826,In_674);
or U4490 (N_4490,In_125,In_1053);
nand U4491 (N_4491,In_593,In_584);
nand U4492 (N_4492,In_1545,In_1592);
nand U4493 (N_4493,In_1014,In_313);
and U4494 (N_4494,In_2161,In_1101);
xor U4495 (N_4495,In_1711,In_525);
xor U4496 (N_4496,In_1885,In_488);
nor U4497 (N_4497,In_908,In_874);
nor U4498 (N_4498,In_699,In_1130);
nand U4499 (N_4499,In_1145,In_2313);
and U4500 (N_4500,In_778,In_1002);
or U4501 (N_4501,In_2282,In_1981);
xor U4502 (N_4502,In_893,In_1384);
or U4503 (N_4503,In_572,In_1940);
and U4504 (N_4504,In_1260,In_2336);
xor U4505 (N_4505,In_1764,In_1017);
xor U4506 (N_4506,In_525,In_743);
nand U4507 (N_4507,In_415,In_668);
and U4508 (N_4508,In_1383,In_590);
nand U4509 (N_4509,In_1600,In_1280);
and U4510 (N_4510,In_1133,In_2017);
and U4511 (N_4511,In_1631,In_1352);
and U4512 (N_4512,In_1159,In_1735);
and U4513 (N_4513,In_1999,In_852);
nand U4514 (N_4514,In_204,In_47);
nor U4515 (N_4515,In_1925,In_573);
xor U4516 (N_4516,In_796,In_1878);
or U4517 (N_4517,In_1772,In_630);
or U4518 (N_4518,In_613,In_554);
xnor U4519 (N_4519,In_307,In_2467);
nand U4520 (N_4520,In_1562,In_1772);
or U4521 (N_4521,In_1069,In_2326);
nand U4522 (N_4522,In_1471,In_1978);
or U4523 (N_4523,In_2048,In_428);
and U4524 (N_4524,In_1457,In_218);
nor U4525 (N_4525,In_890,In_357);
and U4526 (N_4526,In_1373,In_19);
and U4527 (N_4527,In_1497,In_2221);
and U4528 (N_4528,In_686,In_1763);
nand U4529 (N_4529,In_1000,In_117);
and U4530 (N_4530,In_1541,In_1995);
and U4531 (N_4531,In_2179,In_1225);
and U4532 (N_4532,In_1491,In_1265);
nand U4533 (N_4533,In_1242,In_1225);
nand U4534 (N_4534,In_1580,In_1687);
xnor U4535 (N_4535,In_1409,In_2048);
nor U4536 (N_4536,In_2291,In_1057);
nand U4537 (N_4537,In_2238,In_2135);
or U4538 (N_4538,In_688,In_2321);
xor U4539 (N_4539,In_1615,In_903);
xor U4540 (N_4540,In_1905,In_2144);
and U4541 (N_4541,In_809,In_724);
xor U4542 (N_4542,In_1701,In_1549);
nand U4543 (N_4543,In_2317,In_138);
or U4544 (N_4544,In_1184,In_887);
nand U4545 (N_4545,In_931,In_1819);
or U4546 (N_4546,In_340,In_2089);
nor U4547 (N_4547,In_1306,In_1420);
nand U4548 (N_4548,In_1290,In_966);
xor U4549 (N_4549,In_2113,In_826);
and U4550 (N_4550,In_1909,In_2212);
nor U4551 (N_4551,In_2271,In_1675);
or U4552 (N_4552,In_1544,In_595);
nor U4553 (N_4553,In_242,In_758);
or U4554 (N_4554,In_374,In_861);
nand U4555 (N_4555,In_1211,In_646);
nor U4556 (N_4556,In_491,In_1672);
or U4557 (N_4557,In_401,In_1128);
xnor U4558 (N_4558,In_2101,In_533);
nor U4559 (N_4559,In_2200,In_1835);
or U4560 (N_4560,In_1510,In_1503);
nand U4561 (N_4561,In_1810,In_227);
nor U4562 (N_4562,In_2022,In_2095);
and U4563 (N_4563,In_360,In_1167);
and U4564 (N_4564,In_772,In_516);
or U4565 (N_4565,In_213,In_2096);
and U4566 (N_4566,In_280,In_1278);
nand U4567 (N_4567,In_957,In_367);
xnor U4568 (N_4568,In_747,In_1057);
nand U4569 (N_4569,In_1627,In_491);
and U4570 (N_4570,In_308,In_620);
or U4571 (N_4571,In_1397,In_1436);
nor U4572 (N_4572,In_167,In_1856);
nor U4573 (N_4573,In_1138,In_1377);
nand U4574 (N_4574,In_2397,In_1417);
and U4575 (N_4575,In_1561,In_97);
xor U4576 (N_4576,In_742,In_1705);
or U4577 (N_4577,In_36,In_1191);
or U4578 (N_4578,In_2482,In_1681);
nor U4579 (N_4579,In_61,In_385);
or U4580 (N_4580,In_690,In_2433);
or U4581 (N_4581,In_1990,In_1695);
nand U4582 (N_4582,In_1778,In_786);
xor U4583 (N_4583,In_1449,In_1805);
xor U4584 (N_4584,In_881,In_1387);
xnor U4585 (N_4585,In_56,In_907);
nand U4586 (N_4586,In_34,In_293);
nor U4587 (N_4587,In_1336,In_964);
and U4588 (N_4588,In_1143,In_521);
and U4589 (N_4589,In_1774,In_1593);
or U4590 (N_4590,In_1001,In_904);
nand U4591 (N_4591,In_37,In_2284);
nor U4592 (N_4592,In_2105,In_2089);
nand U4593 (N_4593,In_1663,In_380);
nor U4594 (N_4594,In_1719,In_185);
nand U4595 (N_4595,In_1259,In_1117);
nor U4596 (N_4596,In_1750,In_1535);
nor U4597 (N_4597,In_870,In_1111);
or U4598 (N_4598,In_200,In_2059);
nor U4599 (N_4599,In_2303,In_951);
or U4600 (N_4600,In_2447,In_1873);
xor U4601 (N_4601,In_883,In_55);
nand U4602 (N_4602,In_513,In_264);
nor U4603 (N_4603,In_1164,In_849);
xnor U4604 (N_4604,In_903,In_86);
and U4605 (N_4605,In_2374,In_251);
and U4606 (N_4606,In_174,In_1578);
xnor U4607 (N_4607,In_1640,In_2318);
xnor U4608 (N_4608,In_2303,In_1119);
xor U4609 (N_4609,In_1175,In_610);
and U4610 (N_4610,In_1982,In_1307);
or U4611 (N_4611,In_175,In_1565);
and U4612 (N_4612,In_327,In_1050);
nor U4613 (N_4613,In_1964,In_835);
and U4614 (N_4614,In_350,In_2341);
and U4615 (N_4615,In_1421,In_1273);
nor U4616 (N_4616,In_2494,In_2419);
and U4617 (N_4617,In_1689,In_769);
xnor U4618 (N_4618,In_631,In_1317);
xor U4619 (N_4619,In_55,In_196);
nor U4620 (N_4620,In_443,In_485);
nor U4621 (N_4621,In_1228,In_711);
and U4622 (N_4622,In_2370,In_1859);
and U4623 (N_4623,In_1621,In_1275);
and U4624 (N_4624,In_645,In_458);
and U4625 (N_4625,In_985,In_788);
nor U4626 (N_4626,In_260,In_1728);
nor U4627 (N_4627,In_2113,In_2287);
nand U4628 (N_4628,In_113,In_1613);
or U4629 (N_4629,In_1768,In_1316);
nor U4630 (N_4630,In_484,In_1341);
and U4631 (N_4631,In_1074,In_630);
xnor U4632 (N_4632,In_815,In_543);
xor U4633 (N_4633,In_1645,In_948);
nand U4634 (N_4634,In_1495,In_1672);
and U4635 (N_4635,In_194,In_1744);
and U4636 (N_4636,In_161,In_1309);
nand U4637 (N_4637,In_885,In_2463);
and U4638 (N_4638,In_1957,In_2111);
nor U4639 (N_4639,In_1391,In_14);
nand U4640 (N_4640,In_2093,In_430);
nand U4641 (N_4641,In_1878,In_372);
xor U4642 (N_4642,In_1854,In_143);
or U4643 (N_4643,In_1836,In_188);
or U4644 (N_4644,In_2479,In_1738);
nor U4645 (N_4645,In_204,In_846);
and U4646 (N_4646,In_1934,In_136);
or U4647 (N_4647,In_1951,In_1088);
and U4648 (N_4648,In_310,In_1547);
or U4649 (N_4649,In_356,In_806);
or U4650 (N_4650,In_1820,In_1419);
nand U4651 (N_4651,In_1903,In_930);
nor U4652 (N_4652,In_1205,In_1873);
nand U4653 (N_4653,In_1185,In_480);
or U4654 (N_4654,In_1457,In_2256);
nand U4655 (N_4655,In_1303,In_1400);
and U4656 (N_4656,In_1861,In_356);
nand U4657 (N_4657,In_2365,In_1802);
and U4658 (N_4658,In_1934,In_2191);
and U4659 (N_4659,In_195,In_897);
or U4660 (N_4660,In_1625,In_454);
and U4661 (N_4661,In_2026,In_122);
nor U4662 (N_4662,In_565,In_2266);
xor U4663 (N_4663,In_1871,In_2238);
and U4664 (N_4664,In_99,In_2132);
nand U4665 (N_4665,In_1942,In_2243);
and U4666 (N_4666,In_1015,In_233);
or U4667 (N_4667,In_2148,In_1667);
nor U4668 (N_4668,In_1279,In_570);
or U4669 (N_4669,In_853,In_732);
nor U4670 (N_4670,In_1673,In_808);
nand U4671 (N_4671,In_118,In_673);
nand U4672 (N_4672,In_2421,In_2286);
or U4673 (N_4673,In_543,In_1372);
or U4674 (N_4674,In_1381,In_1152);
nand U4675 (N_4675,In_205,In_2261);
nand U4676 (N_4676,In_629,In_999);
nor U4677 (N_4677,In_932,In_1303);
or U4678 (N_4678,In_1557,In_29);
xnor U4679 (N_4679,In_756,In_2245);
and U4680 (N_4680,In_1098,In_1116);
and U4681 (N_4681,In_337,In_1209);
nand U4682 (N_4682,In_383,In_1945);
and U4683 (N_4683,In_2133,In_2024);
and U4684 (N_4684,In_897,In_1682);
and U4685 (N_4685,In_655,In_1872);
or U4686 (N_4686,In_456,In_109);
or U4687 (N_4687,In_2021,In_1899);
xnor U4688 (N_4688,In_221,In_1929);
and U4689 (N_4689,In_979,In_2459);
and U4690 (N_4690,In_941,In_137);
nand U4691 (N_4691,In_1481,In_248);
or U4692 (N_4692,In_1049,In_999);
nor U4693 (N_4693,In_1732,In_404);
or U4694 (N_4694,In_138,In_2286);
or U4695 (N_4695,In_312,In_832);
or U4696 (N_4696,In_1572,In_2322);
nand U4697 (N_4697,In_2205,In_1769);
nand U4698 (N_4698,In_1793,In_1925);
nand U4699 (N_4699,In_1207,In_2272);
xor U4700 (N_4700,In_1431,In_1911);
and U4701 (N_4701,In_1483,In_145);
nor U4702 (N_4702,In_2373,In_1414);
nor U4703 (N_4703,In_1440,In_2084);
nor U4704 (N_4704,In_981,In_351);
or U4705 (N_4705,In_1265,In_1713);
nor U4706 (N_4706,In_218,In_1723);
and U4707 (N_4707,In_135,In_114);
xor U4708 (N_4708,In_1378,In_1253);
and U4709 (N_4709,In_1429,In_1788);
nand U4710 (N_4710,In_1122,In_2082);
or U4711 (N_4711,In_1799,In_2442);
and U4712 (N_4712,In_1722,In_325);
nor U4713 (N_4713,In_736,In_1401);
nand U4714 (N_4714,In_1833,In_1463);
and U4715 (N_4715,In_1287,In_1501);
nand U4716 (N_4716,In_464,In_1865);
nand U4717 (N_4717,In_107,In_325);
and U4718 (N_4718,In_1379,In_1694);
xor U4719 (N_4719,In_2051,In_2164);
nor U4720 (N_4720,In_1878,In_650);
and U4721 (N_4721,In_1411,In_1819);
and U4722 (N_4722,In_1667,In_302);
or U4723 (N_4723,In_557,In_402);
and U4724 (N_4724,In_2281,In_851);
nand U4725 (N_4725,In_185,In_1301);
and U4726 (N_4726,In_1438,In_1809);
nand U4727 (N_4727,In_920,In_606);
nand U4728 (N_4728,In_1699,In_2451);
or U4729 (N_4729,In_578,In_2315);
or U4730 (N_4730,In_2465,In_2227);
nand U4731 (N_4731,In_1135,In_1103);
nand U4732 (N_4732,In_812,In_64);
xor U4733 (N_4733,In_911,In_1727);
xor U4734 (N_4734,In_1807,In_1779);
nor U4735 (N_4735,In_890,In_137);
nor U4736 (N_4736,In_2217,In_2456);
nand U4737 (N_4737,In_1522,In_181);
and U4738 (N_4738,In_1513,In_235);
or U4739 (N_4739,In_976,In_1618);
nand U4740 (N_4740,In_1500,In_1647);
nor U4741 (N_4741,In_2402,In_1772);
nor U4742 (N_4742,In_1141,In_899);
nor U4743 (N_4743,In_2101,In_2267);
nand U4744 (N_4744,In_921,In_1961);
and U4745 (N_4745,In_1484,In_200);
and U4746 (N_4746,In_839,In_2477);
or U4747 (N_4747,In_2001,In_354);
and U4748 (N_4748,In_1262,In_5);
nand U4749 (N_4749,In_626,In_1772);
or U4750 (N_4750,In_1834,In_124);
or U4751 (N_4751,In_1005,In_2061);
and U4752 (N_4752,In_1739,In_1361);
and U4753 (N_4753,In_1662,In_530);
xor U4754 (N_4754,In_2013,In_98);
and U4755 (N_4755,In_1197,In_1072);
nor U4756 (N_4756,In_1473,In_1459);
and U4757 (N_4757,In_2007,In_1672);
or U4758 (N_4758,In_1041,In_1108);
and U4759 (N_4759,In_929,In_1753);
or U4760 (N_4760,In_1052,In_1955);
nor U4761 (N_4761,In_1476,In_989);
or U4762 (N_4762,In_963,In_1147);
and U4763 (N_4763,In_601,In_1729);
and U4764 (N_4764,In_51,In_955);
and U4765 (N_4765,In_2371,In_216);
nand U4766 (N_4766,In_2228,In_1461);
nor U4767 (N_4767,In_1587,In_873);
xnor U4768 (N_4768,In_1266,In_2115);
nor U4769 (N_4769,In_2278,In_2193);
xnor U4770 (N_4770,In_14,In_1498);
and U4771 (N_4771,In_1876,In_1692);
nor U4772 (N_4772,In_1766,In_2207);
xnor U4773 (N_4773,In_269,In_1721);
and U4774 (N_4774,In_979,In_823);
and U4775 (N_4775,In_1388,In_325);
nand U4776 (N_4776,In_1882,In_1096);
and U4777 (N_4777,In_698,In_575);
and U4778 (N_4778,In_2344,In_730);
nand U4779 (N_4779,In_807,In_745);
or U4780 (N_4780,In_958,In_1265);
or U4781 (N_4781,In_1742,In_1829);
xnor U4782 (N_4782,In_2317,In_87);
nand U4783 (N_4783,In_1448,In_960);
and U4784 (N_4784,In_1019,In_1974);
xnor U4785 (N_4785,In_2445,In_117);
and U4786 (N_4786,In_169,In_1917);
or U4787 (N_4787,In_2058,In_1586);
nand U4788 (N_4788,In_307,In_1438);
nor U4789 (N_4789,In_418,In_438);
nand U4790 (N_4790,In_892,In_2188);
and U4791 (N_4791,In_1403,In_1795);
or U4792 (N_4792,In_2018,In_716);
nand U4793 (N_4793,In_1589,In_2003);
nor U4794 (N_4794,In_1839,In_2284);
nand U4795 (N_4795,In_1120,In_191);
and U4796 (N_4796,In_534,In_1831);
nor U4797 (N_4797,In_1814,In_857);
and U4798 (N_4798,In_709,In_993);
or U4799 (N_4799,In_412,In_1261);
and U4800 (N_4800,In_309,In_391);
nor U4801 (N_4801,In_2164,In_2103);
and U4802 (N_4802,In_1727,In_2439);
or U4803 (N_4803,In_2375,In_2104);
nor U4804 (N_4804,In_685,In_972);
nor U4805 (N_4805,In_1388,In_2400);
nand U4806 (N_4806,In_626,In_2338);
and U4807 (N_4807,In_1440,In_1150);
or U4808 (N_4808,In_1657,In_1961);
or U4809 (N_4809,In_643,In_796);
or U4810 (N_4810,In_717,In_544);
nand U4811 (N_4811,In_1301,In_35);
or U4812 (N_4812,In_1199,In_1692);
and U4813 (N_4813,In_1867,In_1350);
nand U4814 (N_4814,In_1182,In_2404);
or U4815 (N_4815,In_483,In_2164);
nand U4816 (N_4816,In_867,In_1942);
nand U4817 (N_4817,In_222,In_2232);
nand U4818 (N_4818,In_728,In_2014);
nor U4819 (N_4819,In_497,In_1540);
nor U4820 (N_4820,In_1801,In_462);
or U4821 (N_4821,In_1955,In_1477);
xor U4822 (N_4822,In_856,In_1038);
xor U4823 (N_4823,In_1333,In_1164);
and U4824 (N_4824,In_28,In_1654);
and U4825 (N_4825,In_906,In_1302);
nand U4826 (N_4826,In_1646,In_1044);
xnor U4827 (N_4827,In_1957,In_654);
nand U4828 (N_4828,In_1601,In_118);
xnor U4829 (N_4829,In_1068,In_430);
or U4830 (N_4830,In_1904,In_144);
nor U4831 (N_4831,In_1443,In_1575);
or U4832 (N_4832,In_1503,In_996);
or U4833 (N_4833,In_517,In_873);
nand U4834 (N_4834,In_1990,In_643);
xnor U4835 (N_4835,In_1007,In_197);
nand U4836 (N_4836,In_1601,In_413);
nor U4837 (N_4837,In_1219,In_1048);
xor U4838 (N_4838,In_1094,In_1741);
or U4839 (N_4839,In_534,In_1873);
xor U4840 (N_4840,In_1358,In_1563);
nor U4841 (N_4841,In_1001,In_1510);
or U4842 (N_4842,In_48,In_445);
or U4843 (N_4843,In_1153,In_131);
nand U4844 (N_4844,In_2052,In_1532);
nor U4845 (N_4845,In_2170,In_1579);
and U4846 (N_4846,In_719,In_344);
nor U4847 (N_4847,In_206,In_1895);
xor U4848 (N_4848,In_2461,In_1547);
xnor U4849 (N_4849,In_1239,In_107);
or U4850 (N_4850,In_481,In_240);
nand U4851 (N_4851,In_1483,In_1153);
nor U4852 (N_4852,In_2066,In_2306);
and U4853 (N_4853,In_341,In_1381);
and U4854 (N_4854,In_795,In_2153);
or U4855 (N_4855,In_334,In_119);
or U4856 (N_4856,In_1456,In_1682);
xor U4857 (N_4857,In_1363,In_671);
nor U4858 (N_4858,In_265,In_1992);
and U4859 (N_4859,In_2374,In_1436);
xnor U4860 (N_4860,In_2491,In_2414);
xnor U4861 (N_4861,In_797,In_2007);
nand U4862 (N_4862,In_669,In_1688);
or U4863 (N_4863,In_1417,In_946);
nand U4864 (N_4864,In_2288,In_211);
nor U4865 (N_4865,In_352,In_229);
and U4866 (N_4866,In_1156,In_529);
nand U4867 (N_4867,In_2342,In_568);
and U4868 (N_4868,In_672,In_1449);
xor U4869 (N_4869,In_920,In_2498);
nand U4870 (N_4870,In_2104,In_1457);
nand U4871 (N_4871,In_490,In_146);
nand U4872 (N_4872,In_413,In_201);
or U4873 (N_4873,In_924,In_1304);
nor U4874 (N_4874,In_925,In_234);
and U4875 (N_4875,In_1709,In_880);
or U4876 (N_4876,In_480,In_401);
or U4877 (N_4877,In_1875,In_848);
nor U4878 (N_4878,In_844,In_401);
and U4879 (N_4879,In_1797,In_1069);
nor U4880 (N_4880,In_611,In_224);
and U4881 (N_4881,In_394,In_1134);
nor U4882 (N_4882,In_1020,In_1461);
xor U4883 (N_4883,In_428,In_1897);
nor U4884 (N_4884,In_2056,In_1713);
xor U4885 (N_4885,In_1477,In_1964);
xor U4886 (N_4886,In_86,In_851);
nor U4887 (N_4887,In_1238,In_1081);
nand U4888 (N_4888,In_1132,In_2320);
and U4889 (N_4889,In_1587,In_334);
nand U4890 (N_4890,In_955,In_2458);
xnor U4891 (N_4891,In_1358,In_2026);
xnor U4892 (N_4892,In_1935,In_2006);
xor U4893 (N_4893,In_1464,In_651);
and U4894 (N_4894,In_897,In_2029);
nor U4895 (N_4895,In_1970,In_155);
nand U4896 (N_4896,In_230,In_1239);
and U4897 (N_4897,In_1785,In_953);
and U4898 (N_4898,In_1314,In_498);
or U4899 (N_4899,In_2385,In_1729);
nor U4900 (N_4900,In_2364,In_1485);
or U4901 (N_4901,In_1671,In_149);
or U4902 (N_4902,In_2263,In_310);
or U4903 (N_4903,In_2450,In_1254);
and U4904 (N_4904,In_1234,In_1444);
and U4905 (N_4905,In_2233,In_1292);
xnor U4906 (N_4906,In_2374,In_1468);
and U4907 (N_4907,In_508,In_227);
nor U4908 (N_4908,In_1577,In_1752);
xor U4909 (N_4909,In_2045,In_673);
or U4910 (N_4910,In_1809,In_188);
or U4911 (N_4911,In_893,In_1518);
nor U4912 (N_4912,In_1860,In_1103);
or U4913 (N_4913,In_106,In_1602);
nor U4914 (N_4914,In_14,In_1357);
nor U4915 (N_4915,In_993,In_649);
nand U4916 (N_4916,In_1498,In_977);
or U4917 (N_4917,In_674,In_14);
and U4918 (N_4918,In_1374,In_1245);
xor U4919 (N_4919,In_1439,In_2339);
and U4920 (N_4920,In_1708,In_1502);
or U4921 (N_4921,In_2284,In_1944);
xor U4922 (N_4922,In_1718,In_2495);
nor U4923 (N_4923,In_498,In_1807);
nor U4924 (N_4924,In_2455,In_1673);
and U4925 (N_4925,In_21,In_175);
or U4926 (N_4926,In_738,In_1381);
xor U4927 (N_4927,In_428,In_2426);
nor U4928 (N_4928,In_1655,In_2060);
xor U4929 (N_4929,In_974,In_1010);
nand U4930 (N_4930,In_1920,In_306);
or U4931 (N_4931,In_1895,In_342);
nand U4932 (N_4932,In_530,In_2365);
and U4933 (N_4933,In_1649,In_2146);
xor U4934 (N_4934,In_877,In_2263);
xnor U4935 (N_4935,In_1133,In_1907);
nand U4936 (N_4936,In_611,In_305);
nor U4937 (N_4937,In_1404,In_1411);
xor U4938 (N_4938,In_90,In_647);
and U4939 (N_4939,In_1699,In_1782);
nand U4940 (N_4940,In_185,In_2118);
nor U4941 (N_4941,In_2211,In_368);
nor U4942 (N_4942,In_1029,In_319);
xnor U4943 (N_4943,In_590,In_1986);
and U4944 (N_4944,In_2299,In_858);
nor U4945 (N_4945,In_555,In_1300);
or U4946 (N_4946,In_1792,In_2358);
and U4947 (N_4947,In_2306,In_1977);
xor U4948 (N_4948,In_1559,In_800);
or U4949 (N_4949,In_967,In_1196);
and U4950 (N_4950,In_750,In_1711);
xnor U4951 (N_4951,In_1358,In_901);
nor U4952 (N_4952,In_1646,In_66);
nand U4953 (N_4953,In_1216,In_909);
or U4954 (N_4954,In_2207,In_482);
nor U4955 (N_4955,In_58,In_866);
nand U4956 (N_4956,In_2442,In_185);
nor U4957 (N_4957,In_201,In_736);
or U4958 (N_4958,In_838,In_363);
nor U4959 (N_4959,In_363,In_2328);
and U4960 (N_4960,In_922,In_84);
nor U4961 (N_4961,In_235,In_766);
nor U4962 (N_4962,In_1249,In_655);
nand U4963 (N_4963,In_1629,In_795);
and U4964 (N_4964,In_81,In_90);
and U4965 (N_4965,In_2292,In_1298);
xor U4966 (N_4966,In_317,In_1884);
nor U4967 (N_4967,In_499,In_1587);
and U4968 (N_4968,In_907,In_2417);
and U4969 (N_4969,In_875,In_2185);
and U4970 (N_4970,In_1357,In_1833);
xnor U4971 (N_4971,In_2016,In_1455);
and U4972 (N_4972,In_1698,In_235);
nand U4973 (N_4973,In_893,In_959);
nand U4974 (N_4974,In_1352,In_1570);
nand U4975 (N_4975,In_1368,In_794);
or U4976 (N_4976,In_2032,In_1789);
and U4977 (N_4977,In_2395,In_2247);
nor U4978 (N_4978,In_1201,In_481);
nor U4979 (N_4979,In_1750,In_900);
nor U4980 (N_4980,In_2144,In_1993);
or U4981 (N_4981,In_60,In_2475);
xor U4982 (N_4982,In_2497,In_1257);
xnor U4983 (N_4983,In_1230,In_10);
xor U4984 (N_4984,In_818,In_684);
xnor U4985 (N_4985,In_1208,In_498);
xnor U4986 (N_4986,In_545,In_810);
nor U4987 (N_4987,In_1082,In_189);
and U4988 (N_4988,In_951,In_1849);
nand U4989 (N_4989,In_2048,In_2232);
nor U4990 (N_4990,In_813,In_2285);
and U4991 (N_4991,In_498,In_602);
nor U4992 (N_4992,In_1219,In_1253);
and U4993 (N_4993,In_2437,In_1755);
xor U4994 (N_4994,In_610,In_174);
nand U4995 (N_4995,In_1075,In_1951);
xor U4996 (N_4996,In_546,In_1734);
xnor U4997 (N_4997,In_1552,In_2070);
nand U4998 (N_4998,In_271,In_689);
xnor U4999 (N_4999,In_1090,In_1086);
or U5000 (N_5000,In_2481,In_181);
xor U5001 (N_5001,In_1279,In_1437);
nor U5002 (N_5002,In_1137,In_1982);
or U5003 (N_5003,In_1902,In_1646);
nand U5004 (N_5004,In_1141,In_1906);
nor U5005 (N_5005,In_223,In_1900);
and U5006 (N_5006,In_58,In_1964);
or U5007 (N_5007,In_1985,In_188);
and U5008 (N_5008,In_2450,In_504);
or U5009 (N_5009,In_2413,In_2188);
or U5010 (N_5010,In_1571,In_167);
and U5011 (N_5011,In_573,In_2232);
nor U5012 (N_5012,In_1627,In_814);
nor U5013 (N_5013,In_1989,In_892);
and U5014 (N_5014,In_17,In_744);
or U5015 (N_5015,In_134,In_1184);
xor U5016 (N_5016,In_1225,In_1356);
nor U5017 (N_5017,In_997,In_1279);
nand U5018 (N_5018,In_1329,In_606);
nand U5019 (N_5019,In_502,In_1794);
xor U5020 (N_5020,In_1617,In_616);
and U5021 (N_5021,In_1926,In_1302);
xnor U5022 (N_5022,In_925,In_2428);
or U5023 (N_5023,In_606,In_651);
or U5024 (N_5024,In_22,In_288);
and U5025 (N_5025,In_1352,In_1943);
and U5026 (N_5026,In_1647,In_599);
nand U5027 (N_5027,In_2205,In_379);
xor U5028 (N_5028,In_946,In_2099);
nand U5029 (N_5029,In_1225,In_944);
xnor U5030 (N_5030,In_1436,In_1021);
or U5031 (N_5031,In_1263,In_559);
xnor U5032 (N_5032,In_305,In_2107);
and U5033 (N_5033,In_2420,In_466);
xor U5034 (N_5034,In_1032,In_187);
and U5035 (N_5035,In_2052,In_2292);
or U5036 (N_5036,In_41,In_476);
or U5037 (N_5037,In_2349,In_7);
nor U5038 (N_5038,In_1039,In_1755);
and U5039 (N_5039,In_1008,In_372);
xor U5040 (N_5040,In_556,In_440);
and U5041 (N_5041,In_1606,In_808);
or U5042 (N_5042,In_1396,In_1678);
nor U5043 (N_5043,In_2454,In_2124);
xor U5044 (N_5044,In_711,In_1679);
nor U5045 (N_5045,In_298,In_348);
and U5046 (N_5046,In_958,In_432);
or U5047 (N_5047,In_1371,In_321);
or U5048 (N_5048,In_274,In_2302);
or U5049 (N_5049,In_358,In_1624);
and U5050 (N_5050,In_218,In_1334);
nor U5051 (N_5051,In_1188,In_607);
nor U5052 (N_5052,In_1089,In_764);
or U5053 (N_5053,In_1454,In_2336);
or U5054 (N_5054,In_2097,In_1589);
nor U5055 (N_5055,In_1672,In_1528);
or U5056 (N_5056,In_2268,In_768);
xnor U5057 (N_5057,In_872,In_618);
or U5058 (N_5058,In_2236,In_835);
and U5059 (N_5059,In_1653,In_310);
or U5060 (N_5060,In_2093,In_2130);
nand U5061 (N_5061,In_2249,In_891);
nand U5062 (N_5062,In_2328,In_1213);
and U5063 (N_5063,In_1868,In_2090);
nor U5064 (N_5064,In_1945,In_913);
and U5065 (N_5065,In_503,In_1818);
xor U5066 (N_5066,In_1858,In_1404);
nor U5067 (N_5067,In_777,In_1516);
nand U5068 (N_5068,In_2161,In_2444);
nand U5069 (N_5069,In_148,In_1579);
nor U5070 (N_5070,In_1455,In_280);
and U5071 (N_5071,In_2450,In_2314);
xor U5072 (N_5072,In_1171,In_2147);
or U5073 (N_5073,In_991,In_1374);
nor U5074 (N_5074,In_1629,In_1754);
nor U5075 (N_5075,In_2371,In_275);
and U5076 (N_5076,In_115,In_1683);
and U5077 (N_5077,In_2469,In_976);
or U5078 (N_5078,In_700,In_914);
nor U5079 (N_5079,In_1310,In_728);
and U5080 (N_5080,In_1310,In_2079);
xnor U5081 (N_5081,In_153,In_456);
xnor U5082 (N_5082,In_755,In_53);
xor U5083 (N_5083,In_2422,In_1004);
xor U5084 (N_5084,In_1205,In_1401);
and U5085 (N_5085,In_2154,In_187);
xor U5086 (N_5086,In_315,In_1185);
nand U5087 (N_5087,In_1778,In_392);
and U5088 (N_5088,In_1494,In_367);
or U5089 (N_5089,In_890,In_315);
xor U5090 (N_5090,In_633,In_122);
or U5091 (N_5091,In_686,In_2022);
nor U5092 (N_5092,In_1440,In_43);
xnor U5093 (N_5093,In_1778,In_1401);
nand U5094 (N_5094,In_1443,In_1303);
or U5095 (N_5095,In_2317,In_76);
nand U5096 (N_5096,In_161,In_1332);
nor U5097 (N_5097,In_178,In_1820);
nand U5098 (N_5098,In_1987,In_1842);
and U5099 (N_5099,In_2255,In_2380);
and U5100 (N_5100,In_835,In_1825);
and U5101 (N_5101,In_452,In_1777);
or U5102 (N_5102,In_1391,In_1437);
nand U5103 (N_5103,In_2319,In_1522);
nor U5104 (N_5104,In_174,In_717);
xnor U5105 (N_5105,In_1382,In_2349);
nor U5106 (N_5106,In_907,In_1194);
xnor U5107 (N_5107,In_242,In_2005);
nand U5108 (N_5108,In_1551,In_1086);
xor U5109 (N_5109,In_578,In_614);
xor U5110 (N_5110,In_1882,In_2098);
nand U5111 (N_5111,In_227,In_1737);
xnor U5112 (N_5112,In_756,In_1057);
and U5113 (N_5113,In_1793,In_1563);
nand U5114 (N_5114,In_493,In_356);
nand U5115 (N_5115,In_1763,In_36);
or U5116 (N_5116,In_1515,In_561);
or U5117 (N_5117,In_1783,In_1722);
xor U5118 (N_5118,In_660,In_1806);
or U5119 (N_5119,In_1597,In_684);
nor U5120 (N_5120,In_2056,In_206);
or U5121 (N_5121,In_1144,In_2127);
and U5122 (N_5122,In_1314,In_281);
or U5123 (N_5123,In_318,In_320);
xor U5124 (N_5124,In_1106,In_1181);
nor U5125 (N_5125,In_1462,In_790);
and U5126 (N_5126,In_2050,In_1494);
nand U5127 (N_5127,In_1296,In_2195);
or U5128 (N_5128,In_2162,In_306);
xor U5129 (N_5129,In_2166,In_2270);
and U5130 (N_5130,In_1835,In_878);
nor U5131 (N_5131,In_812,In_1251);
and U5132 (N_5132,In_505,In_2367);
nor U5133 (N_5133,In_2101,In_1364);
and U5134 (N_5134,In_1732,In_2337);
nor U5135 (N_5135,In_1995,In_526);
xnor U5136 (N_5136,In_8,In_2491);
and U5137 (N_5137,In_1630,In_1521);
nor U5138 (N_5138,In_584,In_663);
nor U5139 (N_5139,In_2209,In_1414);
or U5140 (N_5140,In_622,In_2477);
nor U5141 (N_5141,In_1387,In_87);
xnor U5142 (N_5142,In_2454,In_629);
nand U5143 (N_5143,In_1752,In_624);
nand U5144 (N_5144,In_1748,In_1426);
nand U5145 (N_5145,In_1565,In_436);
nand U5146 (N_5146,In_304,In_1275);
xnor U5147 (N_5147,In_2359,In_2490);
or U5148 (N_5148,In_8,In_1019);
nor U5149 (N_5149,In_256,In_1558);
nand U5150 (N_5150,In_1634,In_2059);
and U5151 (N_5151,In_2202,In_458);
and U5152 (N_5152,In_237,In_138);
xnor U5153 (N_5153,In_1743,In_776);
nor U5154 (N_5154,In_216,In_295);
xnor U5155 (N_5155,In_1996,In_2122);
xnor U5156 (N_5156,In_778,In_1992);
xnor U5157 (N_5157,In_2220,In_361);
and U5158 (N_5158,In_44,In_1202);
or U5159 (N_5159,In_810,In_2379);
or U5160 (N_5160,In_331,In_838);
xor U5161 (N_5161,In_402,In_317);
nand U5162 (N_5162,In_1258,In_1604);
and U5163 (N_5163,In_1665,In_1069);
nor U5164 (N_5164,In_259,In_1349);
and U5165 (N_5165,In_1018,In_1191);
xnor U5166 (N_5166,In_529,In_2472);
and U5167 (N_5167,In_609,In_1982);
and U5168 (N_5168,In_2488,In_1162);
xor U5169 (N_5169,In_650,In_325);
xor U5170 (N_5170,In_148,In_361);
or U5171 (N_5171,In_2319,In_1091);
and U5172 (N_5172,In_2218,In_1960);
and U5173 (N_5173,In_1854,In_99);
nand U5174 (N_5174,In_814,In_2148);
and U5175 (N_5175,In_1186,In_346);
or U5176 (N_5176,In_1449,In_448);
nand U5177 (N_5177,In_500,In_362);
xnor U5178 (N_5178,In_1937,In_879);
nand U5179 (N_5179,In_1809,In_1599);
nor U5180 (N_5180,In_2355,In_2462);
or U5181 (N_5181,In_2490,In_1933);
or U5182 (N_5182,In_744,In_2407);
and U5183 (N_5183,In_876,In_1182);
xor U5184 (N_5184,In_195,In_306);
and U5185 (N_5185,In_211,In_1018);
xnor U5186 (N_5186,In_59,In_2472);
xnor U5187 (N_5187,In_258,In_344);
xor U5188 (N_5188,In_2280,In_593);
xor U5189 (N_5189,In_1106,In_883);
nand U5190 (N_5190,In_681,In_819);
nor U5191 (N_5191,In_505,In_809);
nor U5192 (N_5192,In_366,In_313);
nor U5193 (N_5193,In_135,In_2373);
nor U5194 (N_5194,In_538,In_1284);
nand U5195 (N_5195,In_1616,In_1214);
and U5196 (N_5196,In_1850,In_2344);
xnor U5197 (N_5197,In_890,In_1853);
nor U5198 (N_5198,In_1010,In_788);
and U5199 (N_5199,In_2406,In_363);
and U5200 (N_5200,In_1656,In_655);
or U5201 (N_5201,In_643,In_2124);
and U5202 (N_5202,In_1291,In_2493);
nand U5203 (N_5203,In_1291,In_1833);
and U5204 (N_5204,In_2371,In_2168);
xor U5205 (N_5205,In_18,In_2188);
nor U5206 (N_5206,In_861,In_1354);
and U5207 (N_5207,In_1739,In_1189);
xnor U5208 (N_5208,In_1656,In_746);
and U5209 (N_5209,In_1450,In_2451);
nand U5210 (N_5210,In_1651,In_358);
nand U5211 (N_5211,In_2391,In_1302);
and U5212 (N_5212,In_784,In_2320);
xor U5213 (N_5213,In_2366,In_1646);
and U5214 (N_5214,In_703,In_2174);
nand U5215 (N_5215,In_357,In_2485);
nand U5216 (N_5216,In_767,In_1492);
nor U5217 (N_5217,In_2430,In_2357);
nand U5218 (N_5218,In_1602,In_2055);
xnor U5219 (N_5219,In_1765,In_1133);
nand U5220 (N_5220,In_1833,In_1105);
nand U5221 (N_5221,In_773,In_2461);
xor U5222 (N_5222,In_1258,In_2225);
nand U5223 (N_5223,In_2167,In_1318);
or U5224 (N_5224,In_2062,In_650);
nand U5225 (N_5225,In_294,In_46);
nand U5226 (N_5226,In_1795,In_1196);
nand U5227 (N_5227,In_2023,In_2157);
and U5228 (N_5228,In_353,In_845);
nand U5229 (N_5229,In_2094,In_2318);
and U5230 (N_5230,In_358,In_700);
or U5231 (N_5231,In_1253,In_1740);
nor U5232 (N_5232,In_2166,In_1085);
nor U5233 (N_5233,In_1179,In_1766);
or U5234 (N_5234,In_2365,In_586);
nand U5235 (N_5235,In_1783,In_508);
nand U5236 (N_5236,In_380,In_1363);
xor U5237 (N_5237,In_1714,In_393);
and U5238 (N_5238,In_1073,In_738);
or U5239 (N_5239,In_701,In_330);
nor U5240 (N_5240,In_1304,In_1572);
xor U5241 (N_5241,In_1478,In_576);
or U5242 (N_5242,In_310,In_66);
nor U5243 (N_5243,In_1842,In_847);
nor U5244 (N_5244,In_1789,In_1941);
or U5245 (N_5245,In_868,In_1128);
and U5246 (N_5246,In_607,In_2351);
nand U5247 (N_5247,In_378,In_1884);
nor U5248 (N_5248,In_942,In_2325);
or U5249 (N_5249,In_2001,In_2162);
nand U5250 (N_5250,In_504,In_333);
xnor U5251 (N_5251,In_1811,In_965);
or U5252 (N_5252,In_516,In_1703);
nor U5253 (N_5253,In_1500,In_676);
and U5254 (N_5254,In_928,In_872);
nor U5255 (N_5255,In_1000,In_865);
nand U5256 (N_5256,In_2009,In_1486);
nand U5257 (N_5257,In_1839,In_139);
or U5258 (N_5258,In_598,In_405);
and U5259 (N_5259,In_523,In_1088);
nand U5260 (N_5260,In_82,In_2221);
xor U5261 (N_5261,In_436,In_349);
nor U5262 (N_5262,In_1507,In_1901);
nand U5263 (N_5263,In_1649,In_2419);
or U5264 (N_5264,In_2195,In_1724);
xor U5265 (N_5265,In_674,In_1784);
xnor U5266 (N_5266,In_640,In_1708);
nor U5267 (N_5267,In_2339,In_883);
xnor U5268 (N_5268,In_1029,In_1680);
or U5269 (N_5269,In_1257,In_1968);
and U5270 (N_5270,In_384,In_472);
and U5271 (N_5271,In_463,In_1910);
or U5272 (N_5272,In_2255,In_540);
and U5273 (N_5273,In_63,In_1527);
nand U5274 (N_5274,In_1517,In_1074);
nor U5275 (N_5275,In_199,In_1004);
nor U5276 (N_5276,In_1053,In_1618);
and U5277 (N_5277,In_620,In_834);
xor U5278 (N_5278,In_2056,In_2023);
or U5279 (N_5279,In_55,In_836);
nand U5280 (N_5280,In_823,In_2403);
nand U5281 (N_5281,In_1166,In_1313);
nor U5282 (N_5282,In_695,In_591);
or U5283 (N_5283,In_1066,In_2083);
nor U5284 (N_5284,In_1890,In_692);
or U5285 (N_5285,In_2020,In_2427);
xnor U5286 (N_5286,In_527,In_1275);
or U5287 (N_5287,In_2039,In_2396);
and U5288 (N_5288,In_1772,In_2308);
xor U5289 (N_5289,In_1179,In_627);
nand U5290 (N_5290,In_1140,In_724);
or U5291 (N_5291,In_1634,In_1827);
nand U5292 (N_5292,In_1668,In_598);
xor U5293 (N_5293,In_1285,In_1184);
or U5294 (N_5294,In_1791,In_1649);
nor U5295 (N_5295,In_178,In_533);
nor U5296 (N_5296,In_745,In_101);
nor U5297 (N_5297,In_895,In_2261);
xnor U5298 (N_5298,In_1260,In_1351);
and U5299 (N_5299,In_1384,In_2044);
and U5300 (N_5300,In_2453,In_1730);
nor U5301 (N_5301,In_1207,In_299);
and U5302 (N_5302,In_1823,In_1523);
nor U5303 (N_5303,In_1791,In_1966);
or U5304 (N_5304,In_1085,In_999);
and U5305 (N_5305,In_634,In_151);
nor U5306 (N_5306,In_609,In_1091);
or U5307 (N_5307,In_1029,In_1554);
nand U5308 (N_5308,In_1547,In_2242);
and U5309 (N_5309,In_177,In_767);
and U5310 (N_5310,In_1297,In_1222);
and U5311 (N_5311,In_1504,In_1836);
nor U5312 (N_5312,In_1097,In_1051);
xnor U5313 (N_5313,In_1415,In_2431);
and U5314 (N_5314,In_2046,In_2357);
xnor U5315 (N_5315,In_105,In_1912);
xnor U5316 (N_5316,In_1364,In_750);
xor U5317 (N_5317,In_670,In_913);
or U5318 (N_5318,In_896,In_803);
or U5319 (N_5319,In_2433,In_1805);
xor U5320 (N_5320,In_488,In_2233);
nand U5321 (N_5321,In_1147,In_539);
nand U5322 (N_5322,In_1641,In_2188);
or U5323 (N_5323,In_1835,In_1884);
xor U5324 (N_5324,In_1785,In_1156);
and U5325 (N_5325,In_1134,In_874);
nand U5326 (N_5326,In_1782,In_395);
nor U5327 (N_5327,In_1250,In_1215);
xnor U5328 (N_5328,In_2474,In_2048);
nand U5329 (N_5329,In_559,In_1218);
xnor U5330 (N_5330,In_2384,In_347);
nand U5331 (N_5331,In_2152,In_1913);
nor U5332 (N_5332,In_2104,In_879);
nor U5333 (N_5333,In_1891,In_134);
nor U5334 (N_5334,In_760,In_2107);
or U5335 (N_5335,In_2381,In_1733);
nand U5336 (N_5336,In_331,In_633);
nand U5337 (N_5337,In_1466,In_83);
xor U5338 (N_5338,In_1841,In_293);
nand U5339 (N_5339,In_51,In_109);
and U5340 (N_5340,In_278,In_1424);
or U5341 (N_5341,In_1924,In_2190);
and U5342 (N_5342,In_777,In_1042);
nor U5343 (N_5343,In_2242,In_1943);
and U5344 (N_5344,In_74,In_2257);
and U5345 (N_5345,In_1245,In_1929);
nand U5346 (N_5346,In_1989,In_1203);
or U5347 (N_5347,In_862,In_361);
nand U5348 (N_5348,In_1199,In_1608);
nand U5349 (N_5349,In_1121,In_1365);
or U5350 (N_5350,In_1199,In_1878);
nand U5351 (N_5351,In_1545,In_2328);
and U5352 (N_5352,In_1829,In_2182);
nand U5353 (N_5353,In_1879,In_7);
nand U5354 (N_5354,In_1513,In_1183);
and U5355 (N_5355,In_1011,In_1436);
nand U5356 (N_5356,In_430,In_2226);
and U5357 (N_5357,In_1365,In_366);
or U5358 (N_5358,In_1937,In_1618);
nor U5359 (N_5359,In_504,In_2236);
xnor U5360 (N_5360,In_1980,In_1263);
nand U5361 (N_5361,In_147,In_578);
nor U5362 (N_5362,In_1445,In_1273);
nand U5363 (N_5363,In_237,In_1530);
or U5364 (N_5364,In_2005,In_2168);
xor U5365 (N_5365,In_1716,In_2491);
and U5366 (N_5366,In_104,In_2405);
or U5367 (N_5367,In_1140,In_1450);
or U5368 (N_5368,In_1605,In_52);
and U5369 (N_5369,In_862,In_1658);
nand U5370 (N_5370,In_2109,In_547);
xnor U5371 (N_5371,In_713,In_1396);
or U5372 (N_5372,In_360,In_2003);
nor U5373 (N_5373,In_31,In_2251);
or U5374 (N_5374,In_1421,In_161);
and U5375 (N_5375,In_1743,In_1086);
or U5376 (N_5376,In_1079,In_712);
nor U5377 (N_5377,In_1497,In_1512);
nor U5378 (N_5378,In_78,In_1123);
nor U5379 (N_5379,In_747,In_2003);
and U5380 (N_5380,In_909,In_401);
nor U5381 (N_5381,In_615,In_953);
xnor U5382 (N_5382,In_2155,In_1320);
xor U5383 (N_5383,In_1399,In_1865);
nand U5384 (N_5384,In_1046,In_1828);
and U5385 (N_5385,In_2291,In_695);
xor U5386 (N_5386,In_1924,In_2041);
or U5387 (N_5387,In_1518,In_534);
or U5388 (N_5388,In_715,In_1992);
or U5389 (N_5389,In_188,In_2148);
xnor U5390 (N_5390,In_74,In_1056);
nor U5391 (N_5391,In_990,In_450);
or U5392 (N_5392,In_2016,In_947);
nand U5393 (N_5393,In_671,In_1393);
nor U5394 (N_5394,In_2196,In_971);
nand U5395 (N_5395,In_49,In_1956);
or U5396 (N_5396,In_2227,In_224);
xor U5397 (N_5397,In_76,In_2450);
nand U5398 (N_5398,In_2004,In_1278);
nand U5399 (N_5399,In_1622,In_1158);
and U5400 (N_5400,In_2154,In_1203);
or U5401 (N_5401,In_2095,In_424);
xnor U5402 (N_5402,In_1174,In_783);
xor U5403 (N_5403,In_2019,In_57);
or U5404 (N_5404,In_1719,In_115);
and U5405 (N_5405,In_564,In_2119);
xor U5406 (N_5406,In_1293,In_796);
or U5407 (N_5407,In_2305,In_2304);
xor U5408 (N_5408,In_1830,In_44);
or U5409 (N_5409,In_1424,In_1142);
xor U5410 (N_5410,In_2456,In_1935);
nand U5411 (N_5411,In_1691,In_1025);
xnor U5412 (N_5412,In_1121,In_2120);
nand U5413 (N_5413,In_2081,In_2466);
nand U5414 (N_5414,In_843,In_1069);
or U5415 (N_5415,In_1549,In_1089);
nand U5416 (N_5416,In_664,In_67);
and U5417 (N_5417,In_2240,In_290);
and U5418 (N_5418,In_1009,In_1717);
and U5419 (N_5419,In_1164,In_191);
nor U5420 (N_5420,In_807,In_747);
xor U5421 (N_5421,In_100,In_1451);
and U5422 (N_5422,In_345,In_2421);
and U5423 (N_5423,In_779,In_530);
xor U5424 (N_5424,In_1754,In_1648);
and U5425 (N_5425,In_2164,In_2236);
xnor U5426 (N_5426,In_159,In_1028);
nor U5427 (N_5427,In_1326,In_1535);
nor U5428 (N_5428,In_2063,In_2242);
or U5429 (N_5429,In_2451,In_525);
xnor U5430 (N_5430,In_182,In_136);
or U5431 (N_5431,In_2118,In_275);
nor U5432 (N_5432,In_425,In_1659);
xnor U5433 (N_5433,In_2333,In_2189);
or U5434 (N_5434,In_498,In_287);
nand U5435 (N_5435,In_781,In_1015);
nand U5436 (N_5436,In_1937,In_931);
xnor U5437 (N_5437,In_2239,In_1211);
nand U5438 (N_5438,In_927,In_1954);
nand U5439 (N_5439,In_1027,In_1144);
xnor U5440 (N_5440,In_1820,In_2088);
nand U5441 (N_5441,In_1223,In_342);
or U5442 (N_5442,In_651,In_641);
or U5443 (N_5443,In_305,In_1025);
xnor U5444 (N_5444,In_912,In_2166);
nor U5445 (N_5445,In_662,In_2144);
or U5446 (N_5446,In_353,In_290);
and U5447 (N_5447,In_2373,In_2414);
xor U5448 (N_5448,In_1978,In_2412);
and U5449 (N_5449,In_1159,In_1263);
nand U5450 (N_5450,In_1466,In_1599);
nand U5451 (N_5451,In_1107,In_832);
nand U5452 (N_5452,In_59,In_1037);
xnor U5453 (N_5453,In_1072,In_176);
xor U5454 (N_5454,In_911,In_1201);
or U5455 (N_5455,In_1441,In_824);
or U5456 (N_5456,In_1838,In_2406);
and U5457 (N_5457,In_1284,In_865);
and U5458 (N_5458,In_1683,In_2341);
xnor U5459 (N_5459,In_647,In_1247);
nand U5460 (N_5460,In_1135,In_672);
nand U5461 (N_5461,In_707,In_1633);
nor U5462 (N_5462,In_139,In_1594);
or U5463 (N_5463,In_1292,In_2377);
nand U5464 (N_5464,In_21,In_2112);
nand U5465 (N_5465,In_2486,In_1083);
nor U5466 (N_5466,In_1973,In_882);
nor U5467 (N_5467,In_857,In_852);
and U5468 (N_5468,In_2279,In_890);
or U5469 (N_5469,In_1560,In_165);
nor U5470 (N_5470,In_1779,In_1040);
xnor U5471 (N_5471,In_1564,In_1513);
nand U5472 (N_5472,In_1674,In_1589);
xnor U5473 (N_5473,In_1103,In_1807);
and U5474 (N_5474,In_218,In_2170);
nand U5475 (N_5475,In_1547,In_1949);
or U5476 (N_5476,In_2342,In_1102);
nor U5477 (N_5477,In_2396,In_1067);
nand U5478 (N_5478,In_252,In_1930);
or U5479 (N_5479,In_1058,In_2209);
and U5480 (N_5480,In_715,In_2462);
or U5481 (N_5481,In_2475,In_1924);
nand U5482 (N_5482,In_391,In_686);
nor U5483 (N_5483,In_2183,In_1077);
nand U5484 (N_5484,In_328,In_1525);
nand U5485 (N_5485,In_728,In_1011);
nand U5486 (N_5486,In_1876,In_1773);
nand U5487 (N_5487,In_1963,In_2340);
and U5488 (N_5488,In_1901,In_103);
nand U5489 (N_5489,In_859,In_732);
nand U5490 (N_5490,In_902,In_2229);
xnor U5491 (N_5491,In_1313,In_19);
or U5492 (N_5492,In_1314,In_761);
nor U5493 (N_5493,In_626,In_210);
or U5494 (N_5494,In_784,In_2411);
nand U5495 (N_5495,In_1036,In_260);
or U5496 (N_5496,In_2087,In_2124);
nand U5497 (N_5497,In_1018,In_10);
nand U5498 (N_5498,In_700,In_1691);
nand U5499 (N_5499,In_1528,In_1529);
xnor U5500 (N_5500,In_596,In_784);
xor U5501 (N_5501,In_2180,In_1055);
and U5502 (N_5502,In_204,In_2079);
xnor U5503 (N_5503,In_245,In_2457);
and U5504 (N_5504,In_1665,In_1105);
xor U5505 (N_5505,In_2186,In_173);
nor U5506 (N_5506,In_1252,In_2116);
or U5507 (N_5507,In_863,In_1757);
nor U5508 (N_5508,In_1361,In_2002);
xnor U5509 (N_5509,In_1467,In_1586);
or U5510 (N_5510,In_689,In_1134);
nand U5511 (N_5511,In_675,In_1737);
nand U5512 (N_5512,In_673,In_1712);
nor U5513 (N_5513,In_1420,In_243);
and U5514 (N_5514,In_1265,In_1419);
or U5515 (N_5515,In_985,In_1046);
nor U5516 (N_5516,In_674,In_2159);
or U5517 (N_5517,In_52,In_1162);
and U5518 (N_5518,In_1082,In_536);
or U5519 (N_5519,In_29,In_81);
or U5520 (N_5520,In_480,In_2256);
nand U5521 (N_5521,In_248,In_517);
or U5522 (N_5522,In_572,In_1198);
nand U5523 (N_5523,In_677,In_1307);
nor U5524 (N_5524,In_1362,In_1326);
and U5525 (N_5525,In_2378,In_1570);
nor U5526 (N_5526,In_214,In_1545);
and U5527 (N_5527,In_2404,In_1258);
nor U5528 (N_5528,In_1530,In_2142);
and U5529 (N_5529,In_337,In_263);
and U5530 (N_5530,In_1148,In_128);
xor U5531 (N_5531,In_735,In_2443);
nor U5532 (N_5532,In_324,In_334);
nor U5533 (N_5533,In_1895,In_1362);
and U5534 (N_5534,In_981,In_1841);
or U5535 (N_5535,In_2399,In_1109);
xnor U5536 (N_5536,In_541,In_2456);
nand U5537 (N_5537,In_1813,In_1642);
nor U5538 (N_5538,In_1737,In_542);
nor U5539 (N_5539,In_908,In_309);
nand U5540 (N_5540,In_1548,In_1804);
xnor U5541 (N_5541,In_1904,In_2456);
and U5542 (N_5542,In_751,In_2130);
nor U5543 (N_5543,In_1715,In_2460);
nor U5544 (N_5544,In_2451,In_1486);
xor U5545 (N_5545,In_439,In_2234);
or U5546 (N_5546,In_1561,In_1433);
nand U5547 (N_5547,In_1461,In_2433);
or U5548 (N_5548,In_1610,In_77);
or U5549 (N_5549,In_450,In_1099);
nor U5550 (N_5550,In_1851,In_942);
nor U5551 (N_5551,In_1189,In_1730);
nand U5552 (N_5552,In_553,In_2090);
and U5553 (N_5553,In_725,In_842);
or U5554 (N_5554,In_1607,In_1566);
nand U5555 (N_5555,In_1113,In_2108);
nand U5556 (N_5556,In_2363,In_1274);
and U5557 (N_5557,In_1287,In_1175);
xor U5558 (N_5558,In_1882,In_633);
nand U5559 (N_5559,In_823,In_334);
nand U5560 (N_5560,In_1574,In_677);
or U5561 (N_5561,In_2396,In_31);
nand U5562 (N_5562,In_1487,In_2214);
and U5563 (N_5563,In_1882,In_2292);
xor U5564 (N_5564,In_1413,In_545);
or U5565 (N_5565,In_1487,In_1020);
and U5566 (N_5566,In_200,In_1952);
or U5567 (N_5567,In_1958,In_2113);
or U5568 (N_5568,In_767,In_1293);
and U5569 (N_5569,In_528,In_306);
nand U5570 (N_5570,In_1867,In_115);
or U5571 (N_5571,In_2420,In_55);
nor U5572 (N_5572,In_1561,In_2051);
xnor U5573 (N_5573,In_1746,In_21);
nand U5574 (N_5574,In_2467,In_1028);
xor U5575 (N_5575,In_1861,In_716);
xor U5576 (N_5576,In_2151,In_323);
and U5577 (N_5577,In_1804,In_2130);
or U5578 (N_5578,In_599,In_66);
nor U5579 (N_5579,In_55,In_1297);
nor U5580 (N_5580,In_2286,In_558);
or U5581 (N_5581,In_1635,In_2190);
and U5582 (N_5582,In_2098,In_954);
xor U5583 (N_5583,In_108,In_1452);
or U5584 (N_5584,In_571,In_974);
and U5585 (N_5585,In_1148,In_1210);
nand U5586 (N_5586,In_1909,In_2285);
and U5587 (N_5587,In_1511,In_1462);
xnor U5588 (N_5588,In_1506,In_1216);
xnor U5589 (N_5589,In_548,In_2270);
xor U5590 (N_5590,In_531,In_1281);
nand U5591 (N_5591,In_1525,In_2320);
or U5592 (N_5592,In_1503,In_1605);
nor U5593 (N_5593,In_2189,In_2370);
nand U5594 (N_5594,In_975,In_1271);
and U5595 (N_5595,In_2056,In_258);
and U5596 (N_5596,In_2274,In_1352);
nor U5597 (N_5597,In_1652,In_2040);
and U5598 (N_5598,In_1949,In_1286);
nand U5599 (N_5599,In_1286,In_212);
xnor U5600 (N_5600,In_2181,In_309);
xor U5601 (N_5601,In_377,In_2408);
xnor U5602 (N_5602,In_1068,In_330);
or U5603 (N_5603,In_433,In_257);
and U5604 (N_5604,In_1693,In_7);
nor U5605 (N_5605,In_1247,In_1890);
and U5606 (N_5606,In_1364,In_347);
and U5607 (N_5607,In_385,In_120);
and U5608 (N_5608,In_1018,In_1751);
xor U5609 (N_5609,In_1539,In_534);
and U5610 (N_5610,In_257,In_869);
nand U5611 (N_5611,In_897,In_1317);
nand U5612 (N_5612,In_85,In_740);
and U5613 (N_5613,In_2149,In_2359);
or U5614 (N_5614,In_124,In_430);
and U5615 (N_5615,In_2490,In_988);
xnor U5616 (N_5616,In_1324,In_215);
and U5617 (N_5617,In_522,In_888);
xor U5618 (N_5618,In_1351,In_5);
or U5619 (N_5619,In_112,In_662);
nand U5620 (N_5620,In_855,In_180);
xor U5621 (N_5621,In_91,In_1693);
nor U5622 (N_5622,In_2344,In_770);
or U5623 (N_5623,In_1053,In_2082);
or U5624 (N_5624,In_2398,In_1034);
nand U5625 (N_5625,In_409,In_2493);
xor U5626 (N_5626,In_1305,In_2174);
xor U5627 (N_5627,In_850,In_1350);
xor U5628 (N_5628,In_1282,In_482);
nand U5629 (N_5629,In_220,In_340);
nand U5630 (N_5630,In_660,In_862);
or U5631 (N_5631,In_1336,In_1083);
nand U5632 (N_5632,In_2221,In_2340);
nor U5633 (N_5633,In_933,In_1156);
nand U5634 (N_5634,In_1407,In_1072);
nor U5635 (N_5635,In_708,In_92);
or U5636 (N_5636,In_739,In_1970);
xnor U5637 (N_5637,In_2016,In_348);
and U5638 (N_5638,In_2199,In_2478);
xor U5639 (N_5639,In_642,In_2279);
and U5640 (N_5640,In_1521,In_2193);
or U5641 (N_5641,In_2293,In_1641);
or U5642 (N_5642,In_1409,In_2052);
nand U5643 (N_5643,In_1309,In_1067);
nand U5644 (N_5644,In_1375,In_1985);
xnor U5645 (N_5645,In_1243,In_334);
and U5646 (N_5646,In_921,In_972);
xor U5647 (N_5647,In_189,In_2192);
or U5648 (N_5648,In_2022,In_2430);
or U5649 (N_5649,In_2441,In_2421);
nand U5650 (N_5650,In_321,In_710);
nor U5651 (N_5651,In_1649,In_216);
nor U5652 (N_5652,In_1368,In_225);
xnor U5653 (N_5653,In_737,In_590);
nor U5654 (N_5654,In_1838,In_1509);
and U5655 (N_5655,In_299,In_312);
nor U5656 (N_5656,In_2435,In_268);
xnor U5657 (N_5657,In_910,In_866);
nand U5658 (N_5658,In_1471,In_1637);
and U5659 (N_5659,In_148,In_555);
nand U5660 (N_5660,In_1919,In_489);
and U5661 (N_5661,In_865,In_250);
and U5662 (N_5662,In_2302,In_1606);
and U5663 (N_5663,In_1,In_127);
xor U5664 (N_5664,In_1774,In_465);
nand U5665 (N_5665,In_1716,In_2051);
nand U5666 (N_5666,In_1093,In_1145);
xor U5667 (N_5667,In_1195,In_722);
xor U5668 (N_5668,In_1091,In_60);
nand U5669 (N_5669,In_1718,In_1588);
nand U5670 (N_5670,In_1554,In_268);
nor U5671 (N_5671,In_46,In_1860);
and U5672 (N_5672,In_535,In_1448);
and U5673 (N_5673,In_2083,In_2280);
nand U5674 (N_5674,In_1310,In_739);
or U5675 (N_5675,In_1345,In_2034);
nor U5676 (N_5676,In_305,In_1242);
xor U5677 (N_5677,In_958,In_1167);
nand U5678 (N_5678,In_2167,In_959);
xnor U5679 (N_5679,In_1481,In_303);
xnor U5680 (N_5680,In_2297,In_1298);
or U5681 (N_5681,In_1373,In_779);
or U5682 (N_5682,In_2025,In_710);
nand U5683 (N_5683,In_155,In_1315);
nand U5684 (N_5684,In_835,In_1372);
xor U5685 (N_5685,In_820,In_1267);
nor U5686 (N_5686,In_314,In_776);
nand U5687 (N_5687,In_717,In_1858);
xnor U5688 (N_5688,In_882,In_720);
nand U5689 (N_5689,In_390,In_360);
xnor U5690 (N_5690,In_2369,In_954);
xor U5691 (N_5691,In_1032,In_1746);
nor U5692 (N_5692,In_2213,In_1372);
nand U5693 (N_5693,In_1000,In_1842);
or U5694 (N_5694,In_1540,In_1976);
or U5695 (N_5695,In_903,In_1756);
xor U5696 (N_5696,In_484,In_908);
nor U5697 (N_5697,In_969,In_549);
and U5698 (N_5698,In_2314,In_1415);
nor U5699 (N_5699,In_627,In_968);
nor U5700 (N_5700,In_1662,In_1937);
nand U5701 (N_5701,In_153,In_2354);
and U5702 (N_5702,In_118,In_2093);
and U5703 (N_5703,In_2379,In_1421);
xor U5704 (N_5704,In_1576,In_339);
xor U5705 (N_5705,In_1275,In_1154);
nand U5706 (N_5706,In_382,In_596);
xnor U5707 (N_5707,In_2428,In_2248);
and U5708 (N_5708,In_1573,In_1814);
and U5709 (N_5709,In_604,In_2021);
or U5710 (N_5710,In_2119,In_2113);
nand U5711 (N_5711,In_291,In_817);
and U5712 (N_5712,In_1553,In_1358);
or U5713 (N_5713,In_2124,In_1532);
or U5714 (N_5714,In_1461,In_1749);
or U5715 (N_5715,In_1017,In_2368);
or U5716 (N_5716,In_263,In_2256);
and U5717 (N_5717,In_1550,In_1068);
nor U5718 (N_5718,In_2088,In_1885);
and U5719 (N_5719,In_1341,In_1468);
nand U5720 (N_5720,In_2134,In_406);
and U5721 (N_5721,In_1693,In_119);
and U5722 (N_5722,In_1588,In_1442);
nor U5723 (N_5723,In_170,In_598);
nor U5724 (N_5724,In_667,In_421);
nand U5725 (N_5725,In_1586,In_601);
xnor U5726 (N_5726,In_1095,In_916);
nor U5727 (N_5727,In_1320,In_265);
nor U5728 (N_5728,In_469,In_1033);
nand U5729 (N_5729,In_2031,In_289);
nor U5730 (N_5730,In_599,In_830);
nand U5731 (N_5731,In_732,In_738);
nand U5732 (N_5732,In_1704,In_2004);
and U5733 (N_5733,In_867,In_1542);
nor U5734 (N_5734,In_1193,In_596);
or U5735 (N_5735,In_1823,In_1063);
xnor U5736 (N_5736,In_2485,In_1788);
nor U5737 (N_5737,In_2358,In_1519);
or U5738 (N_5738,In_1825,In_675);
nand U5739 (N_5739,In_661,In_2118);
and U5740 (N_5740,In_2007,In_1511);
xnor U5741 (N_5741,In_1674,In_1868);
nand U5742 (N_5742,In_554,In_1569);
nand U5743 (N_5743,In_945,In_172);
nand U5744 (N_5744,In_77,In_326);
nand U5745 (N_5745,In_344,In_2383);
and U5746 (N_5746,In_1089,In_600);
nor U5747 (N_5747,In_1663,In_643);
and U5748 (N_5748,In_1971,In_790);
and U5749 (N_5749,In_1601,In_2314);
xnor U5750 (N_5750,In_62,In_1040);
nand U5751 (N_5751,In_1049,In_1956);
nand U5752 (N_5752,In_614,In_821);
nand U5753 (N_5753,In_1111,In_1728);
nor U5754 (N_5754,In_1283,In_1775);
xor U5755 (N_5755,In_174,In_1669);
and U5756 (N_5756,In_51,In_934);
and U5757 (N_5757,In_268,In_933);
and U5758 (N_5758,In_2067,In_851);
and U5759 (N_5759,In_1320,In_88);
nor U5760 (N_5760,In_587,In_101);
and U5761 (N_5761,In_2252,In_1824);
or U5762 (N_5762,In_1407,In_962);
nor U5763 (N_5763,In_777,In_2060);
xor U5764 (N_5764,In_656,In_562);
xor U5765 (N_5765,In_2195,In_2359);
and U5766 (N_5766,In_2123,In_172);
or U5767 (N_5767,In_2402,In_1398);
or U5768 (N_5768,In_722,In_883);
nor U5769 (N_5769,In_1903,In_354);
xor U5770 (N_5770,In_897,In_1742);
nor U5771 (N_5771,In_20,In_2064);
nor U5772 (N_5772,In_673,In_1713);
xor U5773 (N_5773,In_582,In_1115);
or U5774 (N_5774,In_1582,In_271);
or U5775 (N_5775,In_1182,In_2067);
nand U5776 (N_5776,In_2249,In_2289);
nor U5777 (N_5777,In_226,In_1894);
and U5778 (N_5778,In_1204,In_2435);
or U5779 (N_5779,In_563,In_2166);
nor U5780 (N_5780,In_1680,In_2438);
nand U5781 (N_5781,In_1728,In_144);
and U5782 (N_5782,In_991,In_848);
nand U5783 (N_5783,In_2294,In_982);
and U5784 (N_5784,In_1765,In_2461);
or U5785 (N_5785,In_1934,In_1400);
and U5786 (N_5786,In_1419,In_449);
and U5787 (N_5787,In_1994,In_1066);
or U5788 (N_5788,In_898,In_376);
or U5789 (N_5789,In_1789,In_642);
xnor U5790 (N_5790,In_1732,In_1840);
or U5791 (N_5791,In_1744,In_2325);
or U5792 (N_5792,In_2335,In_2241);
nor U5793 (N_5793,In_1752,In_1607);
nand U5794 (N_5794,In_340,In_292);
xor U5795 (N_5795,In_314,In_1491);
nand U5796 (N_5796,In_2476,In_2337);
nand U5797 (N_5797,In_1386,In_1112);
nand U5798 (N_5798,In_1733,In_368);
or U5799 (N_5799,In_89,In_2204);
nand U5800 (N_5800,In_559,In_1601);
nand U5801 (N_5801,In_2115,In_291);
and U5802 (N_5802,In_2158,In_40);
and U5803 (N_5803,In_942,In_2153);
xnor U5804 (N_5804,In_1612,In_1374);
or U5805 (N_5805,In_722,In_1767);
nor U5806 (N_5806,In_65,In_2343);
xnor U5807 (N_5807,In_1181,In_1305);
xor U5808 (N_5808,In_101,In_813);
xor U5809 (N_5809,In_1589,In_2147);
nand U5810 (N_5810,In_148,In_2184);
and U5811 (N_5811,In_436,In_333);
nor U5812 (N_5812,In_244,In_2291);
xor U5813 (N_5813,In_1752,In_150);
nor U5814 (N_5814,In_712,In_1375);
xnor U5815 (N_5815,In_2042,In_215);
nand U5816 (N_5816,In_1608,In_2028);
or U5817 (N_5817,In_1324,In_1322);
and U5818 (N_5818,In_780,In_383);
xnor U5819 (N_5819,In_157,In_1603);
or U5820 (N_5820,In_1976,In_2353);
or U5821 (N_5821,In_1383,In_1869);
and U5822 (N_5822,In_266,In_610);
xor U5823 (N_5823,In_701,In_1696);
xor U5824 (N_5824,In_113,In_515);
nand U5825 (N_5825,In_138,In_1045);
nor U5826 (N_5826,In_1353,In_1467);
and U5827 (N_5827,In_62,In_1855);
nand U5828 (N_5828,In_1219,In_2411);
or U5829 (N_5829,In_1357,In_1418);
nor U5830 (N_5830,In_2042,In_23);
nand U5831 (N_5831,In_2071,In_690);
nor U5832 (N_5832,In_857,In_2203);
and U5833 (N_5833,In_1387,In_1111);
nor U5834 (N_5834,In_177,In_224);
nor U5835 (N_5835,In_1817,In_2140);
nand U5836 (N_5836,In_1805,In_260);
nand U5837 (N_5837,In_256,In_1363);
nand U5838 (N_5838,In_1592,In_1492);
xor U5839 (N_5839,In_231,In_161);
nand U5840 (N_5840,In_414,In_2423);
nor U5841 (N_5841,In_1485,In_225);
or U5842 (N_5842,In_1230,In_919);
nor U5843 (N_5843,In_1138,In_589);
nor U5844 (N_5844,In_392,In_115);
nand U5845 (N_5845,In_155,In_768);
xnor U5846 (N_5846,In_1692,In_1065);
xnor U5847 (N_5847,In_546,In_2230);
nor U5848 (N_5848,In_1834,In_899);
xnor U5849 (N_5849,In_1327,In_1287);
nor U5850 (N_5850,In_15,In_1481);
and U5851 (N_5851,In_654,In_44);
nor U5852 (N_5852,In_260,In_1481);
and U5853 (N_5853,In_2348,In_174);
xnor U5854 (N_5854,In_57,In_98);
nor U5855 (N_5855,In_305,In_2251);
xnor U5856 (N_5856,In_125,In_1195);
and U5857 (N_5857,In_117,In_225);
nor U5858 (N_5858,In_2238,In_754);
or U5859 (N_5859,In_1309,In_413);
nor U5860 (N_5860,In_331,In_280);
xnor U5861 (N_5861,In_1836,In_1869);
or U5862 (N_5862,In_2139,In_2037);
and U5863 (N_5863,In_2350,In_1444);
xnor U5864 (N_5864,In_1176,In_166);
xnor U5865 (N_5865,In_724,In_1212);
and U5866 (N_5866,In_397,In_1537);
nor U5867 (N_5867,In_1240,In_2334);
or U5868 (N_5868,In_232,In_1176);
nand U5869 (N_5869,In_499,In_1934);
xnor U5870 (N_5870,In_718,In_1967);
or U5871 (N_5871,In_2058,In_2076);
xor U5872 (N_5872,In_1151,In_765);
nand U5873 (N_5873,In_123,In_213);
and U5874 (N_5874,In_240,In_788);
xnor U5875 (N_5875,In_1060,In_2069);
nor U5876 (N_5876,In_2344,In_1718);
or U5877 (N_5877,In_1075,In_1287);
nand U5878 (N_5878,In_2108,In_1376);
or U5879 (N_5879,In_193,In_1071);
nor U5880 (N_5880,In_1465,In_179);
or U5881 (N_5881,In_287,In_1452);
or U5882 (N_5882,In_558,In_1835);
or U5883 (N_5883,In_2011,In_158);
nand U5884 (N_5884,In_770,In_1718);
xor U5885 (N_5885,In_1774,In_1102);
and U5886 (N_5886,In_666,In_1581);
and U5887 (N_5887,In_1891,In_326);
nand U5888 (N_5888,In_1436,In_2290);
or U5889 (N_5889,In_1855,In_2220);
xnor U5890 (N_5890,In_1462,In_2264);
xor U5891 (N_5891,In_982,In_416);
nand U5892 (N_5892,In_2329,In_2412);
or U5893 (N_5893,In_1915,In_843);
or U5894 (N_5894,In_1016,In_834);
and U5895 (N_5895,In_216,In_2369);
or U5896 (N_5896,In_2398,In_201);
xor U5897 (N_5897,In_1409,In_2155);
nor U5898 (N_5898,In_1311,In_1985);
or U5899 (N_5899,In_1203,In_97);
and U5900 (N_5900,In_111,In_1901);
and U5901 (N_5901,In_2345,In_1773);
xnor U5902 (N_5902,In_330,In_1764);
or U5903 (N_5903,In_2129,In_1857);
nor U5904 (N_5904,In_861,In_233);
and U5905 (N_5905,In_868,In_1509);
xnor U5906 (N_5906,In_1864,In_577);
nand U5907 (N_5907,In_1313,In_1217);
xnor U5908 (N_5908,In_1553,In_2318);
nand U5909 (N_5909,In_1747,In_1455);
and U5910 (N_5910,In_857,In_1287);
and U5911 (N_5911,In_1632,In_307);
nor U5912 (N_5912,In_825,In_1399);
and U5913 (N_5913,In_1698,In_527);
nand U5914 (N_5914,In_513,In_2115);
xor U5915 (N_5915,In_1585,In_1225);
xor U5916 (N_5916,In_1405,In_2181);
nand U5917 (N_5917,In_1109,In_391);
or U5918 (N_5918,In_28,In_2076);
nand U5919 (N_5919,In_903,In_2002);
nor U5920 (N_5920,In_312,In_1654);
or U5921 (N_5921,In_585,In_1411);
nand U5922 (N_5922,In_1467,In_1790);
nand U5923 (N_5923,In_1970,In_2286);
xor U5924 (N_5924,In_2064,In_1390);
or U5925 (N_5925,In_28,In_1837);
and U5926 (N_5926,In_488,In_1965);
xnor U5927 (N_5927,In_2388,In_405);
nor U5928 (N_5928,In_153,In_1726);
nor U5929 (N_5929,In_22,In_144);
nor U5930 (N_5930,In_439,In_1878);
nor U5931 (N_5931,In_1801,In_1992);
or U5932 (N_5932,In_2145,In_1799);
nor U5933 (N_5933,In_1094,In_62);
and U5934 (N_5934,In_455,In_115);
nand U5935 (N_5935,In_326,In_820);
xor U5936 (N_5936,In_1436,In_2326);
xor U5937 (N_5937,In_655,In_1176);
or U5938 (N_5938,In_2357,In_831);
or U5939 (N_5939,In_2306,In_1898);
nand U5940 (N_5940,In_2332,In_750);
nand U5941 (N_5941,In_1952,In_1844);
xor U5942 (N_5942,In_1543,In_2025);
nor U5943 (N_5943,In_2066,In_933);
xnor U5944 (N_5944,In_1220,In_203);
xor U5945 (N_5945,In_1580,In_1707);
nand U5946 (N_5946,In_2044,In_1952);
and U5947 (N_5947,In_1980,In_733);
or U5948 (N_5948,In_1534,In_1863);
nand U5949 (N_5949,In_82,In_2410);
and U5950 (N_5950,In_995,In_40);
nand U5951 (N_5951,In_2043,In_666);
xnor U5952 (N_5952,In_1630,In_1006);
xor U5953 (N_5953,In_545,In_1880);
xnor U5954 (N_5954,In_1839,In_1265);
nand U5955 (N_5955,In_938,In_1626);
or U5956 (N_5956,In_1657,In_966);
nand U5957 (N_5957,In_1400,In_490);
nand U5958 (N_5958,In_1603,In_860);
or U5959 (N_5959,In_153,In_175);
and U5960 (N_5960,In_700,In_142);
nand U5961 (N_5961,In_767,In_636);
xnor U5962 (N_5962,In_1255,In_2120);
nor U5963 (N_5963,In_1309,In_271);
or U5964 (N_5964,In_2390,In_1648);
xnor U5965 (N_5965,In_692,In_1963);
nand U5966 (N_5966,In_2120,In_2154);
nor U5967 (N_5967,In_1666,In_830);
and U5968 (N_5968,In_1442,In_1162);
nor U5969 (N_5969,In_400,In_1948);
and U5970 (N_5970,In_2313,In_1697);
and U5971 (N_5971,In_336,In_1416);
nand U5972 (N_5972,In_2197,In_605);
and U5973 (N_5973,In_2214,In_197);
xor U5974 (N_5974,In_932,In_1924);
nor U5975 (N_5975,In_2180,In_231);
and U5976 (N_5976,In_1737,In_287);
xor U5977 (N_5977,In_2128,In_1901);
nor U5978 (N_5978,In_584,In_1085);
nand U5979 (N_5979,In_2365,In_1439);
xnor U5980 (N_5980,In_818,In_1924);
nor U5981 (N_5981,In_158,In_205);
or U5982 (N_5982,In_2436,In_2192);
and U5983 (N_5983,In_2184,In_612);
nand U5984 (N_5984,In_817,In_1122);
nand U5985 (N_5985,In_708,In_79);
or U5986 (N_5986,In_2090,In_2322);
and U5987 (N_5987,In_871,In_1722);
xor U5988 (N_5988,In_715,In_586);
or U5989 (N_5989,In_1254,In_1795);
nand U5990 (N_5990,In_1072,In_1293);
or U5991 (N_5991,In_1036,In_1516);
nor U5992 (N_5992,In_1567,In_400);
or U5993 (N_5993,In_573,In_594);
xnor U5994 (N_5994,In_1885,In_1419);
nand U5995 (N_5995,In_350,In_1281);
nand U5996 (N_5996,In_536,In_1149);
or U5997 (N_5997,In_1525,In_1636);
and U5998 (N_5998,In_709,In_1721);
xnor U5999 (N_5999,In_2296,In_2370);
nand U6000 (N_6000,In_422,In_2415);
and U6001 (N_6001,In_2051,In_1048);
xnor U6002 (N_6002,In_2125,In_1385);
nor U6003 (N_6003,In_735,In_2131);
nand U6004 (N_6004,In_1046,In_2466);
nand U6005 (N_6005,In_21,In_791);
or U6006 (N_6006,In_1897,In_1879);
nor U6007 (N_6007,In_1562,In_2317);
xor U6008 (N_6008,In_1815,In_510);
or U6009 (N_6009,In_1071,In_2004);
and U6010 (N_6010,In_512,In_144);
and U6011 (N_6011,In_467,In_171);
xnor U6012 (N_6012,In_1703,In_1535);
xor U6013 (N_6013,In_525,In_198);
nor U6014 (N_6014,In_395,In_437);
nor U6015 (N_6015,In_871,In_554);
and U6016 (N_6016,In_1553,In_2183);
and U6017 (N_6017,In_1970,In_2058);
nand U6018 (N_6018,In_1495,In_2042);
xnor U6019 (N_6019,In_552,In_811);
xnor U6020 (N_6020,In_1892,In_1012);
or U6021 (N_6021,In_2388,In_1192);
and U6022 (N_6022,In_1204,In_2393);
or U6023 (N_6023,In_123,In_1713);
nand U6024 (N_6024,In_669,In_1543);
nand U6025 (N_6025,In_265,In_2457);
nor U6026 (N_6026,In_749,In_2217);
nand U6027 (N_6027,In_576,In_664);
nor U6028 (N_6028,In_2488,In_1991);
nor U6029 (N_6029,In_2011,In_637);
and U6030 (N_6030,In_502,In_94);
nor U6031 (N_6031,In_481,In_139);
or U6032 (N_6032,In_1062,In_2233);
or U6033 (N_6033,In_2419,In_1986);
nand U6034 (N_6034,In_218,In_2468);
nand U6035 (N_6035,In_1201,In_1506);
or U6036 (N_6036,In_744,In_2427);
nand U6037 (N_6037,In_1177,In_601);
xnor U6038 (N_6038,In_763,In_1722);
and U6039 (N_6039,In_2062,In_517);
nor U6040 (N_6040,In_1038,In_866);
and U6041 (N_6041,In_1198,In_811);
or U6042 (N_6042,In_1924,In_83);
nor U6043 (N_6043,In_720,In_495);
or U6044 (N_6044,In_1506,In_1787);
xnor U6045 (N_6045,In_2349,In_2374);
and U6046 (N_6046,In_766,In_1982);
nand U6047 (N_6047,In_2013,In_1235);
nand U6048 (N_6048,In_924,In_1716);
and U6049 (N_6049,In_1704,In_562);
or U6050 (N_6050,In_1692,In_2308);
and U6051 (N_6051,In_346,In_1178);
nand U6052 (N_6052,In_2009,In_2260);
xor U6053 (N_6053,In_941,In_1199);
and U6054 (N_6054,In_1181,In_470);
nor U6055 (N_6055,In_357,In_299);
and U6056 (N_6056,In_2413,In_308);
or U6057 (N_6057,In_983,In_2174);
or U6058 (N_6058,In_2032,In_700);
and U6059 (N_6059,In_947,In_1258);
xor U6060 (N_6060,In_473,In_1777);
nand U6061 (N_6061,In_237,In_2380);
nand U6062 (N_6062,In_1568,In_850);
or U6063 (N_6063,In_102,In_589);
xnor U6064 (N_6064,In_1881,In_690);
xor U6065 (N_6065,In_2170,In_1817);
and U6066 (N_6066,In_2330,In_877);
and U6067 (N_6067,In_534,In_1047);
or U6068 (N_6068,In_488,In_232);
nor U6069 (N_6069,In_2127,In_1944);
nand U6070 (N_6070,In_1850,In_16);
or U6071 (N_6071,In_1200,In_1807);
xor U6072 (N_6072,In_2474,In_1391);
or U6073 (N_6073,In_817,In_2367);
nor U6074 (N_6074,In_124,In_1946);
nor U6075 (N_6075,In_661,In_40);
xnor U6076 (N_6076,In_1850,In_1400);
or U6077 (N_6077,In_707,In_1952);
or U6078 (N_6078,In_1599,In_562);
xor U6079 (N_6079,In_1989,In_1085);
nor U6080 (N_6080,In_611,In_120);
nand U6081 (N_6081,In_1202,In_1871);
nor U6082 (N_6082,In_1905,In_507);
nor U6083 (N_6083,In_2371,In_2445);
xnor U6084 (N_6084,In_85,In_1070);
nand U6085 (N_6085,In_663,In_1105);
xnor U6086 (N_6086,In_522,In_1254);
and U6087 (N_6087,In_819,In_1042);
nand U6088 (N_6088,In_983,In_600);
and U6089 (N_6089,In_1162,In_1319);
and U6090 (N_6090,In_1878,In_42);
and U6091 (N_6091,In_747,In_1218);
and U6092 (N_6092,In_1441,In_1517);
xor U6093 (N_6093,In_306,In_411);
nor U6094 (N_6094,In_190,In_2152);
xnor U6095 (N_6095,In_1636,In_820);
and U6096 (N_6096,In_1791,In_1416);
or U6097 (N_6097,In_1175,In_85);
xnor U6098 (N_6098,In_837,In_915);
xor U6099 (N_6099,In_1567,In_1462);
nand U6100 (N_6100,In_1437,In_1572);
xor U6101 (N_6101,In_63,In_1785);
xor U6102 (N_6102,In_426,In_30);
xnor U6103 (N_6103,In_290,In_2475);
nand U6104 (N_6104,In_1804,In_564);
and U6105 (N_6105,In_1546,In_2051);
xnor U6106 (N_6106,In_2460,In_654);
nand U6107 (N_6107,In_28,In_1982);
nor U6108 (N_6108,In_1611,In_2129);
xor U6109 (N_6109,In_1462,In_1805);
nand U6110 (N_6110,In_2099,In_1910);
or U6111 (N_6111,In_1315,In_990);
nor U6112 (N_6112,In_1106,In_2284);
nand U6113 (N_6113,In_2017,In_2163);
nor U6114 (N_6114,In_2429,In_1662);
or U6115 (N_6115,In_2193,In_1178);
nand U6116 (N_6116,In_717,In_88);
xor U6117 (N_6117,In_1335,In_675);
or U6118 (N_6118,In_327,In_2332);
and U6119 (N_6119,In_438,In_672);
xnor U6120 (N_6120,In_2273,In_1488);
nor U6121 (N_6121,In_1849,In_1787);
nor U6122 (N_6122,In_1162,In_1443);
nand U6123 (N_6123,In_762,In_996);
xnor U6124 (N_6124,In_1584,In_398);
and U6125 (N_6125,In_2158,In_700);
xor U6126 (N_6126,In_986,In_1395);
xnor U6127 (N_6127,In_1056,In_230);
nand U6128 (N_6128,In_834,In_1808);
xnor U6129 (N_6129,In_764,In_2347);
or U6130 (N_6130,In_1634,In_305);
nand U6131 (N_6131,In_1971,In_2141);
and U6132 (N_6132,In_1403,In_1067);
nor U6133 (N_6133,In_1026,In_1993);
xnor U6134 (N_6134,In_2184,In_956);
or U6135 (N_6135,In_2255,In_2249);
nor U6136 (N_6136,In_1001,In_1781);
and U6137 (N_6137,In_1952,In_566);
nand U6138 (N_6138,In_1116,In_904);
and U6139 (N_6139,In_1338,In_219);
nor U6140 (N_6140,In_1789,In_446);
or U6141 (N_6141,In_1813,In_1080);
xnor U6142 (N_6142,In_69,In_2085);
or U6143 (N_6143,In_1677,In_0);
and U6144 (N_6144,In_428,In_531);
nor U6145 (N_6145,In_893,In_1705);
nor U6146 (N_6146,In_1357,In_2374);
and U6147 (N_6147,In_2406,In_2011);
or U6148 (N_6148,In_1168,In_1425);
nor U6149 (N_6149,In_385,In_49);
xnor U6150 (N_6150,In_1911,In_1821);
or U6151 (N_6151,In_1372,In_1082);
or U6152 (N_6152,In_481,In_121);
nor U6153 (N_6153,In_2087,In_1132);
nor U6154 (N_6154,In_1926,In_1523);
and U6155 (N_6155,In_2177,In_1148);
and U6156 (N_6156,In_2340,In_1430);
nand U6157 (N_6157,In_341,In_2162);
xnor U6158 (N_6158,In_116,In_32);
and U6159 (N_6159,In_2070,In_49);
and U6160 (N_6160,In_704,In_2482);
nand U6161 (N_6161,In_1774,In_1193);
and U6162 (N_6162,In_1335,In_2329);
or U6163 (N_6163,In_2145,In_467);
nor U6164 (N_6164,In_1887,In_2127);
or U6165 (N_6165,In_1206,In_1508);
xnor U6166 (N_6166,In_1564,In_1947);
nor U6167 (N_6167,In_86,In_2199);
xnor U6168 (N_6168,In_262,In_1997);
nand U6169 (N_6169,In_827,In_258);
xnor U6170 (N_6170,In_101,In_2381);
or U6171 (N_6171,In_2469,In_929);
nor U6172 (N_6172,In_517,In_2058);
xor U6173 (N_6173,In_174,In_2228);
or U6174 (N_6174,In_1466,In_1242);
nor U6175 (N_6175,In_1726,In_1177);
and U6176 (N_6176,In_302,In_823);
and U6177 (N_6177,In_1413,In_1732);
nand U6178 (N_6178,In_1330,In_283);
nor U6179 (N_6179,In_935,In_1909);
or U6180 (N_6180,In_504,In_989);
nand U6181 (N_6181,In_2127,In_1332);
or U6182 (N_6182,In_736,In_141);
nor U6183 (N_6183,In_943,In_1132);
or U6184 (N_6184,In_948,In_2442);
or U6185 (N_6185,In_1193,In_1234);
and U6186 (N_6186,In_2130,In_1784);
nor U6187 (N_6187,In_1513,In_217);
xor U6188 (N_6188,In_895,In_393);
or U6189 (N_6189,In_1556,In_2165);
nor U6190 (N_6190,In_1503,In_2422);
nor U6191 (N_6191,In_1654,In_1138);
nor U6192 (N_6192,In_1120,In_718);
xnor U6193 (N_6193,In_2484,In_2372);
nor U6194 (N_6194,In_1282,In_388);
nor U6195 (N_6195,In_166,In_931);
nand U6196 (N_6196,In_1297,In_1788);
and U6197 (N_6197,In_1521,In_1181);
and U6198 (N_6198,In_1053,In_2158);
and U6199 (N_6199,In_528,In_57);
and U6200 (N_6200,In_939,In_613);
xor U6201 (N_6201,In_499,In_1914);
nor U6202 (N_6202,In_960,In_956);
xnor U6203 (N_6203,In_2232,In_2227);
or U6204 (N_6204,In_2373,In_1390);
nand U6205 (N_6205,In_1152,In_488);
or U6206 (N_6206,In_147,In_200);
nand U6207 (N_6207,In_1039,In_955);
or U6208 (N_6208,In_1342,In_2429);
xor U6209 (N_6209,In_1125,In_1547);
and U6210 (N_6210,In_246,In_378);
nand U6211 (N_6211,In_929,In_892);
or U6212 (N_6212,In_2027,In_1653);
nor U6213 (N_6213,In_1734,In_901);
xnor U6214 (N_6214,In_1368,In_1222);
and U6215 (N_6215,In_2176,In_1774);
xor U6216 (N_6216,In_2130,In_1621);
xor U6217 (N_6217,In_1311,In_125);
xor U6218 (N_6218,In_831,In_771);
and U6219 (N_6219,In_2149,In_1362);
and U6220 (N_6220,In_57,In_2054);
nand U6221 (N_6221,In_2371,In_986);
or U6222 (N_6222,In_1416,In_986);
and U6223 (N_6223,In_2406,In_811);
nand U6224 (N_6224,In_2264,In_2242);
and U6225 (N_6225,In_1331,In_2443);
or U6226 (N_6226,In_2158,In_2424);
nand U6227 (N_6227,In_1197,In_828);
xor U6228 (N_6228,In_2049,In_289);
xnor U6229 (N_6229,In_2483,In_1765);
nand U6230 (N_6230,In_315,In_102);
nand U6231 (N_6231,In_1300,In_1560);
nor U6232 (N_6232,In_377,In_316);
and U6233 (N_6233,In_933,In_2408);
nor U6234 (N_6234,In_419,In_1371);
nand U6235 (N_6235,In_912,In_579);
nor U6236 (N_6236,In_1205,In_232);
xor U6237 (N_6237,In_993,In_453);
and U6238 (N_6238,In_1741,In_724);
xor U6239 (N_6239,In_423,In_478);
and U6240 (N_6240,In_779,In_2110);
or U6241 (N_6241,In_97,In_1219);
and U6242 (N_6242,In_973,In_863);
xor U6243 (N_6243,In_856,In_983);
nor U6244 (N_6244,In_2255,In_2456);
nor U6245 (N_6245,In_1812,In_1804);
nor U6246 (N_6246,In_373,In_2144);
or U6247 (N_6247,In_375,In_1203);
nor U6248 (N_6248,In_2104,In_1723);
nand U6249 (N_6249,In_490,In_1677);
nor U6250 (N_6250,N_3843,N_3506);
or U6251 (N_6251,N_3238,N_5556);
nor U6252 (N_6252,N_1413,N_1583);
or U6253 (N_6253,N_3092,N_93);
nor U6254 (N_6254,N_1173,N_4999);
or U6255 (N_6255,N_6081,N_435);
and U6256 (N_6256,N_2340,N_2023);
and U6257 (N_6257,N_1677,N_1490);
nand U6258 (N_6258,N_6128,N_2859);
nand U6259 (N_6259,N_2891,N_5810);
and U6260 (N_6260,N_5306,N_4804);
nand U6261 (N_6261,N_4249,N_1889);
or U6262 (N_6262,N_2950,N_3138);
or U6263 (N_6263,N_4780,N_5377);
and U6264 (N_6264,N_3760,N_5059);
nand U6265 (N_6265,N_3701,N_2805);
and U6266 (N_6266,N_430,N_3959);
and U6267 (N_6267,N_3008,N_1547);
or U6268 (N_6268,N_5041,N_3046);
nand U6269 (N_6269,N_1638,N_3421);
nand U6270 (N_6270,N_2296,N_1942);
xor U6271 (N_6271,N_5,N_4374);
nand U6272 (N_6272,N_799,N_5955);
nand U6273 (N_6273,N_913,N_529);
nor U6274 (N_6274,N_140,N_5993);
nand U6275 (N_6275,N_40,N_4868);
nor U6276 (N_6276,N_3482,N_1189);
or U6277 (N_6277,N_2188,N_3490);
or U6278 (N_6278,N_2815,N_3463);
nor U6279 (N_6279,N_5359,N_4363);
and U6280 (N_6280,N_901,N_4049);
or U6281 (N_6281,N_5990,N_1176);
nand U6282 (N_6282,N_5658,N_2000);
nor U6283 (N_6283,N_2982,N_4176);
and U6284 (N_6284,N_619,N_1251);
nor U6285 (N_6285,N_5011,N_876);
xnor U6286 (N_6286,N_2534,N_5326);
or U6287 (N_6287,N_4264,N_3938);
nand U6288 (N_6288,N_4972,N_2562);
or U6289 (N_6289,N_625,N_271);
and U6290 (N_6290,N_1577,N_2223);
nand U6291 (N_6291,N_2772,N_5651);
and U6292 (N_6292,N_229,N_1842);
or U6293 (N_6293,N_347,N_6090);
xor U6294 (N_6294,N_2084,N_4193);
xor U6295 (N_6295,N_2732,N_2002);
xnor U6296 (N_6296,N_5272,N_896);
xnor U6297 (N_6297,N_2569,N_5594);
xor U6298 (N_6298,N_2013,N_1603);
and U6299 (N_6299,N_4278,N_1010);
nand U6300 (N_6300,N_1626,N_792);
or U6301 (N_6301,N_5974,N_1211);
xor U6302 (N_6302,N_6199,N_3708);
xor U6303 (N_6303,N_2680,N_5816);
or U6304 (N_6304,N_1962,N_426);
or U6305 (N_6305,N_818,N_3095);
xor U6306 (N_6306,N_2789,N_233);
or U6307 (N_6307,N_1556,N_1804);
nand U6308 (N_6308,N_2908,N_1641);
nor U6309 (N_6309,N_1148,N_584);
nand U6310 (N_6310,N_488,N_2739);
and U6311 (N_6311,N_3732,N_2215);
xnor U6312 (N_6312,N_2916,N_310);
and U6313 (N_6313,N_1769,N_3408);
nand U6314 (N_6314,N_976,N_2216);
or U6315 (N_6315,N_5561,N_4867);
and U6316 (N_6316,N_4639,N_4001);
or U6317 (N_6317,N_2328,N_4813);
nor U6318 (N_6318,N_3560,N_4325);
nand U6319 (N_6319,N_3700,N_4471);
nand U6320 (N_6320,N_1389,N_3153);
and U6321 (N_6321,N_3278,N_1508);
nand U6322 (N_6322,N_2498,N_5058);
or U6323 (N_6323,N_3699,N_4940);
nand U6324 (N_6324,N_3897,N_1921);
nor U6325 (N_6325,N_1614,N_5464);
nand U6326 (N_6326,N_4633,N_1798);
nand U6327 (N_6327,N_5918,N_1534);
xor U6328 (N_6328,N_1482,N_2454);
nor U6329 (N_6329,N_2494,N_6115);
or U6330 (N_6330,N_3478,N_1639);
or U6331 (N_6331,N_956,N_5111);
nor U6332 (N_6332,N_2261,N_3289);
nand U6333 (N_6333,N_2374,N_4463);
nor U6334 (N_6334,N_6159,N_2400);
and U6335 (N_6335,N_1347,N_1179);
xor U6336 (N_6336,N_4918,N_4606);
xnor U6337 (N_6337,N_2074,N_3099);
xor U6338 (N_6338,N_3185,N_1270);
nor U6339 (N_6339,N_2723,N_4225);
nor U6340 (N_6340,N_2055,N_5767);
or U6341 (N_6341,N_4583,N_4305);
and U6342 (N_6342,N_4259,N_1372);
and U6343 (N_6343,N_3829,N_4263);
nand U6344 (N_6344,N_507,N_3369);
nand U6345 (N_6345,N_1784,N_4162);
nand U6346 (N_6346,N_1339,N_348);
xnor U6347 (N_6347,N_5803,N_3895);
nand U6348 (N_6348,N_3671,N_5087);
nor U6349 (N_6349,N_5074,N_977);
nor U6350 (N_6350,N_1916,N_5590);
and U6351 (N_6351,N_27,N_5134);
or U6352 (N_6352,N_2049,N_739);
xnor U6353 (N_6353,N_3413,N_2128);
and U6354 (N_6354,N_2260,N_2620);
or U6355 (N_6355,N_3676,N_5657);
xor U6356 (N_6356,N_4369,N_5690);
or U6357 (N_6357,N_2862,N_5614);
nand U6358 (N_6358,N_159,N_5686);
nor U6359 (N_6359,N_113,N_4923);
or U6360 (N_6360,N_1119,N_4292);
or U6361 (N_6361,N_6204,N_2967);
or U6362 (N_6362,N_615,N_5329);
and U6363 (N_6363,N_1289,N_87);
xor U6364 (N_6364,N_5380,N_3140);
nor U6365 (N_6365,N_389,N_5739);
nand U6366 (N_6366,N_2721,N_1852);
and U6367 (N_6367,N_5700,N_2780);
nor U6368 (N_6368,N_5897,N_2966);
nand U6369 (N_6369,N_4543,N_5519);
xnor U6370 (N_6370,N_700,N_1535);
or U6371 (N_6371,N_4159,N_2095);
nor U6372 (N_6372,N_342,N_2190);
xnor U6373 (N_6373,N_3129,N_5741);
nor U6374 (N_6374,N_3821,N_474);
nand U6375 (N_6375,N_5917,N_1532);
and U6376 (N_6376,N_2647,N_2194);
nand U6377 (N_6377,N_4073,N_320);
and U6378 (N_6378,N_3545,N_2842);
or U6379 (N_6379,N_1878,N_4320);
nor U6380 (N_6380,N_3859,N_668);
or U6381 (N_6381,N_6154,N_3541);
or U6382 (N_6382,N_3476,N_765);
and U6383 (N_6383,N_349,N_6150);
xnor U6384 (N_6384,N_5900,N_610);
xor U6385 (N_6385,N_1805,N_4146);
nor U6386 (N_6386,N_51,N_1409);
nand U6387 (N_6387,N_156,N_3668);
xor U6388 (N_6388,N_3941,N_2821);
nor U6389 (N_6389,N_3537,N_3287);
or U6390 (N_6390,N_1651,N_2272);
and U6391 (N_6391,N_3691,N_3343);
xor U6392 (N_6392,N_64,N_1129);
nand U6393 (N_6393,N_2621,N_44);
or U6394 (N_6394,N_1445,N_5886);
and U6395 (N_6395,N_4796,N_3515);
nand U6396 (N_6396,N_5819,N_3192);
xnor U6397 (N_6397,N_2129,N_3164);
or U6398 (N_6398,N_83,N_1733);
nor U6399 (N_6399,N_5332,N_2477);
nor U6400 (N_6400,N_6216,N_1034);
xor U6401 (N_6401,N_4569,N_1764);
nor U6402 (N_6402,N_6135,N_407);
nor U6403 (N_6403,N_1366,N_4085);
or U6404 (N_6404,N_2973,N_5777);
or U6405 (N_6405,N_2380,N_1067);
nor U6406 (N_6406,N_4290,N_5112);
or U6407 (N_6407,N_5082,N_6210);
or U6408 (N_6408,N_1407,N_560);
xor U6409 (N_6409,N_3266,N_4879);
xor U6410 (N_6410,N_5562,N_4476);
nand U6411 (N_6411,N_3686,N_692);
or U6412 (N_6412,N_3063,N_3646);
nor U6413 (N_6413,N_106,N_2742);
xor U6414 (N_6414,N_2849,N_2524);
nand U6415 (N_6415,N_4704,N_939);
and U6416 (N_6416,N_6231,N_1054);
nor U6417 (N_6417,N_5608,N_6003);
nand U6418 (N_6418,N_4957,N_1674);
nand U6419 (N_6419,N_290,N_4641);
xor U6420 (N_6420,N_4321,N_5143);
or U6421 (N_6421,N_3911,N_3122);
nand U6422 (N_6422,N_1090,N_774);
nor U6423 (N_6423,N_2236,N_5707);
xnor U6424 (N_6424,N_3399,N_5487);
nor U6425 (N_6425,N_5890,N_4803);
xnor U6426 (N_6426,N_5798,N_3009);
xor U6427 (N_6427,N_871,N_3228);
nor U6428 (N_6428,N_2635,N_2965);
xor U6429 (N_6429,N_2545,N_237);
nor U6430 (N_6430,N_5766,N_3749);
xor U6431 (N_6431,N_751,N_3587);
nand U6432 (N_6432,N_2535,N_6059);
nand U6433 (N_6433,N_4198,N_168);
or U6434 (N_6434,N_3487,N_4179);
and U6435 (N_6435,N_2774,N_5737);
or U6436 (N_6436,N_5928,N_975);
xor U6437 (N_6437,N_4802,N_5845);
and U6438 (N_6438,N_1205,N_4618);
xnor U6439 (N_6439,N_2082,N_2786);
nand U6440 (N_6440,N_6075,N_4514);
or U6441 (N_6441,N_3499,N_5335);
nand U6442 (N_6442,N_2096,N_5175);
and U6443 (N_6443,N_2111,N_3147);
nand U6444 (N_6444,N_6104,N_2040);
xor U6445 (N_6445,N_2760,N_4040);
and U6446 (N_6446,N_5314,N_5239);
xnor U6447 (N_6447,N_2605,N_3933);
and U6448 (N_6448,N_6108,N_635);
or U6449 (N_6449,N_577,N_1304);
nand U6450 (N_6450,N_2764,N_1660);
xor U6451 (N_6451,N_4283,N_831);
or U6452 (N_6452,N_1790,N_2905);
xnor U6453 (N_6453,N_48,N_3398);
nor U6454 (N_6454,N_4980,N_2998);
and U6455 (N_6455,N_427,N_1106);
or U6456 (N_6456,N_941,N_752);
nor U6457 (N_6457,N_1196,N_5467);
nand U6458 (N_6458,N_3524,N_2008);
or U6459 (N_6459,N_1448,N_5480);
or U6460 (N_6460,N_5217,N_583);
nor U6461 (N_6461,N_727,N_1871);
xor U6462 (N_6462,N_5310,N_5781);
nor U6463 (N_6463,N_1507,N_721);
or U6464 (N_6464,N_2432,N_3172);
nor U6465 (N_6465,N_3241,N_3738);
nand U6466 (N_6466,N_101,N_1337);
and U6467 (N_6467,N_5482,N_4693);
xnor U6468 (N_6468,N_2897,N_2738);
or U6469 (N_6469,N_2991,N_5303);
nand U6470 (N_6470,N_3724,N_190);
and U6471 (N_6471,N_1588,N_5746);
nor U6472 (N_6472,N_1446,N_3272);
xor U6473 (N_6473,N_3324,N_3341);
or U6474 (N_6474,N_4845,N_578);
or U6475 (N_6475,N_2172,N_3096);
nand U6476 (N_6476,N_4974,N_1938);
and U6477 (N_6477,N_3376,N_3719);
or U6478 (N_6478,N_911,N_5876);
nand U6479 (N_6479,N_1743,N_4554);
xor U6480 (N_6480,N_5761,N_6226);
xor U6481 (N_6481,N_1041,N_1057);
nor U6482 (N_6482,N_3458,N_1715);
nor U6483 (N_6483,N_1308,N_2943);
or U6484 (N_6484,N_3932,N_6246);
and U6485 (N_6485,N_708,N_1455);
and U6486 (N_6486,N_5277,N_714);
or U6487 (N_6487,N_1517,N_2389);
nand U6488 (N_6488,N_6225,N_3202);
or U6489 (N_6489,N_3828,N_2441);
xnor U6490 (N_6490,N_2480,N_4860);
nand U6491 (N_6491,N_5297,N_3437);
xor U6492 (N_6492,N_1462,N_2748);
or U6493 (N_6493,N_5585,N_2689);
nand U6494 (N_6494,N_2708,N_4828);
and U6495 (N_6495,N_1736,N_5232);
nor U6496 (N_6496,N_461,N_3423);
and U6497 (N_6497,N_3893,N_5525);
nand U6498 (N_6498,N_3705,N_1134);
nor U6499 (N_6499,N_3525,N_3687);
xor U6500 (N_6500,N_4344,N_5696);
xor U6501 (N_6501,N_2561,N_3851);
nor U6502 (N_6502,N_1653,N_1201);
nand U6503 (N_6503,N_4169,N_3277);
nor U6504 (N_6504,N_2343,N_1404);
nor U6505 (N_6505,N_894,N_1716);
nor U6506 (N_6506,N_6234,N_3247);
xnor U6507 (N_6507,N_3345,N_3579);
nand U6508 (N_6508,N_6060,N_2066);
nor U6509 (N_6509,N_1744,N_2078);
nor U6510 (N_6510,N_1021,N_2895);
nor U6511 (N_6511,N_4748,N_3470);
and U6512 (N_6512,N_332,N_4635);
xor U6513 (N_6513,N_2985,N_2624);
xor U6514 (N_6514,N_4032,N_3349);
or U6515 (N_6515,N_1786,N_183);
nand U6516 (N_6516,N_1515,N_3330);
nor U6517 (N_6517,N_3471,N_4869);
xor U6518 (N_6518,N_431,N_3226);
nand U6519 (N_6519,N_4960,N_4334);
xor U6520 (N_6520,N_2176,N_4063);
xnor U6521 (N_6521,N_2458,N_2134);
and U6522 (N_6522,N_4136,N_1607);
or U6523 (N_6523,N_5709,N_1964);
or U6524 (N_6524,N_2338,N_5397);
and U6525 (N_6525,N_1321,N_4938);
and U6526 (N_6526,N_3607,N_5252);
or U6527 (N_6527,N_4781,N_3081);
and U6528 (N_6528,N_5991,N_4757);
xor U6529 (N_6529,N_734,N_4392);
or U6530 (N_6530,N_198,N_2779);
nor U6531 (N_6531,N_5345,N_3703);
and U6532 (N_6532,N_722,N_5906);
or U6533 (N_6533,N_5904,N_4586);
xnor U6534 (N_6534,N_4042,N_3294);
nor U6535 (N_6535,N_1777,N_5193);
or U6536 (N_6536,N_5527,N_2807);
nor U6537 (N_6537,N_2553,N_2923);
and U6538 (N_6538,N_5455,N_2077);
or U6539 (N_6539,N_2204,N_5206);
nor U6540 (N_6540,N_2718,N_5593);
and U6541 (N_6541,N_2045,N_6176);
or U6542 (N_6542,N_5754,N_549);
nor U6543 (N_6543,N_1390,N_4562);
or U6544 (N_6544,N_151,N_4516);
nor U6545 (N_6545,N_4665,N_2875);
nand U6546 (N_6546,N_1331,N_637);
nand U6547 (N_6547,N_4791,N_6228);
xor U6548 (N_6548,N_5508,N_5638);
or U6549 (N_6549,N_5178,N_5718);
or U6550 (N_6550,N_3556,N_2184);
nor U6551 (N_6551,N_3880,N_1579);
nor U6552 (N_6552,N_4673,N_2207);
xor U6553 (N_6553,N_3675,N_4642);
nand U6554 (N_6554,N_4445,N_3683);
nor U6555 (N_6555,N_5174,N_5901);
nor U6556 (N_6556,N_1081,N_4440);
and U6557 (N_6557,N_268,N_987);
nand U6558 (N_6558,N_4150,N_2335);
nor U6559 (N_6559,N_5829,N_2657);
and U6560 (N_6560,N_5828,N_5615);
nand U6561 (N_6561,N_810,N_5850);
xnor U6562 (N_6562,N_2741,N_7);
nor U6563 (N_6563,N_3335,N_3455);
nand U6564 (N_6564,N_1381,N_1548);
or U6565 (N_6565,N_5428,N_3130);
nor U6566 (N_6566,N_2039,N_477);
xor U6567 (N_6567,N_793,N_4973);
nor U6568 (N_6568,N_5610,N_2366);
xor U6569 (N_6569,N_2823,N_2877);
nand U6570 (N_6570,N_966,N_1511);
nand U6571 (N_6571,N_6100,N_5858);
nor U6572 (N_6572,N_4409,N_3281);
nor U6573 (N_6573,N_3769,N_1305);
nand U6574 (N_6574,N_1088,N_2163);
nand U6575 (N_6575,N_798,N_386);
nor U6576 (N_6576,N_5211,N_2566);
nor U6577 (N_6577,N_3855,N_656);
nor U6578 (N_6578,N_6137,N_2878);
nand U6579 (N_6579,N_2556,N_4911);
or U6580 (N_6580,N_2714,N_105);
nand U6581 (N_6581,N_5348,N_2051);
xor U6582 (N_6582,N_1433,N_5465);
xnor U6583 (N_6583,N_2012,N_1049);
and U6584 (N_6584,N_3778,N_1735);
nand U6585 (N_6585,N_4667,N_4664);
or U6586 (N_6586,N_5870,N_2161);
nor U6587 (N_6587,N_4393,N_45);
nor U6588 (N_6588,N_4731,N_4446);
xor U6589 (N_6589,N_6052,N_6054);
nor U6590 (N_6590,N_2722,N_4276);
nor U6591 (N_6591,N_1818,N_1279);
nor U6592 (N_6592,N_4462,N_2479);
nand U6593 (N_6593,N_4189,N_2349);
nor U6594 (N_6594,N_2080,N_3826);
or U6595 (N_6595,N_1956,N_5756);
or U6596 (N_6596,N_4466,N_3543);
nor U6597 (N_6597,N_981,N_2928);
and U6598 (N_6598,N_150,N_5507);
xor U6599 (N_6599,N_1874,N_3093);
and U6600 (N_6600,N_4338,N_5064);
or U6601 (N_6601,N_1913,N_1354);
and U6602 (N_6602,N_266,N_444);
xor U6603 (N_6603,N_5823,N_1685);
nand U6604 (N_6604,N_2579,N_2578);
nor U6605 (N_6605,N_5836,N_224);
xnor U6606 (N_6606,N_3242,N_621);
nor U6607 (N_6607,N_5745,N_3114);
or U6608 (N_6608,N_2469,N_445);
xnor U6609 (N_6609,N_686,N_523);
xor U6610 (N_6610,N_4453,N_3726);
xor U6611 (N_6611,N_4257,N_3088);
xor U6612 (N_6612,N_861,N_4082);
and U6613 (N_6613,N_314,N_5156);
nor U6614 (N_6614,N_665,N_4906);
or U6615 (N_6615,N_5595,N_1812);
or U6616 (N_6616,N_804,N_1949);
xor U6617 (N_6617,N_849,N_5555);
and U6618 (N_6618,N_3514,N_2440);
or U6619 (N_6619,N_6130,N_3682);
or U6620 (N_6620,N_1615,N_5912);
nor U6621 (N_6621,N_5558,N_3201);
or U6622 (N_6622,N_1906,N_2234);
or U6623 (N_6623,N_3120,N_5056);
nor U6624 (N_6624,N_3190,N_6190);
nor U6625 (N_6625,N_4203,N_1491);
or U6626 (N_6626,N_139,N_5732);
nand U6627 (N_6627,N_1678,N_590);
and U6628 (N_6628,N_1699,N_1611);
or U6629 (N_6629,N_4644,N_3152);
and U6630 (N_6630,N_2658,N_4750);
xnor U6631 (N_6631,N_2590,N_1836);
or U6632 (N_6632,N_2098,N_2397);
nor U6633 (N_6633,N_2761,N_318);
nor U6634 (N_6634,N_3344,N_1862);
nor U6635 (N_6635,N_687,N_2633);
nor U6636 (N_6636,N_3244,N_3797);
or U6637 (N_6637,N_2883,N_4410);
or U6638 (N_6638,N_4324,N_726);
and U6639 (N_6639,N_5811,N_5675);
nor U6640 (N_6640,N_1309,N_4336);
nor U6641 (N_6641,N_1568,N_2818);
nor U6642 (N_6642,N_1095,N_5855);
and U6643 (N_6643,N_3755,N_3022);
nand U6644 (N_6644,N_4795,N_3663);
or U6645 (N_6645,N_1165,N_3605);
nor U6646 (N_6646,N_1099,N_344);
nor U6647 (N_6647,N_2568,N_4502);
xnor U6648 (N_6648,N_1450,N_120);
nand U6649 (N_6649,N_416,N_2220);
xnor U6650 (N_6650,N_1145,N_4937);
xnor U6651 (N_6651,N_5568,N_542);
nand U6652 (N_6652,N_628,N_5450);
or U6653 (N_6653,N_1600,N_2915);
or U6654 (N_6654,N_3271,N_4855);
nand U6655 (N_6655,N_5880,N_4649);
or U6656 (N_6656,N_634,N_3825);
xnor U6657 (N_6657,N_5526,N_5616);
or U6658 (N_6658,N_2911,N_4391);
and U6659 (N_6659,N_3800,N_3417);
or U6660 (N_6660,N_3823,N_4472);
nand U6661 (N_6661,N_3910,N_5559);
and U6662 (N_6662,N_4303,N_2555);
or U6663 (N_6663,N_6151,N_1839);
nand U6664 (N_6664,N_2984,N_3824);
nand U6665 (N_6665,N_2169,N_5418);
and U6666 (N_6666,N_5694,N_6209);
nand U6667 (N_6667,N_5948,N_4547);
nor U6668 (N_6668,N_1073,N_5395);
or U6669 (N_6669,N_1275,N_2268);
or U6670 (N_6670,N_5822,N_3637);
nand U6671 (N_6671,N_3697,N_3613);
xnor U6672 (N_6672,N_4468,N_328);
xor U6673 (N_6673,N_4811,N_4527);
xor U6674 (N_6674,N_3467,N_3213);
nor U6675 (N_6675,N_6085,N_5516);
xnor U6676 (N_6676,N_2197,N_1302);
and U6677 (N_6677,N_4655,N_1524);
nor U6678 (N_6678,N_161,N_3457);
xnor U6679 (N_6679,N_3507,N_5454);
or U6680 (N_6680,N_3384,N_4966);
nand U6681 (N_6681,N_2986,N_3685);
xnor U6682 (N_6682,N_1055,N_775);
nor U6683 (N_6683,N_1139,N_1665);
nor U6684 (N_6684,N_6079,N_2470);
xnor U6685 (N_6685,N_4856,N_4380);
xnor U6686 (N_6686,N_580,N_1545);
nand U6687 (N_6687,N_405,N_2314);
xnor U6688 (N_6688,N_5824,N_3660);
xor U6689 (N_6689,N_3297,N_5931);
xor U6690 (N_6690,N_5153,N_1071);
xor U6691 (N_6691,N_1746,N_3498);
xnor U6692 (N_6692,N_2613,N_814);
or U6693 (N_6693,N_1965,N_5503);
or U6694 (N_6694,N_6141,N_3766);
or U6695 (N_6695,N_3314,N_2563);
nand U6696 (N_6696,N_1108,N_1306);
nand U6697 (N_6697,N_999,N_2370);
and U6698 (N_6698,N_2054,N_1598);
and U6699 (N_6699,N_1555,N_5144);
nor U6700 (N_6700,N_5970,N_4091);
nand U6701 (N_6701,N_3564,N_4946);
nand U6702 (N_6702,N_3805,N_4822);
nor U6703 (N_6703,N_4039,N_4112);
nor U6704 (N_6704,N_1819,N_1877);
and U6705 (N_6705,N_2806,N_1575);
xor U6706 (N_6706,N_1268,N_4261);
nand U6707 (N_6707,N_1719,N_4935);
nand U6708 (N_6708,N_423,N_91);
xnor U6709 (N_6709,N_203,N_5316);
nor U6710 (N_6710,N_4158,N_253);
xor U6711 (N_6711,N_4794,N_829);
nand U6712 (N_6712,N_5612,N_2766);
nor U6713 (N_6713,N_2421,N_5203);
nand U6714 (N_6714,N_3999,N_1032);
xnor U6715 (N_6715,N_5223,N_4018);
and U6716 (N_6716,N_3632,N_585);
nand U6717 (N_6717,N_3364,N_2593);
nor U6718 (N_6718,N_2119,N_690);
nor U6719 (N_6719,N_4931,N_6068);
nor U6720 (N_6720,N_3353,N_4675);
nor U6721 (N_6721,N_125,N_217);
xor U6722 (N_6722,N_669,N_5089);
or U6723 (N_6723,N_4211,N_6146);
nand U6724 (N_6724,N_4242,N_2071);
xnor U6725 (N_6725,N_4055,N_673);
nor U6726 (N_6726,N_5606,N_403);
and U6727 (N_6727,N_6050,N_3742);
or U6728 (N_6728,N_5280,N_5173);
xnor U6729 (N_6729,N_6131,N_3856);
nand U6730 (N_6730,N_929,N_4568);
and U6731 (N_6731,N_1405,N_5892);
or U6732 (N_6732,N_1367,N_4429);
nor U6733 (N_6733,N_2401,N_5945);
nor U6734 (N_6734,N_2158,N_4300);
and U6735 (N_6735,N_4873,N_1834);
nor U6736 (N_6736,N_36,N_3420);
xor U6737 (N_6737,N_5967,N_3763);
or U6738 (N_6738,N_2402,N_1799);
xnor U6739 (N_6739,N_2924,N_3181);
or U6740 (N_6740,N_3368,N_2627);
nor U6741 (N_6741,N_3206,N_6196);
nand U6742 (N_6742,N_1033,N_3979);
or U6743 (N_6743,N_4691,N_3149);
nand U6744 (N_6744,N_5935,N_3098);
nor U6745 (N_6745,N_568,N_3248);
nand U6746 (N_6746,N_350,N_5874);
nor U6747 (N_6747,N_3267,N_5069);
nor U6748 (N_6748,N_408,N_1789);
and U6749 (N_6749,N_4953,N_3552);
xnor U6750 (N_6750,N_2203,N_3581);
and U6751 (N_6751,N_3912,N_2792);
nor U6752 (N_6752,N_616,N_3307);
and U6753 (N_6753,N_5301,N_4266);
xnor U6754 (N_6754,N_6102,N_1996);
nor U6755 (N_6755,N_3061,N_1479);
or U6756 (N_6756,N_1398,N_6160);
nor U6757 (N_6757,N_1585,N_3808);
and U6758 (N_6758,N_3131,N_78);
nor U6759 (N_6759,N_5607,N_5814);
xnor U6760 (N_6760,N_1707,N_1872);
nor U6761 (N_6761,N_1391,N_6213);
and U6762 (N_6762,N_5073,N_1714);
and U6763 (N_6763,N_1867,N_6044);
and U6764 (N_6764,N_267,N_4662);
and U6765 (N_6765,N_5453,N_4698);
or U6766 (N_6766,N_4810,N_2195);
xnor U6767 (N_6767,N_2451,N_5312);
and U6768 (N_6768,N_4221,N_2649);
nor U6769 (N_6769,N_3533,N_6236);
or U6770 (N_6770,N_5406,N_1232);
or U6771 (N_6771,N_5635,N_5177);
xor U6772 (N_6772,N_4279,N_613);
nand U6773 (N_6773,N_4196,N_800);
nor U6774 (N_6774,N_920,N_5565);
nand U6775 (N_6775,N_2381,N_5192);
nand U6776 (N_6776,N_2031,N_2097);
nor U6777 (N_6777,N_3479,N_5802);
or U6778 (N_6778,N_2186,N_5244);
nand U6779 (N_6779,N_6098,N_1948);
or U6780 (N_6780,N_4941,N_32);
and U6781 (N_6781,N_3291,N_345);
or U6782 (N_6782,N_922,N_5806);
or U6783 (N_6783,N_4688,N_5122);
and U6784 (N_6784,N_1571,N_990);
and U6785 (N_6785,N_694,N_4849);
nor U6786 (N_6786,N_593,N_1070);
and U6787 (N_6787,N_5466,N_330);
or U6788 (N_6788,N_1725,N_1986);
nand U6789 (N_6789,N_4298,N_5999);
and U6790 (N_6790,N_323,N_3113);
and U6791 (N_6791,N_3109,N_1094);
xor U6792 (N_6792,N_3102,N_3258);
xnor U6793 (N_6793,N_2075,N_5403);
xor U6794 (N_6794,N_3971,N_2804);
and U6795 (N_6795,N_2539,N_5976);
xnor U6796 (N_6796,N_5512,N_3084);
nor U6797 (N_6797,N_3787,N_1376);
xor U6798 (N_6798,N_2587,N_4503);
nand U6799 (N_6799,N_3538,N_5130);
or U6800 (N_6800,N_5542,N_3628);
and U6801 (N_6801,N_3557,N_5431);
nor U6802 (N_6802,N_5270,N_3711);
xnor U6803 (N_6803,N_5549,N_3798);
nor U6804 (N_6804,N_5207,N_2377);
nor U6805 (N_6805,N_3767,N_2887);
and U6806 (N_6806,N_4837,N_2057);
and U6807 (N_6807,N_852,N_4110);
and U6808 (N_6808,N_6033,N_192);
or U6809 (N_6809,N_3956,N_23);
xor U6810 (N_6810,N_3677,N_4829);
or U6811 (N_6811,N_888,N_3178);
and U6812 (N_6812,N_5012,N_6111);
xnor U6813 (N_6813,N_3653,N_2778);
and U6814 (N_6814,N_206,N_732);
xor U6815 (N_6815,N_2735,N_4274);
nand U6816 (N_6816,N_5861,N_4275);
and U6817 (N_6817,N_4859,N_3930);
xnor U6818 (N_6818,N_544,N_70);
xor U6819 (N_6819,N_862,N_2584);
nand U6820 (N_6820,N_3404,N_5300);
nand U6821 (N_6821,N_2017,N_2882);
and U6822 (N_6822,N_1410,N_4928);
or U6823 (N_6823,N_1596,N_789);
or U6824 (N_6824,N_1262,N_5155);
nand U6825 (N_6825,N_4023,N_6171);
nor U6826 (N_6826,N_654,N_791);
and U6827 (N_6827,N_1429,N_3296);
nand U6828 (N_6828,N_3446,N_4760);
nand U6829 (N_6829,N_771,N_4920);
or U6830 (N_6830,N_5472,N_4419);
and U6831 (N_6831,N_6206,N_4775);
nand U6832 (N_6832,N_938,N_264);
or U6833 (N_6833,N_3502,N_4816);
nor U6834 (N_6834,N_5779,N_6061);
and U6835 (N_6835,N_489,N_1737);
nand U6836 (N_6836,N_2294,N_3865);
nor U6837 (N_6837,N_174,N_3508);
nand U6838 (N_6838,N_4782,N_4375);
nand U6839 (N_6839,N_2280,N_1995);
xnor U6840 (N_6840,N_2407,N_526);
nand U6841 (N_6841,N_4681,N_5765);
or U6842 (N_6842,N_2483,N_1778);
and U6843 (N_6843,N_1683,N_17);
nor U6844 (N_6844,N_6122,N_582);
nand U6845 (N_6845,N_2138,N_5347);
nor U6846 (N_6846,N_2614,N_842);
nor U6847 (N_6847,N_2144,N_4854);
nand U6848 (N_6848,N_2690,N_1182);
or U6849 (N_6849,N_1256,N_5922);
nand U6850 (N_6850,N_2061,N_540);
xor U6851 (N_6851,N_6086,N_967);
or U6852 (N_6852,N_1668,N_2425);
nand U6853 (N_6853,N_824,N_1300);
or U6854 (N_6854,N_4602,N_4180);
xor U6855 (N_6855,N_503,N_1346);
nand U6856 (N_6856,N_1606,N_1424);
or U6857 (N_6857,N_4484,N_3916);
nand U6858 (N_6858,N_3175,N_5187);
or U6859 (N_6859,N_5563,N_4708);
xor U6860 (N_6860,N_4988,N_4265);
nand U6861 (N_6861,N_4437,N_983);
and U6862 (N_6862,N_6063,N_891);
nor U6863 (N_6863,N_322,N_2707);
or U6864 (N_6864,N_2210,N_5254);
or U6865 (N_6865,N_2782,N_2258);
nor U6866 (N_6866,N_2114,N_1642);
and U6867 (N_6867,N_2960,N_886);
nor U6868 (N_6868,N_6030,N_4636);
nor U6869 (N_6869,N_827,N_2936);
nor U6870 (N_6870,N_3320,N_3424);
nor U6871 (N_6871,N_5978,N_713);
and U6872 (N_6872,N_1442,N_3813);
and U6873 (N_6873,N_4226,N_3236);
xnor U6874 (N_6874,N_5215,N_3606);
and U6875 (N_6875,N_147,N_3492);
nor U6876 (N_6876,N_3612,N_2156);
nor U6877 (N_6877,N_5677,N_2536);
nand U6878 (N_6878,N_4131,N_3227);
and U6879 (N_6879,N_2299,N_5110);
and U6880 (N_6880,N_5683,N_128);
xnor U6881 (N_6881,N_5020,N_4580);
xor U6882 (N_6882,N_187,N_2147);
or U6883 (N_6883,N_1684,N_1661);
and U6884 (N_6884,N_1151,N_4235);
nand U6885 (N_6885,N_5780,N_3328);
and U6886 (N_6886,N_4851,N_3575);
xor U6887 (N_6887,N_1917,N_3054);
nand U6888 (N_6888,N_2505,N_1865);
or U6889 (N_6889,N_845,N_2745);
or U6890 (N_6890,N_2645,N_6134);
and U6891 (N_6891,N_6223,N_4827);
xor U6892 (N_6892,N_309,N_1385);
nand U6893 (N_6893,N_4390,N_3137);
nor U6894 (N_6894,N_2107,N_6193);
and U6895 (N_6895,N_319,N_1883);
nand U6896 (N_6896,N_3336,N_2944);
and U6897 (N_6897,N_4117,N_927);
xnor U6898 (N_6898,N_4284,N_2275);
and U6899 (N_6899,N_3950,N_2700);
and U6900 (N_6900,N_1489,N_5586);
nor U6901 (N_6901,N_5399,N_5210);
xnor U6902 (N_6902,N_532,N_476);
nand U6903 (N_6903,N_6186,N_467);
nor U6904 (N_6904,N_971,N_2164);
nor U6905 (N_6905,N_10,N_2557);
nand U6906 (N_6906,N_821,N_4553);
or U6907 (N_6907,N_2899,N_5708);
nor U6908 (N_6908,N_2475,N_4550);
nand U6909 (N_6909,N_4113,N_2355);
xnor U6910 (N_6910,N_4894,N_1594);
xnor U6911 (N_6911,N_1415,N_3735);
or U6912 (N_6912,N_2580,N_5665);
xnor U6913 (N_6913,N_6051,N_2448);
or U6914 (N_6914,N_2256,N_5389);
or U6915 (N_6915,N_3981,N_3563);
or U6916 (N_6916,N_5220,N_4608);
and U6917 (N_6917,N_2532,N_2756);
nor U6918 (N_6918,N_6177,N_4993);
nor U6919 (N_6919,N_4798,N_1989);
or U6920 (N_6920,N_3416,N_2113);
or U6921 (N_6921,N_1518,N_2455);
or U6922 (N_6922,N_321,N_473);
nor U6923 (N_6923,N_3633,N_3654);
and U6924 (N_6924,N_1083,N_5118);
or U6925 (N_6925,N_3085,N_5109);
nand U6926 (N_6926,N_3079,N_2378);
and U6927 (N_6927,N_4246,N_3674);
nand U6928 (N_6928,N_2274,N_498);
nand U6929 (N_6929,N_2507,N_1072);
nor U6930 (N_6930,N_6056,N_1024);
or U6931 (N_6931,N_3875,N_4138);
xor U6932 (N_6932,N_3559,N_2832);
nand U6933 (N_6933,N_4721,N_3317);
nand U6934 (N_6934,N_5947,N_460);
or U6935 (N_6935,N_4747,N_6200);
nand U6936 (N_6936,N_4712,N_3638);
or U6937 (N_6937,N_269,N_5513);
and U6938 (N_6938,N_3848,N_1258);
and U6939 (N_6939,N_2948,N_5605);
and U6940 (N_6940,N_5557,N_5979);
or U6941 (N_6941,N_5030,N_5647);
and U6942 (N_6942,N_1125,N_3995);
nor U6943 (N_6943,N_1950,N_2406);
or U6944 (N_6944,N_76,N_11);
or U6945 (N_6945,N_438,N_4711);
or U6946 (N_6946,N_162,N_2698);
nand U6947 (N_6947,N_1881,N_4186);
nand U6948 (N_6948,N_1787,N_2192);
nor U6949 (N_6949,N_5358,N_1136);
nand U6950 (N_6950,N_566,N_4710);
nand U6951 (N_6951,N_2576,N_3362);
and U6952 (N_6952,N_4511,N_3727);
xor U6953 (N_6953,N_991,N_4368);
nor U6954 (N_6954,N_1195,N_986);
nor U6955 (N_6955,N_3045,N_6192);
nor U6956 (N_6956,N_2020,N_4672);
nand U6957 (N_6957,N_3894,N_2531);
nor U6958 (N_6958,N_2285,N_4402);
nor U6959 (N_6959,N_429,N_5603);
nor U6960 (N_6960,N_3182,N_660);
xor U6961 (N_6961,N_2931,N_5019);
or U6962 (N_6962,N_1886,N_607);
and U6963 (N_6963,N_539,N_5592);
and U6964 (N_6964,N_4663,N_5342);
nor U6965 (N_6965,N_696,N_4014);
nand U6966 (N_6966,N_5865,N_2160);
and U6967 (N_6967,N_2787,N_3820);
nor U6968 (N_6968,N_1430,N_2737);
or U6969 (N_6969,N_5653,N_4294);
or U6970 (N_6970,N_5419,N_4744);
nor U6971 (N_6971,N_5863,N_4840);
nor U6972 (N_6972,N_2478,N_5304);
nor U6973 (N_6973,N_5026,N_2496);
or U6974 (N_6974,N_5521,N_5853);
nor U6975 (N_6975,N_3595,N_5214);
or U6976 (N_6976,N_4299,N_256);
or U6977 (N_6977,N_636,N_5124);
xnor U6978 (N_6978,N_4800,N_4912);
nor U6979 (N_6979,N_5097,N_3072);
xnor U6980 (N_6980,N_392,N_6107);
nor U6981 (N_6981,N_2419,N_1933);
and U6982 (N_6982,N_3385,N_5368);
and U6983 (N_6983,N_1546,N_5685);
and U6984 (N_6984,N_781,N_4614);
or U6985 (N_6985,N_308,N_1002);
nor U6986 (N_6986,N_3782,N_787);
xnor U6987 (N_6987,N_5852,N_3354);
nor U6988 (N_6988,N_247,N_1068);
nand U6989 (N_6989,N_5343,N_6048);
xnor U6990 (N_6990,N_4192,N_6152);
or U6991 (N_6991,N_5381,N_2978);
and U6992 (N_6992,N_3234,N_4365);
nor U6993 (N_6993,N_3997,N_782);
xnor U6994 (N_6994,N_2793,N_212);
or U6995 (N_6995,N_2127,N_263);
nor U6996 (N_6996,N_2858,N_5913);
nand U6997 (N_6997,N_3907,N_2206);
or U6998 (N_6998,N_531,N_5813);
xor U6999 (N_6999,N_1713,N_5963);
and U7000 (N_7000,N_1666,N_653);
or U7001 (N_7001,N_110,N_1893);
xor U7002 (N_7002,N_4357,N_1437);
and U7003 (N_7003,N_3090,N_1408);
nor U7004 (N_7004,N_795,N_2784);
or U7005 (N_7005,N_3111,N_2162);
xnor U7006 (N_7006,N_5001,N_3504);
nor U7007 (N_7007,N_2200,N_3936);
nand U7008 (N_7008,N_5599,N_3698);
and U7009 (N_7009,N_2867,N_1187);
xnor U7010 (N_7010,N_3986,N_3873);
nand U7011 (N_7011,N_2315,N_2393);
nand U7012 (N_7012,N_3862,N_3806);
and U7013 (N_7013,N_3485,N_6015);
and U7014 (N_7014,N_417,N_4530);
xnor U7015 (N_7015,N_3517,N_3770);
nand U7016 (N_7016,N_2327,N_2550);
xor U7017 (N_7017,N_2014,N_2424);
and U7018 (N_7018,N_5642,N_1503);
xor U7019 (N_7019,N_4945,N_2444);
nand U7020 (N_7020,N_879,N_5299);
nand U7021 (N_7021,N_1330,N_2522);
xor U7022 (N_7022,N_4054,N_1751);
xor U7023 (N_7023,N_4616,N_2413);
xnor U7024 (N_7024,N_2796,N_595);
nand U7025 (N_7025,N_4718,N_1061);
nand U7026 (N_7026,N_5477,N_1833);
and U7027 (N_7027,N_4491,N_5776);
nor U7028 (N_7028,N_4626,N_2726);
nand U7029 (N_7029,N_2783,N_5084);
xnor U7030 (N_7030,N_4027,N_797);
nand U7031 (N_7031,N_3105,N_4373);
or U7032 (N_7032,N_780,N_3957);
or U7033 (N_7033,N_4254,N_2733);
or U7034 (N_7034,N_5626,N_4570);
or U7035 (N_7035,N_4979,N_5588);
nand U7036 (N_7036,N_3522,N_3834);
nand U7037 (N_7037,N_2249,N_436);
nand U7038 (N_7038,N_379,N_2150);
nor U7039 (N_7039,N_6124,N_1332);
nand U7040 (N_7040,N_1191,N_5539);
nand U7041 (N_7041,N_5621,N_3390);
and U7042 (N_7042,N_4784,N_1808);
xnor U7043 (N_7043,N_6017,N_472);
nand U7044 (N_7044,N_3103,N_3356);
nor U7045 (N_7045,N_5896,N_3108);
nor U7046 (N_7046,N_69,N_1565);
and U7047 (N_7047,N_5769,N_662);
xnor U7048 (N_7048,N_2251,N_802);
xnor U7049 (N_7049,N_1540,N_2289);
nand U7050 (N_7050,N_2293,N_5656);
nor U7051 (N_7051,N_3418,N_3852);
or U7052 (N_7052,N_4949,N_331);
xor U7053 (N_7053,N_1526,N_5502);
nor U7054 (N_7054,N_4643,N_4005);
xnor U7055 (N_7055,N_4329,N_4610);
xor U7056 (N_7056,N_1135,N_4678);
nor U7057 (N_7057,N_5894,N_4188);
or U7058 (N_7058,N_2914,N_1019);
or U7059 (N_7059,N_1365,N_4621);
and U7060 (N_7060,N_5875,N_5140);
or U7061 (N_7061,N_2639,N_1941);
nand U7062 (N_7062,N_4422,N_2493);
nand U7063 (N_7063,N_4343,N_1960);
xnor U7064 (N_7064,N_5421,N_2770);
or U7065 (N_7065,N_260,N_3378);
nor U7066 (N_7066,N_1939,N_4510);
and U7067 (N_7067,N_1229,N_5189);
xnor U7068 (N_7068,N_5649,N_1821);
and U7069 (N_7069,N_3462,N_4362);
or U7070 (N_7070,N_5695,N_895);
nor U7071 (N_7071,N_2990,N_1112);
and U7072 (N_7072,N_846,N_2313);
and U7073 (N_7073,N_2434,N_3407);
or U7074 (N_7074,N_4563,N_3055);
xor U7075 (N_7075,N_49,N_5715);
or U7076 (N_7076,N_18,N_2502);
nand U7077 (N_7077,N_6096,N_748);
xor U7078 (N_7078,N_5279,N_1982);
or U7079 (N_7079,N_1453,N_194);
xor U7080 (N_7080,N_3169,N_2653);
and U7081 (N_7081,N_1796,N_4874);
xor U7082 (N_7082,N_1891,N_961);
nand U7083 (N_7083,N_4322,N_600);
xnor U7084 (N_7084,N_2091,N_724);
or U7085 (N_7085,N_5671,N_4019);
xnor U7086 (N_7086,N_3759,N_3443);
and U7087 (N_7087,N_5749,N_2041);
nor U7088 (N_7088,N_5768,N_2198);
nor U7089 (N_7089,N_5227,N_3007);
xnor U7090 (N_7090,N_5864,N_4377);
nand U7091 (N_7091,N_1863,N_5750);
or U7092 (N_7092,N_4777,N_2814);
or U7093 (N_7093,N_3704,N_1564);
nor U7094 (N_7094,N_3176,N_4615);
xnor U7095 (N_7095,N_3681,N_710);
or U7096 (N_7096,N_204,N_3900);
xnor U7097 (N_7097,N_6132,N_6208);
nand U7098 (N_7098,N_1216,N_62);
or U7099 (N_7099,N_1380,N_4986);
or U7100 (N_7100,N_286,N_5843);
xnor U7101 (N_7101,N_1967,N_482);
or U7102 (N_7102,N_5625,N_4304);
or U7103 (N_7103,N_875,N_5197);
and U7104 (N_7104,N_4490,N_4669);
and U7105 (N_7105,N_1400,N_5426);
nor U7106 (N_7106,N_5313,N_4834);
or U7107 (N_7107,N_1792,N_3642);
xnor U7108 (N_7108,N_2304,N_5025);
nand U7109 (N_7109,N_1656,N_565);
nor U7110 (N_7110,N_4826,N_737);
xnor U7111 (N_7111,N_2912,N_6142);
nand U7112 (N_7112,N_353,N_248);
or U7113 (N_7113,N_1250,N_5325);
nand U7114 (N_7114,N_2662,N_5957);
or U7115 (N_7115,N_5452,N_5591);
nand U7116 (N_7116,N_6248,N_4647);
nand U7117 (N_7117,N_5165,N_1428);
and U7118 (N_7118,N_1144,N_339);
xor U7119 (N_7119,N_34,N_4952);
or U7120 (N_7120,N_5003,N_4984);
and U7121 (N_7121,N_5888,N_2245);
and U7122 (N_7122,N_4423,N_1637);
nand U7123 (N_7123,N_313,N_1521);
nand U7124 (N_7124,N_6215,N_5351);
nor U7125 (N_7125,N_1536,N_2719);
or U7126 (N_7126,N_1709,N_5713);
nor U7127 (N_7127,N_3391,N_4115);
and U7128 (N_7128,N_3756,N_4340);
and U7129 (N_7129,N_4046,N_5470);
xor U7130 (N_7130,N_5921,N_3180);
or U7131 (N_7131,N_2361,N_3426);
and U7132 (N_7132,N_485,N_1452);
and U7133 (N_7133,N_3969,N_6211);
or U7134 (N_7134,N_3585,N_1004);
and U7135 (N_7135,N_4652,N_5320);
and U7136 (N_7136,N_2970,N_4017);
nor U7137 (N_7137,N_2353,N_3669);
nand U7138 (N_7138,N_304,N_1977);
nand U7139 (N_7139,N_3115,N_4120);
nor U7140 (N_7140,N_4465,N_439);
nor U7141 (N_7141,N_3623,N_4291);
xnor U7142 (N_7142,N_915,N_5334);
nor U7143 (N_7143,N_6138,N_806);
nand U7144 (N_7144,N_550,N_2099);
xor U7145 (N_7145,N_3839,N_5129);
xnor U7146 (N_7146,N_3906,N_4994);
nor U7147 (N_7147,N_3217,N_1451);
xnor U7148 (N_7148,N_4222,N_521);
nand U7149 (N_7149,N_909,N_4081);
or U7150 (N_7150,N_3948,N_881);
nand U7151 (N_7151,N_20,N_884);
nand U7152 (N_7152,N_3931,N_2884);
or U7153 (N_7153,N_5613,N_4517);
or U7154 (N_7154,N_779,N_3159);
nor U7155 (N_7155,N_3174,N_4366);
xnor U7156 (N_7156,N_3350,N_3005);
or U7157 (N_7157,N_2239,N_5391);
or U7158 (N_7158,N_3793,N_3908);
nor U7159 (N_7159,N_2920,N_4389);
xor U7160 (N_7160,N_2855,N_2347);
and U7161 (N_7161,N_1896,N_5105);
nor U7162 (N_7162,N_1123,N_5523);
and U7163 (N_7163,N_1748,N_2901);
xnor U7164 (N_7164,N_77,N_4414);
nand U7165 (N_7165,N_2375,N_3879);
nor U7166 (N_7166,N_2961,N_4258);
nand U7167 (N_7167,N_942,N_441);
xnor U7168 (N_7168,N_5068,N_2615);
xnor U7169 (N_7169,N_3562,N_6026);
nor U7170 (N_7170,N_2050,N_6049);
xnor U7171 (N_7171,N_2473,N_333);
nor U7172 (N_7172,N_2069,N_5719);
or U7173 (N_7173,N_754,N_5436);
nor U7174 (N_7174,N_3038,N_3899);
xor U7175 (N_7175,N_2546,N_1045);
or U7176 (N_7176,N_3342,N_796);
nand U7177 (N_7177,N_2972,N_1770);
or U7178 (N_7178,N_3167,N_475);
and U7179 (N_7179,N_5633,N_4551);
xnor U7180 (N_7180,N_1120,N_362);
nand U7181 (N_7181,N_358,N_1999);
or U7182 (N_7182,N_4758,N_2809);
xor U7183 (N_7183,N_3847,N_601);
or U7184 (N_7184,N_3662,N_1698);
nor U7185 (N_7185,N_2351,N_618);
nor U7186 (N_7186,N_208,N_434);
xor U7187 (N_7187,N_841,N_3565);
nand U7188 (N_7188,N_1931,N_1008);
nor U7189 (N_7189,N_259,N_4730);
or U7190 (N_7190,N_3136,N_2980);
nand U7191 (N_7191,N_4243,N_4560);
or U7192 (N_7192,N_1097,N_1213);
xnor U7193 (N_7193,N_2907,N_5854);
nand U7194 (N_7194,N_327,N_1416);
xnor U7195 (N_7195,N_3225,N_3526);
nor U7196 (N_7196,N_1846,N_373);
nand U7197 (N_7197,N_1037,N_2812);
and U7198 (N_7198,N_501,N_85);
xnor U7199 (N_7199,N_376,N_1411);
and U7200 (N_7200,N_2957,N_2552);
nor U7201 (N_7201,N_1449,N_254);
nand U7202 (N_7202,N_4376,N_5891);
nor U7203 (N_7203,N_3447,N_3622);
xor U7204 (N_7204,N_1814,N_413);
nand U7205 (N_7205,N_5005,N_251);
xnor U7206 (N_7206,N_5293,N_1899);
and U7207 (N_7207,N_1898,N_4455);
xor U7208 (N_7208,N_5483,N_1895);
or U7209 (N_7209,N_4701,N_3222);
or U7210 (N_7210,N_3001,N_6179);
xor U7211 (N_7211,N_2900,N_4342);
nor U7212 (N_7212,N_3953,N_4917);
xnor U7213 (N_7213,N_5036,N_4053);
nor U7214 (N_7214,N_517,N_1364);
xor U7215 (N_7215,N_2131,N_2811);
nor U7216 (N_7216,N_3733,N_1295);
or U7217 (N_7217,N_5908,N_627);
nor U7218 (N_7218,N_262,N_5654);
nand U7219 (N_7219,N_2829,N_5341);
and U7220 (N_7220,N_1077,N_214);
and U7221 (N_7221,N_5693,N_3315);
nor U7222 (N_7222,N_1652,N_693);
nand U7223 (N_7223,N_916,N_984);
or U7224 (N_7224,N_1695,N_288);
and U7225 (N_7225,N_459,N_3963);
nand U7226 (N_7226,N_5728,N_4101);
or U7227 (N_7227,N_4540,N_1689);
or U7228 (N_7228,N_3112,N_5029);
nor U7229 (N_7229,N_5205,N_2610);
and U7230 (N_7230,N_6140,N_1188);
or U7231 (N_7231,N_4026,N_5720);
xnor U7232 (N_7232,N_381,N_2238);
xnor U7233 (N_7233,N_5940,N_1040);
nor U7234 (N_7234,N_969,N_3496);
or U7235 (N_7235,N_3276,N_340);
or U7236 (N_7236,N_5567,N_5186);
nor U7237 (N_7237,N_52,N_4405);
nand U7238 (N_7238,N_337,N_2819);
and U7239 (N_7239,N_4349,N_3667);
xnor U7240 (N_7240,N_3684,N_5002);
and U7241 (N_7241,N_5812,N_480);
or U7242 (N_7242,N_4601,N_868);
nor U7243 (N_7243,N_3070,N_3275);
xnor U7244 (N_7244,N_1163,N_1207);
or U7245 (N_7245,N_3381,N_4064);
nor U7246 (N_7246,N_324,N_1046);
xor U7247 (N_7247,N_928,N_3540);
nor U7248 (N_7248,N_1307,N_2857);
xnor U7249 (N_7249,N_4020,N_1785);
nor U7250 (N_7250,N_6022,N_6224);
or U7251 (N_7251,N_5322,N_4594);
and U7252 (N_7252,N_5914,N_847);
and U7253 (N_7253,N_1820,N_5311);
and U7254 (N_7254,N_1440,N_3154);
or U7255 (N_7255,N_826,N_2034);
or U7256 (N_7256,N_1421,N_5509);
nand U7257 (N_7257,N_465,N_2319);
and U7258 (N_7258,N_2660,N_1954);
nor U7259 (N_7259,N_4552,N_3477);
xor U7260 (N_7260,N_3494,N_2115);
nand U7261 (N_7261,N_3857,N_1082);
and U7262 (N_7262,N_1171,N_4341);
xor U7263 (N_7263,N_5363,N_5423);
or U7264 (N_7264,N_5065,N_3942);
nor U7265 (N_7265,N_4950,N_889);
xnor U7266 (N_7266,N_2705,N_231);
and U7267 (N_7267,N_4401,N_2063);
nand U7268 (N_7268,N_4004,N_3338);
or U7269 (N_7269,N_1458,N_1966);
and U7270 (N_7270,N_6099,N_4885);
xnor U7271 (N_7271,N_1052,N_5576);
nor U7272 (N_7272,N_4598,N_1753);
nand U7273 (N_7273,N_640,N_1829);
nor U7274 (N_7274,N_4908,N_2170);
nor U7275 (N_7275,N_4267,N_5841);
nor U7276 (N_7276,N_4558,N_1905);
nand U7277 (N_7277,N_311,N_1396);
nor U7278 (N_7278,N_5015,N_2865);
and U7279 (N_7279,N_4722,N_450);
nand U7280 (N_7280,N_2442,N_612);
or U7281 (N_7281,N_3994,N_2669);
xnor U7282 (N_7282,N_4306,N_481);
xor U7283 (N_7283,N_1612,N_767);
nor U7284 (N_7284,N_494,N_4603);
or U7285 (N_7285,N_4769,N_4281);
nand U7286 (N_7286,N_3425,N_1610);
xor U7287 (N_7287,N_1645,N_2693);
and U7288 (N_7288,N_3913,N_4077);
nor U7289 (N_7289,N_589,N_5353);
nand U7290 (N_7290,N_2515,N_57);
nor U7291 (N_7291,N_756,N_1890);
and U7292 (N_7292,N_3251,N_3128);
xor U7293 (N_7293,N_2484,N_3827);
and U7294 (N_7294,N_2130,N_624);
xnor U7295 (N_7295,N_377,N_6057);
or U7296 (N_7296,N_4135,N_2684);
or U7297 (N_7297,N_3597,N_1732);
and U7298 (N_7298,N_4133,N_5449);
nor U7299 (N_7299,N_2364,N_418);
nor U7300 (N_7300,N_4092,N_394);
xor U7301 (N_7301,N_4417,N_1866);
or U7302 (N_7302,N_2360,N_2330);
and U7303 (N_7303,N_5018,N_2003);
nand U7304 (N_7304,N_2331,N_4924);
and U7305 (N_7305,N_4487,N_4738);
and U7306 (N_7306,N_4907,N_4763);
nand U7307 (N_7307,N_4536,N_6007);
nor U7308 (N_7308,N_5054,N_1423);
and U7309 (N_7309,N_552,N_3799);
nand U7310 (N_7310,N_4161,N_5496);
nor U7311 (N_7311,N_58,N_3219);
xor U7312 (N_7312,N_2962,N_1159);
nand U7313 (N_7313,N_1955,N_4345);
xor U7314 (N_7314,N_3752,N_1174);
nor U7315 (N_7315,N_5302,N_42);
nor U7316 (N_7316,N_1851,N_1779);
nand U7317 (N_7317,N_5139,N_6066);
and U7318 (N_7318,N_196,N_2445);
xor U7319 (N_7319,N_3068,N_703);
xor U7320 (N_7320,N_2898,N_2449);
nor U7321 (N_7321,N_646,N_3702);
nor U7322 (N_7322,N_2659,N_5183);
nand U7323 (N_7323,N_2762,N_4838);
and U7324 (N_7324,N_6198,N_4831);
and U7325 (N_7325,N_5088,N_3567);
or U7326 (N_7326,N_1311,N_1476);
or U7327 (N_7327,N_5673,N_4149);
nand U7328 (N_7328,N_2619,N_218);
xor U7329 (N_7329,N_907,N_574);
nand U7330 (N_7330,N_2287,N_6064);
nor U7331 (N_7331,N_4631,N_3532);
xor U7332 (N_7332,N_4713,N_4887);
xor U7333 (N_7333,N_1537,N_5962);
or U7334 (N_7334,N_2088,N_2676);
nor U7335 (N_7335,N_2585,N_3285);
or U7336 (N_7336,N_3791,N_283);
nand U7337 (N_7337,N_5774,N_5730);
or U7338 (N_7338,N_1080,N_950);
and U7339 (N_7339,N_6071,N_2874);
and U7340 (N_7340,N_4420,N_4861);
or U7341 (N_7341,N_397,N_1658);
or U7342 (N_7342,N_2006,N_1036);
nand U7343 (N_7343,N_3572,N_1314);
xor U7344 (N_7344,N_1399,N_4444);
and U7345 (N_7345,N_2835,N_1255);
nor U7346 (N_7346,N_3445,N_2426);
or U7347 (N_7347,N_3832,N_4532);
nor U7348 (N_7348,N_5460,N_623);
or U7349 (N_7349,N_5543,N_2112);
and U7350 (N_7350,N_6187,N_3661);
and U7351 (N_7351,N_1375,N_3132);
or U7352 (N_7352,N_3694,N_5757);
nor U7353 (N_7353,N_6156,N_5932);
xnor U7354 (N_7354,N_1039,N_4862);
and U7355 (N_7355,N_4111,N_1238);
or U7356 (N_7356,N_5237,N_4773);
or U7357 (N_7357,N_496,N_555);
xnor U7358 (N_7358,N_4723,N_1573);
nand U7359 (N_7359,N_3069,N_3757);
and U7360 (N_7360,N_3996,N_2999);
nand U7361 (N_7361,N_500,N_4571);
and U7362 (N_7362,N_1859,N_954);
xnor U7363 (N_7363,N_3394,N_4452);
nor U7364 (N_7364,N_3905,N_5415);
xnor U7365 (N_7365,N_2262,N_5792);
and U7366 (N_7366,N_5023,N_3918);
and U7367 (N_7367,N_2324,N_249);
nor U7368 (N_7368,N_3789,N_2981);
xor U7369 (N_7369,N_3925,N_3734);
xnor U7370 (N_7370,N_3592,N_4280);
nand U7371 (N_7371,N_3998,N_4137);
nand U7372 (N_7372,N_4821,N_853);
nor U7373 (N_7373,N_6080,N_126);
nand U7374 (N_7374,N_5385,N_235);
or U7375 (N_7375,N_246,N_1122);
nand U7376 (N_7376,N_6221,N_2225);
and U7377 (N_7377,N_4461,N_1680);
xnor U7378 (N_7378,N_5387,N_176);
xor U7379 (N_7379,N_3569,N_6031);
nand U7380 (N_7380,N_1850,N_4565);
nand U7381 (N_7381,N_177,N_1597);
nand U7382 (N_7382,N_3198,N_4537);
xnor U7383 (N_7383,N_1297,N_2196);
xor U7384 (N_7384,N_1738,N_2085);
xor U7385 (N_7385,N_1075,N_3892);
xnor U7386 (N_7386,N_1107,N_1879);
nand U7387 (N_7387,N_2797,N_5758);
xor U7388 (N_7388,N_3074,N_5602);
and U7389 (N_7389,N_3878,N_1224);
or U7390 (N_7390,N_1544,N_556);
and U7391 (N_7391,N_5924,N_4533);
and U7392 (N_7392,N_5204,N_280);
and U7393 (N_7393,N_1772,N_338);
nand U7394 (N_7394,N_2840,N_1551);
and U7395 (N_7395,N_4745,N_1840);
nand U7396 (N_7396,N_4561,N_3489);
xnor U7397 (N_7397,N_527,N_2607);
nor U7398 (N_7398,N_3372,N_3280);
xor U7399 (N_7399,N_2759,N_2116);
and U7400 (N_7400,N_3065,N_1760);
or U7401 (N_7401,N_2191,N_5862);
nor U7402 (N_7402,N_2543,N_3018);
and U7403 (N_7403,N_3776,N_4269);
and U7404 (N_7404,N_3580,N_581);
and U7405 (N_7405,N_1694,N_2180);
or U7406 (N_7406,N_5632,N_3926);
nand U7407 (N_7407,N_5773,N_6217);
xnor U7408 (N_7408,N_3549,N_643);
or U7409 (N_7409,N_4021,N_4823);
nand U7410 (N_7410,N_3230,N_2237);
nand U7411 (N_7411,N_3311,N_2930);
nor U7412 (N_7412,N_5131,N_5224);
xnor U7413 (N_7413,N_2094,N_5624);
xnor U7414 (N_7414,N_5532,N_6175);
nor U7415 (N_7415,N_5052,N_3548);
and U7416 (N_7416,N_641,N_2093);
and U7417 (N_7417,N_2437,N_412);
nand U7418 (N_7418,N_2860,N_4286);
or U7419 (N_7419,N_6028,N_2126);
nand U7420 (N_7420,N_1682,N_1312);
nand U7421 (N_7421,N_4739,N_5236);
nor U7422 (N_7422,N_179,N_3361);
nor U7423 (N_7423,N_2356,N_3388);
xnor U7424 (N_7424,N_677,N_5997);
nor U7425 (N_7425,N_210,N_530);
nand U7426 (N_7426,N_2489,N_4916);
nor U7427 (N_7427,N_2670,N_4129);
nor U7428 (N_7428,N_2342,N_546);
or U7429 (N_7429,N_1884,N_2277);
xor U7430 (N_7430,N_404,N_3133);
xnor U7431 (N_7431,N_6038,N_2269);
xor U7432 (N_7432,N_5388,N_4735);
xor U7433 (N_7433,N_276,N_5246);
nand U7434 (N_7434,N_3475,N_4692);
or U7435 (N_7435,N_4467,N_5681);
xor U7436 (N_7436,N_3867,N_1180);
or U7437 (N_7437,N_4088,N_5851);
or U7438 (N_7438,N_3774,N_2211);
and U7439 (N_7439,N_1360,N_5043);
nand U7440 (N_7440,N_422,N_3039);
xor U7441 (N_7441,N_6084,N_5044);
or U7442 (N_7442,N_1828,N_1649);
nand U7443 (N_7443,N_3125,N_1504);
and U7444 (N_7444,N_1936,N_56);
xor U7445 (N_7445,N_4238,N_1473);
nor U7446 (N_7446,N_1704,N_242);
and U7447 (N_7447,N_2118,N_364);
xor U7448 (N_7448,N_3783,N_3619);
and U7449 (N_7449,N_3473,N_3728);
nor U7450 (N_7450,N_1478,N_4600);
or U7451 (N_7451,N_5401,N_3511);
nor U7452 (N_7452,N_154,N_1981);
nand U7453 (N_7453,N_369,N_5241);
xor U7454 (N_7454,N_3240,N_5944);
or U7455 (N_7455,N_458,N_5771);
nor U7456 (N_7456,N_1117,N_3983);
nand U7457 (N_7457,N_1734,N_2443);
or U7458 (N_7458,N_3481,N_5136);
xnor U7459 (N_7459,N_6087,N_2433);
or U7460 (N_7460,N_6074,N_6165);
or U7461 (N_7461,N_2744,N_3984);
xnor U7462 (N_7462,N_5511,N_202);
nor U7463 (N_7463,N_453,N_1480);
or U7464 (N_7464,N_1252,N_1726);
xnor U7465 (N_7465,N_3067,N_943);
xnor U7466 (N_7466,N_452,N_2);
nor U7467 (N_7467,N_5941,N_516);
and U7468 (N_7468,N_2595,N_885);
xor U7469 (N_7469,N_4164,N_866);
and U7470 (N_7470,N_2674,N_2971);
or U7471 (N_7471,N_2504,N_3604);
and U7472 (N_7472,N_4932,N_2749);
or U7473 (N_7473,N_3853,N_2520);
nor U7474 (N_7474,N_5080,N_84);
and U7475 (N_7475,N_2729,N_3029);
nor U7476 (N_7476,N_6078,N_4774);
and U7477 (N_7477,N_1340,N_843);
and U7478 (N_7478,N_5628,N_3578);
and U7479 (N_7479,N_4696,N_2148);
or U7480 (N_7480,N_2217,N_6118);
xnor U7481 (N_7481,N_599,N_3403);
nor U7482 (N_7482,N_5101,N_8);
xnor U7483 (N_7483,N_4287,N_3056);
nor U7484 (N_7484,N_2025,N_1324);
or U7485 (N_7485,N_2508,N_4103);
and U7486 (N_7486,N_1918,N_170);
nor U7487 (N_7487,N_437,N_3713);
or U7488 (N_7488,N_3472,N_1362);
and U7489 (N_7489,N_3245,N_6219);
nand U7490 (N_7490,N_1897,N_5382);
or U7491 (N_7491,N_5373,N_3626);
nand U7492 (N_7492,N_3505,N_3322);
nor U7493 (N_7493,N_4347,N_6214);
nor U7494 (N_7494,N_1512,N_519);
xor U7495 (N_7495,N_801,N_5296);
or U7496 (N_7496,N_755,N_5212);
nand U7497 (N_7497,N_2954,N_2142);
xor U7498 (N_7498,N_1892,N_2765);
or U7499 (N_7499,N_3561,N_2358);
and U7500 (N_7500,N_107,N_109);
nand U7501 (N_7501,N_3142,N_5476);
xnor U7502 (N_7502,N_4134,N_4);
xor U7503 (N_7503,N_5710,N_4628);
or U7504 (N_7504,N_2540,N_3110);
and U7505 (N_7505,N_6178,N_4872);
nor U7506 (N_7506,N_33,N_5235);
or U7507 (N_7507,N_155,N_3166);
and U7508 (N_7508,N_3707,N_1543);
and U7509 (N_7509,N_3024,N_213);
xnor U7510 (N_7510,N_4740,N_1023);
or U7511 (N_7511,N_163,N_2661);
nand U7512 (N_7512,N_1657,N_2153);
xor U7513 (N_7513,N_433,N_3246);
nor U7514 (N_7514,N_289,N_2652);
xnor U7515 (N_7515,N_227,N_5226);
nand U7516 (N_7516,N_551,N_1269);
and U7517 (N_7517,N_1284,N_2308);
xor U7518 (N_7518,N_4990,N_1015);
and U7519 (N_7519,N_209,N_1826);
nand U7520 (N_7520,N_1970,N_630);
or U7521 (N_7521,N_2668,N_5035);
or U7522 (N_7522,N_4897,N_4220);
xnor U7523 (N_7523,N_4677,N_2416);
or U7524 (N_7524,N_2109,N_3405);
nand U7525 (N_7525,N_2232,N_4519);
or U7526 (N_7526,N_1757,N_4155);
and U7527 (N_7527,N_4430,N_3051);
nor U7528 (N_7528,N_4309,N_1940);
nor U7529 (N_7529,N_3725,N_1563);
or U7530 (N_7530,N_3721,N_2880);
or U7531 (N_7531,N_4943,N_1029);
nor U7532 (N_7532,N_773,N_2334);
or U7533 (N_7533,N_4556,N_2810);
nor U7534 (N_7534,N_5600,N_4964);
and U7535 (N_7535,N_4871,N_5276);
nor U7536 (N_7536,N_3058,N_605);
or U7537 (N_7537,N_3710,N_772);
or U7538 (N_7538,N_1043,N_121);
nor U7539 (N_7539,N_4447,N_5644);
xor U7540 (N_7540,N_1142,N_5062);
or U7541 (N_7541,N_82,N_1847);
or U7542 (N_7542,N_4689,N_6116);
nor U7543 (N_7543,N_497,N_469);
xor U7544 (N_7544,N_2724,N_4223);
and U7545 (N_7545,N_3831,N_558);
xor U7546 (N_7546,N_5000,N_869);
xor U7547 (N_7547,N_591,N_2450);
nor U7548 (N_7548,N_6189,N_3512);
nand U7549 (N_7549,N_6201,N_1317);
and U7550 (N_7550,N_2873,N_440);
nor U7551 (N_7551,N_4936,N_2934);
nand U7552 (N_7552,N_2666,N_2438);
xnor U7553 (N_7553,N_4852,N_6065);
or U7554 (N_7554,N_2953,N_1983);
or U7555 (N_7555,N_5045,N_3670);
and U7556 (N_7556,N_5895,N_2687);
and U7557 (N_7557,N_1853,N_4379);
nor U7558 (N_7558,N_1747,N_736);
and U7559 (N_7559,N_21,N_1788);
or U7560 (N_7560,N_1617,N_2053);
nor U7561 (N_7561,N_2630,N_4574);
nand U7562 (N_7562,N_2935,N_5799);
xor U7563 (N_7563,N_2871,N_1185);
nor U7564 (N_7564,N_4501,N_6169);
and U7565 (N_7565,N_3264,N_1098);
xor U7566 (N_7566,N_2987,N_3215);
and U7567 (N_7567,N_47,N_5128);
nor U7568 (N_7568,N_191,N_3574);
nand U7569 (N_7569,N_6127,N_4311);
nor U7570 (N_7570,N_4577,N_1240);
nor U7571 (N_7571,N_1114,N_2910);
and U7572 (N_7572,N_5597,N_3744);
nor U7573 (N_7573,N_6164,N_763);
or U7574 (N_7574,N_1992,N_633);
or U7575 (N_7575,N_360,N_2273);
and U7576 (N_7576,N_4591,N_5903);
and U7577 (N_7577,N_2436,N_2664);
nor U7578 (N_7578,N_3516,N_3118);
xor U7579 (N_7579,N_1781,N_3960);
xor U7580 (N_7580,N_3210,N_30);
nand U7581 (N_7581,N_2850,N_2672);
or U7582 (N_7582,N_2740,N_702);
and U7583 (N_7583,N_4153,N_1219);
xor U7584 (N_7584,N_4156,N_3785);
and U7585 (N_7585,N_2104,N_5770);
nor U7586 (N_7586,N_4480,N_4297);
xnor U7587 (N_7587,N_315,N_2746);
and U7588 (N_7588,N_2151,N_856);
and U7589 (N_7589,N_4607,N_211);
nand U7590 (N_7590,N_4022,N_6184);
xor U7591 (N_7591,N_1178,N_5150);
or U7592 (N_7592,N_4442,N_4301);
nand U7593 (N_7593,N_4754,N_2199);
and U7594 (N_7594,N_3571,N_5569);
and U7595 (N_7595,N_3334,N_5135);
and U7596 (N_7596,N_1885,N_2992);
xor U7597 (N_7597,N_1431,N_2165);
nand U7598 (N_7598,N_3644,N_1621);
and U7599 (N_7599,N_2311,N_5856);
nand U7600 (N_7600,N_4114,N_4612);
nand U7601 (N_7601,N_1858,N_5053);
nor U7602 (N_7602,N_758,N_698);
nand U7603 (N_7603,N_731,N_4128);
nand U7604 (N_7604,N_5936,N_195);
and U7605 (N_7605,N_1854,N_642);
or U7606 (N_7606,N_2575,N_4890);
nand U7607 (N_7607,N_1745,N_5169);
or U7608 (N_7608,N_296,N_2022);
or U7609 (N_7609,N_1461,N_1773);
nand U7610 (N_7610,N_1225,N_1092);
or U7611 (N_7611,N_1670,N_4729);
and U7612 (N_7612,N_3620,N_1470);
nand U7613 (N_7613,N_4208,N_1249);
and U7614 (N_7614,N_1140,N_1669);
nand U7615 (N_7615,N_4413,N_6110);
nor U7616 (N_7616,N_487,N_4165);
xnor U7617 (N_7617,N_2994,N_2231);
xor U7618 (N_7618,N_4534,N_3468);
or U7619 (N_7619,N_136,N_2932);
xnor U7620 (N_7620,N_957,N_1358);
nor U7621 (N_7621,N_5099,N_2208);
xor U7622 (N_7622,N_3119,N_2246);
and U7623 (N_7623,N_396,N_778);
nor U7624 (N_7624,N_4518,N_3442);
or U7625 (N_7625,N_674,N_1338);
xor U7626 (N_7626,N_2157,N_2824);
xor U7627 (N_7627,N_5222,N_2890);
and U7628 (N_7628,N_61,N_4939);
nor U7629 (N_7629,N_5027,N_2675);
nor U7630 (N_7630,N_5589,N_4199);
or U7631 (N_7631,N_6091,N_4566);
nand U7632 (N_7632,N_2560,N_5463);
or U7633 (N_7633,N_5827,N_3441);
or U7634 (N_7634,N_1793,N_4460);
nand U7635 (N_7635,N_2902,N_3);
xor U7636 (N_7636,N_424,N_5315);
nand U7637 (N_7637,N_3161,N_4302);
nor U7638 (N_7638,N_3233,N_834);
nand U7639 (N_7639,N_5294,N_5618);
and U7640 (N_7640,N_1475,N_2975);
nor U7641 (N_7641,N_695,N_4378);
or U7642 (N_7642,N_4024,N_5412);
and U7643 (N_7643,N_6013,N_2457);
or U7644 (N_7644,N_92,N_6016);
or U7645 (N_7645,N_1217,N_3057);
or U7646 (N_7646,N_2601,N_2622);
or U7647 (N_7647,N_4228,N_1342);
nand U7648 (N_7648,N_4958,N_199);
or U7649 (N_7649,N_5764,N_5795);
or U7650 (N_7650,N_4451,N_5196);
xor U7651 (N_7651,N_657,N_2514);
and U7652 (N_7652,N_4637,N_457);
and U7653 (N_7653,N_2715,N_2010);
or U7654 (N_7654,N_4883,N_3943);
nand U7655 (N_7655,N_3430,N_5885);
nand U7656 (N_7656,N_4197,N_5126);
xor U7657 (N_7657,N_2282,N_3329);
or U7658 (N_7658,N_2598,N_3751);
and U7659 (N_7659,N_124,N_104);
or U7660 (N_7660,N_5840,N_6046);
nand U7661 (N_7661,N_1348,N_3377);
and U7662 (N_7662,N_1394,N_3939);
nand U7663 (N_7663,N_4969,N_1795);
nor U7664 (N_7664,N_3794,N_1065);
nand U7665 (N_7665,N_2817,N_1717);
or U7666 (N_7666,N_3833,N_5514);
nor U7667 (N_7667,N_3527,N_4756);
and U7668 (N_7668,N_79,N_3436);
and U7669 (N_7669,N_935,N_2423);
and U7670 (N_7670,N_2773,N_357);
xnor U7671 (N_7671,N_1101,N_2896);
or U7672 (N_7672,N_5154,N_172);
nand U7673 (N_7673,N_1943,N_3835);
xnor U7674 (N_7674,N_2529,N_4328);
or U7675 (N_7675,N_4214,N_738);
nand U7676 (N_7676,N_4436,N_3249);
nand U7677 (N_7677,N_1740,N_2286);
nand U7678 (N_7678,N_3097,N_5216);
nand U7679 (N_7679,N_2713,N_1477);
or U7680 (N_7680,N_219,N_3214);
and U7681 (N_7681,N_1752,N_3365);
and U7682 (N_7682,N_753,N_3903);
nor U7683 (N_7683,N_4317,N_5014);
and U7684 (N_7684,N_5545,N_4100);
xor U7685 (N_7685,N_1259,N_3503);
or U7686 (N_7686,N_5832,N_946);
and U7687 (N_7687,N_1014,N_5553);
nand U7688 (N_7688,N_4525,N_3053);
or U7689 (N_7689,N_1809,N_2643);
xor U7690 (N_7690,N_5704,N_4000);
nand U7691 (N_7691,N_2446,N_4331);
nand U7692 (N_7692,N_5095,N_6000);
nand U7693 (N_7693,N_2411,N_1782);
and U7694 (N_7694,N_840,N_936);
or U7695 (N_7695,N_279,N_1910);
or U7696 (N_7696,N_5550,N_1634);
or U7697 (N_7697,N_3016,N_2337);
nor U7698 (N_7698,N_19,N_1553);
nand U7699 (N_7699,N_1285,N_5744);
nand U7700 (N_7700,N_2788,N_4168);
xnor U7701 (N_7701,N_860,N_3295);
xnor U7702 (N_7702,N_1506,N_3881);
nand U7703 (N_7703,N_2974,N_1110);
xor U7704 (N_7704,N_6133,N_2288);
and U7705 (N_7705,N_5339,N_3568);
nor U7706 (N_7706,N_65,N_2089);
xor U7707 (N_7707,N_2803,N_2847);
and U7708 (N_7708,N_1912,N_974);
nand U7709 (N_7709,N_5170,N_5652);
nand U7710 (N_7710,N_1806,N_5826);
nor U7711 (N_7711,N_524,N_663);
and U7712 (N_7712,N_4080,N_3253);
or U7713 (N_7713,N_1402,N_1558);
nand U7714 (N_7714,N_5481,N_6227);
nor U7715 (N_7715,N_4832,N_5250);
and U7716 (N_7716,N_632,N_3017);
and U7717 (N_7717,N_3465,N_5981);
and U7718 (N_7718,N_1903,N_4227);
nor U7719 (N_7719,N_2919,N_3992);
and U7720 (N_7720,N_2367,N_4676);
or U7721 (N_7721,N_557,N_3768);
nor U7722 (N_7722,N_1945,N_2362);
nand U7723 (N_7723,N_5727,N_5179);
or U7724 (N_7724,N_536,N_4865);
xnor U7725 (N_7725,N_1439,N_2597);
or U7726 (N_7726,N_4801,N_2298);
or U7727 (N_7727,N_1377,N_4578);
nand U7728 (N_7728,N_2491,N_6036);
or U7729 (N_7729,N_2720,N_4808);
nor U7730 (N_7730,N_817,N_1013);
and U7731 (N_7731,N_1710,N_4190);
xnor U7732 (N_7732,N_2462,N_1200);
or U7733 (N_7733,N_2570,N_4038);
xor U7734 (N_7734,N_41,N_1248);
xnor U7735 (N_7735,N_3896,N_4256);
and U7736 (N_7736,N_2679,N_4833);
or U7737 (N_7737,N_5763,N_2955);
and U7738 (N_7738,N_4853,N_3401);
or U7739 (N_7739,N_4079,N_2701);
nand U7740 (N_7740,N_5634,N_5522);
nand U7741 (N_7741,N_2276,N_5547);
or U7742 (N_7742,N_6095,N_171);
or U7743 (N_7743,N_1290,N_4231);
or U7744 (N_7744,N_1647,N_1595);
or U7745 (N_7745,N_807,N_241);
xnor U7746 (N_7746,N_2105,N_4705);
nor U7747 (N_7747,N_5552,N_1294);
nor U7748 (N_7748,N_1313,N_5221);
nand U7749 (N_7749,N_1622,N_4268);
and U7750 (N_7750,N_3928,N_1727);
and U7751 (N_7751,N_5160,N_3599);
nand U7752 (N_7752,N_4323,N_1667);
nor U7753 (N_7753,N_932,N_844);
nor U7754 (N_7754,N_1209,N_3909);
xor U7755 (N_7755,N_658,N_4216);
or U7756 (N_7756,N_648,N_3841);
nand U7757 (N_7757,N_3389,N_1247);
or U7758 (N_7758,N_5740,N_5384);
xnor U7759 (N_7759,N_5458,N_112);
or U7760 (N_7760,N_2513,N_6197);
and U7761 (N_7761,N_603,N_3651);
and U7762 (N_7762,N_2382,N_4087);
and U7763 (N_7763,N_3340,N_341);
nand U7764 (N_7764,N_129,N_1968);
nand U7765 (N_7765,N_3898,N_5361);
nand U7766 (N_7766,N_3173,N_3965);
xor U7767 (N_7767,N_5949,N_4090);
nand U7768 (N_7768,N_6212,N_1234);
xnor U7769 (N_7769,N_1497,N_5698);
xnor U7770 (N_7770,N_4929,N_5489);
xor U7771 (N_7771,N_2471,N_4910);
and U7772 (N_7772,N_4043,N_1501);
nor U7773 (N_7773,N_4399,N_2339);
nand U7774 (N_7774,N_1326,N_142);
nand U7775 (N_7775,N_4844,N_2644);
nor U7776 (N_7776,N_6239,N_5066);
nor U7777 (N_7777,N_5723,N_676);
and U7778 (N_7778,N_786,N_3431);
and U7779 (N_7779,N_2979,N_1454);
and U7780 (N_7780,N_2834,N_937);
nand U7781 (N_7781,N_3890,N_6245);
or U7782 (N_7782,N_3459,N_538);
nor U7783 (N_7783,N_997,N_3570);
and U7784 (N_7784,N_90,N_1172);
nand U7785 (N_7785,N_3034,N_4590);
xnor U7786 (N_7786,N_3510,N_5376);
xnor U7787 (N_7787,N_5357,N_711);
nand U7788 (N_7788,N_4576,N_2178);
nor U7789 (N_7789,N_4927,N_6202);
nand U7790 (N_7790,N_1154,N_4668);
nand U7791 (N_7791,N_4241,N_1296);
nand U7792 (N_7792,N_4426,N_5486);
or U7793 (N_7793,N_4439,N_4147);
nor U7794 (N_7794,N_6018,N_3209);
xnor U7795 (N_7795,N_4121,N_3600);
and U7796 (N_7796,N_5637,N_5838);
xnor U7797 (N_7797,N_1550,N_2688);
or U7798 (N_7798,N_15,N_5243);
nand U7799 (N_7799,N_3659,N_1529);
nand U7800 (N_7800,N_1919,N_3902);
and U7801 (N_7801,N_5048,N_5262);
or U7802 (N_7802,N_1133,N_3982);
nand U7803 (N_7803,N_1298,N_3429);
xnor U7804 (N_7804,N_3195,N_5009);
nor U7805 (N_7805,N_1426,N_2879);
nor U7806 (N_7806,N_3534,N_3737);
nand U7807 (N_7807,N_378,N_4930);
nor U7808 (N_7808,N_5682,N_995);
and U7809 (N_7809,N_4037,N_2062);
and U7810 (N_7810,N_5146,N_1137);
nand U7811 (N_7811,N_2252,N_5871);
or U7812 (N_7812,N_4360,N_5942);
and U7813 (N_7813,N_1447,N_3989);
and U7814 (N_7814,N_4846,N_1803);
and U7815 (N_7815,N_2348,N_1432);
or U7816 (N_7816,N_2801,N_4308);
nand U7817 (N_7817,N_5620,N_4212);
nor U7818 (N_7818,N_5240,N_4640);
nand U7819 (N_7819,N_2242,N_3802);
and U7820 (N_7820,N_5506,N_4012);
or U7821 (N_7821,N_1085,N_1499);
xnor U7822 (N_7822,N_3321,N_2558);
xor U7823 (N_7823,N_5494,N_370);
xnor U7824 (N_7824,N_5712,N_3593);
and U7825 (N_7825,N_1281,N_4154);
nand U7826 (N_7826,N_3229,N_5995);
and U7827 (N_7827,N_5485,N_979);
xnor U7828 (N_7828,N_4609,N_3427);
nor U7829 (N_7829,N_6034,N_185);
and U7830 (N_7830,N_5916,N_4764);
and U7831 (N_7831,N_3151,N_2408);
nor U7832 (N_7832,N_5907,N_2227);
nand U7833 (N_7833,N_5267,N_4734);
and U7834 (N_7834,N_604,N_2281);
nand U7835 (N_7835,N_2519,N_5929);
xor U7836 (N_7836,N_265,N_232);
nand U7837 (N_7837,N_561,N_4746);
xnor U7838 (N_7838,N_3269,N_5711);
xor U7839 (N_7839,N_5574,N_1780);
nor U7840 (N_7840,N_5983,N_3203);
xor U7841 (N_7841,N_5168,N_2892);
and U7842 (N_7842,N_5445,N_1001);
nand U7843 (N_7843,N_5528,N_2516);
xnor U7844 (N_7844,N_6006,N_6004);
nor U7845 (N_7845,N_4753,N_2284);
xor U7846 (N_7846,N_1807,N_2869);
and U7847 (N_7847,N_5572,N_5943);
or U7848 (N_7848,N_2021,N_3860);
or U7849 (N_7849,N_244,N_5479);
or U7850 (N_7850,N_3904,N_1810);
nor U7851 (N_7851,N_2785,N_216);
xor U7852 (N_7852,N_5960,N_5275);
and U7853 (N_7853,N_4634,N_114);
xor U7854 (N_7854,N_6183,N_2692);
nand U7855 (N_7855,N_1204,N_5442);
nand U7856 (N_7856,N_4572,N_3690);
and U7857 (N_7857,N_2390,N_614);
xnor U7858 (N_7858,N_4388,N_1894);
and U7859 (N_7859,N_514,N_4415);
and U7860 (N_7860,N_1990,N_2177);
xnor U7861 (N_7861,N_728,N_5042);
xor U7862 (N_7862,N_127,N_463);
nand U7863 (N_7863,N_6148,N_980);
xor U7864 (N_7864,N_6181,N_2845);
nor U7865 (N_7865,N_2267,N_622);
or U7866 (N_7866,N_4470,N_3116);
nor U7867 (N_7867,N_1241,N_4499);
nand U7868 (N_7868,N_3331,N_2588);
nor U7869 (N_7869,N_6158,N_2617);
nand U7870 (N_7870,N_3435,N_836);
xor U7871 (N_7871,N_959,N_4481);
or U7872 (N_7872,N_5360,N_3889);
and U7873 (N_7873,N_4107,N_410);
nor U7874 (N_7874,N_3598,N_1522);
and U7875 (N_7875,N_2640,N_3935);
or U7876 (N_7876,N_5731,N_4866);
xor U7877 (N_7877,N_4250,N_670);
or U7878 (N_7878,N_305,N_2725);
and U7879 (N_7879,N_2106,N_1459);
and U7880 (N_7880,N_5444,N_1242);
nor U7881 (N_7881,N_3501,N_3484);
nand U7882 (N_7882,N_448,N_2683);
and U7883 (N_7883,N_2702,N_1006);
nand U7884 (N_7884,N_3591,N_1465);
or U7885 (N_7885,N_88,N_5689);
and U7886 (N_7886,N_2291,N_464);
xor U7887 (N_7887,N_5091,N_2447);
xor U7888 (N_7888,N_5786,N_5669);
and U7889 (N_7889,N_2290,N_39);
or U7890 (N_7890,N_4902,N_2174);
nor U7891 (N_7891,N_3500,N_3987);
or U7892 (N_7892,N_4477,N_960);
nand U7893 (N_7893,N_1352,N_5788);
or U7894 (N_7894,N_3784,N_2682);
nor U7895 (N_7895,N_4523,N_1);
or U7896 (N_7896,N_5028,N_1822);
and U7897 (N_7897,N_2011,N_3000);
and U7898 (N_7898,N_3629,N_3888);
nand U7899 (N_7899,N_4433,N_2881);
and U7900 (N_7900,N_5116,N_4058);
and U7901 (N_7901,N_3083,N_1498);
or U7902 (N_7902,N_3031,N_5021);
nor U7903 (N_7903,N_1206,N_3170);
nand U7904 (N_7904,N_4915,N_456);
nor U7905 (N_7905,N_2510,N_513);
nor U7906 (N_7906,N_5959,N_2776);
nor U7907 (N_7907,N_5281,N_873);
or U7908 (N_7908,N_5266,N_4483);
xnor U7909 (N_7909,N_5724,N_2427);
or U7910 (N_7910,N_3375,N_4508);
xor U7911 (N_7911,N_1888,N_3231);
and U7912 (N_7912,N_1318,N_1457);
nand U7913 (N_7913,N_2422,N_1800);
nand U7914 (N_7914,N_380,N_6020);
or U7915 (N_7915,N_3347,N_6103);
or U7916 (N_7916,N_270,N_6125);
xnor U7917 (N_7917,N_822,N_3746);
xnor U7918 (N_7918,N_4977,N_130);
xnor U7919 (N_7919,N_1463,N_5367);
and U7920 (N_7920,N_4010,N_2876);
or U7921 (N_7921,N_5825,N_3914);
or U7922 (N_7922,N_1584,N_6242);
or U7923 (N_7923,N_4167,N_6243);
nand U7924 (N_7924,N_1978,N_1908);
xor U7925 (N_7925,N_5882,N_5679);
or U7926 (N_7926,N_2608,N_2181);
nand U7927 (N_7927,N_5504,N_116);
or U7928 (N_7928,N_1197,N_1692);
nor U7929 (N_7929,N_1848,N_1175);
or U7930 (N_7930,N_730,N_451);
nor U7931 (N_7931,N_1349,N_2379);
or U7932 (N_7932,N_2918,N_71);
nor U7933 (N_7933,N_2065,N_3400);
nor U7934 (N_7934,N_3650,N_3104);
nand U7935 (N_7935,N_5167,N_2428);
and U7936 (N_7936,N_828,N_228);
and U7937 (N_7937,N_5548,N_2399);
or U7938 (N_7938,N_5430,N_3589);
and U7939 (N_7939,N_4955,N_5413);
nor U7940 (N_7940,N_744,N_2292);
or U7941 (N_7941,N_4277,N_3196);
and U7942 (N_7942,N_3370,N_4295);
nand U7943 (N_7943,N_2567,N_3299);
nand U7944 (N_7944,N_1468,N_3615);
and U7945 (N_7945,N_1513,N_5354);
and U7946 (N_7946,N_4878,N_650);
xor U7947 (N_7947,N_2038,N_4660);
and U7948 (N_7948,N_1031,N_145);
nand U7949 (N_7949,N_5778,N_6005);
and U7950 (N_7950,N_1026,N_4736);
and U7951 (N_7951,N_419,N_4172);
or U7952 (N_7952,N_55,N_1994);
nor U7953 (N_7953,N_5055,N_3165);
or U7954 (N_7954,N_1273,N_1469);
or U7955 (N_7955,N_5107,N_1466);
nand U7956 (N_7956,N_4529,N_5583);
or U7957 (N_7957,N_6170,N_5499);
and U7958 (N_7958,N_1693,N_5427);
nand U7959 (N_7959,N_5490,N_6053);
nor U7960 (N_7960,N_5581,N_5703);
or U7961 (N_7961,N_3419,N_3712);
nand U7962 (N_7962,N_4975,N_2637);
and U7963 (N_7963,N_401,N_504);
or U7964 (N_7964,N_287,N_4327);
and U7965 (N_7965,N_1952,N_4157);
and U7966 (N_7966,N_387,N_5405);
xor U7967 (N_7967,N_6032,N_3263);
and U7968 (N_7968,N_3080,N_4858);
nor U7969 (N_7969,N_2500,N_5285);
and U7970 (N_7970,N_5208,N_2485);
nor U7971 (N_7971,N_1369,N_1756);
and U7972 (N_7972,N_1422,N_2028);
and U7973 (N_7973,N_4880,N_1370);
nand U7974 (N_7974,N_5793,N_5560);
and U7975 (N_7975,N_5533,N_3844);
or U7976 (N_7976,N_2430,N_1310);
and U7977 (N_7977,N_5433,N_462);
nor U7978 (N_7978,N_1500,N_1162);
nand U7979 (N_7979,N_543,N_2549);
xor U7980 (N_7980,N_6235,N_1816);
or U7981 (N_7981,N_4771,N_934);
xnor U7982 (N_7982,N_6162,N_132);
or U7983 (N_7983,N_4513,N_277);
xor U7984 (N_7984,N_3211,N_3071);
nand U7985 (N_7985,N_3306,N_3566);
nand U7986 (N_7986,N_3513,N_4474);
and U7987 (N_7987,N_4742,N_2415);
or U7988 (N_7988,N_3148,N_335);
nand U7989 (N_7989,N_3917,N_5985);
xnor U7990 (N_7990,N_1775,N_5231);
and U7991 (N_7991,N_2956,N_2717);
nand U7992 (N_7992,N_1237,N_2346);
or U7993 (N_7993,N_4755,N_1533);
nor U7994 (N_7994,N_4914,N_2222);
and U7995 (N_7995,N_905,N_1663);
xnor U7996 (N_7996,N_2602,N_3415);
xor U7997 (N_7997,N_3438,N_5120);
or U7998 (N_7998,N_1190,N_749);
xor U7999 (N_7999,N_4387,N_4622);
nand U8000 (N_8000,N_3189,N_3357);
nor U8001 (N_8001,N_4875,N_6123);
nand U8002 (N_8002,N_4732,N_5251);
nor U8003 (N_8003,N_506,N_4857);
nand U8004 (N_8004,N_3954,N_1604);
and U8005 (N_8005,N_6,N_4118);
or U8006 (N_8006,N_3731,N_2583);
xnor U8007 (N_8007,N_6043,N_4683);
nor U8008 (N_8008,N_5166,N_3139);
nor U8009 (N_8009,N_4097,N_4109);
and U8010 (N_8010,N_4076,N_1525);
and U8011 (N_8011,N_3257,N_2101);
and U8012 (N_8012,N_3645,N_2667);
or U8013 (N_8013,N_4638,N_863);
xor U8014 (N_8014,N_4089,N_3777);
and U8015 (N_8015,N_5033,N_2332);
nor U8016 (N_8016,N_158,N_3450);
nor U8017 (N_8017,N_3609,N_5909);
xnor U8018 (N_8018,N_6163,N_3316);
nand U8019 (N_8019,N_1644,N_300);
nand U8020 (N_8020,N_2139,N_3052);
or U8021 (N_8021,N_5659,N_5622);
or U8022 (N_8022,N_4720,N_4438);
xor U8023 (N_8023,N_2544,N_768);
and U8024 (N_8024,N_4790,N_3013);
nor U8025 (N_8025,N_2695,N_1047);
xnor U8026 (N_8026,N_5468,N_4316);
or U8027 (N_8027,N_4933,N_5691);
nand U8028 (N_8028,N_2547,N_3882);
or U8029 (N_8029,N_363,N_2392);
nand U8030 (N_8030,N_1066,N_4700);
nor U8031 (N_8031,N_609,N_3680);
nand U8032 (N_8032,N_5072,N_399);
nand U8033 (N_8033,N_343,N_5879);
and U8034 (N_8034,N_3454,N_6106);
nor U8035 (N_8035,N_1143,N_5081);
or U8036 (N_8036,N_5424,N_4485);
or U8037 (N_8037,N_4094,N_1567);
and U8038 (N_8038,N_5447,N_4956);
or U8039 (N_8039,N_5225,N_5611);
xnor U8040 (N_8040,N_2592,N_2110);
nand U8041 (N_8041,N_2320,N_2754);
nand U8042 (N_8042,N_5034,N_651);
and U8043 (N_8043,N_2452,N_1953);
or U8044 (N_8044,N_5317,N_117);
or U8045 (N_8045,N_4948,N_6055);
and U8046 (N_8046,N_188,N_4307);
and U8047 (N_8047,N_2616,N_5668);
nand U8048 (N_8048,N_4166,N_4727);
or U8049 (N_8049,N_1635,N_5804);
nor U8050 (N_8050,N_5842,N_1060);
xnor U8051 (N_8051,N_5643,N_2439);
and U8052 (N_8052,N_2228,N_96);
xnor U8053 (N_8053,N_1438,N_4384);
nand U8054 (N_8054,N_4175,N_5934);
nand U8055 (N_8055,N_1749,N_1301);
or U8056 (N_8056,N_4954,N_3535);
or U8057 (N_8057,N_3060,N_3945);
nand U8058 (N_8058,N_3952,N_5037);
and U8059 (N_8059,N_1492,N_2270);
and U8060 (N_8060,N_2482,N_5133);
xor U8061 (N_8061,N_3184,N_5965);
and U8062 (N_8062,N_6117,N_830);
or U8063 (N_8063,N_5738,N_2730);
nor U8064 (N_8064,N_240,N_3990);
or U8065 (N_8065,N_3955,N_2059);
and U8066 (N_8066,N_4084,N_562);
nor U8067 (N_8067,N_1944,N_75);
nor U8068 (N_8068,N_4797,N_4992);
or U8069 (N_8069,N_6094,N_3947);
nor U8070 (N_8070,N_14,N_1811);
nor U8071 (N_8071,N_1721,N_193);
or U8072 (N_8072,N_1672,N_94);
nand U8073 (N_8073,N_2467,N_4123);
and U8074 (N_8074,N_4500,N_4047);
nand U8075 (N_8075,N_1124,N_2839);
xnor U8076 (N_8076,N_515,N_4717);
nor U8077 (N_8077,N_1801,N_4170);
xnor U8078 (N_8078,N_1214,N_4962);
nor U8079 (N_8079,N_1198,N_2387);
xor U8080 (N_8080,N_1113,N_3678);
or U8081 (N_8081,N_3665,N_1922);
xnor U8082 (N_8082,N_3883,N_697);
and U8083 (N_8083,N_2357,N_5258);
nor U8084 (N_8084,N_5818,N_5383);
nor U8085 (N_8085,N_3845,N_629);
nand U8086 (N_8086,N_137,N_5349);
and U8087 (N_8087,N_4666,N_1257);
or U8088 (N_8088,N_2384,N_3754);
and U8089 (N_8089,N_4752,N_4724);
xor U8090 (N_8090,N_1345,N_384);
nor U8091 (N_8091,N_2323,N_1958);
xor U8092 (N_8092,N_3332,N_1690);
nand U8093 (N_8093,N_2395,N_608);
and U8094 (N_8094,N_645,N_4824);
or U8095 (N_8095,N_3874,N_2968);
nand U8096 (N_8096,N_316,N_4333);
nand U8097 (N_8097,N_2316,N_770);
nor U8098 (N_8098,N_3048,N_5194);
xnor U8099 (N_8099,N_3288,N_4160);
nor U8100 (N_8100,N_898,N_6097);
nand U8101 (N_8101,N_1254,N_1629);
xnor U8102 (N_8102,N_3313,N_5604);
nor U8103 (N_8103,N_5868,N_5163);
xnor U8104 (N_8104,N_4062,N_3688);
nand U8105 (N_8105,N_735,N_4625);
nand U8106 (N_8106,N_63,N_3588);
or U8107 (N_8107,N_200,N_2295);
or U8108 (N_8108,N_3301,N_3961);
or U8109 (N_8109,N_2007,N_4003);
nand U8110 (N_8110,N_3497,N_5939);
and U8111 (N_8111,N_4028,N_2253);
or U8112 (N_8112,N_3358,N_6144);
and U8113 (N_8113,N_3836,N_1152);
xnor U8114 (N_8114,N_239,N_4318);
or U8115 (N_8115,N_3991,N_2604);
nor U8116 (N_8116,N_5469,N_2322);
nor U8117 (N_8117,N_5645,N_5650);
or U8118 (N_8118,N_3863,N_3590);
and U8119 (N_8119,N_3491,N_3652);
nand U8120 (N_8120,N_4884,N_5328);
nand U8121 (N_8121,N_5287,N_3940);
nand U8122 (N_8122,N_5093,N_805);
xor U8123 (N_8123,N_1514,N_4864);
xnor U8124 (N_8124,N_3043,N_414);
nor U8125 (N_8125,N_4078,N_4575);
and U8126 (N_8126,N_6101,N_167);
nand U8127 (N_8127,N_3387,N_5833);
nand U8128 (N_8128,N_3876,N_4002);
nor U8129 (N_8129,N_2641,N_1210);
or U8130 (N_8130,N_5352,N_4033);
and U8131 (N_8131,N_631,N_2618);
and U8132 (N_8132,N_5159,N_4737);
nand U8133 (N_8133,N_3814,N_998);
nand U8134 (N_8134,N_5751,N_3237);
nand U8135 (N_8135,N_2853,N_717);
nor U8136 (N_8136,N_893,N_4889);
nand U8137 (N_8137,N_5725,N_602);
nand U8138 (N_8138,N_103,N_5378);
nand U8139 (N_8139,N_3601,N_2173);
and U8140 (N_8140,N_3434,N_2603);
and U8141 (N_8141,N_2029,N_1711);
and U8142 (N_8142,N_5667,N_2820);
and U8143 (N_8143,N_5040,N_2141);
xor U8144 (N_8144,N_1813,N_1762);
xnor U8145 (N_8145,N_2743,N_2836);
and U8146 (N_8146,N_5692,N_4127);
nor U8147 (N_8147,N_3624,N_2240);
nor U8148 (N_8148,N_499,N_1169);
or U8149 (N_8149,N_3536,N_2537);
and U8150 (N_8150,N_5392,N_2391);
xnor U8151 (N_8151,N_4434,N_2777);
or U8152 (N_8152,N_2125,N_4593);
and U8153 (N_8153,N_5307,N_5008);
nand U8154 (N_8154,N_1648,N_3666);
or U8155 (N_8155,N_3877,N_3155);
nor U8156 (N_8156,N_4564,N_1181);
xor U8157 (N_8157,N_1194,N_5051);
xor U8158 (N_8158,N_1609,N_1580);
and U8159 (N_8159,N_5448,N_1768);
xor U8160 (N_8160,N_4041,N_4177);
nor U8161 (N_8161,N_4970,N_1387);
and U8162 (N_8162,N_3714,N_3293);
or U8163 (N_8163,N_2037,N_4901);
nand U8164 (N_8164,N_2247,N_1837);
xnor U8165 (N_8165,N_4779,N_43);
nand U8166 (N_8166,N_892,N_617);
nor U8167 (N_8167,N_4074,N_1156);
nand U8168 (N_8168,N_760,N_1287);
nand U8169 (N_8169,N_1681,N_1718);
xor U8170 (N_8170,N_5492,N_5432);
xor U8171 (N_8171,N_1303,N_5954);
and U8172 (N_8172,N_5374,N_6002);
xnor U8173 (N_8173,N_3395,N_97);
and U8174 (N_8174,N_6058,N_2140);
and U8175 (N_8175,N_3748,N_1932);
and U8176 (N_8176,N_1030,N_1319);
nor U8177 (N_8177,N_1823,N_4597);
or U8178 (N_8178,N_699,N_5049);
nor U8179 (N_8179,N_1914,N_1168);
nand U8180 (N_8180,N_1924,N_505);
or U8181 (N_8181,N_1776,N_2048);
nor U8182 (N_8182,N_4535,N_5815);
and U8183 (N_8183,N_3014,N_945);
or U8184 (N_8184,N_5061,N_2769);
or U8185 (N_8185,N_2861,N_152);
nor U8186 (N_8186,N_3200,N_2837);
nor U8187 (N_8187,N_5435,N_5398);
xor U8188 (N_8188,N_1243,N_2352);
nand U8189 (N_8189,N_4585,N_5181);
or U8190 (N_8190,N_2183,N_189);
xor U8191 (N_8191,N_5759,N_1328);
nor U8192 (N_8192,N_2359,N_292);
nand U8193 (N_8193,N_644,N_295);
xor U8194 (N_8194,N_3042,N_5261);
xor U8195 (N_8195,N_1280,N_5753);
and U8196 (N_8196,N_1766,N_5966);
nor U8197 (N_8197,N_1951,N_5846);
or U8198 (N_8198,N_2068,N_3801);
nor U8199 (N_8199,N_4905,N_2036);
or U8200 (N_8200,N_5333,N_3530);
xor U8201 (N_8201,N_572,N_234);
nand U8202 (N_8202,N_1817,N_4805);
xor U8203 (N_8203,N_1003,N_483);
xor U8204 (N_8204,N_1467,N_1488);
xor U8205 (N_8205,N_135,N_2302);
or U8206 (N_8206,N_1602,N_2179);
xor U8207 (N_8207,N_2711,N_1794);
nor U8208 (N_8208,N_5180,N_383);
nand U8209 (N_8209,N_5402,N_1427);
xnor U8210 (N_8210,N_825,N_5789);
or U8211 (N_8211,N_1702,N_3346);
xnor U8212 (N_8212,N_3312,N_2060);
or U8213 (N_8213,N_1322,N_5230);
nor U8214 (N_8214,N_1102,N_223);
or U8215 (N_8215,N_2453,N_5596);
nand U8216 (N_8216,N_678,N_4371);
nor U8217 (N_8217,N_968,N_5078);
and U8218 (N_8218,N_2305,N_6203);
nand U8219 (N_8219,N_2663,N_4716);
or U8220 (N_8220,N_4686,N_2167);
xor U8221 (N_8221,N_5672,N_1633);
and U8222 (N_8222,N_2202,N_3011);
or U8223 (N_8223,N_3729,N_1763);
or U8224 (N_8224,N_2466,N_4207);
or U8225 (N_8225,N_783,N_3764);
and U8226 (N_8226,N_4348,N_6136);
or U8227 (N_8227,N_3788,N_1767);
nor U8228 (N_8228,N_1186,N_525);
and U8229 (N_8229,N_4194,N_1283);
or U8230 (N_8230,N_5076,N_4959);
xnor U8231 (N_8231,N_5010,N_359);
xnor U8232 (N_8232,N_5271,N_4715);
xor U8233 (N_8233,N_4119,N_374);
and U8234 (N_8234,N_3284,N_1264);
and U8235 (N_8235,N_3393,N_5269);
and U8236 (N_8236,N_1729,N_4421);
and U8237 (N_8237,N_5716,N_2750);
or U8238 (N_8238,N_5085,N_2512);
and U8239 (N_8239,N_1576,N_4843);
or U8240 (N_8240,N_4661,N_2396);
nor U8241 (N_8241,N_1505,N_230);
xnor U8242 (N_8242,N_2226,N_2019);
nor U8243 (N_8243,N_3327,N_5760);
or U8244 (N_8244,N_1705,N_4818);
nor U8245 (N_8245,N_1118,N_2166);
or U8246 (N_8246,N_6147,N_6072);
and U8247 (N_8247,N_3143,N_1623);
or U8248 (N_8248,N_867,N_1487);
and U8249 (N_8249,N_4173,N_1035);
nand U8250 (N_8250,N_1265,N_4944);
nand U8251 (N_8251,N_3693,N_883);
nand U8252 (N_8252,N_285,N_947);
nor U8253 (N_8253,N_1581,N_2940);
or U8254 (N_8254,N_2808,N_425);
xor U8255 (N_8255,N_4215,N_1783);
nand U8256 (N_8256,N_2673,N_3547);
nor U8257 (N_8257,N_4351,N_4605);
and U8258 (N_8258,N_2459,N_5396);
nand U8259 (N_8259,N_1662,N_5722);
xor U8260 (N_8260,N_3692,N_2102);
or U8261 (N_8261,N_4449,N_2727);
nand U8262 (N_8262,N_902,N_3583);
or U8263 (N_8263,N_5229,N_4116);
nand U8264 (N_8264,N_5125,N_4367);
or U8265 (N_8265,N_3106,N_5938);
nor U8266 (N_8266,N_3025,N_2548);
or U8267 (N_8267,N_301,N_1074);
nand U8268 (N_8268,N_809,N_4083);
nand U8269 (N_8269,N_528,N_4926);
and U8270 (N_8270,N_1016,N_2303);
nor U8271 (N_8271,N_2712,N_5952);
nor U8272 (N_8272,N_4702,N_2938);
or U8273 (N_8273,N_5984,N_647);
nand U8274 (N_8274,N_1084,N_1327);
or U8275 (N_8275,N_5331,N_534);
nor U8276 (N_8276,N_442,N_454);
nand U8277 (N_8277,N_917,N_3036);
xnor U8278 (N_8278,N_2005,N_3366);
or U8279 (N_8279,N_3286,N_2710);
and U8280 (N_8280,N_620,N_2336);
and U8281 (N_8281,N_134,N_1947);
nand U8282 (N_8282,N_3270,N_1132);
and U8283 (N_8283,N_2988,N_1830);
xor U8284 (N_8284,N_1907,N_5869);
nand U8285 (N_8285,N_897,N_4903);
nand U8286 (N_8286,N_6035,N_3374);
xnor U8287 (N_8287,N_854,N_3985);
nand U8288 (N_8288,N_6182,N_4925);
or U8289 (N_8289,N_415,N_3232);
nor U8290 (N_8290,N_2032,N_3643);
nand U8291 (N_8291,N_1538,N_4515);
nor U8292 (N_8292,N_2798,N_398);
nand U8293 (N_8293,N_933,N_215);
and U8294 (N_8294,N_3292,N_761);
nand U8295 (N_8295,N_5540,N_1334);
nand U8296 (N_8296,N_5290,N_4913);
xnor U8297 (N_8297,N_3412,N_6045);
nand U8298 (N_8298,N_3934,N_5587);
nor U8299 (N_8299,N_2154,N_4248);
nor U8300 (N_8300,N_4789,N_169);
nor U8301 (N_8301,N_5953,N_1825);
or U8302 (N_8302,N_291,N_2844);
xor U8303 (N_8303,N_1382,N_2868);
and U8304 (N_8304,N_2699,N_1590);
and U8305 (N_8305,N_5283,N_3380);
and U8306 (N_8306,N_3923,N_3252);
or U8307 (N_8307,N_3337,N_2056);
xnor U8308 (N_8308,N_1927,N_1997);
or U8309 (N_8309,N_274,N_5291);
nor U8310 (N_8310,N_3614,N_6155);
xor U8311 (N_8311,N_2492,N_1923);
and U8312 (N_8312,N_2952,N_4695);
or U8313 (N_8313,N_2121,N_2405);
nand U8314 (N_8314,N_5372,N_3870);
nand U8315 (N_8315,N_4555,N_6232);
and U8316 (N_8316,N_4124,N_1131);
nor U8317 (N_8317,N_1835,N_5520);
nand U8318 (N_8318,N_1388,N_3488);
nand U8319 (N_8319,N_5670,N_880);
nand U8320 (N_8320,N_3223,N_1038);
and U8321 (N_8321,N_1227,N_1193);
or U8322 (N_8322,N_4218,N_6173);
or U8323 (N_8323,N_3304,N_5141);
nand U8324 (N_8324,N_5742,N_865);
and U8325 (N_8325,N_649,N_3168);
or U8326 (N_8326,N_1343,N_2827);
xnor U8327 (N_8327,N_3193,N_5971);
nor U8328 (N_8328,N_3636,N_325);
nor U8329 (N_8329,N_281,N_4289);
and U8330 (N_8330,N_1076,N_1620);
and U8331 (N_8331,N_275,N_518);
or U8332 (N_8332,N_3946,N_3922);
xnor U8333 (N_8333,N_4183,N_5138);
nor U8334 (N_8334,N_1161,N_2625);
nor U8335 (N_8335,N_3809,N_5535);
or U8336 (N_8336,N_5161,N_5987);
nor U8337 (N_8337,N_1857,N_1316);
and U8338 (N_8338,N_4418,N_5185);
xnor U8339 (N_8339,N_352,N_3679);
or U8340 (N_8340,N_4425,N_4895);
nor U8341 (N_8341,N_4489,N_3323);
or U8342 (N_8342,N_3861,N_3647);
nand U8343 (N_8343,N_5640,N_4579);
nor U8344 (N_8344,N_5488,N_3124);
or U8345 (N_8345,N_95,N_3145);
and U8346 (N_8346,N_1572,N_2265);
xor U8347 (N_8347,N_3469,N_2753);
nor U8348 (N_8348,N_197,N_6143);
nor U8349 (N_8349,N_2354,N_1368);
xor U8350 (N_8350,N_4787,N_2926);
nor U8351 (N_8351,N_5094,N_1271);
nor U8352 (N_8352,N_3974,N_652);
or U8353 (N_8353,N_3204,N_4498);
nor U8354 (N_8354,N_4488,N_4684);
nand U8355 (N_8355,N_5057,N_4394);
and U8356 (N_8356,N_2124,N_3558);
nand U8357 (N_8357,N_4182,N_3183);
nor U8358 (N_8358,N_4888,N_6047);
nor U8359 (N_8359,N_1208,N_3461);
nor U8360 (N_8360,N_1166,N_1350);
and U8361 (N_8361,N_1720,N_2951);
xor U8362 (N_8362,N_5199,N_874);
nor U8363 (N_8363,N_747,N_3546);
and U8364 (N_8364,N_4876,N_3255);
and U8365 (N_8365,N_5200,N_2417);
or U8366 (N_8366,N_3409,N_2864);
and U8367 (N_8367,N_3924,N_3027);
xnor U8368 (N_8368,N_3780,N_2648);
nor U8369 (N_8369,N_4354,N_1226);
and U8370 (N_8370,N_5609,N_5794);
nor U8371 (N_8371,N_4892,N_5784);
and U8372 (N_8372,N_4185,N_1632);
or U8373 (N_8373,N_2465,N_2628);
nand U8374 (N_8374,N_2086,N_1741);
and U8375 (N_8375,N_6241,N_5837);
nor U8376 (N_8376,N_688,N_1627);
nand U8377 (N_8377,N_4213,N_5092);
xnor U8378 (N_8378,N_466,N_1018);
xnor U8379 (N_8379,N_3160,N_4195);
or U8380 (N_8380,N_3804,N_4714);
xor U8381 (N_8381,N_769,N_207);
xnor U8382 (N_8382,N_3002,N_491);
nor U8383 (N_8383,N_2278,N_4237);
or U8384 (N_8384,N_746,N_2219);
xor U8385 (N_8385,N_5013,N_661);
and U8386 (N_8386,N_3586,N_743);
or U8387 (N_8387,N_3696,N_4694);
or U8388 (N_8388,N_864,N_1420);
xor U8389 (N_8389,N_2866,N_4982);
nand U8390 (N_8390,N_3740,N_757);
nor U8391 (N_8391,N_2218,N_2243);
nor U8392 (N_8392,N_186,N_4687);
or U8393 (N_8393,N_16,N_5162);
xnor U8394 (N_8394,N_4174,N_679);
nor U8395 (N_8395,N_5086,N_2015);
nor U8396 (N_8396,N_4531,N_1519);
nor U8397 (N_8397,N_3262,N_5176);
xor U8398 (N_8398,N_3224,N_2736);
or U8399 (N_8399,N_4130,N_5505);
and U8400 (N_8400,N_5245,N_5117);
xnor U8401 (N_8401,N_4095,N_5151);
nor U8402 (N_8402,N_4184,N_5456);
or U8403 (N_8403,N_35,N_3150);
xor U8404 (N_8404,N_4229,N_2264);
xor U8405 (N_8405,N_1979,N_2636);
and U8406 (N_8406,N_1436,N_5762);
nand U8407 (N_8407,N_1593,N_4061);
nand U8408 (N_8408,N_691,N_2841);
nand U8409 (N_8409,N_2431,N_1731);
xnor U8410 (N_8410,N_5305,N_3869);
and U8411 (N_8411,N_3871,N_2523);
or U8412 (N_8412,N_5016,N_6011);
and U8413 (N_8413,N_5772,N_2235);
and U8414 (N_8414,N_2476,N_2410);
nand U8415 (N_8415,N_4521,N_5877);
xnor U8416 (N_8416,N_3015,N_3584);
nand U8417 (N_8417,N_1855,N_278);
nand U8418 (N_8418,N_5787,N_4224);
nor U8419 (N_8419,N_5439,N_293);
nor U8420 (N_8420,N_1838,N_4359);
and U8421 (N_8421,N_6077,N_3265);
or U8422 (N_8422,N_479,N_3850);
nor U8423 (N_8423,N_3279,N_2344);
nor U8424 (N_8424,N_1984,N_4069);
xor U8425 (N_8425,N_5324,N_1233);
and U8426 (N_8426,N_6027,N_6120);
or U8427 (N_8427,N_2755,N_478);
and U8428 (N_8428,N_4427,N_3762);
nand U8429 (N_8429,N_312,N_1673);
or U8430 (N_8430,N_930,N_2939);
nor U8431 (N_8431,N_5248,N_4493);
and U8432 (N_8432,N_2886,N_5337);
and U8433 (N_8433,N_182,N_5038);
and U8434 (N_8434,N_81,N_67);
and U8435 (N_8435,N_5551,N_2229);
xnor U8436 (N_8436,N_4815,N_1961);
nor U8437 (N_8437,N_5648,N_3087);
and U8438 (N_8438,N_54,N_5736);
nor U8439 (N_8439,N_2716,N_522);
and U8440 (N_8440,N_4479,N_3550);
nand U8441 (N_8441,N_1616,N_5071);
nor U8442 (N_8442,N_5951,N_1231);
or U8443 (N_8443,N_4850,N_5617);
nand U8444 (N_8444,N_2205,N_2488);
nor U8445 (N_8445,N_3523,N_5493);
xor U8446 (N_8446,N_5394,N_996);
nand U8447 (N_8447,N_1158,N_3673);
nor U8448 (N_8448,N_2703,N_923);
or U8449 (N_8449,N_5872,N_5699);
nor U8450 (N_8450,N_6037,N_2541);
nor U8451 (N_8451,N_2137,N_3309);
or U8452 (N_8452,N_6088,N_5510);
and U8453 (N_8453,N_5655,N_1202);
nand U8454 (N_8454,N_4759,N_2058);
and U8455 (N_8455,N_2838,N_2963);
and U8456 (N_8456,N_98,N_1192);
and U8457 (N_8457,N_238,N_2872);
or U8458 (N_8458,N_1230,N_1774);
or U8459 (N_8459,N_6174,N_1485);
and U8460 (N_8460,N_512,N_4262);
or U8461 (N_8461,N_5860,N_3440);
nor U8462 (N_8462,N_973,N_1245);
nor U8463 (N_8463,N_4482,N_1414);
nor U8464 (N_8464,N_4595,N_1472);
or U8465 (N_8465,N_3460,N_6195);
nor U8466 (N_8466,N_1434,N_3243);
nand U8467 (N_8467,N_5958,N_6172);
xnor U8468 (N_8468,N_3282,N_4408);
nand U8469 (N_8469,N_576,N_6167);
xor U8470 (N_8470,N_306,N_5238);
nand U8471 (N_8471,N_102,N_5429);
nor U8472 (N_8472,N_4108,N_5319);
nor U8473 (N_8473,N_5898,N_4011);
nor U8474 (N_8474,N_2927,N_1406);
and U8475 (N_8475,N_1676,N_1530);
nor U8476 (N_8476,N_447,N_2168);
nand U8477 (N_8477,N_4582,N_5989);
nand U8478 (N_8478,N_37,N_4339);
nand U8479 (N_8479,N_3771,N_1282);
or U8480 (N_8480,N_4008,N_794);
xnor U8481 (N_8481,N_382,N_2609);
nor U8482 (N_8482,N_6129,N_5500);
xor U8483 (N_8483,N_3958,N_4163);
nand U8484 (N_8484,N_2795,N_1419);
nor U8485 (N_8485,N_3576,N_258);
or U8486 (N_8486,N_683,N_3188);
nor U8487 (N_8487,N_4406,N_4706);
and U8488 (N_8488,N_5462,N_5714);
nand U8489 (N_8489,N_667,N_5119);
and U8490 (N_8490,N_1591,N_3765);
or U8491 (N_8491,N_3842,N_2087);
and U8492 (N_8492,N_4680,N_390);
and U8493 (N_8493,N_5598,N_2654);
nor U8494 (N_8494,N_2209,N_982);
or U8495 (N_8495,N_1613,N_4904);
nand U8496 (N_8496,N_5198,N_5726);
nand U8497 (N_8497,N_2632,N_133);
xnor U8498 (N_8498,N_3386,N_5063);
or U8499 (N_8499,N_2977,N_1998);
xor U8500 (N_8500,N_5253,N_6073);
nor U8501 (N_8501,N_908,N_3716);
or U8502 (N_8502,N_4658,N_5529);
nand U8503 (N_8503,N_2650,N_2995);
nand U8504 (N_8504,N_3840,N_912);
nand U8505 (N_8505,N_5975,N_575);
nor U8506 (N_8506,N_1115,N_5318);
nor U8507 (N_8507,N_5096,N_5743);
nand U8508 (N_8508,N_5973,N_205);
or U8509 (N_8509,N_3141,N_3866);
or U8510 (N_8510,N_1435,N_4842);
nor U8511 (N_8511,N_2026,N_1481);
xnor U8512 (N_8512,N_4495,N_2813);
and U8513 (N_8513,N_6222,N_1363);
and U8514 (N_8514,N_3026,N_567);
or U8515 (N_8515,N_6145,N_5820);
nand U8516 (N_8516,N_1876,N_3382);
nand U8517 (N_8517,N_5687,N_3885);
nand U8518 (N_8518,N_5498,N_3977);
xor U8519 (N_8519,N_1708,N_707);
and U8520 (N_8520,N_4051,N_3915);
and U8521 (N_8521,N_4152,N_3004);
and U8522 (N_8522,N_3635,N_4059);
or U8523 (N_8523,N_5702,N_2751);
nand U8524 (N_8524,N_5077,N_5546);
nor U8525 (N_8525,N_5257,N_5202);
nand U8526 (N_8526,N_1355,N_2318);
nor U8527 (N_8527,N_1502,N_2634);
nand U8528 (N_8528,N_1157,N_74);
nand U8529 (N_8529,N_5004,N_1221);
or U8530 (N_8530,N_1560,N_2255);
and U8531 (N_8531,N_3608,N_3706);
nand U8532 (N_8532,N_3554,N_3720);
and U8533 (N_8533,N_2030,N_2136);
xor U8534 (N_8534,N_1153,N_3235);
and U8535 (N_8535,N_951,N_1988);
and U8536 (N_8536,N_1212,N_2909);
and U8537 (N_8537,N_6014,N_1261);
and U8538 (N_8538,N_2694,N_4896);
nor U8539 (N_8539,N_5219,N_962);
or U8540 (N_8540,N_31,N_4370);
nand U8541 (N_8541,N_2499,N_2047);
and U8542 (N_8542,N_5790,N_2373);
xnor U8543 (N_8543,N_5664,N_4512);
or U8544 (N_8544,N_2103,N_1797);
xnor U8545 (N_8545,N_2271,N_1315);
nor U8546 (N_8546,N_2171,N_4356);
and U8547 (N_8547,N_5735,N_38);
or U8548 (N_8548,N_455,N_26);
or U8549 (N_8549,N_925,N_3392);
xnor U8550 (N_8550,N_2317,N_2333);
xor U8551 (N_8551,N_2503,N_3967);
and U8552 (N_8552,N_2230,N_1841);
and U8553 (N_8553,N_148,N_5370);
nor U8554 (N_8554,N_3171,N_1417);
nor U8555 (N_8555,N_5927,N_4835);
nor U8556 (N_8556,N_2363,N_2135);
or U8557 (N_8557,N_4494,N_2525);
or U8558 (N_8558,N_5844,N_2903);
nand U8559 (N_8559,N_4407,N_5213);
and U8560 (N_8560,N_1934,N_816);
or U8561 (N_8561,N_1909,N_4052);
nor U8562 (N_8562,N_2283,N_4624);
or U8563 (N_8563,N_2573,N_1650);
xor U8564 (N_8564,N_5544,N_718);
or U8565 (N_8565,N_5835,N_2418);
nor U8566 (N_8566,N_4030,N_1486);
nand U8567 (N_8567,N_6010,N_5848);
xnor U8568 (N_8568,N_3962,N_5972);
nor U8569 (N_8569,N_2108,N_3352);
and U8570 (N_8570,N_3495,N_6041);
and U8571 (N_8571,N_5619,N_4459);
nand U8572 (N_8572,N_509,N_4690);
or U8573 (N_8573,N_2213,N_3290);
and U8574 (N_8574,N_5098,N_2591);
xnor U8575 (N_8575,N_2300,N_5808);
xor U8576 (N_8576,N_1091,N_2463);
nor U8577 (N_8577,N_201,N_606);
or U8578 (N_8578,N_2889,N_944);
nand U8579 (N_8579,N_671,N_1887);
nor U8580 (N_8580,N_5573,N_4337);
and U8581 (N_8581,N_6188,N_4921);
nand U8582 (N_8582,N_80,N_2582);
xnor U8583 (N_8583,N_1624,N_3020);
nor U8584 (N_8584,N_4627,N_3100);
and U8585 (N_8585,N_1510,N_1845);
or U8586 (N_8586,N_6039,N_4352);
nand U8587 (N_8587,N_985,N_9);
nor U8588 (N_8588,N_4096,N_1655);
nand U8589 (N_8589,N_2326,N_149);
xnor U8590 (N_8590,N_1272,N_1570);
xor U8591 (N_8591,N_4505,N_3837);
nand U8592 (N_8592,N_284,N_2388);
xor U8593 (N_8593,N_4171,N_5623);
or U8594 (N_8594,N_1079,N_3283);
nand U8595 (N_8595,N_4592,N_486);
nor U8596 (N_8596,N_3779,N_3649);
and U8597 (N_8597,N_5102,N_4272);
and U8598 (N_8598,N_1109,N_2257);
nor U8599 (N_8599,N_4335,N_1920);
or U8600 (N_8600,N_5680,N_3672);
nand U8601 (N_8601,N_4400,N_2468);
or U8602 (N_8602,N_597,N_1849);
xor U8603 (N_8603,N_2825,N_6001);
or U8604 (N_8604,N_3411,N_6092);
nor U8605 (N_8605,N_3035,N_2132);
or U8606 (N_8606,N_2885,N_4767);
or U8607 (N_8607,N_4234,N_823);
and U8608 (N_8608,N_1935,N_5007);
nor U8609 (N_8609,N_4353,N_2383);
nor U8610 (N_8610,N_4983,N_2937);
nor U8611 (N_8611,N_1005,N_3772);
xnor U8612 (N_8612,N_3973,N_5263);
or U8613 (N_8613,N_4424,N_3520);
and U8614 (N_8614,N_3308,N_4599);
nand U8615 (N_8615,N_1687,N_5366);
nor U8616 (N_8616,N_5580,N_5409);
or U8617 (N_8617,N_988,N_3221);
nor U8618 (N_8618,N_4381,N_705);
xor U8619 (N_8619,N_2521,N_3076);
or U8620 (N_8620,N_4239,N_5295);
nor U8621 (N_8621,N_1147,N_3539);
nor U8622 (N_8622,N_5478,N_4210);
and U8623 (N_8623,N_3406,N_4765);
or U8624 (N_8624,N_3300,N_3256);
and U8625 (N_8625,N_3887,N_2833);
or U8626 (N_8626,N_4922,N_4839);
nand U8627 (N_8627,N_2233,N_2922);
or U8628 (N_8628,N_1495,N_811);
nand U8629 (N_8629,N_675,N_3397);
nand U8630 (N_8630,N_3807,N_432);
nor U8631 (N_8631,N_2959,N_66);
nand U8632 (N_8632,N_2894,N_1089);
xnor U8633 (N_8633,N_1754,N_5782);
and U8634 (N_8634,N_2852,N_5362);
nor U8635 (N_8635,N_1000,N_2461);
nand U8636 (N_8636,N_5721,N_3658);
xnor U8637 (N_8637,N_921,N_1959);
or U8638 (N_8638,N_6067,N_993);
nand U8639 (N_8639,N_3157,N_2517);
nor U8640 (N_8640,N_138,N_1116);
and U8641 (N_8641,N_6218,N_3021);
xnor U8642 (N_8642,N_2594,N_165);
xor U8643 (N_8643,N_1299,N_2946);
and U8644 (N_8644,N_400,N_3641);
nand U8645 (N_8645,N_4520,N_2767);
xnor U8646 (N_8646,N_406,N_3444);
and U8647 (N_8647,N_5282,N_1724);
nand U8648 (N_8648,N_4232,N_3745);
nor U8649 (N_8649,N_368,N_1379);
nor U8650 (N_8650,N_5400,N_877);
xnor U8651 (N_8651,N_4772,N_520);
and U8652 (N_8652,N_5915,N_6249);
xor U8653 (N_8653,N_3486,N_5515);
xnor U8654 (N_8654,N_2947,N_890);
nand U8655 (N_8655,N_5090,N_2487);
xor U8656 (N_8656,N_5336,N_4448);
nand U8657 (N_8657,N_2870,N_4204);
nor U8658 (N_8658,N_1523,N_236);
xnor U8659 (N_8659,N_4065,N_1601);
or U8660 (N_8660,N_5964,N_5441);
or U8661 (N_8661,N_3089,N_1126);
nand U8662 (N_8662,N_3205,N_5286);
nand U8663 (N_8663,N_4122,N_4139);
and U8664 (N_8664,N_5884,N_5039);
nand U8665 (N_8665,N_2969,N_4623);
xor U8666 (N_8666,N_1022,N_355);
and U8667 (N_8667,N_2146,N_6247);
xor U8668 (N_8668,N_3617,N_5079);
nor U8669 (N_8669,N_5946,N_3050);
xnor U8670 (N_8670,N_3179,N_1104);
nor U8671 (N_8671,N_1824,N_4596);
nor U8672 (N_8672,N_4326,N_855);
xor U8673 (N_8673,N_3753,N_1963);
nand U8674 (N_8674,N_1742,N_1659);
xor U8675 (N_8675,N_3980,N_4244);
nand U8676 (N_8676,N_742,N_5218);
nor U8677 (N_8677,N_3059,N_5375);
nor U8678 (N_8678,N_5705,N_1750);
or U8679 (N_8679,N_5327,N_2123);
nor U8680 (N_8680,N_3811,N_1549);
or U8681 (N_8681,N_6180,N_1062);
or U8682 (N_8682,N_4031,N_4581);
nor U8683 (N_8683,N_719,N_3616);
nand U8684 (N_8684,N_5113,N_3373);
nor U8685 (N_8685,N_5996,N_4464);
nand U8686 (N_8686,N_3156,N_4271);
or U8687 (N_8687,N_1700,N_5831);
nand U8688 (N_8688,N_598,N_1869);
or U8689 (N_8689,N_5147,N_1359);
nor U8690 (N_8690,N_4251,N_4650);
or U8691 (N_8691,N_4025,N_5115);
and U8692 (N_8692,N_850,N_2372);
nor U8693 (N_8693,N_3884,N_1578);
nor U8694 (N_8694,N_1671,N_119);
or U8695 (N_8695,N_1286,N_4066);
and U8696 (N_8696,N_53,N_5564);
xor U8697 (N_8697,N_2221,N_5371);
xnor U8698 (N_8698,N_4741,N_859);
and U8699 (N_8699,N_1048,N_785);
nor U8700 (N_8700,N_1069,N_6083);
nand U8701 (N_8701,N_3396,N_4486);
and U8702 (N_8702,N_2685,N_2816);
or U8703 (N_8703,N_5461,N_5249);
or U8704 (N_8704,N_1815,N_6207);
and U8705 (N_8705,N_3864,N_815);
or U8706 (N_8706,N_5145,N_4557);
and U8707 (N_8707,N_3610,N_6244);
or U8708 (N_8708,N_5582,N_4679);
nand U8709 (N_8709,N_5157,N_115);
and U8710 (N_8710,N_1228,N_2989);
and U8711 (N_8711,N_1288,N_5830);
or U8712 (N_8712,N_1260,N_4522);
nor U8713 (N_8713,N_1589,N_4310);
or U8714 (N_8714,N_3621,N_639);
or U8715 (N_8715,N_446,N_1758);
and U8716 (N_8716,N_6229,N_5601);
nor U8717 (N_8717,N_1017,N_5531);
or U8718 (N_8718,N_4685,N_2996);
or U8719 (N_8719,N_1044,N_4473);
nor U8720 (N_8720,N_4443,N_2474);
or U8721 (N_8721,N_547,N_906);
nand U8722 (N_8722,N_2064,N_4253);
nand U8723 (N_8723,N_559,N_1691);
nand U8724 (N_8724,N_5438,N_1516);
nor U8725 (N_8725,N_4762,N_4783);
or U8726 (N_8726,N_1141,N_3023);
xor U8727 (N_8727,N_1870,N_4997);
or U8728 (N_8728,N_6023,N_2035);
or U8729 (N_8729,N_3466,N_1050);
or U8730 (N_8730,N_1911,N_3594);
xor U8731 (N_8731,N_4807,N_1861);
nor U8732 (N_8732,N_5017,N_131);
xnor U8733 (N_8733,N_759,N_2530);
nor U8734 (N_8734,N_3044,N_2414);
or U8735 (N_8735,N_725,N_5242);
xor U8736 (N_8736,N_122,N_4245);
xnor U8737 (N_8737,N_3655,N_5676);
nor U8738 (N_8738,N_6089,N_2651);
nor U8739 (N_8739,N_5404,N_3717);
nand U8740 (N_8740,N_2709,N_5497);
or U8741 (N_8741,N_1561,N_3318);
nor U8742 (N_8742,N_5050,N_5631);
nor U8743 (N_8743,N_3325,N_6166);
and U8744 (N_8744,N_3422,N_6205);
or U8745 (N_8745,N_3868,N_2763);
or U8746 (N_8746,N_586,N_1630);
nand U8747 (N_8747,N_3966,N_3988);
nor U8748 (N_8748,N_4611,N_4314);
xnor U8749 (N_8749,N_4725,N_3073);
nor U8750 (N_8750,N_4358,N_220);
or U8751 (N_8751,N_5889,N_2757);
nand U8752 (N_8752,N_2301,N_3414);
xor U8753 (N_8753,N_3456,N_2831);
or U8754 (N_8754,N_5866,N_3086);
and U8755 (N_8755,N_6237,N_6168);
nand U8756 (N_8756,N_4504,N_554);
and U8757 (N_8757,N_3920,N_3449);
or U8758 (N_8758,N_1266,N_178);
and U8759 (N_8759,N_5800,N_3003);
and U8760 (N_8760,N_729,N_4332);
nor U8761 (N_8761,N_1276,N_5660);
xnor U8762 (N_8762,N_2564,N_12);
or U8763 (N_8763,N_924,N_2964);
nor U8764 (N_8764,N_4786,N_5639);
nand U8765 (N_8765,N_4589,N_5697);
xor U8766 (N_8766,N_4726,N_594);
xnor U8767 (N_8767,N_2577,N_2073);
xor U8768 (N_8768,N_537,N_5393);
nor U8769 (N_8769,N_3858,N_1679);
nor U8770 (N_8770,N_3775,N_4454);
or U8771 (N_8771,N_2259,N_2307);
and U8772 (N_8772,N_5534,N_1873);
and U8773 (N_8773,N_1460,N_1441);
nor U8774 (N_8774,N_2043,N_4719);
nand U8775 (N_8775,N_2385,N_1378);
xnor U8776 (N_8776,N_680,N_5265);
and U8777 (N_8777,N_2070,N_3428);
and U8778 (N_8778,N_1972,N_1864);
nor U8779 (N_8779,N_3305,N_5930);
nand U8780 (N_8780,N_2846,N_3758);
xnor U8781 (N_8781,N_704,N_2244);
nand U8782 (N_8782,N_25,N_5195);
nor U8783 (N_8783,N_1020,N_833);
and U8784 (N_8784,N_5070,N_5164);
or U8785 (N_8785,N_1528,N_4987);
xor U8786 (N_8786,N_2574,N_4456);
xor U8787 (N_8787,N_4893,N_812);
and U8788 (N_8788,N_3976,N_4965);
and U8789 (N_8789,N_4143,N_4330);
nand U8790 (N_8790,N_5474,N_2768);
nor U8791 (N_8791,N_3631,N_723);
or U8792 (N_8792,N_3972,N_5390);
nor U8793 (N_8793,N_1028,N_1064);
or U8794 (N_8794,N_2120,N_784);
and U8795 (N_8795,N_1011,N_2929);
nor U8796 (N_8796,N_4057,N_3212);
nor U8797 (N_8797,N_1712,N_4542);
nand U8798 (N_8798,N_2345,N_2155);
and U8799 (N_8799,N_5537,N_1494);
or U8800 (N_8800,N_336,N_2904);
xnor U8801 (N_8801,N_1336,N_6009);
nand U8802 (N_8802,N_3573,N_3921);
nand U8803 (N_8803,N_6012,N_2623);
or U8804 (N_8804,N_2843,N_5184);
and U8805 (N_8805,N_2090,N_3348);
nand U8806 (N_8806,N_1293,N_659);
nor U8807 (N_8807,N_4544,N_1484);
nand U8808 (N_8808,N_2983,N_1138);
and U8809 (N_8809,N_4125,N_3186);
nand U8810 (N_8810,N_5060,N_1220);
and U8811 (N_8811,N_4015,N_2092);
xnor U8812 (N_8812,N_5308,N_3453);
xor U8813 (N_8813,N_573,N_1223);
or U8814 (N_8814,N_3363,N_5982);
nor U8815 (N_8815,N_4674,N_918);
xor U8816 (N_8816,N_3816,N_672);
or U8817 (N_8817,N_851,N_1274);
nand U8818 (N_8818,N_4428,N_2033);
and U8819 (N_8819,N_346,N_4707);
nand U8820 (N_8820,N_3975,N_4703);
and U8821 (N_8821,N_1646,N_6040);
nor U8822 (N_8822,N_1056,N_6153);
xor U8823 (N_8823,N_1443,N_1383);
xor U8824 (N_8824,N_4282,N_4104);
and U8825 (N_8825,N_1827,N_4209);
and U8826 (N_8826,N_402,N_2009);
and U8827 (N_8827,N_4411,N_5536);
nand U8828 (N_8828,N_5408,N_4006);
nand U8829 (N_8829,N_3220,N_4397);
and U8830 (N_8830,N_3208,N_953);
or U8831 (N_8831,N_4206,N_391);
xor U8832 (N_8832,N_428,N_5437);
nor U8833 (N_8833,N_2596,N_1562);
nor U8834 (N_8834,N_4098,N_2589);
xor U8835 (N_8835,N_6230,N_4247);
xnor U8836 (N_8836,N_4431,N_1755);
and U8837 (N_8837,N_2044,N_5994);
xnor U8838 (N_8838,N_1856,N_5148);
or U8839 (N_8839,N_1093,N_1105);
and U8840 (N_8840,N_4070,N_914);
or U8841 (N_8841,N_2266,N_361);
or U8842 (N_8842,N_1688,N_1985);
or U8843 (N_8843,N_4646,N_24);
nor U8844 (N_8844,N_4697,N_2027);
or U8845 (N_8845,N_3634,N_1582);
and U8846 (N_8846,N_4545,N_4383);
nand U8847 (N_8847,N_2854,N_1730);
and U8848 (N_8848,N_1215,N_900);
and U8849 (N_8849,N_2263,N_294);
nand U8850 (N_8850,N_5541,N_3786);
and U8851 (N_8851,N_1619,N_3310);
nor U8852 (N_8852,N_3551,N_5688);
nand U8853 (N_8853,N_4507,N_3886);
or U8854 (N_8854,N_2572,N_2933);
and U8855 (N_8855,N_3519,N_4632);
and U8856 (N_8856,N_1608,N_715);
and U8857 (N_8857,N_5344,N_4548);
and U8858 (N_8858,N_3012,N_5867);
nand U8859 (N_8859,N_776,N_1974);
xnor U8860 (N_8860,N_2152,N_4778);
or U8861 (N_8861,N_1357,N_3207);
and U8862 (N_8862,N_1246,N_1739);
nand U8863 (N_8863,N_4656,N_1146);
and U8864 (N_8864,N_3656,N_4541);
nand U8865 (N_8865,N_5259,N_1860);
nand U8866 (N_8866,N_3064,N_4995);
nand U8867 (N_8867,N_4202,N_1631);
nand U8868 (N_8868,N_1103,N_813);
and U8869 (N_8869,N_4659,N_1403);
nand U8870 (N_8870,N_4539,N_5775);
or U8871 (N_8871,N_1127,N_2481);
and U8872 (N_8872,N_684,N_490);
or U8873 (N_8873,N_3822,N_317);
nor U8874 (N_8874,N_1184,N_1087);
nand U8875 (N_8875,N_2527,N_303);
or U8876 (N_8876,N_788,N_225);
xnor U8877 (N_8877,N_60,N_6062);
and U8878 (N_8878,N_535,N_411);
nand U8879 (N_8879,N_2368,N_1901);
nand U8880 (N_8880,N_5919,N_1539);
and U8881 (N_8881,N_4971,N_2941);
or U8882 (N_8882,N_443,N_3817);
xor U8883 (N_8883,N_2100,N_2681);
and U8884 (N_8884,N_4528,N_2004);
nand U8885 (N_8885,N_3077,N_3854);
and U8886 (N_8886,N_6019,N_1344);
xnor U8887 (N_8887,N_4619,N_2312);
xnor U8888 (N_8888,N_1569,N_2279);
xnor U8889 (N_8889,N_2341,N_4178);
xor U8890 (N_8890,N_1902,N_6149);
nor U8891 (N_8891,N_626,N_2863);
nand U8892 (N_8892,N_4361,N_4825);
or U8893 (N_8893,N_3718,N_2528);
nor U8894 (N_8894,N_4841,N_5641);
nor U8895 (N_8895,N_221,N_5108);
or U8896 (N_8896,N_3937,N_4886);
nor U8897 (N_8897,N_250,N_1868);
and U8898 (N_8898,N_1496,N_371);
nor U8899 (N_8899,N_3949,N_1925);
nand U8900 (N_8900,N_1554,N_1027);
or U8901 (N_8901,N_5925,N_50);
nand U8902 (N_8902,N_4382,N_1149);
and U8903 (N_8903,N_4785,N_4255);
nand U8904 (N_8904,N_3006,N_4029);
nand U8905 (N_8905,N_46,N_3041);
and U8906 (N_8906,N_100,N_4629);
nand U8907 (N_8907,N_2731,N_2412);
xor U8908 (N_8908,N_664,N_1111);
nand U8909 (N_8909,N_5575,N_1164);
xor U8910 (N_8910,N_3993,N_803);
xnor U8911 (N_8911,N_4273,N_160);
or U8912 (N_8912,N_3075,N_1235);
nor U8913 (N_8913,N_5260,N_3135);
and U8914 (N_8914,N_4478,N_2752);
nor U8915 (N_8915,N_111,N_166);
xor U8916 (N_8916,N_2706,N_144);
xnor U8917 (N_8917,N_2486,N_1474);
xor U8918 (N_8918,N_5674,N_2371);
or U8919 (N_8919,N_5149,N_510);
and U8920 (N_8920,N_1086,N_2212);
nor U8921 (N_8921,N_2799,N_2696);
and U8922 (N_8922,N_3849,N_356);
or U8923 (N_8923,N_3339,N_1096);
or U8924 (N_8924,N_1915,N_1203);
xnor U8925 (N_8925,N_243,N_1761);
and U8926 (N_8926,N_3518,N_4458);
nand U8927 (N_8927,N_3689,N_2686);
nand U8928 (N_8928,N_6076,N_740);
nand U8929 (N_8929,N_5627,N_153);
and U8930 (N_8930,N_4217,N_4457);
or U8931 (N_8931,N_1574,N_3483);
xnor U8932 (N_8932,N_553,N_4035);
xnor U8933 (N_8933,N_5142,N_3146);
or U8934 (N_8934,N_1353,N_2586);
and U8935 (N_8935,N_5288,N_750);
nor U8936 (N_8936,N_5733,N_4385);
xor U8937 (N_8937,N_4492,N_5104);
xnor U8938 (N_8938,N_1361,N_3360);
nand U8939 (N_8939,N_4102,N_3736);
nor U8940 (N_8940,N_5182,N_4870);
nor U8941 (N_8941,N_5410,N_5446);
or U8942 (N_8942,N_872,N_3439);
and U8943 (N_8943,N_1063,N_3818);
or U8944 (N_8944,N_5330,N_4820);
xnor U8945 (N_8945,N_143,N_3033);
or U8946 (N_8946,N_4141,N_4526);
and U8947 (N_8947,N_2631,N_502);
xnor U8948 (N_8948,N_492,N_1053);
nand U8949 (N_8949,N_298,N_28);
nand U8950 (N_8950,N_4148,N_3032);
xnor U8951 (N_8951,N_5274,N_255);
nor U8952 (N_8952,N_4086,N_638);
nand U8953 (N_8953,N_1012,N_4009);
nand U8954 (N_8954,N_2117,N_3402);
or U8955 (N_8955,N_4236,N_3101);
nand U8956 (N_8956,N_1542,N_3796);
nand U8957 (N_8957,N_372,N_5443);
nand U8958 (N_8958,N_3216,N_6126);
xnor U8959 (N_8959,N_1456,N_4093);
nor U8960 (N_8960,N_5309,N_3531);
nand U8961 (N_8961,N_2942,N_3750);
or U8962 (N_8962,N_682,N_5323);
nand U8963 (N_8963,N_2350,N_4496);
nor U8964 (N_8964,N_5801,N_2822);
or U8965 (N_8965,N_6191,N_926);
and U8966 (N_8966,N_4709,N_882);
xor U8967 (N_8967,N_2329,N_2325);
xor U8968 (N_8968,N_2791,N_4899);
xor U8969 (N_8969,N_2214,N_3529);
nor U8970 (N_8970,N_3919,N_4293);
and U8971 (N_8971,N_5579,N_173);
nand U8972 (N_8972,N_2565,N_3037);
nand U8973 (N_8973,N_1628,N_6194);
and U8974 (N_8974,N_1393,N_6114);
and U8975 (N_8975,N_334,N_5137);
and U8976 (N_8976,N_5980,N_468);
xnor U8977 (N_8977,N_3199,N_5662);
or U8978 (N_8978,N_5937,N_4506);
and U8979 (N_8979,N_5356,N_2800);
nor U8980 (N_8980,N_1218,N_6021);
xor U8981 (N_8981,N_3970,N_4814);
or U8982 (N_8982,N_4285,N_511);
or U8983 (N_8983,N_5284,N_1759);
xnor U8984 (N_8984,N_4034,N_1980);
xnor U8985 (N_8985,N_1333,N_4350);
or U8986 (N_8986,N_4233,N_4201);
nand U8987 (N_8987,N_5887,N_99);
nor U8988 (N_8988,N_2526,N_2403);
or U8989 (N_8989,N_6025,N_5158);
or U8990 (N_8990,N_4951,N_5457);
or U8991 (N_8991,N_3218,N_4509);
nand U8992 (N_8992,N_2734,N_1640);
or U8993 (N_8993,N_5475,N_2420);
nor U8994 (N_8994,N_870,N_2501);
or U8995 (N_8995,N_4766,N_1531);
and U8996 (N_8996,N_2945,N_3452);
and U8997 (N_8997,N_2917,N_5338);
nand U8998 (N_8998,N_3082,N_4007);
or U8999 (N_8999,N_3657,N_4898);
xnor U9000 (N_9000,N_5114,N_5684);
and U9001 (N_9001,N_4648,N_326);
xor U9002 (N_9002,N_3410,N_5847);
or U9003 (N_9003,N_994,N_5734);
nand U9004 (N_9004,N_5190,N_3715);
nand U9005 (N_9005,N_3964,N_2046);
nand U9006 (N_9006,N_4630,N_2830);
nor U9007 (N_9007,N_5933,N_1384);
xor U9008 (N_9008,N_4792,N_3062);
nand U9009 (N_9009,N_3047,N_689);
and U9010 (N_9010,N_701,N_4877);
nor U9011 (N_9011,N_5859,N_1397);
nor U9012 (N_9012,N_1170,N_1236);
nand U9013 (N_9013,N_1464,N_952);
xor U9014 (N_9014,N_2254,N_3030);
xor U9015 (N_9015,N_1418,N_3250);
nor U9016 (N_9016,N_5422,N_899);
and U9017 (N_9017,N_2851,N_5047);
or U9018 (N_9018,N_6029,N_5986);
nor U9019 (N_9019,N_3739,N_5121);
or U9020 (N_9020,N_2310,N_3367);
nor U9021 (N_9021,N_3274,N_4793);
and U9022 (N_9022,N_4934,N_420);
xnor U9023 (N_9023,N_4140,N_5796);
and U9024 (N_9024,N_2297,N_3239);
nand U9025 (N_9025,N_409,N_3639);
nor U9026 (N_9026,N_5022,N_4142);
and U9027 (N_9027,N_904,N_4048);
nand U9028 (N_9028,N_5255,N_4881);
nor U9029 (N_9029,N_4830,N_588);
nand U9030 (N_9030,N_3951,N_2321);
nor U9031 (N_9031,N_4395,N_2559);
xnor U9032 (N_9032,N_1520,N_1605);
nor U9033 (N_9033,N_2182,N_5321);
nor U9034 (N_9034,N_878,N_59);
and U9035 (N_9035,N_5103,N_764);
xnor U9036 (N_9036,N_1155,N_5785);
nand U9037 (N_9037,N_1957,N_297);
or U9038 (N_9038,N_4985,N_4651);
nor U9039 (N_9039,N_4976,N_931);
or U9040 (N_9040,N_4806,N_4145);
and U9041 (N_9041,N_5524,N_5910);
or U9042 (N_9042,N_5883,N_5834);
and U9043 (N_9043,N_1971,N_5666);
and U9044 (N_9044,N_820,N_2072);
or U9045 (N_9045,N_3158,N_4067);
and U9046 (N_9046,N_1728,N_3298);
xnor U9047 (N_9047,N_3582,N_6024);
nor U9048 (N_9048,N_4013,N_835);
nand U9049 (N_9049,N_2001,N_3741);
nand U9050 (N_9050,N_4968,N_1831);
and U9051 (N_9051,N_2309,N_1483);
and U9052 (N_9052,N_5171,N_3049);
nand U9053 (N_9053,N_5471,N_307);
nor U9054 (N_9054,N_5629,N_3602);
nor U9055 (N_9055,N_2076,N_3603);
or U9056 (N_9056,N_4819,N_2376);
and U9057 (N_9057,N_6082,N_1675);
nor U9058 (N_9058,N_4989,N_712);
and U9059 (N_9059,N_3191,N_5075);
nor U9060 (N_9060,N_919,N_141);
nand U9061 (N_9061,N_4475,N_5420);
or U9062 (N_9062,N_1832,N_5067);
and U9063 (N_9063,N_5292,N_1351);
nand U9064 (N_9064,N_2958,N_302);
nor U9065 (N_9065,N_3302,N_5849);
nand U9066 (N_9066,N_1239,N_257);
nor U9067 (N_9067,N_2600,N_4404);
xnor U9068 (N_9068,N_493,N_4909);
and U9069 (N_9069,N_5209,N_2906);
nor U9070 (N_9070,N_5046,N_6161);
or U9071 (N_9071,N_5517,N_2571);
nand U9072 (N_9072,N_3117,N_2997);
nor U9073 (N_9073,N_68,N_2435);
and U9074 (N_9074,N_4099,N_3123);
nor U9075 (N_9075,N_354,N_123);
and U9076 (N_9076,N_4036,N_4126);
nand U9077 (N_9077,N_157,N_6070);
nand U9078 (N_9078,N_1042,N_2888);
and U9079 (N_9079,N_5701,N_978);
or U9080 (N_9080,N_2542,N_2775);
xor U9081 (N_9081,N_5821,N_1636);
and U9082 (N_9082,N_5032,N_1244);
or U9083 (N_9083,N_4978,N_4497);
xnor U9084 (N_9084,N_1643,N_2250);
or U9085 (N_9085,N_848,N_5501);
xnor U9086 (N_9086,N_5234,N_5518);
nand U9087 (N_9087,N_4761,N_2642);
nand U9088 (N_9088,N_1278,N_2826);
or U9089 (N_9089,N_2691,N_4847);
xnor U9090 (N_9090,N_4403,N_3695);
nor U9091 (N_9091,N_1559,N_5584);
nor U9092 (N_9092,N_4996,N_5992);
or U9093 (N_9093,N_175,N_4900);
nor U9094 (N_9094,N_3010,N_858);
or U9095 (N_9095,N_2241,N_5298);
xnor U9096 (N_9096,N_1009,N_3795);
or U9097 (N_9097,N_4106,N_1051);
and U9098 (N_9098,N_1625,N_184);
and U9099 (N_9099,N_4682,N_5571);
xor U9100 (N_9100,N_2042,N_1696);
xnor U9101 (N_9101,N_6069,N_3464);
or U9102 (N_9102,N_3091,N_385);
xnor U9103 (N_9103,N_5264,N_5636);
nor U9104 (N_9104,N_261,N_6139);
or U9105 (N_9105,N_5024,N_1937);
or U9106 (N_9106,N_6112,N_5873);
nand U9107 (N_9107,N_3944,N_2083);
and U9108 (N_9108,N_6093,N_2193);
xnor U9109 (N_9109,N_5706,N_2018);
or U9110 (N_9110,N_1471,N_2024);
nor U9111 (N_9111,N_2306,N_5440);
and U9112 (N_9112,N_2704,N_3773);
or U9113 (N_9113,N_5484,N_3555);
nor U9114 (N_9114,N_3891,N_1586);
nor U9115 (N_9115,N_5961,N_5956);
nor U9116 (N_9116,N_4981,N_587);
nand U9117 (N_9117,N_4538,N_2976);
nand U9118 (N_9118,N_5554,N_4657);
or U9119 (N_9119,N_837,N_1222);
xor U9120 (N_9120,N_1392,N_5364);
nand U9121 (N_9121,N_245,N_2509);
nand U9122 (N_9122,N_1618,N_4817);
xor U9123 (N_9123,N_4967,N_181);
nor U9124 (N_9124,N_5350,N_4963);
xor U9125 (N_9125,N_73,N_596);
or U9126 (N_9126,N_2159,N_1928);
nand U9127 (N_9127,N_887,N_3259);
nor U9128 (N_9128,N_5817,N_5414);
xnor U9129 (N_9129,N_1926,N_5365);
or U9130 (N_9130,N_4751,N_3333);
nor U9131 (N_9131,N_1991,N_940);
xor U9132 (N_9132,N_2394,N_4132);
xnor U9133 (N_9133,N_808,N_5899);
xnor U9134 (N_9134,N_5950,N_2771);
or U9135 (N_9135,N_5247,N_1167);
nand U9136 (N_9136,N_4260,N_2646);
xnor U9137 (N_9137,N_1975,N_365);
xnor U9138 (N_9138,N_5630,N_3121);
nand U9139 (N_9139,N_1701,N_5797);
xnor U9140 (N_9140,N_1900,N_6185);
nor U9141 (N_9141,N_351,N_5538);
nor U9142 (N_9142,N_6233,N_839);
nor U9143 (N_9143,N_367,N_2052);
nand U9144 (N_9144,N_329,N_164);
xnor U9145 (N_9145,N_4056,N_2149);
xor U9146 (N_9146,N_1880,N_3596);
or U9147 (N_9147,N_992,N_3521);
nand U9148 (N_9148,N_3611,N_4836);
nor U9149 (N_9149,N_375,N_2925);
nand U9150 (N_9150,N_706,N_3544);
nand U9151 (N_9151,N_6008,N_3761);
nor U9152 (N_9152,N_4072,N_5717);
nor U9153 (N_9153,N_3803,N_89);
xor U9154 (N_9154,N_948,N_1875);
or U9155 (N_9155,N_4587,N_222);
nand U9156 (N_9156,N_790,N_2224);
and U9157 (N_9157,N_5083,N_1253);
and U9158 (N_9158,N_118,N_5578);
nor U9159 (N_9159,N_1771,N_3303);
or U9160 (N_9160,N_3326,N_3144);
nor U9161 (N_9161,N_2656,N_4776);
nor U9162 (N_9162,N_2921,N_1277);
and U9163 (N_9163,N_3493,N_3066);
or U9164 (N_9164,N_3709,N_766);
and U9165 (N_9165,N_4670,N_1291);
or U9166 (N_9166,N_4016,N_3747);
nand U9167 (N_9167,N_1425,N_1843);
nor U9168 (N_9168,N_4733,N_838);
and U9169 (N_9169,N_2606,N_1791);
xnor U9170 (N_9170,N_5256,N_508);
and U9171 (N_9171,N_1007,N_72);
nand U9172 (N_9172,N_970,N_533);
or U9173 (N_9173,N_4671,N_4919);
or U9174 (N_9174,N_3542,N_5006);
nor U9175 (N_9175,N_1723,N_4386);
nand U9176 (N_9176,N_5451,N_4219);
xnor U9177 (N_9177,N_2802,N_3648);
xnor U9178 (N_9178,N_1150,N_4546);
xnor U9179 (N_9179,N_1706,N_3040);
nand U9180 (N_9180,N_989,N_4270);
xnor U9181 (N_9181,N_3815,N_5857);
or U9182 (N_9182,N_4559,N_3379);
or U9183 (N_9183,N_3553,N_949);
nor U9184 (N_9184,N_1412,N_681);
nor U9185 (N_9185,N_3451,N_1664);
and U9186 (N_9186,N_4524,N_5473);
and U9187 (N_9187,N_5661,N_5729);
or U9188 (N_9188,N_5191,N_1371);
xnor U9189 (N_9189,N_2081,N_903);
and U9190 (N_9190,N_2511,N_6121);
xnor U9191 (N_9191,N_5346,N_1509);
xnor U9192 (N_9192,N_3319,N_832);
or U9193 (N_9193,N_3812,N_541);
nor U9194 (N_9194,N_4604,N_5988);
or U9195 (N_9195,N_5369,N_958);
nor U9196 (N_9196,N_6119,N_3819);
or U9197 (N_9197,N_252,N_2856);
or U9198 (N_9198,N_2665,N_2495);
and U9199 (N_9199,N_564,N_299);
and U9200 (N_9200,N_6042,N_4181);
xnor U9201 (N_9201,N_1686,N_1292);
xnor U9202 (N_9202,N_1557,N_2460);
and U9203 (N_9203,N_1976,N_4312);
nand U9204 (N_9204,N_1329,N_4450);
and U9205 (N_9205,N_3260,N_4355);
xor U9206 (N_9206,N_5998,N_3723);
xor U9207 (N_9207,N_5188,N_3528);
xor U9208 (N_9208,N_1100,N_3927);
and U9209 (N_9209,N_579,N_3355);
nor U9210 (N_9210,N_388,N_0);
and U9211 (N_9211,N_4187,N_4045);
nand U9212 (N_9212,N_5839,N_1177);
nand U9213 (N_9213,N_2581,N_4050);
xnor U9214 (N_9214,N_3351,N_5416);
or U9215 (N_9215,N_1946,N_6220);
nand U9216 (N_9216,N_592,N_3781);
or U9217 (N_9217,N_709,N_1325);
and U9218 (N_9218,N_3019,N_3625);
xnor U9219 (N_9219,N_2629,N_1722);
or U9220 (N_9220,N_3194,N_4891);
nor U9221 (N_9221,N_5355,N_965);
and U9222 (N_9222,N_2122,N_273);
or U9223 (N_9223,N_5881,N_4252);
nor U9224 (N_9224,N_545,N_5566);
or U9225 (N_9225,N_3126,N_1552);
nand U9226 (N_9226,N_3722,N_3094);
nand U9227 (N_9227,N_5491,N_2747);
nor U9228 (N_9228,N_3730,N_5172);
nand U9229 (N_9229,N_4205,N_5278);
nand U9230 (N_9230,N_4728,N_5386);
xor U9231 (N_9231,N_1059,N_3664);
xnor U9232 (N_9232,N_2187,N_964);
nor U9233 (N_9233,N_685,N_2067);
nor U9234 (N_9234,N_6238,N_1973);
or U9235 (N_9235,N_1929,N_2949);
or U9236 (N_9236,N_484,N_4863);
or U9237 (N_9237,N_3432,N_4412);
nand U9238 (N_9238,N_4809,N_3273);
and U9239 (N_9239,N_1058,N_3261);
xnor U9240 (N_9240,N_5411,N_571);
and U9241 (N_9241,N_5495,N_4200);
and U9242 (N_9242,N_3371,N_4191);
and U9243 (N_9243,N_2781,N_180);
xor U9244 (N_9244,N_3078,N_716);
and U9245 (N_9245,N_3127,N_29);
or U9246 (N_9246,N_2533,N_548);
nor U9247 (N_9247,N_393,N_5807);
and U9248 (N_9248,N_3134,N_449);
or U9249 (N_9249,N_1493,N_955);
nand U9250 (N_9250,N_2185,N_5340);
nand U9251 (N_9251,N_1323,N_1882);
xor U9252 (N_9252,N_2133,N_1969);
xor U9253 (N_9253,N_146,N_4044);
xor U9254 (N_9254,N_655,N_1930);
nand U9255 (N_9255,N_5748,N_2365);
or U9256 (N_9256,N_4469,N_495);
nand U9257 (N_9257,N_3448,N_3509);
nand U9258 (N_9258,N_1703,N_4432);
and U9259 (N_9259,N_5791,N_4770);
nor U9260 (N_9260,N_4288,N_4998);
or U9261 (N_9261,N_1802,N_2993);
nand U9262 (N_9262,N_1444,N_4144);
nand U9263 (N_9263,N_2913,N_4315);
xor U9264 (N_9264,N_4653,N_4068);
or U9265 (N_9265,N_4567,N_5893);
nor U9266 (N_9266,N_563,N_3846);
or U9267 (N_9267,N_1697,N_4319);
nor U9268 (N_9268,N_395,N_2655);
or U9269 (N_9269,N_5969,N_972);
nor U9270 (N_9270,N_108,N_1199);
or U9271 (N_9271,N_5926,N_2497);
and U9272 (N_9272,N_5805,N_470);
or U9273 (N_9273,N_3107,N_3838);
nand U9274 (N_9274,N_3901,N_3187);
nand U9275 (N_9275,N_5905,N_2404);
nor U9276 (N_9276,N_4588,N_1335);
xor U9277 (N_9277,N_733,N_4573);
or U9278 (N_9278,N_86,N_1904);
xnor U9279 (N_9279,N_4617,N_3577);
or U9280 (N_9280,N_6240,N_2456);
nand U9281 (N_9281,N_4435,N_2538);
nor U9282 (N_9282,N_4768,N_5379);
nand U9283 (N_9283,N_1395,N_5407);
and U9284 (N_9284,N_5123,N_366);
xor U9285 (N_9285,N_963,N_5106);
or U9286 (N_9286,N_4991,N_2079);
and U9287 (N_9287,N_2848,N_5233);
xnor U9288 (N_9288,N_1341,N_1401);
nand U9289 (N_9289,N_4372,N_5902);
or U9290 (N_9290,N_4396,N_3177);
xnor U9291 (N_9291,N_2143,N_3640);
or U9292 (N_9292,N_4296,N_4398);
and U9293 (N_9293,N_2612,N_4240);
or U9294 (N_9294,N_4416,N_3810);
xor U9295 (N_9295,N_1374,N_3028);
xnor U9296 (N_9296,N_2490,N_4151);
nor U9297 (N_9297,N_2828,N_4230);
nor U9298 (N_9298,N_2398,N_226);
xnor U9299 (N_9299,N_4313,N_1587);
nand U9300 (N_9300,N_1599,N_1078);
nor U9301 (N_9301,N_4060,N_1386);
nor U9302 (N_9302,N_4788,N_1160);
xnor U9303 (N_9303,N_3163,N_4799);
and U9304 (N_9304,N_741,N_2386);
nor U9305 (N_9305,N_5459,N_1356);
xnor U9306 (N_9306,N_4749,N_3630);
and U9307 (N_9307,N_1987,N_5920);
or U9308 (N_9308,N_2671,N_4441);
and U9309 (N_9309,N_5747,N_4620);
or U9310 (N_9310,N_4075,N_4882);
and U9311 (N_9311,N_272,N_13);
xnor U9312 (N_9312,N_720,N_745);
xor U9313 (N_9313,N_2175,N_3792);
or U9314 (N_9314,N_611,N_5755);
xnor U9315 (N_9315,N_6157,N_2697);
and U9316 (N_9316,N_1844,N_910);
and U9317 (N_9317,N_2189,N_2409);
and U9318 (N_9318,N_777,N_1592);
or U9319 (N_9319,N_1541,N_4961);
or U9320 (N_9320,N_421,N_2893);
and U9321 (N_9321,N_1566,N_3359);
and U9322 (N_9322,N_5031,N_4699);
nand U9323 (N_9323,N_5678,N_3627);
nand U9324 (N_9324,N_22,N_569);
nor U9325 (N_9325,N_1527,N_5201);
nand U9326 (N_9326,N_4848,N_5132);
nor U9327 (N_9327,N_2790,N_2472);
nand U9328 (N_9328,N_2464,N_2016);
or U9329 (N_9329,N_2626,N_2728);
nor U9330 (N_9330,N_819,N_6109);
nor U9331 (N_9331,N_5417,N_3474);
nand U9332 (N_9332,N_4743,N_5425);
xor U9333 (N_9333,N_2638,N_4364);
or U9334 (N_9334,N_5152,N_5289);
nor U9335 (N_9335,N_5530,N_3790);
xor U9336 (N_9336,N_1654,N_1128);
and U9337 (N_9337,N_5911,N_5663);
xnor U9338 (N_9338,N_3480,N_3830);
nand U9339 (N_9339,N_3978,N_1130);
nand U9340 (N_9340,N_2611,N_762);
nor U9341 (N_9341,N_4645,N_5878);
or U9342 (N_9342,N_4105,N_3433);
nor U9343 (N_9343,N_6113,N_2248);
nor U9344 (N_9344,N_4942,N_3162);
xnor U9345 (N_9345,N_5809,N_4947);
nor U9346 (N_9346,N_1183,N_1993);
and U9347 (N_9347,N_2677,N_2678);
and U9348 (N_9348,N_2506,N_2554);
and U9349 (N_9349,N_5570,N_1765);
nor U9350 (N_9350,N_5273,N_1121);
nor U9351 (N_9351,N_2599,N_5783);
nor U9352 (N_9352,N_1320,N_471);
or U9353 (N_9353,N_1025,N_4812);
nand U9354 (N_9354,N_3743,N_5752);
and U9355 (N_9355,N_2369,N_4071);
nor U9356 (N_9356,N_1267,N_2794);
and U9357 (N_9357,N_4346,N_2518);
xnor U9358 (N_9358,N_5434,N_4549);
nor U9359 (N_9359,N_3268,N_1373);
or U9360 (N_9360,N_3254,N_3968);
xnor U9361 (N_9361,N_666,N_5977);
xnor U9362 (N_9362,N_6105,N_3383);
nor U9363 (N_9363,N_3872,N_2758);
or U9364 (N_9364,N_5577,N_3618);
or U9365 (N_9365,N_4613,N_5968);
nor U9366 (N_9366,N_4584,N_5268);
xor U9367 (N_9367,N_5228,N_2145);
nand U9368 (N_9368,N_570,N_4654);
or U9369 (N_9369,N_857,N_5100);
nor U9370 (N_9370,N_3929,N_282);
and U9371 (N_9371,N_5646,N_2551);
and U9372 (N_9372,N_5923,N_3197);
xnor U9373 (N_9373,N_2201,N_5127);
and U9374 (N_9374,N_1263,N_2429);
nand U9375 (N_9375,N_4812,N_3192);
and U9376 (N_9376,N_1480,N_4657);
xor U9377 (N_9377,N_2020,N_1131);
nand U9378 (N_9378,N_5573,N_1041);
or U9379 (N_9379,N_5641,N_186);
xnor U9380 (N_9380,N_1189,N_2718);
xnor U9381 (N_9381,N_2444,N_1487);
xor U9382 (N_9382,N_5558,N_848);
and U9383 (N_9383,N_389,N_810);
or U9384 (N_9384,N_2778,N_3128);
xor U9385 (N_9385,N_3446,N_773);
nand U9386 (N_9386,N_5559,N_5291);
nor U9387 (N_9387,N_3899,N_1303);
nor U9388 (N_9388,N_1301,N_1630);
nand U9389 (N_9389,N_1114,N_4496);
nor U9390 (N_9390,N_3194,N_3101);
nor U9391 (N_9391,N_2805,N_4783);
nand U9392 (N_9392,N_1863,N_4578);
or U9393 (N_9393,N_296,N_655);
nand U9394 (N_9394,N_13,N_1354);
and U9395 (N_9395,N_3754,N_4974);
xnor U9396 (N_9396,N_109,N_4071);
nand U9397 (N_9397,N_5548,N_6154);
nor U9398 (N_9398,N_3291,N_1859);
xnor U9399 (N_9399,N_945,N_131);
xor U9400 (N_9400,N_3398,N_4727);
or U9401 (N_9401,N_5250,N_135);
and U9402 (N_9402,N_4623,N_2502);
nor U9403 (N_9403,N_1461,N_6208);
xor U9404 (N_9404,N_3722,N_4093);
nor U9405 (N_9405,N_1907,N_2727);
and U9406 (N_9406,N_5472,N_3791);
or U9407 (N_9407,N_1120,N_2522);
or U9408 (N_9408,N_76,N_3799);
or U9409 (N_9409,N_2836,N_745);
or U9410 (N_9410,N_5912,N_5807);
xnor U9411 (N_9411,N_92,N_2360);
and U9412 (N_9412,N_607,N_1630);
nand U9413 (N_9413,N_6215,N_2451);
xor U9414 (N_9414,N_5525,N_262);
or U9415 (N_9415,N_1661,N_6023);
nor U9416 (N_9416,N_842,N_5988);
or U9417 (N_9417,N_5199,N_1923);
nor U9418 (N_9418,N_2086,N_2770);
nor U9419 (N_9419,N_6192,N_3511);
and U9420 (N_9420,N_1048,N_583);
and U9421 (N_9421,N_963,N_5794);
and U9422 (N_9422,N_5420,N_6082);
or U9423 (N_9423,N_3002,N_2554);
and U9424 (N_9424,N_5023,N_2246);
nand U9425 (N_9425,N_1192,N_4230);
nor U9426 (N_9426,N_929,N_1376);
xor U9427 (N_9427,N_4680,N_1241);
nor U9428 (N_9428,N_5460,N_1786);
or U9429 (N_9429,N_3935,N_589);
nand U9430 (N_9430,N_1007,N_1594);
nor U9431 (N_9431,N_2046,N_124);
nand U9432 (N_9432,N_4381,N_5270);
nor U9433 (N_9433,N_1138,N_1767);
nor U9434 (N_9434,N_1117,N_2966);
nand U9435 (N_9435,N_4576,N_2846);
nand U9436 (N_9436,N_1455,N_874);
nor U9437 (N_9437,N_5217,N_4325);
nand U9438 (N_9438,N_3734,N_5904);
or U9439 (N_9439,N_512,N_3420);
nand U9440 (N_9440,N_1271,N_2539);
and U9441 (N_9441,N_3791,N_5848);
nor U9442 (N_9442,N_3378,N_819);
nor U9443 (N_9443,N_1213,N_875);
and U9444 (N_9444,N_648,N_226);
and U9445 (N_9445,N_4719,N_1415);
and U9446 (N_9446,N_1672,N_1345);
or U9447 (N_9447,N_1533,N_4025);
and U9448 (N_9448,N_1255,N_4192);
and U9449 (N_9449,N_1938,N_5962);
nand U9450 (N_9450,N_922,N_233);
or U9451 (N_9451,N_5859,N_5276);
and U9452 (N_9452,N_312,N_5663);
or U9453 (N_9453,N_1304,N_3358);
nand U9454 (N_9454,N_2166,N_1161);
and U9455 (N_9455,N_3146,N_4583);
nor U9456 (N_9456,N_3736,N_3256);
xor U9457 (N_9457,N_1433,N_5184);
and U9458 (N_9458,N_6062,N_4708);
nor U9459 (N_9459,N_5435,N_613);
nand U9460 (N_9460,N_4079,N_1184);
nand U9461 (N_9461,N_4057,N_77);
nor U9462 (N_9462,N_1203,N_3887);
nand U9463 (N_9463,N_3980,N_1496);
nand U9464 (N_9464,N_4545,N_1380);
and U9465 (N_9465,N_1603,N_5309);
and U9466 (N_9466,N_6020,N_5364);
and U9467 (N_9467,N_3402,N_4765);
and U9468 (N_9468,N_4412,N_5256);
xnor U9469 (N_9469,N_5683,N_5402);
xnor U9470 (N_9470,N_3451,N_2999);
nor U9471 (N_9471,N_6068,N_5462);
nand U9472 (N_9472,N_2682,N_4388);
nand U9473 (N_9473,N_2245,N_1490);
nor U9474 (N_9474,N_1239,N_1447);
and U9475 (N_9475,N_1898,N_72);
and U9476 (N_9476,N_5810,N_2075);
or U9477 (N_9477,N_6070,N_2043);
and U9478 (N_9478,N_5920,N_2018);
nor U9479 (N_9479,N_3638,N_617);
and U9480 (N_9480,N_100,N_4140);
or U9481 (N_9481,N_1295,N_722);
nand U9482 (N_9482,N_5117,N_1568);
and U9483 (N_9483,N_3361,N_6098);
and U9484 (N_9484,N_3691,N_674);
nand U9485 (N_9485,N_2013,N_3603);
or U9486 (N_9486,N_3447,N_2953);
or U9487 (N_9487,N_5942,N_4915);
xor U9488 (N_9488,N_984,N_2562);
or U9489 (N_9489,N_2586,N_4885);
xnor U9490 (N_9490,N_94,N_3490);
nor U9491 (N_9491,N_1515,N_6099);
and U9492 (N_9492,N_1613,N_730);
nand U9493 (N_9493,N_4092,N_3111);
and U9494 (N_9494,N_3723,N_3228);
nor U9495 (N_9495,N_3984,N_4970);
or U9496 (N_9496,N_3130,N_3084);
and U9497 (N_9497,N_6179,N_3219);
nor U9498 (N_9498,N_3751,N_4177);
nor U9499 (N_9499,N_5355,N_1229);
nor U9500 (N_9500,N_4200,N_3105);
xor U9501 (N_9501,N_6064,N_477);
nor U9502 (N_9502,N_1990,N_5654);
nor U9503 (N_9503,N_2862,N_253);
nor U9504 (N_9504,N_6237,N_2550);
and U9505 (N_9505,N_1810,N_5241);
nand U9506 (N_9506,N_1101,N_2640);
or U9507 (N_9507,N_2678,N_3767);
or U9508 (N_9508,N_5950,N_2730);
or U9509 (N_9509,N_1435,N_5556);
nand U9510 (N_9510,N_2991,N_4367);
nand U9511 (N_9511,N_5772,N_5513);
xor U9512 (N_9512,N_4665,N_5339);
xor U9513 (N_9513,N_2700,N_603);
and U9514 (N_9514,N_246,N_2291);
nor U9515 (N_9515,N_2960,N_4137);
xnor U9516 (N_9516,N_4582,N_2442);
xor U9517 (N_9517,N_2745,N_2020);
and U9518 (N_9518,N_1709,N_982);
and U9519 (N_9519,N_6192,N_4974);
nor U9520 (N_9520,N_6199,N_4754);
and U9521 (N_9521,N_2756,N_2815);
xnor U9522 (N_9522,N_3768,N_2447);
nor U9523 (N_9523,N_699,N_5788);
nand U9524 (N_9524,N_2249,N_5844);
nand U9525 (N_9525,N_5815,N_198);
xor U9526 (N_9526,N_2299,N_3563);
nand U9527 (N_9527,N_3987,N_4472);
nor U9528 (N_9528,N_1736,N_1384);
or U9529 (N_9529,N_5399,N_4688);
nor U9530 (N_9530,N_3493,N_2106);
nand U9531 (N_9531,N_3810,N_2834);
and U9532 (N_9532,N_702,N_4787);
nor U9533 (N_9533,N_26,N_2536);
or U9534 (N_9534,N_1390,N_5136);
or U9535 (N_9535,N_1798,N_1116);
or U9536 (N_9536,N_958,N_2891);
nand U9537 (N_9537,N_3532,N_1849);
nand U9538 (N_9538,N_707,N_3080);
and U9539 (N_9539,N_366,N_5971);
and U9540 (N_9540,N_1168,N_354);
nand U9541 (N_9541,N_3055,N_2060);
and U9542 (N_9542,N_2217,N_405);
and U9543 (N_9543,N_4450,N_5070);
or U9544 (N_9544,N_3400,N_5987);
and U9545 (N_9545,N_267,N_4151);
nand U9546 (N_9546,N_4531,N_382);
or U9547 (N_9547,N_950,N_6024);
and U9548 (N_9548,N_4270,N_4103);
or U9549 (N_9549,N_1402,N_244);
or U9550 (N_9550,N_406,N_818);
nor U9551 (N_9551,N_1223,N_3338);
nand U9552 (N_9552,N_4173,N_5318);
nor U9553 (N_9553,N_1070,N_2191);
xnor U9554 (N_9554,N_2566,N_2233);
nor U9555 (N_9555,N_5363,N_4380);
and U9556 (N_9556,N_2436,N_5014);
nand U9557 (N_9557,N_4301,N_4451);
or U9558 (N_9558,N_286,N_2975);
or U9559 (N_9559,N_698,N_1301);
nor U9560 (N_9560,N_1821,N_633);
nor U9561 (N_9561,N_3819,N_4353);
and U9562 (N_9562,N_4740,N_3394);
or U9563 (N_9563,N_454,N_2497);
xnor U9564 (N_9564,N_1098,N_1181);
nand U9565 (N_9565,N_49,N_5485);
xnor U9566 (N_9566,N_1467,N_3115);
and U9567 (N_9567,N_1035,N_5862);
nor U9568 (N_9568,N_4852,N_222);
nor U9569 (N_9569,N_6172,N_3157);
or U9570 (N_9570,N_1650,N_226);
and U9571 (N_9571,N_4555,N_3686);
or U9572 (N_9572,N_5619,N_526);
xor U9573 (N_9573,N_868,N_5799);
nor U9574 (N_9574,N_4814,N_4913);
nand U9575 (N_9575,N_284,N_1846);
nor U9576 (N_9576,N_3806,N_1463);
and U9577 (N_9577,N_520,N_3957);
and U9578 (N_9578,N_3566,N_439);
and U9579 (N_9579,N_3364,N_4067);
nor U9580 (N_9580,N_1025,N_1443);
or U9581 (N_9581,N_3247,N_6161);
and U9582 (N_9582,N_3819,N_4256);
xnor U9583 (N_9583,N_754,N_288);
xor U9584 (N_9584,N_1175,N_5906);
and U9585 (N_9585,N_2525,N_15);
xnor U9586 (N_9586,N_1873,N_2765);
nor U9587 (N_9587,N_3529,N_3934);
or U9588 (N_9588,N_2420,N_5088);
xnor U9589 (N_9589,N_3833,N_1780);
nand U9590 (N_9590,N_2249,N_2552);
or U9591 (N_9591,N_3190,N_421);
nand U9592 (N_9592,N_4400,N_1554);
xor U9593 (N_9593,N_5717,N_3869);
nor U9594 (N_9594,N_2243,N_2802);
nand U9595 (N_9595,N_154,N_1029);
xnor U9596 (N_9596,N_5699,N_1703);
and U9597 (N_9597,N_1962,N_4155);
xnor U9598 (N_9598,N_5029,N_3497);
nor U9599 (N_9599,N_3222,N_1887);
nor U9600 (N_9600,N_2057,N_4660);
or U9601 (N_9601,N_5068,N_403);
nor U9602 (N_9602,N_6071,N_5032);
xnor U9603 (N_9603,N_213,N_2823);
nor U9604 (N_9604,N_380,N_1943);
nand U9605 (N_9605,N_4440,N_3893);
nor U9606 (N_9606,N_3697,N_5755);
and U9607 (N_9607,N_4518,N_566);
nor U9608 (N_9608,N_1256,N_600);
nand U9609 (N_9609,N_4039,N_1367);
xnor U9610 (N_9610,N_4420,N_1444);
and U9611 (N_9611,N_111,N_6037);
nor U9612 (N_9612,N_5215,N_388);
nor U9613 (N_9613,N_777,N_3391);
and U9614 (N_9614,N_601,N_53);
and U9615 (N_9615,N_2911,N_3762);
xnor U9616 (N_9616,N_5536,N_3325);
or U9617 (N_9617,N_5232,N_4600);
xor U9618 (N_9618,N_2560,N_876);
nor U9619 (N_9619,N_2612,N_3027);
nor U9620 (N_9620,N_828,N_3976);
nand U9621 (N_9621,N_3255,N_5659);
nor U9622 (N_9622,N_3002,N_1565);
nand U9623 (N_9623,N_6013,N_56);
xor U9624 (N_9624,N_1783,N_2587);
or U9625 (N_9625,N_661,N_863);
nand U9626 (N_9626,N_166,N_3579);
nand U9627 (N_9627,N_6047,N_3216);
xor U9628 (N_9628,N_3179,N_2321);
xnor U9629 (N_9629,N_4646,N_3297);
nor U9630 (N_9630,N_2409,N_5532);
nor U9631 (N_9631,N_1114,N_3792);
and U9632 (N_9632,N_4189,N_5675);
and U9633 (N_9633,N_2749,N_2402);
nand U9634 (N_9634,N_4800,N_4452);
nor U9635 (N_9635,N_75,N_226);
xnor U9636 (N_9636,N_2396,N_3400);
nor U9637 (N_9637,N_5892,N_5226);
nand U9638 (N_9638,N_5085,N_1606);
or U9639 (N_9639,N_4658,N_5169);
nor U9640 (N_9640,N_562,N_4077);
and U9641 (N_9641,N_4502,N_452);
nor U9642 (N_9642,N_4369,N_785);
and U9643 (N_9643,N_2357,N_394);
xnor U9644 (N_9644,N_1589,N_2713);
and U9645 (N_9645,N_5452,N_1255);
nand U9646 (N_9646,N_704,N_3577);
or U9647 (N_9647,N_1189,N_5910);
nor U9648 (N_9648,N_3471,N_211);
or U9649 (N_9649,N_434,N_1661);
and U9650 (N_9650,N_5493,N_4991);
or U9651 (N_9651,N_2965,N_5536);
xnor U9652 (N_9652,N_6167,N_1497);
or U9653 (N_9653,N_4974,N_3340);
and U9654 (N_9654,N_5144,N_1862);
and U9655 (N_9655,N_6044,N_5372);
nand U9656 (N_9656,N_2970,N_4657);
nand U9657 (N_9657,N_1562,N_3061);
nor U9658 (N_9658,N_6188,N_5476);
xnor U9659 (N_9659,N_2877,N_5856);
and U9660 (N_9660,N_3578,N_6194);
or U9661 (N_9661,N_5092,N_5160);
and U9662 (N_9662,N_5660,N_845);
nand U9663 (N_9663,N_775,N_5191);
xor U9664 (N_9664,N_848,N_5005);
nand U9665 (N_9665,N_5994,N_5031);
xor U9666 (N_9666,N_1015,N_3298);
and U9667 (N_9667,N_4642,N_2928);
or U9668 (N_9668,N_96,N_63);
nor U9669 (N_9669,N_1786,N_6072);
nor U9670 (N_9670,N_1346,N_3768);
nand U9671 (N_9671,N_3337,N_5081);
nor U9672 (N_9672,N_2461,N_5531);
and U9673 (N_9673,N_4534,N_2082);
nor U9674 (N_9674,N_3347,N_3840);
nor U9675 (N_9675,N_34,N_6166);
xor U9676 (N_9676,N_3583,N_5523);
xnor U9677 (N_9677,N_4804,N_5874);
and U9678 (N_9678,N_2828,N_1366);
or U9679 (N_9679,N_4446,N_310);
or U9680 (N_9680,N_3669,N_5310);
nor U9681 (N_9681,N_937,N_2611);
or U9682 (N_9682,N_3987,N_4550);
and U9683 (N_9683,N_4295,N_6108);
nand U9684 (N_9684,N_5674,N_5912);
nor U9685 (N_9685,N_2443,N_4394);
nand U9686 (N_9686,N_4380,N_311);
xnor U9687 (N_9687,N_2065,N_4680);
or U9688 (N_9688,N_3709,N_3646);
nor U9689 (N_9689,N_5709,N_1185);
nor U9690 (N_9690,N_5584,N_609);
and U9691 (N_9691,N_5244,N_1694);
nand U9692 (N_9692,N_1377,N_1965);
xor U9693 (N_9693,N_1079,N_2179);
nor U9694 (N_9694,N_4041,N_2082);
xnor U9695 (N_9695,N_1436,N_3811);
xnor U9696 (N_9696,N_2857,N_4559);
nand U9697 (N_9697,N_5862,N_6002);
or U9698 (N_9698,N_3420,N_1175);
nor U9699 (N_9699,N_5040,N_4233);
or U9700 (N_9700,N_4161,N_3068);
and U9701 (N_9701,N_823,N_5329);
and U9702 (N_9702,N_5691,N_6249);
and U9703 (N_9703,N_284,N_3545);
nand U9704 (N_9704,N_1780,N_503);
xnor U9705 (N_9705,N_1565,N_2420);
nor U9706 (N_9706,N_2889,N_226);
nand U9707 (N_9707,N_5439,N_735);
or U9708 (N_9708,N_2517,N_2851);
or U9709 (N_9709,N_3317,N_1118);
nand U9710 (N_9710,N_5785,N_3001);
xor U9711 (N_9711,N_3856,N_2749);
nor U9712 (N_9712,N_5790,N_6143);
xnor U9713 (N_9713,N_2948,N_4926);
xnor U9714 (N_9714,N_3017,N_20);
xor U9715 (N_9715,N_1704,N_2344);
nor U9716 (N_9716,N_6234,N_2608);
xor U9717 (N_9717,N_3358,N_4759);
nand U9718 (N_9718,N_307,N_6186);
nand U9719 (N_9719,N_312,N_880);
or U9720 (N_9720,N_2468,N_2352);
nor U9721 (N_9721,N_85,N_4635);
and U9722 (N_9722,N_1434,N_1238);
nor U9723 (N_9723,N_2257,N_4527);
or U9724 (N_9724,N_589,N_1490);
nor U9725 (N_9725,N_2096,N_2104);
xnor U9726 (N_9726,N_4732,N_5173);
xor U9727 (N_9727,N_922,N_1952);
nor U9728 (N_9728,N_3543,N_5059);
or U9729 (N_9729,N_3423,N_1565);
or U9730 (N_9730,N_2592,N_2559);
or U9731 (N_9731,N_3737,N_3819);
or U9732 (N_9732,N_842,N_5836);
and U9733 (N_9733,N_3995,N_2847);
and U9734 (N_9734,N_5151,N_619);
and U9735 (N_9735,N_711,N_2175);
xor U9736 (N_9736,N_1696,N_420);
nand U9737 (N_9737,N_5761,N_4365);
or U9738 (N_9738,N_145,N_3843);
xnor U9739 (N_9739,N_1979,N_175);
nand U9740 (N_9740,N_4226,N_2893);
nand U9741 (N_9741,N_3563,N_3653);
xnor U9742 (N_9742,N_2918,N_2845);
xor U9743 (N_9743,N_5102,N_5783);
or U9744 (N_9744,N_4980,N_4819);
nand U9745 (N_9745,N_2275,N_3858);
nand U9746 (N_9746,N_875,N_2930);
or U9747 (N_9747,N_1598,N_5143);
and U9748 (N_9748,N_4979,N_3506);
or U9749 (N_9749,N_1755,N_2127);
and U9750 (N_9750,N_522,N_4722);
or U9751 (N_9751,N_2314,N_3926);
xor U9752 (N_9752,N_4103,N_2775);
xnor U9753 (N_9753,N_4337,N_2115);
nor U9754 (N_9754,N_4302,N_755);
or U9755 (N_9755,N_1980,N_2570);
nand U9756 (N_9756,N_885,N_31);
and U9757 (N_9757,N_1186,N_4989);
xnor U9758 (N_9758,N_4083,N_5286);
or U9759 (N_9759,N_4302,N_3355);
xor U9760 (N_9760,N_2501,N_2235);
nor U9761 (N_9761,N_5772,N_3927);
nand U9762 (N_9762,N_2671,N_586);
and U9763 (N_9763,N_5084,N_2023);
and U9764 (N_9764,N_1807,N_3987);
and U9765 (N_9765,N_5240,N_5660);
xnor U9766 (N_9766,N_5626,N_1231);
and U9767 (N_9767,N_2984,N_4429);
or U9768 (N_9768,N_5125,N_3294);
or U9769 (N_9769,N_4157,N_1842);
xnor U9770 (N_9770,N_2868,N_4274);
nand U9771 (N_9771,N_3249,N_5885);
nor U9772 (N_9772,N_1651,N_4342);
or U9773 (N_9773,N_5383,N_623);
xnor U9774 (N_9774,N_3293,N_4943);
and U9775 (N_9775,N_463,N_3199);
and U9776 (N_9776,N_5566,N_5866);
nor U9777 (N_9777,N_921,N_5416);
nand U9778 (N_9778,N_4126,N_594);
and U9779 (N_9779,N_131,N_5405);
nor U9780 (N_9780,N_2977,N_2312);
and U9781 (N_9781,N_4575,N_18);
and U9782 (N_9782,N_2072,N_1928);
and U9783 (N_9783,N_4888,N_5928);
and U9784 (N_9784,N_2302,N_1227);
xor U9785 (N_9785,N_5229,N_2651);
nand U9786 (N_9786,N_2122,N_3622);
nor U9787 (N_9787,N_540,N_1500);
and U9788 (N_9788,N_3710,N_4936);
xnor U9789 (N_9789,N_537,N_1730);
nor U9790 (N_9790,N_5219,N_5899);
nand U9791 (N_9791,N_1592,N_5181);
xnor U9792 (N_9792,N_1606,N_2164);
nor U9793 (N_9793,N_5013,N_6064);
nand U9794 (N_9794,N_4311,N_5334);
and U9795 (N_9795,N_6153,N_3917);
and U9796 (N_9796,N_3809,N_1227);
xnor U9797 (N_9797,N_4026,N_4175);
xnor U9798 (N_9798,N_5702,N_350);
or U9799 (N_9799,N_4326,N_1010);
nor U9800 (N_9800,N_674,N_5267);
xnor U9801 (N_9801,N_3278,N_5345);
nor U9802 (N_9802,N_4526,N_6165);
nor U9803 (N_9803,N_6073,N_4108);
nand U9804 (N_9804,N_5019,N_2847);
or U9805 (N_9805,N_2355,N_3285);
xnor U9806 (N_9806,N_3592,N_4120);
and U9807 (N_9807,N_953,N_1803);
xnor U9808 (N_9808,N_1078,N_3480);
nand U9809 (N_9809,N_5023,N_4694);
xor U9810 (N_9810,N_4385,N_1450);
nand U9811 (N_9811,N_1975,N_6053);
or U9812 (N_9812,N_1336,N_3535);
or U9813 (N_9813,N_4449,N_3162);
and U9814 (N_9814,N_949,N_1230);
or U9815 (N_9815,N_3058,N_4993);
or U9816 (N_9816,N_1586,N_654);
nand U9817 (N_9817,N_4578,N_3724);
and U9818 (N_9818,N_3327,N_3924);
or U9819 (N_9819,N_1027,N_320);
xnor U9820 (N_9820,N_4155,N_4393);
nor U9821 (N_9821,N_2185,N_2248);
nand U9822 (N_9822,N_4575,N_5811);
or U9823 (N_9823,N_1892,N_6138);
nor U9824 (N_9824,N_4789,N_6168);
xnor U9825 (N_9825,N_3791,N_6058);
nand U9826 (N_9826,N_1383,N_1522);
and U9827 (N_9827,N_1432,N_3363);
or U9828 (N_9828,N_1672,N_2765);
and U9829 (N_9829,N_1627,N_6159);
nand U9830 (N_9830,N_5392,N_4493);
or U9831 (N_9831,N_4163,N_6008);
or U9832 (N_9832,N_3920,N_2359);
nand U9833 (N_9833,N_3411,N_908);
and U9834 (N_9834,N_5059,N_4533);
nand U9835 (N_9835,N_5126,N_706);
or U9836 (N_9836,N_4349,N_2101);
or U9837 (N_9837,N_1566,N_3769);
nand U9838 (N_9838,N_5483,N_4997);
or U9839 (N_9839,N_1572,N_4138);
nor U9840 (N_9840,N_3218,N_4680);
and U9841 (N_9841,N_1344,N_1534);
and U9842 (N_9842,N_5484,N_2712);
nor U9843 (N_9843,N_1348,N_908);
xnor U9844 (N_9844,N_2137,N_5428);
nor U9845 (N_9845,N_69,N_2816);
nand U9846 (N_9846,N_5223,N_4121);
and U9847 (N_9847,N_5174,N_2206);
or U9848 (N_9848,N_3523,N_1595);
or U9849 (N_9849,N_3570,N_4499);
nor U9850 (N_9850,N_2753,N_4031);
nand U9851 (N_9851,N_5156,N_4142);
and U9852 (N_9852,N_1244,N_5652);
nor U9853 (N_9853,N_455,N_407);
xnor U9854 (N_9854,N_4204,N_415);
or U9855 (N_9855,N_787,N_5902);
nor U9856 (N_9856,N_818,N_1465);
nand U9857 (N_9857,N_1073,N_410);
nor U9858 (N_9858,N_4041,N_1480);
and U9859 (N_9859,N_2112,N_4353);
xor U9860 (N_9860,N_5459,N_5321);
nand U9861 (N_9861,N_553,N_3007);
nor U9862 (N_9862,N_3287,N_3575);
nand U9863 (N_9863,N_5837,N_1950);
xnor U9864 (N_9864,N_94,N_5946);
and U9865 (N_9865,N_1213,N_3524);
and U9866 (N_9866,N_488,N_2518);
nor U9867 (N_9867,N_2029,N_2287);
or U9868 (N_9868,N_471,N_3190);
xor U9869 (N_9869,N_4420,N_3232);
or U9870 (N_9870,N_3495,N_5002);
and U9871 (N_9871,N_3657,N_4819);
nor U9872 (N_9872,N_869,N_551);
and U9873 (N_9873,N_4112,N_5922);
nor U9874 (N_9874,N_160,N_107);
xnor U9875 (N_9875,N_4235,N_3232);
nand U9876 (N_9876,N_1278,N_4814);
xnor U9877 (N_9877,N_2770,N_1391);
and U9878 (N_9878,N_1193,N_2410);
or U9879 (N_9879,N_4650,N_2203);
xor U9880 (N_9880,N_4160,N_1454);
nor U9881 (N_9881,N_47,N_463);
and U9882 (N_9882,N_3471,N_1143);
nand U9883 (N_9883,N_4507,N_3841);
nor U9884 (N_9884,N_1990,N_3562);
or U9885 (N_9885,N_4749,N_5404);
nor U9886 (N_9886,N_5689,N_1582);
nand U9887 (N_9887,N_3476,N_2115);
nor U9888 (N_9888,N_807,N_2403);
nand U9889 (N_9889,N_2969,N_5747);
nor U9890 (N_9890,N_3253,N_5478);
nand U9891 (N_9891,N_3709,N_3121);
xor U9892 (N_9892,N_3985,N_4712);
or U9893 (N_9893,N_4816,N_952);
nand U9894 (N_9894,N_5353,N_4304);
xnor U9895 (N_9895,N_684,N_4553);
xor U9896 (N_9896,N_5084,N_1730);
or U9897 (N_9897,N_5282,N_5602);
xnor U9898 (N_9898,N_2532,N_5108);
nor U9899 (N_9899,N_4348,N_1831);
or U9900 (N_9900,N_3480,N_1639);
and U9901 (N_9901,N_2485,N_5450);
nand U9902 (N_9902,N_4307,N_1491);
xnor U9903 (N_9903,N_393,N_5332);
nand U9904 (N_9904,N_2142,N_3368);
and U9905 (N_9905,N_1371,N_5065);
nand U9906 (N_9906,N_6022,N_6082);
xor U9907 (N_9907,N_3140,N_822);
xor U9908 (N_9908,N_455,N_1376);
nor U9909 (N_9909,N_3422,N_4519);
nor U9910 (N_9910,N_5806,N_1080);
or U9911 (N_9911,N_5280,N_3601);
and U9912 (N_9912,N_4033,N_136);
nand U9913 (N_9913,N_2367,N_1580);
xnor U9914 (N_9914,N_5312,N_4713);
xnor U9915 (N_9915,N_94,N_5810);
nand U9916 (N_9916,N_3729,N_3356);
nand U9917 (N_9917,N_5871,N_4634);
xor U9918 (N_9918,N_4839,N_4292);
nand U9919 (N_9919,N_5611,N_3127);
and U9920 (N_9920,N_3381,N_1443);
or U9921 (N_9921,N_6029,N_2121);
nand U9922 (N_9922,N_5040,N_3776);
nand U9923 (N_9923,N_1816,N_3146);
nor U9924 (N_9924,N_4396,N_4467);
xor U9925 (N_9925,N_3080,N_1089);
xor U9926 (N_9926,N_1145,N_2063);
nor U9927 (N_9927,N_2366,N_2948);
nor U9928 (N_9928,N_4295,N_3590);
nand U9929 (N_9929,N_1766,N_5106);
xor U9930 (N_9930,N_1912,N_5325);
and U9931 (N_9931,N_4255,N_5482);
and U9932 (N_9932,N_2242,N_5296);
nand U9933 (N_9933,N_3773,N_5461);
nor U9934 (N_9934,N_2825,N_4027);
xnor U9935 (N_9935,N_1015,N_4605);
and U9936 (N_9936,N_695,N_1668);
nand U9937 (N_9937,N_465,N_4153);
nor U9938 (N_9938,N_1044,N_1138);
or U9939 (N_9939,N_1174,N_3812);
or U9940 (N_9940,N_4337,N_2713);
and U9941 (N_9941,N_4094,N_1450);
xor U9942 (N_9942,N_3675,N_820);
xor U9943 (N_9943,N_4887,N_3995);
or U9944 (N_9944,N_70,N_4447);
xor U9945 (N_9945,N_3737,N_2505);
and U9946 (N_9946,N_2904,N_2054);
nand U9947 (N_9947,N_17,N_4682);
or U9948 (N_9948,N_963,N_3428);
nand U9949 (N_9949,N_3167,N_5090);
nand U9950 (N_9950,N_538,N_2013);
nor U9951 (N_9951,N_1671,N_44);
nand U9952 (N_9952,N_5811,N_4630);
xor U9953 (N_9953,N_2552,N_4071);
and U9954 (N_9954,N_4863,N_5420);
and U9955 (N_9955,N_3356,N_3862);
xor U9956 (N_9956,N_3548,N_1823);
nand U9957 (N_9957,N_788,N_2688);
and U9958 (N_9958,N_5038,N_3826);
and U9959 (N_9959,N_6224,N_3667);
nor U9960 (N_9960,N_177,N_5294);
nor U9961 (N_9961,N_926,N_1227);
xor U9962 (N_9962,N_1056,N_1570);
or U9963 (N_9963,N_2199,N_3645);
xnor U9964 (N_9964,N_3569,N_3987);
xnor U9965 (N_9965,N_5391,N_846);
nor U9966 (N_9966,N_3801,N_5952);
xor U9967 (N_9967,N_5722,N_2047);
nor U9968 (N_9968,N_3279,N_6066);
or U9969 (N_9969,N_247,N_711);
or U9970 (N_9970,N_2325,N_3732);
nand U9971 (N_9971,N_3892,N_5724);
nor U9972 (N_9972,N_4849,N_6248);
and U9973 (N_9973,N_1334,N_3388);
nand U9974 (N_9974,N_5008,N_2278);
nand U9975 (N_9975,N_261,N_4587);
nor U9976 (N_9976,N_492,N_2449);
and U9977 (N_9977,N_4400,N_612);
nor U9978 (N_9978,N_2061,N_4364);
or U9979 (N_9979,N_2448,N_4367);
xnor U9980 (N_9980,N_1752,N_4669);
xor U9981 (N_9981,N_4898,N_3889);
nor U9982 (N_9982,N_2845,N_1669);
or U9983 (N_9983,N_2112,N_1675);
xnor U9984 (N_9984,N_2457,N_2710);
xnor U9985 (N_9985,N_3991,N_1047);
xnor U9986 (N_9986,N_678,N_1672);
or U9987 (N_9987,N_1017,N_1014);
and U9988 (N_9988,N_2573,N_3416);
nand U9989 (N_9989,N_817,N_167);
nor U9990 (N_9990,N_1450,N_5290);
xnor U9991 (N_9991,N_3601,N_3207);
nand U9992 (N_9992,N_1240,N_3256);
and U9993 (N_9993,N_86,N_3176);
nor U9994 (N_9994,N_3726,N_1636);
nand U9995 (N_9995,N_1790,N_1701);
nand U9996 (N_9996,N_1560,N_5399);
nand U9997 (N_9997,N_4983,N_3047);
xor U9998 (N_9998,N_1045,N_2663);
nor U9999 (N_9999,N_3354,N_4684);
or U10000 (N_10000,N_927,N_616);
or U10001 (N_10001,N_5383,N_5920);
nor U10002 (N_10002,N_5279,N_1020);
or U10003 (N_10003,N_5970,N_631);
nor U10004 (N_10004,N_510,N_5010);
nor U10005 (N_10005,N_1297,N_5157);
xnor U10006 (N_10006,N_4776,N_5719);
nor U10007 (N_10007,N_1397,N_5514);
nand U10008 (N_10008,N_1141,N_3349);
xnor U10009 (N_10009,N_237,N_4314);
xor U10010 (N_10010,N_135,N_2999);
and U10011 (N_10011,N_2679,N_4228);
nor U10012 (N_10012,N_169,N_1273);
and U10013 (N_10013,N_3539,N_4221);
nand U10014 (N_10014,N_6202,N_1847);
xnor U10015 (N_10015,N_317,N_4217);
or U10016 (N_10016,N_5921,N_4590);
and U10017 (N_10017,N_470,N_3605);
nand U10018 (N_10018,N_812,N_1010);
and U10019 (N_10019,N_5739,N_6229);
nor U10020 (N_10020,N_3778,N_652);
or U10021 (N_10021,N_5314,N_2555);
or U10022 (N_10022,N_5896,N_4571);
xor U10023 (N_10023,N_5434,N_465);
nor U10024 (N_10024,N_1034,N_1478);
nand U10025 (N_10025,N_1620,N_2166);
or U10026 (N_10026,N_3836,N_901);
xnor U10027 (N_10027,N_4777,N_1774);
and U10028 (N_10028,N_2401,N_484);
xnor U10029 (N_10029,N_2207,N_5614);
nor U10030 (N_10030,N_3491,N_877);
xor U10031 (N_10031,N_4075,N_753);
nand U10032 (N_10032,N_4139,N_634);
nand U10033 (N_10033,N_5992,N_1423);
nand U10034 (N_10034,N_5168,N_3071);
or U10035 (N_10035,N_1477,N_1755);
or U10036 (N_10036,N_1095,N_444);
nand U10037 (N_10037,N_3256,N_838);
nor U10038 (N_10038,N_5988,N_1626);
or U10039 (N_10039,N_786,N_1583);
nor U10040 (N_10040,N_3874,N_4331);
xnor U10041 (N_10041,N_3729,N_118);
and U10042 (N_10042,N_1679,N_1304);
xnor U10043 (N_10043,N_1694,N_1330);
nor U10044 (N_10044,N_5688,N_3083);
nor U10045 (N_10045,N_3280,N_1036);
or U10046 (N_10046,N_1464,N_1148);
and U10047 (N_10047,N_4717,N_2264);
nand U10048 (N_10048,N_2889,N_2561);
and U10049 (N_10049,N_1276,N_746);
nor U10050 (N_10050,N_5480,N_5235);
and U10051 (N_10051,N_5814,N_2398);
nor U10052 (N_10052,N_4682,N_2662);
xnor U10053 (N_10053,N_2192,N_2776);
nor U10054 (N_10054,N_5886,N_4892);
nor U10055 (N_10055,N_1175,N_3596);
and U10056 (N_10056,N_1991,N_745);
xnor U10057 (N_10057,N_1327,N_174);
xnor U10058 (N_10058,N_2141,N_1097);
or U10059 (N_10059,N_333,N_2613);
nor U10060 (N_10060,N_1092,N_564);
nand U10061 (N_10061,N_6135,N_2710);
xor U10062 (N_10062,N_162,N_2456);
nor U10063 (N_10063,N_1118,N_967);
and U10064 (N_10064,N_1637,N_2287);
or U10065 (N_10065,N_5944,N_931);
nand U10066 (N_10066,N_4887,N_1241);
nand U10067 (N_10067,N_3575,N_3230);
nand U10068 (N_10068,N_1553,N_188);
xor U10069 (N_10069,N_5469,N_5496);
nand U10070 (N_10070,N_2785,N_431);
xor U10071 (N_10071,N_3035,N_2031);
and U10072 (N_10072,N_2378,N_6113);
or U10073 (N_10073,N_3752,N_466);
xnor U10074 (N_10074,N_1005,N_1044);
and U10075 (N_10075,N_3641,N_636);
or U10076 (N_10076,N_393,N_367);
xnor U10077 (N_10077,N_4519,N_190);
nand U10078 (N_10078,N_4156,N_2827);
or U10079 (N_10079,N_1587,N_3192);
nand U10080 (N_10080,N_1554,N_2506);
and U10081 (N_10081,N_2781,N_1605);
and U10082 (N_10082,N_3980,N_121);
nand U10083 (N_10083,N_2805,N_2725);
xor U10084 (N_10084,N_3601,N_2697);
xor U10085 (N_10085,N_2974,N_434);
xnor U10086 (N_10086,N_267,N_346);
and U10087 (N_10087,N_102,N_1766);
or U10088 (N_10088,N_3757,N_5190);
nand U10089 (N_10089,N_2453,N_2242);
or U10090 (N_10090,N_3310,N_5719);
and U10091 (N_10091,N_4219,N_5630);
and U10092 (N_10092,N_3478,N_6026);
and U10093 (N_10093,N_178,N_3737);
nor U10094 (N_10094,N_5374,N_238);
nor U10095 (N_10095,N_4580,N_950);
or U10096 (N_10096,N_2922,N_233);
nand U10097 (N_10097,N_4708,N_2320);
xnor U10098 (N_10098,N_4596,N_3474);
nor U10099 (N_10099,N_198,N_2708);
or U10100 (N_10100,N_3224,N_2920);
or U10101 (N_10101,N_5857,N_4116);
or U10102 (N_10102,N_948,N_5156);
and U10103 (N_10103,N_587,N_5168);
nor U10104 (N_10104,N_4325,N_5358);
and U10105 (N_10105,N_1605,N_1337);
and U10106 (N_10106,N_4338,N_699);
nor U10107 (N_10107,N_4627,N_3834);
xnor U10108 (N_10108,N_1828,N_370);
nand U10109 (N_10109,N_3665,N_4388);
and U10110 (N_10110,N_1880,N_6112);
xor U10111 (N_10111,N_2469,N_350);
and U10112 (N_10112,N_1227,N_5965);
and U10113 (N_10113,N_1510,N_5939);
nand U10114 (N_10114,N_20,N_4078);
xor U10115 (N_10115,N_224,N_5298);
xor U10116 (N_10116,N_3890,N_3755);
or U10117 (N_10117,N_1526,N_494);
nand U10118 (N_10118,N_4887,N_5980);
nor U10119 (N_10119,N_55,N_635);
or U10120 (N_10120,N_262,N_28);
nor U10121 (N_10121,N_406,N_5316);
or U10122 (N_10122,N_5836,N_1179);
and U10123 (N_10123,N_6218,N_5895);
or U10124 (N_10124,N_4171,N_907);
or U10125 (N_10125,N_2729,N_2364);
xnor U10126 (N_10126,N_1944,N_5073);
xor U10127 (N_10127,N_4460,N_538);
xor U10128 (N_10128,N_2327,N_2817);
nand U10129 (N_10129,N_2454,N_1945);
nor U10130 (N_10130,N_2626,N_2850);
and U10131 (N_10131,N_4874,N_2520);
nor U10132 (N_10132,N_910,N_889);
nor U10133 (N_10133,N_2373,N_6173);
and U10134 (N_10134,N_2567,N_1872);
nand U10135 (N_10135,N_4327,N_885);
and U10136 (N_10136,N_1649,N_2821);
xor U10137 (N_10137,N_1856,N_5518);
or U10138 (N_10138,N_4514,N_5236);
and U10139 (N_10139,N_3653,N_487);
and U10140 (N_10140,N_932,N_1103);
nand U10141 (N_10141,N_5821,N_1176);
or U10142 (N_10142,N_4610,N_4398);
xor U10143 (N_10143,N_168,N_6117);
or U10144 (N_10144,N_3036,N_5366);
nand U10145 (N_10145,N_1944,N_1468);
xor U10146 (N_10146,N_3187,N_5012);
xor U10147 (N_10147,N_3187,N_479);
nor U10148 (N_10148,N_2945,N_2739);
xor U10149 (N_10149,N_1715,N_1299);
xor U10150 (N_10150,N_620,N_3245);
and U10151 (N_10151,N_2187,N_2996);
xor U10152 (N_10152,N_1283,N_1282);
xnor U10153 (N_10153,N_2396,N_3298);
and U10154 (N_10154,N_5777,N_846);
or U10155 (N_10155,N_987,N_1460);
and U10156 (N_10156,N_6127,N_4662);
xor U10157 (N_10157,N_6034,N_4790);
or U10158 (N_10158,N_4837,N_1735);
and U10159 (N_10159,N_3844,N_788);
and U10160 (N_10160,N_3976,N_5404);
xor U10161 (N_10161,N_4582,N_2245);
nor U10162 (N_10162,N_3967,N_2405);
nor U10163 (N_10163,N_3521,N_4809);
nand U10164 (N_10164,N_4845,N_265);
or U10165 (N_10165,N_4592,N_5148);
nor U10166 (N_10166,N_5738,N_1381);
nor U10167 (N_10167,N_3910,N_5765);
nand U10168 (N_10168,N_3613,N_4384);
nor U10169 (N_10169,N_3540,N_477);
or U10170 (N_10170,N_3872,N_2336);
xnor U10171 (N_10171,N_494,N_2461);
nand U10172 (N_10172,N_1688,N_5199);
and U10173 (N_10173,N_5234,N_3432);
nand U10174 (N_10174,N_1958,N_1518);
nand U10175 (N_10175,N_3747,N_3934);
nor U10176 (N_10176,N_547,N_5830);
xor U10177 (N_10177,N_5152,N_1762);
nor U10178 (N_10178,N_4326,N_3031);
xor U10179 (N_10179,N_5751,N_5254);
and U10180 (N_10180,N_3744,N_2054);
or U10181 (N_10181,N_4629,N_4411);
or U10182 (N_10182,N_2320,N_2439);
and U10183 (N_10183,N_2847,N_5091);
nand U10184 (N_10184,N_5092,N_5);
nor U10185 (N_10185,N_4616,N_5849);
and U10186 (N_10186,N_3334,N_2216);
nand U10187 (N_10187,N_154,N_5754);
or U10188 (N_10188,N_4255,N_4892);
nand U10189 (N_10189,N_1649,N_1890);
nor U10190 (N_10190,N_5683,N_188);
xnor U10191 (N_10191,N_3705,N_1539);
xnor U10192 (N_10192,N_5527,N_744);
and U10193 (N_10193,N_2957,N_4675);
and U10194 (N_10194,N_3294,N_953);
nor U10195 (N_10195,N_5619,N_2842);
xnor U10196 (N_10196,N_4067,N_6046);
or U10197 (N_10197,N_4194,N_2258);
nand U10198 (N_10198,N_3463,N_2805);
nand U10199 (N_10199,N_2935,N_5369);
nor U10200 (N_10200,N_1376,N_5246);
or U10201 (N_10201,N_5605,N_3482);
and U10202 (N_10202,N_4757,N_1102);
nand U10203 (N_10203,N_6035,N_1295);
or U10204 (N_10204,N_4928,N_4023);
and U10205 (N_10205,N_2273,N_3587);
and U10206 (N_10206,N_2140,N_1566);
nor U10207 (N_10207,N_5286,N_1187);
and U10208 (N_10208,N_5971,N_5945);
and U10209 (N_10209,N_4475,N_3828);
nor U10210 (N_10210,N_300,N_2445);
nand U10211 (N_10211,N_2451,N_620);
xnor U10212 (N_10212,N_2763,N_2441);
nor U10213 (N_10213,N_6195,N_5744);
and U10214 (N_10214,N_4139,N_511);
nand U10215 (N_10215,N_2019,N_3521);
nand U10216 (N_10216,N_902,N_165);
or U10217 (N_10217,N_2047,N_1207);
and U10218 (N_10218,N_3691,N_2689);
nand U10219 (N_10219,N_1780,N_4732);
nand U10220 (N_10220,N_4060,N_5447);
nor U10221 (N_10221,N_3790,N_1866);
xnor U10222 (N_10222,N_5388,N_2333);
and U10223 (N_10223,N_3158,N_210);
nand U10224 (N_10224,N_3592,N_3378);
and U10225 (N_10225,N_1282,N_2253);
or U10226 (N_10226,N_1357,N_5111);
nand U10227 (N_10227,N_5459,N_6174);
xor U10228 (N_10228,N_3062,N_209);
xnor U10229 (N_10229,N_3314,N_5641);
or U10230 (N_10230,N_3747,N_2977);
and U10231 (N_10231,N_4180,N_1588);
xnor U10232 (N_10232,N_2142,N_4190);
and U10233 (N_10233,N_690,N_6070);
or U10234 (N_10234,N_4334,N_4283);
or U10235 (N_10235,N_5462,N_4761);
xor U10236 (N_10236,N_1564,N_1199);
nor U10237 (N_10237,N_1461,N_1643);
or U10238 (N_10238,N_4684,N_4698);
nor U10239 (N_10239,N_5645,N_4658);
xor U10240 (N_10240,N_3392,N_11);
nor U10241 (N_10241,N_1087,N_2187);
nor U10242 (N_10242,N_4748,N_1675);
and U10243 (N_10243,N_6110,N_3952);
xnor U10244 (N_10244,N_145,N_1005);
xor U10245 (N_10245,N_2471,N_4636);
xor U10246 (N_10246,N_5735,N_2740);
or U10247 (N_10247,N_408,N_416);
nor U10248 (N_10248,N_3139,N_3534);
nor U10249 (N_10249,N_172,N_4499);
xor U10250 (N_10250,N_142,N_723);
or U10251 (N_10251,N_3459,N_4472);
nand U10252 (N_10252,N_5422,N_4696);
nor U10253 (N_10253,N_5400,N_3018);
nor U10254 (N_10254,N_1416,N_1531);
or U10255 (N_10255,N_1158,N_4355);
nand U10256 (N_10256,N_3495,N_2847);
nor U10257 (N_10257,N_3813,N_3297);
xnor U10258 (N_10258,N_2558,N_942);
xor U10259 (N_10259,N_268,N_4907);
or U10260 (N_10260,N_2023,N_3475);
and U10261 (N_10261,N_3898,N_1238);
or U10262 (N_10262,N_1505,N_6233);
nand U10263 (N_10263,N_5107,N_4970);
nor U10264 (N_10264,N_6094,N_1653);
and U10265 (N_10265,N_3102,N_4230);
or U10266 (N_10266,N_1258,N_2897);
xnor U10267 (N_10267,N_208,N_789);
nand U10268 (N_10268,N_2442,N_772);
and U10269 (N_10269,N_875,N_3610);
and U10270 (N_10270,N_5123,N_3179);
or U10271 (N_10271,N_1419,N_5237);
or U10272 (N_10272,N_3685,N_5783);
nand U10273 (N_10273,N_5838,N_6001);
and U10274 (N_10274,N_4066,N_2327);
nor U10275 (N_10275,N_2048,N_4077);
xor U10276 (N_10276,N_211,N_5350);
xnor U10277 (N_10277,N_1638,N_3506);
nor U10278 (N_10278,N_3365,N_532);
and U10279 (N_10279,N_1943,N_742);
and U10280 (N_10280,N_5907,N_2484);
and U10281 (N_10281,N_1757,N_440);
nand U10282 (N_10282,N_1496,N_1910);
or U10283 (N_10283,N_3152,N_210);
nand U10284 (N_10284,N_887,N_1660);
xor U10285 (N_10285,N_4078,N_3916);
nand U10286 (N_10286,N_3704,N_4186);
nand U10287 (N_10287,N_1268,N_810);
nand U10288 (N_10288,N_2167,N_5482);
and U10289 (N_10289,N_2685,N_1670);
or U10290 (N_10290,N_5841,N_5278);
nor U10291 (N_10291,N_3036,N_2434);
and U10292 (N_10292,N_4771,N_1824);
xor U10293 (N_10293,N_5892,N_5536);
nand U10294 (N_10294,N_755,N_3571);
and U10295 (N_10295,N_3388,N_5649);
and U10296 (N_10296,N_5559,N_579);
nor U10297 (N_10297,N_1702,N_3842);
and U10298 (N_10298,N_4484,N_3160);
xor U10299 (N_10299,N_3994,N_4696);
or U10300 (N_10300,N_1367,N_267);
nand U10301 (N_10301,N_2121,N_82);
nor U10302 (N_10302,N_3145,N_2601);
or U10303 (N_10303,N_5386,N_2759);
nor U10304 (N_10304,N_1217,N_694);
xnor U10305 (N_10305,N_5386,N_3124);
xor U10306 (N_10306,N_5597,N_768);
or U10307 (N_10307,N_2222,N_682);
xor U10308 (N_10308,N_2832,N_4158);
nor U10309 (N_10309,N_2809,N_5264);
xnor U10310 (N_10310,N_1701,N_4447);
and U10311 (N_10311,N_458,N_5055);
and U10312 (N_10312,N_1661,N_2926);
and U10313 (N_10313,N_3968,N_554);
nor U10314 (N_10314,N_19,N_6013);
and U10315 (N_10315,N_5992,N_3337);
nand U10316 (N_10316,N_989,N_5407);
or U10317 (N_10317,N_4065,N_798);
or U10318 (N_10318,N_2928,N_3584);
nor U10319 (N_10319,N_2845,N_6177);
nand U10320 (N_10320,N_4484,N_1822);
or U10321 (N_10321,N_2244,N_5217);
and U10322 (N_10322,N_93,N_2706);
nor U10323 (N_10323,N_5480,N_2669);
nor U10324 (N_10324,N_6229,N_4576);
nor U10325 (N_10325,N_576,N_1729);
xnor U10326 (N_10326,N_4738,N_3344);
nor U10327 (N_10327,N_2938,N_544);
nor U10328 (N_10328,N_2915,N_4983);
or U10329 (N_10329,N_2415,N_3254);
xnor U10330 (N_10330,N_3750,N_452);
or U10331 (N_10331,N_455,N_3915);
nor U10332 (N_10332,N_250,N_278);
nand U10333 (N_10333,N_5776,N_6085);
and U10334 (N_10334,N_362,N_1528);
or U10335 (N_10335,N_304,N_3812);
nor U10336 (N_10336,N_963,N_5951);
or U10337 (N_10337,N_4943,N_5388);
nor U10338 (N_10338,N_4383,N_6200);
xnor U10339 (N_10339,N_2024,N_2593);
and U10340 (N_10340,N_4391,N_336);
or U10341 (N_10341,N_4401,N_2767);
nand U10342 (N_10342,N_447,N_1717);
xnor U10343 (N_10343,N_1449,N_2759);
nand U10344 (N_10344,N_2082,N_4028);
nand U10345 (N_10345,N_2496,N_1073);
or U10346 (N_10346,N_4001,N_5204);
nor U10347 (N_10347,N_5848,N_760);
xor U10348 (N_10348,N_4638,N_5157);
nor U10349 (N_10349,N_4806,N_2534);
or U10350 (N_10350,N_581,N_4535);
nand U10351 (N_10351,N_604,N_620);
nor U10352 (N_10352,N_3899,N_1827);
nand U10353 (N_10353,N_3445,N_5158);
or U10354 (N_10354,N_439,N_2979);
or U10355 (N_10355,N_5116,N_5218);
xnor U10356 (N_10356,N_927,N_3767);
xor U10357 (N_10357,N_5409,N_1427);
xnor U10358 (N_10358,N_3148,N_5027);
xor U10359 (N_10359,N_5190,N_6080);
or U10360 (N_10360,N_5101,N_1027);
nor U10361 (N_10361,N_1148,N_3722);
and U10362 (N_10362,N_5831,N_5859);
nand U10363 (N_10363,N_6079,N_996);
or U10364 (N_10364,N_3325,N_1215);
nor U10365 (N_10365,N_1890,N_911);
nor U10366 (N_10366,N_4739,N_1410);
or U10367 (N_10367,N_416,N_4145);
or U10368 (N_10368,N_236,N_1083);
nor U10369 (N_10369,N_5367,N_3858);
xor U10370 (N_10370,N_2078,N_445);
and U10371 (N_10371,N_2641,N_5038);
nor U10372 (N_10372,N_1616,N_5184);
nor U10373 (N_10373,N_4565,N_5847);
nand U10374 (N_10374,N_3170,N_2087);
and U10375 (N_10375,N_1382,N_4569);
xnor U10376 (N_10376,N_4918,N_5669);
and U10377 (N_10377,N_3304,N_4157);
nand U10378 (N_10378,N_4047,N_2582);
nand U10379 (N_10379,N_3379,N_5599);
nor U10380 (N_10380,N_1633,N_4975);
or U10381 (N_10381,N_1220,N_5913);
xnor U10382 (N_10382,N_4070,N_4900);
nand U10383 (N_10383,N_2792,N_4009);
nand U10384 (N_10384,N_2159,N_5423);
nand U10385 (N_10385,N_639,N_6185);
nand U10386 (N_10386,N_691,N_4264);
and U10387 (N_10387,N_4803,N_665);
or U10388 (N_10388,N_3647,N_2107);
nand U10389 (N_10389,N_931,N_4391);
and U10390 (N_10390,N_5677,N_1425);
nand U10391 (N_10391,N_1516,N_1280);
and U10392 (N_10392,N_5103,N_5332);
xor U10393 (N_10393,N_5411,N_1796);
xnor U10394 (N_10394,N_3907,N_550);
nand U10395 (N_10395,N_450,N_4950);
or U10396 (N_10396,N_1902,N_1313);
or U10397 (N_10397,N_4709,N_5657);
or U10398 (N_10398,N_787,N_990);
or U10399 (N_10399,N_1464,N_1452);
nand U10400 (N_10400,N_6194,N_5294);
nand U10401 (N_10401,N_5617,N_893);
xor U10402 (N_10402,N_2385,N_3265);
and U10403 (N_10403,N_5371,N_718);
and U10404 (N_10404,N_3990,N_3486);
or U10405 (N_10405,N_4302,N_5291);
nand U10406 (N_10406,N_5872,N_2912);
nand U10407 (N_10407,N_4654,N_1238);
nand U10408 (N_10408,N_1451,N_5648);
nor U10409 (N_10409,N_1624,N_1051);
xor U10410 (N_10410,N_702,N_6026);
xor U10411 (N_10411,N_4800,N_4369);
and U10412 (N_10412,N_5025,N_5803);
nor U10413 (N_10413,N_2015,N_5392);
and U10414 (N_10414,N_3340,N_5386);
nor U10415 (N_10415,N_5637,N_4216);
and U10416 (N_10416,N_2647,N_2492);
xor U10417 (N_10417,N_471,N_4734);
xnor U10418 (N_10418,N_819,N_1688);
nand U10419 (N_10419,N_695,N_805);
nor U10420 (N_10420,N_2950,N_5663);
or U10421 (N_10421,N_2443,N_806);
and U10422 (N_10422,N_3047,N_1873);
and U10423 (N_10423,N_1493,N_2630);
or U10424 (N_10424,N_5460,N_3858);
nand U10425 (N_10425,N_4965,N_2393);
and U10426 (N_10426,N_4845,N_1378);
nand U10427 (N_10427,N_3043,N_3637);
xor U10428 (N_10428,N_3108,N_3410);
and U10429 (N_10429,N_252,N_2739);
or U10430 (N_10430,N_6053,N_531);
nand U10431 (N_10431,N_4341,N_5329);
and U10432 (N_10432,N_3462,N_2773);
or U10433 (N_10433,N_2061,N_5029);
and U10434 (N_10434,N_2553,N_1437);
and U10435 (N_10435,N_2772,N_67);
xnor U10436 (N_10436,N_3354,N_4727);
xor U10437 (N_10437,N_2188,N_1853);
or U10438 (N_10438,N_6121,N_4455);
xnor U10439 (N_10439,N_5910,N_5365);
xor U10440 (N_10440,N_134,N_5171);
and U10441 (N_10441,N_758,N_5116);
or U10442 (N_10442,N_4934,N_3707);
nand U10443 (N_10443,N_5477,N_3296);
nor U10444 (N_10444,N_5250,N_502);
nor U10445 (N_10445,N_1384,N_21);
nand U10446 (N_10446,N_5946,N_657);
or U10447 (N_10447,N_2793,N_1808);
and U10448 (N_10448,N_5798,N_2802);
nor U10449 (N_10449,N_3441,N_3235);
nor U10450 (N_10450,N_1476,N_1626);
or U10451 (N_10451,N_2479,N_2586);
xnor U10452 (N_10452,N_3960,N_5298);
nor U10453 (N_10453,N_1311,N_3256);
nor U10454 (N_10454,N_4850,N_5782);
nand U10455 (N_10455,N_3639,N_1897);
xor U10456 (N_10456,N_2970,N_2079);
and U10457 (N_10457,N_367,N_2334);
nor U10458 (N_10458,N_5642,N_295);
nand U10459 (N_10459,N_3314,N_3500);
xnor U10460 (N_10460,N_4037,N_2225);
nand U10461 (N_10461,N_599,N_1624);
xnor U10462 (N_10462,N_6153,N_260);
or U10463 (N_10463,N_244,N_4838);
and U10464 (N_10464,N_2366,N_3191);
xor U10465 (N_10465,N_4513,N_3963);
xor U10466 (N_10466,N_1486,N_2053);
nor U10467 (N_10467,N_33,N_3990);
nand U10468 (N_10468,N_2445,N_325);
nand U10469 (N_10469,N_2851,N_5194);
xor U10470 (N_10470,N_2373,N_4987);
nand U10471 (N_10471,N_1859,N_1629);
nor U10472 (N_10472,N_3492,N_5915);
nor U10473 (N_10473,N_3296,N_808);
or U10474 (N_10474,N_6149,N_4579);
xnor U10475 (N_10475,N_3623,N_4143);
or U10476 (N_10476,N_6019,N_3737);
nor U10477 (N_10477,N_836,N_90);
nand U10478 (N_10478,N_3764,N_4081);
and U10479 (N_10479,N_5921,N_6014);
nand U10480 (N_10480,N_1984,N_2337);
and U10481 (N_10481,N_3936,N_3038);
nor U10482 (N_10482,N_2822,N_1415);
xor U10483 (N_10483,N_3062,N_3176);
and U10484 (N_10484,N_589,N_4933);
xnor U10485 (N_10485,N_1491,N_5041);
nor U10486 (N_10486,N_2445,N_3480);
or U10487 (N_10487,N_148,N_5038);
or U10488 (N_10488,N_3502,N_3779);
xor U10489 (N_10489,N_81,N_4869);
xnor U10490 (N_10490,N_3445,N_1582);
nand U10491 (N_10491,N_1318,N_2169);
or U10492 (N_10492,N_4621,N_3958);
or U10493 (N_10493,N_1330,N_4004);
nor U10494 (N_10494,N_1576,N_2846);
and U10495 (N_10495,N_844,N_566);
or U10496 (N_10496,N_1873,N_6214);
and U10497 (N_10497,N_4628,N_3934);
and U10498 (N_10498,N_4950,N_4749);
nor U10499 (N_10499,N_2508,N_3224);
and U10500 (N_10500,N_4052,N_2650);
and U10501 (N_10501,N_3976,N_954);
and U10502 (N_10502,N_1391,N_5969);
nor U10503 (N_10503,N_4803,N_5401);
and U10504 (N_10504,N_5575,N_3865);
or U10505 (N_10505,N_3896,N_4746);
and U10506 (N_10506,N_1882,N_4513);
nor U10507 (N_10507,N_1362,N_1188);
nor U10508 (N_10508,N_632,N_4447);
or U10509 (N_10509,N_875,N_3343);
nand U10510 (N_10510,N_2589,N_4172);
and U10511 (N_10511,N_5795,N_4566);
or U10512 (N_10512,N_4432,N_124);
and U10513 (N_10513,N_170,N_888);
or U10514 (N_10514,N_2177,N_412);
or U10515 (N_10515,N_1620,N_4824);
xnor U10516 (N_10516,N_1742,N_4373);
nand U10517 (N_10517,N_4433,N_5004);
or U10518 (N_10518,N_1489,N_6039);
and U10519 (N_10519,N_875,N_4866);
or U10520 (N_10520,N_472,N_5318);
nand U10521 (N_10521,N_5635,N_3392);
nor U10522 (N_10522,N_4149,N_4879);
nand U10523 (N_10523,N_319,N_4165);
and U10524 (N_10524,N_3162,N_4743);
xnor U10525 (N_10525,N_2832,N_1486);
or U10526 (N_10526,N_1101,N_3028);
nor U10527 (N_10527,N_4146,N_2099);
or U10528 (N_10528,N_3474,N_458);
nor U10529 (N_10529,N_3068,N_5661);
or U10530 (N_10530,N_615,N_3658);
and U10531 (N_10531,N_2457,N_4747);
and U10532 (N_10532,N_743,N_1820);
nor U10533 (N_10533,N_227,N_2248);
or U10534 (N_10534,N_5932,N_2165);
and U10535 (N_10535,N_4810,N_3782);
nor U10536 (N_10536,N_162,N_872);
xnor U10537 (N_10537,N_2130,N_1925);
and U10538 (N_10538,N_4344,N_5420);
nand U10539 (N_10539,N_1342,N_2005);
nor U10540 (N_10540,N_2315,N_5256);
and U10541 (N_10541,N_122,N_2257);
and U10542 (N_10542,N_1905,N_3852);
or U10543 (N_10543,N_4454,N_5332);
and U10544 (N_10544,N_760,N_2607);
nand U10545 (N_10545,N_2747,N_646);
nand U10546 (N_10546,N_2079,N_1165);
or U10547 (N_10547,N_1932,N_3508);
xor U10548 (N_10548,N_5549,N_868);
nand U10549 (N_10549,N_4687,N_2681);
nor U10550 (N_10550,N_70,N_2159);
nor U10551 (N_10551,N_2827,N_4388);
nand U10552 (N_10552,N_1216,N_2337);
or U10553 (N_10553,N_5752,N_2738);
or U10554 (N_10554,N_4986,N_6130);
xor U10555 (N_10555,N_3677,N_4304);
or U10556 (N_10556,N_4992,N_3552);
and U10557 (N_10557,N_509,N_5065);
nor U10558 (N_10558,N_4153,N_4846);
nand U10559 (N_10559,N_5447,N_560);
and U10560 (N_10560,N_50,N_377);
nand U10561 (N_10561,N_3802,N_6098);
and U10562 (N_10562,N_2565,N_4443);
and U10563 (N_10563,N_3415,N_2903);
nand U10564 (N_10564,N_1134,N_1802);
or U10565 (N_10565,N_37,N_1731);
and U10566 (N_10566,N_679,N_561);
or U10567 (N_10567,N_1582,N_2442);
and U10568 (N_10568,N_2418,N_79);
or U10569 (N_10569,N_2805,N_1989);
xnor U10570 (N_10570,N_2517,N_3336);
nor U10571 (N_10571,N_3886,N_2040);
xor U10572 (N_10572,N_5628,N_965);
nand U10573 (N_10573,N_2493,N_1892);
or U10574 (N_10574,N_5748,N_4443);
or U10575 (N_10575,N_4616,N_5715);
nor U10576 (N_10576,N_3222,N_2105);
and U10577 (N_10577,N_100,N_623);
and U10578 (N_10578,N_4062,N_739);
or U10579 (N_10579,N_4219,N_2738);
and U10580 (N_10580,N_4212,N_6142);
nor U10581 (N_10581,N_3270,N_2252);
or U10582 (N_10582,N_1003,N_1802);
or U10583 (N_10583,N_2848,N_2510);
or U10584 (N_10584,N_5669,N_1524);
xor U10585 (N_10585,N_4629,N_5287);
or U10586 (N_10586,N_5727,N_3189);
nor U10587 (N_10587,N_3809,N_811);
xnor U10588 (N_10588,N_1773,N_1052);
and U10589 (N_10589,N_658,N_2550);
xor U10590 (N_10590,N_4377,N_3755);
or U10591 (N_10591,N_3409,N_706);
and U10592 (N_10592,N_3439,N_2744);
or U10593 (N_10593,N_3363,N_2443);
or U10594 (N_10594,N_5376,N_1634);
and U10595 (N_10595,N_1343,N_2835);
or U10596 (N_10596,N_3377,N_1668);
nand U10597 (N_10597,N_517,N_4019);
and U10598 (N_10598,N_4187,N_5420);
nand U10599 (N_10599,N_449,N_4325);
and U10600 (N_10600,N_4568,N_4670);
nor U10601 (N_10601,N_1348,N_875);
nand U10602 (N_10602,N_5119,N_2678);
nor U10603 (N_10603,N_2774,N_4317);
nor U10604 (N_10604,N_5074,N_2002);
nand U10605 (N_10605,N_850,N_4484);
or U10606 (N_10606,N_5358,N_4568);
and U10607 (N_10607,N_4030,N_607);
nor U10608 (N_10608,N_2385,N_5894);
xor U10609 (N_10609,N_1367,N_1564);
xor U10610 (N_10610,N_2222,N_1514);
or U10611 (N_10611,N_4936,N_2574);
nor U10612 (N_10612,N_6228,N_6063);
and U10613 (N_10613,N_5965,N_2258);
xnor U10614 (N_10614,N_484,N_5808);
or U10615 (N_10615,N_1301,N_4350);
nand U10616 (N_10616,N_4379,N_1256);
or U10617 (N_10617,N_1755,N_3254);
or U10618 (N_10618,N_3665,N_4613);
and U10619 (N_10619,N_4168,N_417);
xnor U10620 (N_10620,N_1462,N_2805);
nand U10621 (N_10621,N_4968,N_5704);
nand U10622 (N_10622,N_4572,N_4067);
nor U10623 (N_10623,N_362,N_2961);
or U10624 (N_10624,N_3725,N_6025);
xor U10625 (N_10625,N_5535,N_480);
and U10626 (N_10626,N_5234,N_4493);
nand U10627 (N_10627,N_885,N_3118);
and U10628 (N_10628,N_2697,N_3854);
nand U10629 (N_10629,N_5236,N_3932);
nor U10630 (N_10630,N_2243,N_4392);
nor U10631 (N_10631,N_5650,N_3516);
nor U10632 (N_10632,N_2588,N_4181);
xnor U10633 (N_10633,N_3397,N_3707);
nor U10634 (N_10634,N_3960,N_4049);
and U10635 (N_10635,N_398,N_4657);
xnor U10636 (N_10636,N_2021,N_1909);
and U10637 (N_10637,N_3970,N_1033);
nor U10638 (N_10638,N_3782,N_4383);
or U10639 (N_10639,N_2355,N_5931);
nand U10640 (N_10640,N_5357,N_5650);
nand U10641 (N_10641,N_2204,N_5258);
or U10642 (N_10642,N_5712,N_6094);
nand U10643 (N_10643,N_5430,N_5246);
xor U10644 (N_10644,N_3446,N_5592);
or U10645 (N_10645,N_6163,N_3589);
nor U10646 (N_10646,N_6001,N_2365);
xnor U10647 (N_10647,N_1896,N_52);
xor U10648 (N_10648,N_252,N_4906);
and U10649 (N_10649,N_977,N_4881);
or U10650 (N_10650,N_2063,N_720);
and U10651 (N_10651,N_1923,N_5718);
xnor U10652 (N_10652,N_4738,N_3278);
or U10653 (N_10653,N_1198,N_3057);
or U10654 (N_10654,N_1004,N_2843);
nor U10655 (N_10655,N_417,N_622);
and U10656 (N_10656,N_2752,N_1611);
and U10657 (N_10657,N_5896,N_3819);
xor U10658 (N_10658,N_2189,N_41);
nand U10659 (N_10659,N_2866,N_3433);
nand U10660 (N_10660,N_3839,N_269);
or U10661 (N_10661,N_469,N_147);
xor U10662 (N_10662,N_5894,N_0);
or U10663 (N_10663,N_3294,N_4173);
and U10664 (N_10664,N_6009,N_3531);
nor U10665 (N_10665,N_1525,N_4501);
nor U10666 (N_10666,N_1831,N_509);
and U10667 (N_10667,N_4820,N_1608);
or U10668 (N_10668,N_3605,N_3143);
nor U10669 (N_10669,N_1250,N_4952);
or U10670 (N_10670,N_3591,N_1613);
nor U10671 (N_10671,N_1419,N_288);
or U10672 (N_10672,N_3298,N_3280);
nor U10673 (N_10673,N_3006,N_3737);
nor U10674 (N_10674,N_2080,N_5662);
and U10675 (N_10675,N_2550,N_2747);
xor U10676 (N_10676,N_4708,N_2345);
or U10677 (N_10677,N_450,N_615);
nor U10678 (N_10678,N_72,N_6139);
nor U10679 (N_10679,N_6054,N_228);
and U10680 (N_10680,N_6149,N_463);
xnor U10681 (N_10681,N_2448,N_2646);
nor U10682 (N_10682,N_1305,N_4139);
or U10683 (N_10683,N_3120,N_3130);
nand U10684 (N_10684,N_5651,N_2543);
nand U10685 (N_10685,N_1924,N_1737);
and U10686 (N_10686,N_3265,N_1332);
or U10687 (N_10687,N_614,N_1852);
nor U10688 (N_10688,N_3861,N_430);
or U10689 (N_10689,N_2545,N_5360);
nand U10690 (N_10690,N_2218,N_902);
or U10691 (N_10691,N_664,N_5945);
or U10692 (N_10692,N_1905,N_72);
xnor U10693 (N_10693,N_5272,N_4072);
xnor U10694 (N_10694,N_2128,N_4752);
or U10695 (N_10695,N_1901,N_4558);
xnor U10696 (N_10696,N_1336,N_4967);
nand U10697 (N_10697,N_3552,N_4801);
and U10698 (N_10698,N_3691,N_5983);
or U10699 (N_10699,N_5438,N_1956);
nand U10700 (N_10700,N_3346,N_4340);
nor U10701 (N_10701,N_3644,N_5833);
and U10702 (N_10702,N_3855,N_2229);
or U10703 (N_10703,N_345,N_4880);
xnor U10704 (N_10704,N_368,N_4100);
or U10705 (N_10705,N_125,N_5631);
nand U10706 (N_10706,N_4556,N_2755);
xor U10707 (N_10707,N_5405,N_1316);
nor U10708 (N_10708,N_4834,N_685);
or U10709 (N_10709,N_2274,N_109);
or U10710 (N_10710,N_628,N_4287);
nand U10711 (N_10711,N_1960,N_4210);
nor U10712 (N_10712,N_6198,N_1707);
or U10713 (N_10713,N_1666,N_5370);
nor U10714 (N_10714,N_4880,N_4620);
and U10715 (N_10715,N_3473,N_235);
and U10716 (N_10716,N_141,N_712);
nor U10717 (N_10717,N_3627,N_5870);
nand U10718 (N_10718,N_145,N_6142);
nor U10719 (N_10719,N_462,N_4156);
or U10720 (N_10720,N_2197,N_4845);
or U10721 (N_10721,N_3879,N_4520);
and U10722 (N_10722,N_639,N_5926);
xor U10723 (N_10723,N_4767,N_4288);
xor U10724 (N_10724,N_3881,N_4675);
nor U10725 (N_10725,N_5517,N_2926);
nor U10726 (N_10726,N_2483,N_2087);
or U10727 (N_10727,N_1633,N_5625);
xnor U10728 (N_10728,N_1623,N_3102);
or U10729 (N_10729,N_1688,N_5784);
nor U10730 (N_10730,N_127,N_6000);
nand U10731 (N_10731,N_5393,N_1163);
or U10732 (N_10732,N_617,N_4826);
xor U10733 (N_10733,N_4964,N_1113);
xnor U10734 (N_10734,N_5533,N_2233);
and U10735 (N_10735,N_5076,N_598);
xnor U10736 (N_10736,N_2419,N_1715);
and U10737 (N_10737,N_4490,N_588);
and U10738 (N_10738,N_5968,N_5960);
nor U10739 (N_10739,N_6146,N_2597);
or U10740 (N_10740,N_3671,N_5336);
nor U10741 (N_10741,N_3889,N_463);
nand U10742 (N_10742,N_5596,N_6173);
nand U10743 (N_10743,N_3348,N_838);
or U10744 (N_10744,N_3360,N_2107);
nand U10745 (N_10745,N_4813,N_3153);
or U10746 (N_10746,N_4684,N_5633);
nand U10747 (N_10747,N_414,N_875);
xor U10748 (N_10748,N_703,N_5744);
nand U10749 (N_10749,N_3230,N_4339);
nor U10750 (N_10750,N_4473,N_4167);
or U10751 (N_10751,N_5279,N_766);
and U10752 (N_10752,N_4754,N_6220);
nor U10753 (N_10753,N_247,N_1841);
nor U10754 (N_10754,N_3503,N_1406);
or U10755 (N_10755,N_3128,N_3414);
nand U10756 (N_10756,N_2000,N_4318);
and U10757 (N_10757,N_1937,N_3041);
xnor U10758 (N_10758,N_5095,N_5847);
nor U10759 (N_10759,N_5872,N_4540);
nand U10760 (N_10760,N_2104,N_5809);
nor U10761 (N_10761,N_2744,N_2026);
xor U10762 (N_10762,N_6204,N_1752);
or U10763 (N_10763,N_1107,N_4777);
xor U10764 (N_10764,N_6148,N_700);
nand U10765 (N_10765,N_5484,N_911);
nor U10766 (N_10766,N_3384,N_5302);
nand U10767 (N_10767,N_2639,N_3217);
xor U10768 (N_10768,N_976,N_2000);
and U10769 (N_10769,N_3270,N_1183);
xnor U10770 (N_10770,N_1285,N_3343);
or U10771 (N_10771,N_6249,N_283);
nor U10772 (N_10772,N_5272,N_2601);
and U10773 (N_10773,N_4236,N_1445);
or U10774 (N_10774,N_4642,N_3909);
xor U10775 (N_10775,N_531,N_1201);
and U10776 (N_10776,N_1215,N_3172);
or U10777 (N_10777,N_4630,N_5689);
nor U10778 (N_10778,N_62,N_2981);
nor U10779 (N_10779,N_3045,N_704);
xor U10780 (N_10780,N_5623,N_4722);
nand U10781 (N_10781,N_682,N_3431);
nand U10782 (N_10782,N_364,N_321);
and U10783 (N_10783,N_3805,N_5049);
xor U10784 (N_10784,N_3919,N_134);
or U10785 (N_10785,N_6103,N_603);
or U10786 (N_10786,N_1888,N_344);
xnor U10787 (N_10787,N_4890,N_1731);
and U10788 (N_10788,N_5270,N_2316);
xnor U10789 (N_10789,N_1479,N_1453);
nand U10790 (N_10790,N_5751,N_3121);
or U10791 (N_10791,N_2158,N_1938);
nor U10792 (N_10792,N_4946,N_3902);
nand U10793 (N_10793,N_4102,N_4722);
and U10794 (N_10794,N_1483,N_82);
nor U10795 (N_10795,N_1040,N_2241);
or U10796 (N_10796,N_3967,N_2464);
and U10797 (N_10797,N_3231,N_1710);
xor U10798 (N_10798,N_466,N_5071);
and U10799 (N_10799,N_4490,N_3120);
nand U10800 (N_10800,N_1547,N_3403);
nand U10801 (N_10801,N_2520,N_379);
nor U10802 (N_10802,N_546,N_787);
nor U10803 (N_10803,N_4147,N_3515);
nor U10804 (N_10804,N_1785,N_4904);
and U10805 (N_10805,N_1616,N_4188);
or U10806 (N_10806,N_5355,N_4122);
or U10807 (N_10807,N_3114,N_3199);
xnor U10808 (N_10808,N_5346,N_3955);
nand U10809 (N_10809,N_5140,N_1033);
xor U10810 (N_10810,N_4471,N_2951);
and U10811 (N_10811,N_574,N_5322);
nand U10812 (N_10812,N_577,N_748);
or U10813 (N_10813,N_2332,N_4848);
nand U10814 (N_10814,N_1228,N_18);
nand U10815 (N_10815,N_2396,N_3468);
or U10816 (N_10816,N_4363,N_3242);
nand U10817 (N_10817,N_1977,N_1415);
nand U10818 (N_10818,N_3084,N_1644);
and U10819 (N_10819,N_3215,N_2801);
nand U10820 (N_10820,N_5551,N_4934);
or U10821 (N_10821,N_4807,N_4412);
nand U10822 (N_10822,N_2609,N_5748);
xor U10823 (N_10823,N_2626,N_2265);
and U10824 (N_10824,N_993,N_5047);
nand U10825 (N_10825,N_3064,N_5337);
xor U10826 (N_10826,N_2996,N_1895);
and U10827 (N_10827,N_889,N_230);
and U10828 (N_10828,N_5145,N_4580);
nand U10829 (N_10829,N_2345,N_5454);
xnor U10830 (N_10830,N_5207,N_4951);
or U10831 (N_10831,N_4294,N_326);
or U10832 (N_10832,N_2952,N_2326);
xor U10833 (N_10833,N_1462,N_2014);
xor U10834 (N_10834,N_2625,N_6113);
nand U10835 (N_10835,N_2377,N_3416);
nand U10836 (N_10836,N_3845,N_5621);
and U10837 (N_10837,N_2562,N_5941);
nor U10838 (N_10838,N_5891,N_724);
xnor U10839 (N_10839,N_4066,N_4928);
nor U10840 (N_10840,N_3515,N_884);
nand U10841 (N_10841,N_139,N_4016);
xnor U10842 (N_10842,N_5945,N_736);
and U10843 (N_10843,N_5880,N_3926);
nand U10844 (N_10844,N_3907,N_5150);
xor U10845 (N_10845,N_847,N_3362);
nor U10846 (N_10846,N_4947,N_3002);
nor U10847 (N_10847,N_1587,N_3202);
nor U10848 (N_10848,N_3133,N_1110);
and U10849 (N_10849,N_5294,N_6242);
xor U10850 (N_10850,N_3014,N_1844);
xor U10851 (N_10851,N_322,N_3482);
and U10852 (N_10852,N_2902,N_5891);
or U10853 (N_10853,N_690,N_4982);
nand U10854 (N_10854,N_587,N_2344);
xnor U10855 (N_10855,N_5765,N_2886);
and U10856 (N_10856,N_5912,N_1943);
nor U10857 (N_10857,N_5435,N_4812);
and U10858 (N_10858,N_4398,N_1182);
and U10859 (N_10859,N_4173,N_576);
nand U10860 (N_10860,N_3630,N_4178);
nand U10861 (N_10861,N_3026,N_4673);
or U10862 (N_10862,N_3127,N_6081);
nor U10863 (N_10863,N_5987,N_603);
or U10864 (N_10864,N_5656,N_6196);
and U10865 (N_10865,N_1300,N_3658);
or U10866 (N_10866,N_1948,N_4574);
and U10867 (N_10867,N_394,N_720);
nand U10868 (N_10868,N_4885,N_6127);
nand U10869 (N_10869,N_3,N_3438);
nor U10870 (N_10870,N_3096,N_3053);
or U10871 (N_10871,N_5791,N_2065);
nor U10872 (N_10872,N_164,N_1304);
xor U10873 (N_10873,N_4372,N_3331);
and U10874 (N_10874,N_4433,N_2106);
xor U10875 (N_10875,N_1329,N_4693);
or U10876 (N_10876,N_2218,N_2387);
xor U10877 (N_10877,N_1199,N_5354);
nor U10878 (N_10878,N_1621,N_5863);
or U10879 (N_10879,N_2339,N_5859);
and U10880 (N_10880,N_1010,N_2952);
or U10881 (N_10881,N_2178,N_5461);
nand U10882 (N_10882,N_6128,N_3821);
nand U10883 (N_10883,N_3485,N_3343);
or U10884 (N_10884,N_751,N_1111);
xor U10885 (N_10885,N_1800,N_2811);
or U10886 (N_10886,N_4672,N_2027);
or U10887 (N_10887,N_4796,N_2597);
and U10888 (N_10888,N_3822,N_2505);
or U10889 (N_10889,N_1907,N_4114);
nand U10890 (N_10890,N_2871,N_3465);
or U10891 (N_10891,N_2835,N_3147);
or U10892 (N_10892,N_6035,N_3478);
nand U10893 (N_10893,N_4464,N_4868);
xnor U10894 (N_10894,N_1032,N_3104);
and U10895 (N_10895,N_2522,N_4790);
and U10896 (N_10896,N_6239,N_6161);
nand U10897 (N_10897,N_5097,N_1947);
or U10898 (N_10898,N_4472,N_3186);
and U10899 (N_10899,N_4345,N_630);
or U10900 (N_10900,N_4706,N_2958);
or U10901 (N_10901,N_4444,N_3430);
nor U10902 (N_10902,N_950,N_3474);
nand U10903 (N_10903,N_4658,N_4951);
and U10904 (N_10904,N_4009,N_5544);
and U10905 (N_10905,N_1836,N_2042);
or U10906 (N_10906,N_1946,N_1031);
nand U10907 (N_10907,N_6186,N_4683);
xor U10908 (N_10908,N_4938,N_5965);
nor U10909 (N_10909,N_4743,N_3407);
xor U10910 (N_10910,N_3188,N_5424);
xnor U10911 (N_10911,N_5024,N_270);
and U10912 (N_10912,N_3205,N_1929);
or U10913 (N_10913,N_1887,N_5901);
and U10914 (N_10914,N_5096,N_674);
nor U10915 (N_10915,N_3728,N_1803);
xnor U10916 (N_10916,N_5379,N_4034);
and U10917 (N_10917,N_5122,N_2860);
nand U10918 (N_10918,N_940,N_3531);
nor U10919 (N_10919,N_5338,N_881);
xnor U10920 (N_10920,N_3145,N_6067);
or U10921 (N_10921,N_5712,N_3639);
nand U10922 (N_10922,N_5021,N_3917);
or U10923 (N_10923,N_5280,N_3776);
or U10924 (N_10924,N_3069,N_3672);
and U10925 (N_10925,N_1184,N_1651);
xor U10926 (N_10926,N_537,N_3078);
or U10927 (N_10927,N_337,N_988);
xor U10928 (N_10928,N_1905,N_1848);
xor U10929 (N_10929,N_1076,N_4347);
xnor U10930 (N_10930,N_562,N_576);
xnor U10931 (N_10931,N_3472,N_5011);
xor U10932 (N_10932,N_2781,N_5978);
and U10933 (N_10933,N_16,N_4333);
xor U10934 (N_10934,N_2545,N_4931);
nor U10935 (N_10935,N_1919,N_767);
xnor U10936 (N_10936,N_290,N_5842);
xor U10937 (N_10937,N_2892,N_4839);
or U10938 (N_10938,N_3427,N_2844);
and U10939 (N_10939,N_4543,N_722);
nor U10940 (N_10940,N_3738,N_4837);
xor U10941 (N_10941,N_5995,N_5303);
and U10942 (N_10942,N_3788,N_5742);
xor U10943 (N_10943,N_3711,N_167);
nand U10944 (N_10944,N_1550,N_4405);
xor U10945 (N_10945,N_687,N_2725);
nor U10946 (N_10946,N_6006,N_4857);
nand U10947 (N_10947,N_721,N_1594);
nand U10948 (N_10948,N_604,N_290);
or U10949 (N_10949,N_2492,N_6064);
nand U10950 (N_10950,N_1273,N_3120);
or U10951 (N_10951,N_3481,N_3645);
nor U10952 (N_10952,N_5585,N_6019);
and U10953 (N_10953,N_6083,N_2216);
nand U10954 (N_10954,N_631,N_5934);
nor U10955 (N_10955,N_1612,N_852);
or U10956 (N_10956,N_1448,N_3660);
xnor U10957 (N_10957,N_5098,N_5688);
nand U10958 (N_10958,N_5828,N_608);
nand U10959 (N_10959,N_1956,N_2755);
or U10960 (N_10960,N_264,N_6118);
and U10961 (N_10961,N_3386,N_5510);
or U10962 (N_10962,N_1269,N_2446);
nand U10963 (N_10963,N_5880,N_4089);
xnor U10964 (N_10964,N_1311,N_5471);
nor U10965 (N_10965,N_4300,N_1046);
nand U10966 (N_10966,N_5115,N_2843);
and U10967 (N_10967,N_4825,N_5495);
xnor U10968 (N_10968,N_2622,N_4858);
and U10969 (N_10969,N_1404,N_3054);
or U10970 (N_10970,N_5227,N_322);
xnor U10971 (N_10971,N_2409,N_3291);
nand U10972 (N_10972,N_1823,N_1846);
nand U10973 (N_10973,N_4727,N_3315);
nand U10974 (N_10974,N_2413,N_1695);
xor U10975 (N_10975,N_1201,N_5666);
and U10976 (N_10976,N_3347,N_201);
nand U10977 (N_10977,N_742,N_106);
or U10978 (N_10978,N_5105,N_4497);
nor U10979 (N_10979,N_1367,N_4549);
nor U10980 (N_10980,N_4040,N_3827);
and U10981 (N_10981,N_1750,N_5161);
nand U10982 (N_10982,N_199,N_4615);
and U10983 (N_10983,N_5619,N_5881);
or U10984 (N_10984,N_697,N_4867);
or U10985 (N_10985,N_5301,N_2029);
nor U10986 (N_10986,N_3597,N_4250);
nor U10987 (N_10987,N_699,N_96);
nor U10988 (N_10988,N_4987,N_2100);
nor U10989 (N_10989,N_4941,N_2604);
xnor U10990 (N_10990,N_5535,N_1743);
and U10991 (N_10991,N_2005,N_5934);
xnor U10992 (N_10992,N_5958,N_1065);
xnor U10993 (N_10993,N_1822,N_906);
xnor U10994 (N_10994,N_643,N_3655);
nor U10995 (N_10995,N_3756,N_5515);
nand U10996 (N_10996,N_4500,N_5956);
nand U10997 (N_10997,N_3517,N_223);
or U10998 (N_10998,N_3305,N_6015);
and U10999 (N_10999,N_1206,N_4439);
xor U11000 (N_11000,N_4939,N_815);
nor U11001 (N_11001,N_1281,N_957);
or U11002 (N_11002,N_5810,N_3542);
and U11003 (N_11003,N_5249,N_1535);
nand U11004 (N_11004,N_2555,N_4494);
nand U11005 (N_11005,N_3362,N_5608);
and U11006 (N_11006,N_1549,N_5825);
and U11007 (N_11007,N_6005,N_5383);
or U11008 (N_11008,N_4304,N_1051);
and U11009 (N_11009,N_4695,N_1397);
or U11010 (N_11010,N_2748,N_5696);
nand U11011 (N_11011,N_6225,N_5160);
xor U11012 (N_11012,N_2146,N_1801);
nand U11013 (N_11013,N_96,N_2931);
xnor U11014 (N_11014,N_3997,N_4701);
or U11015 (N_11015,N_1959,N_4308);
or U11016 (N_11016,N_3135,N_5099);
and U11017 (N_11017,N_5713,N_2441);
nor U11018 (N_11018,N_3004,N_1294);
or U11019 (N_11019,N_1474,N_719);
and U11020 (N_11020,N_1415,N_1490);
nor U11021 (N_11021,N_4764,N_1893);
and U11022 (N_11022,N_719,N_4955);
xnor U11023 (N_11023,N_4299,N_352);
and U11024 (N_11024,N_576,N_3600);
nor U11025 (N_11025,N_5950,N_2022);
or U11026 (N_11026,N_5582,N_2963);
and U11027 (N_11027,N_5060,N_2890);
xor U11028 (N_11028,N_232,N_5267);
or U11029 (N_11029,N_4386,N_3813);
or U11030 (N_11030,N_1297,N_5396);
xor U11031 (N_11031,N_4245,N_5776);
nor U11032 (N_11032,N_1793,N_829);
xor U11033 (N_11033,N_473,N_121);
nor U11034 (N_11034,N_3902,N_1983);
nand U11035 (N_11035,N_328,N_2099);
nor U11036 (N_11036,N_5643,N_5255);
and U11037 (N_11037,N_4638,N_5958);
xnor U11038 (N_11038,N_1022,N_1894);
nor U11039 (N_11039,N_3415,N_1402);
nand U11040 (N_11040,N_5,N_5624);
nor U11041 (N_11041,N_3043,N_4940);
and U11042 (N_11042,N_3570,N_1716);
nor U11043 (N_11043,N_1331,N_2187);
xor U11044 (N_11044,N_2668,N_5093);
nor U11045 (N_11045,N_1924,N_4058);
nand U11046 (N_11046,N_5092,N_223);
nand U11047 (N_11047,N_1622,N_2110);
nand U11048 (N_11048,N_277,N_3422);
and U11049 (N_11049,N_2522,N_1269);
or U11050 (N_11050,N_4475,N_1626);
and U11051 (N_11051,N_2328,N_4916);
xor U11052 (N_11052,N_2121,N_125);
and U11053 (N_11053,N_5528,N_1740);
nor U11054 (N_11054,N_3461,N_4702);
or U11055 (N_11055,N_4170,N_2431);
nand U11056 (N_11056,N_5569,N_2770);
or U11057 (N_11057,N_5903,N_163);
or U11058 (N_11058,N_6084,N_6219);
and U11059 (N_11059,N_3368,N_1254);
xnor U11060 (N_11060,N_1381,N_2267);
xor U11061 (N_11061,N_486,N_3856);
nor U11062 (N_11062,N_380,N_2566);
xor U11063 (N_11063,N_2176,N_1403);
and U11064 (N_11064,N_2765,N_2340);
and U11065 (N_11065,N_2989,N_6087);
or U11066 (N_11066,N_5372,N_5014);
nand U11067 (N_11067,N_2560,N_1242);
nand U11068 (N_11068,N_782,N_3007);
nor U11069 (N_11069,N_4778,N_5500);
nor U11070 (N_11070,N_5248,N_2306);
and U11071 (N_11071,N_2587,N_3315);
xor U11072 (N_11072,N_6025,N_3237);
nor U11073 (N_11073,N_1505,N_3805);
or U11074 (N_11074,N_4123,N_5229);
or U11075 (N_11075,N_411,N_5017);
and U11076 (N_11076,N_817,N_3454);
nor U11077 (N_11077,N_2285,N_73);
nand U11078 (N_11078,N_5374,N_5532);
nand U11079 (N_11079,N_1241,N_961);
and U11080 (N_11080,N_5280,N_1045);
nand U11081 (N_11081,N_3375,N_2145);
xnor U11082 (N_11082,N_3940,N_5182);
nand U11083 (N_11083,N_3496,N_5924);
nor U11084 (N_11084,N_4372,N_5957);
nor U11085 (N_11085,N_5880,N_2748);
nor U11086 (N_11086,N_1370,N_4944);
xnor U11087 (N_11087,N_3445,N_3715);
or U11088 (N_11088,N_1107,N_1249);
xor U11089 (N_11089,N_5057,N_295);
and U11090 (N_11090,N_3196,N_3627);
nand U11091 (N_11091,N_4360,N_467);
or U11092 (N_11092,N_209,N_6162);
nand U11093 (N_11093,N_3341,N_3267);
nor U11094 (N_11094,N_4682,N_5525);
and U11095 (N_11095,N_940,N_5959);
or U11096 (N_11096,N_4351,N_706);
or U11097 (N_11097,N_4995,N_2528);
xnor U11098 (N_11098,N_687,N_1492);
xnor U11099 (N_11099,N_1577,N_4769);
nand U11100 (N_11100,N_131,N_3558);
or U11101 (N_11101,N_4710,N_5607);
xnor U11102 (N_11102,N_260,N_2289);
xor U11103 (N_11103,N_5969,N_3645);
and U11104 (N_11104,N_3350,N_2183);
nand U11105 (N_11105,N_1173,N_5861);
or U11106 (N_11106,N_2431,N_1503);
nor U11107 (N_11107,N_3902,N_2131);
nor U11108 (N_11108,N_146,N_1231);
xnor U11109 (N_11109,N_3256,N_5287);
or U11110 (N_11110,N_4648,N_4125);
xor U11111 (N_11111,N_6184,N_1296);
nand U11112 (N_11112,N_2786,N_3682);
nand U11113 (N_11113,N_260,N_3687);
or U11114 (N_11114,N_3494,N_5818);
nand U11115 (N_11115,N_717,N_1994);
or U11116 (N_11116,N_656,N_1566);
and U11117 (N_11117,N_797,N_6142);
or U11118 (N_11118,N_6020,N_1710);
or U11119 (N_11119,N_2213,N_2795);
and U11120 (N_11120,N_5953,N_4132);
nand U11121 (N_11121,N_2419,N_3866);
xor U11122 (N_11122,N_855,N_5513);
and U11123 (N_11123,N_6109,N_4340);
xor U11124 (N_11124,N_4028,N_1764);
xnor U11125 (N_11125,N_3250,N_4110);
xnor U11126 (N_11126,N_4076,N_4231);
nand U11127 (N_11127,N_4506,N_2774);
nand U11128 (N_11128,N_6030,N_5671);
or U11129 (N_11129,N_984,N_3247);
and U11130 (N_11130,N_408,N_4580);
xnor U11131 (N_11131,N_515,N_385);
nand U11132 (N_11132,N_4,N_3837);
or U11133 (N_11133,N_708,N_2973);
nor U11134 (N_11134,N_4437,N_5375);
nor U11135 (N_11135,N_4292,N_4571);
or U11136 (N_11136,N_5699,N_762);
nor U11137 (N_11137,N_1458,N_486);
nor U11138 (N_11138,N_3151,N_4581);
and U11139 (N_11139,N_4554,N_3019);
or U11140 (N_11140,N_4891,N_3199);
xnor U11141 (N_11141,N_4319,N_1174);
xnor U11142 (N_11142,N_5241,N_1358);
nand U11143 (N_11143,N_3681,N_3877);
nor U11144 (N_11144,N_2604,N_5769);
nand U11145 (N_11145,N_4125,N_3079);
or U11146 (N_11146,N_5041,N_3249);
or U11147 (N_11147,N_250,N_3696);
xnor U11148 (N_11148,N_1186,N_3373);
or U11149 (N_11149,N_5380,N_546);
and U11150 (N_11150,N_1184,N_4851);
nor U11151 (N_11151,N_5432,N_3178);
or U11152 (N_11152,N_2099,N_6017);
nand U11153 (N_11153,N_3892,N_1095);
nand U11154 (N_11154,N_3801,N_2270);
nand U11155 (N_11155,N_298,N_974);
nand U11156 (N_11156,N_3014,N_2655);
and U11157 (N_11157,N_1624,N_5433);
nor U11158 (N_11158,N_6064,N_6045);
xnor U11159 (N_11159,N_1413,N_2259);
and U11160 (N_11160,N_4109,N_595);
nor U11161 (N_11161,N_1145,N_1717);
nand U11162 (N_11162,N_3720,N_3144);
xor U11163 (N_11163,N_5603,N_2446);
or U11164 (N_11164,N_2646,N_1015);
or U11165 (N_11165,N_5480,N_6006);
nand U11166 (N_11166,N_4672,N_6153);
and U11167 (N_11167,N_456,N_1430);
nor U11168 (N_11168,N_2707,N_1770);
nand U11169 (N_11169,N_1591,N_892);
and U11170 (N_11170,N_2727,N_1948);
nand U11171 (N_11171,N_5291,N_4752);
or U11172 (N_11172,N_2920,N_829);
or U11173 (N_11173,N_4597,N_1715);
nand U11174 (N_11174,N_5866,N_950);
or U11175 (N_11175,N_4982,N_3449);
nand U11176 (N_11176,N_1663,N_2122);
nand U11177 (N_11177,N_625,N_1191);
nor U11178 (N_11178,N_4593,N_5864);
xor U11179 (N_11179,N_5303,N_5667);
and U11180 (N_11180,N_2525,N_6050);
and U11181 (N_11181,N_3029,N_1852);
or U11182 (N_11182,N_4786,N_80);
nor U11183 (N_11183,N_5834,N_3497);
nor U11184 (N_11184,N_2409,N_811);
nand U11185 (N_11185,N_1873,N_3800);
xor U11186 (N_11186,N_3163,N_144);
or U11187 (N_11187,N_5345,N_1453);
xor U11188 (N_11188,N_2300,N_4023);
xnor U11189 (N_11189,N_402,N_2928);
nand U11190 (N_11190,N_3676,N_1853);
nor U11191 (N_11191,N_661,N_473);
and U11192 (N_11192,N_4195,N_1834);
and U11193 (N_11193,N_1314,N_6043);
and U11194 (N_11194,N_1397,N_5333);
or U11195 (N_11195,N_668,N_534);
or U11196 (N_11196,N_1843,N_537);
and U11197 (N_11197,N_4581,N_3232);
or U11198 (N_11198,N_5798,N_236);
or U11199 (N_11199,N_4216,N_4245);
nand U11200 (N_11200,N_3943,N_2250);
xor U11201 (N_11201,N_4618,N_1580);
nand U11202 (N_11202,N_1229,N_2054);
xor U11203 (N_11203,N_5967,N_1367);
nand U11204 (N_11204,N_5293,N_346);
and U11205 (N_11205,N_1737,N_2758);
nand U11206 (N_11206,N_4032,N_6223);
and U11207 (N_11207,N_4563,N_962);
nand U11208 (N_11208,N_1437,N_609);
or U11209 (N_11209,N_6042,N_4286);
or U11210 (N_11210,N_4075,N_5154);
xnor U11211 (N_11211,N_523,N_6100);
or U11212 (N_11212,N_431,N_4880);
nor U11213 (N_11213,N_808,N_5166);
xor U11214 (N_11214,N_3414,N_3584);
or U11215 (N_11215,N_2537,N_5346);
xnor U11216 (N_11216,N_4940,N_4887);
or U11217 (N_11217,N_3046,N_431);
nand U11218 (N_11218,N_4493,N_5382);
and U11219 (N_11219,N_1721,N_5491);
xnor U11220 (N_11220,N_877,N_77);
and U11221 (N_11221,N_2655,N_1894);
nor U11222 (N_11222,N_867,N_1829);
xor U11223 (N_11223,N_3853,N_4436);
xor U11224 (N_11224,N_5691,N_2660);
nand U11225 (N_11225,N_4683,N_2838);
or U11226 (N_11226,N_2990,N_2837);
or U11227 (N_11227,N_178,N_1545);
and U11228 (N_11228,N_1458,N_3310);
xnor U11229 (N_11229,N_3893,N_4915);
and U11230 (N_11230,N_1101,N_363);
or U11231 (N_11231,N_6048,N_1014);
xnor U11232 (N_11232,N_3574,N_2336);
nor U11233 (N_11233,N_5637,N_274);
xnor U11234 (N_11234,N_5012,N_3539);
and U11235 (N_11235,N_6173,N_5120);
xor U11236 (N_11236,N_1182,N_6165);
nor U11237 (N_11237,N_5970,N_3846);
xnor U11238 (N_11238,N_3002,N_2615);
nor U11239 (N_11239,N_4668,N_2480);
or U11240 (N_11240,N_5243,N_3671);
and U11241 (N_11241,N_2395,N_5277);
or U11242 (N_11242,N_5381,N_2694);
nor U11243 (N_11243,N_2968,N_630);
nand U11244 (N_11244,N_1095,N_5352);
nand U11245 (N_11245,N_3253,N_1244);
and U11246 (N_11246,N_2764,N_287);
and U11247 (N_11247,N_1831,N_4521);
nand U11248 (N_11248,N_6012,N_3051);
nand U11249 (N_11249,N_6107,N_4307);
or U11250 (N_11250,N_1367,N_3110);
nor U11251 (N_11251,N_2850,N_3412);
nand U11252 (N_11252,N_3427,N_4096);
and U11253 (N_11253,N_3312,N_5639);
or U11254 (N_11254,N_1114,N_5833);
and U11255 (N_11255,N_2634,N_3240);
and U11256 (N_11256,N_5491,N_833);
or U11257 (N_11257,N_1540,N_2590);
nor U11258 (N_11258,N_2592,N_1584);
nand U11259 (N_11259,N_4451,N_643);
nand U11260 (N_11260,N_5623,N_2584);
xor U11261 (N_11261,N_1672,N_996);
and U11262 (N_11262,N_4521,N_5021);
xor U11263 (N_11263,N_2425,N_3954);
nand U11264 (N_11264,N_863,N_879);
xnor U11265 (N_11265,N_2149,N_802);
and U11266 (N_11266,N_326,N_5212);
and U11267 (N_11267,N_4009,N_1198);
and U11268 (N_11268,N_95,N_6022);
nand U11269 (N_11269,N_1816,N_3837);
nor U11270 (N_11270,N_1757,N_323);
or U11271 (N_11271,N_2557,N_1547);
or U11272 (N_11272,N_3957,N_5719);
or U11273 (N_11273,N_1136,N_1066);
or U11274 (N_11274,N_6096,N_2577);
nor U11275 (N_11275,N_2512,N_107);
and U11276 (N_11276,N_1775,N_595);
xnor U11277 (N_11277,N_4881,N_1757);
and U11278 (N_11278,N_951,N_1583);
xor U11279 (N_11279,N_3911,N_2983);
xnor U11280 (N_11280,N_4611,N_667);
xor U11281 (N_11281,N_5136,N_1595);
xor U11282 (N_11282,N_6016,N_4034);
or U11283 (N_11283,N_270,N_5158);
or U11284 (N_11284,N_1733,N_2002);
xnor U11285 (N_11285,N_5432,N_518);
nor U11286 (N_11286,N_3999,N_4652);
nand U11287 (N_11287,N_5095,N_5019);
and U11288 (N_11288,N_1363,N_4259);
and U11289 (N_11289,N_2462,N_845);
or U11290 (N_11290,N_5645,N_3587);
xor U11291 (N_11291,N_4321,N_4798);
and U11292 (N_11292,N_102,N_3634);
nor U11293 (N_11293,N_1776,N_591);
xnor U11294 (N_11294,N_365,N_130);
nor U11295 (N_11295,N_5194,N_3809);
nand U11296 (N_11296,N_3201,N_5109);
nor U11297 (N_11297,N_1656,N_355);
xnor U11298 (N_11298,N_3746,N_4441);
nor U11299 (N_11299,N_175,N_2644);
and U11300 (N_11300,N_2900,N_690);
nand U11301 (N_11301,N_1959,N_856);
nor U11302 (N_11302,N_5827,N_2513);
and U11303 (N_11303,N_5702,N_0);
and U11304 (N_11304,N_3008,N_2607);
nand U11305 (N_11305,N_4745,N_1307);
nor U11306 (N_11306,N_1350,N_2809);
nand U11307 (N_11307,N_1060,N_3842);
or U11308 (N_11308,N_798,N_2139);
or U11309 (N_11309,N_4722,N_5740);
nor U11310 (N_11310,N_4273,N_4104);
nor U11311 (N_11311,N_369,N_5090);
xor U11312 (N_11312,N_971,N_3468);
nand U11313 (N_11313,N_2377,N_4126);
and U11314 (N_11314,N_1710,N_1341);
xor U11315 (N_11315,N_4258,N_3851);
nor U11316 (N_11316,N_1041,N_5425);
xnor U11317 (N_11317,N_4256,N_3855);
or U11318 (N_11318,N_373,N_890);
and U11319 (N_11319,N_3091,N_382);
nand U11320 (N_11320,N_4225,N_772);
and U11321 (N_11321,N_2110,N_2216);
nand U11322 (N_11322,N_2782,N_1347);
nor U11323 (N_11323,N_749,N_179);
and U11324 (N_11324,N_759,N_2693);
and U11325 (N_11325,N_949,N_557);
and U11326 (N_11326,N_1536,N_1650);
nand U11327 (N_11327,N_5948,N_549);
xor U11328 (N_11328,N_2185,N_4972);
and U11329 (N_11329,N_1532,N_5208);
nand U11330 (N_11330,N_6041,N_3651);
nand U11331 (N_11331,N_2476,N_5932);
nor U11332 (N_11332,N_828,N_4559);
nor U11333 (N_11333,N_493,N_4366);
and U11334 (N_11334,N_4742,N_6176);
nand U11335 (N_11335,N_2741,N_5191);
nor U11336 (N_11336,N_3132,N_3803);
and U11337 (N_11337,N_3074,N_4842);
nand U11338 (N_11338,N_2609,N_4616);
nor U11339 (N_11339,N_3219,N_2346);
and U11340 (N_11340,N_4941,N_3495);
and U11341 (N_11341,N_3216,N_421);
or U11342 (N_11342,N_1284,N_5710);
nor U11343 (N_11343,N_2994,N_2648);
or U11344 (N_11344,N_3345,N_2933);
nand U11345 (N_11345,N_2810,N_2111);
nor U11346 (N_11346,N_1219,N_2584);
nor U11347 (N_11347,N_3469,N_4866);
nor U11348 (N_11348,N_1526,N_5012);
or U11349 (N_11349,N_1300,N_3722);
nor U11350 (N_11350,N_5563,N_1205);
and U11351 (N_11351,N_4114,N_3565);
xnor U11352 (N_11352,N_3228,N_5833);
or U11353 (N_11353,N_36,N_5569);
and U11354 (N_11354,N_3670,N_3244);
or U11355 (N_11355,N_1862,N_4186);
and U11356 (N_11356,N_1682,N_4765);
nand U11357 (N_11357,N_2954,N_2165);
nor U11358 (N_11358,N_2,N_4345);
and U11359 (N_11359,N_5242,N_5439);
xor U11360 (N_11360,N_2141,N_4507);
nor U11361 (N_11361,N_6007,N_632);
and U11362 (N_11362,N_1572,N_554);
or U11363 (N_11363,N_3730,N_1383);
xor U11364 (N_11364,N_1068,N_6217);
xnor U11365 (N_11365,N_1188,N_772);
nand U11366 (N_11366,N_3306,N_1785);
nor U11367 (N_11367,N_296,N_3674);
xnor U11368 (N_11368,N_219,N_4093);
nand U11369 (N_11369,N_4626,N_452);
nor U11370 (N_11370,N_5879,N_4752);
or U11371 (N_11371,N_3228,N_3215);
xnor U11372 (N_11372,N_4095,N_139);
nor U11373 (N_11373,N_2177,N_1523);
nor U11374 (N_11374,N_3227,N_5307);
xor U11375 (N_11375,N_5036,N_5368);
nand U11376 (N_11376,N_2109,N_1937);
nor U11377 (N_11377,N_2556,N_1833);
and U11378 (N_11378,N_2399,N_6127);
xor U11379 (N_11379,N_1440,N_3594);
nand U11380 (N_11380,N_4256,N_5006);
xor U11381 (N_11381,N_612,N_4412);
nand U11382 (N_11382,N_1331,N_4471);
or U11383 (N_11383,N_2910,N_1125);
xnor U11384 (N_11384,N_3519,N_477);
or U11385 (N_11385,N_1354,N_4616);
xor U11386 (N_11386,N_4606,N_3017);
nor U11387 (N_11387,N_589,N_5756);
and U11388 (N_11388,N_5610,N_2730);
nor U11389 (N_11389,N_6182,N_5091);
and U11390 (N_11390,N_3207,N_884);
xor U11391 (N_11391,N_5760,N_3542);
xnor U11392 (N_11392,N_5973,N_690);
or U11393 (N_11393,N_5988,N_4749);
or U11394 (N_11394,N_2433,N_3701);
or U11395 (N_11395,N_2814,N_5853);
nand U11396 (N_11396,N_4889,N_140);
xnor U11397 (N_11397,N_2592,N_810);
xnor U11398 (N_11398,N_5464,N_1362);
and U11399 (N_11399,N_2939,N_5712);
and U11400 (N_11400,N_5819,N_5026);
and U11401 (N_11401,N_3344,N_2631);
or U11402 (N_11402,N_1948,N_6227);
and U11403 (N_11403,N_876,N_172);
and U11404 (N_11404,N_5067,N_1329);
xor U11405 (N_11405,N_5533,N_3574);
nand U11406 (N_11406,N_305,N_3540);
or U11407 (N_11407,N_5845,N_1019);
nand U11408 (N_11408,N_3067,N_4057);
and U11409 (N_11409,N_3202,N_464);
nand U11410 (N_11410,N_1121,N_2868);
nor U11411 (N_11411,N_5402,N_2085);
xor U11412 (N_11412,N_4300,N_4169);
and U11413 (N_11413,N_5006,N_1149);
or U11414 (N_11414,N_6004,N_6168);
xnor U11415 (N_11415,N_3225,N_4646);
nor U11416 (N_11416,N_6017,N_4539);
and U11417 (N_11417,N_4492,N_5150);
nand U11418 (N_11418,N_1717,N_2010);
nor U11419 (N_11419,N_5375,N_5408);
nand U11420 (N_11420,N_1839,N_1274);
or U11421 (N_11421,N_5328,N_5726);
or U11422 (N_11422,N_498,N_1432);
nand U11423 (N_11423,N_3180,N_5924);
and U11424 (N_11424,N_3705,N_4551);
or U11425 (N_11425,N_1316,N_1966);
and U11426 (N_11426,N_4644,N_1824);
or U11427 (N_11427,N_5250,N_1779);
and U11428 (N_11428,N_1957,N_191);
or U11429 (N_11429,N_1563,N_5606);
nand U11430 (N_11430,N_3356,N_4570);
xor U11431 (N_11431,N_3759,N_2282);
xnor U11432 (N_11432,N_5691,N_6191);
nor U11433 (N_11433,N_2942,N_4273);
or U11434 (N_11434,N_3423,N_189);
xor U11435 (N_11435,N_3547,N_2201);
and U11436 (N_11436,N_1996,N_1312);
nand U11437 (N_11437,N_3332,N_4468);
xor U11438 (N_11438,N_5873,N_3766);
or U11439 (N_11439,N_2245,N_490);
nand U11440 (N_11440,N_334,N_3813);
and U11441 (N_11441,N_3066,N_662);
xnor U11442 (N_11442,N_101,N_2264);
nor U11443 (N_11443,N_3388,N_696);
and U11444 (N_11444,N_4156,N_3761);
nand U11445 (N_11445,N_79,N_5579);
nand U11446 (N_11446,N_806,N_3683);
nor U11447 (N_11447,N_1128,N_4023);
nor U11448 (N_11448,N_1113,N_5360);
nand U11449 (N_11449,N_33,N_2927);
and U11450 (N_11450,N_1489,N_3026);
xor U11451 (N_11451,N_2327,N_2782);
nand U11452 (N_11452,N_5809,N_467);
xnor U11453 (N_11453,N_2313,N_4696);
nor U11454 (N_11454,N_5746,N_1286);
xnor U11455 (N_11455,N_3644,N_3226);
nand U11456 (N_11456,N_1335,N_2593);
xnor U11457 (N_11457,N_5045,N_5356);
and U11458 (N_11458,N_4336,N_5976);
nor U11459 (N_11459,N_1746,N_654);
or U11460 (N_11460,N_446,N_3285);
nor U11461 (N_11461,N_2102,N_5233);
and U11462 (N_11462,N_1157,N_1128);
nand U11463 (N_11463,N_6025,N_2425);
nor U11464 (N_11464,N_657,N_6131);
nand U11465 (N_11465,N_773,N_4256);
xor U11466 (N_11466,N_5223,N_1986);
nand U11467 (N_11467,N_811,N_4822);
and U11468 (N_11468,N_5023,N_96);
and U11469 (N_11469,N_891,N_3222);
and U11470 (N_11470,N_3824,N_117);
nand U11471 (N_11471,N_2076,N_43);
xor U11472 (N_11472,N_2611,N_758);
or U11473 (N_11473,N_4317,N_266);
nor U11474 (N_11474,N_368,N_5071);
xnor U11475 (N_11475,N_3060,N_4872);
nor U11476 (N_11476,N_2903,N_1862);
nand U11477 (N_11477,N_6063,N_3115);
or U11478 (N_11478,N_2651,N_6223);
nor U11479 (N_11479,N_5843,N_2280);
and U11480 (N_11480,N_3013,N_1616);
and U11481 (N_11481,N_370,N_4355);
nand U11482 (N_11482,N_4664,N_1603);
or U11483 (N_11483,N_5954,N_2887);
xnor U11484 (N_11484,N_2763,N_4601);
and U11485 (N_11485,N_3646,N_4298);
nor U11486 (N_11486,N_4770,N_2811);
nand U11487 (N_11487,N_3181,N_4248);
xnor U11488 (N_11488,N_1004,N_1620);
or U11489 (N_11489,N_5846,N_1141);
nand U11490 (N_11490,N_647,N_4970);
and U11491 (N_11491,N_742,N_2083);
xnor U11492 (N_11492,N_884,N_1395);
nand U11493 (N_11493,N_3870,N_361);
xnor U11494 (N_11494,N_3717,N_1948);
xor U11495 (N_11495,N_782,N_4835);
nor U11496 (N_11496,N_3094,N_3406);
nand U11497 (N_11497,N_3036,N_2002);
or U11498 (N_11498,N_216,N_4187);
xnor U11499 (N_11499,N_3845,N_6076);
and U11500 (N_11500,N_1141,N_248);
and U11501 (N_11501,N_2488,N_4641);
xor U11502 (N_11502,N_2424,N_4403);
xnor U11503 (N_11503,N_1349,N_5035);
nand U11504 (N_11504,N_810,N_175);
and U11505 (N_11505,N_3141,N_4421);
xnor U11506 (N_11506,N_2563,N_76);
xnor U11507 (N_11507,N_1558,N_4816);
nand U11508 (N_11508,N_3685,N_3863);
and U11509 (N_11509,N_3519,N_2354);
or U11510 (N_11510,N_4462,N_627);
nand U11511 (N_11511,N_1321,N_6177);
and U11512 (N_11512,N_710,N_5930);
or U11513 (N_11513,N_4589,N_3765);
xor U11514 (N_11514,N_5871,N_3449);
and U11515 (N_11515,N_506,N_1639);
or U11516 (N_11516,N_3025,N_5598);
nand U11517 (N_11517,N_5760,N_4669);
nand U11518 (N_11518,N_5573,N_1013);
xnor U11519 (N_11519,N_5907,N_3447);
or U11520 (N_11520,N_298,N_6006);
and U11521 (N_11521,N_1824,N_719);
nor U11522 (N_11522,N_4568,N_3156);
and U11523 (N_11523,N_1111,N_5895);
xor U11524 (N_11524,N_4182,N_4776);
xor U11525 (N_11525,N_1833,N_2311);
xor U11526 (N_11526,N_5199,N_2299);
xnor U11527 (N_11527,N_5866,N_564);
xnor U11528 (N_11528,N_1659,N_4128);
nor U11529 (N_11529,N_279,N_2029);
nor U11530 (N_11530,N_2079,N_635);
xor U11531 (N_11531,N_4277,N_4971);
xor U11532 (N_11532,N_4085,N_1429);
xor U11533 (N_11533,N_4357,N_4660);
or U11534 (N_11534,N_2038,N_1286);
and U11535 (N_11535,N_1099,N_2996);
xor U11536 (N_11536,N_2859,N_2450);
or U11537 (N_11537,N_6013,N_1550);
nand U11538 (N_11538,N_3549,N_1602);
or U11539 (N_11539,N_2895,N_5959);
or U11540 (N_11540,N_648,N_4033);
nand U11541 (N_11541,N_1368,N_3752);
nand U11542 (N_11542,N_3904,N_120);
nor U11543 (N_11543,N_3462,N_2127);
nor U11544 (N_11544,N_1497,N_4596);
xnor U11545 (N_11545,N_1240,N_5385);
xnor U11546 (N_11546,N_4837,N_933);
nor U11547 (N_11547,N_2674,N_232);
nand U11548 (N_11548,N_3879,N_2089);
and U11549 (N_11549,N_383,N_1417);
or U11550 (N_11550,N_2797,N_983);
or U11551 (N_11551,N_2007,N_2361);
nand U11552 (N_11552,N_4320,N_2930);
nor U11553 (N_11553,N_1386,N_5770);
xor U11554 (N_11554,N_5594,N_3897);
xor U11555 (N_11555,N_2803,N_5771);
nor U11556 (N_11556,N_2658,N_1853);
nand U11557 (N_11557,N_4380,N_4157);
or U11558 (N_11558,N_1602,N_415);
nor U11559 (N_11559,N_2065,N_1407);
xnor U11560 (N_11560,N_5371,N_230);
and U11561 (N_11561,N_528,N_4664);
and U11562 (N_11562,N_1119,N_2698);
or U11563 (N_11563,N_3389,N_4677);
nand U11564 (N_11564,N_1373,N_6157);
or U11565 (N_11565,N_873,N_4377);
xor U11566 (N_11566,N_4948,N_1260);
nor U11567 (N_11567,N_1937,N_2850);
and U11568 (N_11568,N_3208,N_5977);
xnor U11569 (N_11569,N_3019,N_44);
nor U11570 (N_11570,N_1473,N_5943);
and U11571 (N_11571,N_2489,N_3486);
nor U11572 (N_11572,N_4035,N_5831);
nor U11573 (N_11573,N_4186,N_3939);
or U11574 (N_11574,N_4467,N_2128);
xor U11575 (N_11575,N_5451,N_2337);
nand U11576 (N_11576,N_5886,N_4813);
or U11577 (N_11577,N_793,N_1690);
nand U11578 (N_11578,N_3083,N_2999);
xnor U11579 (N_11579,N_835,N_5793);
xnor U11580 (N_11580,N_5924,N_2648);
or U11581 (N_11581,N_4856,N_4000);
and U11582 (N_11582,N_5110,N_3427);
xor U11583 (N_11583,N_89,N_491);
nand U11584 (N_11584,N_972,N_4378);
and U11585 (N_11585,N_2277,N_3396);
nand U11586 (N_11586,N_3607,N_4721);
and U11587 (N_11587,N_4766,N_1834);
and U11588 (N_11588,N_6157,N_2438);
and U11589 (N_11589,N_2173,N_3768);
nor U11590 (N_11590,N_1750,N_3222);
and U11591 (N_11591,N_1223,N_3246);
and U11592 (N_11592,N_4649,N_4150);
and U11593 (N_11593,N_4863,N_4007);
or U11594 (N_11594,N_3499,N_1853);
and U11595 (N_11595,N_4850,N_6030);
and U11596 (N_11596,N_3136,N_2052);
nor U11597 (N_11597,N_852,N_6111);
nor U11598 (N_11598,N_5128,N_3339);
and U11599 (N_11599,N_4339,N_5992);
nor U11600 (N_11600,N_384,N_449);
xnor U11601 (N_11601,N_2345,N_3801);
or U11602 (N_11602,N_6095,N_4632);
xor U11603 (N_11603,N_3866,N_3209);
or U11604 (N_11604,N_5530,N_4037);
or U11605 (N_11605,N_1123,N_744);
and U11606 (N_11606,N_5676,N_4436);
nand U11607 (N_11607,N_609,N_3799);
or U11608 (N_11608,N_2098,N_1011);
xor U11609 (N_11609,N_1037,N_1668);
or U11610 (N_11610,N_3108,N_2977);
and U11611 (N_11611,N_3077,N_3353);
or U11612 (N_11612,N_2158,N_1243);
and U11613 (N_11613,N_922,N_6161);
xnor U11614 (N_11614,N_3332,N_4449);
and U11615 (N_11615,N_1743,N_4775);
nand U11616 (N_11616,N_4076,N_2054);
nor U11617 (N_11617,N_755,N_5264);
and U11618 (N_11618,N_4963,N_5553);
or U11619 (N_11619,N_238,N_3075);
or U11620 (N_11620,N_5488,N_1869);
nand U11621 (N_11621,N_134,N_3060);
nor U11622 (N_11622,N_4255,N_5957);
nor U11623 (N_11623,N_4047,N_2801);
and U11624 (N_11624,N_1642,N_2462);
and U11625 (N_11625,N_2502,N_2027);
xor U11626 (N_11626,N_1877,N_1523);
nor U11627 (N_11627,N_740,N_18);
nand U11628 (N_11628,N_3895,N_4452);
xor U11629 (N_11629,N_3368,N_1030);
nand U11630 (N_11630,N_4526,N_905);
nand U11631 (N_11631,N_4544,N_541);
xor U11632 (N_11632,N_2293,N_1416);
nand U11633 (N_11633,N_1534,N_4667);
or U11634 (N_11634,N_2800,N_2325);
nor U11635 (N_11635,N_5738,N_5770);
or U11636 (N_11636,N_3661,N_433);
nor U11637 (N_11637,N_4326,N_2569);
nor U11638 (N_11638,N_3774,N_856);
nor U11639 (N_11639,N_3777,N_2748);
xor U11640 (N_11640,N_1988,N_3061);
and U11641 (N_11641,N_5862,N_2712);
or U11642 (N_11642,N_2272,N_5783);
xnor U11643 (N_11643,N_5354,N_5379);
nand U11644 (N_11644,N_2965,N_5073);
nand U11645 (N_11645,N_4605,N_2896);
nand U11646 (N_11646,N_4652,N_4843);
and U11647 (N_11647,N_1617,N_3248);
and U11648 (N_11648,N_2495,N_1368);
or U11649 (N_11649,N_966,N_1388);
xor U11650 (N_11650,N_4113,N_2304);
or U11651 (N_11651,N_5163,N_2918);
and U11652 (N_11652,N_3211,N_5134);
xor U11653 (N_11653,N_1696,N_4605);
xor U11654 (N_11654,N_4416,N_509);
xnor U11655 (N_11655,N_4738,N_5387);
xor U11656 (N_11656,N_3315,N_4844);
nor U11657 (N_11657,N_787,N_2976);
or U11658 (N_11658,N_3115,N_5585);
xnor U11659 (N_11659,N_3716,N_4212);
nand U11660 (N_11660,N_1427,N_671);
nand U11661 (N_11661,N_4532,N_5624);
nor U11662 (N_11662,N_4955,N_2695);
nand U11663 (N_11663,N_2068,N_5002);
nand U11664 (N_11664,N_65,N_1255);
and U11665 (N_11665,N_2720,N_4946);
or U11666 (N_11666,N_5076,N_1892);
nand U11667 (N_11667,N_5550,N_2642);
xnor U11668 (N_11668,N_535,N_2814);
and U11669 (N_11669,N_3212,N_1835);
and U11670 (N_11670,N_843,N_3448);
or U11671 (N_11671,N_778,N_5548);
or U11672 (N_11672,N_1105,N_6036);
xor U11673 (N_11673,N_4754,N_3390);
nand U11674 (N_11674,N_5513,N_578);
or U11675 (N_11675,N_1455,N_2876);
and U11676 (N_11676,N_3263,N_2978);
nor U11677 (N_11677,N_4680,N_5907);
or U11678 (N_11678,N_5582,N_3072);
xor U11679 (N_11679,N_2200,N_3042);
nor U11680 (N_11680,N_1149,N_5752);
xnor U11681 (N_11681,N_5598,N_6015);
and U11682 (N_11682,N_5650,N_3092);
or U11683 (N_11683,N_4482,N_2360);
nor U11684 (N_11684,N_1534,N_2490);
nor U11685 (N_11685,N_3975,N_3755);
and U11686 (N_11686,N_6243,N_1501);
and U11687 (N_11687,N_2767,N_6238);
xor U11688 (N_11688,N_5296,N_4610);
xnor U11689 (N_11689,N_4823,N_4425);
and U11690 (N_11690,N_6143,N_4696);
xnor U11691 (N_11691,N_376,N_762);
and U11692 (N_11692,N_4093,N_66);
nand U11693 (N_11693,N_994,N_405);
nand U11694 (N_11694,N_3248,N_735);
and U11695 (N_11695,N_5763,N_3588);
nor U11696 (N_11696,N_1099,N_1275);
xor U11697 (N_11697,N_1880,N_1670);
nor U11698 (N_11698,N_1016,N_3864);
nor U11699 (N_11699,N_2890,N_2023);
or U11700 (N_11700,N_1001,N_3543);
and U11701 (N_11701,N_5773,N_5128);
nor U11702 (N_11702,N_2704,N_3898);
xor U11703 (N_11703,N_154,N_4961);
nand U11704 (N_11704,N_1551,N_46);
or U11705 (N_11705,N_3058,N_4503);
nor U11706 (N_11706,N_2974,N_2581);
nand U11707 (N_11707,N_512,N_962);
and U11708 (N_11708,N_2913,N_2609);
xnor U11709 (N_11709,N_4953,N_5372);
nor U11710 (N_11710,N_4623,N_5707);
nand U11711 (N_11711,N_2664,N_4058);
nor U11712 (N_11712,N_4499,N_5817);
or U11713 (N_11713,N_1882,N_5793);
xor U11714 (N_11714,N_4008,N_3271);
or U11715 (N_11715,N_717,N_2226);
and U11716 (N_11716,N_1006,N_2284);
and U11717 (N_11717,N_5380,N_3036);
nor U11718 (N_11718,N_3948,N_4558);
and U11719 (N_11719,N_4257,N_4116);
nor U11720 (N_11720,N_4232,N_5100);
nor U11721 (N_11721,N_2646,N_3102);
nor U11722 (N_11722,N_4908,N_3436);
or U11723 (N_11723,N_944,N_3757);
and U11724 (N_11724,N_4212,N_680);
nand U11725 (N_11725,N_5992,N_3099);
xnor U11726 (N_11726,N_4007,N_5370);
or U11727 (N_11727,N_3972,N_1582);
nor U11728 (N_11728,N_1349,N_1219);
xor U11729 (N_11729,N_2378,N_1247);
nand U11730 (N_11730,N_5761,N_2070);
or U11731 (N_11731,N_2127,N_5761);
or U11732 (N_11732,N_437,N_1407);
xnor U11733 (N_11733,N_1598,N_119);
and U11734 (N_11734,N_3933,N_942);
xor U11735 (N_11735,N_2969,N_636);
or U11736 (N_11736,N_5820,N_4645);
nor U11737 (N_11737,N_5950,N_6177);
nor U11738 (N_11738,N_4791,N_4131);
or U11739 (N_11739,N_3187,N_1017);
and U11740 (N_11740,N_3776,N_5570);
xor U11741 (N_11741,N_475,N_3908);
nand U11742 (N_11742,N_4420,N_31);
and U11743 (N_11743,N_4749,N_1325);
nor U11744 (N_11744,N_2566,N_2977);
xor U11745 (N_11745,N_3871,N_3900);
nor U11746 (N_11746,N_3861,N_5612);
nor U11747 (N_11747,N_1929,N_5971);
and U11748 (N_11748,N_4875,N_1076);
nand U11749 (N_11749,N_5326,N_218);
and U11750 (N_11750,N_3847,N_1198);
nand U11751 (N_11751,N_2897,N_5296);
and U11752 (N_11752,N_4529,N_5214);
and U11753 (N_11753,N_3563,N_4469);
xnor U11754 (N_11754,N_4048,N_5363);
xor U11755 (N_11755,N_3887,N_1102);
nor U11756 (N_11756,N_1846,N_4046);
nand U11757 (N_11757,N_4854,N_2800);
nand U11758 (N_11758,N_365,N_261);
and U11759 (N_11759,N_1633,N_2421);
or U11760 (N_11760,N_2841,N_3034);
nand U11761 (N_11761,N_2490,N_2118);
or U11762 (N_11762,N_5605,N_60);
and U11763 (N_11763,N_5358,N_5101);
nor U11764 (N_11764,N_1654,N_630);
xor U11765 (N_11765,N_5478,N_5817);
nand U11766 (N_11766,N_3125,N_3773);
xor U11767 (N_11767,N_2142,N_3409);
or U11768 (N_11768,N_1353,N_3563);
or U11769 (N_11769,N_3879,N_4076);
nand U11770 (N_11770,N_2668,N_5639);
or U11771 (N_11771,N_1956,N_3657);
nor U11772 (N_11772,N_2744,N_1765);
xor U11773 (N_11773,N_1271,N_3021);
nand U11774 (N_11774,N_5299,N_2896);
xnor U11775 (N_11775,N_2542,N_839);
or U11776 (N_11776,N_3716,N_4307);
and U11777 (N_11777,N_2163,N_4010);
xor U11778 (N_11778,N_1577,N_5641);
and U11779 (N_11779,N_2158,N_3166);
and U11780 (N_11780,N_2274,N_2242);
nor U11781 (N_11781,N_1140,N_3477);
and U11782 (N_11782,N_2462,N_320);
xor U11783 (N_11783,N_3603,N_3199);
nor U11784 (N_11784,N_44,N_4431);
and U11785 (N_11785,N_2569,N_4472);
xnor U11786 (N_11786,N_943,N_2399);
and U11787 (N_11787,N_5117,N_183);
xor U11788 (N_11788,N_1491,N_3805);
or U11789 (N_11789,N_4013,N_4620);
or U11790 (N_11790,N_4185,N_3617);
nor U11791 (N_11791,N_5534,N_5223);
nand U11792 (N_11792,N_5736,N_554);
xnor U11793 (N_11793,N_520,N_2604);
and U11794 (N_11794,N_580,N_1206);
or U11795 (N_11795,N_3059,N_5130);
xor U11796 (N_11796,N_2360,N_4040);
nand U11797 (N_11797,N_677,N_2496);
nor U11798 (N_11798,N_1144,N_4763);
xnor U11799 (N_11799,N_3249,N_552);
and U11800 (N_11800,N_3689,N_5204);
nand U11801 (N_11801,N_5578,N_2829);
nand U11802 (N_11802,N_4712,N_3832);
or U11803 (N_11803,N_3550,N_2218);
and U11804 (N_11804,N_4143,N_3083);
and U11805 (N_11805,N_292,N_609);
or U11806 (N_11806,N_1139,N_3040);
nand U11807 (N_11807,N_5177,N_1163);
and U11808 (N_11808,N_5381,N_5363);
nor U11809 (N_11809,N_5998,N_4960);
nand U11810 (N_11810,N_5672,N_2532);
xor U11811 (N_11811,N_1720,N_1592);
and U11812 (N_11812,N_3732,N_3885);
and U11813 (N_11813,N_124,N_1845);
nand U11814 (N_11814,N_5386,N_135);
xnor U11815 (N_11815,N_1003,N_221);
nor U11816 (N_11816,N_2146,N_6146);
nor U11817 (N_11817,N_5286,N_4355);
or U11818 (N_11818,N_2666,N_3638);
and U11819 (N_11819,N_3060,N_891);
nand U11820 (N_11820,N_3746,N_2032);
or U11821 (N_11821,N_3831,N_5616);
or U11822 (N_11822,N_1510,N_4701);
xor U11823 (N_11823,N_2596,N_2331);
xnor U11824 (N_11824,N_2715,N_4020);
and U11825 (N_11825,N_4632,N_1833);
or U11826 (N_11826,N_4199,N_5478);
and U11827 (N_11827,N_5562,N_1519);
or U11828 (N_11828,N_1382,N_2023);
and U11829 (N_11829,N_1042,N_3560);
or U11830 (N_11830,N_3431,N_5270);
nand U11831 (N_11831,N_5673,N_3270);
nand U11832 (N_11832,N_6088,N_2587);
xor U11833 (N_11833,N_743,N_5707);
nand U11834 (N_11834,N_4321,N_631);
and U11835 (N_11835,N_42,N_3247);
or U11836 (N_11836,N_349,N_4524);
or U11837 (N_11837,N_4165,N_2379);
and U11838 (N_11838,N_1652,N_203);
xnor U11839 (N_11839,N_837,N_1562);
xor U11840 (N_11840,N_3963,N_2004);
nor U11841 (N_11841,N_6165,N_5437);
or U11842 (N_11842,N_3271,N_3663);
nor U11843 (N_11843,N_5353,N_348);
nand U11844 (N_11844,N_3599,N_3793);
nand U11845 (N_11845,N_3116,N_683);
nor U11846 (N_11846,N_2878,N_5207);
nor U11847 (N_11847,N_4245,N_5219);
and U11848 (N_11848,N_3508,N_2790);
or U11849 (N_11849,N_5769,N_5095);
nand U11850 (N_11850,N_5561,N_1528);
xnor U11851 (N_11851,N_2347,N_2179);
xnor U11852 (N_11852,N_275,N_6045);
or U11853 (N_11853,N_5505,N_2335);
nand U11854 (N_11854,N_5082,N_413);
nand U11855 (N_11855,N_5608,N_6135);
and U11856 (N_11856,N_6171,N_1862);
or U11857 (N_11857,N_4192,N_1067);
and U11858 (N_11858,N_4202,N_4482);
xnor U11859 (N_11859,N_1321,N_5042);
or U11860 (N_11860,N_2017,N_4602);
nand U11861 (N_11861,N_2165,N_171);
xor U11862 (N_11862,N_93,N_2885);
and U11863 (N_11863,N_1892,N_557);
nand U11864 (N_11864,N_6191,N_5989);
xnor U11865 (N_11865,N_3142,N_2774);
nor U11866 (N_11866,N_4499,N_2832);
nand U11867 (N_11867,N_2027,N_643);
or U11868 (N_11868,N_1692,N_4747);
nor U11869 (N_11869,N_870,N_3286);
xnor U11870 (N_11870,N_489,N_6132);
nand U11871 (N_11871,N_3907,N_5032);
and U11872 (N_11872,N_5579,N_6097);
nand U11873 (N_11873,N_3164,N_1828);
nand U11874 (N_11874,N_574,N_1191);
xor U11875 (N_11875,N_1144,N_1427);
and U11876 (N_11876,N_612,N_4670);
nor U11877 (N_11877,N_365,N_911);
xor U11878 (N_11878,N_3424,N_358);
nor U11879 (N_11879,N_1449,N_1015);
nor U11880 (N_11880,N_1864,N_3623);
and U11881 (N_11881,N_1738,N_305);
xor U11882 (N_11882,N_3805,N_5093);
and U11883 (N_11883,N_2966,N_997);
xnor U11884 (N_11884,N_3920,N_1227);
nand U11885 (N_11885,N_3803,N_1210);
or U11886 (N_11886,N_701,N_4100);
nor U11887 (N_11887,N_4935,N_1048);
or U11888 (N_11888,N_2217,N_2284);
or U11889 (N_11889,N_5230,N_5066);
and U11890 (N_11890,N_3514,N_1628);
and U11891 (N_11891,N_6146,N_573);
or U11892 (N_11892,N_4903,N_2358);
nor U11893 (N_11893,N_6052,N_3800);
and U11894 (N_11894,N_1537,N_1193);
or U11895 (N_11895,N_2228,N_5095);
or U11896 (N_11896,N_2333,N_5996);
and U11897 (N_11897,N_2871,N_320);
xor U11898 (N_11898,N_2165,N_3743);
nand U11899 (N_11899,N_5610,N_1958);
xnor U11900 (N_11900,N_5817,N_1105);
xor U11901 (N_11901,N_101,N_6139);
or U11902 (N_11902,N_4919,N_5770);
or U11903 (N_11903,N_6165,N_1547);
or U11904 (N_11904,N_2365,N_6028);
or U11905 (N_11905,N_3641,N_799);
or U11906 (N_11906,N_4314,N_4655);
and U11907 (N_11907,N_5443,N_4031);
nor U11908 (N_11908,N_6182,N_5892);
nor U11909 (N_11909,N_3231,N_686);
and U11910 (N_11910,N_604,N_133);
nor U11911 (N_11911,N_4676,N_3869);
and U11912 (N_11912,N_1501,N_682);
or U11913 (N_11913,N_250,N_1640);
and U11914 (N_11914,N_6120,N_316);
nand U11915 (N_11915,N_2096,N_4499);
nor U11916 (N_11916,N_1868,N_429);
nand U11917 (N_11917,N_1037,N_3554);
or U11918 (N_11918,N_2193,N_1325);
and U11919 (N_11919,N_5388,N_2046);
nand U11920 (N_11920,N_6106,N_1172);
nand U11921 (N_11921,N_1447,N_3807);
nand U11922 (N_11922,N_4046,N_607);
and U11923 (N_11923,N_5685,N_1684);
nor U11924 (N_11924,N_3323,N_3913);
or U11925 (N_11925,N_5724,N_4892);
xor U11926 (N_11926,N_715,N_1456);
nor U11927 (N_11927,N_2099,N_5115);
and U11928 (N_11928,N_5645,N_3099);
and U11929 (N_11929,N_5397,N_4222);
nor U11930 (N_11930,N_1790,N_3197);
nand U11931 (N_11931,N_1896,N_3688);
or U11932 (N_11932,N_5869,N_3134);
xnor U11933 (N_11933,N_5777,N_5020);
and U11934 (N_11934,N_1245,N_5748);
nand U11935 (N_11935,N_1250,N_4342);
nor U11936 (N_11936,N_3295,N_1013);
nor U11937 (N_11937,N_1111,N_4456);
and U11938 (N_11938,N_3105,N_2941);
xor U11939 (N_11939,N_574,N_4626);
nand U11940 (N_11940,N_137,N_5620);
and U11941 (N_11941,N_3436,N_190);
nor U11942 (N_11942,N_886,N_3257);
and U11943 (N_11943,N_4563,N_1074);
nor U11944 (N_11944,N_5009,N_4390);
and U11945 (N_11945,N_59,N_5757);
and U11946 (N_11946,N_958,N_4390);
nor U11947 (N_11947,N_1228,N_3702);
or U11948 (N_11948,N_2824,N_5939);
or U11949 (N_11949,N_2212,N_94);
xnor U11950 (N_11950,N_1875,N_2742);
or U11951 (N_11951,N_750,N_6231);
xor U11952 (N_11952,N_939,N_5922);
xnor U11953 (N_11953,N_3289,N_1465);
or U11954 (N_11954,N_4364,N_4396);
or U11955 (N_11955,N_5603,N_3605);
or U11956 (N_11956,N_2602,N_5643);
nor U11957 (N_11957,N_4592,N_3047);
nand U11958 (N_11958,N_5940,N_324);
xnor U11959 (N_11959,N_895,N_5346);
nor U11960 (N_11960,N_2407,N_6215);
nand U11961 (N_11961,N_393,N_2219);
nand U11962 (N_11962,N_1115,N_2948);
nor U11963 (N_11963,N_662,N_3607);
or U11964 (N_11964,N_2989,N_3416);
xor U11965 (N_11965,N_1612,N_5597);
or U11966 (N_11966,N_395,N_900);
nor U11967 (N_11967,N_3569,N_4325);
or U11968 (N_11968,N_1176,N_1855);
xnor U11969 (N_11969,N_497,N_110);
nand U11970 (N_11970,N_2105,N_6059);
nor U11971 (N_11971,N_917,N_5478);
nor U11972 (N_11972,N_3727,N_3198);
nor U11973 (N_11973,N_43,N_80);
xnor U11974 (N_11974,N_5203,N_6245);
nor U11975 (N_11975,N_1104,N_5247);
nor U11976 (N_11976,N_2322,N_2000);
and U11977 (N_11977,N_484,N_2747);
or U11978 (N_11978,N_88,N_2786);
and U11979 (N_11979,N_5117,N_4608);
xnor U11980 (N_11980,N_5766,N_203);
xnor U11981 (N_11981,N_1658,N_362);
or U11982 (N_11982,N_6101,N_2741);
and U11983 (N_11983,N_6003,N_3413);
xor U11984 (N_11984,N_3140,N_3831);
xor U11985 (N_11985,N_753,N_4248);
xnor U11986 (N_11986,N_2841,N_6107);
nand U11987 (N_11987,N_3121,N_1878);
xnor U11988 (N_11988,N_4139,N_2559);
nand U11989 (N_11989,N_2665,N_5159);
nor U11990 (N_11990,N_4696,N_27);
nor U11991 (N_11991,N_4145,N_6012);
or U11992 (N_11992,N_191,N_3812);
nand U11993 (N_11993,N_4774,N_4781);
or U11994 (N_11994,N_1509,N_5336);
and U11995 (N_11995,N_2607,N_3273);
nand U11996 (N_11996,N_2473,N_464);
nand U11997 (N_11997,N_5337,N_1658);
and U11998 (N_11998,N_4968,N_4053);
xnor U11999 (N_11999,N_752,N_5939);
and U12000 (N_12000,N_5551,N_3888);
xor U12001 (N_12001,N_929,N_1916);
xnor U12002 (N_12002,N_5445,N_4358);
and U12003 (N_12003,N_620,N_4926);
or U12004 (N_12004,N_2557,N_1277);
nand U12005 (N_12005,N_1068,N_2369);
or U12006 (N_12006,N_2014,N_4581);
nor U12007 (N_12007,N_3966,N_3544);
or U12008 (N_12008,N_385,N_1929);
and U12009 (N_12009,N_3470,N_6066);
nor U12010 (N_12010,N_1213,N_2070);
nor U12011 (N_12011,N_4980,N_4371);
and U12012 (N_12012,N_3323,N_6203);
nand U12013 (N_12013,N_4795,N_3522);
and U12014 (N_12014,N_1216,N_2333);
and U12015 (N_12015,N_5433,N_3326);
nor U12016 (N_12016,N_5989,N_3556);
or U12017 (N_12017,N_2496,N_5269);
or U12018 (N_12018,N_591,N_3439);
or U12019 (N_12019,N_5495,N_5699);
nor U12020 (N_12020,N_4245,N_2041);
or U12021 (N_12021,N_5981,N_963);
or U12022 (N_12022,N_3367,N_1953);
xor U12023 (N_12023,N_1516,N_1200);
and U12024 (N_12024,N_839,N_2295);
or U12025 (N_12025,N_5177,N_4361);
nand U12026 (N_12026,N_3943,N_5092);
nor U12027 (N_12027,N_1014,N_3325);
or U12028 (N_12028,N_679,N_5521);
and U12029 (N_12029,N_1521,N_3733);
and U12030 (N_12030,N_4933,N_5734);
xor U12031 (N_12031,N_439,N_3445);
and U12032 (N_12032,N_4606,N_2426);
nand U12033 (N_12033,N_3799,N_3315);
xor U12034 (N_12034,N_1176,N_2130);
nand U12035 (N_12035,N_5697,N_1809);
nand U12036 (N_12036,N_5521,N_1082);
and U12037 (N_12037,N_5874,N_6001);
or U12038 (N_12038,N_2500,N_2929);
nor U12039 (N_12039,N_1241,N_2945);
nand U12040 (N_12040,N_231,N_6021);
nor U12041 (N_12041,N_216,N_2044);
and U12042 (N_12042,N_2615,N_3214);
nand U12043 (N_12043,N_619,N_4948);
nand U12044 (N_12044,N_1851,N_3660);
nand U12045 (N_12045,N_3609,N_1941);
xnor U12046 (N_12046,N_5381,N_2309);
xor U12047 (N_12047,N_2325,N_5193);
and U12048 (N_12048,N_4775,N_2860);
nor U12049 (N_12049,N_3628,N_5239);
nor U12050 (N_12050,N_4165,N_4302);
nor U12051 (N_12051,N_3276,N_1920);
nor U12052 (N_12052,N_2754,N_1433);
nor U12053 (N_12053,N_504,N_1409);
xor U12054 (N_12054,N_5131,N_2703);
or U12055 (N_12055,N_2472,N_1438);
and U12056 (N_12056,N_2531,N_2680);
or U12057 (N_12057,N_5686,N_475);
xnor U12058 (N_12058,N_1802,N_2590);
or U12059 (N_12059,N_6017,N_5074);
nor U12060 (N_12060,N_4262,N_43);
xor U12061 (N_12061,N_3084,N_4312);
and U12062 (N_12062,N_5002,N_6181);
nor U12063 (N_12063,N_4485,N_5749);
xnor U12064 (N_12064,N_972,N_3271);
or U12065 (N_12065,N_446,N_6);
nor U12066 (N_12066,N_3092,N_3095);
and U12067 (N_12067,N_2556,N_5124);
and U12068 (N_12068,N_5881,N_5446);
or U12069 (N_12069,N_3963,N_4331);
and U12070 (N_12070,N_717,N_4649);
xor U12071 (N_12071,N_354,N_1430);
or U12072 (N_12072,N_5882,N_2702);
nor U12073 (N_12073,N_2028,N_2844);
or U12074 (N_12074,N_2778,N_6062);
or U12075 (N_12075,N_1948,N_3134);
and U12076 (N_12076,N_1072,N_5861);
nand U12077 (N_12077,N_4592,N_5951);
xnor U12078 (N_12078,N_1730,N_1742);
xnor U12079 (N_12079,N_2966,N_4595);
xor U12080 (N_12080,N_2465,N_539);
xnor U12081 (N_12081,N_6082,N_697);
xor U12082 (N_12082,N_5632,N_508);
and U12083 (N_12083,N_4062,N_1980);
or U12084 (N_12084,N_2229,N_1860);
nor U12085 (N_12085,N_881,N_284);
xor U12086 (N_12086,N_2740,N_5377);
or U12087 (N_12087,N_1011,N_797);
nand U12088 (N_12088,N_2425,N_1972);
or U12089 (N_12089,N_3922,N_2193);
nor U12090 (N_12090,N_85,N_1114);
or U12091 (N_12091,N_6139,N_2942);
or U12092 (N_12092,N_6178,N_2380);
or U12093 (N_12093,N_2044,N_1599);
nor U12094 (N_12094,N_5834,N_6136);
or U12095 (N_12095,N_3102,N_5861);
nand U12096 (N_12096,N_6222,N_2604);
and U12097 (N_12097,N_5326,N_5645);
xnor U12098 (N_12098,N_4699,N_4697);
nor U12099 (N_12099,N_4551,N_2522);
nor U12100 (N_12100,N_3227,N_2923);
or U12101 (N_12101,N_4136,N_2460);
nor U12102 (N_12102,N_4287,N_2743);
nand U12103 (N_12103,N_4618,N_635);
xor U12104 (N_12104,N_3128,N_4540);
nand U12105 (N_12105,N_6068,N_634);
nor U12106 (N_12106,N_5773,N_5591);
nor U12107 (N_12107,N_3624,N_2297);
or U12108 (N_12108,N_100,N_2796);
nor U12109 (N_12109,N_3426,N_5849);
nor U12110 (N_12110,N_4115,N_61);
or U12111 (N_12111,N_2662,N_3194);
or U12112 (N_12112,N_563,N_5608);
nor U12113 (N_12113,N_760,N_2781);
or U12114 (N_12114,N_2249,N_2277);
xor U12115 (N_12115,N_5206,N_5941);
and U12116 (N_12116,N_42,N_78);
nor U12117 (N_12117,N_5084,N_1906);
and U12118 (N_12118,N_2868,N_5484);
xnor U12119 (N_12119,N_1115,N_4938);
and U12120 (N_12120,N_6008,N_949);
nor U12121 (N_12121,N_2895,N_5622);
xor U12122 (N_12122,N_25,N_3482);
or U12123 (N_12123,N_1747,N_5072);
and U12124 (N_12124,N_670,N_2490);
or U12125 (N_12125,N_3306,N_1620);
and U12126 (N_12126,N_4161,N_4721);
xnor U12127 (N_12127,N_5410,N_2957);
xnor U12128 (N_12128,N_5996,N_2078);
or U12129 (N_12129,N_4470,N_755);
xnor U12130 (N_12130,N_555,N_4308);
nor U12131 (N_12131,N_2172,N_2851);
xnor U12132 (N_12132,N_449,N_5083);
nor U12133 (N_12133,N_2588,N_4429);
nand U12134 (N_12134,N_901,N_145);
nor U12135 (N_12135,N_3431,N_5331);
nor U12136 (N_12136,N_4148,N_2956);
or U12137 (N_12137,N_3931,N_4394);
and U12138 (N_12138,N_1945,N_3414);
nor U12139 (N_12139,N_1450,N_1671);
xnor U12140 (N_12140,N_3336,N_5514);
xor U12141 (N_12141,N_2771,N_3592);
and U12142 (N_12142,N_3929,N_2701);
and U12143 (N_12143,N_3097,N_5463);
nor U12144 (N_12144,N_4871,N_5691);
and U12145 (N_12145,N_5078,N_3636);
xnor U12146 (N_12146,N_2948,N_895);
nand U12147 (N_12147,N_4804,N_1962);
or U12148 (N_12148,N_3791,N_6155);
or U12149 (N_12149,N_4724,N_4026);
nand U12150 (N_12150,N_3162,N_6206);
or U12151 (N_12151,N_3693,N_2554);
and U12152 (N_12152,N_5012,N_2950);
or U12153 (N_12153,N_5221,N_2984);
nand U12154 (N_12154,N_1576,N_917);
and U12155 (N_12155,N_1797,N_2369);
nand U12156 (N_12156,N_5440,N_834);
and U12157 (N_12157,N_2549,N_248);
and U12158 (N_12158,N_2182,N_5558);
or U12159 (N_12159,N_4209,N_4180);
or U12160 (N_12160,N_2305,N_4177);
nor U12161 (N_12161,N_5769,N_3616);
nor U12162 (N_12162,N_2796,N_3854);
and U12163 (N_12163,N_2877,N_150);
xnor U12164 (N_12164,N_1215,N_5046);
nor U12165 (N_12165,N_6073,N_1440);
nand U12166 (N_12166,N_692,N_647);
and U12167 (N_12167,N_5471,N_3686);
xnor U12168 (N_12168,N_4589,N_1459);
xnor U12169 (N_12169,N_4265,N_816);
and U12170 (N_12170,N_4112,N_1085);
nand U12171 (N_12171,N_5331,N_5803);
and U12172 (N_12172,N_25,N_5093);
nor U12173 (N_12173,N_5869,N_1812);
nand U12174 (N_12174,N_5885,N_10);
xnor U12175 (N_12175,N_658,N_639);
nor U12176 (N_12176,N_1626,N_1501);
nand U12177 (N_12177,N_958,N_1922);
nand U12178 (N_12178,N_3283,N_1712);
or U12179 (N_12179,N_215,N_3717);
nand U12180 (N_12180,N_6044,N_4252);
xnor U12181 (N_12181,N_1876,N_415);
and U12182 (N_12182,N_4600,N_3985);
xor U12183 (N_12183,N_5758,N_4254);
nand U12184 (N_12184,N_1136,N_669);
and U12185 (N_12185,N_5494,N_3293);
or U12186 (N_12186,N_2116,N_6090);
nand U12187 (N_12187,N_5282,N_5067);
or U12188 (N_12188,N_4234,N_4575);
xor U12189 (N_12189,N_5320,N_2685);
xnor U12190 (N_12190,N_586,N_2695);
nand U12191 (N_12191,N_4817,N_3311);
xor U12192 (N_12192,N_3666,N_1851);
and U12193 (N_12193,N_2574,N_3276);
and U12194 (N_12194,N_222,N_4634);
or U12195 (N_12195,N_5108,N_5433);
nand U12196 (N_12196,N_1565,N_4809);
or U12197 (N_12197,N_4341,N_4201);
nor U12198 (N_12198,N_1570,N_595);
xnor U12199 (N_12199,N_1736,N_4707);
nor U12200 (N_12200,N_4591,N_4762);
nor U12201 (N_12201,N_384,N_108);
nand U12202 (N_12202,N_4503,N_435);
or U12203 (N_12203,N_261,N_5816);
or U12204 (N_12204,N_5881,N_3861);
nor U12205 (N_12205,N_6198,N_1868);
xor U12206 (N_12206,N_4879,N_4990);
nor U12207 (N_12207,N_1839,N_1569);
or U12208 (N_12208,N_3785,N_1951);
nor U12209 (N_12209,N_585,N_3246);
nor U12210 (N_12210,N_3274,N_4876);
xor U12211 (N_12211,N_335,N_4661);
and U12212 (N_12212,N_5473,N_3831);
nor U12213 (N_12213,N_5957,N_1217);
or U12214 (N_12214,N_1903,N_4008);
xor U12215 (N_12215,N_3607,N_2385);
xor U12216 (N_12216,N_1511,N_5778);
or U12217 (N_12217,N_5179,N_2174);
or U12218 (N_12218,N_3660,N_1216);
nor U12219 (N_12219,N_5425,N_2549);
nand U12220 (N_12220,N_105,N_5432);
xor U12221 (N_12221,N_6102,N_432);
nand U12222 (N_12222,N_4603,N_2964);
and U12223 (N_12223,N_1137,N_6226);
nand U12224 (N_12224,N_1787,N_79);
nor U12225 (N_12225,N_2345,N_1013);
nor U12226 (N_12226,N_2246,N_5462);
or U12227 (N_12227,N_613,N_807);
nand U12228 (N_12228,N_1835,N_1178);
xnor U12229 (N_12229,N_2595,N_687);
nand U12230 (N_12230,N_3905,N_2437);
xor U12231 (N_12231,N_54,N_5167);
nand U12232 (N_12232,N_3285,N_1227);
nor U12233 (N_12233,N_989,N_155);
nor U12234 (N_12234,N_2574,N_6059);
xnor U12235 (N_12235,N_3084,N_433);
or U12236 (N_12236,N_6048,N_4499);
and U12237 (N_12237,N_1564,N_664);
nand U12238 (N_12238,N_112,N_3765);
nand U12239 (N_12239,N_4693,N_1132);
or U12240 (N_12240,N_2667,N_787);
and U12241 (N_12241,N_1295,N_1416);
nor U12242 (N_12242,N_4939,N_5116);
xnor U12243 (N_12243,N_1162,N_4798);
nor U12244 (N_12244,N_3894,N_4670);
or U12245 (N_12245,N_261,N_4870);
xor U12246 (N_12246,N_3743,N_4353);
nand U12247 (N_12247,N_4291,N_1000);
nor U12248 (N_12248,N_1131,N_328);
or U12249 (N_12249,N_1783,N_1555);
xnor U12250 (N_12250,N_3301,N_6200);
or U12251 (N_12251,N_6218,N_1855);
nand U12252 (N_12252,N_2092,N_305);
nor U12253 (N_12253,N_4854,N_5000);
nand U12254 (N_12254,N_83,N_4991);
nor U12255 (N_12255,N_1223,N_3438);
and U12256 (N_12256,N_122,N_5357);
and U12257 (N_12257,N_4352,N_1619);
nor U12258 (N_12258,N_1822,N_1841);
and U12259 (N_12259,N_1174,N_1334);
and U12260 (N_12260,N_6092,N_197);
and U12261 (N_12261,N_4752,N_4299);
and U12262 (N_12262,N_374,N_3359);
xnor U12263 (N_12263,N_2634,N_32);
and U12264 (N_12264,N_2508,N_510);
and U12265 (N_12265,N_175,N_5078);
and U12266 (N_12266,N_2701,N_4625);
or U12267 (N_12267,N_5438,N_591);
xor U12268 (N_12268,N_2650,N_1432);
xor U12269 (N_12269,N_2603,N_2840);
xnor U12270 (N_12270,N_4247,N_2265);
xor U12271 (N_12271,N_1403,N_4002);
nand U12272 (N_12272,N_590,N_1198);
xor U12273 (N_12273,N_3564,N_200);
and U12274 (N_12274,N_1108,N_4981);
and U12275 (N_12275,N_4269,N_5967);
nand U12276 (N_12276,N_4585,N_3388);
or U12277 (N_12277,N_3283,N_2448);
or U12278 (N_12278,N_5230,N_1290);
nor U12279 (N_12279,N_4370,N_4968);
xor U12280 (N_12280,N_414,N_1735);
xor U12281 (N_12281,N_3407,N_696);
and U12282 (N_12282,N_4167,N_1014);
nor U12283 (N_12283,N_4988,N_3541);
nand U12284 (N_12284,N_2884,N_1834);
nor U12285 (N_12285,N_4985,N_1425);
xnor U12286 (N_12286,N_2608,N_4908);
nor U12287 (N_12287,N_2497,N_2511);
and U12288 (N_12288,N_110,N_3807);
nand U12289 (N_12289,N_1363,N_5086);
nand U12290 (N_12290,N_4619,N_4506);
and U12291 (N_12291,N_4938,N_5906);
nor U12292 (N_12292,N_4115,N_5481);
nor U12293 (N_12293,N_205,N_2774);
and U12294 (N_12294,N_5437,N_1744);
nand U12295 (N_12295,N_5121,N_3182);
or U12296 (N_12296,N_2784,N_5406);
xor U12297 (N_12297,N_3549,N_2506);
xnor U12298 (N_12298,N_3816,N_3839);
nand U12299 (N_12299,N_1504,N_5341);
nor U12300 (N_12300,N_1462,N_4246);
nor U12301 (N_12301,N_1052,N_1005);
nand U12302 (N_12302,N_2625,N_1981);
or U12303 (N_12303,N_5863,N_5680);
nor U12304 (N_12304,N_4542,N_2809);
nand U12305 (N_12305,N_156,N_4301);
xor U12306 (N_12306,N_4537,N_4750);
nor U12307 (N_12307,N_3911,N_5564);
nand U12308 (N_12308,N_5179,N_5195);
and U12309 (N_12309,N_3614,N_1649);
nor U12310 (N_12310,N_5323,N_4452);
and U12311 (N_12311,N_4854,N_2333);
nand U12312 (N_12312,N_2791,N_4457);
and U12313 (N_12313,N_5063,N_469);
nor U12314 (N_12314,N_1685,N_1627);
nand U12315 (N_12315,N_2830,N_4557);
nand U12316 (N_12316,N_2835,N_4530);
nor U12317 (N_12317,N_3235,N_1402);
nor U12318 (N_12318,N_4318,N_657);
xor U12319 (N_12319,N_3877,N_124);
nand U12320 (N_12320,N_3578,N_3639);
or U12321 (N_12321,N_4626,N_301);
nand U12322 (N_12322,N_5239,N_5820);
xnor U12323 (N_12323,N_2306,N_3775);
and U12324 (N_12324,N_2049,N_2883);
xor U12325 (N_12325,N_2049,N_4949);
nand U12326 (N_12326,N_5647,N_4353);
and U12327 (N_12327,N_3978,N_5269);
xnor U12328 (N_12328,N_3859,N_6218);
and U12329 (N_12329,N_5063,N_1019);
nor U12330 (N_12330,N_3730,N_480);
or U12331 (N_12331,N_3713,N_5666);
xor U12332 (N_12332,N_2446,N_5008);
nand U12333 (N_12333,N_147,N_3901);
nand U12334 (N_12334,N_1333,N_3046);
and U12335 (N_12335,N_2947,N_415);
nor U12336 (N_12336,N_5767,N_1760);
xnor U12337 (N_12337,N_2409,N_2662);
xnor U12338 (N_12338,N_2512,N_2103);
nor U12339 (N_12339,N_2984,N_5723);
xor U12340 (N_12340,N_3650,N_5923);
xnor U12341 (N_12341,N_5477,N_2253);
or U12342 (N_12342,N_1835,N_5571);
nor U12343 (N_12343,N_5931,N_1222);
xor U12344 (N_12344,N_3709,N_1978);
or U12345 (N_12345,N_2451,N_3660);
nor U12346 (N_12346,N_864,N_5821);
and U12347 (N_12347,N_796,N_5260);
or U12348 (N_12348,N_893,N_3381);
nor U12349 (N_12349,N_1138,N_5909);
nor U12350 (N_12350,N_4642,N_3949);
and U12351 (N_12351,N_1169,N_175);
nor U12352 (N_12352,N_1172,N_1079);
nand U12353 (N_12353,N_1890,N_4136);
xnor U12354 (N_12354,N_845,N_974);
or U12355 (N_12355,N_848,N_2260);
nand U12356 (N_12356,N_4421,N_5091);
and U12357 (N_12357,N_4983,N_3405);
or U12358 (N_12358,N_163,N_4078);
xnor U12359 (N_12359,N_2710,N_2085);
or U12360 (N_12360,N_4493,N_4239);
or U12361 (N_12361,N_2596,N_551);
xnor U12362 (N_12362,N_3897,N_1061);
nand U12363 (N_12363,N_5578,N_3386);
or U12364 (N_12364,N_2345,N_3147);
nor U12365 (N_12365,N_5060,N_130);
nor U12366 (N_12366,N_1421,N_1661);
or U12367 (N_12367,N_853,N_1862);
nand U12368 (N_12368,N_5416,N_3033);
nand U12369 (N_12369,N_3562,N_2333);
nor U12370 (N_12370,N_5844,N_2001);
nand U12371 (N_12371,N_414,N_3475);
nor U12372 (N_12372,N_1007,N_2981);
nor U12373 (N_12373,N_1404,N_2231);
xnor U12374 (N_12374,N_3348,N_4720);
nor U12375 (N_12375,N_5311,N_4667);
nor U12376 (N_12376,N_981,N_1208);
xnor U12377 (N_12377,N_3854,N_3303);
and U12378 (N_12378,N_3479,N_4766);
and U12379 (N_12379,N_1975,N_2711);
and U12380 (N_12380,N_858,N_324);
and U12381 (N_12381,N_1607,N_1376);
and U12382 (N_12382,N_1684,N_3877);
nor U12383 (N_12383,N_5047,N_2889);
and U12384 (N_12384,N_1003,N_214);
nor U12385 (N_12385,N_5463,N_2463);
and U12386 (N_12386,N_3877,N_4875);
and U12387 (N_12387,N_4259,N_1224);
nand U12388 (N_12388,N_300,N_3345);
or U12389 (N_12389,N_5190,N_1810);
nand U12390 (N_12390,N_960,N_5333);
xor U12391 (N_12391,N_1354,N_646);
nor U12392 (N_12392,N_1732,N_5818);
and U12393 (N_12393,N_4774,N_2505);
or U12394 (N_12394,N_1177,N_3194);
and U12395 (N_12395,N_3982,N_360);
or U12396 (N_12396,N_1926,N_2770);
and U12397 (N_12397,N_2956,N_1283);
xor U12398 (N_12398,N_3431,N_3123);
xnor U12399 (N_12399,N_5197,N_3782);
nor U12400 (N_12400,N_5039,N_4151);
nor U12401 (N_12401,N_2689,N_1672);
xor U12402 (N_12402,N_2892,N_4577);
xor U12403 (N_12403,N_764,N_4021);
nor U12404 (N_12404,N_1708,N_5841);
xnor U12405 (N_12405,N_3727,N_3249);
or U12406 (N_12406,N_1192,N_1694);
or U12407 (N_12407,N_5165,N_205);
or U12408 (N_12408,N_873,N_230);
nand U12409 (N_12409,N_3042,N_489);
nand U12410 (N_12410,N_5791,N_5114);
or U12411 (N_12411,N_4645,N_4850);
or U12412 (N_12412,N_2753,N_4390);
or U12413 (N_12413,N_4764,N_5016);
and U12414 (N_12414,N_5215,N_2486);
xor U12415 (N_12415,N_2003,N_665);
xnor U12416 (N_12416,N_5229,N_650);
xnor U12417 (N_12417,N_2415,N_2094);
xor U12418 (N_12418,N_1414,N_1224);
and U12419 (N_12419,N_5404,N_3362);
nand U12420 (N_12420,N_4331,N_6187);
and U12421 (N_12421,N_494,N_896);
or U12422 (N_12422,N_5186,N_2022);
nor U12423 (N_12423,N_1120,N_1323);
xnor U12424 (N_12424,N_5714,N_5402);
and U12425 (N_12425,N_5274,N_290);
and U12426 (N_12426,N_969,N_4329);
nor U12427 (N_12427,N_6200,N_5391);
or U12428 (N_12428,N_5219,N_5861);
and U12429 (N_12429,N_3310,N_2418);
nor U12430 (N_12430,N_5115,N_964);
nor U12431 (N_12431,N_246,N_2259);
nand U12432 (N_12432,N_5119,N_5958);
nor U12433 (N_12433,N_4468,N_3637);
or U12434 (N_12434,N_880,N_2622);
and U12435 (N_12435,N_3343,N_5737);
and U12436 (N_12436,N_2693,N_2869);
or U12437 (N_12437,N_2126,N_5428);
nor U12438 (N_12438,N_5814,N_4348);
nand U12439 (N_12439,N_2047,N_2986);
or U12440 (N_12440,N_4503,N_252);
nand U12441 (N_12441,N_4308,N_3275);
and U12442 (N_12442,N_2945,N_2010);
nand U12443 (N_12443,N_6188,N_2916);
nand U12444 (N_12444,N_3324,N_5393);
and U12445 (N_12445,N_2655,N_3287);
nand U12446 (N_12446,N_1533,N_215);
or U12447 (N_12447,N_5141,N_2460);
nand U12448 (N_12448,N_5801,N_1072);
and U12449 (N_12449,N_518,N_770);
or U12450 (N_12450,N_2678,N_853);
and U12451 (N_12451,N_5821,N_1660);
nand U12452 (N_12452,N_1665,N_1215);
nor U12453 (N_12453,N_4266,N_4851);
and U12454 (N_12454,N_2916,N_390);
and U12455 (N_12455,N_5507,N_4492);
or U12456 (N_12456,N_325,N_3261);
nor U12457 (N_12457,N_1366,N_745);
xnor U12458 (N_12458,N_3942,N_993);
and U12459 (N_12459,N_5157,N_3069);
and U12460 (N_12460,N_2092,N_2481);
nor U12461 (N_12461,N_313,N_3978);
nand U12462 (N_12462,N_418,N_303);
xnor U12463 (N_12463,N_3592,N_613);
and U12464 (N_12464,N_4645,N_1416);
nand U12465 (N_12465,N_3451,N_137);
nor U12466 (N_12466,N_1165,N_992);
and U12467 (N_12467,N_3948,N_4800);
nand U12468 (N_12468,N_2640,N_5837);
nand U12469 (N_12469,N_5088,N_4039);
nand U12470 (N_12470,N_911,N_5588);
nor U12471 (N_12471,N_5733,N_2982);
xor U12472 (N_12472,N_1712,N_1540);
nor U12473 (N_12473,N_1621,N_286);
or U12474 (N_12474,N_3385,N_2758);
xor U12475 (N_12475,N_4052,N_4220);
nand U12476 (N_12476,N_3756,N_1044);
and U12477 (N_12477,N_1301,N_787);
nor U12478 (N_12478,N_4850,N_4483);
and U12479 (N_12479,N_1656,N_4288);
xnor U12480 (N_12480,N_6073,N_4443);
or U12481 (N_12481,N_3807,N_3440);
xnor U12482 (N_12482,N_3443,N_3435);
nor U12483 (N_12483,N_4467,N_5856);
or U12484 (N_12484,N_5796,N_3635);
nand U12485 (N_12485,N_4924,N_3253);
or U12486 (N_12486,N_2487,N_4514);
nand U12487 (N_12487,N_5931,N_2357);
nor U12488 (N_12488,N_400,N_2634);
nor U12489 (N_12489,N_5359,N_4023);
and U12490 (N_12490,N_3636,N_1435);
or U12491 (N_12491,N_4783,N_3224);
xor U12492 (N_12492,N_2387,N_830);
or U12493 (N_12493,N_5757,N_4094);
xor U12494 (N_12494,N_4327,N_5628);
and U12495 (N_12495,N_1053,N_3927);
and U12496 (N_12496,N_222,N_2477);
and U12497 (N_12497,N_5862,N_4139);
or U12498 (N_12498,N_522,N_4162);
or U12499 (N_12499,N_5840,N_1742);
nand U12500 (N_12500,N_6987,N_7575);
nor U12501 (N_12501,N_11967,N_8097);
nor U12502 (N_12502,N_8431,N_8759);
and U12503 (N_12503,N_10764,N_11398);
or U12504 (N_12504,N_10968,N_12204);
and U12505 (N_12505,N_11606,N_7699);
and U12506 (N_12506,N_11055,N_8117);
nor U12507 (N_12507,N_12337,N_12143);
or U12508 (N_12508,N_9075,N_10782);
nor U12509 (N_12509,N_9096,N_11850);
nor U12510 (N_12510,N_7022,N_10237);
nor U12511 (N_12511,N_6337,N_11065);
xor U12512 (N_12512,N_11081,N_8495);
xor U12513 (N_12513,N_7994,N_11527);
nor U12514 (N_12514,N_8567,N_9407);
xnor U12515 (N_12515,N_9135,N_9117);
nor U12516 (N_12516,N_10308,N_9121);
nor U12517 (N_12517,N_9528,N_8150);
nand U12518 (N_12518,N_7050,N_6674);
nor U12519 (N_12519,N_11474,N_10527);
and U12520 (N_12520,N_11135,N_8357);
nand U12521 (N_12521,N_7724,N_8995);
and U12522 (N_12522,N_11202,N_10479);
nor U12523 (N_12523,N_12127,N_8068);
nand U12524 (N_12524,N_9197,N_8436);
nor U12525 (N_12525,N_8813,N_10869);
xnor U12526 (N_12526,N_9378,N_7784);
xor U12527 (N_12527,N_8943,N_11704);
xnor U12528 (N_12528,N_9425,N_11936);
xor U12529 (N_12529,N_9515,N_7058);
nand U12530 (N_12530,N_11825,N_9364);
xnor U12531 (N_12531,N_9835,N_9230);
xor U12532 (N_12532,N_10844,N_7770);
nand U12533 (N_12533,N_10459,N_10695);
nand U12534 (N_12534,N_8365,N_8289);
nand U12535 (N_12535,N_7509,N_10273);
or U12536 (N_12536,N_11532,N_11289);
nor U12537 (N_12537,N_12488,N_11663);
xor U12538 (N_12538,N_11777,N_6372);
xnor U12539 (N_12539,N_9661,N_11981);
xor U12540 (N_12540,N_9258,N_11024);
and U12541 (N_12541,N_11662,N_9449);
nor U12542 (N_12542,N_7074,N_12300);
or U12543 (N_12543,N_11915,N_6681);
nand U12544 (N_12544,N_9306,N_11833);
nor U12545 (N_12545,N_7277,N_8958);
xor U12546 (N_12546,N_11493,N_9108);
xnor U12547 (N_12547,N_8184,N_7079);
and U12548 (N_12548,N_9134,N_8213);
or U12549 (N_12549,N_10142,N_6954);
or U12550 (N_12550,N_11929,N_8796);
xnor U12551 (N_12551,N_9426,N_8073);
xnor U12552 (N_12552,N_6883,N_6630);
or U12553 (N_12553,N_8816,N_11178);
and U12554 (N_12554,N_11014,N_11690);
nand U12555 (N_12555,N_9721,N_11297);
nand U12556 (N_12556,N_6426,N_9332);
xnor U12557 (N_12557,N_9756,N_12291);
nand U12558 (N_12558,N_9138,N_7213);
nand U12559 (N_12559,N_10955,N_11896);
xor U12560 (N_12560,N_12429,N_9583);
nand U12561 (N_12561,N_7665,N_11802);
and U12562 (N_12562,N_8059,N_9260);
nor U12563 (N_12563,N_8901,N_10430);
nor U12564 (N_12564,N_7025,N_8680);
nand U12565 (N_12565,N_10461,N_7250);
or U12566 (N_12566,N_7227,N_12314);
and U12567 (N_12567,N_9119,N_10973);
nand U12568 (N_12568,N_8502,N_11807);
nand U12569 (N_12569,N_7670,N_9019);
nor U12570 (N_12570,N_6633,N_9485);
nor U12571 (N_12571,N_7864,N_7568);
nor U12572 (N_12572,N_8610,N_10948);
and U12573 (N_12573,N_9857,N_8657);
xor U12574 (N_12574,N_6367,N_11630);
nor U12575 (N_12575,N_9503,N_9251);
nor U12576 (N_12576,N_10601,N_8626);
xor U12577 (N_12577,N_6490,N_7194);
and U12578 (N_12578,N_10903,N_7734);
xor U12579 (N_12579,N_9939,N_7481);
nand U12580 (N_12580,N_11190,N_7020);
nand U12581 (N_12581,N_7092,N_6658);
or U12582 (N_12582,N_12355,N_6469);
nor U12583 (N_12583,N_6381,N_10553);
xnor U12584 (N_12584,N_11550,N_12255);
nand U12585 (N_12585,N_7122,N_7732);
nand U12586 (N_12586,N_11449,N_11684);
nand U12587 (N_12587,N_9326,N_10696);
nor U12588 (N_12588,N_10128,N_8472);
and U12589 (N_12589,N_11084,N_9816);
nor U12590 (N_12590,N_11218,N_11914);
or U12591 (N_12591,N_8999,N_10211);
nor U12592 (N_12592,N_10954,N_10909);
or U12593 (N_12593,N_7212,N_7334);
nor U12594 (N_12594,N_10737,N_7660);
nand U12595 (N_12595,N_8849,N_8772);
nand U12596 (N_12596,N_6645,N_6439);
xnor U12597 (N_12597,N_12360,N_6877);
nand U12598 (N_12598,N_12330,N_10173);
nand U12599 (N_12599,N_9546,N_8486);
xnor U12600 (N_12600,N_6753,N_10453);
and U12601 (N_12601,N_9151,N_6431);
or U12602 (N_12602,N_7725,N_8276);
or U12603 (N_12603,N_11245,N_11443);
nor U12604 (N_12604,N_12059,N_7842);
nand U12605 (N_12605,N_8799,N_10428);
nand U12606 (N_12606,N_7901,N_6863);
nor U12607 (N_12607,N_7570,N_11828);
or U12608 (N_12608,N_10230,N_11219);
nor U12609 (N_12609,N_8028,N_8722);
nand U12610 (N_12610,N_11234,N_8527);
and U12611 (N_12611,N_12113,N_11043);
or U12612 (N_12612,N_9498,N_9808);
nand U12613 (N_12613,N_6548,N_9871);
nand U12614 (N_12614,N_7633,N_10834);
or U12615 (N_12615,N_9545,N_7309);
and U12616 (N_12616,N_8955,N_12106);
or U12617 (N_12617,N_11384,N_9133);
or U12618 (N_12618,N_11291,N_8423);
nor U12619 (N_12619,N_8079,N_7240);
xnor U12620 (N_12620,N_11912,N_6557);
nor U12621 (N_12621,N_9214,N_6796);
and U12622 (N_12622,N_7877,N_9368);
or U12623 (N_12623,N_6972,N_7367);
xnor U12624 (N_12624,N_7905,N_12240);
xor U12625 (N_12625,N_6566,N_7011);
nand U12626 (N_12626,N_8092,N_10987);
or U12627 (N_12627,N_11045,N_8319);
xnor U12628 (N_12628,N_11950,N_11293);
or U12629 (N_12629,N_8043,N_8784);
or U12630 (N_12630,N_7483,N_12088);
or U12631 (N_12631,N_10106,N_10496);
and U12632 (N_12632,N_7121,N_8936);
nor U12633 (N_12633,N_11191,N_9352);
and U12634 (N_12634,N_6653,N_6483);
and U12635 (N_12635,N_9313,N_11714);
and U12636 (N_12636,N_12420,N_9366);
nand U12637 (N_12637,N_12254,N_12116);
nand U12638 (N_12638,N_10557,N_8854);
xor U12639 (N_12639,N_8204,N_10191);
nor U12640 (N_12640,N_9596,N_12168);
and U12641 (N_12641,N_9188,N_12220);
nand U12642 (N_12642,N_7314,N_10049);
and U12643 (N_12643,N_9113,N_6870);
nor U12644 (N_12644,N_11327,N_11491);
or U12645 (N_12645,N_11926,N_12152);
nand U12646 (N_12646,N_11283,N_12378);
nor U12647 (N_12647,N_9310,N_8393);
xnor U12648 (N_12648,N_7101,N_9249);
and U12649 (N_12649,N_11332,N_8424);
nor U12650 (N_12650,N_12008,N_7142);
or U12651 (N_12651,N_7005,N_10202);
xnor U12652 (N_12652,N_12262,N_11296);
nor U12653 (N_12653,N_6886,N_9376);
or U12654 (N_12654,N_10370,N_6656);
and U12655 (N_12655,N_8435,N_10139);
nor U12656 (N_12656,N_9571,N_7696);
and U12657 (N_12657,N_6599,N_9698);
and U12658 (N_12658,N_8636,N_10295);
nor U12659 (N_12659,N_11287,N_9496);
or U12660 (N_12660,N_12323,N_7581);
xor U12661 (N_12661,N_7669,N_9719);
nor U12662 (N_12662,N_12099,N_9938);
and U12663 (N_12663,N_7698,N_6628);
and U12664 (N_12664,N_7681,N_6510);
or U12665 (N_12665,N_12258,N_10243);
xor U12666 (N_12666,N_9115,N_8199);
xnor U12667 (N_12667,N_10085,N_10424);
or U12668 (N_12668,N_10422,N_10267);
or U12669 (N_12669,N_9143,N_7221);
and U12670 (N_12670,N_7263,N_11204);
xnor U12671 (N_12671,N_6890,N_8866);
or U12672 (N_12672,N_7517,N_11356);
xor U12673 (N_12673,N_7590,N_12375);
nand U12674 (N_12674,N_10187,N_7223);
nor U12675 (N_12675,N_7152,N_11688);
and U12676 (N_12676,N_9293,N_7645);
or U12677 (N_12677,N_6934,N_11700);
nor U12678 (N_12678,N_9131,N_9463);
and U12679 (N_12679,N_9829,N_11539);
xnor U12680 (N_12680,N_10227,N_10642);
nor U12681 (N_12681,N_7835,N_10417);
nand U12682 (N_12682,N_11280,N_7700);
xor U12683 (N_12683,N_9632,N_6986);
nor U12684 (N_12684,N_9412,N_11972);
xnor U12685 (N_12685,N_8152,N_7392);
and U12686 (N_12686,N_10916,N_10238);
nor U12687 (N_12687,N_9123,N_9103);
xor U12688 (N_12688,N_12095,N_7723);
nor U12689 (N_12689,N_9098,N_12159);
or U12690 (N_12690,N_8130,N_10821);
or U12691 (N_12691,N_8447,N_10153);
nor U12692 (N_12692,N_9387,N_8053);
xnor U12693 (N_12693,N_7515,N_8571);
xnor U12694 (N_12694,N_7053,N_7084);
xor U12695 (N_12695,N_11778,N_6375);
and U12696 (N_12696,N_8157,N_11567);
nand U12697 (N_12697,N_9041,N_8815);
nor U12698 (N_12698,N_6563,N_9850);
nor U12699 (N_12699,N_11028,N_11042);
xor U12700 (N_12700,N_7261,N_7709);
and U12701 (N_12701,N_9691,N_11713);
xor U12702 (N_12702,N_11795,N_8056);
and U12703 (N_12703,N_10577,N_6787);
nand U12704 (N_12704,N_12174,N_8604);
nor U12705 (N_12705,N_12303,N_12273);
and U12706 (N_12706,N_7939,N_9591);
xnor U12707 (N_12707,N_12440,N_7322);
and U12708 (N_12708,N_9551,N_9811);
nor U12709 (N_12709,N_8003,N_10311);
and U12710 (N_12710,N_9985,N_8081);
nor U12711 (N_12711,N_7695,N_9956);
or U12712 (N_12712,N_11397,N_7520);
nor U12713 (N_12713,N_6290,N_7416);
and U12714 (N_12714,N_10068,N_9475);
or U12715 (N_12715,N_10051,N_10907);
xnor U12716 (N_12716,N_7693,N_11895);
nor U12717 (N_12717,N_7529,N_7503);
or U12718 (N_12718,N_7694,N_9071);
and U12719 (N_12719,N_8774,N_9641);
and U12720 (N_12720,N_8290,N_6725);
nor U12721 (N_12721,N_9962,N_7762);
or U12722 (N_12722,N_8463,N_9490);
nand U12723 (N_12723,N_12069,N_12126);
or U12724 (N_12724,N_7739,N_10827);
nor U12725 (N_12725,N_8453,N_7801);
nand U12726 (N_12726,N_7916,N_12012);
xor U12727 (N_12727,N_11412,N_8979);
xnor U12728 (N_12728,N_8175,N_7903);
and U12729 (N_12729,N_8932,N_7598);
and U12730 (N_12730,N_9552,N_12237);
and U12731 (N_12731,N_8616,N_6379);
xor U12732 (N_12732,N_8906,N_7546);
xor U12733 (N_12733,N_10998,N_8197);
nand U12734 (N_12734,N_8889,N_7411);
xor U12735 (N_12735,N_8253,N_6974);
xnor U12736 (N_12736,N_10621,N_12402);
nor U12737 (N_12737,N_12392,N_6727);
or U12738 (N_12738,N_11726,N_11908);
or U12739 (N_12739,N_8539,N_7655);
nand U12740 (N_12740,N_9921,N_11920);
xor U12741 (N_12741,N_8761,N_10358);
nor U12742 (N_12742,N_11852,N_8650);
nand U12743 (N_12743,N_11371,N_8538);
or U12744 (N_12744,N_12413,N_10426);
or U12745 (N_12745,N_7430,N_9064);
and U12746 (N_12746,N_6983,N_8893);
xor U12747 (N_12747,N_10975,N_7539);
and U12748 (N_12748,N_12002,N_10645);
or U12749 (N_12749,N_6866,N_6559);
nand U12750 (N_12750,N_11607,N_8509);
xor U12751 (N_12751,N_8376,N_10419);
or U12752 (N_12752,N_7764,N_8855);
nor U12753 (N_12753,N_6688,N_9150);
or U12754 (N_12754,N_6925,N_7181);
nor U12755 (N_12755,N_6635,N_7313);
nor U12756 (N_12756,N_8755,N_12217);
and U12757 (N_12757,N_11945,N_6466);
nand U12758 (N_12758,N_7863,N_8069);
or U12759 (N_12759,N_6542,N_11946);
nor U12760 (N_12760,N_6419,N_12064);
nor U12761 (N_12761,N_10061,N_11007);
nand U12762 (N_12762,N_11983,N_10590);
xnor U12763 (N_12763,N_7302,N_9862);
nand U12764 (N_12764,N_8550,N_11576);
xor U12765 (N_12765,N_6835,N_7021);
nand U12766 (N_12766,N_11438,N_6506);
nand U12767 (N_12767,N_11281,N_10905);
or U12768 (N_12768,N_6931,N_10515);
and U12769 (N_12769,N_9421,N_9038);
nand U12770 (N_12770,N_7034,N_11783);
or U12771 (N_12771,N_7118,N_9523);
and U12772 (N_12772,N_9981,N_6670);
xor U12773 (N_12773,N_11054,N_12162);
and U12774 (N_12774,N_9036,N_12144);
and U12775 (N_12775,N_8768,N_7138);
nor U12776 (N_12776,N_9062,N_7950);
nand U12777 (N_12777,N_8649,N_8615);
nand U12778 (N_12778,N_7549,N_8421);
nand U12779 (N_12779,N_6701,N_8205);
nor U12780 (N_12780,N_10162,N_10258);
or U12781 (N_12781,N_6301,N_12053);
nor U12782 (N_12782,N_12470,N_9001);
xnor U12783 (N_12783,N_6749,N_11038);
and U12784 (N_12784,N_6932,N_6823);
and U12785 (N_12785,N_6640,N_8648);
and U12786 (N_12786,N_6370,N_8731);
nor U12787 (N_12787,N_9093,N_6343);
nand U12788 (N_12788,N_7648,N_7913);
xnor U12789 (N_12789,N_11413,N_9281);
or U12790 (N_12790,N_6945,N_7596);
nor U12791 (N_12791,N_9029,N_8929);
nand U12792 (N_12792,N_11520,N_7757);
xnor U12793 (N_12793,N_9454,N_7679);
nor U12794 (N_12794,N_11685,N_10159);
or U12795 (N_12795,N_9331,N_8168);
xor U12796 (N_12796,N_8656,N_11615);
or U12797 (N_12797,N_8320,N_9580);
and U12798 (N_12798,N_9502,N_12032);
nand U12799 (N_12799,N_7871,N_8831);
nand U12800 (N_12800,N_8349,N_9320);
or U12801 (N_12801,N_7941,N_7512);
and U12802 (N_12802,N_12308,N_11667);
or U12803 (N_12803,N_9003,N_11057);
or U12804 (N_12804,N_11166,N_11757);
nand U12805 (N_12805,N_8040,N_12453);
xor U12806 (N_12806,N_10836,N_9520);
or U12807 (N_12807,N_11011,N_10081);
nand U12808 (N_12808,N_6486,N_8544);
nand U12809 (N_12809,N_6321,N_11127);
or U12810 (N_12810,N_11987,N_9586);
and U12811 (N_12811,N_8261,N_11435);
and U12812 (N_12812,N_11102,N_10890);
nor U12813 (N_12813,N_10993,N_8194);
nor U12814 (N_12814,N_12007,N_9484);
or U12815 (N_12815,N_7333,N_6554);
nand U12816 (N_12816,N_6963,N_8008);
and U12817 (N_12817,N_10190,N_11686);
and U12818 (N_12818,N_11486,N_11032);
nand U12819 (N_12819,N_7288,N_9012);
or U12820 (N_12820,N_10877,N_9955);
or U12821 (N_12821,N_9902,N_11149);
xnor U12822 (N_12822,N_6316,N_10866);
or U12823 (N_12823,N_9457,N_7867);
nand U12824 (N_12824,N_9276,N_10565);
and U12825 (N_12825,N_9238,N_7667);
and U12826 (N_12826,N_9741,N_6671);
nand U12827 (N_12827,N_11411,N_11818);
nand U12828 (N_12828,N_10130,N_10390);
xnor U12829 (N_12829,N_10562,N_7720);
and U12830 (N_12830,N_11565,N_7834);
or U12831 (N_12831,N_8835,N_6643);
nor U12832 (N_12832,N_9349,N_12370);
nand U12833 (N_12833,N_12349,N_7673);
or U12834 (N_12834,N_10271,N_9400);
xnor U12835 (N_12835,N_11571,N_8853);
nand U12836 (N_12836,N_12114,N_8852);
and U12837 (N_12837,N_9726,N_11814);
and U12838 (N_12838,N_11592,N_9101);
or U12839 (N_12839,N_6371,N_11910);
or U12840 (N_12840,N_8129,N_9157);
nor U12841 (N_12841,N_9519,N_12456);
nor U12842 (N_12842,N_8569,N_9162);
or U12843 (N_12843,N_12476,N_7358);
or U12844 (N_12844,N_12421,N_8823);
nor U12845 (N_12845,N_11703,N_11484);
xnor U12846 (N_12846,N_11931,N_9898);
xor U12847 (N_12847,N_6806,N_10962);
or U12848 (N_12848,N_6341,N_6523);
or U12849 (N_12849,N_11259,N_6784);
and U12850 (N_12850,N_11473,N_6752);
or U12851 (N_12851,N_11430,N_9876);
nand U12852 (N_12852,N_12381,N_10058);
nor U12853 (N_12853,N_6276,N_8914);
nor U12854 (N_12854,N_8283,N_8167);
nand U12855 (N_12855,N_9774,N_11151);
nand U12856 (N_12856,N_9507,N_8337);
and U12857 (N_12857,N_8325,N_12350);
nor U12858 (N_12858,N_9290,N_6982);
nor U12859 (N_12859,N_7294,N_8543);
nor U12860 (N_12860,N_10701,N_9236);
and U12861 (N_12861,N_9911,N_11722);
nand U12862 (N_12862,N_8444,N_7295);
nor U12863 (N_12863,N_6973,N_8187);
or U12864 (N_12864,N_11720,N_11596);
xnor U12865 (N_12865,N_7153,N_7767);
nor U12866 (N_12866,N_10352,N_11803);
or U12867 (N_12867,N_6838,N_9055);
nand U12868 (N_12868,N_8702,N_10674);
or U12869 (N_12869,N_9705,N_8726);
xnor U12870 (N_12870,N_8153,N_9164);
and U12871 (N_12871,N_9799,N_6481);
or U12872 (N_12872,N_11209,N_10514);
nand U12873 (N_12873,N_11035,N_10923);
nor U12874 (N_12874,N_7935,N_8333);
nand U12875 (N_12875,N_9713,N_11712);
nand U12876 (N_12876,N_11605,N_12347);
nor U12877 (N_12877,N_9779,N_6757);
and U12878 (N_12878,N_11088,N_7131);
nor U12879 (N_12879,N_7792,N_7637);
xor U12880 (N_12880,N_7861,N_8050);
and U12881 (N_12881,N_9935,N_12425);
xnor U12882 (N_12882,N_12183,N_11897);
xnor U12883 (N_12883,N_9148,N_6418);
and U12884 (N_12884,N_11153,N_9766);
nor U12885 (N_12885,N_7113,N_11086);
nor U12886 (N_12886,N_9934,N_12487);
nand U12887 (N_12887,N_11309,N_11436);
and U12888 (N_12888,N_6434,N_11258);
or U12889 (N_12889,N_9609,N_7253);
and U12890 (N_12890,N_7530,N_8006);
xnor U12891 (N_12891,N_12187,N_10414);
xor U12892 (N_12892,N_8925,N_7752);
nor U12893 (N_12893,N_7771,N_6637);
xor U12894 (N_12894,N_12417,N_8907);
nor U12895 (N_12895,N_8264,N_10495);
and U12896 (N_12896,N_8963,N_6444);
nor U12897 (N_12897,N_12416,N_10828);
and U12898 (N_12898,N_9652,N_6606);
nand U12899 (N_12899,N_6257,N_7028);
nor U12900 (N_12900,N_10756,N_10961);
xor U12901 (N_12901,N_10855,N_7356);
nand U12902 (N_12902,N_9220,N_9777);
xnor U12903 (N_12903,N_11919,N_7066);
nor U12904 (N_12904,N_8501,N_11847);
or U12905 (N_12905,N_9289,N_7843);
nand U12906 (N_12906,N_11229,N_10133);
nor U12907 (N_12907,N_7711,N_10730);
nor U12908 (N_12908,N_11938,N_11104);
nor U12909 (N_12909,N_11008,N_10145);
or U12910 (N_12910,N_8978,N_8260);
xor U12911 (N_12911,N_10926,N_9600);
xor U12912 (N_12912,N_11797,N_12361);
xnor U12913 (N_12913,N_7249,N_9428);
nor U12914 (N_12914,N_8181,N_7957);
and U12915 (N_12915,N_12110,N_11900);
nor U12916 (N_12916,N_8678,N_6509);
and U12917 (N_12917,N_9217,N_6858);
xnor U12918 (N_12918,N_10879,N_12139);
nor U12919 (N_12919,N_7988,N_9971);
nand U12920 (N_12920,N_8491,N_11124);
and U12921 (N_12921,N_6765,N_10574);
nor U12922 (N_12922,N_11964,N_9644);
nor U12923 (N_12923,N_8787,N_12023);
nand U12924 (N_12924,N_11528,N_8652);
nand U12925 (N_12925,N_7866,N_7773);
nand U12926 (N_12926,N_7692,N_11740);
nand U12927 (N_12927,N_11325,N_11590);
xor U12928 (N_12928,N_8824,N_7032);
and U12929 (N_12929,N_10210,N_7737);
xor U12930 (N_12930,N_6978,N_10681);
xor U12931 (N_12931,N_7875,N_8669);
or U12932 (N_12932,N_6334,N_8860);
nand U12933 (N_12933,N_9063,N_7558);
nand U12934 (N_12934,N_12184,N_8467);
and U12935 (N_12935,N_7977,N_8315);
nand U12936 (N_12936,N_11957,N_8668);
xnor U12937 (N_12937,N_7403,N_10491);
and U12938 (N_12938,N_11587,N_10024);
and U12939 (N_12939,N_7576,N_6297);
nor U12940 (N_12940,N_9852,N_7970);
xor U12941 (N_12941,N_8331,N_8352);
or U12942 (N_12942,N_11425,N_8448);
and U12943 (N_12943,N_12197,N_10952);
and U12944 (N_12944,N_9703,N_7146);
or U12945 (N_12945,N_8126,N_8875);
or U12946 (N_12946,N_11534,N_8944);
and U12947 (N_12947,N_7386,N_10194);
and U12948 (N_12948,N_6501,N_8859);
nand U12949 (N_12949,N_10945,N_8520);
and U12950 (N_12950,N_11133,N_9834);
and U12951 (N_12951,N_7218,N_12015);
and U12952 (N_12952,N_6284,N_9288);
nand U12953 (N_12953,N_12075,N_10249);
nor U12954 (N_12954,N_10279,N_11303);
nand U12955 (N_12955,N_8977,N_7824);
nand U12956 (N_12956,N_11171,N_9690);
xor U12957 (N_12957,N_6496,N_9683);
and U12958 (N_12958,N_10092,N_10792);
nand U12959 (N_12959,N_6780,N_9184);
nor U12960 (N_12960,N_10611,N_8640);
and U12961 (N_12961,N_6785,N_8957);
or U12962 (N_12962,N_11480,N_7346);
and U12963 (N_12963,N_7758,N_8471);
xor U12964 (N_12964,N_9562,N_11516);
or U12965 (N_12965,N_10676,N_10829);
or U12966 (N_12966,N_8177,N_8517);
and U12967 (N_12967,N_12316,N_9040);
and U12968 (N_12968,N_6848,N_8601);
or U12969 (N_12969,N_11215,N_7488);
xor U12970 (N_12970,N_9822,N_6853);
xnor U12971 (N_12971,N_12047,N_10113);
and U12972 (N_12972,N_8113,N_8840);
and U12973 (N_12973,N_7252,N_9088);
xnor U12974 (N_12974,N_9851,N_10337);
nand U12975 (N_12975,N_11854,N_7004);
and U12976 (N_12976,N_9044,N_12105);
and U12977 (N_12977,N_9754,N_11706);
or U12978 (N_12978,N_9870,N_11786);
nand U12979 (N_12979,N_9043,N_7039);
nor U12980 (N_12980,N_11119,N_9073);
nor U12981 (N_12981,N_9727,N_8255);
xnor U12982 (N_12982,N_9453,N_8387);
or U12983 (N_12983,N_7271,N_11760);
or U12984 (N_12984,N_11591,N_8727);
or U12985 (N_12985,N_9518,N_10144);
nor U12986 (N_12986,N_8545,N_11136);
nand U12987 (N_12987,N_12387,N_9124);
and U12988 (N_12988,N_9893,N_8525);
nor U12989 (N_12989,N_7583,N_11198);
and U12990 (N_12990,N_10920,N_9970);
nor U12991 (N_12991,N_7810,N_11101);
nor U12992 (N_12992,N_6894,N_7465);
or U12993 (N_12993,N_8207,N_7310);
nor U12994 (N_12994,N_8735,N_11792);
or U12995 (N_12995,N_7373,N_10885);
xor U12996 (N_12996,N_8653,N_11562);
nand U12997 (N_12997,N_11622,N_11745);
or U12998 (N_12998,N_10541,N_8821);
and U12999 (N_12999,N_9599,N_10825);
xor U13000 (N_13000,N_6867,N_11147);
xor U13001 (N_13001,N_8710,N_6369);
xor U13002 (N_13002,N_9460,N_7371);
xor U13003 (N_13003,N_9606,N_9536);
or U13004 (N_13004,N_10341,N_6634);
or U13005 (N_13005,N_9350,N_9452);
or U13006 (N_13006,N_10137,N_10623);
and U13007 (N_13007,N_7143,N_10765);
and U13008 (N_13008,N_8535,N_8679);
nand U13009 (N_13009,N_10080,N_7231);
xnor U13010 (N_13010,N_9399,N_11793);
xnor U13011 (N_13011,N_12092,N_9418);
nor U13012 (N_13012,N_10534,N_10462);
xnor U13013 (N_13013,N_12063,N_12119);
xnor U13014 (N_13014,N_7653,N_9176);
or U13015 (N_13015,N_9805,N_9990);
nand U13016 (N_13016,N_9190,N_7907);
xor U13017 (N_13017,N_11305,N_11231);
nor U13018 (N_13018,N_11079,N_9798);
xor U13019 (N_13019,N_12382,N_12054);
nor U13020 (N_13020,N_9607,N_8847);
or U13021 (N_13021,N_7013,N_10849);
nor U13022 (N_13022,N_12109,N_9333);
and U13023 (N_13023,N_7608,N_10738);
and U13024 (N_13024,N_7363,N_12028);
and U13025 (N_13025,N_6900,N_7287);
xor U13026 (N_13026,N_7216,N_9890);
nand U13027 (N_13027,N_8627,N_9000);
nor U13028 (N_13028,N_11246,N_8512);
or U13029 (N_13029,N_8766,N_11482);
and U13030 (N_13030,N_10433,N_10779);
and U13031 (N_13031,N_7427,N_10010);
nand U13032 (N_13032,N_9226,N_8872);
and U13033 (N_13033,N_9027,N_8432);
and U13034 (N_13034,N_6377,N_8286);
and U13035 (N_13035,N_9855,N_10704);
nor U13036 (N_13036,N_8803,N_6685);
or U13037 (N_13037,N_7697,N_6463);
nand U13038 (N_13038,N_8599,N_9576);
or U13039 (N_13039,N_8725,N_8138);
nand U13040 (N_13040,N_9988,N_8381);
xnor U13041 (N_13041,N_10427,N_7006);
or U13042 (N_13042,N_6829,N_9628);
nand U13043 (N_13043,N_7380,N_9964);
nand U13044 (N_13044,N_10861,N_7639);
nand U13045 (N_13045,N_7029,N_9380);
xor U13046 (N_13046,N_10294,N_11140);
and U13047 (N_13047,N_10075,N_9321);
or U13048 (N_13048,N_10192,N_11588);
and U13049 (N_13049,N_11865,N_9780);
or U13050 (N_13050,N_6650,N_6353);
or U13051 (N_13051,N_6440,N_10285);
xor U13052 (N_13052,N_7836,N_6811);
and U13053 (N_13053,N_9601,N_6411);
and U13054 (N_13054,N_11942,N_6511);
or U13055 (N_13055,N_11775,N_8593);
or U13056 (N_13056,N_9068,N_9383);
xnor U13057 (N_13057,N_6995,N_10015);
and U13058 (N_13058,N_9612,N_10437);
and U13059 (N_13059,N_9894,N_9104);
nand U13060 (N_13060,N_11376,N_10739);
nand U13061 (N_13061,N_10027,N_8733);
or U13062 (N_13062,N_6346,N_10763);
xnor U13063 (N_13063,N_7301,N_7087);
nand U13064 (N_13064,N_7541,N_11358);
nor U13065 (N_13065,N_12085,N_11352);
nor U13066 (N_13066,N_6465,N_7329);
or U13067 (N_13067,N_7148,N_7279);
nand U13068 (N_13068,N_7200,N_6741);
xnor U13069 (N_13069,N_10841,N_10118);
and U13070 (N_13070,N_10356,N_6468);
and U13071 (N_13071,N_9759,N_7147);
xnor U13072 (N_13072,N_9737,N_11187);
and U13073 (N_13073,N_12005,N_10780);
xnor U13074 (N_13074,N_9299,N_7414);
or U13075 (N_13075,N_9587,N_7384);
nand U13076 (N_13076,N_10473,N_10691);
and U13077 (N_13077,N_6578,N_9836);
xnor U13078 (N_13078,N_11122,N_11611);
nand U13079 (N_13079,N_9720,N_12141);
nand U13080 (N_13080,N_11235,N_11469);
and U13081 (N_13081,N_11566,N_9023);
nand U13082 (N_13082,N_9813,N_9567);
xor U13083 (N_13083,N_7401,N_7353);
and U13084 (N_13084,N_9327,N_6362);
and U13085 (N_13085,N_11432,N_11991);
xor U13086 (N_13086,N_12253,N_11374);
xor U13087 (N_13087,N_12169,N_7788);
nand U13088 (N_13088,N_6907,N_7811);
and U13089 (N_13089,N_7335,N_11761);
xnor U13090 (N_13090,N_11403,N_6275);
nor U13091 (N_13091,N_8674,N_7543);
or U13092 (N_13092,N_9608,N_11570);
xnor U13093 (N_13093,N_8613,N_8555);
and U13094 (N_13094,N_8004,N_8306);
or U13095 (N_13095,N_8715,N_6748);
nor U13096 (N_13096,N_10588,N_10689);
nor U13097 (N_13097,N_7183,N_6664);
nand U13098 (N_13098,N_7973,N_11838);
xnor U13099 (N_13099,N_6852,N_8721);
or U13100 (N_13100,N_7874,N_10537);
xor U13101 (N_13101,N_12292,N_11978);
or U13102 (N_13102,N_8402,N_11314);
and U13103 (N_13103,N_6956,N_8104);
and U13104 (N_13104,N_6941,N_8347);
and U13105 (N_13105,N_6289,N_11072);
xnor U13106 (N_13106,N_8115,N_6891);
or U13107 (N_13107,N_11940,N_10291);
nand U13108 (N_13108,N_11426,N_11800);
or U13109 (N_13109,N_10421,N_8494);
xnor U13110 (N_13110,N_7425,N_10454);
nor U13111 (N_13111,N_11660,N_7270);
or U13112 (N_13112,N_11409,N_8924);
xnor U13113 (N_13113,N_9992,N_11697);
nand U13114 (N_13114,N_10203,N_6473);
nor U13115 (N_13115,N_11173,N_8927);
nor U13116 (N_13116,N_12394,N_9618);
xor U13117 (N_13117,N_11909,N_10797);
nor U13118 (N_13118,N_11820,N_7439);
or U13119 (N_13119,N_9298,N_9061);
and U13120 (N_13120,N_11971,N_8108);
xor U13121 (N_13121,N_8506,N_7354);
and U13122 (N_13122,N_7691,N_12084);
and U13123 (N_13123,N_11969,N_10893);
nand U13124 (N_13124,N_10725,N_8166);
or U13125 (N_13125,N_9611,N_8921);
xnor U13126 (N_13126,N_10355,N_8714);
nand U13127 (N_13127,N_10316,N_8987);
or U13128 (N_13128,N_11621,N_10157);
and U13129 (N_13129,N_10528,N_6998);
xor U13130 (N_13130,N_9508,N_11393);
and U13131 (N_13131,N_6743,N_11018);
xnor U13132 (N_13132,N_11274,N_7554);
or U13133 (N_13133,N_12430,N_11646);
nor U13134 (N_13134,N_11666,N_7680);
or U13135 (N_13135,N_10630,N_8666);
or U13136 (N_13136,N_9464,N_9139);
or U13137 (N_13137,N_7330,N_11742);
nand U13138 (N_13138,N_11804,N_12409);
or U13139 (N_13139,N_12020,N_9729);
xor U13140 (N_13140,N_10659,N_11597);
or U13141 (N_13141,N_12228,N_7870);
xnor U13142 (N_13142,N_9677,N_11346);
or U13143 (N_13143,N_6885,N_7248);
nor U13144 (N_13144,N_9370,N_10372);
nor U13145 (N_13145,N_7951,N_12408);
or U13146 (N_13146,N_6282,N_6397);
or U13147 (N_13147,N_9838,N_11682);
xor U13148 (N_13148,N_9959,N_8949);
and U13149 (N_13149,N_6383,N_9919);
nand U13150 (N_13150,N_7009,N_7436);
xnor U13151 (N_13151,N_8737,N_11462);
or U13152 (N_13152,N_6544,N_6846);
or U13153 (N_13153,N_9560,N_8080);
or U13154 (N_13154,N_9328,N_9173);
or U13155 (N_13155,N_11157,N_11442);
xnor U13156 (N_13156,N_8546,N_11354);
xor U13157 (N_13157,N_7001,N_10147);
and U13158 (N_13158,N_10759,N_11734);
or U13159 (N_13159,N_9769,N_6423);
and U13160 (N_13160,N_11117,N_8176);
nor U13161 (N_13161,N_11600,N_7315);
nor U13162 (N_13162,N_6647,N_8488);
nor U13163 (N_13163,N_7462,N_10042);
nor U13164 (N_13164,N_6564,N_7266);
xnor U13165 (N_13165,N_7306,N_11694);
or U13166 (N_13166,N_7890,N_10361);
or U13167 (N_13167,N_10530,N_10573);
or U13168 (N_13168,N_10062,N_9840);
and U13169 (N_13169,N_8894,N_8102);
nand U13170 (N_13170,N_7379,N_11970);
nor U13171 (N_13171,N_10902,N_7735);
nor U13172 (N_13172,N_6839,N_10149);
nand U13173 (N_13173,N_7328,N_7246);
nand U13174 (N_13174,N_11519,N_12432);
or U13175 (N_13175,N_7895,N_9848);
or U13176 (N_13176,N_11139,N_6560);
and U13177 (N_13177,N_7573,N_10852);
xnor U13178 (N_13178,N_8985,N_6617);
nand U13179 (N_13179,N_6756,N_8795);
xnor U13180 (N_13180,N_7477,N_10761);
nor U13181 (N_13181,N_12200,N_10098);
and U13182 (N_13182,N_7292,N_9736);
nor U13183 (N_13183,N_10912,N_11790);
or U13184 (N_13184,N_11155,N_10066);
and U13185 (N_13185,N_11064,N_6504);
nor U13186 (N_13186,N_8976,N_12158);
or U13187 (N_13187,N_9666,N_10303);
nor U13188 (N_13188,N_7684,N_9353);
nor U13189 (N_13189,N_6642,N_9787);
and U13190 (N_13190,N_8235,N_11873);
or U13191 (N_13191,N_7601,N_7803);
or U13192 (N_13192,N_12275,N_12401);
or U13193 (N_13193,N_11750,N_7617);
nand U13194 (N_13194,N_7360,N_10654);
and U13195 (N_13195,N_6804,N_10972);
nor U13196 (N_13196,N_11944,N_11886);
nand U13197 (N_13197,N_10593,N_6988);
xnor U13198 (N_13198,N_6952,N_7892);
nor U13199 (N_13199,N_12079,N_12118);
nor U13200 (N_13200,N_7927,N_11575);
or U13201 (N_13201,N_12399,N_8046);
nor U13202 (N_13202,N_6296,N_8973);
xor U13203 (N_13203,N_7882,N_9575);
or U13204 (N_13204,N_9402,N_11062);
xnor U13205 (N_13205,N_12490,N_9155);
and U13206 (N_13206,N_9152,N_7272);
nand U13207 (N_13207,N_7872,N_12438);
xnor U13208 (N_13208,N_9648,N_9486);
and U13209 (N_13209,N_8469,N_11956);
nor U13210 (N_13210,N_7236,N_9125);
nand U13211 (N_13211,N_11888,N_8523);
xnor U13212 (N_13212,N_7099,N_12358);
nor U13213 (N_13213,N_7638,N_10043);
or U13214 (N_13214,N_9237,N_8696);
nor U13215 (N_13215,N_7320,N_11771);
or U13216 (N_13216,N_7589,N_7209);
xor U13217 (N_13217,N_12319,N_7420);
nor U13218 (N_13218,N_6292,N_8497);
nor U13219 (N_13219,N_8992,N_6428);
nand U13220 (N_13220,N_6604,N_8420);
nand U13221 (N_13221,N_8293,N_12186);
xnor U13222 (N_13222,N_7990,N_12481);
xor U13223 (N_13223,N_10722,N_6345);
nand U13224 (N_13224,N_6906,N_11827);
or U13225 (N_13225,N_8296,N_9841);
and U13226 (N_13226,N_12414,N_12444);
xor U13227 (N_13227,N_8838,N_6684);
xor U13228 (N_13228,N_11031,N_6662);
nand U13229 (N_13229,N_6521,N_10788);
nor U13230 (N_13230,N_11067,N_7676);
nor U13231 (N_13231,N_11732,N_9009);
and U13232 (N_13232,N_6935,N_9267);
nor U13233 (N_13233,N_11959,N_8595);
nand U13234 (N_13234,N_10174,N_8960);
nand U13235 (N_13235,N_9414,N_8686);
or U13236 (N_13236,N_9330,N_7398);
or U13237 (N_13237,N_10956,N_7959);
or U13238 (N_13238,N_7721,N_6320);
and U13239 (N_13239,N_8672,N_11979);
xnor U13240 (N_13240,N_6879,N_7467);
nor U13241 (N_13241,N_6502,N_12250);
or U13242 (N_13242,N_9621,N_10476);
nand U13243 (N_13243,N_11767,N_6857);
and U13244 (N_13244,N_10165,N_7164);
nand U13245 (N_13245,N_6812,N_10538);
nand U13246 (N_13246,N_7881,N_9248);
nor U13247 (N_13247,N_9126,N_10896);
nand U13248 (N_13248,N_8611,N_11513);
nor U13249 (N_13249,N_8763,N_9651);
nand U13250 (N_13250,N_6689,N_8089);
nand U13251 (N_13251,N_10994,N_6842);
nor U13252 (N_13252,N_11195,N_11687);
and U13253 (N_13253,N_7308,N_11415);
nand U13254 (N_13254,N_6953,N_9171);
nor U13255 (N_13255,N_6478,N_7703);
and U13256 (N_13256,N_10030,N_8297);
and U13257 (N_13257,N_10216,N_11019);
nor U13258 (N_13258,N_8266,N_8941);
xnor U13259 (N_13259,N_9905,N_8189);
and U13260 (N_13260,N_7136,N_9127);
nor U13261 (N_13261,N_6442,N_11999);
nor U13262 (N_13262,N_10499,N_7938);
nor U13263 (N_13263,N_6930,N_7055);
nor U13264 (N_13264,N_11806,N_10647);
nor U13265 (N_13265,N_12437,N_8948);
nand U13266 (N_13266,N_9912,N_10999);
or U13267 (N_13267,N_7873,N_6339);
xor U13268 (N_13268,N_11526,N_12207);
or U13269 (N_13269,N_11779,N_7133);
nand U13270 (N_13270,N_10140,N_10591);
xor U13271 (N_13271,N_11811,N_9982);
nor U13272 (N_13272,N_6903,N_9926);
or U13273 (N_13273,N_10980,N_11784);
or U13274 (N_13274,N_9059,N_11216);
and U13275 (N_13275,N_11743,N_10406);
or U13276 (N_13276,N_11525,N_7305);
xnor U13277 (N_13277,N_9205,N_9904);
and U13278 (N_13278,N_7311,N_11390);
nor U13279 (N_13279,N_7170,N_9847);
nor U13280 (N_13280,N_9639,N_7201);
nor U13281 (N_13281,N_9160,N_6484);
or U13282 (N_13282,N_8342,N_6357);
nand U13283 (N_13283,N_6691,N_11934);
or U13284 (N_13284,N_7753,N_7975);
xor U13285 (N_13285,N_7915,N_10362);
xor U13286 (N_13286,N_7713,N_7860);
or U13287 (N_13287,N_9116,N_8776);
xor U13288 (N_13288,N_10839,N_9297);
nor U13289 (N_13289,N_10632,N_6547);
and U13290 (N_13290,N_9441,N_12026);
and U13291 (N_13291,N_8839,N_7585);
xnor U13292 (N_13292,N_9655,N_9932);
xnor U13293 (N_13293,N_11680,N_7054);
nor U13294 (N_13294,N_11949,N_11370);
nand U13295 (N_13295,N_8556,N_11906);
nor U13296 (N_13296,N_7490,N_7602);
or U13297 (N_13297,N_11132,N_7355);
nor U13298 (N_13298,N_11976,N_10600);
and U13299 (N_13299,N_6287,N_11692);
and U13300 (N_13300,N_11744,N_8389);
or U13301 (N_13301,N_9526,N_10667);
nand U13302 (N_13302,N_11481,N_6609);
or U13303 (N_13303,N_9708,N_12182);
or U13304 (N_13304,N_7369,N_6269);
nor U13305 (N_13305,N_11210,N_10005);
nor U13306 (N_13306,N_10921,N_8049);
nor U13307 (N_13307,N_6639,N_7972);
and U13308 (N_13308,N_10607,N_6325);
xnor U13309 (N_13309,N_6965,N_8018);
xor U13310 (N_13310,N_9296,N_7466);
or U13311 (N_13311,N_8756,N_10072);
nor U13312 (N_13312,N_12014,N_11419);
nor U13313 (N_13313,N_11458,N_8781);
and U13314 (N_13314,N_8459,N_10385);
nor U13315 (N_13315,N_7091,N_7502);
xor U13316 (N_13316,N_11808,N_9301);
or U13317 (N_13317,N_8620,N_9573);
nor U13318 (N_13318,N_7532,N_6844);
or U13319 (N_13319,N_8883,N_8094);
nor U13320 (N_13320,N_6920,N_8262);
nor U13321 (N_13321,N_7285,N_8479);
nand U13322 (N_13322,N_8474,N_10296);
nand U13323 (N_13323,N_12301,N_7613);
nor U13324 (N_13324,N_12138,N_10107);
xor U13325 (N_13325,N_9615,N_6655);
or U13326 (N_13326,N_11005,N_8201);
or U13327 (N_13327,N_9471,N_6576);
or U13328 (N_13328,N_8863,N_6649);
or U13329 (N_13329,N_12277,N_9887);
xnor U13330 (N_13330,N_9856,N_7002);
or U13331 (N_13331,N_8098,N_7631);
nor U13332 (N_13332,N_10323,N_11844);
or U13333 (N_13333,N_12364,N_7173);
and U13334 (N_13334,N_9558,N_6713);
xnor U13335 (N_13335,N_9384,N_8341);
nor U13336 (N_13336,N_11095,N_9757);
or U13337 (N_13337,N_7898,N_6958);
and U13338 (N_13338,N_11375,N_7106);
xor U13339 (N_13339,N_7778,N_9080);
or U13340 (N_13340,N_8323,N_10447);
or U13341 (N_13341,N_9070,N_6507);
xor U13342 (N_13342,N_12142,N_7666);
nor U13343 (N_13343,N_8429,N_7434);
and U13344 (N_13344,N_11294,N_10497);
nand U13345 (N_13345,N_11333,N_9271);
or U13346 (N_13346,N_7160,N_10166);
nor U13347 (N_13347,N_10241,N_10487);
nand U13348 (N_13348,N_7545,N_10800);
nor U13349 (N_13349,N_7683,N_11021);
xor U13350 (N_13350,N_8573,N_8589);
xor U13351 (N_13351,N_10953,N_7664);
xor U13352 (N_13352,N_6408,N_8843);
xor U13353 (N_13353,N_8114,N_10122);
xnor U13354 (N_13354,N_6278,N_10215);
or U13355 (N_13355,N_12468,N_7088);
nand U13356 (N_13356,N_10131,N_10287);
nor U13357 (N_13357,N_8614,N_8990);
xnor U13358 (N_13358,N_10331,N_8234);
and U13359 (N_13359,N_10096,N_11199);
or U13360 (N_13360,N_6595,N_7999);
and U13361 (N_13361,N_8247,N_7855);
nand U13362 (N_13362,N_11175,N_11441);
or U13363 (N_13363,N_9500,N_11099);
or U13364 (N_13364,N_9739,N_8536);
and U13365 (N_13365,N_7629,N_10698);
xor U13366 (N_13366,N_10682,N_12034);
and U13367 (N_13367,N_10136,N_7996);
nand U13368 (N_13368,N_12148,N_7954);
or U13369 (N_13369,N_9482,N_9900);
or U13370 (N_13370,N_12344,N_11203);
or U13371 (N_13371,N_9032,N_11834);
xor U13372 (N_13372,N_9588,N_6526);
xnor U13373 (N_13373,N_10490,N_10320);
nor U13374 (N_13374,N_6310,N_6892);
xnor U13375 (N_13375,N_7189,N_9594);
nor U13376 (N_13376,N_7616,N_11379);
or U13377 (N_13377,N_6966,N_6850);
and U13378 (N_13378,N_10321,N_8482);
nor U13379 (N_13379,N_12044,N_9410);
nand U13380 (N_13380,N_11353,N_6937);
and U13381 (N_13381,N_7712,N_8962);
nand U13382 (N_13382,N_8915,N_9047);
or U13383 (N_13383,N_11623,N_12227);
and U13384 (N_13384,N_9335,N_6702);
xnor U13385 (N_13385,N_9050,N_6543);
nor U13386 (N_13386,N_9514,N_8285);
nand U13387 (N_13387,N_10143,N_8065);
nor U13388 (N_13388,N_6365,N_7198);
nand U13389 (N_13389,N_7175,N_6690);
and U13390 (N_13390,N_6326,N_7451);
and U13391 (N_13391,N_10608,N_8612);
nor U13392 (N_13392,N_8685,N_8087);
nand U13393 (N_13393,N_6406,N_8603);
nand U13394 (N_13394,N_8946,N_7443);
xnor U13395 (N_13395,N_10185,N_10348);
nand U13396 (N_13396,N_8370,N_9554);
and U13397 (N_13397,N_9849,N_9640);
nand U13398 (N_13398,N_7442,N_12377);
nand U13399 (N_13399,N_6709,N_10100);
xor U13400 (N_13400,N_7251,N_9405);
or U13401 (N_13401,N_7923,N_11241);
nand U13402 (N_13402,N_10851,N_10257);
nor U13403 (N_13403,N_11313,N_8980);
or U13404 (N_13404,N_9709,N_7678);
nor U13405 (N_13405,N_11222,N_10079);
nand U13406 (N_13406,N_10868,N_12463);
xnor U13407 (N_13407,N_6311,N_12196);
xor U13408 (N_13408,N_7257,N_6924);
nor U13409 (N_13409,N_6626,N_7981);
or U13410 (N_13410,N_12108,N_12261);
xnor U13411 (N_13411,N_12293,N_7191);
xor U13412 (N_13412,N_12386,N_11100);
nand U13413 (N_13413,N_11323,N_12011);
nor U13414 (N_13414,N_9234,N_6435);
nand U13415 (N_13415,N_12279,N_6263);
xnor U13416 (N_13416,N_7967,N_12242);
and U13417 (N_13417,N_9316,N_11013);
and U13418 (N_13418,N_10398,N_10726);
xnor U13419 (N_13419,N_9345,N_10314);
nand U13420 (N_13420,N_11478,N_7254);
and U13421 (N_13421,N_6518,N_8190);
nand U13422 (N_13422,N_9147,N_11815);
nand U13423 (N_13423,N_10325,N_11475);
xor U13424 (N_13424,N_11465,N_11372);
and U13425 (N_13425,N_6928,N_10013);
or U13426 (N_13426,N_7592,N_11986);
or U13427 (N_13427,N_6266,N_7510);
nand U13428 (N_13428,N_10205,N_9060);
nand U13429 (N_13429,N_9178,N_11911);
nor U13430 (N_13430,N_11840,N_8373);
nand U13431 (N_13431,N_12120,N_8797);
xnor U13432 (N_13432,N_11051,N_9844);
nand U13433 (N_13433,N_10171,N_12195);
or U13434 (N_13434,N_8576,N_9553);
nand U13435 (N_13435,N_12326,N_6340);
and U13436 (N_13436,N_12190,N_10924);
or U13437 (N_13437,N_8367,N_10509);
or U13438 (N_13438,N_9413,N_11418);
nor U13439 (N_13439,N_11017,N_11144);
nand U13440 (N_13440,N_10288,N_7922);
or U13441 (N_13441,N_6261,N_7461);
nand U13442 (N_13442,N_10913,N_9314);
nor U13443 (N_13443,N_12278,N_7162);
and U13444 (N_13444,N_8967,N_10648);
or U13445 (N_13445,N_11034,N_6352);
xor U13446 (N_13446,N_12380,N_12170);
xnor U13447 (N_13447,N_9504,N_12333);
or U13448 (N_13448,N_8238,N_7458);
nor U13449 (N_13449,N_7031,N_9863);
nor U13450 (N_13450,N_7793,N_10714);
or U13451 (N_13451,N_10281,N_6555);
or U13452 (N_13452,N_12327,N_7018);
nor U13453 (N_13453,N_8500,N_8662);
and U13454 (N_13454,N_10471,N_8384);
and U13455 (N_13455,N_12405,N_6392);
or U13456 (N_13456,N_12471,N_10411);
nor U13457 (N_13457,N_10633,N_11508);
nand U13458 (N_13458,N_6536,N_12443);
nor U13459 (N_13459,N_9768,N_9801);
and U13460 (N_13460,N_8625,N_7652);
nor U13461 (N_13461,N_6898,N_10762);
and U13462 (N_13462,N_7043,N_10265);
nand U13463 (N_13463,N_11787,N_10052);
nor U13464 (N_13464,N_12410,N_12016);
nand U13465 (N_13465,N_9246,N_9168);
xnor U13466 (N_13466,N_7220,N_8740);
nand U13467 (N_13467,N_11537,N_8440);
nand U13468 (N_13468,N_10097,N_10875);
nand U13469 (N_13469,N_6376,N_12495);
or U13470 (N_13470,N_7500,N_11781);
xnor U13471 (N_13471,N_7704,N_8180);
and U13472 (N_13472,N_6793,N_8154);
and U13473 (N_13473,N_10041,N_10860);
or U13474 (N_13474,N_8375,N_8033);
or U13475 (N_13475,N_7896,N_8443);
xor U13476 (N_13476,N_10802,N_12469);
and U13477 (N_13477,N_8220,N_11867);
xnor U13478 (N_13478,N_12031,N_12122);
and U13479 (N_13479,N_10120,N_9817);
nand U13480 (N_13480,N_11301,N_9633);
xnor U13481 (N_13481,N_10450,N_7542);
nand U13482 (N_13482,N_6968,N_7010);
nand U13483 (N_13483,N_11197,N_10713);
nor U13484 (N_13484,N_12097,N_9182);
xor U13485 (N_13485,N_7657,N_11489);
nor U13486 (N_13486,N_7832,N_8993);
or U13487 (N_13487,N_8439,N_9022);
and U13488 (N_13488,N_11614,N_11595);
xor U13489 (N_13489,N_8836,N_9516);
or U13490 (N_13490,N_8058,N_6789);
xnor U13491 (N_13491,N_10888,N_7471);
and U13492 (N_13492,N_8076,N_12193);
xnor U13493 (N_13493,N_6939,N_7786);
or U13494 (N_13494,N_7141,N_11046);
nand U13495 (N_13495,N_6819,N_8931);
or U13496 (N_13496,N_10235,N_11001);
and U13497 (N_13497,N_8136,N_11930);
xnor U13498 (N_13498,N_9356,N_8842);
xor U13499 (N_13499,N_7199,N_7127);
nand U13500 (N_13500,N_8382,N_7960);
nor U13501 (N_13501,N_6794,N_10665);
nand U13502 (N_13502,N_10498,N_7687);
xnor U13503 (N_13503,N_8552,N_8075);
nand U13504 (N_13504,N_12100,N_6260);
xor U13505 (N_13505,N_9707,N_7419);
nor U13506 (N_13506,N_6387,N_8100);
or U13507 (N_13507,N_11529,N_10091);
and U13508 (N_13508,N_12045,N_7989);
or U13509 (N_13509,N_9395,N_10439);
nor U13510 (N_13510,N_10401,N_9680);
nand U13511 (N_13511,N_10489,N_7326);
nand U13512 (N_13512,N_7258,N_8257);
or U13513 (N_13513,N_9363,N_11541);
nor U13514 (N_13514,N_11286,N_9225);
xor U13515 (N_13515,N_12331,N_9091);
xnor U13516 (N_13516,N_8704,N_6860);
nand U13517 (N_13517,N_10798,N_7124);
xnor U13518 (N_13518,N_10583,N_12172);
nor U13519 (N_13519,N_8345,N_10857);
nor U13520 (N_13520,N_11373,N_10340);
nor U13521 (N_13521,N_10108,N_6868);
nand U13522 (N_13522,N_8404,N_11421);
and U13523 (N_13523,N_10634,N_11962);
xnor U13524 (N_13524,N_11092,N_7069);
or U13525 (N_13525,N_8158,N_7457);
nand U13526 (N_13526,N_9753,N_9744);
xnor U13527 (N_13527,N_8584,N_9002);
and U13528 (N_13528,N_11901,N_6385);
and U13529 (N_13529,N_7618,N_11564);
nand U13530 (N_13530,N_6382,N_9362);
nor U13531 (N_13531,N_9883,N_7850);
or U13532 (N_13532,N_9051,N_8379);
nor U13533 (N_13533,N_9398,N_9309);
xor U13534 (N_13534,N_12131,N_6910);
nor U13535 (N_13535,N_6707,N_6319);
xor U13536 (N_13536,N_10025,N_7045);
and U13537 (N_13537,N_7300,N_11796);
xor U13538 (N_13538,N_7574,N_9892);
nand U13539 (N_13539,N_8877,N_7557);
and U13540 (N_13540,N_10429,N_11832);
nand U13541 (N_13541,N_6855,N_10115);
and U13542 (N_13542,N_11242,N_9305);
and U13543 (N_13543,N_6686,N_10615);
or U13544 (N_13544,N_10225,N_9037);
nor U13545 (N_13545,N_10720,N_10522);
xnor U13546 (N_13546,N_7551,N_11027);
xor U13547 (N_13547,N_10180,N_10709);
and U13548 (N_13548,N_8478,N_12477);
nand U13549 (N_13549,N_10679,N_9386);
xnor U13550 (N_13550,N_11445,N_7137);
nand U13551 (N_13551,N_11984,N_8391);
and U13552 (N_13552,N_10283,N_12135);
xnor U13553 (N_13553,N_10938,N_9548);
or U13554 (N_13554,N_7255,N_9401);
and U13555 (N_13555,N_6977,N_7582);
and U13556 (N_13556,N_8806,N_7159);
nor U13557 (N_13557,N_12156,N_6495);
or U13558 (N_13558,N_8338,N_6768);
or U13559 (N_13559,N_9033,N_6550);
nor U13560 (N_13560,N_10155,N_7454);
nand U13561 (N_13561,N_6298,N_10028);
nor U13562 (N_13562,N_10505,N_8558);
nand U13563 (N_13563,N_8118,N_10606);
nand U13564 (N_13564,N_6438,N_10721);
nor U13565 (N_13565,N_11872,N_8119);
and U13566 (N_13566,N_9187,N_12199);
xnor U13567 (N_13567,N_8771,N_10470);
nand U13568 (N_13568,N_9136,N_7324);
and U13569 (N_13569,N_8277,N_9284);
nand U13570 (N_13570,N_10978,N_9081);
or U13571 (N_13571,N_12161,N_12248);
and U13572 (N_13572,N_10576,N_12208);
nor U13573 (N_13573,N_11997,N_11612);
and U13574 (N_13574,N_11764,N_10239);
xnor U13575 (N_13575,N_6747,N_7230);
nand U13576 (N_13576,N_11955,N_9250);
or U13577 (N_13577,N_8216,N_7347);
or U13578 (N_13578,N_7378,N_11626);
nor U13579 (N_13579,N_8346,N_7849);
or U13580 (N_13580,N_10313,N_9625);
nor U13581 (N_13581,N_11025,N_11399);
nor U13582 (N_13582,N_12260,N_8991);
nor U13583 (N_13583,N_8372,N_7564);
xor U13584 (N_13584,N_11517,N_6971);
or U13585 (N_13585,N_11603,N_8994);
xor U13586 (N_13586,N_10663,N_6916);
nor U13587 (N_13587,N_10880,N_11243);
nand U13588 (N_13588,N_12078,N_7747);
or U13589 (N_13589,N_8749,N_7887);
nand U13590 (N_13590,N_8718,N_9517);
xor U13591 (N_13591,N_7115,N_7911);
xnor U13592 (N_13592,N_9701,N_11431);
and U13593 (N_13593,N_11702,N_9657);
nor U13594 (N_13594,N_11681,N_8203);
or U13595 (N_13595,N_6460,N_12365);
xor U13596 (N_13596,N_9922,N_11735);
nor U13597 (N_13597,N_6981,N_10660);
nand U13598 (N_13598,N_9438,N_9896);
nor U13599 (N_13599,N_7862,N_11068);
nor U13600 (N_13600,N_10942,N_11693);
and U13601 (N_13601,N_7195,N_11499);
xor U13602 (N_13602,N_7269,N_11096);
nor U13603 (N_13603,N_10209,N_9142);
or U13604 (N_13604,N_12145,N_8147);
or U13605 (N_13605,N_8947,N_11217);
xnor U13606 (N_13606,N_6482,N_7415);
nand U13607 (N_13607,N_11675,N_12281);
and U13608 (N_13608,N_7740,N_8896);
or U13609 (N_13609,N_9731,N_11857);
nor U13610 (N_13610,N_6492,N_7580);
and U13611 (N_13611,N_10333,N_11272);
nor U13612 (N_13612,N_11330,N_7125);
or U13613 (N_13613,N_6788,N_6663);
or U13614 (N_13614,N_8037,N_6742);
and U13615 (N_13615,N_7744,N_10464);
nor U13616 (N_13616,N_7432,N_10324);
or U13617 (N_13617,N_9396,N_12334);
and U13618 (N_13618,N_6746,N_6629);
and U13619 (N_13619,N_8422,N_11039);
xor U13620 (N_13620,N_7603,N_6347);
nor U13621 (N_13621,N_8123,N_7178);
xor U13622 (N_13622,N_10511,N_6413);
nor U13623 (N_13623,N_10507,N_11460);
nand U13624 (N_13624,N_10664,N_9877);
or U13625 (N_13625,N_11533,N_8164);
and U13626 (N_13626,N_11824,N_12134);
nor U13627 (N_13627,N_9952,N_11581);
or U13628 (N_13628,N_8857,N_7182);
and U13629 (N_13629,N_12389,N_6668);
nor U13630 (N_13630,N_7857,N_9845);
or U13631 (N_13631,N_6731,N_6608);
nand U13632 (N_13632,N_7297,N_10892);
xnor U13633 (N_13633,N_8528,N_9860);
xnor U13634 (N_13634,N_11583,N_9465);
nor U13635 (N_13635,N_9888,N_9149);
xnor U13636 (N_13636,N_7484,N_7452);
nor U13637 (N_13637,N_10653,N_11574);
and U13638 (N_13638,N_10169,N_11366);
or U13639 (N_13639,N_8408,N_10022);
or U13640 (N_13640,N_12052,N_11608);
or U13641 (N_13641,N_11989,N_8047);
nor U13642 (N_13642,N_6616,N_11251);
nand U13643 (N_13643,N_9750,N_8504);
xnor U13644 (N_13644,N_10812,N_7591);
or U13645 (N_13645,N_9415,N_7130);
nor U13646 (N_13646,N_6470,N_10526);
xnor U13647 (N_13647,N_12266,N_7070);
nand U13648 (N_13648,N_9268,N_7112);
or U13649 (N_13649,N_9420,N_9198);
or U13650 (N_13650,N_7341,N_9057);
nor U13651 (N_13651,N_7225,N_12050);
nor U13652 (N_13652,N_7547,N_12060);
nor U13653 (N_13653,N_8661,N_9282);
and U13654 (N_13654,N_8935,N_8335);
and U13655 (N_13655,N_11334,N_9828);
and U13656 (N_13656,N_11657,N_11963);
nor U13657 (N_13657,N_10889,N_6726);
xnor U13658 (N_13658,N_8029,N_8621);
nand U13659 (N_13659,N_10393,N_10561);
and U13660 (N_13660,N_11876,N_7800);
and U13661 (N_13661,N_7634,N_10415);
nor U13662 (N_13662,N_10078,N_8570);
or U13663 (N_13663,N_10843,N_10266);
xor U13664 (N_13664,N_7410,N_8256);
nand U13665 (N_13665,N_8531,N_10803);
or U13666 (N_13666,N_12385,N_7976);
xor U13667 (N_13667,N_9976,N_9021);
xnor U13668 (N_13668,N_9656,N_7594);
and U13669 (N_13669,N_6718,N_9595);
xnor U13670 (N_13670,N_7318,N_8898);
or U13671 (N_13671,N_6315,N_9195);
xor U13672 (N_13672,N_9166,N_6600);
nor U13673 (N_13673,N_7192,N_10794);
nand U13674 (N_13674,N_9315,N_8363);
nand U13675 (N_13675,N_8817,N_9202);
nor U13676 (N_13676,N_9634,N_8940);
nand U13677 (N_13677,N_7119,N_11211);
xor U13678 (N_13678,N_9889,N_7211);
nand U13679 (N_13679,N_10304,N_10019);
xor U13680 (N_13680,N_12442,N_8807);
nand U13681 (N_13681,N_9031,N_11213);
or U13682 (N_13682,N_6862,N_7956);
xnor U13683 (N_13683,N_9106,N_8581);
and U13684 (N_13684,N_11036,N_11733);
nand U13685 (N_13685,N_10455,N_9762);
or U13686 (N_13686,N_8850,N_8753);
nand U13687 (N_13687,N_7840,N_9186);
and U13688 (N_13688,N_8083,N_10589);
and U13689 (N_13689,N_8997,N_11463);
and U13690 (N_13690,N_6449,N_10883);
nand U13691 (N_13691,N_8070,N_11162);
nand U13692 (N_13692,N_10148,N_10925);
nand U13693 (N_13693,N_12307,N_9789);
xor U13694 (N_13694,N_7262,N_11176);
nand U13695 (N_13695,N_6530,N_10138);
or U13696 (N_13696,N_8630,N_8972);
and U13697 (N_13697,N_8461,N_8462);
xor U13698 (N_13698,N_10486,N_6433);
or U13699 (N_13699,N_10104,N_9107);
nand U13700 (N_13700,N_10158,N_11150);
nand U13701 (N_13701,N_9767,N_9319);
and U13702 (N_13702,N_10350,N_8631);
and U13703 (N_13703,N_6524,N_7710);
nor U13704 (N_13704,N_7132,N_11401);
and U13705 (N_13705,N_10000,N_10077);
or U13706 (N_13706,N_10110,N_10742);
and U13707 (N_13707,N_8001,N_8396);
xor U13708 (N_13708,N_11009,N_11278);
nand U13709 (N_13709,N_9853,N_7885);
and U13710 (N_13710,N_11185,N_11716);
nand U13711 (N_13711,N_9846,N_12192);
and U13712 (N_13712,N_12321,N_8908);
nor U13713 (N_13713,N_10736,N_7486);
and U13714 (N_13714,N_12009,N_7813);
xnor U13715 (N_13715,N_6700,N_8279);
and U13716 (N_13716,N_10347,N_11026);
or U13717 (N_13717,N_9385,N_8019);
xor U13718 (N_13718,N_12188,N_9130);
or U13719 (N_13719,N_6286,N_6450);
nor U13720 (N_13720,N_12270,N_8689);
nor U13721 (N_13721,N_7408,N_10605);
or U13722 (N_13722,N_11268,N_8275);
or U13723 (N_13723,N_8551,N_10772);
or U13724 (N_13724,N_7041,N_12010);
nand U13725 (N_13725,N_10388,N_11193);
or U13726 (N_13726,N_8522,N_9626);
nand U13727 (N_13727,N_11543,N_7886);
or U13728 (N_13728,N_11770,N_10586);
nor U13729 (N_13729,N_10031,N_6329);
xor U13730 (N_13730,N_6687,N_11337);
xnor U13731 (N_13731,N_8568,N_12022);
nand U13732 (N_13732,N_11799,N_8172);
nand U13733 (N_13733,N_11887,N_10706);
nand U13734 (N_13734,N_9812,N_9991);
or U13735 (N_13735,N_6488,N_6349);
xor U13736 (N_13736,N_6856,N_7876);
xnor U13737 (N_13737,N_9443,N_7469);
xor U13738 (N_13738,N_7733,N_6638);
and U13739 (N_13739,N_9764,N_8913);
nand U13740 (N_13740,N_8223,N_7234);
and U13741 (N_13741,N_11466,N_9244);
or U13742 (N_13742,N_10374,N_8916);
nand U13743 (N_13743,N_10261,N_7949);
or U13744 (N_13744,N_7743,N_9807);
xor U13745 (N_13745,N_7948,N_12271);
xnor U13746 (N_13746,N_10823,N_11831);
nand U13747 (N_13747,N_8895,N_9539);
xor U13748 (N_13748,N_9346,N_9561);
or U13749 (N_13749,N_8879,N_6989);
and U13750 (N_13750,N_8575,N_7422);
nand U13751 (N_13751,N_10217,N_6610);
or U13752 (N_13752,N_10229,N_9466);
nor U13753 (N_13753,N_11456,N_8224);
xor U13754 (N_13754,N_10760,N_10791);
and U13755 (N_13755,N_7978,N_7858);
nand U13756 (N_13756,N_8304,N_8191);
xnor U13757 (N_13757,N_8562,N_11288);
or U13758 (N_13758,N_12407,N_11003);
or U13759 (N_13759,N_10817,N_6889);
nor U13760 (N_13760,N_10572,N_8369);
or U13761 (N_13761,N_6990,N_6498);
xor U13762 (N_13762,N_6800,N_10201);
nor U13763 (N_13763,N_10971,N_9958);
nand U13764 (N_13764,N_10741,N_10423);
and U13765 (N_13765,N_7128,N_8903);
and U13766 (N_13766,N_7569,N_6350);
and U13767 (N_13767,N_9487,N_7260);
nand U13768 (N_13768,N_6736,N_7780);
xor U13769 (N_13769,N_7015,N_9947);
and U13770 (N_13770,N_11192,N_8281);
nor U13771 (N_13771,N_10207,N_9662);
nand U13772 (N_13772,N_9424,N_10017);
nand U13773 (N_13773,N_9369,N_8812);
or U13774 (N_13774,N_12215,N_6625);
and U13775 (N_13775,N_9501,N_8687);
nor U13776 (N_13776,N_7362,N_11467);
and U13777 (N_13777,N_11240,N_7979);
and U13778 (N_13778,N_10517,N_9392);
nand U13779 (N_13779,N_8134,N_11721);
nor U13780 (N_13780,N_6445,N_11924);
and U13781 (N_13781,N_6730,N_11315);
xor U13782 (N_13782,N_11648,N_11654);
nand U13783 (N_13783,N_12289,N_12339);
nand U13784 (N_13784,N_6795,N_10293);
xor U13785 (N_13785,N_9359,N_9348);
and U13786 (N_13786,N_9642,N_8057);
xor U13787 (N_13787,N_12205,N_8841);
nand U13788 (N_13788,N_11507,N_11883);
nor U13789 (N_13789,N_6424,N_11794);
xnor U13790 (N_13790,N_12366,N_9878);
and U13791 (N_13791,N_8825,N_8143);
or U13792 (N_13792,N_11542,N_12234);
xnor U13793 (N_13793,N_8193,N_10006);
or U13794 (N_13794,N_10636,N_7897);
and U13795 (N_13795,N_8961,N_11253);
xor U13796 (N_13796,N_11841,N_8388);
nor U13797 (N_13797,N_11273,N_10680);
xnor U13798 (N_13798,N_8905,N_11711);
and U13799 (N_13799,N_7036,N_12264);
nand U13800 (N_13800,N_12313,N_10690);
or U13801 (N_13801,N_7931,N_9913);
xnor U13802 (N_13802,N_10582,N_7232);
nor U13803 (N_13803,N_8259,N_10809);
and U13804 (N_13804,N_8039,N_6926);
and U13805 (N_13805,N_9696,N_6596);
nand U13806 (N_13806,N_12268,N_12341);
or U13807 (N_13807,N_7980,N_12263);
and U13808 (N_13808,N_6453,N_9439);
nand U13809 (N_13809,N_12367,N_7659);
nand U13810 (N_13810,N_8642,N_9435);
or U13811 (N_13811,N_7117,N_11016);
or U13812 (N_13812,N_12290,N_9963);
nor U13813 (N_13813,N_6936,N_8487);
nor U13814 (N_13814,N_8869,N_7537);
xnor U13815 (N_13815,N_6888,N_9676);
nand U13816 (N_13816,N_9949,N_10472);
nand U13817 (N_13817,N_10790,N_10629);
nor U13818 (N_13818,N_11822,N_11226);
nand U13819 (N_13819,N_6778,N_6476);
or U13820 (N_13820,N_12472,N_11454);
nand U13821 (N_13821,N_11593,N_12103);
xor U13822 (N_13822,N_11355,N_11350);
nor U13823 (N_13823,N_9200,N_7418);
nor U13824 (N_13824,N_7933,N_6436);
nor U13825 (N_13825,N_9827,N_10232);
nor U13826 (N_13826,N_8470,N_8892);
or U13827 (N_13827,N_8326,N_7438);
nor U13828 (N_13828,N_9620,N_8996);
and U13829 (N_13829,N_8712,N_8208);
xnor U13830 (N_13830,N_7080,N_10708);
nor U13831 (N_13831,N_8110,N_10666);
xnor U13832 (N_13832,N_8125,N_7437);
and U13833 (N_13833,N_6636,N_9476);
nor U13834 (N_13834,N_12465,N_6591);
nor U13835 (N_13835,N_11363,N_8101);
nor U13836 (N_13836,N_6412,N_8454);
nor U13837 (N_13837,N_7961,N_9751);
nand U13838 (N_13838,N_10766,N_11429);
and U13839 (N_13839,N_6590,N_7073);
and U13840 (N_13840,N_6579,N_11966);
or U13841 (N_13841,N_8899,N_6872);
xnor U13842 (N_13842,N_9207,N_11661);
xnor U13843 (N_13843,N_6425,N_10050);
xor U13844 (N_13844,N_7998,N_10349);
nand U13845 (N_13845,N_11741,N_9944);
or U13846 (N_13846,N_7965,N_12096);
nor U13847 (N_13847,N_11503,N_10029);
nor U13848 (N_13848,N_9530,N_6391);
nand U13849 (N_13849,N_11317,N_8427);
xnor U13850 (N_13850,N_8739,N_10087);
and U13851 (N_13851,N_8561,N_7940);
nand U13852 (N_13852,N_11408,N_9663);
and U13853 (N_13853,N_8051,N_10644);
xnor U13854 (N_13854,N_11679,N_11228);
nor U13855 (N_13855,N_7370,N_9566);
and U13856 (N_13856,N_12485,N_8209);
nand U13857 (N_13857,N_7610,N_9474);
and U13858 (N_13858,N_11167,N_11339);
nor U13859 (N_13859,N_8729,N_6694);
nor U13860 (N_13860,N_10740,N_10932);
nand U13861 (N_13861,N_8414,N_8267);
and U13862 (N_13862,N_9417,N_7395);
and U13863 (N_13863,N_9461,N_6740);
nor U13864 (N_13864,N_12209,N_10189);
nor U13865 (N_13865,N_7224,N_8748);
and U13866 (N_13866,N_11158,N_7755);
and U13867 (N_13867,N_12311,N_10199);
and U13868 (N_13868,N_6880,N_12081);
nand U13869 (N_13869,N_8061,N_12077);
nor U13870 (N_13870,N_11077,N_11238);
nand U13871 (N_13871,N_12393,N_9193);
nand U13872 (N_13872,N_6582,N_10806);
or U13873 (N_13873,N_10055,N_12494);
and U13874 (N_13874,N_9791,N_11609);
nand U13875 (N_13875,N_10816,N_9444);
and U13876 (N_13876,N_9995,N_10531);
nand U13877 (N_13877,N_8891,N_7774);
or U13878 (N_13878,N_10618,N_9506);
and U13879 (N_13879,N_10219,N_6611);
xor U13880 (N_13880,N_11189,N_12460);
and U13881 (N_13881,N_9858,N_12224);
and U13882 (N_13882,N_8752,N_11265);
and U13883 (N_13883,N_8005,N_6399);
xnor U13884 (N_13884,N_9540,N_10255);
nand U13885 (N_13885,N_6979,N_12219);
nor U13886 (N_13886,N_8311,N_12383);
xnor U13887 (N_13887,N_11907,N_10193);
xnor U13888 (N_13888,N_6961,N_6732);
or U13889 (N_13889,N_11701,N_9940);
or U13890 (N_13890,N_11584,N_11990);
nor U13891 (N_13891,N_6472,N_11302);
and U13892 (N_13892,N_6938,N_10410);
or U13893 (N_13893,N_12104,N_8142);
nand U13894 (N_13894,N_7846,N_8691);
nand U13895 (N_13895,N_7827,N_6299);
nor U13896 (N_13896,N_7756,N_8515);
or U13897 (N_13897,N_8121,N_6805);
nor U13898 (N_13898,N_12448,N_10911);
and U13899 (N_13899,N_6627,N_8398);
nor U13900 (N_13900,N_7016,N_11407);
xor U13901 (N_13901,N_10457,N_9434);
and U13902 (N_13902,N_10789,N_9472);
and U13903 (N_13903,N_6631,N_11066);
or U13904 (N_13904,N_12322,N_10967);
xnor U13905 (N_13905,N_8699,N_8273);
and U13906 (N_13906,N_7473,N_7528);
nor U13907 (N_13907,N_10757,N_6462);
or U13908 (N_13908,N_8442,N_7226);
or U13909 (N_13909,N_7805,N_6519);
nand U13910 (N_13910,N_7030,N_12274);
xnor U13911 (N_13911,N_11365,N_9341);
nand U13912 (N_13912,N_10547,N_11396);
nor U13913 (N_13913,N_8900,N_7331);
nor U13914 (N_13914,N_8984,N_11108);
nand U13915 (N_13915,N_8132,N_7172);
or U13916 (N_13916,N_10524,N_8361);
nand U13917 (N_13917,N_9531,N_9650);
and U13918 (N_13918,N_8532,N_9647);
nor U13919 (N_13919,N_12166,N_12445);
and U13920 (N_13920,N_7636,N_10156);
and U13921 (N_13921,N_11319,N_9819);
nand U13922 (N_13922,N_8651,N_11097);
xor U13923 (N_13923,N_7794,N_12046);
xnor U13924 (N_13924,N_10343,N_10628);
nand U13925 (N_13925,N_9264,N_9678);
xor U13926 (N_13926,N_9603,N_6908);
xor U13927 (N_13927,N_11451,N_11050);
nor U13928 (N_13928,N_11758,N_10071);
or U13929 (N_13929,N_12305,N_10141);
xnor U13930 (N_13930,N_6494,N_12194);
and U13931 (N_13931,N_10309,N_8221);
nor U13932 (N_13932,N_9243,N_9627);
nand U13933 (N_13933,N_7751,N_12041);
and U13934 (N_13934,N_6792,N_10824);
or U13935 (N_13935,N_6363,N_7932);
nand U13936 (N_13936,N_6467,N_6619);
nand U13937 (N_13937,N_9724,N_10298);
xor U13938 (N_13938,N_11329,N_10867);
xor U13939 (N_13939,N_7785,N_11378);
xor U13940 (N_13940,N_9614,N_7507);
and U13941 (N_13941,N_8230,N_9513);
xor U13942 (N_13942,N_10604,N_6553);
xnor U13943 (N_13943,N_9884,N_7597);
or U13944 (N_13944,N_10554,N_11357);
nand U13945 (N_13945,N_12160,N_11665);
xor U13946 (N_13946,N_8305,N_6927);
or U13947 (N_13947,N_8378,N_9903);
and U13948 (N_13948,N_11405,N_6864);
or U13949 (N_13949,N_9431,N_7241);
nor U13950 (N_13950,N_6336,N_12173);
or U13951 (N_13951,N_11670,N_8042);
nand U13952 (N_13952,N_7468,N_8280);
xor U13953 (N_13953,N_12302,N_10056);
and U13954 (N_13954,N_6430,N_9072);
nor U13955 (N_13955,N_8745,N_9765);
and U13956 (N_13956,N_7802,N_9240);
or U13957 (N_13957,N_10124,N_10035);
or U13958 (N_13958,N_11947,N_10724);
nand U13959 (N_13959,N_11601,N_6531);
nor U13960 (N_13960,N_8405,N_9685);
xnor U13961 (N_13961,N_8785,N_12243);
nor U13962 (N_13962,N_9016,N_6309);
nand U13963 (N_13963,N_10163,N_7716);
xnor U13964 (N_13964,N_11316,N_7040);
nand U13965 (N_13965,N_7847,N_12343);
and U13966 (N_13966,N_9718,N_8090);
xor U13967 (N_13967,N_8165,N_7062);
xor U13968 (N_13968,N_12296,N_6929);
xnor U13969 (N_13969,N_9524,N_9491);
or U13970 (N_13970,N_6666,N_7779);
or U13971 (N_13971,N_10109,N_10745);
nor U13972 (N_13972,N_11640,N_6791);
xor U13973 (N_13973,N_7103,N_8348);
or U13974 (N_13974,N_6834,N_11112);
nor U13975 (N_13975,N_12286,N_9725);
nand U13976 (N_13976,N_7587,N_9242);
and U13977 (N_13977,N_10172,N_10246);
nand U13978 (N_13978,N_8728,N_7942);
or U13979 (N_13979,N_7086,N_12210);
nor U13980 (N_13980,N_9074,N_10409);
and U13981 (N_13981,N_8272,N_7833);
or U13982 (N_13982,N_7605,N_7731);
nor U13983 (N_13983,N_11427,N_10434);
or U13984 (N_13984,N_7000,N_10715);
nand U13985 (N_13985,N_9083,N_6720);
and U13986 (N_13986,N_7063,N_11208);
or U13987 (N_13987,N_9035,N_11678);
nand U13988 (N_13988,N_10918,N_12091);
nor U13989 (N_13989,N_6911,N_10569);
and U13990 (N_13990,N_7348,N_10596);
or U13991 (N_13991,N_9429,N_9493);
or U13992 (N_13992,N_12422,N_9110);
nand U13993 (N_13993,N_11120,N_8671);
nor U13994 (N_13994,N_10639,N_12351);
or U13995 (N_13995,N_11049,N_11109);
xnor U13996 (N_13996,N_8162,N_7566);
nand U13997 (N_13997,N_10856,N_7807);
or U13998 (N_13998,N_9542,N_10862);
or U13999 (N_13999,N_6955,N_12423);
and U14000 (N_14000,N_8588,N_6409);
or U14001 (N_14001,N_8217,N_9212);
and U14002 (N_14002,N_11083,N_10981);
and U14003 (N_14003,N_10196,N_9477);
xnor U14004 (N_14004,N_6847,N_9382);
and U14005 (N_14005,N_11858,N_7578);
nor U14006 (N_14006,N_10413,N_12241);
nor U14007 (N_14007,N_6516,N_11531);
nor U14008 (N_14008,N_7766,N_11300);
and U14009 (N_14009,N_7433,N_7934);
nand U14010 (N_14010,N_11782,N_11917);
and U14011 (N_14011,N_11080,N_8742);
nor U14012 (N_14012,N_11705,N_10188);
nor U14013 (N_14013,N_7883,N_9960);
nor U14014 (N_14014,N_10269,N_11220);
nor U14015 (N_14015,N_6950,N_9653);
nand U14016 (N_14016,N_8918,N_6845);
xnor U14017 (N_14017,N_9082,N_8598);
or U14018 (N_14018,N_10012,N_7093);
and U14019 (N_14019,N_10876,N_11033);
xor U14020 (N_14020,N_9979,N_8403);
nand U14021 (N_14021,N_12150,N_8862);
or U14022 (N_14022,N_8186,N_6758);
nor U14023 (N_14023,N_7120,N_9978);
nor U14024 (N_14024,N_8754,N_6914);
and U14025 (N_14025,N_7238,N_10884);
nor U14026 (N_14026,N_8291,N_10598);
nand U14027 (N_14027,N_8211,N_7706);
xnor U14028 (N_14028,N_8481,N_7856);
nand U14029 (N_14029,N_10542,N_10383);
nor U14030 (N_14030,N_10151,N_8791);
nand U14031 (N_14031,N_8583,N_8024);
or U14032 (N_14032,N_11958,N_6809);
xor U14033 (N_14033,N_9914,N_6342);
and U14034 (N_14034,N_8228,N_11842);
and U14035 (N_14035,N_9775,N_8318);
nand U14036 (N_14036,N_9933,N_10904);
xnor U14037 (N_14037,N_12473,N_10581);
nand U14038 (N_14038,N_10099,N_8292);
nand U14039 (N_14039,N_7985,N_10276);
xnor U14040 (N_14040,N_11131,N_11263);
and U14041 (N_14041,N_8269,N_9304);
or U14042 (N_14042,N_11170,N_6404);
or U14043 (N_14043,N_9972,N_8591);
nand U14044 (N_14044,N_6335,N_10477);
nand U14045 (N_14045,N_9045,N_11110);
and U14046 (N_14046,N_10226,N_9915);
xor U14047 (N_14047,N_9818,N_9917);
xnor U14048 (N_14048,N_10546,N_8665);
nor U14049 (N_14049,N_11856,N_10446);
and U14050 (N_14050,N_11659,N_11545);
or U14051 (N_14051,N_11362,N_7562);
nor U14052 (N_14052,N_10094,N_7604);
nor U14053 (N_14053,N_6313,N_12441);
nand U14054 (N_14054,N_8484,N_10894);
nor U14055 (N_14055,N_10334,N_6770);
and U14056 (N_14056,N_12310,N_9745);
nor U14057 (N_14057,N_10396,N_8084);
nand U14058 (N_14058,N_6471,N_10046);
and U14059 (N_14059,N_10539,N_9419);
nor U14060 (N_14060,N_12165,N_7491);
nand U14061 (N_14061,N_8499,N_10502);
and U14062 (N_14062,N_10516,N_11691);
nor U14063 (N_14063,N_9391,N_9916);
or U14064 (N_14064,N_9968,N_7188);
and U14065 (N_14065,N_7944,N_9602);
or U14066 (N_14066,N_11890,N_7424);
or U14067 (N_14067,N_9020,N_7026);
or U14068 (N_14068,N_10521,N_6695);
or U14069 (N_14069,N_11328,N_10731);
or U14070 (N_14070,N_8066,N_11184);
or U14071 (N_14071,N_6457,N_8232);
nand U14072 (N_14072,N_9265,N_8808);
nand U14073 (N_14073,N_10964,N_10186);
or U14074 (N_14074,N_10488,N_8743);
nor U14075 (N_14075,N_8928,N_10734);
or U14076 (N_14076,N_8392,N_7763);
nand U14077 (N_14077,N_12093,N_12201);
xor U14078 (N_14078,N_6728,N_11809);
and U14079 (N_14079,N_6253,N_10672);
and U14080 (N_14080,N_10959,N_12128);
xnor U14081 (N_14081,N_6940,N_11159);
nor U14082 (N_14082,N_6571,N_8540);
or U14083 (N_14083,N_12019,N_6771);
nor U14084 (N_14084,N_10801,N_8329);
and U14085 (N_14085,N_11340,N_10960);
nor U14086 (N_14086,N_12036,N_6259);
nor U14087 (N_14087,N_11672,N_7479);
or U14088 (N_14088,N_12464,N_10686);
and U14089 (N_14089,N_8880,N_9842);
and U14090 (N_14090,N_11433,N_8249);
or U14091 (N_14091,N_10206,N_8851);
or U14092 (N_14092,N_10947,N_11853);
or U14093 (N_14093,N_7790,N_9280);
and U14094 (N_14094,N_6830,N_9312);
or U14095 (N_14095,N_8214,N_8206);
nor U14096 (N_14096,N_9442,N_10786);
nand U14097 (N_14097,N_9379,N_10060);
nand U14098 (N_14098,N_10887,N_9067);
xor U14099 (N_14099,N_11424,N_6841);
nor U14100 (N_14100,N_7480,N_10638);
nor U14101 (N_14101,N_9692,N_8188);
nor U14102 (N_14102,N_9999,N_8246);
and U14103 (N_14103,N_7741,N_6705);
nand U14104 (N_14104,N_8968,N_10958);
or U14105 (N_14105,N_7995,N_11103);
xor U14106 (N_14106,N_10262,N_6996);
xor U14107 (N_14107,N_8802,N_6272);
and U14108 (N_14108,N_11801,N_9322);
xnor U14109 (N_14109,N_12496,N_6587);
xor U14110 (N_14110,N_8951,N_11642);
nand U14111 (N_14111,N_7244,N_12155);
xor U14112 (N_14112,N_7769,N_6782);
nor U14113 (N_14113,N_9886,N_10838);
nand U14114 (N_14114,N_12450,N_10768);
or U14115 (N_14115,N_8124,N_11650);
xor U14116 (N_14116,N_10212,N_7100);
and U14117 (N_14117,N_7056,N_11579);
nand U14118 (N_14118,N_10927,N_6960);
or U14119 (N_14119,N_10631,N_7145);
nand U14120 (N_14120,N_11558,N_7702);
nor U14121 (N_14121,N_9144,N_12324);
xnor U14122 (N_14122,N_7446,N_10332);
and U14123 (N_14123,N_6386,N_9445);
xnor U14124 (N_14124,N_6717,N_10983);
and U14125 (N_14125,N_8777,N_11282);
or U14126 (N_14126,N_8786,N_10550);
and U14127 (N_14127,N_10103,N_6366);
nand U14128 (N_14128,N_8547,N_6328);
nand U14129 (N_14129,N_9228,N_8480);
nand U14130 (N_14130,N_11129,N_8541);
nor U14131 (N_14131,N_8409,N_12037);
or U14132 (N_14132,N_9864,N_7495);
and U14133 (N_14133,N_10699,N_12478);
nand U14134 (N_14134,N_8377,N_10743);
nand U14135 (N_14135,N_7761,N_6515);
nor U14136 (N_14136,N_11785,N_11837);
and U14137 (N_14137,N_7048,N_11098);
nand U14138 (N_14138,N_11164,N_9773);
and U14139 (N_14139,N_7496,N_9946);
or U14140 (N_14140,N_8950,N_11056);
xor U14141 (N_14141,N_9255,N_11568);
nand U14142 (N_14142,N_7619,N_9570);
nand U14143 (N_14143,N_7478,N_8038);
and U14144 (N_14144,N_7409,N_12452);
xnor U14145 (N_14145,N_8579,N_7705);
xnor U14146 (N_14146,N_7499,N_7184);
nor U14147 (N_14147,N_8072,N_7368);
xnor U14148 (N_14148,N_7114,N_8750);
nand U14149 (N_14149,N_7003,N_12039);
or U14150 (N_14150,N_11613,N_8779);
nand U14151 (N_14151,N_9245,N_11748);
nand U14152 (N_14152,N_7428,N_12235);
xnor U14153 (N_14153,N_11118,N_9802);
or U14154 (N_14154,N_7738,N_6520);
or U14155 (N_14155,N_9549,N_11342);
or U14156 (N_14156,N_7372,N_11470);
or U14157 (N_14157,N_10274,N_8010);
or U14158 (N_14158,N_10395,N_12030);
xor U14159 (N_14159,N_8793,N_10086);
nand U14160 (N_14160,N_12229,N_9755);
and U14161 (N_14161,N_9308,N_12280);
and U14162 (N_14162,N_7556,N_7900);
nor U14163 (N_14163,N_9221,N_11450);
xnor U14164 (N_14164,N_10627,N_9867);
nand U14165 (N_14165,N_7718,N_9233);
xnor U14166 (N_14166,N_6583,N_10845);
and U14167 (N_14167,N_6338,N_7276);
xnor U14168 (N_14168,N_10014,N_6307);
or U14169 (N_14169,N_10045,N_10771);
xnor U14170 (N_14170,N_7193,N_11040);
or U14171 (N_14171,N_10864,N_10897);
nand U14172 (N_14172,N_6374,N_8313);
nand U14173 (N_14173,N_8151,N_10617);
nand U14174 (N_14174,N_10532,N_11037);
or U14175 (N_14175,N_10435,N_11255);
and U14176 (N_14176,N_10379,N_9682);
or U14177 (N_14177,N_7413,N_11863);
xor U14178 (N_14178,N_10065,N_8582);
or U14179 (N_14179,N_8633,N_11932);
or U14180 (N_14180,N_10449,N_10609);
or U14181 (N_14181,N_6533,N_9710);
or U14182 (N_14182,N_8336,N_9432);
or U14183 (N_14183,N_7991,N_7782);
and U14184 (N_14184,N_10256,N_7983);
or U14185 (N_14185,N_7799,N_6621);
and U14186 (N_14186,N_7374,N_8475);
or U14187 (N_14187,N_11819,N_6760);
nand U14188 (N_14188,N_8412,N_11152);
nor U14189 (N_14189,N_11312,N_10512);
nand U14190 (N_14190,N_12102,N_9637);
nand U14191 (N_14191,N_7550,N_10443);
nor U14192 (N_14192,N_10377,N_10846);
nor U14193 (N_14193,N_7686,N_9266);
nand U14194 (N_14194,N_11121,N_7719);
or U14195 (N_14195,N_8663,N_10930);
or U14196 (N_14196,N_7839,N_10878);
or U14197 (N_14197,N_10774,N_7375);
and U14198 (N_14198,N_10369,N_6474);
xor U14199 (N_14199,N_9585,N_10982);
nand U14200 (N_14200,N_12090,N_7831);
nand U14201 (N_14201,N_10152,N_10671);
nand U14202 (N_14202,N_9910,N_10850);
and U14203 (N_14203,N_10063,N_7516);
or U14204 (N_14204,N_10747,N_11514);
nor U14205 (N_14205,N_6948,N_10040);
nand U14206 (N_14206,N_11168,N_11879);
or U14207 (N_14207,N_12006,N_11428);
and U14208 (N_14208,N_9806,N_10282);
nand U14209 (N_14209,N_6415,N_10910);
and U14210 (N_14210,N_10566,N_7586);
nor U14211 (N_14211,N_6762,N_9278);
xor U14212 (N_14212,N_11821,N_10405);
and U14213 (N_14213,N_9592,N_12043);
or U14214 (N_14214,N_9645,N_10767);
and U14215 (N_14215,N_7728,N_11143);
nor U14216 (N_14216,N_10871,N_9712);
or U14217 (N_14217,N_12269,N_7964);
nand U14218 (N_14218,N_9740,N_10520);
nand U14219 (N_14219,N_6288,N_11249);
nand U14220 (N_14220,N_7327,N_9028);
nor U14221 (N_14221,N_10560,N_12176);
xor U14222 (N_14222,N_8353,N_7841);
nand U14223 (N_14223,N_10326,N_8912);
or U14224 (N_14224,N_8169,N_7155);
and U14225 (N_14225,N_6355,N_11860);
nand U14226 (N_14226,N_10778,N_8981);
nor U14227 (N_14227,N_10039,N_12388);
nand U14228 (N_14228,N_12265,N_10963);
xnor U14229 (N_14229,N_9132,N_7065);
nor U14230 (N_14230,N_8473,N_7595);
nor U14231 (N_14231,N_6485,N_11180);
and U14232 (N_14232,N_12446,N_10123);
xor U14233 (N_14233,N_9227,N_8563);
or U14234 (N_14234,N_6539,N_10360);
xnor U14235 (N_14235,N_9185,N_12418);
nor U14236 (N_14236,N_6323,N_9206);
nand U14237 (N_14237,N_6306,N_6273);
nand U14238 (N_14238,N_9323,N_8064);
nor U14239 (N_14239,N_7098,N_8744);
nor U14240 (N_14240,N_12492,N_8133);
and U14241 (N_14241,N_8628,N_9622);
and U14242 (N_14242,N_8930,N_9782);
and U14243 (N_14243,N_7456,N_10523);
and U14244 (N_14244,N_8452,N_9532);
nor U14245 (N_14245,N_7804,N_9172);
and U14246 (N_14246,N_8635,N_9574);
nor U14247 (N_14247,N_6803,N_6715);
nor U14248 (N_14248,N_7215,N_6665);
nor U14249 (N_14249,N_10614,N_7614);
nor U14250 (N_14250,N_11130,N_8282);
and U14251 (N_14251,N_11710,N_6822);
xnor U14252 (N_14252,N_6452,N_8455);
and U14253 (N_14253,N_7925,N_8885);
and U14254 (N_14254,N_9665,N_7336);
or U14255 (N_14255,N_9629,N_9374);
and U14256 (N_14256,N_10093,N_8438);
and U14257 (N_14257,N_11299,N_11496);
nor U14258 (N_14258,N_12137,N_11891);
and U14259 (N_14259,N_6255,N_7787);
xor U14260 (N_14260,N_7376,N_9231);
xnor U14261 (N_14261,N_8861,N_6570);
or U14262 (N_14262,N_9654,N_10286);
xnor U14263 (N_14263,N_11071,N_7555);
and U14264 (N_14264,N_9792,N_10872);
nor U14265 (N_14265,N_10933,N_8178);
and U14266 (N_14266,N_6429,N_7635);
nand U14267 (N_14267,N_6489,N_8233);
nor U14268 (N_14268,N_10442,N_11123);
xor U14269 (N_14269,N_7014,N_11078);
or U14270 (N_14270,N_9145,N_8161);
or U14271 (N_14271,N_12177,N_11618);
and U14272 (N_14272,N_11023,N_9467);
nor U14273 (N_14273,N_8489,N_6875);
or U14274 (N_14274,N_8959,N_8606);
nor U14275 (N_14275,N_6779,N_8736);
xnor U14276 (N_14276,N_7388,N_12080);
nand U14277 (N_14277,N_8560,N_6295);
and U14278 (N_14278,N_10263,N_10847);
and U14279 (N_14279,N_11629,N_8364);
or U14280 (N_14280,N_6767,N_9832);
and U14281 (N_14281,N_12185,N_6333);
or U14282 (N_14282,N_10328,N_8105);
or U14283 (N_14283,N_9120,N_7672);
xor U14284 (N_14284,N_7291,N_11765);
or U14285 (N_14285,N_10444,N_10977);
or U14286 (N_14286,N_6594,N_8183);
and U14287 (N_14287,N_11902,N_8450);
or U14288 (N_14288,N_7061,N_10944);
xnor U14289 (N_14289,N_8173,N_11154);
xor U14290 (N_14290,N_7612,N_10160);
nand U14291 (N_14291,N_6921,N_7812);
and U14292 (N_14292,N_12164,N_7781);
nor U14293 (N_14293,N_7242,N_6592);
nor U14294 (N_14294,N_7222,N_10111);
nor U14295 (N_14295,N_6305,N_11206);
nand U14296 (N_14296,N_10900,N_8886);
nand U14297 (N_14297,N_8328,N_11656);
nand U14298 (N_14298,N_12282,N_7749);
or U14299 (N_14299,N_8826,N_7730);
nand U14300 (N_14300,N_7624,N_9795);
nand U14301 (N_14301,N_8271,N_6871);
xor U14302 (N_14302,N_6775,N_8622);
or U14303 (N_14303,N_8012,N_8933);
nand U14304 (N_14304,N_11326,N_11160);
nand U14305 (N_14305,N_12256,N_8574);
or U14306 (N_14306,N_12214,N_10164);
nor U14307 (N_14307,N_7060,N_11580);
or U14308 (N_14308,N_10848,N_7844);
xor U14309 (N_14309,N_6648,N_11239);
nand U14310 (N_14310,N_8112,N_8966);
nor U14311 (N_14311,N_10367,N_6535);
nand U14312 (N_14312,N_7924,N_9597);
nor U14313 (N_14313,N_8458,N_7205);
and U14314 (N_14314,N_10656,N_10578);
nand U14315 (N_14315,N_7464,N_12489);
xnor U14316 (N_14316,N_9544,N_12055);
xor U14317 (N_14317,N_7256,N_10456);
or U14318 (N_14318,N_10808,N_8878);
nand U14319 (N_14319,N_6697,N_6813);
or U14320 (N_14320,N_9533,N_6538);
xor U14321 (N_14321,N_9393,N_9209);
nand U14322 (N_14322,N_9925,N_8758);
xnor U14323 (N_14323,N_7316,N_12223);
nor U14324 (N_14324,N_11439,N_11015);
or U14325 (N_14325,N_10397,N_9295);
or U14326 (N_14326,N_8374,N_12089);
nand U14327 (N_14327,N_11434,N_10445);
xor U14328 (N_14328,N_9957,N_8566);
nand U14329 (N_14329,N_9303,N_10807);
nor U14330 (N_14330,N_6432,N_9311);
and U14331 (N_14331,N_8394,N_7140);
nand U14332 (N_14332,N_11250,N_10254);
xnor U14333 (N_14333,N_10819,N_10504);
nor U14334 (N_14334,N_12404,N_8048);
nand U14335 (N_14335,N_9572,N_12338);
or U14336 (N_14336,N_9929,N_10270);
and U14337 (N_14337,N_7075,N_6946);
and U14338 (N_14338,N_10175,N_9263);
and U14339 (N_14339,N_6384,N_10048);
nor U14340 (N_14340,N_9681,N_7880);
nor U14341 (N_14341,N_8195,N_8025);
and U14342 (N_14342,N_7144,N_12163);
or U14343 (N_14343,N_7879,N_9158);
xnor U14344 (N_14344,N_6763,N_10950);
and U14345 (N_14345,N_6477,N_9930);
and U14346 (N_14346,N_8009,N_9598);
nor U14347 (N_14347,N_11138,N_11633);
or U14348 (N_14348,N_7567,N_7830);
xor U14349 (N_14349,N_9728,N_12397);
nand U14350 (N_14350,N_10669,N_11826);
or U14351 (N_14351,N_8730,N_11134);
nand U14352 (N_14352,N_8312,N_10074);
or U14353 (N_14353,N_9758,N_9797);
and U14354 (N_14354,N_10485,N_8145);
nor U14355 (N_14355,N_10290,N_7853);
nor U14356 (N_14356,N_6918,N_7963);
xor U14357 (N_14357,N_9307,N_12245);
or U14358 (N_14358,N_10662,N_10567);
or U14359 (N_14359,N_11729,N_10381);
or U14360 (N_14360,N_7493,N_8871);
or U14361 (N_14361,N_12203,N_10503);
nand U14362 (N_14362,N_10317,N_7312);
or U14363 (N_14363,N_12368,N_9450);
xor U14364 (N_14364,N_6947,N_9577);
nor U14365 (N_14365,N_8667,N_7385);
xnor U14366 (N_14366,N_11169,N_10354);
xor U14367 (N_14367,N_9122,N_9584);
nand U14368 (N_14368,N_8011,N_8770);
and U14369 (N_14369,N_10675,N_9394);
and U14370 (N_14370,N_9285,N_6356);
nand U14371 (N_14371,N_6710,N_6601);
or U14372 (N_14372,N_9079,N_11214);
nand U14373 (N_14373,N_10931,N_8054);
nor U14374 (N_14374,N_10533,N_6999);
nor U14375 (N_14375,N_12298,N_7868);
xor U14376 (N_14376,N_10865,N_9752);
xnor U14377 (N_14377,N_10463,N_7982);
nand U14378 (N_14378,N_6354,N_7622);
xnor U14379 (N_14379,N_9937,N_9659);
xor U14380 (N_14380,N_10832,N_10556);
nand U14381 (N_14381,N_8140,N_9056);
nand U14382 (N_14382,N_11998,N_9804);
or U14383 (N_14383,N_11497,N_9196);
and U14384 (N_14384,N_7273,N_8548);
nor U14385 (N_14385,N_8302,N_9997);
or U14386 (N_14386,N_10253,N_11417);
or U14387 (N_14387,N_6909,N_6577);
nand U14388 (N_14388,N_6651,N_10268);
or U14389 (N_14389,N_8242,N_7952);
nor U14390 (N_14390,N_6302,N_9279);
xnor U14391 (N_14391,N_9259,N_8496);
and U14392 (N_14392,N_11643,N_9529);
and U14393 (N_14393,N_10705,N_9406);
xnor U14394 (N_14394,N_8366,N_10366);
and U14395 (N_14395,N_7245,N_10555);
or U14396 (N_14396,N_6922,N_8078);
xnor U14397 (N_14397,N_11759,N_7492);
and U14398 (N_14398,N_11982,N_8530);
or U14399 (N_14399,N_7526,N_10548);
nand U14400 (N_14400,N_11647,N_9868);
or U14401 (N_14401,N_7777,N_11544);
and U14402 (N_14402,N_7798,N_12222);
and U14403 (N_14403,N_8945,N_11731);
and U14404 (N_14404,N_6994,N_8032);
nand U14405 (N_14405,N_11207,N_8811);
nand U14406 (N_14406,N_9525,N_11925);
nor U14407 (N_14407,N_8174,N_12384);
or U14408 (N_14408,N_6558,N_12001);
xor U14409 (N_14409,N_8882,N_9403);
and U14410 (N_14410,N_11472,N_7214);
and U14411 (N_14411,N_8778,N_12189);
nor U14412 (N_14412,N_12225,N_7342);
nand U14413 (N_14413,N_11810,N_11882);
or U14414 (N_14414,N_9325,N_10937);
or U14415 (N_14415,N_10218,N_7620);
nand U14416 (N_14416,N_11683,N_7229);
or U14417 (N_14417,N_8982,N_10213);
or U14418 (N_14418,N_9427,N_8659);
nand U14419 (N_14419,N_7540,N_7821);
and U14420 (N_14420,N_10053,N_7024);
and U14421 (N_14421,N_7247,N_7974);
xor U14422 (N_14422,N_9742,N_12226);
xnor U14423 (N_14423,N_8000,N_11585);
or U14424 (N_14424,N_8911,N_9163);
xnor U14425 (N_14425,N_8683,N_11954);
and U14426 (N_14426,N_10830,N_11653);
nand U14427 (N_14427,N_10735,N_7390);
nand U14428 (N_14428,N_7102,N_10387);
xnor U14429 (N_14429,N_6459,N_6913);
or U14430 (N_14430,N_10776,N_6373);
nand U14431 (N_14431,N_9660,N_10339);
nor U14432 (N_14432,N_10264,N_7463);
nand U14433 (N_14433,N_9994,N_7281);
nor U14434 (N_14434,N_8196,N_10831);
nand U14435 (N_14435,N_10150,N_11090);
nor U14436 (N_14436,N_6293,N_11829);
xnor U14437 (N_14437,N_9697,N_9292);
nor U14438 (N_14438,N_9975,N_9229);
or U14439 (N_14439,N_9907,N_9747);
or U14440 (N_14440,N_8034,N_11855);
xor U14441 (N_14441,N_10979,N_7037);
nand U14442 (N_14442,N_10277,N_12048);
nor U14443 (N_14443,N_9716,N_10312);
and U14444 (N_14444,N_10891,N_7497);
and U14445 (N_14445,N_11553,N_7169);
and U14446 (N_14446,N_9011,N_6615);
or U14447 (N_14447,N_7109,N_10023);
nand U14448 (N_14448,N_6368,N_6252);
or U14449 (N_14449,N_6514,N_10330);
nand U14450 (N_14450,N_7482,N_11200);
xor U14451 (N_14451,N_9291,N_7407);
xnor U14452 (N_14452,N_10506,N_12372);
nand U14453 (N_14453,N_11619,N_11980);
nand U14454 (N_14454,N_9748,N_9923);
nor U14455 (N_14455,N_10602,N_11689);
nand U14456 (N_14456,N_7611,N_6603);
and U14457 (N_14457,N_6887,N_9833);
nor U14458 (N_14458,N_9875,N_7139);
nand U14459 (N_14459,N_11115,N_7626);
and U14460 (N_14460,N_9318,N_9865);
nand U14461 (N_14461,N_7521,N_7609);
nand U14462 (N_14462,N_7332,N_12419);
and U14463 (N_14463,N_6455,N_7417);
and U14464 (N_14464,N_12191,N_7268);
or U14465 (N_14465,N_12299,N_7280);
nand U14466 (N_14466,N_11943,N_12395);
or U14467 (N_14467,N_7382,N_10635);
or U14468 (N_14468,N_11589,N_10233);
and U14469 (N_14469,N_8897,N_6586);
nand U14470 (N_14470,N_9671,N_8294);
and U14471 (N_14471,N_10221,N_9881);
nor U14472 (N_14472,N_12345,N_11739);
nand U14473 (N_14473,N_12058,N_11501);
or U14474 (N_14474,N_7404,N_10752);
and U14475 (N_14475,N_11012,N_7621);
nand U14476 (N_14476,N_8027,N_8017);
nor U14477 (N_14477,N_11749,N_6869);
nor U14478 (N_14478,N_7082,N_7239);
nor U14479 (N_14479,N_10359,N_11256);
xor U14480 (N_14480,N_11789,N_9389);
xor U14481 (N_14481,N_10076,N_7627);
nand U14482 (N_14482,N_11927,N_8585);
and U14483 (N_14483,N_9408,N_8243);
xnor U14484 (N_14484,N_10289,N_6364);
or U14485 (N_14485,N_9686,N_6598);
or U14486 (N_14486,N_9437,N_6251);
nor U14487 (N_14487,N_9998,N_10480);
or U14488 (N_14488,N_9649,N_6962);
or U14489 (N_14489,N_6456,N_7893);
nand U14490 (N_14490,N_9336,N_7350);
and U14491 (N_14491,N_9820,N_11389);
or U14492 (N_14492,N_8446,N_10116);
xnor U14493 (N_14493,N_10833,N_6790);
and U14494 (N_14494,N_10815,N_10908);
nor U14495 (N_14495,N_6711,N_12202);
or U14496 (N_14496,N_9275,N_6984);
nand U14497 (N_14497,N_7083,N_10946);
xnor U14498 (N_14498,N_9277,N_11502);
nand U14499 (N_14499,N_10895,N_6300);
xor U14500 (N_14500,N_12221,N_7078);
nor U14501 (N_14501,N_7323,N_7366);
and U14502 (N_14502,N_10976,N_11406);
xor U14503 (N_14503,N_6420,N_9565);
and U14504 (N_14504,N_9809,N_10300);
and U14505 (N_14505,N_7852,N_11903);
xor U14506 (N_14506,N_12403,N_9569);
nor U14507 (N_14507,N_7177,N_8031);
and U14508 (N_14508,N_7869,N_6497);
xor U14509 (N_14509,N_11165,N_12426);
nand U14510 (N_14510,N_11916,N_7848);
or U14511 (N_14511,N_8013,N_6777);
xor U14512 (N_14512,N_10683,N_9547);
nor U14513 (N_14513,N_11237,N_8091);
nand U14514 (N_14514,N_12073,N_12013);
or U14515 (N_14515,N_9761,N_8597);
xnor U14516 (N_14516,N_9986,N_6781);
xnor U14517 (N_14517,N_11022,N_12171);
nor U14518 (N_14518,N_10009,N_11968);
and U14519 (N_14519,N_11321,N_11000);
nand U14520 (N_14520,N_7822,N_11063);
nor U14521 (N_14521,N_7588,N_8219);
or U14522 (N_14522,N_11885,N_10997);
or U14523 (N_14523,N_11446,N_6843);
and U14524 (N_14524,N_12346,N_12071);
and U14525 (N_14525,N_9006,N_9076);
nor U14526 (N_14526,N_8965,N_6818);
and U14527 (N_14527,N_7450,N_7514);
xnor U14528 (N_14528,N_6264,N_8225);
xnor U14529 (N_14529,N_8200,N_10729);
or U14530 (N_14530,N_11459,N_10881);
and U14531 (N_14531,N_8171,N_9966);
and U14532 (N_14532,N_9153,N_12312);
and U14533 (N_14533,N_12017,N_11874);
or U14534 (N_14534,N_12458,N_8534);
nand U14535 (N_14535,N_9054,N_7943);
nor U14536 (N_14536,N_11993,N_9695);
nand U14537 (N_14537,N_11540,N_9784);
nand U14538 (N_14538,N_8131,N_9224);
nand U14539 (N_14539,N_9839,N_12062);
nor U14540 (N_14540,N_7364,N_10204);
and U14541 (N_14541,N_11367,N_9534);
and U14542 (N_14542,N_7444,N_9969);
or U14543 (N_14543,N_11695,N_9451);
nand U14544 (N_14544,N_8644,N_9675);
and U14545 (N_14545,N_7920,N_12070);
nor U14546 (N_14546,N_10969,N_11380);
xor U14547 (N_14547,N_8144,N_10220);
and U14548 (N_14548,N_9830,N_6737);
or U14549 (N_14549,N_8887,N_7814);
nor U14550 (N_14550,N_6831,N_7397);
nand U14551 (N_14551,N_10003,N_8380);
or U14552 (N_14552,N_8909,N_10777);
or U14553 (N_14553,N_8416,N_12466);
or U14554 (N_14554,N_9058,N_11455);
and U14555 (N_14555,N_11347,N_10306);
xor U14556 (N_14556,N_10612,N_9936);
nand U14557 (N_14557,N_11058,N_11074);
nor U14558 (N_14558,N_10391,N_12061);
and U14559 (N_14559,N_9563,N_9953);
nand U14560 (N_14560,N_6322,N_7997);
nor U14561 (N_14561,N_7210,N_11599);
nor U14562 (N_14562,N_7165,N_11453);
and U14563 (N_14563,N_9479,N_6820);
and U14564 (N_14564,N_10536,N_7423);
nand U14565 (N_14565,N_6410,N_6545);
and U14566 (N_14566,N_11723,N_7217);
nand U14567 (N_14567,N_6458,N_7707);
or U14568 (N_14568,N_10127,N_11498);
xnor U14569 (N_14569,N_9543,N_11530);
nand U14570 (N_14570,N_10088,N_11073);
nand U14571 (N_14571,N_12003,N_10467);
or U14572 (N_14572,N_9961,N_12467);
nand U14573 (N_14573,N_11414,N_6672);
nand U14574 (N_14574,N_11194,N_11252);
or U14575 (N_14575,N_7962,N_10719);
or U14576 (N_14576,N_12066,N_11674);
nor U14577 (N_14577,N_11113,N_7865);
xor U14578 (N_14578,N_10974,N_8954);
xor U14579 (N_14579,N_6815,N_6970);
nand U14580 (N_14580,N_6402,N_8634);
nand U14581 (N_14581,N_10684,N_6817);
nor U14582 (N_14582,N_10378,N_12149);
and U14583 (N_14583,N_8287,N_10826);
nand U14584 (N_14584,N_12040,N_7538);
xnor U14585 (N_14585,N_7919,N_9089);
nor U14586 (N_14586,N_9983,N_10222);
xor U14587 (N_14587,N_11320,N_6783);
or U14588 (N_14588,N_9192,N_11582);
nor U14589 (N_14589,N_6714,N_6654);
nand U14590 (N_14590,N_9670,N_7179);
or U14591 (N_14591,N_6865,N_9783);
nor U14592 (N_14592,N_7447,N_7052);
or U14593 (N_14593,N_9092,N_9749);
nand U14594 (N_14594,N_10919,N_6873);
nor U14595 (N_14595,N_7647,N_7651);
nand U14596 (N_14596,N_11416,N_9694);
xor U14597 (N_14597,N_9733,N_6447);
nor U14598 (N_14598,N_9714,N_8417);
nand U14599 (N_14599,N_9505,N_10223);
or U14600 (N_14600,N_9497,N_9159);
nand U14601 (N_14601,N_8014,N_10244);
or U14602 (N_14602,N_7275,N_9509);
and U14603 (N_14603,N_10114,N_7259);
xnor U14604 (N_14604,N_7319,N_7993);
xnor U14605 (N_14605,N_12067,N_7197);
or U14606 (N_14606,N_8986,N_10125);
xnor U14607 (N_14607,N_8468,N_9252);
or U14608 (N_14608,N_10436,N_9882);
xnor U14609 (N_14609,N_9446,N_10985);
and U14610 (N_14610,N_8681,N_10368);
and U14611 (N_14611,N_12411,N_8314);
or U14612 (N_14612,N_8537,N_10327);
nand U14613 (N_14613,N_12239,N_9381);
xor U14614 (N_14614,N_12353,N_11719);
or U14615 (N_14615,N_11602,N_7460);
nand U14616 (N_14616,N_11148,N_6414);
nor U14617 (N_14617,N_6967,N_9340);
xor U14618 (N_14618,N_11922,N_8596);
or U14619 (N_14619,N_7399,N_9873);
xnor U14620 (N_14620,N_9462,N_8970);
or U14621 (N_14621,N_9538,N_6772);
nor U14622 (N_14622,N_11059,N_6997);
or U14623 (N_14623,N_7357,N_8397);
nor U14624 (N_14624,N_8085,N_9165);
nor U14625 (N_14625,N_9247,N_9941);
or U14626 (N_14626,N_8938,N_11586);
nand U14627 (N_14627,N_11029,N_11322);
nor U14628 (N_14628,N_9024,N_7064);
nand U14629 (N_14629,N_8418,N_11752);
nor U14630 (N_14630,N_8864,N_11142);
nand U14631 (N_14631,N_12356,N_7531);
nand U14632 (N_14632,N_12086,N_6574);
nand U14633 (N_14633,N_11992,N_8624);
or U14634 (N_14634,N_6786,N_9007);
xor U14635 (N_14635,N_10657,N_9646);
nand U14636 (N_14636,N_7818,N_11351);
nor U14637 (N_14637,N_7623,N_10570);
nand U14638 (N_14638,N_9980,N_12427);
or U14639 (N_14639,N_8155,N_9489);
nor U14640 (N_14640,N_7768,N_7688);
or U14641 (N_14641,N_9734,N_10493);
xnor U14642 (N_14642,N_10465,N_12284);
or U14643 (N_14643,N_11535,N_10182);
or U14644 (N_14644,N_8760,N_6267);
nor U14645 (N_14645,N_9102,N_11554);
nor U14646 (N_14646,N_7359,N_10431);
or U14647 (N_14647,N_7349,N_6378);
and U14648 (N_14648,N_8339,N_12359);
nand U14649 (N_14649,N_10901,N_6416);
or U14650 (N_14650,N_8592,N_10384);
xor U14651 (N_14651,N_9824,N_8222);
nor U14652 (N_14652,N_9179,N_9564);
xnor U14653 (N_14653,N_8705,N_8401);
nor U14654 (N_14654,N_8605,N_10198);
nor U14655 (N_14655,N_6723,N_7116);
and U14656 (N_14656,N_11275,N_6814);
nand U14657 (N_14657,N_8713,N_9199);
and U14658 (N_14658,N_10389,N_7498);
xnor U14659 (N_14659,N_7156,N_7185);
and U14660 (N_14660,N_11805,N_10482);
nor U14661 (N_14661,N_8356,N_11227);
xor U14662 (N_14662,N_11625,N_12285);
nor U14663 (N_14663,N_7361,N_9239);
nor U14664 (N_14664,N_7899,N_9097);
xor U14665 (N_14665,N_10059,N_11973);
and U14666 (N_14666,N_6417,N_12336);
nand U14667 (N_14667,N_9631,N_10408);
nor U14668 (N_14668,N_10858,N_10727);
or U14669 (N_14669,N_6652,N_11552);
or U14670 (N_14670,N_6318,N_8594);
nor U14671 (N_14671,N_8428,N_10915);
or U14672 (N_14672,N_10718,N_11557);
nor U14673 (N_14673,N_11965,N_11107);
nor U14674 (N_14674,N_9954,N_11382);
and U14675 (N_14675,N_11006,N_7449);
nor U14676 (N_14676,N_10146,N_8284);
nor U14677 (N_14677,N_11269,N_9763);
and U14678 (N_14678,N_9430,N_6575);
xnor U14679 (N_14679,N_11223,N_8675);
and U14680 (N_14680,N_10643,N_10032);
xnor U14681 (N_14681,N_6503,N_6522);
nor U14682 (N_14682,N_7508,N_6632);
and U14683 (N_14683,N_6899,N_11391);
or U14684 (N_14684,N_12447,N_8873);
nand U14685 (N_14685,N_12129,N_10197);
or U14686 (N_14686,N_8179,N_7628);
nor U14687 (N_14687,N_8814,N_8846);
or U14688 (N_14688,N_11341,N_10886);
nand U14689 (N_14689,N_8503,N_10278);
xor U14690 (N_14690,N_11948,N_7727);
or U14691 (N_14691,N_12363,N_12087);
or U14692 (N_14692,N_8044,N_7928);
or U14693 (N_14693,N_9112,N_9433);
nand U14694 (N_14694,N_10716,N_11628);
nand U14695 (N_14695,N_12376,N_10240);
or U14696 (N_14696,N_12304,N_10519);
nor U14697 (N_14697,N_11996,N_10818);
xnor U14698 (N_14698,N_7917,N_6359);
nand U14699 (N_14699,N_11728,N_7754);
nor U14700 (N_14700,N_11386,N_9556);
nand U14701 (N_14701,N_8263,N_11645);
xnor U14702 (N_14702,N_9177,N_7243);
xnor U14703 (N_14703,N_9170,N_8226);
nand U14704 (N_14704,N_11935,N_7552);
nor U14705 (N_14705,N_7823,N_6573);
or U14706 (N_14706,N_7203,N_10121);
nor U14707 (N_14707,N_9175,N_7094);
nand U14708 (N_14708,N_11836,N_8362);
nand U14709 (N_14709,N_7089,N_9770);
or U14710 (N_14710,N_11780,N_8870);
xnor U14711 (N_14711,N_8623,N_9568);
nor U14712 (N_14712,N_6618,N_9371);
nor U14713 (N_14713,N_10622,N_8830);
xor U14714 (N_14714,N_7808,N_10034);
xor U14715 (N_14715,N_8818,N_9996);
or U14716 (N_14716,N_8160,N_12206);
or U14717 (N_14717,N_12390,N_7750);
or U14718 (N_14718,N_8492,N_6721);
or U14719 (N_14719,N_7742,N_6703);
nor U14720 (N_14720,N_12257,N_10723);
nor U14721 (N_14721,N_6400,N_11044);
nand U14722 (N_14722,N_8820,N_7527);
and U14723 (N_14723,N_9141,N_10751);
xor U14724 (N_14724,N_7937,N_6614);
and U14725 (N_14725,N_7987,N_6593);
nand U14726 (N_14726,N_8237,N_8434);
nand U14727 (N_14727,N_6396,N_9099);
nor U14728 (N_14728,N_8239,N_11921);
or U14729 (N_14729,N_8516,N_8829);
nand U14730 (N_14730,N_6769,N_6712);
and U14731 (N_14731,N_9948,N_6677);
xor U14732 (N_14732,N_8244,N_8399);
or U14733 (N_14733,N_6568,N_9984);
or U14734 (N_14734,N_7921,N_8738);
xor U14735 (N_14735,N_6854,N_9987);
xnor U14736 (N_14736,N_10469,N_6669);
xor U14737 (N_14737,N_10928,N_9711);
nor U14738 (N_14738,N_11360,N_8804);
and U14739 (N_14739,N_7344,N_6851);
and U14740 (N_14740,N_7912,N_10452);
xor U14741 (N_14741,N_12493,N_12498);
nor U14742 (N_14742,N_7838,N_9702);
and U14743 (N_14743,N_11423,N_8095);
and U14744 (N_14744,N_9494,N_8810);
nor U14745 (N_14745,N_12288,N_9771);
and U14746 (N_14746,N_10067,N_8572);
xnor U14747 (N_14747,N_10494,N_11381);
or U14748 (N_14748,N_7649,N_8055);
xnor U14749 (N_14749,N_9610,N_9559);
nor U14750 (N_14750,N_7845,N_10345);
or U14751 (N_14751,N_11512,N_8390);
xor U14752 (N_14752,N_6569,N_7286);
nor U14753 (N_14753,N_6876,N_11392);
nor U14754 (N_14754,N_9459,N_6422);
nor U14755 (N_14755,N_11224,N_8456);
nand U14756 (N_14756,N_10805,N_9901);
xnor U14757 (N_14757,N_12125,N_11937);
and U14758 (N_14758,N_8419,N_12153);
nor U14759 (N_14759,N_8135,N_8406);
nor U14760 (N_14760,N_10748,N_10854);
xnor U14761 (N_14761,N_11010,N_11457);
and U14762 (N_14762,N_8641,N_9723);
and U14763 (N_14763,N_8215,N_11676);
nor U14764 (N_14764,N_8868,N_7445);
nand U14765 (N_14765,N_6675,N_7176);
and U14766 (N_14766,N_7154,N_11292);
and U14767 (N_14767,N_10168,N_9895);
or U14768 (N_14768,N_10898,N_11763);
or U14769 (N_14769,N_9201,N_8410);
nor U14770 (N_14770,N_8590,N_11492);
nand U14771 (N_14771,N_12146,N_6896);
and U14772 (N_14772,N_11487,N_11141);
and U14773 (N_14773,N_8514,N_9146);
or U14774 (N_14774,N_7157,N_11461);
nor U14775 (N_14775,N_11995,N_11878);
nand U14776 (N_14776,N_7455,N_6933);
and U14777 (N_14777,N_9216,N_9590);
nor U14778 (N_14778,N_6724,N_10746);
xor U14779 (N_14779,N_11791,N_8310);
xor U14780 (N_14780,N_10936,N_7298);
nor U14781 (N_14781,N_9253,N_6722);
or U14782 (N_14782,N_6680,N_9687);
nand U14783 (N_14783,N_7966,N_10813);
or U14784 (N_14784,N_10371,N_9825);
or U14785 (N_14785,N_9375,N_8557);
xor U14786 (N_14786,N_8700,N_10376);
xnor U14787 (N_14787,N_7544,N_6527);
nand U14788 (N_14788,N_8407,N_7663);
and U14789 (N_14789,N_8697,N_7519);
nand U14790 (N_14790,N_8248,N_10440);
or U14791 (N_14791,N_11444,N_11845);
xor U14792 (N_14792,N_6698,N_8241);
nor U14793 (N_14793,N_11875,N_7476);
nor U14794 (N_14794,N_6849,N_8792);
xnor U14795 (N_14795,N_6816,N_8460);
and U14796 (N_14796,N_6734,N_12038);
nand U14797 (N_14797,N_12018,N_8819);
and U14798 (N_14798,N_11551,N_6699);
nor U14799 (N_14799,N_9522,N_11849);
nor U14800 (N_14800,N_10957,N_8023);
xor U14801 (N_14801,N_7815,N_12027);
nor U14802 (N_14802,N_7971,N_12021);
nand U14803 (N_14803,N_7969,N_9114);
xnor U14804 (N_14804,N_9699,N_8554);
xor U14805 (N_14805,N_6766,N_8952);
or U14806 (N_14806,N_10795,N_7806);
or U14807 (N_14807,N_10650,N_7017);
and U14808 (N_14808,N_11851,N_11724);
nand U14809 (N_14809,N_6623,N_7429);
and U14810 (N_14810,N_11093,N_10571);
nand U14811 (N_14811,N_7149,N_12342);
or U14812 (N_14812,N_12057,N_9351);
nor U14813 (N_14813,N_8321,N_11048);
xnor U14814 (N_14814,N_8586,N_9630);
or U14815 (N_14815,N_10859,N_7187);
nand U14816 (N_14816,N_6893,N_7393);
xor U14817 (N_14817,N_9510,N_6395);
xnor U14818 (N_14818,N_11627,N_7820);
xor U14819 (N_14819,N_6464,N_9034);
nor U14820 (N_14820,N_11556,N_8146);
nand U14821 (N_14821,N_9617,N_10949);
xnor U14822 (N_14822,N_10773,N_9397);
nor U14823 (N_14823,N_7760,N_11610);
nand U14824 (N_14824,N_10432,N_9361);
or U14825 (N_14825,N_12216,N_7391);
and U14826 (N_14826,N_9931,N_8437);
xnor U14827 (N_14827,N_7690,N_10250);
and U14828 (N_14828,N_9329,N_10640);
or U14829 (N_14829,N_8646,N_11509);
xor U14830 (N_14830,N_8022,N_6281);
or U14831 (N_14831,N_9065,N_7776);
or U14832 (N_14832,N_8619,N_10687);
xor U14833 (N_14833,N_8711,N_8677);
nand U14834 (N_14834,N_6528,N_11177);
xnor U14835 (N_14835,N_11485,N_12374);
or U14836 (N_14836,N_11137,N_11085);
xor U14837 (N_14837,N_9664,N_11644);
or U14838 (N_14838,N_9967,N_9950);
xnor U14839 (N_14839,N_8498,N_7459);
nor U14840 (N_14840,N_9095,N_8783);
nor U14841 (N_14841,N_10692,N_9679);
and U14842 (N_14842,N_10594,N_8359);
nor U14843 (N_14843,N_6390,N_10132);
xor U14844 (N_14844,N_7077,N_8430);
and U14845 (N_14845,N_7394,N_12251);
or U14846 (N_14846,N_6837,N_8299);
and U14847 (N_14847,N_9874,N_8974);
xnor U14848 (N_14848,N_10492,N_11866);
xor U14849 (N_14849,N_8477,N_6810);
nand U14850 (N_14850,N_12424,N_10822);
xor U14851 (N_14851,N_11338,N_8542);
and U14852 (N_14852,N_9235,N_9455);
xor U14853 (N_14853,N_10501,N_10064);
and U14854 (N_14854,N_9105,N_7168);
nand U14855 (N_14855,N_12180,N_12098);
xnor U14856 (N_14856,N_7968,N_11668);
xnor U14857 (N_14857,N_9480,N_12130);
and U14858 (N_14858,N_6361,N_8805);
and U14859 (N_14859,N_12491,N_11385);
or U14860 (N_14860,N_11182,N_12147);
nor U14861 (N_14861,N_9360,N_9582);
xor U14862 (N_14862,N_10167,N_9579);
nand U14863 (N_14863,N_8717,N_9837);
and U14864 (N_14864,N_9730,N_6902);
and U14865 (N_14865,N_12246,N_7406);
nor U14866 (N_14866,N_11402,N_9973);
nor U14867 (N_14867,N_11069,N_12231);
xor U14868 (N_14868,N_11308,N_8163);
nor U14869 (N_14869,N_6581,N_6682);
nor U14870 (N_14870,N_7400,N_7736);
nor U14871 (N_14871,N_12178,N_10117);
xnor U14872 (N_14872,N_11812,N_8969);
nand U14873 (N_14873,N_6660,N_7936);
or U14874 (N_14874,N_10183,N_8694);
nor U14875 (N_14875,N_10037,N_12232);
or U14876 (N_14876,N_11547,N_6915);
nand U14877 (N_14877,N_10310,N_11420);
or U14878 (N_14878,N_9069,N_10083);
nand U14879 (N_14879,N_9094,N_6612);
xor U14880 (N_14880,N_8148,N_8953);
or U14881 (N_14881,N_8240,N_11776);
xor U14882 (N_14882,N_6421,N_12136);
and U14883 (N_14883,N_9974,N_9287);
nand U14884 (N_14884,N_11383,N_10835);
and U14885 (N_14885,N_7685,N_7946);
xor U14886 (N_14886,N_8021,N_9488);
or U14887 (N_14887,N_9005,N_9078);
nand U14888 (N_14888,N_12455,N_9636);
and U14889 (N_14889,N_12140,N_10863);
nand U14890 (N_14890,N_7317,N_7654);
nor U14891 (N_14891,N_6549,N_12357);
nand U14892 (N_14892,N_8707,N_9993);
xor U14893 (N_14893,N_8529,N_7090);
nor U14894 (N_14894,N_10392,N_7174);
nor U14895 (N_14895,N_10346,N_9456);
nor U14896 (N_14896,N_7525,N_6572);
or U14897 (N_14897,N_9337,N_9604);
xor U14898 (N_14898,N_9688,N_9635);
xnor U14899 (N_14899,N_11737,N_8062);
nand U14900 (N_14900,N_9241,N_7072);
xnor U14901 (N_14901,N_12065,N_12315);
or U14902 (N_14902,N_11495,N_11698);
nor U14903 (N_14903,N_9483,N_7825);
nand U14904 (N_14904,N_8888,N_7307);
xor U14905 (N_14905,N_8580,N_10545);
nand U14906 (N_14906,N_10394,N_10540);
nand U14907 (N_14907,N_6331,N_6597);
nor U14908 (N_14908,N_10661,N_10990);
or U14909 (N_14909,N_7494,N_7523);
and U14910 (N_14910,N_7396,N_11279);
nand U14911 (N_14911,N_12230,N_6874);
xor U14912 (N_14912,N_12306,N_7107);
and U14913 (N_14913,N_10917,N_12252);
nand U14914 (N_14914,N_9700,N_9859);
and U14915 (N_14915,N_9943,N_10625);
or U14916 (N_14916,N_6912,N_11076);
and U14917 (N_14917,N_11053,N_8035);
xor U14918 (N_14918,N_8519,N_8660);
nand U14919 (N_14919,N_11905,N_11864);
xor U14920 (N_14920,N_11400,N_11212);
xor U14921 (N_14921,N_10991,N_12483);
and U14922 (N_14922,N_8709,N_6613);
or U14923 (N_14923,N_7151,N_10070);
nor U14924 (N_14924,N_11725,N_10707);
or U14925 (N_14925,N_9891,N_8265);
nand U14926 (N_14926,N_7918,N_12461);
or U14927 (N_14927,N_7535,N_8400);
nand U14928 (N_14928,N_10448,N_8045);
or U14929 (N_14929,N_7571,N_6441);
xor U14930 (N_14930,N_7894,N_7501);
nor U14931 (N_14931,N_6588,N_7044);
and U14932 (N_14932,N_7606,N_11898);
xnor U14933 (N_14933,N_7992,N_8288);
and U14934 (N_14934,N_8600,N_8688);
nor U14935 (N_14935,N_11747,N_7854);
and U14936 (N_14936,N_10322,N_11260);
and U14937 (N_14937,N_11488,N_10228);
or U14938 (N_14938,N_10749,N_9623);
nand U14939 (N_14939,N_6380,N_10016);
nand U14940 (N_14940,N_12212,N_9458);
or U14941 (N_14941,N_11699,N_9746);
nand U14942 (N_14942,N_11186,N_8026);
or U14943 (N_14943,N_10252,N_8324);
nor U14944 (N_14944,N_11960,N_7095);
and U14945 (N_14945,N_9821,N_6407);
xor U14946 (N_14946,N_6683,N_11975);
nand U14947 (N_14947,N_7472,N_8159);
nor U14948 (N_14948,N_11620,N_7714);
and U14949 (N_14949,N_11859,N_10697);
nand U14950 (N_14950,N_9137,N_6942);
xnor U14951 (N_14951,N_11928,N_6551);
xor U14952 (N_14952,N_12499,N_10179);
or U14953 (N_14953,N_8466,N_7646);
nor U14954 (N_14954,N_11952,N_6676);
nor U14955 (N_14955,N_7658,N_9365);
and U14956 (N_14956,N_12480,N_9210);
and U14957 (N_14957,N_10641,N_11183);
and U14958 (N_14958,N_8202,N_11464);
and U14959 (N_14959,N_10637,N_6525);
or U14960 (N_14960,N_9367,N_12042);
or U14961 (N_14961,N_11094,N_7650);
xor U14962 (N_14962,N_11262,N_9918);
nor U14963 (N_14963,N_10084,N_8643);
xnor U14964 (N_14964,N_12451,N_11244);
nor U14965 (N_14965,N_8185,N_8301);
or U14966 (N_14966,N_12244,N_11471);
and U14967 (N_14967,N_11506,N_8182);
nor U14968 (N_14968,N_7274,N_10693);
or U14969 (N_14969,N_10842,N_8724);
nand U14970 (N_14970,N_10939,N_6517);
xor U14971 (N_14971,N_8684,N_7906);
and U14972 (N_14972,N_7926,N_6327);
nand U14973 (N_14973,N_6330,N_9776);
xnor U14974 (N_14974,N_6607,N_6622);
and U14975 (N_14975,N_10580,N_11310);
or U14976 (N_14976,N_8128,N_8354);
xor U14977 (N_14977,N_8411,N_7412);
or U14978 (N_14978,N_7625,N_12068);
nand U14979 (N_14979,N_10733,N_8553);
nand U14980 (N_14980,N_8317,N_6840);
nand U14981 (N_14981,N_9638,N_6256);
nand U14982 (N_14982,N_8465,N_11377);
or U14983 (N_14983,N_11348,N_10375);
and U14984 (N_14984,N_6268,N_9977);
or U14985 (N_14985,N_6324,N_11813);
xor U14986 (N_14986,N_8236,N_8451);
or U14987 (N_14987,N_7325,N_8386);
nor U14988 (N_14988,N_8344,N_9481);
nand U14989 (N_14989,N_9785,N_8989);
and U14990 (N_14990,N_10466,N_7563);
or U14991 (N_14991,N_11772,N_7096);
nand U14992 (N_14992,N_7789,N_10307);
nor U14993 (N_14993,N_11306,N_11261);
nand U14994 (N_14994,N_12454,N_7081);
nand U14995 (N_14995,N_9906,N_9377);
xor U14996 (N_14996,N_8082,N_7701);
nor U14997 (N_14997,N_10129,N_7293);
nand U14998 (N_14998,N_8371,N_6644);
xnor U14999 (N_14999,N_9257,N_10259);
xnor U15000 (N_15000,N_10382,N_6348);
or U15001 (N_15001,N_8703,N_11511);
nor U15002 (N_15002,N_12121,N_7474);
nor U15003 (N_15003,N_8828,N_9693);
xnor U15004 (N_15004,N_12457,N_8251);
nor U15005 (N_15005,N_10500,N_8609);
nand U15006 (N_15006,N_6624,N_6254);
and U15007 (N_15007,N_8939,N_7722);
and U15008 (N_15008,N_6279,N_11364);
xor U15009 (N_15009,N_12238,N_12004);
nor U15010 (N_15010,N_6620,N_8937);
nor U15011 (N_15011,N_12362,N_7180);
xnor U15012 (N_15012,N_6744,N_9334);
nand U15013 (N_15013,N_7504,N_6693);
and U15014 (N_15014,N_11746,N_8510);
nand U15015 (N_15015,N_11061,N_6859);
nor U15016 (N_15016,N_11569,N_11637);
or U15017 (N_15017,N_11868,N_11232);
nor U15018 (N_15018,N_10095,N_10102);
nor U15019 (N_15019,N_8638,N_10119);
nor U15020 (N_15020,N_11893,N_7158);
nor U15021 (N_15021,N_7135,N_8856);
nor U15022 (N_15022,N_9232,N_8632);
or U15023 (N_15023,N_6827,N_9372);
nand U15024 (N_15024,N_11345,N_6389);
and U15025 (N_15025,N_11361,N_8751);
nand U15026 (N_15026,N_12320,N_11635);
xnor U15027 (N_15027,N_7085,N_10758);
xnor U15028 (N_15028,N_7365,N_10242);
or U15029 (N_15029,N_9781,N_12167);
or U15030 (N_15030,N_9048,N_10694);
nand U15031 (N_15031,N_12297,N_11468);
and U15032 (N_15032,N_12431,N_6344);
xnor U15033 (N_15033,N_8964,N_11336);
and U15034 (N_15034,N_11561,N_9810);
nand U15035 (N_15035,N_6562,N_10592);
or U15036 (N_15036,N_9495,N_8485);
xnor U15037 (N_15037,N_7190,N_11116);
nand U15038 (N_15038,N_9423,N_7643);
nand U15039 (N_15039,N_7889,N_9436);
and U15040 (N_15040,N_11846,N_11549);
nand U15041 (N_15041,N_6673,N_7607);
and U15042 (N_15042,N_6314,N_7600);
nor U15043 (N_15043,N_8682,N_6657);
nor U15044 (N_15044,N_10882,N_8549);
and U15045 (N_15045,N_12400,N_10438);
and U15046 (N_15046,N_8746,N_6561);
nor U15047 (N_15047,N_10407,N_6508);
xor U15048 (N_15048,N_10038,N_11440);
and U15049 (N_15049,N_8327,N_11479);
xor U15050 (N_15050,N_10585,N_11515);
nand U15051 (N_15051,N_9270,N_7111);
or U15052 (N_15052,N_11664,N_12049);
and U15053 (N_15053,N_8518,N_8507);
xnor U15054 (N_15054,N_10651,N_10785);
or U15055 (N_15055,N_8844,N_9557);
and U15056 (N_15056,N_8093,N_7057);
and U15057 (N_15057,N_8587,N_10236);
and U15058 (N_15058,N_7559,N_8063);
nor U15059 (N_15059,N_12035,N_7632);
xnor U15060 (N_15060,N_10338,N_6250);
xor U15061 (N_15061,N_10112,N_8149);
xnor U15062 (N_15062,N_11881,N_11889);
and U15063 (N_15063,N_7387,N_8513);
xnor U15064 (N_15064,N_12133,N_10404);
nor U15065 (N_15065,N_10154,N_8445);
nor U15066 (N_15066,N_12000,N_12435);
xor U15067 (N_15067,N_6951,N_8701);
and U15068 (N_15068,N_7765,N_9128);
and U15069 (N_15069,N_8762,N_11933);
or U15070 (N_15070,N_10579,N_7914);
nand U15071 (N_15071,N_8210,N_11126);
xnor U15072 (N_15072,N_9965,N_8822);
or U15073 (N_15073,N_10603,N_9416);
and U15074 (N_15074,N_9800,N_9422);
nand U15075 (N_15075,N_6351,N_11041);
or U15076 (N_15076,N_8988,N_8874);
nor U15077 (N_15077,N_11707,N_8629);
xor U15078 (N_15078,N_8300,N_12175);
xnor U15079 (N_15079,N_7071,N_7405);
or U15080 (N_15080,N_8920,N_12439);
xor U15081 (N_15081,N_11087,N_7677);
nor U15082 (N_15082,N_10508,N_7068);
and U15083 (N_15083,N_12024,N_9831);
or U15084 (N_15084,N_7902,N_9550);
nand U15085 (N_15085,N_8192,N_11174);
or U15086 (N_15086,N_10755,N_8734);
xor U15087 (N_15087,N_12354,N_10386);
nor U15088 (N_15088,N_9788,N_12329);
and U15089 (N_15089,N_10544,N_11105);
xnor U15090 (N_15090,N_8041,N_6802);
nor U15091 (N_15091,N_10161,N_7196);
nor U15092 (N_15092,N_6437,N_10564);
and U15093 (N_15093,N_10619,N_9013);
nand U15094 (N_15094,N_7715,N_6832);
and U15095 (N_15095,N_8607,N_11655);
nand U15096 (N_15096,N_7377,N_10989);
nor U15097 (N_15097,N_6448,N_7888);
and U15098 (N_15098,N_10575,N_8218);
and U15099 (N_15099,N_11830,N_7536);
nand U15100 (N_15100,N_6992,N_10234);
or U15101 (N_15101,N_6552,N_11285);
or U15102 (N_15102,N_11447,N_9760);
xor U15103 (N_15103,N_8794,N_6991);
xor U15104 (N_15104,N_10418,N_6312);
and U15105 (N_15105,N_8526,N_10584);
and U15106 (N_15106,N_12474,N_11994);
nand U15107 (N_15107,N_11089,N_10475);
and U15108 (N_15108,N_8837,N_9672);
nor U15109 (N_15109,N_6759,N_10260);
xnor U15110 (N_15110,N_7929,N_11753);
xnor U15111 (N_15111,N_7012,N_8298);
xor U15112 (N_15112,N_7745,N_9826);
nor U15113 (N_15113,N_12236,N_10568);
nand U15114 (N_15114,N_9269,N_8139);
nor U15115 (N_15115,N_10280,N_9717);
nor U15116 (N_15116,N_9735,N_12348);
nand U15117 (N_15117,N_8716,N_9668);
and U15118 (N_15118,N_11172,N_7513);
and U15119 (N_15119,N_9869,N_9404);
nand U15120 (N_15120,N_11146,N_6776);
nor U15121 (N_15121,N_10853,N_10613);
or U15122 (N_15122,N_10820,N_9942);
and U15123 (N_15123,N_6605,N_7237);
xor U15124 (N_15124,N_9448,N_10484);
nand U15125 (N_15125,N_6708,N_10412);
or U15126 (N_15126,N_7289,N_10018);
nand U15127 (N_15127,N_12101,N_10363);
or U15128 (N_15128,N_12154,N_6454);
nand U15129 (N_15129,N_6704,N_11649);
xor U15130 (N_15130,N_9181,N_11862);
nor U15131 (N_15131,N_11572,N_9215);
and U15132 (N_15132,N_10344,N_10329);
nand U15133 (N_15133,N_7615,N_12391);
and U15134 (N_15134,N_12267,N_8141);
and U15135 (N_15135,N_8922,N_12318);
or U15136 (N_15136,N_10416,N_7296);
or U15137 (N_15137,N_9815,N_9343);
nor U15138 (N_15138,N_8060,N_9053);
nand U15139 (N_15139,N_11221,N_10712);
nand U15140 (N_15140,N_10373,N_6285);
nor U15141 (N_15141,N_11652,N_10992);
and U15142 (N_15142,N_8511,N_7381);
nand U15143 (N_15143,N_6729,N_10703);
and U15144 (N_15144,N_11437,N_7644);
xor U15145 (N_15145,N_9706,N_12112);
nand U15146 (N_15146,N_7453,N_7204);
and U15147 (N_15147,N_8769,N_9015);
or U15148 (N_15148,N_11225,N_6589);
and U15149 (N_15149,N_7945,N_8350);
and U15150 (N_15150,N_6585,N_6897);
or U15151 (N_15151,N_9218,N_8274);
or U15152 (N_15152,N_11082,N_9511);
nand U15153 (N_15153,N_6451,N_9793);
nand U15154 (N_15154,N_6754,N_8016);
nor U15155 (N_15155,N_7431,N_8956);
and U15156 (N_15156,N_10986,N_11548);
and U15157 (N_15157,N_7042,N_10996);
nor U15158 (N_15158,N_11696,N_10101);
xnor U15159 (N_15159,N_8505,N_11817);
nor U15160 (N_15160,N_8334,N_6799);
nor U15161 (N_15161,N_8476,N_7910);
nand U15162 (N_15162,N_7284,N_7448);
and U15163 (N_15163,N_11247,N_9017);
and U15164 (N_15164,N_7097,N_11368);
nand U15165 (N_15165,N_9989,N_11617);
or U15166 (N_15166,N_11188,N_6277);
or U15167 (N_15167,N_7682,N_6446);
and U15168 (N_15168,N_9084,N_7668);
xor U15169 (N_15169,N_10995,N_6274);
xor U15170 (N_15170,N_8533,N_12247);
or U15171 (N_15171,N_8464,N_9213);
nor U15172 (N_15172,N_6661,N_9140);
xor U15173 (N_15173,N_8116,N_10929);
or U15174 (N_15174,N_9189,N_12025);
nor U15175 (N_15175,N_8111,N_10090);
nor U15176 (N_15176,N_7027,N_10599);
xor U15177 (N_15177,N_8457,N_9684);
and U15178 (N_15178,N_9473,N_8809);
nand U15179 (N_15179,N_11730,N_7129);
and U15180 (N_15180,N_8764,N_10870);
nor U15181 (N_15181,N_10543,N_9843);
nand U15182 (N_15182,N_10775,N_12497);
or U15183 (N_15183,N_8278,N_10970);
xnor U15184 (N_15184,N_8355,N_10425);
and U15185 (N_15185,N_7816,N_8106);
or U15186 (N_15186,N_9211,N_7489);
xor U15187 (N_15187,N_8693,N_10301);
or U15188 (N_15188,N_10616,N_12396);
xnor U15189 (N_15189,N_8876,N_6750);
or U15190 (N_15190,N_6678,N_8890);
or U15191 (N_15191,N_11248,N_7746);
nand U15192 (N_15192,N_11816,N_11290);
and U15193 (N_15193,N_9527,N_6798);
nor U15194 (N_15194,N_11754,N_8433);
and U15195 (N_15195,N_10134,N_8198);
nand U15196 (N_15196,N_11448,N_10610);
nand U15197 (N_15197,N_11756,N_10796);
nand U15198 (N_15198,N_7829,N_6304);
xnor U15199 (N_15199,N_10200,N_12459);
xnor U15200 (N_15200,N_11669,N_7859);
nand U15201 (N_15201,N_6773,N_6393);
xnor U15202 (N_15202,N_9738,N_8645);
and U15203 (N_15203,N_10224,N_7783);
xnor U15204 (N_15204,N_11604,N_10732);
or U15205 (N_15205,N_10305,N_9909);
xor U15206 (N_15206,N_10668,N_9219);
nor U15207 (N_15207,N_10181,N_10702);
xor U15208 (N_15208,N_12484,N_10284);
or U15209 (N_15209,N_11577,N_8425);
xor U15210 (N_15210,N_10105,N_10004);
nor U15211 (N_15211,N_9254,N_9743);
nor U15212 (N_15212,N_9772,N_10402);
nand U15213 (N_15213,N_7008,N_6975);
or U15214 (N_15214,N_7630,N_8521);
and U15215 (N_15215,N_11521,N_10069);
or U15216 (N_15216,N_9794,N_10036);
nand U15217 (N_15217,N_9286,N_9100);
and U15218 (N_15218,N_11311,N_9732);
nor U15219 (N_15219,N_8848,N_11634);
nand U15220 (N_15220,N_10336,N_9409);
and U15221 (N_15221,N_11727,N_8074);
or U15222 (N_15222,N_11870,N_12157);
and U15223 (N_15223,N_6706,N_7518);
nor U15224 (N_15224,N_9222,N_9026);
nand U15225 (N_15225,N_7485,N_11114);
or U15226 (N_15226,N_7662,N_12340);
xor U15227 (N_15227,N_10799,N_8602);
nand U15228 (N_15228,N_12276,N_10275);
xor U15229 (N_15229,N_7671,N_12428);
xor U15230 (N_15230,N_11839,N_9046);
nor U15231 (N_15231,N_11941,N_6308);
nor U15232 (N_15232,N_9354,N_11974);
nand U15233 (N_15233,N_8845,N_10810);
xor U15234 (N_15234,N_7171,N_11869);
or U15235 (N_15235,N_8340,N_11632);
nor U15236 (N_15236,N_10525,N_10549);
and U15237 (N_15237,N_6943,N_7953);
and U15238 (N_15238,N_9300,N_7511);
xor U15239 (N_15239,N_9283,N_8483);
nand U15240 (N_15240,N_8881,N_6949);
or U15241 (N_15241,N_7290,N_10906);
and U15242 (N_15242,N_10054,N_11639);
xnor U15243 (N_15243,N_8998,N_9085);
nand U15244 (N_15244,N_8919,N_10649);
nor U15245 (N_15245,N_11616,N_7267);
nor U15246 (N_15246,N_11708,N_8706);
or U15247 (N_15247,N_8673,N_10251);
xor U15248 (N_15248,N_7775,N_6360);
and U15249 (N_15249,N_8250,N_8096);
xor U15250 (N_15250,N_9823,N_12033);
nor U15251 (N_15251,N_9920,N_11490);
xor U15252 (N_15252,N_8212,N_6985);
xor U15253 (N_15253,N_10335,N_7343);
xor U15254 (N_15254,N_8695,N_6884);
nand U15255 (N_15255,N_8664,N_8773);
nand U15256 (N_15256,N_11798,N_8449);
or U15257 (N_15257,N_6761,N_8368);
nor U15258 (N_15258,N_7440,N_11196);
or U15259 (N_15259,N_8782,N_11179);
or U15260 (N_15260,N_11953,N_9512);
nand U15261 (N_15261,N_10728,N_10899);
nor U15262 (N_15262,N_8723,N_8698);
nor U15263 (N_15263,N_10342,N_8971);
and U15264 (N_15264,N_10753,N_12317);
nand U15265 (N_15265,N_11335,N_11271);
nor U15266 (N_15266,N_7038,N_7947);
nand U15267 (N_15267,N_10458,N_8790);
and U15268 (N_15268,N_12111,N_11631);
nor U15269 (N_15269,N_6479,N_6716);
nor U15270 (N_15270,N_7851,N_10380);
nand U15271 (N_15271,N_7878,N_11673);
nand U15272 (N_15272,N_10026,N_7264);
and U15273 (N_15273,N_6258,N_7817);
and U15274 (N_15274,N_9880,N_6513);
and U15275 (N_15275,N_12309,N_8358);
nand U15276 (N_15276,N_11977,N_6394);
and U15277 (N_15277,N_7986,N_11536);
xor U15278 (N_15278,N_6398,N_11522);
xor U15279 (N_15279,N_8007,N_7208);
nor U15280 (N_15280,N_7826,N_9087);
nor U15281 (N_15281,N_10837,N_12151);
or U15282 (N_15282,N_8330,N_10940);
or U15283 (N_15283,N_6821,N_7228);
or U15284 (N_15284,N_9555,N_8747);
nand U15285 (N_15285,N_11518,N_8413);
xor U15286 (N_15286,N_11483,N_10400);
and U15287 (N_15287,N_6755,N_8385);
or U15288 (N_15288,N_11918,N_7708);
nor U15289 (N_15289,N_9778,N_11904);
or U15290 (N_15290,N_8827,N_9899);
nand U15291 (N_15291,N_12482,N_9478);
nand U15292 (N_15292,N_11985,N_9885);
xor U15293 (N_15293,N_10474,N_8077);
and U15294 (N_15294,N_11658,N_6719);
xnor U15295 (N_15295,N_9440,N_10011);
xnor U15296 (N_15296,N_8107,N_12436);
and U15297 (N_15297,N_8867,N_7321);
nand U15298 (N_15298,N_6332,N_6667);
nor U15299 (N_15299,N_8067,N_8780);
nand U15300 (N_15300,N_9358,N_12124);
and U15301 (N_15301,N_10658,N_8767);
and U15302 (N_15302,N_7123,N_9339);
nand U15303 (N_15303,N_9004,N_12462);
nand U15304 (N_15304,N_7435,N_9090);
xnor U15305 (N_15305,N_6480,N_8904);
nor U15306 (N_15306,N_7426,N_7572);
nor U15307 (N_15307,N_9535,N_6901);
and U15308 (N_15308,N_6824,N_11410);
xnor U15309 (N_15309,N_10529,N_10840);
nor U15310 (N_15310,N_8252,N_10297);
and U15311 (N_15311,N_7046,N_7908);
or U15312 (N_15312,N_10793,N_12083);
nand U15313 (N_15313,N_9272,N_11264);
and U15314 (N_15314,N_12415,N_9324);
or U15315 (N_15315,N_7930,N_6565);
xnor U15316 (N_15316,N_9447,N_9469);
or U15317 (N_15317,N_9927,N_8926);
or U15318 (N_15318,N_12072,N_11578);
and U15319 (N_15319,N_7340,N_12369);
and U15320 (N_15320,N_10988,N_10711);
xnor U15321 (N_15321,N_12486,N_6532);
nand U15322 (N_15322,N_7593,N_6751);
xnor U15323 (N_15323,N_7402,N_12051);
nand U15324 (N_15324,N_9613,N_8884);
nor U15325 (N_15325,N_8565,N_9872);
nand U15326 (N_15326,N_10710,N_12211);
nor U15327 (N_15327,N_10984,N_11755);
xnor U15328 (N_15328,N_10673,N_8316);
nor U15329 (N_15329,N_8832,N_7475);
xnor U15330 (N_15330,N_10008,N_11884);
and U15331 (N_15331,N_10420,N_8332);
nor U15332 (N_15332,N_6401,N_11106);
xor U15333 (N_15333,N_11156,N_6861);
and U15334 (N_15334,N_12479,N_11877);
nand U15335 (N_15335,N_7809,N_6836);
or U15336 (N_15336,N_6895,N_12406);
nor U15337 (N_15337,N_7674,N_9049);
or U15338 (N_15338,N_10518,N_8654);
xnor U15339 (N_15339,N_7729,N_11422);
or U15340 (N_15340,N_6567,N_6443);
nand U15341 (N_15341,N_11738,N_6993);
and U15342 (N_15342,N_10558,N_11477);
nand U15343 (N_15343,N_11369,N_6405);
or U15344 (N_15344,N_9704,N_9790);
nand U15345 (N_15345,N_8639,N_6919);
nand U15346 (N_15346,N_8676,N_6739);
or U15347 (N_15347,N_7984,N_7278);
and U15348 (N_15348,N_11020,N_8741);
or U15349 (N_15349,N_10047,N_6764);
or U15350 (N_15350,N_7186,N_8765);
or U15351 (N_15351,N_7837,N_10934);
nand U15352 (N_15352,N_10073,N_6904);
and U15353 (N_15353,N_6529,N_8757);
nor U15354 (N_15354,N_11555,N_9273);
and U15355 (N_15355,N_7059,N_11774);
or U15356 (N_15356,N_6317,N_9118);
or U15357 (N_15357,N_8559,N_7795);
or U15358 (N_15358,N_11395,N_6262);
xnor U15359 (N_15359,N_7791,N_8720);
nand U15360 (N_15360,N_8834,N_11004);
nor U15361 (N_15361,N_12218,N_7108);
xor U15362 (N_15362,N_6733,N_10951);
or U15363 (N_15363,N_10966,N_9499);
or U15364 (N_15364,N_6499,N_10646);
or U15365 (N_15365,N_9203,N_9722);
nor U15366 (N_15366,N_9261,N_7337);
or U15367 (N_15367,N_8309,N_7219);
xor U15368 (N_15368,N_12379,N_7689);
or U15369 (N_15369,N_11861,N_7884);
or U15370 (N_15370,N_9042,N_7126);
nand U15371 (N_15371,N_10184,N_9010);
xor U15372 (N_15372,N_9274,N_8800);
or U15373 (N_15373,N_9077,N_9018);
and U15374 (N_15374,N_10688,N_8227);
xnor U15375 (N_15375,N_11677,N_9854);
nor U15376 (N_15376,N_7548,N_10770);
nand U15377 (N_15377,N_8229,N_9169);
nand U15378 (N_15378,N_11344,N_6646);
nand U15379 (N_15379,N_12328,N_11091);
nand U15380 (N_15380,N_7958,N_7909);
nand U15381 (N_15381,N_9897,N_8801);
nand U15382 (N_15382,N_10678,N_10965);
and U15383 (N_15383,N_10007,N_12115);
and U15384 (N_15384,N_10208,N_9338);
or U15385 (N_15385,N_9578,N_6878);
or U15386 (N_15386,N_11145,N_10787);
nand U15387 (N_15387,N_6265,N_10272);
or U15388 (N_15388,N_10483,N_9470);
and U15389 (N_15389,N_10057,N_8127);
nor U15390 (N_15390,N_10351,N_7299);
and U15391 (N_15391,N_9674,N_11343);
nand U15392 (N_15392,N_8170,N_9492);
xnor U15393 (N_15393,N_9667,N_7599);
nor U15394 (N_15394,N_11230,N_11894);
nor U15395 (N_15395,N_10784,N_12181);
nor U15396 (N_15396,N_7035,N_7441);
nand U15397 (N_15397,N_11452,N_9180);
nand U15398 (N_15398,N_9715,N_11762);
and U15399 (N_15399,N_9879,N_8637);
nor U15400 (N_15400,N_6541,N_6774);
or U15401 (N_15401,N_10170,N_7265);
xor U15402 (N_15402,N_11388,N_11892);
nor U15403 (N_15403,N_6556,N_12056);
or U15404 (N_15404,N_8564,N_11052);
or U15405 (N_15405,N_8493,N_8303);
nor U15406 (N_15406,N_6271,N_9262);
nand U15407 (N_15407,N_11318,N_9302);
and U15408 (N_15408,N_12249,N_10744);
or U15409 (N_15409,N_12123,N_11500);
and U15410 (N_15410,N_6584,N_6964);
xnor U15411 (N_15411,N_7007,N_10935);
nor U15412 (N_15412,N_9541,N_7019);
and U15413 (N_15413,N_10403,N_12332);
nor U15414 (N_15414,N_10089,N_12094);
and U15415 (N_15415,N_11843,N_11641);
nand U15416 (N_15416,N_9924,N_7023);
nand U15417 (N_15417,N_7338,N_10769);
nor U15418 (N_15418,N_12283,N_9256);
or U15419 (N_15419,N_7206,N_10652);
nor U15420 (N_15420,N_8270,N_10677);
or U15421 (N_15421,N_11961,N_6602);
xor U15422 (N_15422,N_10126,N_7759);
nand U15423 (N_15423,N_8258,N_7049);
nand U15424 (N_15424,N_6388,N_6491);
xor U15425 (N_15425,N_6881,N_7033);
or U15426 (N_15426,N_8254,N_11766);
or U15427 (N_15427,N_9154,N_8865);
or U15428 (N_15428,N_11913,N_6825);
or U15429 (N_15429,N_10873,N_8923);
nor U15430 (N_15430,N_11047,N_7282);
and U15431 (N_15431,N_7351,N_12434);
nand U15432 (N_15432,N_11769,N_11638);
nand U15433 (N_15433,N_7163,N_7561);
nor U15434 (N_15434,N_12179,N_10315);
nand U15435 (N_15435,N_7345,N_11476);
nor U15436 (N_15436,N_11494,N_7076);
nor U15437 (N_15437,N_9643,N_6905);
nor U15438 (N_15438,N_8231,N_9052);
and U15439 (N_15439,N_11277,N_8690);
nand U15440 (N_15440,N_6659,N_11880);
nor U15441 (N_15441,N_11524,N_9294);
or U15442 (N_15442,N_8719,N_6493);
xor U15443 (N_15443,N_9593,N_12475);
nand U15444 (N_15444,N_7283,N_11505);
nor U15445 (N_15445,N_11717,N_7717);
or U15446 (N_15446,N_10481,N_10620);
nand U15447 (N_15447,N_7067,N_7047);
nand U15448 (N_15448,N_11205,N_9803);
and U15449 (N_15449,N_10783,N_8789);
or U15450 (N_15450,N_11563,N_9619);
xor U15451 (N_15451,N_12433,N_7110);
or U15452 (N_15452,N_9589,N_11671);
and U15453 (N_15453,N_10685,N_10248);
nor U15454 (N_15454,N_10943,N_11324);
and U15455 (N_15455,N_9161,N_9390);
nor U15456 (N_15456,N_6980,N_8109);
or U15457 (N_15457,N_11951,N_8608);
nor U15458 (N_15458,N_6923,N_10176);
xor U15459 (N_15459,N_11773,N_8508);
xnor U15460 (N_15460,N_10563,N_8910);
nor U15461 (N_15461,N_12029,N_8307);
xnor U15462 (N_15462,N_9066,N_11266);
nor U15463 (N_15463,N_9658,N_10135);
nor U15464 (N_15464,N_9111,N_12294);
nor U15465 (N_15465,N_10399,N_6512);
nand U15466 (N_15466,N_9030,N_6641);
xor U15467 (N_15467,N_11270,N_7560);
xor U15468 (N_15468,N_9945,N_7470);
or U15469 (N_15469,N_8858,N_11331);
nor U15470 (N_15470,N_10626,N_10460);
nand U15471 (N_15471,N_9357,N_11276);
nor U15472 (N_15472,N_9317,N_12259);
nor U15473 (N_15473,N_8308,N_6540);
and U15474 (N_15474,N_11070,N_11718);
or U15475 (N_15475,N_7352,N_8088);
nor U15476 (N_15476,N_8732,N_9156);
nand U15477 (N_15477,N_10292,N_8415);
xor U15478 (N_15478,N_9008,N_7796);
or U15479 (N_15479,N_8617,N_11125);
and U15480 (N_15480,N_7656,N_11788);
or U15481 (N_15481,N_11510,N_11284);
nand U15482 (N_15482,N_6969,N_12233);
nand U15483 (N_15483,N_11594,N_9223);
or U15484 (N_15484,N_8658,N_9174);
nand U15485 (N_15485,N_9373,N_10364);
nor U15486 (N_15486,N_6957,N_11768);
and U15487 (N_15487,N_7339,N_8036);
xnor U15488 (N_15488,N_8942,N_6534);
nand U15489 (N_15489,N_6291,N_7641);
nand U15490 (N_15490,N_10510,N_8788);
xnor U15491 (N_15491,N_6797,N_9673);
xnor U15492 (N_15492,N_10214,N_6959);
or U15493 (N_15493,N_11002,N_10781);
and U15494 (N_15494,N_9814,N_10302);
nand U15495 (N_15495,N_11307,N_8975);
and U15496 (N_15496,N_12213,N_11923);
and U15497 (N_15497,N_11560,N_12412);
xnor U15498 (N_15498,N_8156,N_12449);
nor U15499 (N_15499,N_7105,N_9183);
nand U15500 (N_15500,N_6944,N_12074);
xor U15501 (N_15501,N_11387,N_11201);
and U15502 (N_15502,N_8692,N_10318);
or U15503 (N_15503,N_8322,N_8670);
and U15504 (N_15504,N_10551,N_8524);
nor U15505 (N_15505,N_7534,N_6833);
nand U15506 (N_15506,N_12295,N_11181);
nor U15507 (N_15507,N_10559,N_7797);
nor U15508 (N_15508,N_9521,N_9951);
or U15509 (N_15509,N_11871,N_8798);
nor U15510 (N_15510,N_11295,N_9624);
nor U15511 (N_15511,N_7726,N_11538);
xor U15512 (N_15512,N_11939,N_7955);
and U15513 (N_15513,N_10595,N_9468);
or U15514 (N_15514,N_11304,N_7303);
xor U15515 (N_15515,N_10195,N_8647);
nand U15516 (N_15516,N_7579,N_11823);
nor U15517 (N_15517,N_10468,N_11298);
nand U15518 (N_15518,N_7421,N_8775);
and U15519 (N_15519,N_9388,N_11233);
xor U15520 (N_15520,N_8441,N_7553);
xnor U15521 (N_15521,N_10754,N_10587);
nor U15522 (N_15522,N_8618,N_8295);
nand U15523 (N_15523,N_11636,N_11111);
and U15524 (N_15524,N_7389,N_12198);
xnor U15525 (N_15525,N_7675,N_8103);
nand U15526 (N_15526,N_8002,N_7642);
and U15527 (N_15527,N_7235,N_10717);
nor U15528 (N_15528,N_6696,N_11359);
or U15529 (N_15529,N_7748,N_9347);
xor U15530 (N_15530,N_6283,N_7506);
xor U15531 (N_15531,N_7487,N_8383);
and U15532 (N_15532,N_7051,N_11267);
nand U15533 (N_15533,N_8578,N_8360);
nor U15534 (N_15534,N_8122,N_8099);
and U15535 (N_15535,N_6280,N_9908);
nand U15536 (N_15536,N_8071,N_11257);
or U15537 (N_15537,N_10941,N_8983);
or U15538 (N_15538,N_10365,N_10319);
xor U15539 (N_15539,N_9786,N_9861);
and U15540 (N_15540,N_11254,N_9928);
or U15541 (N_15541,N_10814,N_7161);
xor U15542 (N_15542,N_8490,N_10177);
and U15543 (N_15543,N_8030,N_7104);
or U15544 (N_15544,N_10513,N_7584);
nor U15545 (N_15545,N_7533,N_7819);
or U15546 (N_15546,N_10357,N_10535);
and U15547 (N_15547,N_12132,N_9342);
nand U15548 (N_15548,N_8577,N_12082);
nor U15549 (N_15549,N_11624,N_10914);
nand U15550 (N_15550,N_6427,N_12352);
nand U15551 (N_15551,N_6580,N_7233);
and U15552 (N_15552,N_10247,N_7661);
or U15553 (N_15553,N_10245,N_10552);
or U15554 (N_15554,N_10804,N_7304);
xnor U15555 (N_15555,N_6546,N_12272);
nor U15556 (N_15556,N_6537,N_9581);
or U15557 (N_15557,N_11709,N_7134);
xor U15558 (N_15558,N_9129,N_10655);
or U15559 (N_15559,N_10597,N_10231);
and U15560 (N_15560,N_7383,N_12371);
nand U15561 (N_15561,N_9204,N_10700);
nor U15562 (N_15562,N_10922,N_11075);
nor U15563 (N_15563,N_8426,N_11848);
or U15564 (N_15564,N_11559,N_10002);
xnor U15565 (N_15565,N_6745,N_6475);
nand U15566 (N_15566,N_6403,N_6461);
and U15567 (N_15567,N_11236,N_7565);
and U15568 (N_15568,N_7891,N_11751);
nand U15569 (N_15569,N_6303,N_8343);
nand U15570 (N_15570,N_10451,N_11523);
xnor U15571 (N_15571,N_8268,N_10874);
nand U15572 (N_15572,N_8395,N_9537);
and U15573 (N_15573,N_6735,N_6808);
nor U15574 (N_15574,N_6828,N_12287);
xor U15575 (N_15575,N_10044,N_11394);
xnor U15576 (N_15576,N_6976,N_9208);
nor U15577 (N_15577,N_9355,N_9411);
nor U15578 (N_15578,N_11899,N_10478);
and U15579 (N_15579,N_11573,N_9344);
nand U15580 (N_15580,N_8086,N_11404);
and U15581 (N_15581,N_6679,N_10353);
nand U15582 (N_15582,N_7202,N_8917);
and U15583 (N_15583,N_6882,N_8020);
or U15584 (N_15584,N_11736,N_8655);
xor U15585 (N_15585,N_6917,N_11504);
xor U15586 (N_15586,N_7167,N_6294);
nand U15587 (N_15587,N_7522,N_10750);
and U15588 (N_15588,N_10811,N_10033);
xor U15589 (N_15589,N_9616,N_6505);
and U15590 (N_15590,N_9014,N_6801);
and U15591 (N_15591,N_8833,N_6358);
xor U15592 (N_15592,N_10624,N_11835);
xnor U15593 (N_15593,N_6807,N_8052);
or U15594 (N_15594,N_10001,N_9866);
xnor U15595 (N_15595,N_9194,N_6500);
nand U15596 (N_15596,N_7640,N_7505);
and U15597 (N_15597,N_12398,N_9167);
or U15598 (N_15598,N_7577,N_7166);
or U15599 (N_15599,N_7207,N_12373);
xor U15600 (N_15600,N_7828,N_6826);
nor U15601 (N_15601,N_10082,N_11060);
xor U15602 (N_15602,N_11030,N_9109);
and U15603 (N_15603,N_11715,N_7524);
nand U15604 (N_15604,N_9689,N_11546);
xnor U15605 (N_15605,N_7150,N_8351);
xor U15606 (N_15606,N_9039,N_10299);
xor U15607 (N_15607,N_11598,N_6738);
nand U15608 (N_15608,N_11163,N_11161);
nand U15609 (N_15609,N_8708,N_10021);
or U15610 (N_15610,N_12107,N_7904);
and U15611 (N_15611,N_9796,N_12335);
xnor U15612 (N_15612,N_10020,N_9025);
and U15613 (N_15613,N_10441,N_8245);
and U15614 (N_15614,N_9669,N_8902);
nand U15615 (N_15615,N_9605,N_12117);
nand U15616 (N_15616,N_6692,N_12325);
or U15617 (N_15617,N_7772,N_6270);
nor U15618 (N_15618,N_12076,N_11651);
xnor U15619 (N_15619,N_9191,N_11349);
nand U15620 (N_15620,N_8137,N_11988);
nor U15621 (N_15621,N_8934,N_6487);
nand U15622 (N_15622,N_8015,N_9086);
or U15623 (N_15623,N_10178,N_10670);
nand U15624 (N_15624,N_8120,N_11128);
xnor U15625 (N_15625,N_8280,N_9777);
xnor U15626 (N_15626,N_7486,N_9045);
xnor U15627 (N_15627,N_10500,N_7402);
xnor U15628 (N_15628,N_10898,N_6693);
xor U15629 (N_15629,N_8914,N_9624);
or U15630 (N_15630,N_6804,N_7969);
or U15631 (N_15631,N_9659,N_10478);
nand U15632 (N_15632,N_6929,N_11779);
xnor U15633 (N_15633,N_8435,N_11077);
and U15634 (N_15634,N_11129,N_11751);
and U15635 (N_15635,N_9425,N_6381);
or U15636 (N_15636,N_9966,N_7308);
nand U15637 (N_15637,N_9443,N_6423);
or U15638 (N_15638,N_11000,N_10538);
or U15639 (N_15639,N_9601,N_10400);
xnor U15640 (N_15640,N_11192,N_12403);
xnor U15641 (N_15641,N_6892,N_11071);
xnor U15642 (N_15642,N_7796,N_8480);
nor U15643 (N_15643,N_12096,N_9544);
xor U15644 (N_15644,N_10810,N_10400);
or U15645 (N_15645,N_7057,N_11335);
or U15646 (N_15646,N_10871,N_8708);
nor U15647 (N_15647,N_6925,N_7263);
and U15648 (N_15648,N_7411,N_8153);
or U15649 (N_15649,N_9432,N_10719);
and U15650 (N_15650,N_11016,N_9381);
or U15651 (N_15651,N_11677,N_7580);
nor U15652 (N_15652,N_11236,N_11417);
and U15653 (N_15653,N_6710,N_8539);
nor U15654 (N_15654,N_8301,N_7668);
xor U15655 (N_15655,N_11767,N_6371);
nand U15656 (N_15656,N_9307,N_9289);
nor U15657 (N_15657,N_11234,N_7164);
or U15658 (N_15658,N_6785,N_9534);
nor U15659 (N_15659,N_9311,N_9275);
xnor U15660 (N_15660,N_12202,N_11895);
and U15661 (N_15661,N_10933,N_9880);
nor U15662 (N_15662,N_7173,N_9371);
and U15663 (N_15663,N_8676,N_12204);
nor U15664 (N_15664,N_6520,N_6927);
xor U15665 (N_15665,N_10011,N_6748);
xor U15666 (N_15666,N_11510,N_6637);
nand U15667 (N_15667,N_9035,N_10782);
and U15668 (N_15668,N_8501,N_8331);
or U15669 (N_15669,N_6260,N_9747);
xnor U15670 (N_15670,N_9800,N_6563);
and U15671 (N_15671,N_7971,N_6560);
nor U15672 (N_15672,N_8907,N_12230);
nor U15673 (N_15673,N_11391,N_10292);
or U15674 (N_15674,N_9605,N_8211);
and U15675 (N_15675,N_8944,N_7930);
and U15676 (N_15676,N_9590,N_11271);
and U15677 (N_15677,N_10502,N_10856);
nand U15678 (N_15678,N_10165,N_9442);
or U15679 (N_15679,N_7884,N_7688);
or U15680 (N_15680,N_8038,N_9859);
xor U15681 (N_15681,N_7469,N_6742);
or U15682 (N_15682,N_8743,N_7582);
xor U15683 (N_15683,N_11321,N_9416);
nor U15684 (N_15684,N_9342,N_8255);
or U15685 (N_15685,N_10571,N_9847);
nor U15686 (N_15686,N_11788,N_11391);
xor U15687 (N_15687,N_10573,N_12119);
xor U15688 (N_15688,N_11853,N_11785);
and U15689 (N_15689,N_8267,N_6838);
or U15690 (N_15690,N_8669,N_8817);
xor U15691 (N_15691,N_7630,N_10212);
nor U15692 (N_15692,N_11354,N_6827);
nand U15693 (N_15693,N_8775,N_8585);
nand U15694 (N_15694,N_8436,N_8843);
and U15695 (N_15695,N_12308,N_7776);
nand U15696 (N_15696,N_11488,N_11112);
nor U15697 (N_15697,N_11884,N_7885);
and U15698 (N_15698,N_8561,N_8410);
or U15699 (N_15699,N_11448,N_12134);
nor U15700 (N_15700,N_7962,N_10216);
xnor U15701 (N_15701,N_10726,N_11541);
and U15702 (N_15702,N_9027,N_10562);
or U15703 (N_15703,N_9494,N_8177);
nor U15704 (N_15704,N_8644,N_11560);
or U15705 (N_15705,N_7884,N_6314);
and U15706 (N_15706,N_8601,N_9696);
or U15707 (N_15707,N_6317,N_12465);
xnor U15708 (N_15708,N_8118,N_10858);
and U15709 (N_15709,N_11000,N_10727);
nor U15710 (N_15710,N_6885,N_9686);
and U15711 (N_15711,N_6457,N_11563);
xnor U15712 (N_15712,N_9055,N_10543);
xor U15713 (N_15713,N_9864,N_7411);
or U15714 (N_15714,N_10826,N_8625);
or U15715 (N_15715,N_7707,N_12015);
xor U15716 (N_15716,N_8658,N_7018);
nor U15717 (N_15717,N_6596,N_8042);
nor U15718 (N_15718,N_8961,N_6396);
xnor U15719 (N_15719,N_8587,N_11886);
or U15720 (N_15720,N_12149,N_7558);
nand U15721 (N_15721,N_11537,N_11719);
xor U15722 (N_15722,N_12067,N_11475);
and U15723 (N_15723,N_7061,N_10386);
or U15724 (N_15724,N_8128,N_8500);
xor U15725 (N_15725,N_11497,N_9088);
xnor U15726 (N_15726,N_7579,N_6540);
nand U15727 (N_15727,N_8230,N_9451);
and U15728 (N_15728,N_8064,N_9784);
and U15729 (N_15729,N_11853,N_10722);
or U15730 (N_15730,N_8140,N_10278);
and U15731 (N_15731,N_10403,N_10522);
and U15732 (N_15732,N_10613,N_7361);
or U15733 (N_15733,N_10631,N_11222);
and U15734 (N_15734,N_6259,N_8842);
nand U15735 (N_15735,N_11445,N_9903);
or U15736 (N_15736,N_6896,N_10147);
or U15737 (N_15737,N_11591,N_9206);
and U15738 (N_15738,N_6509,N_8465);
and U15739 (N_15739,N_10929,N_9612);
xnor U15740 (N_15740,N_8511,N_7598);
or U15741 (N_15741,N_10532,N_12011);
nand U15742 (N_15742,N_7736,N_8860);
nor U15743 (N_15743,N_9749,N_7748);
or U15744 (N_15744,N_9082,N_6285);
nor U15745 (N_15745,N_12477,N_6708);
and U15746 (N_15746,N_7512,N_9426);
or U15747 (N_15747,N_9699,N_11320);
and U15748 (N_15748,N_12193,N_7562);
or U15749 (N_15749,N_12020,N_6414);
or U15750 (N_15750,N_10469,N_8609);
xor U15751 (N_15751,N_10001,N_8194);
and U15752 (N_15752,N_7816,N_6283);
xnor U15753 (N_15753,N_7067,N_11460);
and U15754 (N_15754,N_11131,N_11247);
nor U15755 (N_15755,N_11348,N_10668);
xnor U15756 (N_15756,N_6706,N_7143);
nand U15757 (N_15757,N_8670,N_6926);
and U15758 (N_15758,N_11874,N_9373);
nand U15759 (N_15759,N_10799,N_11132);
xnor U15760 (N_15760,N_12208,N_10583);
xor U15761 (N_15761,N_11253,N_10386);
nand U15762 (N_15762,N_11812,N_10374);
or U15763 (N_15763,N_7261,N_12335);
nor U15764 (N_15764,N_6884,N_8605);
xnor U15765 (N_15765,N_7544,N_12164);
xnor U15766 (N_15766,N_9009,N_11839);
nor U15767 (N_15767,N_7798,N_10327);
nor U15768 (N_15768,N_6915,N_10083);
and U15769 (N_15769,N_11834,N_9518);
nand U15770 (N_15770,N_11071,N_9969);
nor U15771 (N_15771,N_11771,N_9438);
xor U15772 (N_15772,N_9065,N_11864);
xor U15773 (N_15773,N_8394,N_9864);
nor U15774 (N_15774,N_8086,N_7723);
xor U15775 (N_15775,N_6673,N_9538);
and U15776 (N_15776,N_10124,N_6344);
xor U15777 (N_15777,N_9399,N_7362);
and U15778 (N_15778,N_6463,N_11957);
xor U15779 (N_15779,N_6404,N_9221);
or U15780 (N_15780,N_10279,N_6980);
and U15781 (N_15781,N_6530,N_11166);
and U15782 (N_15782,N_8198,N_8625);
nand U15783 (N_15783,N_11457,N_8377);
and U15784 (N_15784,N_10012,N_11482);
xor U15785 (N_15785,N_6882,N_7069);
xor U15786 (N_15786,N_7578,N_9973);
nor U15787 (N_15787,N_9640,N_11178);
and U15788 (N_15788,N_10404,N_9417);
xnor U15789 (N_15789,N_6744,N_7127);
xnor U15790 (N_15790,N_9030,N_11339);
nor U15791 (N_15791,N_6452,N_7786);
and U15792 (N_15792,N_11922,N_7704);
or U15793 (N_15793,N_7960,N_7407);
or U15794 (N_15794,N_7228,N_7809);
or U15795 (N_15795,N_8738,N_11241);
and U15796 (N_15796,N_8518,N_8241);
or U15797 (N_15797,N_8330,N_6642);
and U15798 (N_15798,N_6563,N_8679);
xor U15799 (N_15799,N_10181,N_6255);
nor U15800 (N_15800,N_10330,N_6643);
nand U15801 (N_15801,N_7684,N_6954);
nor U15802 (N_15802,N_12086,N_11071);
xor U15803 (N_15803,N_10988,N_7648);
xnor U15804 (N_15804,N_8452,N_8878);
or U15805 (N_15805,N_7976,N_6600);
xnor U15806 (N_15806,N_8036,N_10805);
nor U15807 (N_15807,N_6689,N_11262);
or U15808 (N_15808,N_9162,N_12298);
nor U15809 (N_15809,N_7762,N_7823);
or U15810 (N_15810,N_10901,N_10611);
or U15811 (N_15811,N_9283,N_7808);
xnor U15812 (N_15812,N_7065,N_12008);
xnor U15813 (N_15813,N_7962,N_6281);
and U15814 (N_15814,N_11419,N_10710);
and U15815 (N_15815,N_7768,N_11139);
xor U15816 (N_15816,N_9062,N_6968);
or U15817 (N_15817,N_10185,N_8392);
nand U15818 (N_15818,N_9736,N_7864);
or U15819 (N_15819,N_9156,N_10579);
nand U15820 (N_15820,N_6582,N_9173);
nand U15821 (N_15821,N_9105,N_7502);
nor U15822 (N_15822,N_10237,N_12484);
or U15823 (N_15823,N_11022,N_12204);
or U15824 (N_15824,N_11821,N_7186);
nor U15825 (N_15825,N_7109,N_6967);
nor U15826 (N_15826,N_11529,N_10874);
xor U15827 (N_15827,N_7352,N_11051);
nor U15828 (N_15828,N_9212,N_11881);
nor U15829 (N_15829,N_9426,N_10055);
or U15830 (N_15830,N_8844,N_8269);
nand U15831 (N_15831,N_8371,N_7955);
and U15832 (N_15832,N_11202,N_8223);
nor U15833 (N_15833,N_7275,N_11549);
nor U15834 (N_15834,N_8497,N_6856);
or U15835 (N_15835,N_10483,N_7449);
and U15836 (N_15836,N_8930,N_8531);
xor U15837 (N_15837,N_11534,N_6421);
nand U15838 (N_15838,N_9035,N_10106);
and U15839 (N_15839,N_6319,N_9519);
nand U15840 (N_15840,N_11682,N_9830);
xnor U15841 (N_15841,N_7410,N_11669);
nor U15842 (N_15842,N_12281,N_7125);
or U15843 (N_15843,N_7959,N_6522);
xor U15844 (N_15844,N_6594,N_10638);
nand U15845 (N_15845,N_7717,N_8307);
nand U15846 (N_15846,N_9100,N_10035);
and U15847 (N_15847,N_8610,N_8618);
and U15848 (N_15848,N_9805,N_8995);
nand U15849 (N_15849,N_6330,N_11606);
and U15850 (N_15850,N_6665,N_10233);
or U15851 (N_15851,N_7594,N_10248);
xor U15852 (N_15852,N_7908,N_10004);
nor U15853 (N_15853,N_10304,N_8316);
or U15854 (N_15854,N_10360,N_11851);
and U15855 (N_15855,N_10074,N_6440);
nand U15856 (N_15856,N_9721,N_6524);
nand U15857 (N_15857,N_7926,N_7937);
or U15858 (N_15858,N_9650,N_11803);
xor U15859 (N_15859,N_12185,N_8277);
nor U15860 (N_15860,N_7612,N_8154);
or U15861 (N_15861,N_11927,N_10823);
and U15862 (N_15862,N_9129,N_8624);
or U15863 (N_15863,N_8613,N_7951);
or U15864 (N_15864,N_12296,N_10909);
nand U15865 (N_15865,N_10799,N_7092);
and U15866 (N_15866,N_8112,N_8300);
nand U15867 (N_15867,N_8353,N_6612);
xor U15868 (N_15868,N_9221,N_11884);
nand U15869 (N_15869,N_9613,N_11079);
and U15870 (N_15870,N_7140,N_12121);
xnor U15871 (N_15871,N_6813,N_8256);
xnor U15872 (N_15872,N_11389,N_7061);
nor U15873 (N_15873,N_10990,N_10157);
xnor U15874 (N_15874,N_8532,N_11097);
nand U15875 (N_15875,N_8560,N_7104);
nor U15876 (N_15876,N_9874,N_9560);
xnor U15877 (N_15877,N_6927,N_11952);
xor U15878 (N_15878,N_8084,N_8369);
and U15879 (N_15879,N_12173,N_9292);
or U15880 (N_15880,N_8508,N_6755);
xor U15881 (N_15881,N_8895,N_10952);
nor U15882 (N_15882,N_8389,N_7382);
nor U15883 (N_15883,N_8660,N_11665);
nand U15884 (N_15884,N_7320,N_11811);
nor U15885 (N_15885,N_11659,N_8902);
nor U15886 (N_15886,N_8936,N_8299);
and U15887 (N_15887,N_10818,N_6794);
xor U15888 (N_15888,N_9924,N_12380);
xor U15889 (N_15889,N_8606,N_9328);
and U15890 (N_15890,N_12410,N_6326);
xor U15891 (N_15891,N_11723,N_10398);
xnor U15892 (N_15892,N_11868,N_10759);
nor U15893 (N_15893,N_6887,N_10353);
nor U15894 (N_15894,N_6823,N_6547);
xnor U15895 (N_15895,N_9365,N_10815);
xor U15896 (N_15896,N_7997,N_9591);
nand U15897 (N_15897,N_10428,N_11816);
or U15898 (N_15898,N_7913,N_8987);
and U15899 (N_15899,N_10474,N_9480);
or U15900 (N_15900,N_8598,N_7639);
and U15901 (N_15901,N_8387,N_10500);
nand U15902 (N_15902,N_7942,N_12025);
nand U15903 (N_15903,N_8423,N_8244);
nor U15904 (N_15904,N_6668,N_9564);
xnor U15905 (N_15905,N_6821,N_9557);
nor U15906 (N_15906,N_11740,N_9059);
or U15907 (N_15907,N_7945,N_10333);
nand U15908 (N_15908,N_7206,N_7054);
nand U15909 (N_15909,N_11078,N_11704);
nand U15910 (N_15910,N_11182,N_6671);
or U15911 (N_15911,N_7871,N_10324);
xnor U15912 (N_15912,N_6295,N_8150);
nor U15913 (N_15913,N_9181,N_6833);
or U15914 (N_15914,N_10145,N_11532);
xnor U15915 (N_15915,N_8363,N_6746);
or U15916 (N_15916,N_8653,N_12191);
nor U15917 (N_15917,N_7798,N_7424);
and U15918 (N_15918,N_11966,N_12144);
and U15919 (N_15919,N_10155,N_7751);
xnor U15920 (N_15920,N_8844,N_6539);
xor U15921 (N_15921,N_9342,N_10082);
nor U15922 (N_15922,N_6747,N_10181);
xnor U15923 (N_15923,N_7500,N_8908);
or U15924 (N_15924,N_10321,N_10455);
nor U15925 (N_15925,N_9626,N_10851);
nand U15926 (N_15926,N_8986,N_10978);
or U15927 (N_15927,N_7553,N_10100);
nand U15928 (N_15928,N_8237,N_6962);
and U15929 (N_15929,N_9388,N_12022);
nor U15930 (N_15930,N_9388,N_8395);
xor U15931 (N_15931,N_8786,N_10233);
nand U15932 (N_15932,N_7164,N_9934);
xnor U15933 (N_15933,N_10910,N_10545);
and U15934 (N_15934,N_10581,N_6995);
or U15935 (N_15935,N_10831,N_9472);
nor U15936 (N_15936,N_10528,N_10395);
nand U15937 (N_15937,N_8234,N_11696);
and U15938 (N_15938,N_7431,N_7326);
xor U15939 (N_15939,N_8704,N_9114);
nand U15940 (N_15940,N_7225,N_11990);
and U15941 (N_15941,N_10842,N_10027);
nand U15942 (N_15942,N_11294,N_11904);
xor U15943 (N_15943,N_10607,N_11889);
nand U15944 (N_15944,N_9669,N_8464);
nand U15945 (N_15945,N_10352,N_10055);
xor U15946 (N_15946,N_8184,N_11187);
or U15947 (N_15947,N_8434,N_9285);
nor U15948 (N_15948,N_9899,N_9010);
and U15949 (N_15949,N_8443,N_9838);
nor U15950 (N_15950,N_7336,N_7165);
and U15951 (N_15951,N_10007,N_6333);
nand U15952 (N_15952,N_12172,N_6816);
and U15953 (N_15953,N_9253,N_6665);
and U15954 (N_15954,N_11338,N_11210);
or U15955 (N_15955,N_10762,N_10883);
and U15956 (N_15956,N_6681,N_9350);
and U15957 (N_15957,N_9640,N_9976);
or U15958 (N_15958,N_8974,N_11051);
and U15959 (N_15959,N_6949,N_11291);
and U15960 (N_15960,N_6393,N_10069);
and U15961 (N_15961,N_10517,N_11957);
and U15962 (N_15962,N_10364,N_9246);
nor U15963 (N_15963,N_8028,N_10687);
nor U15964 (N_15964,N_9538,N_7190);
nand U15965 (N_15965,N_11312,N_7372);
nor U15966 (N_15966,N_9521,N_6364);
or U15967 (N_15967,N_8845,N_10351);
and U15968 (N_15968,N_11705,N_6380);
or U15969 (N_15969,N_8848,N_7264);
xor U15970 (N_15970,N_6901,N_9244);
xnor U15971 (N_15971,N_12334,N_12177);
nor U15972 (N_15972,N_12295,N_8237);
nand U15973 (N_15973,N_9088,N_7592);
xnor U15974 (N_15974,N_7717,N_7559);
nand U15975 (N_15975,N_9186,N_11313);
nor U15976 (N_15976,N_9858,N_7702);
nand U15977 (N_15977,N_10860,N_8594);
nor U15978 (N_15978,N_7365,N_8528);
xor U15979 (N_15979,N_12268,N_10541);
or U15980 (N_15980,N_8575,N_6814);
xor U15981 (N_15981,N_11051,N_9061);
xnor U15982 (N_15982,N_6818,N_9005);
and U15983 (N_15983,N_11304,N_8334);
nand U15984 (N_15984,N_6464,N_10960);
nor U15985 (N_15985,N_7646,N_7444);
xnor U15986 (N_15986,N_8179,N_8259);
xor U15987 (N_15987,N_6311,N_11637);
nor U15988 (N_15988,N_12348,N_8504);
or U15989 (N_15989,N_7483,N_6647);
or U15990 (N_15990,N_6338,N_9434);
or U15991 (N_15991,N_7091,N_11252);
or U15992 (N_15992,N_9421,N_10092);
xor U15993 (N_15993,N_8403,N_7528);
or U15994 (N_15994,N_7711,N_8744);
xor U15995 (N_15995,N_8807,N_8691);
or U15996 (N_15996,N_12036,N_11433);
nand U15997 (N_15997,N_6648,N_11815);
nor U15998 (N_15998,N_8443,N_8653);
or U15999 (N_15999,N_9146,N_9415);
and U16000 (N_16000,N_9441,N_7188);
nand U16001 (N_16001,N_12063,N_8465);
and U16002 (N_16002,N_12000,N_8383);
and U16003 (N_16003,N_6564,N_8016);
nor U16004 (N_16004,N_10915,N_7912);
and U16005 (N_16005,N_10916,N_6821);
nand U16006 (N_16006,N_11590,N_6550);
nand U16007 (N_16007,N_9622,N_6428);
nor U16008 (N_16008,N_7033,N_9465);
nor U16009 (N_16009,N_10582,N_8789);
or U16010 (N_16010,N_12131,N_11152);
or U16011 (N_16011,N_9424,N_10756);
or U16012 (N_16012,N_10844,N_12346);
xnor U16013 (N_16013,N_7398,N_7908);
xnor U16014 (N_16014,N_11463,N_7793);
or U16015 (N_16015,N_10753,N_9732);
nand U16016 (N_16016,N_9310,N_12433);
nand U16017 (N_16017,N_8832,N_6285);
xnor U16018 (N_16018,N_10858,N_10097);
nand U16019 (N_16019,N_9454,N_12174);
nand U16020 (N_16020,N_7571,N_8149);
nor U16021 (N_16021,N_7174,N_6776);
nor U16022 (N_16022,N_10816,N_10109);
nor U16023 (N_16023,N_8648,N_9582);
and U16024 (N_16024,N_11289,N_8406);
nor U16025 (N_16025,N_6595,N_10903);
nand U16026 (N_16026,N_7201,N_6282);
xor U16027 (N_16027,N_7652,N_12400);
and U16028 (N_16028,N_7111,N_10713);
nand U16029 (N_16029,N_10200,N_7503);
nand U16030 (N_16030,N_10050,N_10954);
and U16031 (N_16031,N_9990,N_11162);
nand U16032 (N_16032,N_11456,N_11481);
or U16033 (N_16033,N_10540,N_11343);
xor U16034 (N_16034,N_7403,N_9258);
and U16035 (N_16035,N_7909,N_11621);
nor U16036 (N_16036,N_10661,N_11473);
or U16037 (N_16037,N_7400,N_7423);
nand U16038 (N_16038,N_6901,N_8650);
and U16039 (N_16039,N_12066,N_12317);
or U16040 (N_16040,N_6421,N_9493);
xnor U16041 (N_16041,N_11903,N_7237);
xnor U16042 (N_16042,N_11983,N_7755);
nand U16043 (N_16043,N_9378,N_6459);
nand U16044 (N_16044,N_10520,N_6973);
and U16045 (N_16045,N_8876,N_6295);
xor U16046 (N_16046,N_6704,N_8851);
xor U16047 (N_16047,N_10193,N_9648);
or U16048 (N_16048,N_10354,N_9607);
and U16049 (N_16049,N_10811,N_8505);
nand U16050 (N_16050,N_10283,N_6870);
nand U16051 (N_16051,N_9067,N_8295);
or U16052 (N_16052,N_10351,N_12214);
and U16053 (N_16053,N_9397,N_11368);
nand U16054 (N_16054,N_11082,N_10027);
and U16055 (N_16055,N_11720,N_10561);
nor U16056 (N_16056,N_9820,N_6893);
or U16057 (N_16057,N_8157,N_7379);
and U16058 (N_16058,N_9008,N_9569);
xor U16059 (N_16059,N_9012,N_10081);
xnor U16060 (N_16060,N_11679,N_11727);
and U16061 (N_16061,N_7684,N_7811);
and U16062 (N_16062,N_12177,N_7390);
nor U16063 (N_16063,N_11742,N_7351);
nand U16064 (N_16064,N_10881,N_9749);
nor U16065 (N_16065,N_6492,N_7681);
or U16066 (N_16066,N_11772,N_9075);
nand U16067 (N_16067,N_11691,N_10705);
nor U16068 (N_16068,N_7891,N_9478);
nor U16069 (N_16069,N_7048,N_9539);
xnor U16070 (N_16070,N_11528,N_9158);
xnor U16071 (N_16071,N_11888,N_7688);
or U16072 (N_16072,N_7201,N_8357);
xnor U16073 (N_16073,N_10334,N_6456);
or U16074 (N_16074,N_7633,N_6536);
or U16075 (N_16075,N_9052,N_8263);
nand U16076 (N_16076,N_7519,N_8096);
and U16077 (N_16077,N_7084,N_6580);
or U16078 (N_16078,N_7435,N_9739);
nand U16079 (N_16079,N_9023,N_9248);
nand U16080 (N_16080,N_12157,N_8930);
nand U16081 (N_16081,N_10558,N_8531);
nand U16082 (N_16082,N_8614,N_7409);
xor U16083 (N_16083,N_8422,N_7822);
nand U16084 (N_16084,N_8692,N_7199);
and U16085 (N_16085,N_11877,N_8568);
or U16086 (N_16086,N_10125,N_12177);
and U16087 (N_16087,N_11003,N_9765);
nor U16088 (N_16088,N_9012,N_7539);
and U16089 (N_16089,N_6662,N_12324);
xnor U16090 (N_16090,N_10006,N_10654);
or U16091 (N_16091,N_10678,N_9435);
nor U16092 (N_16092,N_11013,N_7668);
and U16093 (N_16093,N_10332,N_10222);
and U16094 (N_16094,N_6622,N_7342);
and U16095 (N_16095,N_6568,N_9451);
or U16096 (N_16096,N_7347,N_11120);
nor U16097 (N_16097,N_6736,N_6281);
xor U16098 (N_16098,N_7979,N_8951);
or U16099 (N_16099,N_6683,N_7381);
or U16100 (N_16100,N_10592,N_10210);
or U16101 (N_16101,N_11438,N_12214);
xor U16102 (N_16102,N_11583,N_7229);
or U16103 (N_16103,N_9929,N_9704);
nor U16104 (N_16104,N_8031,N_7128);
nor U16105 (N_16105,N_9270,N_9582);
nand U16106 (N_16106,N_12078,N_9062);
or U16107 (N_16107,N_10459,N_7377);
or U16108 (N_16108,N_10138,N_11730);
nand U16109 (N_16109,N_12481,N_7294);
or U16110 (N_16110,N_10427,N_7716);
and U16111 (N_16111,N_6792,N_12494);
nor U16112 (N_16112,N_9956,N_9367);
nor U16113 (N_16113,N_11157,N_8305);
nor U16114 (N_16114,N_7969,N_8796);
xnor U16115 (N_16115,N_10541,N_8746);
nand U16116 (N_16116,N_9446,N_12073);
xor U16117 (N_16117,N_8196,N_7496);
or U16118 (N_16118,N_9855,N_9820);
and U16119 (N_16119,N_12380,N_7574);
nor U16120 (N_16120,N_7805,N_6954);
or U16121 (N_16121,N_6419,N_10134);
xnor U16122 (N_16122,N_11946,N_7686);
nor U16123 (N_16123,N_6984,N_7254);
nand U16124 (N_16124,N_9772,N_9143);
nand U16125 (N_16125,N_10627,N_11339);
and U16126 (N_16126,N_8733,N_11615);
xor U16127 (N_16127,N_11823,N_8036);
nand U16128 (N_16128,N_12350,N_11610);
and U16129 (N_16129,N_6731,N_10971);
and U16130 (N_16130,N_9813,N_10435);
or U16131 (N_16131,N_6730,N_10797);
nor U16132 (N_16132,N_6747,N_11676);
xor U16133 (N_16133,N_10517,N_7720);
nor U16134 (N_16134,N_7698,N_9023);
xor U16135 (N_16135,N_11439,N_12284);
and U16136 (N_16136,N_7792,N_11684);
and U16137 (N_16137,N_12359,N_7597);
or U16138 (N_16138,N_7745,N_9852);
or U16139 (N_16139,N_11183,N_11251);
and U16140 (N_16140,N_8816,N_12252);
xnor U16141 (N_16141,N_8520,N_7000);
nor U16142 (N_16142,N_8723,N_7767);
xnor U16143 (N_16143,N_11557,N_7860);
xor U16144 (N_16144,N_6562,N_9366);
and U16145 (N_16145,N_8589,N_9343);
or U16146 (N_16146,N_11561,N_7594);
xor U16147 (N_16147,N_9720,N_7529);
or U16148 (N_16148,N_10357,N_11649);
nand U16149 (N_16149,N_6915,N_11491);
and U16150 (N_16150,N_11790,N_11874);
xnor U16151 (N_16151,N_8578,N_9166);
nand U16152 (N_16152,N_9431,N_11140);
and U16153 (N_16153,N_7416,N_6313);
nand U16154 (N_16154,N_11598,N_7013);
nand U16155 (N_16155,N_12347,N_7336);
and U16156 (N_16156,N_8764,N_7521);
or U16157 (N_16157,N_7267,N_8670);
nor U16158 (N_16158,N_9109,N_7623);
or U16159 (N_16159,N_7777,N_12145);
nor U16160 (N_16160,N_8895,N_6411);
and U16161 (N_16161,N_8972,N_11830);
nand U16162 (N_16162,N_10134,N_6971);
and U16163 (N_16163,N_11647,N_12094);
xor U16164 (N_16164,N_11228,N_7657);
and U16165 (N_16165,N_11312,N_8356);
and U16166 (N_16166,N_11097,N_8331);
xor U16167 (N_16167,N_8580,N_9044);
and U16168 (N_16168,N_10517,N_6399);
or U16169 (N_16169,N_6626,N_10526);
nor U16170 (N_16170,N_10014,N_6735);
nor U16171 (N_16171,N_11858,N_10951);
and U16172 (N_16172,N_7582,N_11289);
or U16173 (N_16173,N_10124,N_10623);
or U16174 (N_16174,N_6427,N_9717);
nor U16175 (N_16175,N_12077,N_8778);
nand U16176 (N_16176,N_9017,N_11668);
and U16177 (N_16177,N_12476,N_11771);
nand U16178 (N_16178,N_7490,N_9324);
nand U16179 (N_16179,N_6912,N_10547);
or U16180 (N_16180,N_10842,N_7255);
or U16181 (N_16181,N_10548,N_12373);
nand U16182 (N_16182,N_10058,N_12076);
xnor U16183 (N_16183,N_7752,N_11290);
and U16184 (N_16184,N_9741,N_7391);
nand U16185 (N_16185,N_10202,N_7161);
nor U16186 (N_16186,N_10742,N_7644);
nand U16187 (N_16187,N_10741,N_9604);
or U16188 (N_16188,N_7597,N_10936);
or U16189 (N_16189,N_11048,N_12366);
nor U16190 (N_16190,N_8416,N_6827);
or U16191 (N_16191,N_10254,N_9401);
nand U16192 (N_16192,N_11415,N_11993);
and U16193 (N_16193,N_9900,N_10228);
xnor U16194 (N_16194,N_12474,N_9578);
nand U16195 (N_16195,N_10848,N_12118);
or U16196 (N_16196,N_7715,N_11901);
and U16197 (N_16197,N_12100,N_8838);
and U16198 (N_16198,N_9633,N_6417);
nand U16199 (N_16199,N_11454,N_9299);
and U16200 (N_16200,N_11458,N_8171);
nor U16201 (N_16201,N_11858,N_9708);
xor U16202 (N_16202,N_10963,N_10443);
and U16203 (N_16203,N_11153,N_11023);
nor U16204 (N_16204,N_7225,N_7288);
nand U16205 (N_16205,N_9448,N_10197);
nor U16206 (N_16206,N_7293,N_10087);
nor U16207 (N_16207,N_8498,N_11975);
xor U16208 (N_16208,N_11472,N_10289);
nand U16209 (N_16209,N_8693,N_8832);
xnor U16210 (N_16210,N_7711,N_12208);
xor U16211 (N_16211,N_6622,N_10429);
xnor U16212 (N_16212,N_11801,N_9375);
or U16213 (N_16213,N_8769,N_9545);
nor U16214 (N_16214,N_11109,N_6459);
nand U16215 (N_16215,N_12429,N_10442);
or U16216 (N_16216,N_12434,N_11071);
xor U16217 (N_16217,N_7426,N_12033);
xor U16218 (N_16218,N_8445,N_8013);
or U16219 (N_16219,N_12281,N_7406);
nand U16220 (N_16220,N_9873,N_10264);
nand U16221 (N_16221,N_10151,N_11748);
xor U16222 (N_16222,N_9078,N_6638);
nand U16223 (N_16223,N_8204,N_11562);
xor U16224 (N_16224,N_9396,N_12065);
or U16225 (N_16225,N_9317,N_11720);
nand U16226 (N_16226,N_9304,N_7959);
xnor U16227 (N_16227,N_6443,N_9397);
nand U16228 (N_16228,N_7624,N_8854);
nor U16229 (N_16229,N_7298,N_9936);
or U16230 (N_16230,N_11036,N_7372);
nand U16231 (N_16231,N_8718,N_11854);
nand U16232 (N_16232,N_11394,N_12114);
or U16233 (N_16233,N_9834,N_7868);
nor U16234 (N_16234,N_7488,N_12149);
and U16235 (N_16235,N_6780,N_10804);
or U16236 (N_16236,N_6992,N_12017);
nor U16237 (N_16237,N_10430,N_7955);
nand U16238 (N_16238,N_6410,N_9588);
or U16239 (N_16239,N_8004,N_11291);
nor U16240 (N_16240,N_9217,N_11432);
and U16241 (N_16241,N_7526,N_11546);
and U16242 (N_16242,N_8782,N_8009);
nand U16243 (N_16243,N_11594,N_10218);
xnor U16244 (N_16244,N_9581,N_8638);
nand U16245 (N_16245,N_10331,N_8921);
nand U16246 (N_16246,N_7058,N_7705);
nand U16247 (N_16247,N_11596,N_8557);
nor U16248 (N_16248,N_7104,N_6492);
nor U16249 (N_16249,N_10415,N_11214);
xor U16250 (N_16250,N_11367,N_11929);
xnor U16251 (N_16251,N_7190,N_7566);
or U16252 (N_16252,N_8911,N_7125);
and U16253 (N_16253,N_8019,N_8571);
nand U16254 (N_16254,N_8555,N_10023);
nor U16255 (N_16255,N_8255,N_9577);
and U16256 (N_16256,N_12176,N_12434);
nand U16257 (N_16257,N_9287,N_8432);
xor U16258 (N_16258,N_6592,N_11659);
xnor U16259 (N_16259,N_10544,N_6450);
xnor U16260 (N_16260,N_11347,N_10807);
nor U16261 (N_16261,N_12102,N_6310);
nor U16262 (N_16262,N_10957,N_7733);
nand U16263 (N_16263,N_10928,N_12193);
nand U16264 (N_16264,N_10282,N_9373);
or U16265 (N_16265,N_6855,N_11910);
nor U16266 (N_16266,N_8090,N_10171);
nand U16267 (N_16267,N_6563,N_11949);
nand U16268 (N_16268,N_10380,N_6544);
nor U16269 (N_16269,N_7940,N_7227);
xnor U16270 (N_16270,N_11615,N_11344);
xnor U16271 (N_16271,N_11063,N_11034);
nand U16272 (N_16272,N_10558,N_10984);
nor U16273 (N_16273,N_11411,N_8835);
or U16274 (N_16274,N_7033,N_8750);
or U16275 (N_16275,N_9419,N_9470);
nor U16276 (N_16276,N_8320,N_10927);
xnor U16277 (N_16277,N_11355,N_11966);
nor U16278 (N_16278,N_11098,N_10398);
xnor U16279 (N_16279,N_9545,N_8827);
nor U16280 (N_16280,N_7886,N_11513);
nand U16281 (N_16281,N_9338,N_10833);
and U16282 (N_16282,N_8522,N_11166);
or U16283 (N_16283,N_7173,N_11631);
or U16284 (N_16284,N_9637,N_7272);
nor U16285 (N_16285,N_9194,N_6678);
xor U16286 (N_16286,N_11636,N_8982);
xnor U16287 (N_16287,N_9534,N_9727);
or U16288 (N_16288,N_9500,N_8447);
or U16289 (N_16289,N_12228,N_11915);
or U16290 (N_16290,N_9146,N_6292);
nor U16291 (N_16291,N_8708,N_8392);
nor U16292 (N_16292,N_11600,N_7403);
nor U16293 (N_16293,N_6986,N_9245);
nand U16294 (N_16294,N_8624,N_6994);
or U16295 (N_16295,N_10642,N_11647);
or U16296 (N_16296,N_9081,N_7907);
or U16297 (N_16297,N_6739,N_11354);
or U16298 (N_16298,N_6461,N_11450);
xor U16299 (N_16299,N_10577,N_9167);
nand U16300 (N_16300,N_9745,N_10530);
xor U16301 (N_16301,N_7039,N_7101);
xor U16302 (N_16302,N_11897,N_11569);
or U16303 (N_16303,N_6371,N_11382);
nand U16304 (N_16304,N_8609,N_11399);
nand U16305 (N_16305,N_6758,N_12263);
nand U16306 (N_16306,N_10692,N_11403);
and U16307 (N_16307,N_6565,N_10176);
xor U16308 (N_16308,N_10872,N_7035);
or U16309 (N_16309,N_7853,N_11631);
nand U16310 (N_16310,N_8957,N_12423);
nand U16311 (N_16311,N_7817,N_11223);
nand U16312 (N_16312,N_11383,N_7694);
or U16313 (N_16313,N_11907,N_6530);
or U16314 (N_16314,N_10590,N_11997);
nor U16315 (N_16315,N_12403,N_8985);
nand U16316 (N_16316,N_12106,N_10407);
nand U16317 (N_16317,N_9167,N_10077);
or U16318 (N_16318,N_10751,N_10215);
or U16319 (N_16319,N_9819,N_7651);
xor U16320 (N_16320,N_12149,N_10241);
xor U16321 (N_16321,N_10303,N_10804);
nor U16322 (N_16322,N_9183,N_6888);
or U16323 (N_16323,N_7831,N_10726);
nor U16324 (N_16324,N_9722,N_11633);
nand U16325 (N_16325,N_7154,N_12358);
nor U16326 (N_16326,N_7607,N_7426);
nand U16327 (N_16327,N_10141,N_11622);
nor U16328 (N_16328,N_10943,N_12338);
or U16329 (N_16329,N_9658,N_7479);
nor U16330 (N_16330,N_9217,N_6415);
nand U16331 (N_16331,N_7599,N_6482);
and U16332 (N_16332,N_8486,N_11676);
nand U16333 (N_16333,N_10329,N_9093);
and U16334 (N_16334,N_9068,N_11939);
nand U16335 (N_16335,N_7246,N_11256);
xnor U16336 (N_16336,N_8391,N_11018);
and U16337 (N_16337,N_6713,N_10753);
xnor U16338 (N_16338,N_6329,N_10340);
and U16339 (N_16339,N_10811,N_6927);
or U16340 (N_16340,N_11076,N_6282);
nor U16341 (N_16341,N_9401,N_8357);
nand U16342 (N_16342,N_9937,N_10771);
nand U16343 (N_16343,N_11957,N_8462);
or U16344 (N_16344,N_9387,N_8199);
or U16345 (N_16345,N_11830,N_12431);
nand U16346 (N_16346,N_10568,N_10903);
nand U16347 (N_16347,N_10402,N_9334);
and U16348 (N_16348,N_8381,N_10008);
nand U16349 (N_16349,N_9144,N_7394);
and U16350 (N_16350,N_6685,N_12442);
and U16351 (N_16351,N_12441,N_10217);
or U16352 (N_16352,N_10022,N_6970);
xor U16353 (N_16353,N_11311,N_7375);
nand U16354 (N_16354,N_6682,N_9272);
nand U16355 (N_16355,N_7590,N_12090);
nand U16356 (N_16356,N_8291,N_10546);
xnor U16357 (N_16357,N_8031,N_10060);
or U16358 (N_16358,N_9412,N_7392);
nand U16359 (N_16359,N_7179,N_11117);
or U16360 (N_16360,N_9412,N_8253);
xnor U16361 (N_16361,N_8206,N_10058);
nand U16362 (N_16362,N_10486,N_12129);
nor U16363 (N_16363,N_11665,N_6468);
and U16364 (N_16364,N_8667,N_9098);
nand U16365 (N_16365,N_7631,N_6491);
or U16366 (N_16366,N_7165,N_10142);
nor U16367 (N_16367,N_8585,N_8001);
nor U16368 (N_16368,N_6314,N_10605);
or U16369 (N_16369,N_7980,N_8780);
and U16370 (N_16370,N_10727,N_10227);
nand U16371 (N_16371,N_9155,N_10290);
xor U16372 (N_16372,N_9574,N_9463);
xor U16373 (N_16373,N_8354,N_10420);
xor U16374 (N_16374,N_7450,N_9302);
nor U16375 (N_16375,N_11093,N_12391);
and U16376 (N_16376,N_7518,N_12297);
and U16377 (N_16377,N_6258,N_10055);
and U16378 (N_16378,N_10351,N_6510);
nand U16379 (N_16379,N_11714,N_7460);
xor U16380 (N_16380,N_9981,N_6828);
nor U16381 (N_16381,N_6808,N_8865);
or U16382 (N_16382,N_9026,N_9466);
nor U16383 (N_16383,N_6448,N_11517);
or U16384 (N_16384,N_9301,N_12379);
nor U16385 (N_16385,N_6894,N_9507);
nor U16386 (N_16386,N_9517,N_6829);
and U16387 (N_16387,N_7536,N_12281);
nand U16388 (N_16388,N_10143,N_9610);
or U16389 (N_16389,N_9728,N_7902);
nand U16390 (N_16390,N_11211,N_9435);
or U16391 (N_16391,N_10159,N_10705);
nand U16392 (N_16392,N_11653,N_11114);
xnor U16393 (N_16393,N_11105,N_10508);
or U16394 (N_16394,N_9568,N_12096);
xor U16395 (N_16395,N_6633,N_10158);
nand U16396 (N_16396,N_9644,N_8226);
and U16397 (N_16397,N_10845,N_6465);
xnor U16398 (N_16398,N_12151,N_11832);
xor U16399 (N_16399,N_9156,N_8781);
and U16400 (N_16400,N_12256,N_9200);
or U16401 (N_16401,N_7939,N_7354);
xor U16402 (N_16402,N_7299,N_7915);
nor U16403 (N_16403,N_6886,N_12062);
xnor U16404 (N_16404,N_11517,N_8831);
xor U16405 (N_16405,N_9530,N_8305);
or U16406 (N_16406,N_10556,N_8743);
xor U16407 (N_16407,N_7638,N_12411);
and U16408 (N_16408,N_11668,N_9539);
and U16409 (N_16409,N_8344,N_9741);
nand U16410 (N_16410,N_9193,N_10176);
nand U16411 (N_16411,N_8694,N_9094);
and U16412 (N_16412,N_8183,N_7291);
xnor U16413 (N_16413,N_12491,N_11538);
xor U16414 (N_16414,N_9742,N_9195);
and U16415 (N_16415,N_10657,N_7181);
nand U16416 (N_16416,N_10718,N_9704);
nor U16417 (N_16417,N_9363,N_11295);
and U16418 (N_16418,N_10389,N_10102);
xor U16419 (N_16419,N_8315,N_6667);
and U16420 (N_16420,N_7608,N_7484);
and U16421 (N_16421,N_6988,N_7533);
or U16422 (N_16422,N_6440,N_9080);
nand U16423 (N_16423,N_7831,N_10014);
and U16424 (N_16424,N_9293,N_11906);
nand U16425 (N_16425,N_11662,N_8422);
nand U16426 (N_16426,N_8406,N_11347);
and U16427 (N_16427,N_6623,N_12459);
or U16428 (N_16428,N_11844,N_7564);
nand U16429 (N_16429,N_8995,N_7522);
xnor U16430 (N_16430,N_6823,N_9369);
xnor U16431 (N_16431,N_8418,N_6468);
nand U16432 (N_16432,N_8181,N_9954);
and U16433 (N_16433,N_10382,N_6941);
nor U16434 (N_16434,N_8571,N_7244);
nand U16435 (N_16435,N_9479,N_12070);
xor U16436 (N_16436,N_6711,N_7072);
and U16437 (N_16437,N_6998,N_9676);
nor U16438 (N_16438,N_11301,N_7817);
xor U16439 (N_16439,N_9281,N_10003);
xor U16440 (N_16440,N_7502,N_9566);
or U16441 (N_16441,N_7985,N_6531);
and U16442 (N_16442,N_8864,N_6861);
or U16443 (N_16443,N_10328,N_12315);
nand U16444 (N_16444,N_11355,N_10696);
nand U16445 (N_16445,N_10574,N_11222);
or U16446 (N_16446,N_11937,N_6834);
nand U16447 (N_16447,N_7602,N_11041);
or U16448 (N_16448,N_11831,N_11066);
nand U16449 (N_16449,N_10769,N_8771);
nand U16450 (N_16450,N_9752,N_6559);
nor U16451 (N_16451,N_12377,N_11548);
xnor U16452 (N_16452,N_9914,N_12389);
xnor U16453 (N_16453,N_10762,N_10915);
or U16454 (N_16454,N_7147,N_12043);
nand U16455 (N_16455,N_9707,N_6779);
nand U16456 (N_16456,N_7936,N_11286);
nor U16457 (N_16457,N_8781,N_6951);
xnor U16458 (N_16458,N_6331,N_11978);
nand U16459 (N_16459,N_12301,N_10461);
nor U16460 (N_16460,N_11267,N_6477);
and U16461 (N_16461,N_8534,N_8757);
nor U16462 (N_16462,N_7481,N_9525);
xor U16463 (N_16463,N_7670,N_12363);
nand U16464 (N_16464,N_9868,N_12320);
or U16465 (N_16465,N_7068,N_10683);
nand U16466 (N_16466,N_6439,N_11548);
xnor U16467 (N_16467,N_10710,N_11847);
or U16468 (N_16468,N_8564,N_10249);
nor U16469 (N_16469,N_9472,N_11041);
xor U16470 (N_16470,N_6792,N_8502);
or U16471 (N_16471,N_9591,N_8241);
or U16472 (N_16472,N_7020,N_12242);
nor U16473 (N_16473,N_10713,N_10208);
and U16474 (N_16474,N_8482,N_11991);
or U16475 (N_16475,N_9743,N_7501);
and U16476 (N_16476,N_12309,N_8978);
nor U16477 (N_16477,N_11027,N_6833);
nand U16478 (N_16478,N_8461,N_6581);
xor U16479 (N_16479,N_9122,N_10321);
or U16480 (N_16480,N_9253,N_7309);
and U16481 (N_16481,N_11191,N_6460);
and U16482 (N_16482,N_11967,N_11877);
nand U16483 (N_16483,N_11968,N_10716);
or U16484 (N_16484,N_6930,N_9419);
xor U16485 (N_16485,N_11081,N_7207);
and U16486 (N_16486,N_9309,N_6271);
nand U16487 (N_16487,N_8797,N_11016);
nor U16488 (N_16488,N_6752,N_9604);
xor U16489 (N_16489,N_10575,N_7153);
xnor U16490 (N_16490,N_10491,N_10951);
or U16491 (N_16491,N_10304,N_9978);
xnor U16492 (N_16492,N_8395,N_7189);
or U16493 (N_16493,N_11614,N_7211);
nor U16494 (N_16494,N_10947,N_11132);
and U16495 (N_16495,N_12449,N_10934);
and U16496 (N_16496,N_8356,N_9677);
and U16497 (N_16497,N_8121,N_8742);
and U16498 (N_16498,N_7211,N_7569);
nor U16499 (N_16499,N_6612,N_11392);
nor U16500 (N_16500,N_10152,N_6695);
xnor U16501 (N_16501,N_9244,N_8331);
nor U16502 (N_16502,N_8233,N_10671);
nor U16503 (N_16503,N_7294,N_9555);
xor U16504 (N_16504,N_10457,N_6880);
and U16505 (N_16505,N_7310,N_11298);
nand U16506 (N_16506,N_11405,N_8321);
and U16507 (N_16507,N_12228,N_12085);
and U16508 (N_16508,N_10113,N_8915);
or U16509 (N_16509,N_6428,N_9462);
nor U16510 (N_16510,N_9619,N_10799);
or U16511 (N_16511,N_12473,N_9623);
nand U16512 (N_16512,N_12466,N_10735);
nor U16513 (N_16513,N_7638,N_9996);
nor U16514 (N_16514,N_10176,N_12043);
nor U16515 (N_16515,N_9552,N_10367);
xnor U16516 (N_16516,N_7772,N_11426);
or U16517 (N_16517,N_9380,N_8203);
nor U16518 (N_16518,N_6770,N_11849);
or U16519 (N_16519,N_9766,N_11650);
nor U16520 (N_16520,N_6297,N_10932);
xor U16521 (N_16521,N_11143,N_10389);
nand U16522 (N_16522,N_7455,N_11989);
xnor U16523 (N_16523,N_6333,N_7453);
xnor U16524 (N_16524,N_11745,N_6587);
nand U16525 (N_16525,N_10999,N_11055);
nand U16526 (N_16526,N_8054,N_11503);
and U16527 (N_16527,N_8316,N_11247);
nand U16528 (N_16528,N_9502,N_10662);
xnor U16529 (N_16529,N_9056,N_8147);
nor U16530 (N_16530,N_9728,N_7228);
or U16531 (N_16531,N_7154,N_8004);
or U16532 (N_16532,N_10113,N_7060);
or U16533 (N_16533,N_11799,N_11563);
nand U16534 (N_16534,N_11003,N_12173);
nor U16535 (N_16535,N_7407,N_8205);
or U16536 (N_16536,N_6895,N_11504);
or U16537 (N_16537,N_11267,N_12443);
nand U16538 (N_16538,N_7043,N_8800);
or U16539 (N_16539,N_8894,N_10159);
or U16540 (N_16540,N_8509,N_7480);
nor U16541 (N_16541,N_9927,N_8719);
nor U16542 (N_16542,N_7895,N_7816);
or U16543 (N_16543,N_8203,N_6780);
or U16544 (N_16544,N_8978,N_7393);
and U16545 (N_16545,N_10670,N_7617);
xor U16546 (N_16546,N_7345,N_10231);
nor U16547 (N_16547,N_7292,N_9667);
xnor U16548 (N_16548,N_11685,N_7783);
nand U16549 (N_16549,N_8351,N_6748);
xor U16550 (N_16550,N_9638,N_9511);
and U16551 (N_16551,N_11719,N_12289);
xor U16552 (N_16552,N_6892,N_6642);
nand U16553 (N_16553,N_10823,N_12304);
nor U16554 (N_16554,N_7025,N_7933);
nand U16555 (N_16555,N_7689,N_7980);
nand U16556 (N_16556,N_7057,N_7291);
or U16557 (N_16557,N_6856,N_7914);
nor U16558 (N_16558,N_10236,N_7922);
or U16559 (N_16559,N_10629,N_11107);
or U16560 (N_16560,N_10819,N_10541);
xor U16561 (N_16561,N_8083,N_11216);
or U16562 (N_16562,N_8219,N_8493);
and U16563 (N_16563,N_10361,N_7026);
or U16564 (N_16564,N_8129,N_10424);
xor U16565 (N_16565,N_8021,N_6777);
or U16566 (N_16566,N_6830,N_7693);
or U16567 (N_16567,N_6957,N_10114);
xor U16568 (N_16568,N_9759,N_8531);
nor U16569 (N_16569,N_7966,N_8297);
xnor U16570 (N_16570,N_7328,N_10762);
and U16571 (N_16571,N_8855,N_7064);
nand U16572 (N_16572,N_6796,N_8271);
or U16573 (N_16573,N_7742,N_9743);
xor U16574 (N_16574,N_11306,N_8617);
nand U16575 (N_16575,N_6763,N_6594);
nand U16576 (N_16576,N_7794,N_9974);
and U16577 (N_16577,N_6437,N_11795);
and U16578 (N_16578,N_11441,N_7969);
and U16579 (N_16579,N_8834,N_8233);
nand U16580 (N_16580,N_7352,N_11415);
nor U16581 (N_16581,N_6528,N_9050);
and U16582 (N_16582,N_12082,N_11763);
xnor U16583 (N_16583,N_10958,N_10149);
xnor U16584 (N_16584,N_6310,N_6768);
or U16585 (N_16585,N_11656,N_7111);
or U16586 (N_16586,N_8999,N_9797);
or U16587 (N_16587,N_9458,N_8602);
nor U16588 (N_16588,N_6950,N_9388);
nor U16589 (N_16589,N_8089,N_6656);
or U16590 (N_16590,N_11951,N_12333);
xor U16591 (N_16591,N_9123,N_11573);
nand U16592 (N_16592,N_7719,N_9874);
xor U16593 (N_16593,N_6843,N_11880);
nor U16594 (N_16594,N_9961,N_6339);
nor U16595 (N_16595,N_11992,N_10817);
or U16596 (N_16596,N_11796,N_10331);
nand U16597 (N_16597,N_11167,N_8034);
xnor U16598 (N_16598,N_12365,N_11444);
or U16599 (N_16599,N_8200,N_6644);
xnor U16600 (N_16600,N_11586,N_10150);
and U16601 (N_16601,N_10172,N_10562);
or U16602 (N_16602,N_11031,N_11065);
nor U16603 (N_16603,N_9733,N_12355);
and U16604 (N_16604,N_9464,N_10771);
and U16605 (N_16605,N_8742,N_9705);
nor U16606 (N_16606,N_6762,N_10000);
nand U16607 (N_16607,N_7202,N_8479);
nor U16608 (N_16608,N_6439,N_8174);
xor U16609 (N_16609,N_6851,N_6871);
or U16610 (N_16610,N_8936,N_11048);
and U16611 (N_16611,N_10279,N_9755);
nand U16612 (N_16612,N_10198,N_10532);
nand U16613 (N_16613,N_6518,N_11766);
nor U16614 (N_16614,N_10144,N_7478);
nand U16615 (N_16615,N_10681,N_7277);
and U16616 (N_16616,N_6562,N_10628);
nand U16617 (N_16617,N_9553,N_7992);
and U16618 (N_16618,N_9940,N_10531);
and U16619 (N_16619,N_6837,N_8611);
xor U16620 (N_16620,N_7901,N_12210);
or U16621 (N_16621,N_6889,N_9606);
or U16622 (N_16622,N_10524,N_10157);
or U16623 (N_16623,N_12445,N_8391);
nand U16624 (N_16624,N_8829,N_8037);
or U16625 (N_16625,N_8512,N_10271);
nor U16626 (N_16626,N_8347,N_8765);
or U16627 (N_16627,N_9232,N_8642);
or U16628 (N_16628,N_8040,N_9043);
or U16629 (N_16629,N_10206,N_12391);
xor U16630 (N_16630,N_6934,N_11732);
nor U16631 (N_16631,N_9327,N_8109);
xor U16632 (N_16632,N_11269,N_7779);
or U16633 (N_16633,N_11507,N_10144);
or U16634 (N_16634,N_12048,N_6962);
xor U16635 (N_16635,N_9808,N_8251);
nand U16636 (N_16636,N_7535,N_10038);
and U16637 (N_16637,N_6670,N_8714);
or U16638 (N_16638,N_6790,N_6287);
or U16639 (N_16639,N_12425,N_11301);
or U16640 (N_16640,N_7847,N_12279);
xnor U16641 (N_16641,N_6407,N_8052);
nor U16642 (N_16642,N_6761,N_11262);
and U16643 (N_16643,N_9341,N_11329);
nand U16644 (N_16644,N_8510,N_9175);
or U16645 (N_16645,N_10475,N_6362);
and U16646 (N_16646,N_11392,N_12130);
xor U16647 (N_16647,N_6315,N_10382);
nor U16648 (N_16648,N_11647,N_9739);
and U16649 (N_16649,N_9928,N_9171);
xnor U16650 (N_16650,N_6841,N_9292);
or U16651 (N_16651,N_11275,N_9696);
xor U16652 (N_16652,N_10239,N_7182);
nor U16653 (N_16653,N_8992,N_11606);
and U16654 (N_16654,N_11055,N_7621);
or U16655 (N_16655,N_9787,N_9954);
nor U16656 (N_16656,N_10583,N_8391);
and U16657 (N_16657,N_8046,N_10311);
xor U16658 (N_16658,N_12067,N_9237);
and U16659 (N_16659,N_7221,N_10098);
nor U16660 (N_16660,N_8650,N_7045);
or U16661 (N_16661,N_8173,N_6423);
or U16662 (N_16662,N_12247,N_7859);
or U16663 (N_16663,N_7413,N_10410);
nor U16664 (N_16664,N_6828,N_8568);
nor U16665 (N_16665,N_10975,N_12372);
nand U16666 (N_16666,N_8679,N_10010);
and U16667 (N_16667,N_9788,N_7107);
and U16668 (N_16668,N_11275,N_6599);
xor U16669 (N_16669,N_8477,N_10019);
xor U16670 (N_16670,N_10756,N_11046);
nand U16671 (N_16671,N_6770,N_9663);
nand U16672 (N_16672,N_8506,N_8273);
and U16673 (N_16673,N_11040,N_6779);
and U16674 (N_16674,N_10651,N_11620);
or U16675 (N_16675,N_8926,N_8471);
or U16676 (N_16676,N_9168,N_9943);
nor U16677 (N_16677,N_9914,N_11566);
or U16678 (N_16678,N_8359,N_12197);
and U16679 (N_16679,N_7266,N_6490);
xnor U16680 (N_16680,N_8767,N_10393);
nor U16681 (N_16681,N_7637,N_6417);
xor U16682 (N_16682,N_9253,N_10907);
nand U16683 (N_16683,N_11614,N_7475);
nor U16684 (N_16684,N_9458,N_6554);
xor U16685 (N_16685,N_8380,N_6555);
nor U16686 (N_16686,N_8579,N_9108);
xor U16687 (N_16687,N_10882,N_6701);
xor U16688 (N_16688,N_6838,N_8234);
and U16689 (N_16689,N_7802,N_9076);
and U16690 (N_16690,N_10845,N_10100);
nor U16691 (N_16691,N_6948,N_11645);
nor U16692 (N_16692,N_11756,N_7766);
nand U16693 (N_16693,N_11860,N_10821);
xnor U16694 (N_16694,N_6380,N_9032);
and U16695 (N_16695,N_9835,N_6499);
nand U16696 (N_16696,N_7342,N_11424);
nand U16697 (N_16697,N_9507,N_10056);
xor U16698 (N_16698,N_11218,N_11545);
nand U16699 (N_16699,N_10351,N_10553);
or U16700 (N_16700,N_11461,N_7326);
nor U16701 (N_16701,N_10041,N_6341);
xnor U16702 (N_16702,N_6489,N_12455);
nand U16703 (N_16703,N_9917,N_6429);
nor U16704 (N_16704,N_10888,N_8536);
and U16705 (N_16705,N_8419,N_7390);
and U16706 (N_16706,N_7689,N_10766);
xnor U16707 (N_16707,N_11359,N_7850);
nor U16708 (N_16708,N_8746,N_10056);
or U16709 (N_16709,N_11808,N_10280);
or U16710 (N_16710,N_11991,N_10916);
nand U16711 (N_16711,N_9625,N_9536);
nand U16712 (N_16712,N_7782,N_12484);
nor U16713 (N_16713,N_7639,N_12287);
and U16714 (N_16714,N_8264,N_8592);
nor U16715 (N_16715,N_8251,N_11742);
nand U16716 (N_16716,N_9475,N_8836);
nor U16717 (N_16717,N_8425,N_8604);
and U16718 (N_16718,N_11656,N_11223);
or U16719 (N_16719,N_8190,N_7340);
nand U16720 (N_16720,N_10579,N_9965);
xnor U16721 (N_16721,N_7620,N_9132);
nand U16722 (N_16722,N_8972,N_6838);
nand U16723 (N_16723,N_11047,N_9808);
and U16724 (N_16724,N_11666,N_10135);
and U16725 (N_16725,N_11223,N_10856);
nor U16726 (N_16726,N_11543,N_7095);
or U16727 (N_16727,N_8646,N_11017);
nand U16728 (N_16728,N_8924,N_10782);
nor U16729 (N_16729,N_6751,N_7689);
or U16730 (N_16730,N_11390,N_9699);
nor U16731 (N_16731,N_12260,N_9429);
and U16732 (N_16732,N_8375,N_8337);
or U16733 (N_16733,N_10212,N_10200);
or U16734 (N_16734,N_6276,N_9884);
or U16735 (N_16735,N_8089,N_11520);
nor U16736 (N_16736,N_6574,N_7140);
xor U16737 (N_16737,N_6792,N_7115);
or U16738 (N_16738,N_11817,N_8975);
nand U16739 (N_16739,N_6841,N_8576);
nand U16740 (N_16740,N_11754,N_11032);
and U16741 (N_16741,N_7864,N_11069);
nor U16742 (N_16742,N_9433,N_7989);
nand U16743 (N_16743,N_6814,N_11970);
nor U16744 (N_16744,N_9729,N_11441);
nor U16745 (N_16745,N_6728,N_11002);
nor U16746 (N_16746,N_6827,N_7406);
and U16747 (N_16747,N_10321,N_9069);
nor U16748 (N_16748,N_6310,N_10515);
nand U16749 (N_16749,N_6753,N_7554);
xor U16750 (N_16750,N_11298,N_11881);
nor U16751 (N_16751,N_7664,N_9011);
xor U16752 (N_16752,N_10045,N_9266);
or U16753 (N_16753,N_11449,N_9712);
xnor U16754 (N_16754,N_7533,N_9421);
nand U16755 (N_16755,N_11410,N_7439);
xor U16756 (N_16756,N_10779,N_7235);
nor U16757 (N_16757,N_6403,N_7991);
xnor U16758 (N_16758,N_10573,N_12100);
nor U16759 (N_16759,N_11449,N_11536);
nor U16760 (N_16760,N_8820,N_12370);
and U16761 (N_16761,N_9307,N_7356);
xnor U16762 (N_16762,N_7066,N_12473);
and U16763 (N_16763,N_9675,N_7708);
and U16764 (N_16764,N_10366,N_6362);
nand U16765 (N_16765,N_9449,N_10907);
nor U16766 (N_16766,N_8194,N_8090);
and U16767 (N_16767,N_7964,N_6742);
or U16768 (N_16768,N_6601,N_7972);
nand U16769 (N_16769,N_8691,N_11241);
xnor U16770 (N_16770,N_11368,N_9907);
xnor U16771 (N_16771,N_7411,N_11664);
nor U16772 (N_16772,N_11348,N_11053);
or U16773 (N_16773,N_11845,N_10945);
or U16774 (N_16774,N_11840,N_11711);
or U16775 (N_16775,N_9531,N_7884);
nand U16776 (N_16776,N_9710,N_8510);
nor U16777 (N_16777,N_12204,N_8856);
nor U16778 (N_16778,N_11614,N_10464);
xor U16779 (N_16779,N_9205,N_7686);
xnor U16780 (N_16780,N_9928,N_8977);
xor U16781 (N_16781,N_11997,N_11675);
nor U16782 (N_16782,N_9140,N_6606);
xnor U16783 (N_16783,N_12369,N_7895);
nor U16784 (N_16784,N_10311,N_6471);
nor U16785 (N_16785,N_6780,N_10294);
nor U16786 (N_16786,N_9248,N_12191);
xnor U16787 (N_16787,N_11955,N_9625);
nand U16788 (N_16788,N_11271,N_10370);
and U16789 (N_16789,N_10195,N_11033);
and U16790 (N_16790,N_9532,N_11275);
nor U16791 (N_16791,N_7277,N_11539);
nand U16792 (N_16792,N_8627,N_8311);
or U16793 (N_16793,N_10556,N_11859);
nor U16794 (N_16794,N_9226,N_10305);
and U16795 (N_16795,N_9937,N_10052);
and U16796 (N_16796,N_10934,N_9488);
nand U16797 (N_16797,N_10127,N_6295);
or U16798 (N_16798,N_10000,N_10741);
nand U16799 (N_16799,N_6313,N_6405);
xnor U16800 (N_16800,N_10643,N_9897);
nand U16801 (N_16801,N_6777,N_10631);
or U16802 (N_16802,N_7412,N_10738);
nand U16803 (N_16803,N_11566,N_8338);
or U16804 (N_16804,N_11907,N_10051);
xor U16805 (N_16805,N_10913,N_8449);
and U16806 (N_16806,N_11024,N_8787);
nand U16807 (N_16807,N_10049,N_12190);
and U16808 (N_16808,N_7964,N_8642);
and U16809 (N_16809,N_7783,N_11773);
nand U16810 (N_16810,N_8928,N_11369);
or U16811 (N_16811,N_10359,N_11837);
xor U16812 (N_16812,N_9850,N_9190);
and U16813 (N_16813,N_7141,N_12329);
nand U16814 (N_16814,N_7524,N_11072);
nor U16815 (N_16815,N_9990,N_8573);
or U16816 (N_16816,N_11079,N_10421);
xor U16817 (N_16817,N_11819,N_9378);
and U16818 (N_16818,N_8204,N_12214);
xnor U16819 (N_16819,N_12305,N_9158);
nor U16820 (N_16820,N_9104,N_8873);
or U16821 (N_16821,N_11040,N_8750);
and U16822 (N_16822,N_10900,N_8136);
and U16823 (N_16823,N_9259,N_7754);
and U16824 (N_16824,N_10939,N_11103);
xor U16825 (N_16825,N_7324,N_7377);
nor U16826 (N_16826,N_11462,N_10600);
xnor U16827 (N_16827,N_10149,N_12455);
and U16828 (N_16828,N_6354,N_9953);
or U16829 (N_16829,N_8548,N_12380);
xor U16830 (N_16830,N_7225,N_6317);
or U16831 (N_16831,N_7398,N_9994);
or U16832 (N_16832,N_7088,N_7187);
nor U16833 (N_16833,N_6360,N_7360);
nand U16834 (N_16834,N_10896,N_11302);
nor U16835 (N_16835,N_9490,N_9027);
xor U16836 (N_16836,N_7643,N_9741);
or U16837 (N_16837,N_7288,N_11767);
or U16838 (N_16838,N_10098,N_10909);
and U16839 (N_16839,N_12364,N_8974);
nand U16840 (N_16840,N_12344,N_8348);
nor U16841 (N_16841,N_6793,N_11407);
nand U16842 (N_16842,N_11919,N_9361);
nand U16843 (N_16843,N_11369,N_7499);
nor U16844 (N_16844,N_12382,N_11117);
and U16845 (N_16845,N_8869,N_12071);
nand U16846 (N_16846,N_6943,N_9649);
or U16847 (N_16847,N_7612,N_10698);
or U16848 (N_16848,N_8121,N_11262);
nor U16849 (N_16849,N_11124,N_9669);
or U16850 (N_16850,N_10915,N_6723);
nand U16851 (N_16851,N_11220,N_10202);
nor U16852 (N_16852,N_8406,N_8395);
xor U16853 (N_16853,N_6809,N_8663);
or U16854 (N_16854,N_11842,N_9995);
xnor U16855 (N_16855,N_7151,N_11489);
nand U16856 (N_16856,N_6348,N_10005);
nor U16857 (N_16857,N_9947,N_9497);
or U16858 (N_16858,N_7448,N_11890);
nor U16859 (N_16859,N_11993,N_7805);
xnor U16860 (N_16860,N_7486,N_11377);
or U16861 (N_16861,N_10084,N_10757);
nor U16862 (N_16862,N_11666,N_12140);
or U16863 (N_16863,N_12104,N_11513);
nor U16864 (N_16864,N_11328,N_8766);
xor U16865 (N_16865,N_10181,N_9452);
and U16866 (N_16866,N_12312,N_10451);
nor U16867 (N_16867,N_10915,N_10384);
and U16868 (N_16868,N_8214,N_10108);
and U16869 (N_16869,N_8721,N_11909);
xor U16870 (N_16870,N_12351,N_8001);
nand U16871 (N_16871,N_10225,N_6826);
nor U16872 (N_16872,N_9639,N_6411);
or U16873 (N_16873,N_11470,N_11812);
nand U16874 (N_16874,N_10359,N_11920);
and U16875 (N_16875,N_7316,N_10123);
or U16876 (N_16876,N_6818,N_7559);
xor U16877 (N_16877,N_7002,N_6599);
or U16878 (N_16878,N_10356,N_10546);
nand U16879 (N_16879,N_7306,N_9757);
and U16880 (N_16880,N_8468,N_6607);
nand U16881 (N_16881,N_6582,N_9497);
and U16882 (N_16882,N_11728,N_6900);
and U16883 (N_16883,N_11985,N_9341);
xor U16884 (N_16884,N_10738,N_10831);
or U16885 (N_16885,N_9462,N_6892);
and U16886 (N_16886,N_8429,N_8366);
nand U16887 (N_16887,N_10700,N_12312);
or U16888 (N_16888,N_7123,N_11384);
or U16889 (N_16889,N_10189,N_8669);
xor U16890 (N_16890,N_10226,N_8945);
nor U16891 (N_16891,N_11996,N_10653);
and U16892 (N_16892,N_6403,N_11401);
nand U16893 (N_16893,N_11160,N_10911);
nand U16894 (N_16894,N_10455,N_9280);
or U16895 (N_16895,N_6959,N_9405);
nor U16896 (N_16896,N_10918,N_6924);
and U16897 (N_16897,N_11139,N_11864);
xor U16898 (N_16898,N_7218,N_6574);
and U16899 (N_16899,N_7809,N_12322);
nor U16900 (N_16900,N_7115,N_9798);
xor U16901 (N_16901,N_6307,N_10681);
xnor U16902 (N_16902,N_8147,N_6370);
nand U16903 (N_16903,N_12017,N_8958);
xnor U16904 (N_16904,N_7990,N_10227);
or U16905 (N_16905,N_7993,N_10121);
xor U16906 (N_16906,N_8924,N_10680);
xnor U16907 (N_16907,N_6337,N_8809);
nor U16908 (N_16908,N_8713,N_8915);
nor U16909 (N_16909,N_10554,N_9071);
or U16910 (N_16910,N_9306,N_7812);
and U16911 (N_16911,N_9669,N_6385);
nor U16912 (N_16912,N_8859,N_10930);
nor U16913 (N_16913,N_10759,N_6500);
nor U16914 (N_16914,N_11115,N_9269);
nor U16915 (N_16915,N_8231,N_9449);
or U16916 (N_16916,N_12132,N_10259);
xor U16917 (N_16917,N_12441,N_10422);
or U16918 (N_16918,N_11529,N_11162);
xnor U16919 (N_16919,N_11044,N_9764);
nor U16920 (N_16920,N_10479,N_10686);
nand U16921 (N_16921,N_6285,N_11315);
xor U16922 (N_16922,N_9495,N_8858);
nor U16923 (N_16923,N_12311,N_11650);
or U16924 (N_16924,N_7436,N_8318);
nand U16925 (N_16925,N_8786,N_10083);
and U16926 (N_16926,N_10191,N_6530);
nor U16927 (N_16927,N_10097,N_11547);
nor U16928 (N_16928,N_7746,N_9307);
or U16929 (N_16929,N_10147,N_7067);
xor U16930 (N_16930,N_12412,N_8148);
or U16931 (N_16931,N_7571,N_7442);
or U16932 (N_16932,N_10973,N_7007);
or U16933 (N_16933,N_6547,N_9690);
nand U16934 (N_16934,N_11516,N_11758);
nor U16935 (N_16935,N_9019,N_11343);
xnor U16936 (N_16936,N_10259,N_8110);
and U16937 (N_16937,N_8073,N_7010);
or U16938 (N_16938,N_11369,N_10528);
nand U16939 (N_16939,N_7049,N_7038);
nor U16940 (N_16940,N_7823,N_6986);
xor U16941 (N_16941,N_11415,N_12290);
and U16942 (N_16942,N_10833,N_11531);
nand U16943 (N_16943,N_11254,N_10692);
and U16944 (N_16944,N_7389,N_7928);
nor U16945 (N_16945,N_11292,N_12214);
nor U16946 (N_16946,N_12083,N_11011);
and U16947 (N_16947,N_10848,N_9999);
xor U16948 (N_16948,N_9607,N_7365);
xor U16949 (N_16949,N_10226,N_9894);
nand U16950 (N_16950,N_10141,N_8302);
xnor U16951 (N_16951,N_7522,N_9460);
nor U16952 (N_16952,N_11646,N_11831);
or U16953 (N_16953,N_6830,N_11742);
nor U16954 (N_16954,N_11854,N_9188);
nand U16955 (N_16955,N_10776,N_6729);
nor U16956 (N_16956,N_9843,N_7033);
xnor U16957 (N_16957,N_9774,N_7359);
and U16958 (N_16958,N_9438,N_6783);
and U16959 (N_16959,N_10289,N_9262);
and U16960 (N_16960,N_7439,N_12240);
xnor U16961 (N_16961,N_10472,N_12120);
or U16962 (N_16962,N_12430,N_10172);
nand U16963 (N_16963,N_7917,N_8995);
nor U16964 (N_16964,N_6521,N_7082);
or U16965 (N_16965,N_11346,N_11349);
and U16966 (N_16966,N_6392,N_10353);
nor U16967 (N_16967,N_10132,N_6916);
or U16968 (N_16968,N_6519,N_6984);
or U16969 (N_16969,N_8356,N_11240);
xor U16970 (N_16970,N_7924,N_6523);
nor U16971 (N_16971,N_9578,N_11435);
nor U16972 (N_16972,N_10714,N_8464);
and U16973 (N_16973,N_9568,N_6312);
nor U16974 (N_16974,N_6596,N_7422);
and U16975 (N_16975,N_6290,N_8356);
xnor U16976 (N_16976,N_11715,N_9598);
nand U16977 (N_16977,N_9432,N_11569);
nor U16978 (N_16978,N_11579,N_9327);
or U16979 (N_16979,N_9899,N_10523);
nor U16980 (N_16980,N_11165,N_12165);
and U16981 (N_16981,N_11281,N_10879);
nand U16982 (N_16982,N_8736,N_8576);
xor U16983 (N_16983,N_8698,N_10083);
nor U16984 (N_16984,N_10361,N_12473);
or U16985 (N_16985,N_8240,N_7540);
and U16986 (N_16986,N_6570,N_10748);
xor U16987 (N_16987,N_8444,N_7245);
nor U16988 (N_16988,N_9280,N_9562);
and U16989 (N_16989,N_10083,N_9636);
xor U16990 (N_16990,N_9144,N_9773);
or U16991 (N_16991,N_10765,N_10047);
nor U16992 (N_16992,N_6277,N_11387);
and U16993 (N_16993,N_11707,N_10590);
xnor U16994 (N_16994,N_12207,N_12160);
or U16995 (N_16995,N_11333,N_9873);
xor U16996 (N_16996,N_10474,N_12303);
and U16997 (N_16997,N_11958,N_10083);
or U16998 (N_16998,N_9701,N_8664);
and U16999 (N_16999,N_10029,N_10770);
nand U17000 (N_17000,N_10453,N_8247);
nand U17001 (N_17001,N_8072,N_11160);
nand U17002 (N_17002,N_7002,N_7479);
and U17003 (N_17003,N_12135,N_7019);
xnor U17004 (N_17004,N_7899,N_9749);
xnor U17005 (N_17005,N_6859,N_7765);
and U17006 (N_17006,N_10743,N_11997);
nor U17007 (N_17007,N_7439,N_8362);
or U17008 (N_17008,N_10404,N_6284);
or U17009 (N_17009,N_9713,N_9618);
and U17010 (N_17010,N_8460,N_7169);
and U17011 (N_17011,N_11081,N_11532);
nor U17012 (N_17012,N_10160,N_8761);
and U17013 (N_17013,N_7635,N_7294);
xor U17014 (N_17014,N_6465,N_8300);
nor U17015 (N_17015,N_7235,N_11498);
and U17016 (N_17016,N_8552,N_7027);
or U17017 (N_17017,N_7984,N_8618);
and U17018 (N_17018,N_10632,N_8025);
xor U17019 (N_17019,N_7859,N_8306);
nor U17020 (N_17020,N_10646,N_6790);
and U17021 (N_17021,N_7693,N_7878);
and U17022 (N_17022,N_7195,N_9287);
or U17023 (N_17023,N_11799,N_10680);
and U17024 (N_17024,N_10069,N_9737);
nand U17025 (N_17025,N_10542,N_9905);
nand U17026 (N_17026,N_9512,N_9963);
xnor U17027 (N_17027,N_11838,N_9537);
nor U17028 (N_17028,N_11874,N_9624);
xor U17029 (N_17029,N_12257,N_9802);
nand U17030 (N_17030,N_7851,N_10411);
nor U17031 (N_17031,N_7605,N_7346);
nor U17032 (N_17032,N_7753,N_6728);
and U17033 (N_17033,N_8788,N_12121);
nand U17034 (N_17034,N_12098,N_10424);
nand U17035 (N_17035,N_11574,N_11422);
xor U17036 (N_17036,N_10623,N_9357);
nor U17037 (N_17037,N_9433,N_10126);
xor U17038 (N_17038,N_6278,N_7211);
or U17039 (N_17039,N_6758,N_6819);
and U17040 (N_17040,N_10878,N_9149);
xor U17041 (N_17041,N_10559,N_8160);
and U17042 (N_17042,N_10927,N_8888);
nand U17043 (N_17043,N_6688,N_11452);
nor U17044 (N_17044,N_9083,N_8141);
nor U17045 (N_17045,N_6281,N_11606);
xor U17046 (N_17046,N_7054,N_9009);
xnor U17047 (N_17047,N_11346,N_11169);
nand U17048 (N_17048,N_8442,N_11102);
xor U17049 (N_17049,N_11306,N_8122);
nand U17050 (N_17050,N_11275,N_7960);
and U17051 (N_17051,N_10470,N_7387);
nor U17052 (N_17052,N_11084,N_10376);
and U17053 (N_17053,N_11706,N_10996);
nor U17054 (N_17054,N_8693,N_10864);
nand U17055 (N_17055,N_11397,N_7104);
nand U17056 (N_17056,N_8203,N_7968);
nor U17057 (N_17057,N_9610,N_9208);
nor U17058 (N_17058,N_9168,N_11629);
xor U17059 (N_17059,N_10507,N_8261);
or U17060 (N_17060,N_8604,N_7378);
nor U17061 (N_17061,N_7207,N_9366);
nand U17062 (N_17062,N_10166,N_10414);
xor U17063 (N_17063,N_11736,N_10456);
nor U17064 (N_17064,N_12179,N_10687);
nand U17065 (N_17065,N_11898,N_9177);
nand U17066 (N_17066,N_9896,N_12496);
or U17067 (N_17067,N_10947,N_11402);
or U17068 (N_17068,N_8228,N_10032);
xnor U17069 (N_17069,N_8113,N_11827);
xor U17070 (N_17070,N_12432,N_11107);
nor U17071 (N_17071,N_8061,N_11756);
or U17072 (N_17072,N_10030,N_6889);
nor U17073 (N_17073,N_6723,N_10066);
and U17074 (N_17074,N_11522,N_7862);
nand U17075 (N_17075,N_11687,N_9599);
nand U17076 (N_17076,N_8221,N_10971);
or U17077 (N_17077,N_9088,N_7725);
and U17078 (N_17078,N_6660,N_6665);
and U17079 (N_17079,N_11084,N_9574);
nand U17080 (N_17080,N_11271,N_11436);
nor U17081 (N_17081,N_11806,N_6652);
xnor U17082 (N_17082,N_9725,N_11301);
nor U17083 (N_17083,N_11422,N_9641);
and U17084 (N_17084,N_9846,N_9529);
nor U17085 (N_17085,N_12023,N_10820);
xor U17086 (N_17086,N_11989,N_8506);
and U17087 (N_17087,N_12097,N_7450);
or U17088 (N_17088,N_6308,N_11806);
nand U17089 (N_17089,N_10107,N_7111);
nor U17090 (N_17090,N_6803,N_6334);
nand U17091 (N_17091,N_11841,N_10812);
nor U17092 (N_17092,N_11231,N_10937);
and U17093 (N_17093,N_6260,N_12402);
or U17094 (N_17094,N_10184,N_10219);
and U17095 (N_17095,N_12102,N_9897);
xor U17096 (N_17096,N_7180,N_8476);
nor U17097 (N_17097,N_11051,N_11660);
xor U17098 (N_17098,N_10230,N_8706);
nor U17099 (N_17099,N_6546,N_8490);
nor U17100 (N_17100,N_8878,N_8227);
and U17101 (N_17101,N_11268,N_11848);
and U17102 (N_17102,N_11437,N_7871);
nor U17103 (N_17103,N_8076,N_6741);
nand U17104 (N_17104,N_10377,N_12024);
and U17105 (N_17105,N_9988,N_11807);
nor U17106 (N_17106,N_8023,N_8863);
nor U17107 (N_17107,N_6499,N_6432);
or U17108 (N_17108,N_10046,N_7727);
nand U17109 (N_17109,N_7585,N_8752);
nand U17110 (N_17110,N_10381,N_8005);
xor U17111 (N_17111,N_6825,N_11870);
or U17112 (N_17112,N_10451,N_6438);
nor U17113 (N_17113,N_9415,N_8839);
xnor U17114 (N_17114,N_12126,N_10871);
or U17115 (N_17115,N_9506,N_6643);
or U17116 (N_17116,N_12464,N_11134);
or U17117 (N_17117,N_9569,N_12432);
or U17118 (N_17118,N_8588,N_7596);
or U17119 (N_17119,N_10183,N_10319);
xor U17120 (N_17120,N_7692,N_7375);
nand U17121 (N_17121,N_7023,N_10301);
nand U17122 (N_17122,N_8428,N_9810);
nand U17123 (N_17123,N_10640,N_10809);
or U17124 (N_17124,N_11053,N_8333);
or U17125 (N_17125,N_7552,N_6734);
or U17126 (N_17126,N_9855,N_8541);
nand U17127 (N_17127,N_9172,N_6271);
or U17128 (N_17128,N_8532,N_11815);
nor U17129 (N_17129,N_7830,N_10188);
nand U17130 (N_17130,N_11784,N_7246);
nand U17131 (N_17131,N_6511,N_9824);
xnor U17132 (N_17132,N_12112,N_9491);
or U17133 (N_17133,N_10139,N_9639);
nor U17134 (N_17134,N_7627,N_10078);
and U17135 (N_17135,N_10906,N_9813);
xnor U17136 (N_17136,N_8690,N_9989);
and U17137 (N_17137,N_11672,N_7276);
nand U17138 (N_17138,N_8772,N_6328);
or U17139 (N_17139,N_10384,N_6576);
and U17140 (N_17140,N_11248,N_8889);
nor U17141 (N_17141,N_6361,N_11418);
xnor U17142 (N_17142,N_11975,N_6541);
nand U17143 (N_17143,N_7656,N_10331);
nor U17144 (N_17144,N_10882,N_6557);
and U17145 (N_17145,N_6304,N_6613);
and U17146 (N_17146,N_11906,N_12485);
and U17147 (N_17147,N_7321,N_8578);
xnor U17148 (N_17148,N_7242,N_11715);
xnor U17149 (N_17149,N_8749,N_9633);
nand U17150 (N_17150,N_9178,N_12083);
nor U17151 (N_17151,N_7966,N_10278);
nor U17152 (N_17152,N_7863,N_7441);
nand U17153 (N_17153,N_7310,N_11591);
nor U17154 (N_17154,N_9985,N_11762);
and U17155 (N_17155,N_8434,N_9971);
nand U17156 (N_17156,N_12226,N_7194);
or U17157 (N_17157,N_12241,N_6307);
xnor U17158 (N_17158,N_7047,N_6571);
and U17159 (N_17159,N_7400,N_12327);
xnor U17160 (N_17160,N_7637,N_10690);
nand U17161 (N_17161,N_9382,N_11521);
and U17162 (N_17162,N_7200,N_11380);
or U17163 (N_17163,N_6346,N_8946);
xnor U17164 (N_17164,N_7316,N_9605);
and U17165 (N_17165,N_11545,N_11028);
nand U17166 (N_17166,N_8160,N_11139);
or U17167 (N_17167,N_9660,N_10385);
nand U17168 (N_17168,N_8842,N_11948);
nand U17169 (N_17169,N_9673,N_8239);
and U17170 (N_17170,N_12304,N_9339);
nand U17171 (N_17171,N_11611,N_7488);
nor U17172 (N_17172,N_11544,N_8641);
nand U17173 (N_17173,N_8595,N_12485);
xnor U17174 (N_17174,N_9563,N_10257);
xor U17175 (N_17175,N_9649,N_8480);
nor U17176 (N_17176,N_6643,N_8059);
or U17177 (N_17177,N_11027,N_10661);
xor U17178 (N_17178,N_11578,N_11677);
or U17179 (N_17179,N_11237,N_6898);
or U17180 (N_17180,N_10981,N_8278);
and U17181 (N_17181,N_9832,N_10428);
xor U17182 (N_17182,N_10764,N_7623);
nor U17183 (N_17183,N_8084,N_8886);
nor U17184 (N_17184,N_11938,N_11329);
nor U17185 (N_17185,N_6953,N_6607);
nor U17186 (N_17186,N_8709,N_9570);
nand U17187 (N_17187,N_7339,N_11588);
and U17188 (N_17188,N_9195,N_9682);
and U17189 (N_17189,N_11737,N_8747);
nor U17190 (N_17190,N_8793,N_7963);
or U17191 (N_17191,N_8176,N_6395);
nand U17192 (N_17192,N_8747,N_7529);
xnor U17193 (N_17193,N_7629,N_10240);
or U17194 (N_17194,N_9279,N_6272);
or U17195 (N_17195,N_9457,N_9538);
xnor U17196 (N_17196,N_11679,N_9129);
nand U17197 (N_17197,N_10032,N_7054);
or U17198 (N_17198,N_8929,N_11748);
nor U17199 (N_17199,N_8435,N_6355);
nor U17200 (N_17200,N_9445,N_8689);
xnor U17201 (N_17201,N_10246,N_12317);
nand U17202 (N_17202,N_8531,N_9442);
or U17203 (N_17203,N_10755,N_12340);
nor U17204 (N_17204,N_9625,N_9439);
nor U17205 (N_17205,N_11414,N_8277);
xor U17206 (N_17206,N_12258,N_8500);
or U17207 (N_17207,N_11221,N_6465);
nor U17208 (N_17208,N_11025,N_8365);
nor U17209 (N_17209,N_9735,N_10966);
nor U17210 (N_17210,N_10448,N_11523);
xor U17211 (N_17211,N_10822,N_9616);
xor U17212 (N_17212,N_11053,N_8795);
and U17213 (N_17213,N_8879,N_7722);
nand U17214 (N_17214,N_8153,N_9904);
or U17215 (N_17215,N_9639,N_9805);
xnor U17216 (N_17216,N_7927,N_6751);
nand U17217 (N_17217,N_11761,N_7023);
nand U17218 (N_17218,N_11174,N_7975);
nand U17219 (N_17219,N_11465,N_10387);
xor U17220 (N_17220,N_11916,N_10138);
xnor U17221 (N_17221,N_10528,N_6336);
nor U17222 (N_17222,N_11026,N_11926);
xor U17223 (N_17223,N_7678,N_9779);
xor U17224 (N_17224,N_6358,N_11825);
nand U17225 (N_17225,N_11670,N_7429);
xnor U17226 (N_17226,N_6993,N_9770);
nor U17227 (N_17227,N_12167,N_11203);
nand U17228 (N_17228,N_7667,N_12456);
and U17229 (N_17229,N_7548,N_10549);
or U17230 (N_17230,N_11393,N_6834);
and U17231 (N_17231,N_12377,N_7490);
nand U17232 (N_17232,N_9570,N_9837);
nor U17233 (N_17233,N_7678,N_10157);
and U17234 (N_17234,N_12082,N_8378);
nor U17235 (N_17235,N_9691,N_11317);
or U17236 (N_17236,N_7585,N_11940);
or U17237 (N_17237,N_7776,N_7987);
and U17238 (N_17238,N_9576,N_9896);
and U17239 (N_17239,N_9301,N_7556);
nand U17240 (N_17240,N_6892,N_11336);
xnor U17241 (N_17241,N_7533,N_7333);
nor U17242 (N_17242,N_9878,N_7568);
nor U17243 (N_17243,N_12173,N_10065);
and U17244 (N_17244,N_7648,N_12026);
or U17245 (N_17245,N_8304,N_6510);
nor U17246 (N_17246,N_6337,N_6790);
nand U17247 (N_17247,N_9349,N_9166);
and U17248 (N_17248,N_7452,N_8160);
or U17249 (N_17249,N_6910,N_12308);
xor U17250 (N_17250,N_8455,N_10423);
and U17251 (N_17251,N_7414,N_7632);
nand U17252 (N_17252,N_8236,N_7993);
or U17253 (N_17253,N_6637,N_9705);
nand U17254 (N_17254,N_8561,N_11665);
nor U17255 (N_17255,N_6399,N_6316);
and U17256 (N_17256,N_9752,N_10853);
nor U17257 (N_17257,N_7761,N_11198);
xnor U17258 (N_17258,N_11992,N_6691);
nor U17259 (N_17259,N_6891,N_9253);
xor U17260 (N_17260,N_11614,N_8777);
and U17261 (N_17261,N_7862,N_9763);
or U17262 (N_17262,N_8426,N_8819);
and U17263 (N_17263,N_7040,N_7747);
nor U17264 (N_17264,N_11272,N_9458);
and U17265 (N_17265,N_8140,N_11632);
nor U17266 (N_17266,N_10145,N_11307);
nand U17267 (N_17267,N_10667,N_9308);
nand U17268 (N_17268,N_9788,N_10496);
nor U17269 (N_17269,N_7477,N_8175);
and U17270 (N_17270,N_10509,N_7715);
xnor U17271 (N_17271,N_7240,N_9598);
xnor U17272 (N_17272,N_9698,N_6773);
nand U17273 (N_17273,N_9461,N_10719);
xnor U17274 (N_17274,N_8793,N_9169);
nand U17275 (N_17275,N_11751,N_8347);
or U17276 (N_17276,N_6390,N_9883);
nand U17277 (N_17277,N_6748,N_7396);
nor U17278 (N_17278,N_7191,N_9641);
nor U17279 (N_17279,N_9008,N_10741);
nand U17280 (N_17280,N_8700,N_10119);
or U17281 (N_17281,N_7134,N_10474);
nor U17282 (N_17282,N_6531,N_6466);
and U17283 (N_17283,N_10511,N_7965);
and U17284 (N_17284,N_7396,N_6300);
or U17285 (N_17285,N_6894,N_9027);
and U17286 (N_17286,N_7771,N_7986);
or U17287 (N_17287,N_11274,N_12269);
xnor U17288 (N_17288,N_10914,N_7285);
nor U17289 (N_17289,N_11029,N_11955);
nor U17290 (N_17290,N_10843,N_11735);
or U17291 (N_17291,N_11837,N_7606);
nor U17292 (N_17292,N_9277,N_7016);
or U17293 (N_17293,N_8289,N_9763);
xnor U17294 (N_17294,N_9169,N_10273);
and U17295 (N_17295,N_6491,N_8833);
xor U17296 (N_17296,N_9606,N_6737);
and U17297 (N_17297,N_9533,N_10270);
or U17298 (N_17298,N_9277,N_8527);
or U17299 (N_17299,N_6611,N_9414);
and U17300 (N_17300,N_12194,N_10184);
and U17301 (N_17301,N_7872,N_9870);
nor U17302 (N_17302,N_12060,N_8755);
nand U17303 (N_17303,N_7272,N_11572);
or U17304 (N_17304,N_7125,N_8355);
nor U17305 (N_17305,N_7539,N_10449);
or U17306 (N_17306,N_6258,N_8567);
nand U17307 (N_17307,N_11242,N_10994);
and U17308 (N_17308,N_6479,N_10104);
nor U17309 (N_17309,N_11764,N_9446);
nor U17310 (N_17310,N_11463,N_10804);
xnor U17311 (N_17311,N_10270,N_8894);
or U17312 (N_17312,N_9183,N_9986);
nand U17313 (N_17313,N_11615,N_11069);
and U17314 (N_17314,N_6964,N_7942);
xnor U17315 (N_17315,N_8588,N_6345);
nor U17316 (N_17316,N_6642,N_11607);
nand U17317 (N_17317,N_6940,N_7237);
xnor U17318 (N_17318,N_10931,N_8714);
and U17319 (N_17319,N_10003,N_7831);
xor U17320 (N_17320,N_9995,N_9523);
and U17321 (N_17321,N_12448,N_11255);
and U17322 (N_17322,N_11544,N_6707);
and U17323 (N_17323,N_10500,N_8715);
or U17324 (N_17324,N_9504,N_12019);
nor U17325 (N_17325,N_11660,N_11930);
nor U17326 (N_17326,N_6942,N_10379);
nand U17327 (N_17327,N_8975,N_11021);
and U17328 (N_17328,N_10933,N_7954);
xnor U17329 (N_17329,N_7988,N_6735);
nor U17330 (N_17330,N_12307,N_9682);
xnor U17331 (N_17331,N_6403,N_7610);
and U17332 (N_17332,N_7508,N_7759);
nor U17333 (N_17333,N_9249,N_7866);
or U17334 (N_17334,N_6852,N_10122);
or U17335 (N_17335,N_10668,N_9639);
or U17336 (N_17336,N_11765,N_11321);
or U17337 (N_17337,N_6497,N_10717);
nor U17338 (N_17338,N_8959,N_11599);
and U17339 (N_17339,N_8855,N_9382);
xnor U17340 (N_17340,N_11018,N_9832);
nand U17341 (N_17341,N_8411,N_8470);
or U17342 (N_17342,N_11409,N_9853);
or U17343 (N_17343,N_7015,N_12091);
nand U17344 (N_17344,N_6371,N_10049);
and U17345 (N_17345,N_12311,N_10641);
or U17346 (N_17346,N_7941,N_11068);
nor U17347 (N_17347,N_7677,N_7266);
nand U17348 (N_17348,N_7626,N_9734);
nor U17349 (N_17349,N_8681,N_7216);
xnor U17350 (N_17350,N_12372,N_11215);
nand U17351 (N_17351,N_8128,N_12265);
nand U17352 (N_17352,N_10838,N_11017);
or U17353 (N_17353,N_6462,N_9227);
and U17354 (N_17354,N_11623,N_8217);
nor U17355 (N_17355,N_10238,N_11980);
nor U17356 (N_17356,N_6763,N_8117);
nand U17357 (N_17357,N_7036,N_7353);
and U17358 (N_17358,N_8992,N_10723);
nor U17359 (N_17359,N_9445,N_9229);
and U17360 (N_17360,N_9770,N_10448);
xnor U17361 (N_17361,N_9453,N_8200);
or U17362 (N_17362,N_6551,N_10180);
nor U17363 (N_17363,N_7447,N_9376);
nor U17364 (N_17364,N_10670,N_10491);
xnor U17365 (N_17365,N_9674,N_8627);
nor U17366 (N_17366,N_8131,N_12391);
nor U17367 (N_17367,N_11328,N_11180);
xnor U17368 (N_17368,N_7324,N_6425);
nand U17369 (N_17369,N_9282,N_7061);
or U17370 (N_17370,N_9608,N_6902);
and U17371 (N_17371,N_7154,N_9201);
or U17372 (N_17372,N_8984,N_12014);
nor U17373 (N_17373,N_9510,N_11766);
and U17374 (N_17374,N_7891,N_10949);
or U17375 (N_17375,N_12380,N_11995);
nor U17376 (N_17376,N_9643,N_10004);
or U17377 (N_17377,N_8778,N_11916);
nor U17378 (N_17378,N_7195,N_10774);
nand U17379 (N_17379,N_9306,N_9894);
nand U17380 (N_17380,N_7472,N_8291);
xnor U17381 (N_17381,N_6805,N_10270);
and U17382 (N_17382,N_10575,N_12289);
and U17383 (N_17383,N_9308,N_7274);
nand U17384 (N_17384,N_11433,N_11636);
nand U17385 (N_17385,N_11797,N_11281);
nor U17386 (N_17386,N_10013,N_8961);
and U17387 (N_17387,N_9053,N_7649);
or U17388 (N_17388,N_12255,N_6418);
nand U17389 (N_17389,N_8402,N_7687);
or U17390 (N_17390,N_8405,N_10276);
or U17391 (N_17391,N_10046,N_11558);
or U17392 (N_17392,N_6998,N_10417);
xor U17393 (N_17393,N_8027,N_10281);
and U17394 (N_17394,N_11174,N_8445);
nand U17395 (N_17395,N_8789,N_9496);
xor U17396 (N_17396,N_6366,N_9376);
or U17397 (N_17397,N_12494,N_8632);
nand U17398 (N_17398,N_6662,N_6726);
nand U17399 (N_17399,N_11071,N_12376);
nor U17400 (N_17400,N_7024,N_11942);
nor U17401 (N_17401,N_12075,N_9945);
and U17402 (N_17402,N_10973,N_11677);
nor U17403 (N_17403,N_6344,N_11591);
nor U17404 (N_17404,N_9684,N_11086);
nand U17405 (N_17405,N_10834,N_8812);
nor U17406 (N_17406,N_10037,N_8184);
nand U17407 (N_17407,N_7817,N_7175);
nand U17408 (N_17408,N_7995,N_8256);
nand U17409 (N_17409,N_6908,N_7051);
nor U17410 (N_17410,N_7535,N_6971);
xor U17411 (N_17411,N_7197,N_8228);
nor U17412 (N_17412,N_12167,N_11904);
xor U17413 (N_17413,N_9081,N_9201);
xor U17414 (N_17414,N_9003,N_10960);
nand U17415 (N_17415,N_11915,N_10846);
and U17416 (N_17416,N_10377,N_10564);
nand U17417 (N_17417,N_6877,N_10382);
nor U17418 (N_17418,N_11746,N_8691);
nand U17419 (N_17419,N_7466,N_9702);
xor U17420 (N_17420,N_8295,N_6300);
xor U17421 (N_17421,N_8098,N_8707);
xnor U17422 (N_17422,N_8623,N_7678);
and U17423 (N_17423,N_7943,N_8736);
nor U17424 (N_17424,N_11428,N_9924);
and U17425 (N_17425,N_6913,N_7437);
or U17426 (N_17426,N_7069,N_8041);
nand U17427 (N_17427,N_11171,N_10156);
nand U17428 (N_17428,N_7625,N_9295);
or U17429 (N_17429,N_10628,N_6530);
xor U17430 (N_17430,N_8883,N_11756);
xor U17431 (N_17431,N_8585,N_11184);
nand U17432 (N_17432,N_7345,N_11807);
or U17433 (N_17433,N_10719,N_8036);
xnor U17434 (N_17434,N_9211,N_6907);
nand U17435 (N_17435,N_6714,N_6622);
xor U17436 (N_17436,N_10280,N_11460);
nand U17437 (N_17437,N_10783,N_10972);
nor U17438 (N_17438,N_9122,N_7070);
nor U17439 (N_17439,N_6565,N_11164);
nand U17440 (N_17440,N_8979,N_6445);
and U17441 (N_17441,N_8834,N_11042);
and U17442 (N_17442,N_10883,N_9515);
nand U17443 (N_17443,N_10568,N_8586);
or U17444 (N_17444,N_6413,N_8126);
or U17445 (N_17445,N_11891,N_8933);
nor U17446 (N_17446,N_10294,N_7645);
nor U17447 (N_17447,N_7854,N_8097);
nor U17448 (N_17448,N_6532,N_11436);
nor U17449 (N_17449,N_6350,N_6544);
nand U17450 (N_17450,N_7920,N_10611);
and U17451 (N_17451,N_6595,N_11331);
xor U17452 (N_17452,N_6291,N_11617);
or U17453 (N_17453,N_10615,N_12048);
nor U17454 (N_17454,N_8810,N_11428);
xor U17455 (N_17455,N_12415,N_7333);
or U17456 (N_17456,N_6986,N_10953);
or U17457 (N_17457,N_11370,N_11571);
nand U17458 (N_17458,N_11723,N_11155);
nor U17459 (N_17459,N_9956,N_7445);
xnor U17460 (N_17460,N_8332,N_11249);
xor U17461 (N_17461,N_11765,N_10869);
nor U17462 (N_17462,N_10431,N_10646);
nor U17463 (N_17463,N_9830,N_7435);
nor U17464 (N_17464,N_11626,N_6495);
nor U17465 (N_17465,N_12112,N_11245);
nor U17466 (N_17466,N_11315,N_6572);
and U17467 (N_17467,N_7756,N_6347);
nand U17468 (N_17468,N_12287,N_9373);
and U17469 (N_17469,N_10956,N_11022);
and U17470 (N_17470,N_6763,N_10039);
xor U17471 (N_17471,N_10893,N_8907);
or U17472 (N_17472,N_9034,N_11742);
or U17473 (N_17473,N_12359,N_6876);
nor U17474 (N_17474,N_8013,N_9512);
and U17475 (N_17475,N_9656,N_9714);
xnor U17476 (N_17476,N_8415,N_7447);
and U17477 (N_17477,N_11946,N_9596);
xnor U17478 (N_17478,N_7046,N_9711);
xor U17479 (N_17479,N_10722,N_6857);
and U17480 (N_17480,N_12143,N_12437);
or U17481 (N_17481,N_9221,N_11508);
and U17482 (N_17482,N_11794,N_11693);
nor U17483 (N_17483,N_8741,N_10899);
nor U17484 (N_17484,N_8632,N_8036);
nor U17485 (N_17485,N_8083,N_8667);
nand U17486 (N_17486,N_11415,N_11983);
and U17487 (N_17487,N_8382,N_9338);
nand U17488 (N_17488,N_11480,N_12437);
xor U17489 (N_17489,N_8816,N_11091);
or U17490 (N_17490,N_8757,N_9760);
or U17491 (N_17491,N_6942,N_6788);
nor U17492 (N_17492,N_10282,N_11323);
or U17493 (N_17493,N_7472,N_6921);
xor U17494 (N_17494,N_7701,N_11848);
xor U17495 (N_17495,N_11621,N_11963);
and U17496 (N_17496,N_11097,N_10728);
xor U17497 (N_17497,N_9528,N_11396);
or U17498 (N_17498,N_12108,N_12165);
nand U17499 (N_17499,N_9267,N_7960);
and U17500 (N_17500,N_10911,N_10694);
xor U17501 (N_17501,N_9435,N_10774);
and U17502 (N_17502,N_8058,N_7279);
nand U17503 (N_17503,N_10891,N_8299);
nand U17504 (N_17504,N_10216,N_7069);
or U17505 (N_17505,N_8217,N_10691);
xnor U17506 (N_17506,N_6644,N_11113);
nor U17507 (N_17507,N_9377,N_8516);
nor U17508 (N_17508,N_6905,N_7324);
nand U17509 (N_17509,N_7208,N_11759);
nor U17510 (N_17510,N_6519,N_9874);
nand U17511 (N_17511,N_8035,N_7059);
or U17512 (N_17512,N_6866,N_8196);
xnor U17513 (N_17513,N_9875,N_8991);
and U17514 (N_17514,N_7379,N_11050);
or U17515 (N_17515,N_11918,N_7515);
or U17516 (N_17516,N_12086,N_11874);
nor U17517 (N_17517,N_12370,N_7728);
and U17518 (N_17518,N_8099,N_10443);
nand U17519 (N_17519,N_12420,N_10553);
or U17520 (N_17520,N_7573,N_9577);
or U17521 (N_17521,N_10064,N_9369);
or U17522 (N_17522,N_6482,N_11305);
or U17523 (N_17523,N_7891,N_6545);
or U17524 (N_17524,N_9894,N_8406);
nor U17525 (N_17525,N_11542,N_6527);
and U17526 (N_17526,N_8910,N_8530);
and U17527 (N_17527,N_10398,N_7744);
and U17528 (N_17528,N_11522,N_9265);
and U17529 (N_17529,N_12058,N_10075);
and U17530 (N_17530,N_12135,N_6665);
xor U17531 (N_17531,N_11638,N_11001);
nand U17532 (N_17532,N_7028,N_6717);
and U17533 (N_17533,N_8476,N_7793);
or U17534 (N_17534,N_11104,N_7518);
and U17535 (N_17535,N_8898,N_8346);
xnor U17536 (N_17536,N_9755,N_7446);
nand U17537 (N_17537,N_10832,N_11360);
nand U17538 (N_17538,N_11245,N_10439);
or U17539 (N_17539,N_6287,N_9859);
nand U17540 (N_17540,N_6822,N_6549);
or U17541 (N_17541,N_11357,N_10041);
xor U17542 (N_17542,N_12103,N_8937);
nor U17543 (N_17543,N_11676,N_9431);
and U17544 (N_17544,N_12161,N_6954);
nand U17545 (N_17545,N_12024,N_12015);
nor U17546 (N_17546,N_6588,N_11539);
xnor U17547 (N_17547,N_9964,N_10811);
nand U17548 (N_17548,N_6782,N_7208);
nand U17549 (N_17549,N_9434,N_12339);
nand U17550 (N_17550,N_8041,N_10214);
nor U17551 (N_17551,N_10564,N_10233);
or U17552 (N_17552,N_7356,N_8343);
xnor U17553 (N_17553,N_7011,N_11893);
xor U17554 (N_17554,N_7302,N_9510);
and U17555 (N_17555,N_12317,N_10137);
nand U17556 (N_17556,N_9243,N_7696);
and U17557 (N_17557,N_11274,N_8940);
nand U17558 (N_17558,N_7101,N_12247);
or U17559 (N_17559,N_7293,N_7304);
or U17560 (N_17560,N_6906,N_9967);
nand U17561 (N_17561,N_10509,N_10352);
or U17562 (N_17562,N_10494,N_8215);
xnor U17563 (N_17563,N_6256,N_7429);
nand U17564 (N_17564,N_7514,N_6365);
and U17565 (N_17565,N_8467,N_10446);
xnor U17566 (N_17566,N_9509,N_7267);
nor U17567 (N_17567,N_6521,N_8788);
nand U17568 (N_17568,N_6703,N_12361);
or U17569 (N_17569,N_7675,N_6296);
or U17570 (N_17570,N_9530,N_8951);
and U17571 (N_17571,N_8687,N_7735);
xor U17572 (N_17572,N_8275,N_8335);
or U17573 (N_17573,N_6788,N_8460);
or U17574 (N_17574,N_11332,N_11877);
xor U17575 (N_17575,N_9241,N_7476);
or U17576 (N_17576,N_9481,N_6822);
and U17577 (N_17577,N_6353,N_6271);
nor U17578 (N_17578,N_6798,N_12218);
or U17579 (N_17579,N_10058,N_12217);
xor U17580 (N_17580,N_9832,N_8045);
or U17581 (N_17581,N_7307,N_11676);
nand U17582 (N_17582,N_10945,N_11631);
and U17583 (N_17583,N_6343,N_11865);
nor U17584 (N_17584,N_7531,N_12200);
xnor U17585 (N_17585,N_6273,N_10169);
nor U17586 (N_17586,N_8609,N_7741);
xnor U17587 (N_17587,N_12463,N_6994);
xnor U17588 (N_17588,N_12301,N_9892);
and U17589 (N_17589,N_8686,N_10582);
nor U17590 (N_17590,N_9337,N_7797);
and U17591 (N_17591,N_11600,N_10407);
nor U17592 (N_17592,N_7967,N_10765);
nand U17593 (N_17593,N_9902,N_7569);
xor U17594 (N_17594,N_9390,N_8327);
and U17595 (N_17595,N_12498,N_9221);
nand U17596 (N_17596,N_7938,N_11035);
nand U17597 (N_17597,N_11329,N_11986);
and U17598 (N_17598,N_7564,N_9624);
nor U17599 (N_17599,N_12223,N_12198);
nand U17600 (N_17600,N_7577,N_6789);
nor U17601 (N_17601,N_11712,N_6976);
xnor U17602 (N_17602,N_8694,N_12340);
or U17603 (N_17603,N_10099,N_10233);
and U17604 (N_17604,N_8957,N_11121);
xnor U17605 (N_17605,N_8221,N_7967);
or U17606 (N_17606,N_7472,N_11003);
or U17607 (N_17607,N_11982,N_9519);
nand U17608 (N_17608,N_11021,N_8554);
nor U17609 (N_17609,N_11433,N_11142);
or U17610 (N_17610,N_6404,N_9206);
nor U17611 (N_17611,N_6427,N_8387);
xnor U17612 (N_17612,N_8679,N_11150);
nand U17613 (N_17613,N_11843,N_7454);
or U17614 (N_17614,N_6737,N_11831);
xnor U17615 (N_17615,N_9719,N_8399);
xnor U17616 (N_17616,N_9152,N_11109);
nand U17617 (N_17617,N_7264,N_11045);
and U17618 (N_17618,N_10019,N_7485);
nor U17619 (N_17619,N_11547,N_9774);
nand U17620 (N_17620,N_9160,N_8215);
nor U17621 (N_17621,N_9886,N_6736);
or U17622 (N_17622,N_11810,N_10004);
nand U17623 (N_17623,N_9661,N_6442);
xor U17624 (N_17624,N_7310,N_9348);
and U17625 (N_17625,N_10027,N_7370);
xor U17626 (N_17626,N_11175,N_8211);
nand U17627 (N_17627,N_8995,N_11748);
or U17628 (N_17628,N_9516,N_12436);
nand U17629 (N_17629,N_9818,N_9602);
nor U17630 (N_17630,N_8618,N_7097);
and U17631 (N_17631,N_7408,N_11326);
xnor U17632 (N_17632,N_10532,N_7156);
xnor U17633 (N_17633,N_8319,N_12045);
nor U17634 (N_17634,N_8394,N_6525);
or U17635 (N_17635,N_6796,N_6879);
and U17636 (N_17636,N_6298,N_8967);
xnor U17637 (N_17637,N_12431,N_7262);
nand U17638 (N_17638,N_8269,N_8055);
xnor U17639 (N_17639,N_7937,N_8382);
or U17640 (N_17640,N_12476,N_10505);
nand U17641 (N_17641,N_10478,N_10113);
nor U17642 (N_17642,N_10640,N_7061);
and U17643 (N_17643,N_12154,N_12263);
xnor U17644 (N_17644,N_10729,N_11188);
xnor U17645 (N_17645,N_11103,N_8338);
nand U17646 (N_17646,N_7372,N_10536);
xor U17647 (N_17647,N_12102,N_12204);
and U17648 (N_17648,N_9514,N_7705);
or U17649 (N_17649,N_8562,N_11825);
and U17650 (N_17650,N_11785,N_10741);
or U17651 (N_17651,N_8152,N_11420);
or U17652 (N_17652,N_9470,N_10996);
xnor U17653 (N_17653,N_7624,N_9261);
and U17654 (N_17654,N_8657,N_6512);
xnor U17655 (N_17655,N_8420,N_11656);
nand U17656 (N_17656,N_12376,N_11820);
xor U17657 (N_17657,N_8859,N_9405);
or U17658 (N_17658,N_10331,N_9057);
or U17659 (N_17659,N_8759,N_6719);
or U17660 (N_17660,N_6773,N_6466);
or U17661 (N_17661,N_11277,N_7793);
nor U17662 (N_17662,N_12291,N_9619);
and U17663 (N_17663,N_7283,N_8901);
nand U17664 (N_17664,N_11377,N_12360);
or U17665 (N_17665,N_10354,N_12473);
xnor U17666 (N_17666,N_8077,N_11981);
or U17667 (N_17667,N_11034,N_12325);
nand U17668 (N_17668,N_10503,N_7902);
nor U17669 (N_17669,N_11529,N_11422);
nand U17670 (N_17670,N_11464,N_7761);
or U17671 (N_17671,N_7219,N_6561);
nand U17672 (N_17672,N_10019,N_9196);
or U17673 (N_17673,N_8886,N_7382);
and U17674 (N_17674,N_12235,N_10708);
nand U17675 (N_17675,N_10313,N_9653);
and U17676 (N_17676,N_12362,N_9701);
xor U17677 (N_17677,N_7742,N_11648);
nand U17678 (N_17678,N_7059,N_12469);
nand U17679 (N_17679,N_8614,N_8381);
or U17680 (N_17680,N_8090,N_12059);
and U17681 (N_17681,N_11204,N_12064);
and U17682 (N_17682,N_6812,N_6489);
nor U17683 (N_17683,N_9580,N_8036);
nor U17684 (N_17684,N_12247,N_9097);
nand U17685 (N_17685,N_8619,N_7773);
xor U17686 (N_17686,N_10267,N_6633);
nor U17687 (N_17687,N_7029,N_9378);
and U17688 (N_17688,N_11292,N_9743);
or U17689 (N_17689,N_9955,N_9265);
nor U17690 (N_17690,N_10194,N_6877);
nor U17691 (N_17691,N_10221,N_9634);
nand U17692 (N_17692,N_7509,N_10452);
xnor U17693 (N_17693,N_11937,N_11416);
xnor U17694 (N_17694,N_7846,N_12210);
or U17695 (N_17695,N_11743,N_10827);
and U17696 (N_17696,N_6340,N_8092);
or U17697 (N_17697,N_6272,N_8516);
nor U17698 (N_17698,N_7526,N_11257);
nor U17699 (N_17699,N_6286,N_8551);
and U17700 (N_17700,N_12108,N_10917);
xor U17701 (N_17701,N_12062,N_11993);
or U17702 (N_17702,N_9125,N_11118);
and U17703 (N_17703,N_8042,N_8735);
and U17704 (N_17704,N_10275,N_10019);
nor U17705 (N_17705,N_6886,N_8051);
or U17706 (N_17706,N_8502,N_9461);
nand U17707 (N_17707,N_9006,N_9651);
nor U17708 (N_17708,N_7982,N_7955);
xor U17709 (N_17709,N_10932,N_11090);
and U17710 (N_17710,N_10424,N_10105);
xnor U17711 (N_17711,N_8982,N_8405);
nand U17712 (N_17712,N_6313,N_9064);
xor U17713 (N_17713,N_11899,N_7048);
or U17714 (N_17714,N_6564,N_7593);
xnor U17715 (N_17715,N_7935,N_6872);
nand U17716 (N_17716,N_11383,N_7532);
and U17717 (N_17717,N_12467,N_12073);
xnor U17718 (N_17718,N_12274,N_8178);
nand U17719 (N_17719,N_6459,N_6352);
or U17720 (N_17720,N_9108,N_10729);
or U17721 (N_17721,N_11993,N_8411);
xnor U17722 (N_17722,N_7298,N_6365);
nor U17723 (N_17723,N_7589,N_7992);
xnor U17724 (N_17724,N_10189,N_8195);
and U17725 (N_17725,N_9411,N_11408);
and U17726 (N_17726,N_11482,N_8291);
and U17727 (N_17727,N_12167,N_7812);
and U17728 (N_17728,N_11046,N_11217);
and U17729 (N_17729,N_7566,N_10887);
and U17730 (N_17730,N_8127,N_11297);
nor U17731 (N_17731,N_6255,N_8188);
nor U17732 (N_17732,N_10792,N_7671);
and U17733 (N_17733,N_11527,N_7622);
nand U17734 (N_17734,N_11560,N_11675);
nor U17735 (N_17735,N_9566,N_9722);
and U17736 (N_17736,N_8520,N_11475);
xor U17737 (N_17737,N_9435,N_8871);
nand U17738 (N_17738,N_12061,N_7891);
or U17739 (N_17739,N_11832,N_6761);
and U17740 (N_17740,N_8589,N_10213);
nand U17741 (N_17741,N_6789,N_11623);
or U17742 (N_17742,N_8627,N_6843);
or U17743 (N_17743,N_7049,N_8673);
nor U17744 (N_17744,N_7141,N_7497);
nor U17745 (N_17745,N_9127,N_7032);
and U17746 (N_17746,N_12397,N_8550);
nor U17747 (N_17747,N_11721,N_10571);
nand U17748 (N_17748,N_11510,N_8632);
or U17749 (N_17749,N_11339,N_12482);
xor U17750 (N_17750,N_10298,N_8181);
and U17751 (N_17751,N_10830,N_8725);
or U17752 (N_17752,N_9678,N_7326);
or U17753 (N_17753,N_10695,N_8744);
nor U17754 (N_17754,N_6855,N_6804);
xor U17755 (N_17755,N_9621,N_11160);
or U17756 (N_17756,N_7082,N_6333);
or U17757 (N_17757,N_7144,N_12137);
and U17758 (N_17758,N_11060,N_12187);
and U17759 (N_17759,N_8885,N_9897);
nor U17760 (N_17760,N_9934,N_7916);
nand U17761 (N_17761,N_11108,N_8899);
nand U17762 (N_17762,N_9483,N_11599);
or U17763 (N_17763,N_7127,N_9208);
nand U17764 (N_17764,N_6876,N_11121);
xor U17765 (N_17765,N_10794,N_8281);
and U17766 (N_17766,N_9846,N_11616);
and U17767 (N_17767,N_12154,N_8899);
nor U17768 (N_17768,N_9592,N_11742);
and U17769 (N_17769,N_9610,N_9662);
or U17770 (N_17770,N_11765,N_7887);
and U17771 (N_17771,N_9760,N_6357);
nor U17772 (N_17772,N_10725,N_6533);
nor U17773 (N_17773,N_9654,N_9478);
and U17774 (N_17774,N_7039,N_10735);
nor U17775 (N_17775,N_7879,N_8088);
xnor U17776 (N_17776,N_8903,N_12369);
and U17777 (N_17777,N_7053,N_7326);
xor U17778 (N_17778,N_6446,N_8586);
xor U17779 (N_17779,N_8321,N_11122);
or U17780 (N_17780,N_11829,N_7158);
nand U17781 (N_17781,N_10293,N_11314);
or U17782 (N_17782,N_6487,N_11380);
nand U17783 (N_17783,N_7950,N_12425);
nand U17784 (N_17784,N_7172,N_8298);
nand U17785 (N_17785,N_12277,N_7339);
xor U17786 (N_17786,N_7232,N_7257);
nor U17787 (N_17787,N_7946,N_11130);
and U17788 (N_17788,N_9412,N_10879);
nand U17789 (N_17789,N_6546,N_11156);
nor U17790 (N_17790,N_6449,N_10417);
or U17791 (N_17791,N_6514,N_8826);
xnor U17792 (N_17792,N_10400,N_8667);
or U17793 (N_17793,N_7491,N_9239);
or U17794 (N_17794,N_8131,N_8158);
or U17795 (N_17795,N_8104,N_11107);
xor U17796 (N_17796,N_8617,N_9825);
nand U17797 (N_17797,N_9181,N_8865);
xnor U17798 (N_17798,N_8288,N_12163);
or U17799 (N_17799,N_9246,N_8240);
and U17800 (N_17800,N_6605,N_7564);
and U17801 (N_17801,N_8903,N_8917);
nor U17802 (N_17802,N_10285,N_7799);
xnor U17803 (N_17803,N_9561,N_8636);
nand U17804 (N_17804,N_6591,N_11482);
or U17805 (N_17805,N_8090,N_12419);
or U17806 (N_17806,N_9919,N_10525);
or U17807 (N_17807,N_12193,N_7483);
and U17808 (N_17808,N_7019,N_11622);
nand U17809 (N_17809,N_7042,N_6412);
and U17810 (N_17810,N_9268,N_7597);
nor U17811 (N_17811,N_10273,N_11434);
or U17812 (N_17812,N_7988,N_8761);
or U17813 (N_17813,N_9999,N_7766);
xor U17814 (N_17814,N_11660,N_6726);
or U17815 (N_17815,N_6643,N_6362);
nor U17816 (N_17816,N_6608,N_10283);
nand U17817 (N_17817,N_11633,N_10445);
or U17818 (N_17818,N_12190,N_11120);
and U17819 (N_17819,N_6843,N_6289);
and U17820 (N_17820,N_7512,N_10404);
and U17821 (N_17821,N_8473,N_11906);
and U17822 (N_17822,N_7257,N_11816);
xnor U17823 (N_17823,N_8887,N_8047);
nand U17824 (N_17824,N_11092,N_11742);
or U17825 (N_17825,N_8523,N_10224);
or U17826 (N_17826,N_7476,N_9139);
nand U17827 (N_17827,N_12253,N_6515);
and U17828 (N_17828,N_10265,N_9471);
nor U17829 (N_17829,N_7735,N_10712);
nor U17830 (N_17830,N_7642,N_11272);
xnor U17831 (N_17831,N_10381,N_8957);
xnor U17832 (N_17832,N_7424,N_11826);
nor U17833 (N_17833,N_7215,N_9459);
or U17834 (N_17834,N_7829,N_7639);
xor U17835 (N_17835,N_9739,N_10969);
xor U17836 (N_17836,N_7782,N_8751);
and U17837 (N_17837,N_11451,N_11922);
or U17838 (N_17838,N_7814,N_8322);
or U17839 (N_17839,N_6752,N_9388);
or U17840 (N_17840,N_9549,N_7149);
nand U17841 (N_17841,N_7901,N_12025);
nor U17842 (N_17842,N_8056,N_7878);
nor U17843 (N_17843,N_6553,N_6580);
or U17844 (N_17844,N_9482,N_8173);
and U17845 (N_17845,N_6345,N_8099);
nand U17846 (N_17846,N_11077,N_10220);
nand U17847 (N_17847,N_11709,N_9895);
nor U17848 (N_17848,N_7558,N_10584);
and U17849 (N_17849,N_8834,N_8653);
and U17850 (N_17850,N_12212,N_7815);
xor U17851 (N_17851,N_11257,N_9605);
and U17852 (N_17852,N_9065,N_10156);
xnor U17853 (N_17853,N_9763,N_10455);
nor U17854 (N_17854,N_11378,N_11615);
and U17855 (N_17855,N_8851,N_11501);
xnor U17856 (N_17856,N_10185,N_8536);
or U17857 (N_17857,N_8523,N_11463);
xnor U17858 (N_17858,N_9712,N_6414);
nand U17859 (N_17859,N_10283,N_7513);
and U17860 (N_17860,N_6411,N_10720);
or U17861 (N_17861,N_6513,N_11917);
nor U17862 (N_17862,N_12292,N_7084);
xor U17863 (N_17863,N_9134,N_7982);
or U17864 (N_17864,N_10210,N_10891);
or U17865 (N_17865,N_8675,N_8757);
or U17866 (N_17866,N_9000,N_8422);
nor U17867 (N_17867,N_10945,N_10605);
or U17868 (N_17868,N_9515,N_7399);
nand U17869 (N_17869,N_8728,N_8255);
nand U17870 (N_17870,N_9166,N_11250);
nor U17871 (N_17871,N_9295,N_9261);
and U17872 (N_17872,N_7872,N_9745);
xnor U17873 (N_17873,N_11410,N_9121);
xnor U17874 (N_17874,N_7665,N_7575);
nor U17875 (N_17875,N_12238,N_11802);
and U17876 (N_17876,N_9310,N_12393);
and U17877 (N_17877,N_7378,N_8179);
or U17878 (N_17878,N_8582,N_8000);
nand U17879 (N_17879,N_7698,N_11811);
xor U17880 (N_17880,N_8167,N_9271);
nand U17881 (N_17881,N_10126,N_11476);
and U17882 (N_17882,N_8791,N_10267);
nand U17883 (N_17883,N_6347,N_8898);
or U17884 (N_17884,N_9544,N_11709);
or U17885 (N_17885,N_8206,N_10121);
xor U17886 (N_17886,N_10887,N_9622);
or U17887 (N_17887,N_11333,N_7028);
nand U17888 (N_17888,N_6605,N_9175);
nand U17889 (N_17889,N_11624,N_8542);
nor U17890 (N_17890,N_10208,N_10405);
nand U17891 (N_17891,N_9426,N_10089);
and U17892 (N_17892,N_10266,N_12493);
and U17893 (N_17893,N_10544,N_6281);
or U17894 (N_17894,N_9069,N_7375);
nand U17895 (N_17895,N_7733,N_9013);
and U17896 (N_17896,N_8730,N_10390);
xor U17897 (N_17897,N_7473,N_9422);
xor U17898 (N_17898,N_6989,N_8376);
and U17899 (N_17899,N_9020,N_6516);
xor U17900 (N_17900,N_7627,N_9378);
and U17901 (N_17901,N_11333,N_6455);
and U17902 (N_17902,N_11358,N_7136);
xnor U17903 (N_17903,N_11812,N_8616);
xnor U17904 (N_17904,N_8512,N_9833);
and U17905 (N_17905,N_8633,N_8315);
and U17906 (N_17906,N_6972,N_7394);
nor U17907 (N_17907,N_12089,N_10390);
nor U17908 (N_17908,N_10552,N_7293);
nand U17909 (N_17909,N_8144,N_6683);
nor U17910 (N_17910,N_8281,N_7839);
and U17911 (N_17911,N_12375,N_10465);
nor U17912 (N_17912,N_8479,N_11525);
nand U17913 (N_17913,N_10546,N_8328);
xor U17914 (N_17914,N_7965,N_8102);
xor U17915 (N_17915,N_9565,N_10528);
xnor U17916 (N_17916,N_9156,N_8256);
or U17917 (N_17917,N_10611,N_10327);
nand U17918 (N_17918,N_10483,N_10610);
nor U17919 (N_17919,N_12471,N_8891);
nand U17920 (N_17920,N_8317,N_12098);
nor U17921 (N_17921,N_11714,N_9389);
and U17922 (N_17922,N_12321,N_9853);
nor U17923 (N_17923,N_7938,N_11532);
or U17924 (N_17924,N_7022,N_11859);
and U17925 (N_17925,N_9602,N_7721);
xor U17926 (N_17926,N_11418,N_7338);
nand U17927 (N_17927,N_7440,N_7214);
and U17928 (N_17928,N_8980,N_6456);
xor U17929 (N_17929,N_9727,N_8408);
and U17930 (N_17930,N_7465,N_12209);
xnor U17931 (N_17931,N_9356,N_8249);
xnor U17932 (N_17932,N_6344,N_12391);
nand U17933 (N_17933,N_12077,N_9270);
and U17934 (N_17934,N_6964,N_10974);
or U17935 (N_17935,N_8263,N_8255);
nor U17936 (N_17936,N_12349,N_8601);
or U17937 (N_17937,N_9245,N_6707);
xor U17938 (N_17938,N_7257,N_9681);
nand U17939 (N_17939,N_8178,N_8430);
and U17940 (N_17940,N_7941,N_11525);
xnor U17941 (N_17941,N_11172,N_10554);
nor U17942 (N_17942,N_9790,N_7300);
nor U17943 (N_17943,N_10436,N_7575);
nand U17944 (N_17944,N_9565,N_11998);
nor U17945 (N_17945,N_12149,N_9950);
or U17946 (N_17946,N_9522,N_10270);
nor U17947 (N_17947,N_7624,N_10382);
nor U17948 (N_17948,N_11233,N_8183);
or U17949 (N_17949,N_11601,N_10150);
and U17950 (N_17950,N_11161,N_11054);
or U17951 (N_17951,N_11810,N_7110);
nand U17952 (N_17952,N_11995,N_10581);
and U17953 (N_17953,N_9141,N_8881);
or U17954 (N_17954,N_12078,N_12124);
nand U17955 (N_17955,N_9478,N_7140);
or U17956 (N_17956,N_8086,N_12292);
nor U17957 (N_17957,N_7091,N_7589);
or U17958 (N_17958,N_10959,N_6327);
or U17959 (N_17959,N_11038,N_11123);
nor U17960 (N_17960,N_10144,N_11854);
xor U17961 (N_17961,N_7372,N_11999);
xor U17962 (N_17962,N_7588,N_10769);
xor U17963 (N_17963,N_8912,N_6676);
nor U17964 (N_17964,N_8299,N_8030);
nand U17965 (N_17965,N_6990,N_12303);
xor U17966 (N_17966,N_8567,N_7524);
and U17967 (N_17967,N_12239,N_9956);
xor U17968 (N_17968,N_6902,N_7617);
nor U17969 (N_17969,N_10931,N_6602);
or U17970 (N_17970,N_12010,N_11677);
or U17971 (N_17971,N_7092,N_7014);
and U17972 (N_17972,N_11547,N_8198);
and U17973 (N_17973,N_10482,N_10808);
or U17974 (N_17974,N_11912,N_10870);
nor U17975 (N_17975,N_7418,N_7336);
nand U17976 (N_17976,N_8570,N_6685);
xnor U17977 (N_17977,N_11952,N_10171);
xnor U17978 (N_17978,N_7189,N_8194);
nor U17979 (N_17979,N_7053,N_10207);
nand U17980 (N_17980,N_11810,N_10257);
nor U17981 (N_17981,N_9194,N_10402);
xnor U17982 (N_17982,N_6752,N_8357);
nand U17983 (N_17983,N_11950,N_7853);
and U17984 (N_17984,N_6279,N_9695);
nor U17985 (N_17985,N_8822,N_10279);
and U17986 (N_17986,N_9101,N_10085);
nor U17987 (N_17987,N_8032,N_8554);
and U17988 (N_17988,N_8088,N_8805);
or U17989 (N_17989,N_11743,N_7626);
nor U17990 (N_17990,N_10217,N_8860);
or U17991 (N_17991,N_8471,N_7115);
xnor U17992 (N_17992,N_10989,N_6637);
or U17993 (N_17993,N_8250,N_12254);
nor U17994 (N_17994,N_9409,N_10344);
nand U17995 (N_17995,N_7173,N_11861);
and U17996 (N_17996,N_9623,N_8475);
nand U17997 (N_17997,N_8262,N_10052);
or U17998 (N_17998,N_9034,N_11138);
nor U17999 (N_17999,N_7062,N_7348);
and U18000 (N_18000,N_9179,N_6839);
nor U18001 (N_18001,N_9706,N_10072);
nor U18002 (N_18002,N_8833,N_11380);
nor U18003 (N_18003,N_8872,N_9823);
xor U18004 (N_18004,N_8632,N_10514);
nand U18005 (N_18005,N_10775,N_8080);
or U18006 (N_18006,N_8638,N_8952);
and U18007 (N_18007,N_10804,N_8136);
nor U18008 (N_18008,N_7476,N_9208);
or U18009 (N_18009,N_8775,N_11414);
nor U18010 (N_18010,N_9221,N_10680);
nand U18011 (N_18011,N_12175,N_8458);
xnor U18012 (N_18012,N_10348,N_7098);
xor U18013 (N_18013,N_8984,N_7464);
nor U18014 (N_18014,N_9015,N_7570);
nand U18015 (N_18015,N_8766,N_9614);
or U18016 (N_18016,N_6252,N_11633);
nor U18017 (N_18017,N_11162,N_8966);
or U18018 (N_18018,N_10578,N_8198);
nor U18019 (N_18019,N_6358,N_11208);
nor U18020 (N_18020,N_11604,N_8434);
or U18021 (N_18021,N_7747,N_11068);
nor U18022 (N_18022,N_11709,N_6367);
nand U18023 (N_18023,N_8661,N_7451);
nor U18024 (N_18024,N_9347,N_6373);
and U18025 (N_18025,N_11755,N_10643);
and U18026 (N_18026,N_7620,N_10087);
and U18027 (N_18027,N_10208,N_7185);
nor U18028 (N_18028,N_6525,N_9394);
or U18029 (N_18029,N_10563,N_9259);
nor U18030 (N_18030,N_7662,N_9503);
nand U18031 (N_18031,N_8468,N_11038);
and U18032 (N_18032,N_7071,N_8503);
and U18033 (N_18033,N_12143,N_10192);
nor U18034 (N_18034,N_7507,N_8030);
xor U18035 (N_18035,N_8973,N_11833);
or U18036 (N_18036,N_10316,N_7808);
nor U18037 (N_18037,N_7876,N_10674);
and U18038 (N_18038,N_7823,N_11726);
nand U18039 (N_18039,N_7544,N_7339);
nor U18040 (N_18040,N_11223,N_6504);
xor U18041 (N_18041,N_12431,N_12496);
nor U18042 (N_18042,N_8159,N_8227);
nor U18043 (N_18043,N_8515,N_10407);
or U18044 (N_18044,N_11810,N_11702);
or U18045 (N_18045,N_12317,N_9667);
xor U18046 (N_18046,N_10102,N_6929);
or U18047 (N_18047,N_11039,N_11333);
nor U18048 (N_18048,N_6912,N_12282);
xor U18049 (N_18049,N_8007,N_7985);
xor U18050 (N_18050,N_7007,N_9578);
xnor U18051 (N_18051,N_9625,N_10945);
or U18052 (N_18052,N_7769,N_8017);
and U18053 (N_18053,N_6572,N_7113);
nor U18054 (N_18054,N_9703,N_10028);
nand U18055 (N_18055,N_9696,N_10305);
nand U18056 (N_18056,N_11546,N_10364);
nand U18057 (N_18057,N_10105,N_10094);
nor U18058 (N_18058,N_12429,N_9567);
or U18059 (N_18059,N_11111,N_7545);
and U18060 (N_18060,N_10164,N_8778);
nand U18061 (N_18061,N_9336,N_6971);
nor U18062 (N_18062,N_9477,N_8503);
nand U18063 (N_18063,N_7165,N_9321);
nand U18064 (N_18064,N_10441,N_11606);
xnor U18065 (N_18065,N_11964,N_9516);
or U18066 (N_18066,N_11592,N_8341);
or U18067 (N_18067,N_9807,N_12236);
or U18068 (N_18068,N_11179,N_7014);
nand U18069 (N_18069,N_8187,N_11893);
and U18070 (N_18070,N_8254,N_9972);
and U18071 (N_18071,N_7616,N_11296);
and U18072 (N_18072,N_6604,N_7031);
nor U18073 (N_18073,N_8236,N_7921);
or U18074 (N_18074,N_11059,N_7636);
nand U18075 (N_18075,N_9103,N_9643);
or U18076 (N_18076,N_11130,N_6741);
or U18077 (N_18077,N_10567,N_6941);
nand U18078 (N_18078,N_11721,N_11960);
nand U18079 (N_18079,N_7453,N_7402);
nor U18080 (N_18080,N_11725,N_10508);
or U18081 (N_18081,N_6637,N_8093);
and U18082 (N_18082,N_8633,N_6322);
and U18083 (N_18083,N_9607,N_9619);
or U18084 (N_18084,N_9300,N_8311);
or U18085 (N_18085,N_11748,N_7123);
and U18086 (N_18086,N_7856,N_9722);
xnor U18087 (N_18087,N_9934,N_7068);
and U18088 (N_18088,N_9086,N_11185);
xor U18089 (N_18089,N_6677,N_10161);
nand U18090 (N_18090,N_8398,N_10484);
or U18091 (N_18091,N_9204,N_12407);
and U18092 (N_18092,N_10393,N_8790);
nand U18093 (N_18093,N_8172,N_10190);
nor U18094 (N_18094,N_7787,N_11405);
xnor U18095 (N_18095,N_9456,N_8497);
xor U18096 (N_18096,N_7315,N_9856);
or U18097 (N_18097,N_6633,N_8372);
nand U18098 (N_18098,N_11695,N_7791);
or U18099 (N_18099,N_12156,N_8262);
and U18100 (N_18100,N_10680,N_10538);
nand U18101 (N_18101,N_6516,N_9209);
xnor U18102 (N_18102,N_12383,N_12060);
xor U18103 (N_18103,N_9826,N_7404);
or U18104 (N_18104,N_9522,N_7181);
nand U18105 (N_18105,N_11223,N_7510);
xnor U18106 (N_18106,N_8356,N_6879);
nor U18107 (N_18107,N_12214,N_7395);
nor U18108 (N_18108,N_6801,N_10058);
xor U18109 (N_18109,N_7446,N_10549);
nand U18110 (N_18110,N_9848,N_9778);
nand U18111 (N_18111,N_11275,N_10311);
nor U18112 (N_18112,N_7113,N_9536);
nand U18113 (N_18113,N_6582,N_11893);
nand U18114 (N_18114,N_10115,N_10276);
nand U18115 (N_18115,N_8152,N_11767);
nor U18116 (N_18116,N_6692,N_7549);
and U18117 (N_18117,N_7220,N_9881);
nand U18118 (N_18118,N_6349,N_6556);
xor U18119 (N_18119,N_8306,N_8194);
nand U18120 (N_18120,N_11051,N_9925);
nor U18121 (N_18121,N_7509,N_11194);
nand U18122 (N_18122,N_8898,N_6603);
or U18123 (N_18123,N_7587,N_6988);
nand U18124 (N_18124,N_8667,N_8348);
nor U18125 (N_18125,N_8945,N_8837);
and U18126 (N_18126,N_8744,N_8459);
and U18127 (N_18127,N_8389,N_7320);
and U18128 (N_18128,N_9350,N_9137);
and U18129 (N_18129,N_12470,N_10611);
nand U18130 (N_18130,N_8014,N_11795);
or U18131 (N_18131,N_8099,N_12006);
nor U18132 (N_18132,N_8271,N_7570);
and U18133 (N_18133,N_11095,N_8896);
nand U18134 (N_18134,N_6980,N_7460);
xnor U18135 (N_18135,N_10239,N_8658);
nand U18136 (N_18136,N_8465,N_8601);
or U18137 (N_18137,N_12490,N_8505);
or U18138 (N_18138,N_10066,N_8650);
nand U18139 (N_18139,N_6666,N_9466);
nor U18140 (N_18140,N_7544,N_12138);
or U18141 (N_18141,N_11280,N_10278);
or U18142 (N_18142,N_6453,N_9360);
nor U18143 (N_18143,N_11428,N_8136);
or U18144 (N_18144,N_11738,N_6982);
and U18145 (N_18145,N_8949,N_10810);
or U18146 (N_18146,N_7265,N_6690);
nand U18147 (N_18147,N_12052,N_8855);
xnor U18148 (N_18148,N_8153,N_10197);
nand U18149 (N_18149,N_9416,N_10981);
or U18150 (N_18150,N_11078,N_10611);
nand U18151 (N_18151,N_7704,N_11997);
nand U18152 (N_18152,N_7933,N_9298);
nor U18153 (N_18153,N_11434,N_9848);
nand U18154 (N_18154,N_7416,N_12115);
and U18155 (N_18155,N_6414,N_6618);
xor U18156 (N_18156,N_10141,N_8524);
nor U18157 (N_18157,N_9275,N_12315);
nand U18158 (N_18158,N_12070,N_9176);
xnor U18159 (N_18159,N_6478,N_11593);
xnor U18160 (N_18160,N_6435,N_10425);
xor U18161 (N_18161,N_8237,N_12048);
or U18162 (N_18162,N_12133,N_9580);
and U18163 (N_18163,N_8982,N_11346);
and U18164 (N_18164,N_7008,N_8044);
nor U18165 (N_18165,N_7920,N_11493);
nand U18166 (N_18166,N_8342,N_6276);
or U18167 (N_18167,N_8399,N_7115);
or U18168 (N_18168,N_6710,N_6897);
nand U18169 (N_18169,N_6916,N_9000);
nand U18170 (N_18170,N_10692,N_6666);
nor U18171 (N_18171,N_9469,N_10981);
nand U18172 (N_18172,N_8134,N_10408);
or U18173 (N_18173,N_6691,N_9110);
and U18174 (N_18174,N_8641,N_8721);
nand U18175 (N_18175,N_11470,N_6900);
nand U18176 (N_18176,N_7308,N_9513);
or U18177 (N_18177,N_8371,N_12443);
or U18178 (N_18178,N_6937,N_12409);
or U18179 (N_18179,N_9163,N_10519);
xor U18180 (N_18180,N_11164,N_7032);
or U18181 (N_18181,N_7740,N_11632);
xor U18182 (N_18182,N_11248,N_6432);
nand U18183 (N_18183,N_6380,N_11427);
xnor U18184 (N_18184,N_10654,N_7121);
nor U18185 (N_18185,N_11445,N_9814);
and U18186 (N_18186,N_11358,N_11013);
and U18187 (N_18187,N_11538,N_11282);
and U18188 (N_18188,N_11916,N_8686);
nor U18189 (N_18189,N_11676,N_9764);
and U18190 (N_18190,N_12244,N_7481);
or U18191 (N_18191,N_7917,N_12064);
nand U18192 (N_18192,N_9031,N_8612);
nand U18193 (N_18193,N_7434,N_6337);
and U18194 (N_18194,N_6748,N_7769);
xor U18195 (N_18195,N_7954,N_8841);
nand U18196 (N_18196,N_7198,N_10908);
or U18197 (N_18197,N_6473,N_9967);
nand U18198 (N_18198,N_11955,N_7592);
nand U18199 (N_18199,N_6268,N_6526);
nand U18200 (N_18200,N_10108,N_9079);
and U18201 (N_18201,N_6434,N_9975);
nand U18202 (N_18202,N_9018,N_11116);
nor U18203 (N_18203,N_7607,N_10024);
and U18204 (N_18204,N_11403,N_7771);
nor U18205 (N_18205,N_9918,N_8543);
xnor U18206 (N_18206,N_9088,N_12216);
nand U18207 (N_18207,N_8447,N_10609);
and U18208 (N_18208,N_7782,N_9059);
or U18209 (N_18209,N_8649,N_6452);
and U18210 (N_18210,N_6436,N_11464);
or U18211 (N_18211,N_7726,N_10912);
or U18212 (N_18212,N_6359,N_7339);
or U18213 (N_18213,N_8352,N_10864);
and U18214 (N_18214,N_7183,N_9224);
and U18215 (N_18215,N_8527,N_12435);
and U18216 (N_18216,N_6448,N_10068);
xor U18217 (N_18217,N_12142,N_6884);
xor U18218 (N_18218,N_12005,N_12470);
nor U18219 (N_18219,N_7360,N_12043);
xnor U18220 (N_18220,N_11687,N_9913);
nor U18221 (N_18221,N_8303,N_9932);
nor U18222 (N_18222,N_10750,N_9735);
xor U18223 (N_18223,N_10100,N_6693);
or U18224 (N_18224,N_6985,N_8936);
nand U18225 (N_18225,N_10416,N_11157);
or U18226 (N_18226,N_10167,N_7246);
and U18227 (N_18227,N_6398,N_7618);
nor U18228 (N_18228,N_6585,N_6884);
and U18229 (N_18229,N_8628,N_6368);
nand U18230 (N_18230,N_8499,N_6691);
xor U18231 (N_18231,N_7259,N_10273);
nor U18232 (N_18232,N_10185,N_7731);
and U18233 (N_18233,N_8712,N_12167);
nand U18234 (N_18234,N_6766,N_12348);
xnor U18235 (N_18235,N_9202,N_10470);
xor U18236 (N_18236,N_8773,N_12083);
xnor U18237 (N_18237,N_11492,N_11121);
nor U18238 (N_18238,N_7112,N_11595);
and U18239 (N_18239,N_6697,N_7368);
xnor U18240 (N_18240,N_9121,N_9387);
nor U18241 (N_18241,N_7335,N_9425);
nor U18242 (N_18242,N_8451,N_12377);
or U18243 (N_18243,N_6527,N_8548);
xor U18244 (N_18244,N_6743,N_11332);
nand U18245 (N_18245,N_7723,N_9224);
xor U18246 (N_18246,N_12397,N_10455);
and U18247 (N_18247,N_7251,N_10992);
xnor U18248 (N_18248,N_6578,N_11369);
xnor U18249 (N_18249,N_10230,N_11416);
or U18250 (N_18250,N_9312,N_11338);
or U18251 (N_18251,N_10508,N_7803);
nor U18252 (N_18252,N_8051,N_11673);
xor U18253 (N_18253,N_9129,N_10115);
nor U18254 (N_18254,N_11216,N_8355);
xor U18255 (N_18255,N_8012,N_9387);
nand U18256 (N_18256,N_9623,N_6718);
nand U18257 (N_18257,N_10895,N_8613);
and U18258 (N_18258,N_7803,N_11028);
and U18259 (N_18259,N_8808,N_8532);
xor U18260 (N_18260,N_7940,N_9466);
xnor U18261 (N_18261,N_8991,N_10301);
nand U18262 (N_18262,N_9109,N_6976);
and U18263 (N_18263,N_10995,N_10379);
and U18264 (N_18264,N_11224,N_11956);
nor U18265 (N_18265,N_10027,N_10504);
or U18266 (N_18266,N_10023,N_7499);
nor U18267 (N_18267,N_9822,N_10789);
nand U18268 (N_18268,N_10080,N_6989);
nor U18269 (N_18269,N_10960,N_7569);
nand U18270 (N_18270,N_9786,N_9389);
nor U18271 (N_18271,N_9863,N_12233);
or U18272 (N_18272,N_9152,N_11216);
and U18273 (N_18273,N_12415,N_7038);
nand U18274 (N_18274,N_9778,N_11873);
nor U18275 (N_18275,N_6563,N_11561);
nand U18276 (N_18276,N_7377,N_11763);
nor U18277 (N_18277,N_7416,N_7171);
xnor U18278 (N_18278,N_6939,N_12009);
nand U18279 (N_18279,N_11168,N_7627);
nand U18280 (N_18280,N_8797,N_10642);
or U18281 (N_18281,N_9195,N_8371);
nand U18282 (N_18282,N_8647,N_7720);
nor U18283 (N_18283,N_7471,N_10113);
nand U18284 (N_18284,N_11225,N_8519);
xnor U18285 (N_18285,N_9074,N_12305);
xor U18286 (N_18286,N_7192,N_12367);
nand U18287 (N_18287,N_9662,N_7540);
or U18288 (N_18288,N_6839,N_12435);
and U18289 (N_18289,N_6899,N_6758);
and U18290 (N_18290,N_9051,N_11097);
or U18291 (N_18291,N_10859,N_9088);
xnor U18292 (N_18292,N_7858,N_7375);
and U18293 (N_18293,N_6588,N_7887);
nand U18294 (N_18294,N_8983,N_11741);
and U18295 (N_18295,N_8165,N_11327);
nor U18296 (N_18296,N_10716,N_6605);
nor U18297 (N_18297,N_7508,N_11040);
or U18298 (N_18298,N_7001,N_7352);
or U18299 (N_18299,N_10515,N_12089);
nand U18300 (N_18300,N_8815,N_12336);
and U18301 (N_18301,N_8267,N_8848);
nand U18302 (N_18302,N_6593,N_7927);
or U18303 (N_18303,N_7691,N_11190);
xor U18304 (N_18304,N_11686,N_6902);
nor U18305 (N_18305,N_9679,N_7366);
nand U18306 (N_18306,N_8641,N_9930);
and U18307 (N_18307,N_7865,N_10476);
xnor U18308 (N_18308,N_6782,N_8845);
nor U18309 (N_18309,N_9526,N_11202);
xnor U18310 (N_18310,N_8626,N_8970);
nand U18311 (N_18311,N_7493,N_11161);
or U18312 (N_18312,N_10813,N_10797);
or U18313 (N_18313,N_10184,N_8314);
xnor U18314 (N_18314,N_10540,N_7192);
xor U18315 (N_18315,N_6859,N_6680);
or U18316 (N_18316,N_9724,N_10909);
and U18317 (N_18317,N_12193,N_9958);
nand U18318 (N_18318,N_8269,N_10231);
nor U18319 (N_18319,N_6982,N_11596);
nor U18320 (N_18320,N_9859,N_11214);
and U18321 (N_18321,N_8802,N_7087);
xnor U18322 (N_18322,N_9527,N_9951);
nor U18323 (N_18323,N_8670,N_9955);
nor U18324 (N_18324,N_6820,N_7595);
xnor U18325 (N_18325,N_10132,N_8012);
xnor U18326 (N_18326,N_8567,N_9502);
nor U18327 (N_18327,N_10104,N_9934);
and U18328 (N_18328,N_10624,N_8736);
xor U18329 (N_18329,N_9382,N_10511);
and U18330 (N_18330,N_8546,N_6823);
and U18331 (N_18331,N_11297,N_6574);
and U18332 (N_18332,N_9829,N_7756);
and U18333 (N_18333,N_11570,N_11447);
xor U18334 (N_18334,N_7945,N_7796);
or U18335 (N_18335,N_8356,N_8975);
nor U18336 (N_18336,N_7260,N_12064);
and U18337 (N_18337,N_11791,N_11634);
nand U18338 (N_18338,N_12315,N_8562);
nand U18339 (N_18339,N_11692,N_6861);
and U18340 (N_18340,N_7804,N_7696);
or U18341 (N_18341,N_6683,N_10201);
and U18342 (N_18342,N_12207,N_12478);
and U18343 (N_18343,N_10861,N_11161);
nor U18344 (N_18344,N_10810,N_6304);
xnor U18345 (N_18345,N_6591,N_9956);
xnor U18346 (N_18346,N_9292,N_12383);
or U18347 (N_18347,N_10590,N_8321);
nand U18348 (N_18348,N_8413,N_8769);
nor U18349 (N_18349,N_7842,N_7675);
nor U18350 (N_18350,N_8542,N_9203);
or U18351 (N_18351,N_9244,N_11499);
and U18352 (N_18352,N_10452,N_9394);
nor U18353 (N_18353,N_6560,N_9442);
nor U18354 (N_18354,N_9022,N_9421);
xor U18355 (N_18355,N_9888,N_8503);
or U18356 (N_18356,N_9518,N_9059);
xor U18357 (N_18357,N_9256,N_8029);
and U18358 (N_18358,N_11134,N_9234);
nand U18359 (N_18359,N_10684,N_8229);
nor U18360 (N_18360,N_11115,N_10925);
nand U18361 (N_18361,N_9936,N_10233);
nand U18362 (N_18362,N_9893,N_8991);
nor U18363 (N_18363,N_12191,N_10731);
nand U18364 (N_18364,N_11124,N_11618);
or U18365 (N_18365,N_9421,N_8886);
nand U18366 (N_18366,N_11279,N_7303);
and U18367 (N_18367,N_7457,N_6520);
xor U18368 (N_18368,N_8217,N_7979);
nand U18369 (N_18369,N_7009,N_8636);
nand U18370 (N_18370,N_11578,N_6670);
xnor U18371 (N_18371,N_6562,N_11420);
nand U18372 (N_18372,N_10651,N_7083);
nand U18373 (N_18373,N_10971,N_11343);
nand U18374 (N_18374,N_11551,N_9862);
or U18375 (N_18375,N_12169,N_11705);
and U18376 (N_18376,N_7110,N_8136);
nand U18377 (N_18377,N_9545,N_11961);
and U18378 (N_18378,N_10048,N_6385);
nor U18379 (N_18379,N_9725,N_7685);
and U18380 (N_18380,N_7845,N_7820);
or U18381 (N_18381,N_12496,N_12347);
nand U18382 (N_18382,N_7155,N_8655);
or U18383 (N_18383,N_6688,N_7472);
nand U18384 (N_18384,N_11623,N_6805);
or U18385 (N_18385,N_8306,N_6360);
nor U18386 (N_18386,N_11604,N_8482);
or U18387 (N_18387,N_11401,N_10178);
and U18388 (N_18388,N_10551,N_11004);
nand U18389 (N_18389,N_10364,N_11362);
nor U18390 (N_18390,N_8685,N_7547);
xnor U18391 (N_18391,N_8395,N_11307);
nor U18392 (N_18392,N_10436,N_10547);
and U18393 (N_18393,N_12345,N_10347);
or U18394 (N_18394,N_6572,N_7302);
and U18395 (N_18395,N_6541,N_11887);
nor U18396 (N_18396,N_7305,N_8727);
nand U18397 (N_18397,N_11856,N_10583);
and U18398 (N_18398,N_9298,N_11388);
xor U18399 (N_18399,N_8184,N_6551);
or U18400 (N_18400,N_7585,N_9323);
nand U18401 (N_18401,N_8216,N_9369);
and U18402 (N_18402,N_7899,N_7261);
xnor U18403 (N_18403,N_7476,N_9558);
nand U18404 (N_18404,N_11390,N_10281);
and U18405 (N_18405,N_7025,N_7927);
and U18406 (N_18406,N_6454,N_11349);
and U18407 (N_18407,N_11591,N_6501);
nand U18408 (N_18408,N_8976,N_11078);
or U18409 (N_18409,N_8212,N_8311);
xnor U18410 (N_18410,N_11204,N_6608);
or U18411 (N_18411,N_10594,N_11433);
xor U18412 (N_18412,N_6641,N_11714);
and U18413 (N_18413,N_9073,N_11344);
nor U18414 (N_18414,N_8387,N_8166);
nand U18415 (N_18415,N_12292,N_10880);
xnor U18416 (N_18416,N_8440,N_11742);
or U18417 (N_18417,N_10732,N_7935);
or U18418 (N_18418,N_6684,N_7155);
nand U18419 (N_18419,N_10567,N_11643);
nor U18420 (N_18420,N_9493,N_9028);
nand U18421 (N_18421,N_7364,N_11510);
xnor U18422 (N_18422,N_6647,N_11785);
xnor U18423 (N_18423,N_8548,N_7901);
and U18424 (N_18424,N_8171,N_7672);
xnor U18425 (N_18425,N_11854,N_8638);
nand U18426 (N_18426,N_6589,N_7812);
or U18427 (N_18427,N_8124,N_12146);
or U18428 (N_18428,N_10875,N_11634);
xor U18429 (N_18429,N_12381,N_11989);
or U18430 (N_18430,N_12289,N_11608);
or U18431 (N_18431,N_9860,N_10917);
or U18432 (N_18432,N_7630,N_11024);
nor U18433 (N_18433,N_11006,N_7489);
nor U18434 (N_18434,N_11571,N_7829);
and U18435 (N_18435,N_9049,N_7825);
nor U18436 (N_18436,N_9914,N_12013);
and U18437 (N_18437,N_6428,N_8847);
nand U18438 (N_18438,N_11430,N_6498);
or U18439 (N_18439,N_6522,N_11178);
nor U18440 (N_18440,N_10143,N_6320);
or U18441 (N_18441,N_6977,N_7568);
or U18442 (N_18442,N_11672,N_7804);
xor U18443 (N_18443,N_9113,N_11333);
xnor U18444 (N_18444,N_9022,N_10642);
or U18445 (N_18445,N_9427,N_7791);
nor U18446 (N_18446,N_7046,N_7120);
and U18447 (N_18447,N_10311,N_11926);
xnor U18448 (N_18448,N_8397,N_7882);
or U18449 (N_18449,N_7879,N_7691);
and U18450 (N_18450,N_9829,N_7358);
nor U18451 (N_18451,N_8137,N_8163);
nand U18452 (N_18452,N_11910,N_9522);
nand U18453 (N_18453,N_12189,N_7481);
and U18454 (N_18454,N_9693,N_9350);
xnor U18455 (N_18455,N_9235,N_10116);
and U18456 (N_18456,N_8464,N_6305);
or U18457 (N_18457,N_11998,N_11820);
and U18458 (N_18458,N_8398,N_6892);
and U18459 (N_18459,N_6759,N_7466);
and U18460 (N_18460,N_7195,N_8204);
xor U18461 (N_18461,N_9716,N_10984);
xnor U18462 (N_18462,N_9518,N_12377);
or U18463 (N_18463,N_6944,N_8650);
and U18464 (N_18464,N_11306,N_8039);
xnor U18465 (N_18465,N_7963,N_9935);
nor U18466 (N_18466,N_10695,N_6335);
nand U18467 (N_18467,N_12277,N_8955);
xor U18468 (N_18468,N_12017,N_10895);
nor U18469 (N_18469,N_8677,N_6337);
xor U18470 (N_18470,N_12319,N_8672);
and U18471 (N_18471,N_12092,N_8707);
or U18472 (N_18472,N_10392,N_11468);
xnor U18473 (N_18473,N_12388,N_10877);
nand U18474 (N_18474,N_11914,N_9155);
xor U18475 (N_18475,N_10334,N_6446);
or U18476 (N_18476,N_7902,N_7579);
nor U18477 (N_18477,N_8194,N_10466);
nand U18478 (N_18478,N_11703,N_8952);
xor U18479 (N_18479,N_9206,N_12190);
and U18480 (N_18480,N_8749,N_11133);
nor U18481 (N_18481,N_6549,N_7937);
xor U18482 (N_18482,N_9366,N_10811);
xnor U18483 (N_18483,N_7085,N_10259);
and U18484 (N_18484,N_7816,N_10838);
xnor U18485 (N_18485,N_7823,N_9330);
nand U18486 (N_18486,N_9196,N_7879);
and U18487 (N_18487,N_7141,N_11665);
nand U18488 (N_18488,N_9023,N_12336);
nor U18489 (N_18489,N_6486,N_6916);
xnor U18490 (N_18490,N_12296,N_10236);
and U18491 (N_18491,N_8380,N_7608);
nor U18492 (N_18492,N_8420,N_11354);
xor U18493 (N_18493,N_8589,N_9133);
or U18494 (N_18494,N_10935,N_8606);
nor U18495 (N_18495,N_9917,N_8162);
and U18496 (N_18496,N_7473,N_7266);
nand U18497 (N_18497,N_9708,N_11912);
and U18498 (N_18498,N_11257,N_9947);
or U18499 (N_18499,N_11366,N_11910);
or U18500 (N_18500,N_7446,N_9707);
or U18501 (N_18501,N_9375,N_11878);
xor U18502 (N_18502,N_12374,N_6395);
and U18503 (N_18503,N_12391,N_12027);
xor U18504 (N_18504,N_7036,N_7182);
and U18505 (N_18505,N_6924,N_9985);
or U18506 (N_18506,N_7094,N_6780);
nor U18507 (N_18507,N_7062,N_7995);
xnor U18508 (N_18508,N_8393,N_9147);
and U18509 (N_18509,N_10211,N_8253);
and U18510 (N_18510,N_12448,N_6806);
and U18511 (N_18511,N_9397,N_11044);
xnor U18512 (N_18512,N_9400,N_12410);
nand U18513 (N_18513,N_9931,N_6747);
nand U18514 (N_18514,N_11796,N_7455);
xnor U18515 (N_18515,N_11133,N_12454);
or U18516 (N_18516,N_7293,N_6345);
and U18517 (N_18517,N_6372,N_9595);
or U18518 (N_18518,N_7978,N_9211);
nand U18519 (N_18519,N_9421,N_7951);
or U18520 (N_18520,N_11193,N_10403);
nand U18521 (N_18521,N_6783,N_7193);
xor U18522 (N_18522,N_10941,N_8070);
xnor U18523 (N_18523,N_8117,N_10150);
nand U18524 (N_18524,N_7408,N_9078);
xnor U18525 (N_18525,N_8506,N_10077);
nor U18526 (N_18526,N_6870,N_9024);
or U18527 (N_18527,N_12115,N_9236);
nand U18528 (N_18528,N_7015,N_12323);
nor U18529 (N_18529,N_9383,N_10690);
nand U18530 (N_18530,N_6554,N_8005);
and U18531 (N_18531,N_11662,N_6720);
nand U18532 (N_18532,N_11270,N_9944);
or U18533 (N_18533,N_7823,N_7221);
nand U18534 (N_18534,N_9281,N_7964);
or U18535 (N_18535,N_6550,N_7015);
or U18536 (N_18536,N_10933,N_7193);
and U18537 (N_18537,N_11451,N_10560);
nand U18538 (N_18538,N_10591,N_7332);
nand U18539 (N_18539,N_6775,N_7897);
or U18540 (N_18540,N_8996,N_9979);
nor U18541 (N_18541,N_10463,N_9990);
xnor U18542 (N_18542,N_10246,N_11728);
nand U18543 (N_18543,N_11843,N_11994);
or U18544 (N_18544,N_8370,N_11872);
nand U18545 (N_18545,N_8991,N_12157);
nor U18546 (N_18546,N_8232,N_7975);
or U18547 (N_18547,N_11760,N_11721);
and U18548 (N_18548,N_7118,N_8750);
xor U18549 (N_18549,N_10191,N_10909);
and U18550 (N_18550,N_12266,N_10958);
or U18551 (N_18551,N_6421,N_7246);
nor U18552 (N_18552,N_8091,N_11192);
nor U18553 (N_18553,N_10644,N_12186);
and U18554 (N_18554,N_9229,N_6646);
and U18555 (N_18555,N_11620,N_6496);
nor U18556 (N_18556,N_6817,N_7222);
nor U18557 (N_18557,N_7369,N_8213);
xnor U18558 (N_18558,N_10062,N_9811);
xnor U18559 (N_18559,N_10574,N_11764);
and U18560 (N_18560,N_8334,N_11580);
nor U18561 (N_18561,N_10104,N_7876);
nor U18562 (N_18562,N_7350,N_9144);
nand U18563 (N_18563,N_10058,N_12201);
or U18564 (N_18564,N_7655,N_11711);
and U18565 (N_18565,N_9994,N_10579);
xor U18566 (N_18566,N_10405,N_6286);
nand U18567 (N_18567,N_10711,N_9447);
nand U18568 (N_18568,N_9263,N_7808);
and U18569 (N_18569,N_7910,N_10040);
and U18570 (N_18570,N_6723,N_8986);
nor U18571 (N_18571,N_10672,N_8535);
and U18572 (N_18572,N_8041,N_9449);
or U18573 (N_18573,N_8301,N_10466);
and U18574 (N_18574,N_10490,N_9183);
xnor U18575 (N_18575,N_8351,N_6584);
or U18576 (N_18576,N_11972,N_7622);
nand U18577 (N_18577,N_7499,N_7254);
nor U18578 (N_18578,N_11631,N_10950);
and U18579 (N_18579,N_11971,N_10774);
nor U18580 (N_18580,N_9848,N_11556);
nand U18581 (N_18581,N_8835,N_6659);
nor U18582 (N_18582,N_11191,N_7763);
nand U18583 (N_18583,N_10491,N_9425);
or U18584 (N_18584,N_9459,N_6336);
or U18585 (N_18585,N_6943,N_8875);
and U18586 (N_18586,N_8939,N_8698);
and U18587 (N_18587,N_8054,N_9688);
or U18588 (N_18588,N_9781,N_7998);
nor U18589 (N_18589,N_6714,N_7665);
nand U18590 (N_18590,N_8101,N_12091);
xor U18591 (N_18591,N_11733,N_7725);
nor U18592 (N_18592,N_11276,N_10081);
nor U18593 (N_18593,N_9811,N_10557);
nand U18594 (N_18594,N_9921,N_11654);
nor U18595 (N_18595,N_8732,N_10241);
nand U18596 (N_18596,N_8686,N_7629);
and U18597 (N_18597,N_11496,N_8192);
or U18598 (N_18598,N_7001,N_10102);
nor U18599 (N_18599,N_8729,N_10519);
nand U18600 (N_18600,N_9935,N_6972);
nor U18601 (N_18601,N_7880,N_6410);
xor U18602 (N_18602,N_7451,N_9452);
nor U18603 (N_18603,N_9702,N_9679);
xor U18604 (N_18604,N_9096,N_6696);
nand U18605 (N_18605,N_6654,N_8104);
or U18606 (N_18606,N_6606,N_6429);
nand U18607 (N_18607,N_8720,N_10684);
xor U18608 (N_18608,N_9815,N_7238);
and U18609 (N_18609,N_7951,N_10269);
nor U18610 (N_18610,N_8507,N_7396);
and U18611 (N_18611,N_8563,N_8372);
or U18612 (N_18612,N_11653,N_8673);
xnor U18613 (N_18613,N_10522,N_7749);
xnor U18614 (N_18614,N_7796,N_9486);
or U18615 (N_18615,N_9534,N_10491);
nor U18616 (N_18616,N_12357,N_10477);
xnor U18617 (N_18617,N_11244,N_6487);
xor U18618 (N_18618,N_11253,N_8450);
and U18619 (N_18619,N_10773,N_6429);
xnor U18620 (N_18620,N_6366,N_10491);
nand U18621 (N_18621,N_10544,N_9917);
or U18622 (N_18622,N_8475,N_8533);
nor U18623 (N_18623,N_11845,N_11080);
and U18624 (N_18624,N_7945,N_6446);
xnor U18625 (N_18625,N_9555,N_11280);
nand U18626 (N_18626,N_6267,N_7293);
or U18627 (N_18627,N_10311,N_11848);
and U18628 (N_18628,N_12351,N_8029);
or U18629 (N_18629,N_10295,N_11257);
xnor U18630 (N_18630,N_11726,N_7426);
nor U18631 (N_18631,N_11597,N_10684);
xnor U18632 (N_18632,N_11261,N_7700);
nor U18633 (N_18633,N_11719,N_6341);
and U18634 (N_18634,N_7689,N_6260);
and U18635 (N_18635,N_6769,N_6312);
nor U18636 (N_18636,N_7299,N_12286);
nand U18637 (N_18637,N_12291,N_11172);
nand U18638 (N_18638,N_6483,N_11108);
xnor U18639 (N_18639,N_8514,N_11538);
and U18640 (N_18640,N_7748,N_9703);
nor U18641 (N_18641,N_10177,N_12103);
and U18642 (N_18642,N_8684,N_11967);
xnor U18643 (N_18643,N_11981,N_8110);
nor U18644 (N_18644,N_11379,N_11830);
nand U18645 (N_18645,N_10614,N_11188);
and U18646 (N_18646,N_7562,N_11132);
nor U18647 (N_18647,N_8575,N_9309);
and U18648 (N_18648,N_7511,N_10336);
and U18649 (N_18649,N_7577,N_8659);
nor U18650 (N_18650,N_8047,N_8227);
nor U18651 (N_18651,N_10477,N_9731);
nor U18652 (N_18652,N_9826,N_10665);
and U18653 (N_18653,N_10733,N_10063);
or U18654 (N_18654,N_7309,N_10022);
and U18655 (N_18655,N_6659,N_6874);
nor U18656 (N_18656,N_8973,N_11903);
and U18657 (N_18657,N_10164,N_11344);
xnor U18658 (N_18658,N_12262,N_12384);
xnor U18659 (N_18659,N_7222,N_10856);
or U18660 (N_18660,N_9208,N_7685);
nor U18661 (N_18661,N_6360,N_10526);
nand U18662 (N_18662,N_8829,N_8399);
nor U18663 (N_18663,N_10887,N_8935);
xnor U18664 (N_18664,N_6655,N_9646);
nand U18665 (N_18665,N_10412,N_11654);
or U18666 (N_18666,N_7837,N_8771);
xnor U18667 (N_18667,N_11607,N_6694);
nand U18668 (N_18668,N_11335,N_6309);
nor U18669 (N_18669,N_9031,N_8957);
or U18670 (N_18670,N_10803,N_6733);
nor U18671 (N_18671,N_7198,N_12231);
nand U18672 (N_18672,N_11238,N_7225);
or U18673 (N_18673,N_7649,N_10563);
and U18674 (N_18674,N_9678,N_12050);
xnor U18675 (N_18675,N_7963,N_6531);
xor U18676 (N_18676,N_8252,N_7725);
and U18677 (N_18677,N_11108,N_7657);
xor U18678 (N_18678,N_8906,N_8278);
nor U18679 (N_18679,N_11797,N_10339);
or U18680 (N_18680,N_7316,N_9646);
and U18681 (N_18681,N_8013,N_12134);
nand U18682 (N_18682,N_8416,N_10212);
nand U18683 (N_18683,N_12055,N_8891);
nor U18684 (N_18684,N_6336,N_9409);
nor U18685 (N_18685,N_7153,N_7516);
nand U18686 (N_18686,N_8005,N_7857);
nor U18687 (N_18687,N_9067,N_10206);
or U18688 (N_18688,N_8500,N_9557);
nand U18689 (N_18689,N_11966,N_9360);
nor U18690 (N_18690,N_10706,N_9230);
nand U18691 (N_18691,N_8147,N_9418);
nor U18692 (N_18692,N_9024,N_10131);
xnor U18693 (N_18693,N_7935,N_11302);
or U18694 (N_18694,N_9145,N_12324);
nor U18695 (N_18695,N_10991,N_11149);
and U18696 (N_18696,N_9382,N_9070);
nor U18697 (N_18697,N_12173,N_11710);
or U18698 (N_18698,N_9243,N_11301);
and U18699 (N_18699,N_11961,N_10334);
nand U18700 (N_18700,N_8671,N_11127);
nand U18701 (N_18701,N_11362,N_10698);
or U18702 (N_18702,N_6764,N_6732);
xor U18703 (N_18703,N_9528,N_8053);
or U18704 (N_18704,N_12374,N_12334);
nand U18705 (N_18705,N_6882,N_10652);
nor U18706 (N_18706,N_10721,N_7624);
nand U18707 (N_18707,N_12348,N_11009);
xnor U18708 (N_18708,N_7866,N_11221);
nand U18709 (N_18709,N_12056,N_7191);
xor U18710 (N_18710,N_11703,N_6544);
or U18711 (N_18711,N_9723,N_9712);
xor U18712 (N_18712,N_8301,N_9919);
or U18713 (N_18713,N_10024,N_11381);
nor U18714 (N_18714,N_7321,N_9508);
nand U18715 (N_18715,N_7241,N_7591);
or U18716 (N_18716,N_12273,N_7730);
nand U18717 (N_18717,N_8574,N_11274);
xor U18718 (N_18718,N_7280,N_6796);
nand U18719 (N_18719,N_9845,N_11915);
nand U18720 (N_18720,N_8288,N_11910);
nand U18721 (N_18721,N_8314,N_8240);
nand U18722 (N_18722,N_9559,N_7549);
or U18723 (N_18723,N_8296,N_12480);
or U18724 (N_18724,N_11750,N_7265);
xor U18725 (N_18725,N_11803,N_7920);
nand U18726 (N_18726,N_10377,N_7718);
nor U18727 (N_18727,N_9437,N_7474);
or U18728 (N_18728,N_10621,N_10170);
xnor U18729 (N_18729,N_11497,N_7061);
or U18730 (N_18730,N_7622,N_10382);
and U18731 (N_18731,N_7689,N_11314);
and U18732 (N_18732,N_11937,N_12496);
or U18733 (N_18733,N_6346,N_8673);
or U18734 (N_18734,N_8401,N_7183);
nor U18735 (N_18735,N_12363,N_8268);
nand U18736 (N_18736,N_7461,N_12422);
nor U18737 (N_18737,N_10459,N_10151);
nor U18738 (N_18738,N_11923,N_9621);
nor U18739 (N_18739,N_9070,N_9879);
xnor U18740 (N_18740,N_10081,N_7778);
and U18741 (N_18741,N_6259,N_10199);
xor U18742 (N_18742,N_11254,N_6925);
xor U18743 (N_18743,N_8518,N_11839);
nor U18744 (N_18744,N_10420,N_12326);
xor U18745 (N_18745,N_10376,N_12269);
and U18746 (N_18746,N_7709,N_11252);
and U18747 (N_18747,N_11961,N_8609);
nand U18748 (N_18748,N_6922,N_10777);
xor U18749 (N_18749,N_11870,N_11263);
nand U18750 (N_18750,N_15336,N_17085);
nand U18751 (N_18751,N_14034,N_18678);
nand U18752 (N_18752,N_17486,N_15202);
and U18753 (N_18753,N_15881,N_13468);
or U18754 (N_18754,N_15543,N_12727);
xnor U18755 (N_18755,N_16650,N_15081);
or U18756 (N_18756,N_17441,N_18398);
xor U18757 (N_18757,N_15355,N_15784);
nor U18758 (N_18758,N_13181,N_18008);
and U18759 (N_18759,N_18556,N_14172);
and U18760 (N_18760,N_17054,N_15311);
xnor U18761 (N_18761,N_16319,N_12986);
nand U18762 (N_18762,N_13019,N_17417);
nand U18763 (N_18763,N_18512,N_17806);
xor U18764 (N_18764,N_14335,N_15587);
or U18765 (N_18765,N_13269,N_18221);
and U18766 (N_18766,N_12684,N_12681);
nand U18767 (N_18767,N_14892,N_16617);
and U18768 (N_18768,N_16059,N_18716);
xnor U18769 (N_18769,N_14858,N_16189);
nand U18770 (N_18770,N_13910,N_12651);
nand U18771 (N_18771,N_13616,N_12639);
or U18772 (N_18772,N_13568,N_18536);
nand U18773 (N_18773,N_13835,N_13258);
or U18774 (N_18774,N_17566,N_16000);
nand U18775 (N_18775,N_13675,N_17206);
nand U18776 (N_18776,N_13272,N_17135);
or U18777 (N_18777,N_14065,N_17672);
nand U18778 (N_18778,N_12742,N_18466);
or U18779 (N_18779,N_15124,N_13230);
and U18780 (N_18780,N_15140,N_13368);
or U18781 (N_18781,N_17525,N_17710);
or U18782 (N_18782,N_14743,N_17181);
nand U18783 (N_18783,N_17632,N_13165);
xor U18784 (N_18784,N_17276,N_15668);
nand U18785 (N_18785,N_17930,N_15420);
nor U18786 (N_18786,N_13866,N_16768);
nor U18787 (N_18787,N_16583,N_15327);
and U18788 (N_18788,N_17805,N_16634);
nor U18789 (N_18789,N_17794,N_16034);
and U18790 (N_18790,N_16866,N_17067);
nor U18791 (N_18791,N_16279,N_16602);
xor U18792 (N_18792,N_14063,N_15074);
nand U18793 (N_18793,N_17011,N_17184);
xor U18794 (N_18794,N_13475,N_18063);
or U18795 (N_18795,N_16798,N_14136);
or U18796 (N_18796,N_15883,N_15952);
and U18797 (N_18797,N_14804,N_17694);
xor U18798 (N_18798,N_18577,N_17327);
xnor U18799 (N_18799,N_16401,N_13097);
nor U18800 (N_18800,N_15949,N_16804);
nor U18801 (N_18801,N_16425,N_16789);
or U18802 (N_18802,N_17369,N_13704);
and U18803 (N_18803,N_15623,N_14579);
and U18804 (N_18804,N_18484,N_15706);
and U18805 (N_18805,N_15615,N_12700);
nor U18806 (N_18806,N_13608,N_15203);
or U18807 (N_18807,N_16349,N_17836);
xnor U18808 (N_18808,N_15301,N_14538);
nor U18809 (N_18809,N_17675,N_18724);
nand U18810 (N_18810,N_17972,N_14951);
or U18811 (N_18811,N_14346,N_15445);
nand U18812 (N_18812,N_15839,N_12653);
nor U18813 (N_18813,N_14975,N_16536);
or U18814 (N_18814,N_15964,N_16491);
nor U18815 (N_18815,N_16744,N_16779);
nor U18816 (N_18816,N_17698,N_15474);
or U18817 (N_18817,N_15571,N_14401);
nand U18818 (N_18818,N_14875,N_16274);
or U18819 (N_18819,N_16109,N_18596);
or U18820 (N_18820,N_18696,N_16226);
xnor U18821 (N_18821,N_17303,N_17594);
xor U18822 (N_18822,N_13023,N_17692);
and U18823 (N_18823,N_13476,N_13423);
nor U18824 (N_18824,N_15902,N_16040);
xnor U18825 (N_18825,N_12718,N_14803);
and U18826 (N_18826,N_18178,N_14744);
or U18827 (N_18827,N_17969,N_15528);
xnor U18828 (N_18828,N_13664,N_17822);
nand U18829 (N_18829,N_15376,N_14314);
or U18830 (N_18830,N_14705,N_17765);
and U18831 (N_18831,N_18080,N_13595);
or U18832 (N_18832,N_17134,N_14684);
nor U18833 (N_18833,N_18099,N_16480);
or U18834 (N_18834,N_16568,N_15953);
nand U18835 (N_18835,N_16266,N_13005);
or U18836 (N_18836,N_17111,N_14873);
xnor U18837 (N_18837,N_18426,N_15064);
nor U18838 (N_18838,N_16570,N_15872);
nor U18839 (N_18839,N_16654,N_16879);
nor U18840 (N_18840,N_17921,N_13526);
nand U18841 (N_18841,N_16982,N_15484);
and U18842 (N_18842,N_13759,N_15741);
and U18843 (N_18843,N_15493,N_17670);
xor U18844 (N_18844,N_13401,N_15800);
nor U18845 (N_18845,N_12779,N_13129);
nand U18846 (N_18846,N_14174,N_13139);
nor U18847 (N_18847,N_17693,N_15052);
nand U18848 (N_18848,N_17306,N_14503);
xor U18849 (N_18849,N_14917,N_17496);
xnor U18850 (N_18850,N_15996,N_16312);
and U18851 (N_18851,N_13126,N_15359);
nand U18852 (N_18852,N_15709,N_17947);
xor U18853 (N_18853,N_14874,N_13565);
nand U18854 (N_18854,N_12781,N_16803);
nor U18855 (N_18855,N_13967,N_15895);
nor U18856 (N_18856,N_16557,N_17776);
and U18857 (N_18857,N_17401,N_15176);
xor U18858 (N_18858,N_14637,N_18509);
nor U18859 (N_18859,N_14599,N_14453);
nand U18860 (N_18860,N_14590,N_13862);
xnor U18861 (N_18861,N_13582,N_13335);
or U18862 (N_18862,N_15166,N_17989);
xor U18863 (N_18863,N_18697,N_15280);
xnor U18864 (N_18864,N_16464,N_12909);
xnor U18865 (N_18865,N_13603,N_14671);
nand U18866 (N_18866,N_17816,N_14945);
or U18867 (N_18867,N_12949,N_14282);
nand U18868 (N_18868,N_18390,N_16008);
xnor U18869 (N_18869,N_15849,N_17215);
nand U18870 (N_18870,N_15796,N_16805);
or U18871 (N_18871,N_18587,N_14964);
nand U18872 (N_18872,N_16797,N_15229);
or U18873 (N_18873,N_15554,N_15038);
nand U18874 (N_18874,N_15220,N_14850);
nor U18875 (N_18875,N_17863,N_16415);
nand U18876 (N_18876,N_15450,N_12510);
nor U18877 (N_18877,N_17664,N_15133);
xnor U18878 (N_18878,N_15760,N_14116);
and U18879 (N_18879,N_17137,N_13796);
nor U18880 (N_18880,N_16827,N_18247);
xnor U18881 (N_18881,N_16696,N_16533);
or U18882 (N_18882,N_12674,N_17430);
and U18883 (N_18883,N_16261,N_13597);
nor U18884 (N_18884,N_13617,N_16966);
and U18885 (N_18885,N_17962,N_13605);
nand U18886 (N_18886,N_15876,N_15620);
nor U18887 (N_18887,N_15009,N_15068);
nand U18888 (N_18888,N_16784,N_13869);
nor U18889 (N_18889,N_16537,N_18342);
xor U18890 (N_18890,N_17841,N_15778);
or U18891 (N_18891,N_14275,N_15442);
nand U18892 (N_18892,N_16143,N_15986);
nand U18893 (N_18893,N_15717,N_14552);
nand U18894 (N_18894,N_17032,N_15066);
or U18895 (N_18895,N_16441,N_14851);
and U18896 (N_18896,N_15152,N_17346);
nand U18897 (N_18897,N_13307,N_12736);
nand U18898 (N_18898,N_16010,N_17696);
or U18899 (N_18899,N_13699,N_14774);
nor U18900 (N_18900,N_13052,N_16127);
xnor U18901 (N_18901,N_15008,N_14754);
nor U18902 (N_18902,N_16577,N_17047);
or U18903 (N_18903,N_18481,N_18331);
nor U18904 (N_18904,N_13764,N_12878);
and U18905 (N_18905,N_18538,N_12694);
or U18906 (N_18906,N_16947,N_13263);
nor U18907 (N_18907,N_14623,N_18067);
or U18908 (N_18908,N_15243,N_16519);
nor U18909 (N_18909,N_13594,N_17033);
xor U18910 (N_18910,N_15728,N_17616);
or U18911 (N_18911,N_14058,N_14467);
xnor U18912 (N_18912,N_17803,N_17120);
nor U18913 (N_18913,N_14094,N_13960);
and U18914 (N_18914,N_14510,N_17012);
nand U18915 (N_18915,N_12905,N_16198);
xor U18916 (N_18916,N_18313,N_14361);
nand U18917 (N_18917,N_14595,N_16291);
nand U18918 (N_18918,N_15866,N_15691);
and U18919 (N_18919,N_15901,N_13725);
xnor U18920 (N_18920,N_17813,N_17349);
nor U18921 (N_18921,N_13669,N_15974);
and U18922 (N_18922,N_14281,N_18039);
nor U18923 (N_18923,N_12876,N_12806);
or U18924 (N_18924,N_17270,N_13486);
and U18925 (N_18925,N_15303,N_16373);
or U18926 (N_18926,N_14061,N_13969);
or U18927 (N_18927,N_16306,N_18213);
xor U18928 (N_18928,N_14500,N_17884);
or U18929 (N_18929,N_17622,N_16163);
nor U18930 (N_18930,N_15832,N_14998);
xnor U18931 (N_18931,N_15286,N_17044);
nor U18932 (N_18932,N_18365,N_13337);
nand U18933 (N_18933,N_17384,N_14870);
or U18934 (N_18934,N_15987,N_17371);
or U18935 (N_18935,N_13239,N_17015);
xnor U18936 (N_18936,N_12853,N_17125);
nor U18937 (N_18937,N_15762,N_18263);
and U18938 (N_18938,N_13948,N_15016);
xnor U18939 (N_18939,N_13225,N_18656);
nor U18940 (N_18940,N_13120,N_16815);
nand U18941 (N_18941,N_17634,N_13389);
and U18942 (N_18942,N_18260,N_13000);
nand U18943 (N_18943,N_15221,N_18098);
xor U18944 (N_18944,N_17018,N_13149);
and U18945 (N_18945,N_17296,N_18399);
and U18946 (N_18946,N_18586,N_17518);
xor U18947 (N_18947,N_15393,N_13155);
xnor U18948 (N_18948,N_17530,N_17598);
and U18949 (N_18949,N_12537,N_17416);
or U18950 (N_18950,N_16099,N_12545);
or U18951 (N_18951,N_16594,N_18400);
and U18952 (N_18952,N_17847,N_15062);
or U18953 (N_18953,N_18726,N_17472);
nand U18954 (N_18954,N_17022,N_15567);
and U18955 (N_18955,N_13112,N_14425);
nand U18956 (N_18956,N_18069,N_12560);
nand U18957 (N_18957,N_15156,N_16332);
xnor U18958 (N_18958,N_16292,N_14939);
xnor U18959 (N_18959,N_14539,N_12749);
nand U18960 (N_18960,N_18524,N_14620);
nor U18961 (N_18961,N_14665,N_17885);
nand U18962 (N_18962,N_16812,N_16077);
and U18963 (N_18963,N_17244,N_16014);
xnor U18964 (N_18964,N_18446,N_13164);
and U18965 (N_18965,N_15300,N_18442);
or U18966 (N_18966,N_13163,N_18579);
and U18967 (N_18967,N_15590,N_18294);
and U18968 (N_18968,N_15642,N_15975);
and U18969 (N_18969,N_18224,N_16210);
or U18970 (N_18970,N_18269,N_13183);
and U18971 (N_18971,N_15997,N_18430);
nand U18972 (N_18972,N_16727,N_16453);
xnor U18973 (N_18973,N_18107,N_15310);
xnor U18974 (N_18974,N_18148,N_16635);
or U18975 (N_18975,N_13937,N_18428);
xor U18976 (N_18976,N_17383,N_16755);
or U18977 (N_18977,N_18545,N_15033);
xor U18978 (N_18978,N_12837,N_13657);
nor U18979 (N_18979,N_18103,N_18440);
and U18980 (N_18980,N_17479,N_14662);
or U18981 (N_18981,N_15099,N_16223);
and U18982 (N_18982,N_13557,N_13364);
xnor U18983 (N_18983,N_12557,N_13050);
or U18984 (N_18984,N_13553,N_13416);
or U18985 (N_18985,N_13325,N_14435);
xnor U18986 (N_18986,N_14542,N_12675);
or U18987 (N_18987,N_15856,N_13276);
xor U18988 (N_18988,N_17643,N_15580);
xor U18989 (N_18989,N_16501,N_18258);
nand U18990 (N_18990,N_18163,N_13362);
and U18991 (N_18991,N_18278,N_14965);
nand U18992 (N_18992,N_15805,N_15906);
nand U18993 (N_18993,N_17328,N_16228);
or U18994 (N_18994,N_17907,N_17539);
nor U18995 (N_18995,N_18102,N_17565);
and U18996 (N_18996,N_17176,N_17820);
xor U18997 (N_18997,N_16184,N_16985);
nand U18998 (N_18998,N_16120,N_12609);
or U18999 (N_18999,N_13824,N_15870);
and U19000 (N_19000,N_14265,N_18443);
and U19001 (N_19001,N_14656,N_13914);
nor U19002 (N_19002,N_16217,N_17128);
xnor U19003 (N_19003,N_16710,N_17136);
nand U19004 (N_19004,N_14155,N_18233);
nor U19005 (N_19005,N_14634,N_17993);
and U19006 (N_19006,N_18308,N_16183);
nand U19007 (N_19007,N_14956,N_16336);
xor U19008 (N_19008,N_17285,N_18353);
or U19009 (N_19009,N_14481,N_13624);
nor U19010 (N_19010,N_13190,N_16680);
nor U19011 (N_19011,N_18515,N_16857);
nand U19012 (N_19012,N_17658,N_18271);
nand U19013 (N_19013,N_13237,N_16729);
and U19014 (N_19014,N_18460,N_18548);
nor U19015 (N_19015,N_14857,N_13078);
nand U19016 (N_19016,N_18652,N_16036);
xor U19017 (N_19017,N_15905,N_13949);
xnor U19018 (N_19018,N_14115,N_15602);
nand U19019 (N_19019,N_17524,N_13156);
nor U19020 (N_19020,N_15539,N_15114);
and U19021 (N_19021,N_14801,N_12532);
nand U19022 (N_19022,N_13299,N_16020);
nand U19023 (N_19023,N_18675,N_14954);
and U19024 (N_19024,N_15342,N_15605);
xnor U19025 (N_19025,N_14505,N_17919);
xnor U19026 (N_19026,N_15456,N_16687);
nand U19027 (N_19027,N_14379,N_14853);
xor U19028 (N_19028,N_14869,N_14162);
or U19029 (N_19029,N_15181,N_15281);
nor U19030 (N_19030,N_15757,N_14348);
nor U19031 (N_19031,N_15164,N_14356);
or U19032 (N_19032,N_18074,N_17676);
xnor U19033 (N_19033,N_15212,N_12939);
and U19034 (N_19034,N_15931,N_13130);
xor U19035 (N_19035,N_15419,N_17061);
nor U19036 (N_19036,N_13662,N_17075);
nor U19037 (N_19037,N_18002,N_15654);
or U19038 (N_19038,N_14611,N_12811);
or U19039 (N_19039,N_18635,N_17175);
nor U19040 (N_19040,N_18259,N_13460);
nor U19041 (N_19041,N_17282,N_13038);
nor U19042 (N_19042,N_15955,N_15289);
nor U19043 (N_19043,N_15254,N_12892);
xnor U19044 (N_19044,N_18420,N_18431);
or U19045 (N_19045,N_13111,N_14412);
nand U19046 (N_19046,N_14895,N_15088);
or U19047 (N_19047,N_13905,N_15513);
or U19048 (N_19048,N_13278,N_15846);
nor U19049 (N_19049,N_17552,N_14760);
nor U19050 (N_19050,N_17996,N_16979);
or U19051 (N_19051,N_16502,N_15911);
nor U19052 (N_19052,N_14042,N_16413);
and U19053 (N_19053,N_13903,N_15626);
nand U19054 (N_19054,N_13343,N_17365);
nand U19055 (N_19055,N_15806,N_12777);
or U19056 (N_19056,N_18673,N_15667);
and U19057 (N_19057,N_16846,N_16974);
and U19058 (N_19058,N_14617,N_15957);
nor U19059 (N_19059,N_15461,N_16234);
or U19060 (N_19060,N_15148,N_13970);
and U19061 (N_19061,N_18244,N_17414);
xor U19062 (N_19062,N_15680,N_16745);
and U19063 (N_19063,N_13554,N_15071);
xnor U19064 (N_19064,N_13090,N_15437);
xnor U19065 (N_19065,N_13310,N_17666);
nor U19066 (N_19066,N_16939,N_17899);
xnor U19067 (N_19067,N_15833,N_17515);
xor U19068 (N_19068,N_12670,N_13607);
and U19069 (N_19069,N_18312,N_13196);
nand U19070 (N_19070,N_14609,N_14655);
and U19071 (N_19071,N_16747,N_13426);
nand U19072 (N_19072,N_16007,N_16326);
and U19073 (N_19073,N_12914,N_13712);
nor U19074 (N_19074,N_14716,N_13696);
and U19075 (N_19075,N_14902,N_14734);
or U19076 (N_19076,N_13838,N_17191);
and U19077 (N_19077,N_13178,N_14295);
nand U19078 (N_19078,N_18463,N_13891);
nor U19079 (N_19079,N_16558,N_17062);
or U19080 (N_19080,N_15921,N_17888);
nand U19081 (N_19081,N_14122,N_15818);
nand U19082 (N_19082,N_17465,N_14929);
nor U19083 (N_19083,N_15492,N_15803);
and U19084 (N_19084,N_17412,N_15991);
nor U19085 (N_19085,N_17941,N_13593);
and U19086 (N_19086,N_12542,N_12929);
nor U19087 (N_19087,N_16268,N_16022);
nor U19088 (N_19088,N_17976,N_16324);
xor U19089 (N_19089,N_15003,N_15418);
nor U19090 (N_19090,N_16197,N_14022);
and U19091 (N_19091,N_15549,N_14841);
nor U19092 (N_19092,N_17503,N_17968);
xor U19093 (N_19093,N_16694,N_16090);
or U19094 (N_19094,N_16172,N_16520);
or U19095 (N_19095,N_18168,N_17275);
nand U19096 (N_19096,N_18082,N_17977);
and U19097 (N_19097,N_16607,N_18633);
or U19098 (N_19098,N_14690,N_17261);
nor U19099 (N_19099,N_13806,N_14396);
and U19100 (N_19100,N_15126,N_14859);
and U19101 (N_19101,N_16021,N_14785);
nand U19102 (N_19102,N_16298,N_17209);
nand U19103 (N_19103,N_12592,N_17589);
xor U19104 (N_19104,N_17929,N_16205);
nor U19105 (N_19105,N_16448,N_18638);
nand U19106 (N_19106,N_16574,N_16386);
nand U19107 (N_19107,N_15867,N_16418);
nand U19108 (N_19108,N_14879,N_13311);
and U19109 (N_19109,N_18465,N_17326);
xnor U19110 (N_19110,N_16422,N_13134);
or U19111 (N_19111,N_14181,N_14961);
and U19112 (N_19112,N_14541,N_13701);
and U19113 (N_19113,N_13761,N_14818);
and U19114 (N_19114,N_18270,N_15190);
or U19115 (N_19115,N_17232,N_15248);
or U19116 (N_19116,N_17273,N_13930);
and U19117 (N_19117,N_15622,N_14720);
and U19118 (N_19118,N_15705,N_15368);
xor U19119 (N_19119,N_13706,N_18468);
or U19120 (N_19120,N_15296,N_16961);
nor U19121 (N_19121,N_13997,N_12930);
xnor U19122 (N_19122,N_13037,N_15308);
nor U19123 (N_19123,N_12658,N_18193);
xor U19124 (N_19124,N_13204,N_14313);
or U19125 (N_19125,N_15070,N_13691);
or U19126 (N_19126,N_18181,N_18423);
nor U19127 (N_19127,N_12946,N_13140);
and U19128 (N_19128,N_14193,N_17572);
nor U19129 (N_19129,N_15351,N_13405);
nor U19130 (N_19130,N_17127,N_14697);
xor U19131 (N_19131,N_18530,N_12571);
nor U19132 (N_19132,N_14483,N_17886);
nand U19133 (N_19133,N_17093,N_13938);
nand U19134 (N_19134,N_13179,N_16290);
nand U19135 (N_19135,N_18179,N_17671);
xor U19136 (N_19136,N_13655,N_15625);
or U19137 (N_19137,N_16366,N_17213);
and U19138 (N_19138,N_17819,N_15184);
xor U19139 (N_19139,N_17856,N_13184);
xor U19140 (N_19140,N_14000,N_14202);
nand U19141 (N_19141,N_17667,N_14835);
nand U19142 (N_19142,N_15205,N_17043);
xnor U19143 (N_19143,N_18663,N_15488);
nand U19144 (N_19144,N_18644,N_14571);
or U19145 (N_19145,N_16529,N_15729);
and U19146 (N_19146,N_12981,N_16221);
and U19147 (N_19147,N_12872,N_15476);
nand U19148 (N_19148,N_12903,N_14664);
nor U19149 (N_19149,N_18145,N_17810);
nor U19150 (N_19150,N_16071,N_17741);
nor U19151 (N_19151,N_17619,N_18106);
nor U19152 (N_19152,N_16347,N_18089);
xor U19153 (N_19153,N_13927,N_16883);
nand U19154 (N_19154,N_13397,N_17190);
and U19155 (N_19155,N_13981,N_13461);
xor U19156 (N_19156,N_17751,N_15558);
xor U19157 (N_19157,N_16211,N_13398);
nand U19158 (N_19158,N_13544,N_13413);
xor U19159 (N_19159,N_16934,N_15593);
xnor U19160 (N_19160,N_14137,N_12767);
and U19161 (N_19161,N_17866,N_18417);
and U19162 (N_19162,N_17752,N_15962);
or U19163 (N_19163,N_13943,N_14894);
xor U19164 (N_19164,N_12739,N_14343);
and U19165 (N_19165,N_16585,N_15239);
or U19166 (N_19166,N_12954,N_17592);
nand U19167 (N_19167,N_13809,N_16028);
xor U19168 (N_19168,N_15328,N_15610);
nand U19169 (N_19169,N_13068,N_13737);
nor U19170 (N_19170,N_14217,N_13092);
xor U19171 (N_19171,N_13417,N_18433);
or U19172 (N_19172,N_13986,N_17231);
nor U19173 (N_19173,N_13131,N_16517);
and U19174 (N_19174,N_14863,N_16627);
and U19175 (N_19175,N_18214,N_14771);
or U19176 (N_19176,N_17500,N_13495);
and U19177 (N_19177,N_17734,N_13074);
or U19178 (N_19178,N_15211,N_13465);
nor U19179 (N_19179,N_16683,N_12821);
nand U19180 (N_19180,N_16535,N_13373);
or U19181 (N_19181,N_15394,N_13955);
and U19182 (N_19182,N_18262,N_12549);
and U19183 (N_19183,N_12996,N_17571);
or U19184 (N_19184,N_13464,N_18742);
xor U19185 (N_19185,N_18606,N_12548);
nor U19186 (N_19186,N_17736,N_14935);
nor U19187 (N_19187,N_15791,N_13747);
nand U19188 (N_19188,N_17226,N_17889);
xnor U19189 (N_19189,N_15053,N_16204);
and U19190 (N_19190,N_15319,N_15346);
nor U19191 (N_19191,N_13425,N_14557);
or U19192 (N_19192,N_17626,N_17463);
nand U19193 (N_19193,N_14746,N_15963);
or U19194 (N_19194,N_16791,N_16178);
and U19195 (N_19195,N_18209,N_15125);
nand U19196 (N_19196,N_18616,N_14658);
or U19197 (N_19197,N_12788,N_15193);
nor U19198 (N_19198,N_13133,N_16608);
and U19199 (N_19199,N_15891,N_16658);
xor U19200 (N_19200,N_18232,N_16778);
nor U19201 (N_19201,N_12720,N_17459);
xor U19202 (N_19202,N_17713,N_13715);
and U19203 (N_19203,N_18467,N_16229);
nand U19204 (N_19204,N_18542,N_17251);
nor U19205 (N_19205,N_14632,N_18537);
nand U19206 (N_19206,N_17035,N_16575);
nor U19207 (N_19207,N_14100,N_13451);
xnor U19208 (N_19208,N_15491,N_18482);
xor U19209 (N_19209,N_14526,N_14006);
xor U19210 (N_19210,N_15159,N_18283);
nand U19211 (N_19211,N_13570,N_17586);
nor U19212 (N_19212,N_12623,N_13345);
nor U19213 (N_19213,N_17271,N_12772);
xnor U19214 (N_19214,N_17201,N_17991);
nor U19215 (N_19215,N_16712,N_15504);
nand U19216 (N_19216,N_16233,N_13873);
xor U19217 (N_19217,N_12925,N_14201);
and U19218 (N_19218,N_14173,N_17119);
nand U19219 (N_19219,N_15950,N_17733);
and U19220 (N_19220,N_13539,N_15385);
xor U19221 (N_19221,N_15646,N_12959);
xnor U19222 (N_19222,N_17155,N_18202);
nand U19223 (N_19223,N_15083,N_18007);
or U19224 (N_19224,N_16858,N_14214);
xor U19225 (N_19225,N_15002,N_18329);
or U19226 (N_19226,N_13718,N_13705);
xor U19227 (N_19227,N_14001,N_13409);
nand U19228 (N_19228,N_13114,N_13895);
nand U19229 (N_19229,N_16833,N_16783);
or U19230 (N_19230,N_15725,N_15713);
and U19231 (N_19231,N_16988,N_13500);
or U19232 (N_19232,N_16371,N_15501);
or U19233 (N_19233,N_14408,N_14742);
or U19234 (N_19234,N_12689,N_13638);
nor U19235 (N_19235,N_12828,N_16015);
or U19236 (N_19236,N_12762,N_12603);
xnor U19237 (N_19237,N_14333,N_16390);
nand U19238 (N_19238,N_15892,N_17654);
or U19239 (N_19239,N_13846,N_17957);
or U19240 (N_19240,N_16195,N_15751);
nor U19241 (N_19241,N_14197,N_12522);
and U19242 (N_19242,N_17729,N_14825);
xor U19243 (N_19243,N_15928,N_13572);
nor U19244 (N_19244,N_12822,N_15608);
and U19245 (N_19245,N_16452,N_15802);
xnor U19246 (N_19246,N_14271,N_18087);
or U19247 (N_19247,N_18170,N_13851);
nand U19248 (N_19248,N_18318,N_14989);
xor U19249 (N_19249,N_16307,N_18358);
nor U19250 (N_19250,N_16705,N_12595);
nand U19251 (N_19251,N_13330,N_16081);
xor U19252 (N_19252,N_16528,N_17253);
xnor U19253 (N_19253,N_12566,N_12673);
and U19254 (N_19254,N_12933,N_18637);
nand U19255 (N_19255,N_15115,N_16525);
nand U19256 (N_19256,N_16962,N_12540);
and U19257 (N_19257,N_16175,N_14969);
xor U19258 (N_19258,N_13667,N_15799);
nand U19259 (N_19259,N_16892,N_16854);
xor U19260 (N_19260,N_16042,N_13976);
nand U19261 (N_19261,N_13693,N_15173);
nor U19262 (N_19262,N_15031,N_15186);
nor U19263 (N_19263,N_16875,N_13720);
nor U19264 (N_19264,N_18418,N_13372);
and U19265 (N_19265,N_14203,N_15775);
nand U19266 (N_19266,N_18108,N_13222);
and U19267 (N_19267,N_15250,N_14198);
or U19268 (N_19268,N_18101,N_14554);
and U19269 (N_19269,N_13501,N_18169);
and U19270 (N_19270,N_17728,N_16499);
xnor U19271 (N_19271,N_18184,N_16225);
xnor U19272 (N_19272,N_14199,N_18300);
and U19273 (N_19273,N_14899,N_15916);
xnor U19274 (N_19274,N_17984,N_12818);
nand U19275 (N_19275,N_12813,N_18335);
nand U19276 (N_19276,N_14808,N_17187);
nor U19277 (N_19277,N_18020,N_15556);
xnor U19278 (N_19278,N_13562,N_18014);
xor U19279 (N_19279,N_13722,N_12647);
nor U19280 (N_19280,N_18654,N_17050);
nand U19281 (N_19281,N_14779,N_18590);
nand U19282 (N_19282,N_13527,N_16201);
nand U19283 (N_19283,N_17042,N_12652);
nand U19284 (N_19284,N_13220,N_17084);
nor U19285 (N_19285,N_15683,N_16915);
and U19286 (N_19286,N_15297,N_12597);
xnor U19287 (N_19287,N_16257,N_14532);
or U19288 (N_19288,N_15454,N_12646);
nand U19289 (N_19289,N_14428,N_13219);
or U19290 (N_19290,N_18324,N_17827);
nand U19291 (N_19291,N_15413,N_16484);
and U19292 (N_19292,N_16975,N_14334);
nor U19293 (N_19293,N_14589,N_18688);
and U19294 (N_19294,N_17161,N_13378);
or U19295 (N_19295,N_12526,N_16813);
nor U19296 (N_19296,N_14039,N_16145);
and U19297 (N_19297,N_14066,N_17169);
and U19298 (N_19298,N_17737,N_13259);
nor U19299 (N_19299,N_14733,N_17341);
nor U19300 (N_19300,N_15890,N_14406);
nor U19301 (N_19301,N_15153,N_14648);
and U19302 (N_19302,N_13573,N_18029);
nor U19303 (N_19303,N_15377,N_18248);
or U19304 (N_19304,N_14872,N_14472);
nand U19305 (N_19305,N_15795,N_14904);
or U19306 (N_19306,N_18093,N_13041);
or U19307 (N_19307,N_14423,N_16886);
nand U19308 (N_19308,N_17403,N_14140);
xor U19309 (N_19309,N_16514,N_14298);
or U19310 (N_19310,N_16065,N_12640);
and U19311 (N_19311,N_17230,N_17402);
or U19312 (N_19312,N_18473,N_16835);
and U19313 (N_19313,N_14826,N_15993);
nor U19314 (N_19314,N_15732,N_15143);
or U19315 (N_19315,N_15449,N_15027);
nand U19316 (N_19316,N_12780,N_18677);
and U19317 (N_19317,N_15841,N_18710);
nor U19318 (N_19318,N_15287,N_17274);
nor U19319 (N_19319,N_16993,N_14108);
nor U19320 (N_19320,N_14854,N_12773);
and U19321 (N_19321,N_15487,N_15721);
and U19322 (N_19322,N_13889,N_17659);
or U19323 (N_19323,N_13533,N_13916);
xnor U19324 (N_19324,N_16852,N_17638);
nand U19325 (N_19325,N_17971,N_14507);
nand U19326 (N_19326,N_12596,N_18105);
xor U19327 (N_19327,N_15604,N_15384);
and U19328 (N_19328,N_13040,N_18138);
nand U19329 (N_19329,N_14080,N_14441);
or U19330 (N_19330,N_16118,N_18478);
xor U19331 (N_19331,N_13059,N_13540);
nand U19332 (N_19332,N_15292,N_16110);
and U19333 (N_19333,N_14290,N_13233);
nor U19334 (N_19334,N_13989,N_17257);
xor U19335 (N_19335,N_18483,N_17444);
and U19336 (N_19336,N_13576,N_14688);
nor U19337 (N_19337,N_17718,N_15237);
and U19338 (N_19338,N_17716,N_16329);
or U19339 (N_19339,N_13484,N_12722);
xor U19340 (N_19340,N_14008,N_13320);
nand U19341 (N_19341,N_12799,N_13457);
xor U19342 (N_19342,N_16359,N_14365);
or U19343 (N_19343,N_13289,N_15551);
nor U19344 (N_19344,N_13977,N_18200);
and U19345 (N_19345,N_15309,N_13315);
nand U19346 (N_19346,N_18117,N_16018);
or U19347 (N_19347,N_16467,N_17543);
and U19348 (N_19348,N_17440,N_13614);
nor U19349 (N_19349,N_13795,N_12778);
nor U19350 (N_19350,N_14030,N_17464);
and U19351 (N_19351,N_14639,N_13117);
or U19352 (N_19352,N_18362,N_18421);
or U19353 (N_19353,N_17179,N_16530);
nor U19354 (N_19354,N_15511,N_17668);
or U19355 (N_19355,N_16522,N_14641);
nor U19356 (N_19356,N_13399,N_15877);
nand U19357 (N_19357,N_16513,N_16941);
nand U19358 (N_19358,N_15562,N_15396);
or U19359 (N_19359,N_18160,N_13945);
or U19360 (N_19360,N_14479,N_12869);
and U19361 (N_19361,N_15468,N_16543);
nor U19362 (N_19362,N_16439,N_16426);
nor U19363 (N_19363,N_15619,N_12936);
and U19364 (N_19364,N_12601,N_18059);
or U19365 (N_19365,N_15067,N_17106);
xor U19366 (N_19366,N_12656,N_17677);
nand U19367 (N_19367,N_13575,N_18250);
xnor U19368 (N_19368,N_17364,N_15334);
xnor U19369 (N_19369,N_17014,N_15282);
and U19370 (N_19370,N_16898,N_16345);
nand U19371 (N_19371,N_13631,N_17387);
or U19372 (N_19372,N_12719,N_13432);
and U19373 (N_19373,N_15794,N_13096);
and U19374 (N_19374,N_15269,N_16553);
or U19375 (N_19375,N_15616,N_16730);
nor U19376 (N_19376,N_13670,N_17252);
xor U19377 (N_19377,N_17115,N_15995);
and U19378 (N_19378,N_15294,N_13876);
and U19379 (N_19379,N_16656,N_17476);
nor U19380 (N_19380,N_16026,N_14424);
nor U19381 (N_19381,N_14692,N_12637);
and U19382 (N_19382,N_13803,N_14615);
nor U19383 (N_19383,N_15111,N_15464);
nor U19384 (N_19384,N_13636,N_18653);
and U19385 (N_19385,N_15050,N_14591);
xor U19386 (N_19386,N_14167,N_13656);
or U19387 (N_19387,N_13175,N_16052);
nand U19388 (N_19388,N_16300,N_16763);
nor U19389 (N_19389,N_12507,N_17768);
nand U19390 (N_19390,N_12910,N_12812);
nand U19391 (N_19391,N_18018,N_15041);
xnor U19392 (N_19392,N_17487,N_17347);
and U19393 (N_19393,N_15886,N_16896);
and U19394 (N_19394,N_14135,N_15354);
nand U19395 (N_19395,N_13663,N_12561);
nand U19396 (N_19396,N_13113,N_18547);
nor U19397 (N_19397,N_15565,N_17263);
xnor U19398 (N_19398,N_16069,N_12874);
and U19399 (N_19399,N_18648,N_17354);
and U19400 (N_19400,N_17902,N_15787);
or U19401 (N_19401,N_15739,N_16796);
nand U19402 (N_19402,N_16242,N_14031);
and U19403 (N_19403,N_18227,N_17774);
nand U19404 (N_19404,N_16578,N_17547);
nand U19405 (N_19405,N_13494,N_17732);
and U19406 (N_19406,N_15783,N_13328);
xor U19407 (N_19407,N_13979,N_18268);
xor U19408 (N_19408,N_13192,N_16286);
or U19409 (N_19409,N_17436,N_17635);
and U19410 (N_19410,N_15167,N_17532);
nor U19411 (N_19411,N_12591,N_17195);
nand U19412 (N_19412,N_13223,N_15617);
nor U19413 (N_19413,N_14059,N_15715);
nand U19414 (N_19414,N_16393,N_15525);
xor U19415 (N_19415,N_17240,N_17584);
nor U19416 (N_19416,N_14269,N_16709);
nand U19417 (N_19417,N_18304,N_13009);
and U19418 (N_19418,N_13836,N_15929);
or U19419 (N_19419,N_15665,N_15129);
nand U19420 (N_19420,N_13779,N_17662);
and U19421 (N_19421,N_14139,N_16646);
nand U19422 (N_19422,N_18563,N_17194);
nand U19423 (N_19423,N_18264,N_16837);
nor U19424 (N_19424,N_14786,N_14177);
and U19425 (N_19425,N_15888,N_18643);
nand U19426 (N_19426,N_18683,N_14033);
and U19427 (N_19427,N_14947,N_18600);
xnor U19428 (N_19428,N_14653,N_18005);
xor U19429 (N_19429,N_14013,N_14837);
or U19430 (N_19430,N_12569,N_16055);
and U19431 (N_19431,N_16093,N_14682);
or U19432 (N_19432,N_14291,N_14143);
nor U19433 (N_19433,N_17560,N_17953);
nor U19434 (N_19434,N_13290,N_16644);
or U19435 (N_19435,N_17970,N_15636);
nor U19436 (N_19436,N_13881,N_17482);
or U19437 (N_19437,N_12858,N_13317);
xnor U19438 (N_19438,N_14772,N_15370);
xnor U19439 (N_19439,N_16478,N_13602);
xor U19440 (N_19440,N_14967,N_16062);
nand U19441 (N_19441,N_16460,N_13710);
xnor U19442 (N_19442,N_12676,N_14708);
nor U19443 (N_19443,N_13536,N_12894);
and U19444 (N_19444,N_15258,N_16004);
or U19445 (N_19445,N_14053,N_13138);
nand U19446 (N_19446,N_15776,N_15275);
nand U19447 (N_19447,N_13615,N_18237);
or U19448 (N_19448,N_12562,N_14384);
or U19449 (N_19449,N_16482,N_15655);
xnor U19450 (N_19450,N_14805,N_13407);
and U19451 (N_19451,N_16928,N_16068);
or U19452 (N_19452,N_13428,N_13658);
nand U19453 (N_19453,N_18177,N_18747);
nor U19454 (N_19454,N_13404,N_17222);
nor U19455 (N_19455,N_13733,N_16381);
nand U19456 (N_19456,N_13479,N_17460);
nand U19457 (N_19457,N_15631,N_15107);
nor U19458 (N_19458,N_18631,N_15862);
nand U19459 (N_19459,N_16177,N_16037);
nor U19460 (N_19460,N_17633,N_13649);
or U19461 (N_19461,N_12667,N_13797);
nor U19462 (N_19462,N_15197,N_13157);
and U19463 (N_19463,N_16101,N_18743);
or U19464 (N_19464,N_13377,N_15606);
and U19465 (N_19465,N_17721,N_14728);
or U19466 (N_19466,N_14231,N_17604);
xor U19467 (N_19467,N_12789,N_15836);
xnor U19468 (N_19468,N_17027,N_18140);
nor U19469 (N_19469,N_15588,N_16555);
xor U19470 (N_19470,N_13769,N_15781);
nand U19471 (N_19471,N_15288,N_14638);
or U19472 (N_19472,N_14024,N_14062);
or U19473 (N_19473,N_17150,N_14433);
nor U19474 (N_19474,N_17133,N_13295);
nor U19475 (N_19475,N_17236,N_16016);
or U19476 (N_19476,N_12755,N_16096);
nand U19477 (N_19477,N_15711,N_16188);
xnor U19478 (N_19478,N_16450,N_16094);
nor U19479 (N_19479,N_18535,N_15614);
nand U19480 (N_19480,N_12993,N_12608);
or U19481 (N_19481,N_18060,N_16669);
and U19482 (N_19482,N_13169,N_16046);
nor U19483 (N_19483,N_16389,N_18012);
and U19484 (N_19484,N_16668,N_14186);
or U19485 (N_19485,N_14718,N_16149);
nor U19486 (N_19486,N_15720,N_16440);
nand U19487 (N_19487,N_14321,N_16919);
or U19488 (N_19488,N_13122,N_18083);
and U19489 (N_19489,N_12785,N_16997);
xnor U19490 (N_19490,N_17182,N_15235);
nand U19491 (N_19491,N_16604,N_17909);
nor U19492 (N_19492,N_15224,N_16907);
xnor U19493 (N_19493,N_14619,N_14166);
nor U19494 (N_19494,N_17840,N_13736);
and U19495 (N_19495,N_16991,N_15335);
or U19496 (N_19496,N_13287,N_16356);
xnor U19497 (N_19497,N_17510,N_13067);
nand U19498 (N_19498,N_14337,N_14315);
xor U19499 (N_19499,N_18571,N_12867);
nand U19500 (N_19500,N_17999,N_16534);
or U19501 (N_19501,N_16148,N_17623);
nor U19502 (N_19502,N_17089,N_14011);
nor U19503 (N_19503,N_18497,N_13266);
or U19504 (N_19504,N_16321,N_13523);
and U19505 (N_19505,N_16924,N_13261);
or U19506 (N_19506,N_16706,N_18289);
xor U19507 (N_19507,N_16921,N_14159);
nand U19508 (N_19508,N_18561,N_17312);
nor U19509 (N_19509,N_18076,N_12834);
or U19510 (N_19510,N_16508,N_15817);
or U19511 (N_19511,N_15548,N_16157);
and U19512 (N_19512,N_12814,N_18422);
and U19513 (N_19513,N_16639,N_16642);
nand U19514 (N_19514,N_18393,N_17641);
xnor U19515 (N_19515,N_12882,N_14607);
nor U19516 (N_19516,N_16737,N_16855);
or U19517 (N_19517,N_16249,N_15589);
xor U19518 (N_19518,N_18676,N_17467);
and U19519 (N_19519,N_13877,N_16391);
xor U19520 (N_19520,N_16667,N_15049);
nand U19521 (N_19521,N_15970,N_17488);
xor U19522 (N_19522,N_18496,N_14213);
and U19523 (N_19523,N_14920,N_12805);
or U19524 (N_19524,N_13621,N_15196);
nand U19525 (N_19525,N_14876,N_18709);
and U19526 (N_19526,N_12511,N_17117);
nand U19527 (N_19527,N_12715,N_12696);
nor U19528 (N_19528,N_15072,N_12886);
or U19529 (N_19529,N_12911,N_16679);
nand U19530 (N_19530,N_18095,N_13201);
or U19531 (N_19531,N_17558,N_15339);
or U19532 (N_19532,N_17904,N_14621);
xor U19533 (N_19533,N_16414,N_15013);
and U19534 (N_19534,N_18734,N_13434);
and U19535 (N_19535,N_13752,N_17057);
xor U19536 (N_19536,N_15200,N_14577);
xnor U19537 (N_19537,N_17569,N_14341);
and U19538 (N_19538,N_16963,N_13316);
and U19539 (N_19539,N_14886,N_13843);
nor U19540 (N_19540,N_12659,N_17961);
nand U19541 (N_19541,N_17028,N_17162);
nand U19542 (N_19542,N_14468,N_17845);
nor U19543 (N_19543,N_15026,N_15252);
or U19544 (N_19544,N_14432,N_18553);
and U19545 (N_19545,N_18720,N_12683);
and U19546 (N_19546,N_14888,N_12890);
xnor U19547 (N_19547,N_18667,N_18151);
xnor U19548 (N_19548,N_18343,N_18651);
and U19549 (N_19549,N_12567,N_16105);
and U19550 (N_19550,N_13028,N_17485);
and U19551 (N_19551,N_17843,N_14302);
nor U19552 (N_19552,N_17388,N_16636);
nand U19553 (N_19553,N_15462,N_15559);
nand U19554 (N_19554,N_18305,N_18037);
nor U19555 (N_19555,N_13849,N_12915);
and U19556 (N_19556,N_16243,N_16983);
or U19557 (N_19557,N_17483,N_14457);
nor U19558 (N_19558,N_16159,N_18040);
nand U19559 (N_19559,N_12902,N_15966);
and U19560 (N_19560,N_18256,N_13051);
nor U19561 (N_19561,N_17077,N_12840);
or U19562 (N_19562,N_17691,N_13079);
xnor U19563 (N_19563,N_16045,N_16972);
or U19564 (N_19564,N_13784,N_18301);
or U19565 (N_19565,N_18731,N_12956);
nand U19566 (N_19566,N_15880,N_17258);
xnor U19567 (N_19567,N_13395,N_14349);
xnor U19568 (N_19568,N_16492,N_17427);
xnor U19569 (N_19569,N_17259,N_15889);
xor U19570 (N_19570,N_15285,N_18124);
nand U19571 (N_19571,N_15320,N_17657);
or U19572 (N_19572,N_16301,N_17523);
nand U19573 (N_19573,N_16288,N_14832);
and U19574 (N_19574,N_14484,N_12580);
or U19575 (N_19575,N_18403,N_15215);
nand U19576 (N_19576,N_13929,N_17385);
and U19577 (N_19577,N_16897,N_16331);
nand U19578 (N_19578,N_14212,N_13896);
nor U19579 (N_19579,N_18199,N_15875);
nor U19580 (N_19580,N_14587,N_17129);
and U19581 (N_19581,N_18728,N_14695);
or U19582 (N_19582,N_18714,N_18578);
and U19583 (N_19583,N_16573,N_18325);
and U19584 (N_19584,N_18113,N_18255);
or U19585 (N_19585,N_16255,N_14109);
nor U19586 (N_19586,N_15904,N_14943);
xnor U19587 (N_19587,N_15443,N_14908);
nand U19588 (N_19588,N_18584,N_15274);
or U19589 (N_19589,N_17896,N_13581);
nor U19590 (N_19590,N_18155,N_18494);
nor U19591 (N_19591,N_15871,N_15579);
or U19592 (N_19592,N_13980,N_14289);
or U19593 (N_19593,N_14099,N_15132);
nand U19594 (N_19594,N_13679,N_14101);
nor U19595 (N_19595,N_18010,N_16316);
or U19596 (N_19596,N_14487,N_13991);
nor U19597 (N_19597,N_14669,N_16905);
xor U19598 (N_19598,N_16498,N_17105);
nand U19599 (N_19599,N_15325,N_17753);
and U19600 (N_19600,N_15188,N_13104);
xor U19601 (N_19601,N_12550,N_13815);
and U19602 (N_19602,N_18694,N_14081);
or U19603 (N_19603,N_18079,N_18624);
nand U19604 (N_19604,N_15976,N_12871);
nand U19605 (N_19605,N_15772,N_17661);
xnor U19606 (N_19606,N_18238,N_14355);
or U19607 (N_19607,N_15135,N_15688);
or U19608 (N_19608,N_17562,N_17965);
nand U19609 (N_19609,N_15422,N_13818);
and U19610 (N_19610,N_12520,N_16660);
xor U19611 (N_19611,N_13293,N_13303);
and U19612 (N_19612,N_16275,N_16468);
nor U19613 (N_19613,N_18488,N_14654);
xor U19614 (N_19614,N_17269,N_15843);
and U19615 (N_19615,N_15723,N_16125);
and U19616 (N_19616,N_15343,N_13321);
or U19617 (N_19617,N_16352,N_18411);
nor U19618 (N_19618,N_14234,N_13419);
xor U19619 (N_19619,N_13994,N_16592);
xnor U19620 (N_19620,N_14568,N_13642);
xnor U19621 (N_19621,N_16995,N_15932);
and U19622 (N_19622,N_14748,N_14727);
and U19623 (N_19623,N_15681,N_15318);
nand U19624 (N_19624,N_14154,N_16518);
and U19625 (N_19625,N_13653,N_13437);
and U19626 (N_19626,N_14357,N_18050);
and U19627 (N_19627,N_12509,N_15391);
xor U19628 (N_19628,N_15407,N_13076);
nand U19629 (N_19629,N_16075,N_13816);
or U19630 (N_19630,N_14504,N_16131);
nor U19631 (N_19631,N_14210,N_14466);
and U19632 (N_19632,N_16505,N_15352);
xor U19633 (N_19633,N_13538,N_13284);
or U19634 (N_19634,N_16354,N_18604);
nor U19635 (N_19635,N_15500,N_16841);
nand U19636 (N_19636,N_14543,N_12554);
nand U19637 (N_19637,N_17773,N_15119);
or U19638 (N_19638,N_18458,N_14626);
nor U19639 (N_19639,N_17550,N_13498);
nand U19640 (N_19640,N_14674,N_15857);
or U19641 (N_19641,N_12784,N_12976);
nor U19642 (N_19642,N_12707,N_17687);
and U19643 (N_19643,N_13884,N_13243);
and U19644 (N_19644,N_17373,N_17557);
or U19645 (N_19645,N_17239,N_13548);
nand U19646 (N_19646,N_14310,N_14215);
or U19647 (N_19647,N_15922,N_13951);
and U19648 (N_19648,N_14474,N_17262);
nor U19649 (N_19649,N_16054,N_17630);
xnor U19650 (N_19650,N_16212,N_13618);
and U19651 (N_19651,N_14715,N_16545);
and U19652 (N_19652,N_14912,N_18550);
nor U19653 (N_19653,N_16417,N_15388);
or U19654 (N_19654,N_13268,N_14016);
nor U19655 (N_19655,N_17418,N_18306);
and U19656 (N_19656,N_14687,N_13018);
nand U19657 (N_19657,N_15702,N_17339);
or U19658 (N_19658,N_13279,N_15797);
or U19659 (N_19659,N_18081,N_18309);
nor U19660 (N_19660,N_15000,N_16981);
xnor U19661 (N_19661,N_12961,N_15943);
nor U19662 (N_19662,N_16978,N_15724);
nand U19663 (N_19663,N_15727,N_14736);
and U19664 (N_19664,N_17590,N_13150);
and U19665 (N_19665,N_13931,N_15686);
or U19666 (N_19666,N_15271,N_14238);
nand U19667 (N_19667,N_16652,N_15448);
nor U19668 (N_19668,N_18132,N_14925);
and U19669 (N_19669,N_16616,N_18056);
nor U19670 (N_19670,N_14946,N_12972);
nand U19671 (N_19671,N_18733,N_16017);
and U19672 (N_19672,N_15134,N_15304);
and U19673 (N_19673,N_17871,N_13793);
or U19674 (N_19674,N_15767,N_17100);
nand U19675 (N_19675,N_13577,N_13681);
xor U19676 (N_19676,N_12950,N_14362);
and U19677 (N_19677,N_14597,N_14035);
and U19678 (N_19678,N_16563,N_14578);
nand U19679 (N_19679,N_16265,N_14938);
nand U19680 (N_19680,N_17649,N_15295);
nand U19681 (N_19681,N_13734,N_17172);
or U19682 (N_19682,N_12819,N_13411);
nor U19683 (N_19683,N_15860,N_14891);
xor U19684 (N_19684,N_15985,N_13932);
nand U19685 (N_19685,N_16550,N_16030);
and U19686 (N_19686,N_15972,N_17272);
xnor U19687 (N_19687,N_16295,N_12924);
nor U19688 (N_19688,N_16649,N_16431);
nand U19689 (N_19689,N_14195,N_13822);
and U19690 (N_19690,N_18173,N_17682);
nand U19691 (N_19691,N_18321,N_15858);
nor U19692 (N_19692,N_13677,N_15017);
nand U19693 (N_19693,N_14145,N_17314);
xor U19694 (N_19694,N_14262,N_18684);
and U19695 (N_19695,N_16774,N_15045);
xor U19696 (N_19696,N_18690,N_15908);
or U19697 (N_19697,N_13379,N_15734);
nand U19698 (N_19698,N_14111,N_16405);
and U19699 (N_19699,N_16697,N_18216);
or U19700 (N_19700,N_12565,N_18475);
and U19701 (N_19701,N_17697,N_16200);
nand U19702 (N_19702,N_14451,N_18211);
or U19703 (N_19703,N_16049,N_17433);
or U19704 (N_19704,N_15789,N_16847);
nand U19705 (N_19705,N_14559,N_16860);
and U19706 (N_19706,N_15718,N_13620);
xnor U19707 (N_19707,N_16871,N_16877);
xnor U19708 (N_19708,N_15047,N_15232);
or U19709 (N_19709,N_18505,N_12599);
nor U19710 (N_19710,N_17249,N_13212);
xnor U19711 (N_19711,N_13717,N_16466);
and U19712 (N_19712,N_18030,N_16144);
xor U19713 (N_19713,N_17324,N_17048);
nor U19714 (N_19714,N_16830,N_17878);
and U19715 (N_19715,N_17316,N_17005);
nand U19716 (N_19716,N_16591,N_15284);
or U19717 (N_19717,N_18231,N_17798);
xor U19718 (N_19718,N_17469,N_17858);
xnor U19719 (N_19719,N_16598,N_13442);
or U19720 (N_19720,N_13999,N_14354);
nand U19721 (N_19721,N_17448,N_13569);
xor U19722 (N_19722,N_17702,N_13755);
nor U19723 (N_19723,N_15934,N_17955);
nor U19724 (N_19724,N_17374,N_18048);
nor U19725 (N_19725,N_15840,N_14953);
and U19726 (N_19726,N_13363,N_12584);
xor U19727 (N_19727,N_13987,N_13767);
nand U19728 (N_19728,N_13334,N_18583);
nor U19729 (N_19729,N_16902,N_16053);
nand U19730 (N_19730,N_18075,N_14060);
nor U19731 (N_19731,N_15900,N_15138);
or U19732 (N_19732,N_16025,N_14991);
nor U19733 (N_19733,N_18036,N_14009);
and U19734 (N_19734,N_13232,N_17873);
xnor U19735 (N_19735,N_13908,N_13125);
nand U19736 (N_19736,N_15898,N_16958);
and U19737 (N_19737,N_13893,N_15112);
xnor U19738 (N_19738,N_13053,N_16785);
nand U19739 (N_19739,N_18704,N_14865);
or U19740 (N_19740,N_18626,N_13909);
nand U19741 (N_19741,N_13633,N_14107);
nor U19742 (N_19742,N_16361,N_16432);
or U19743 (N_19743,N_16134,N_14125);
nand U19744 (N_19744,N_13302,N_14124);
nor U19745 (N_19745,N_18071,N_15079);
and U19746 (N_19746,N_14319,N_12615);
nor U19747 (N_19747,N_14927,N_18261);
nand U19748 (N_19748,N_14575,N_14286);
nand U19749 (N_19749,N_14582,N_16711);
nand U19750 (N_19750,N_17065,N_12737);
xnor U19751 (N_19751,N_14471,N_13865);
nand U19752 (N_19752,N_18337,N_12868);
xnor U19753 (N_19753,N_15023,N_14521);
or U19754 (N_19754,N_13918,N_14877);
nand U19755 (N_19755,N_12655,N_13323);
nand U19756 (N_19756,N_12973,N_14570);
xnor U19757 (N_19757,N_16495,N_15251);
nand U19758 (N_19758,N_18444,N_13274);
or U19759 (N_19759,N_15242,N_15570);
nor U19760 (N_19760,N_15046,N_15572);
and U19761 (N_19761,N_15032,N_18220);
nand U19762 (N_19762,N_14072,N_14882);
nand U19763 (N_19763,N_12957,N_15238);
and U19764 (N_19764,N_18085,N_14766);
nand U19765 (N_19765,N_16623,N_18402);
nor U19766 (N_19766,N_15494,N_16500);
nor U19767 (N_19767,N_18511,N_17656);
nand U19768 (N_19768,N_14223,N_18738);
xnor U19769 (N_19769,N_13095,N_17588);
nand U19770 (N_19770,N_15749,N_13735);
nor U19771 (N_19771,N_17450,N_15307);
and U19772 (N_19772,N_14816,N_13744);
xor U19773 (N_19773,N_12671,N_16596);
nor U19774 (N_19774,N_14113,N_15428);
nand U19775 (N_19775,N_13771,N_14820);
nor U19776 (N_19776,N_18500,N_17870);
and U19777 (N_19777,N_18543,N_16271);
nand U19778 (N_19778,N_12863,N_16767);
and U19779 (N_19779,N_17410,N_17735);
xor U19780 (N_19780,N_17183,N_18464);
and U19781 (N_19781,N_17828,N_12964);
or U19782 (N_19782,N_13073,N_13109);
xnor U19783 (N_19783,N_14005,N_16690);
nor U19784 (N_19784,N_13791,N_18116);
nand U19785 (N_19785,N_15123,N_16734);
xnor U19786 (N_19786,N_16771,N_12960);
nor U19787 (N_19787,N_12769,N_14911);
nor U19788 (N_19788,N_18042,N_16104);
nor U19789 (N_19789,N_16141,N_14848);
nand U19790 (N_19790,N_14098,N_18719);
nand U19791 (N_19791,N_17304,N_18739);
or U19792 (N_19792,N_15879,N_13341);
nor U19793 (N_19793,N_17744,N_16064);
or U19794 (N_19794,N_12680,N_18485);
or U19795 (N_19795,N_17358,N_18208);
nand U19796 (N_19796,N_14646,N_14627);
or U19797 (N_19797,N_14997,N_13203);
and U19798 (N_19798,N_17527,N_15899);
nor U19799 (N_19799,N_17924,N_14160);
nor U19800 (N_19800,N_17754,N_14704);
or U19801 (N_19801,N_13438,N_18197);
and U19802 (N_19802,N_14003,N_15007);
nor U19803 (N_19803,N_17395,N_12815);
nor U19804 (N_19804,N_17918,N_18722);
and U19805 (N_19805,N_12517,N_16136);
nor U19806 (N_19806,N_16873,N_15096);
or U19807 (N_19807,N_17481,N_18539);
nor U19808 (N_19808,N_14544,N_15137);
xnor U19809 (N_19809,N_14719,N_18705);
nand U19810 (N_19810,N_15988,N_17366);
and U19811 (N_19811,N_14270,N_16350);
nand U19812 (N_19812,N_18134,N_17131);
nand U19813 (N_19813,N_17108,N_16473);
xnor U19814 (N_19814,N_17350,N_12734);
and U19815 (N_19815,N_18424,N_15809);
xor U19816 (N_19816,N_15087,N_16082);
nand U19817 (N_19817,N_15333,N_13485);
nor U19818 (N_19818,N_12793,N_17860);
or U19819 (N_19819,N_18493,N_14631);
nor U19820 (N_19820,N_15831,N_16693);
nand U19821 (N_19821,N_14222,N_13490);
nor U19822 (N_19822,N_14780,N_13242);
or U19823 (N_19823,N_14392,N_17839);
or U19824 (N_19824,N_15677,N_14037);
nand U19825 (N_19825,N_13961,N_15091);
nor U19826 (N_19826,N_12695,N_16908);
nand U19827 (N_19827,N_14067,N_13511);
xnor U19828 (N_19828,N_18414,N_15130);
nand U19829 (N_19829,N_17544,N_12690);
nor U19830 (N_19830,N_18130,N_15874);
nand U19831 (N_19831,N_18275,N_12817);
nor U19832 (N_19832,N_18416,N_13567);
or U19833 (N_19833,N_13629,N_12792);
nand U19834 (N_19834,N_16323,N_13244);
nor U19835 (N_19835,N_14548,N_15581);
and U19836 (N_19836,N_13588,N_17080);
xnor U19837 (N_19837,N_17782,N_16444);
xor U19838 (N_19838,N_14773,N_16056);
nor U19839 (N_19839,N_15937,N_16999);
xor U19840 (N_19840,N_17151,N_13384);
nor U19841 (N_19841,N_12859,N_14434);
nor U19842 (N_19842,N_15144,N_14502);
nand U19843 (N_19843,N_15097,N_15707);
or U19844 (N_19844,N_17112,N_13151);
and U19845 (N_19845,N_13863,N_14488);
nor U19846 (N_19846,N_14192,N_15028);
and U19847 (N_19847,N_13030,N_14885);
or U19848 (N_19848,N_18245,N_17579);
xnor U19849 (N_19849,N_13071,N_16076);
or U19850 (N_19850,N_13333,N_15766);
xor U19851 (N_19851,N_14528,N_16546);
and U19852 (N_19852,N_17156,N_16114);
nor U19853 (N_19853,N_17895,N_14710);
xor U19854 (N_19854,N_16445,N_17540);
and U19855 (N_19855,N_16357,N_14717);
or U19856 (N_19856,N_16926,N_17379);
nor U19857 (N_19857,N_17790,N_15700);
xor U19858 (N_19858,N_12877,N_13015);
nor U19859 (N_19859,N_15569,N_15349);
nor U19860 (N_19860,N_15042,N_18369);
nand U19861 (N_19861,N_13382,N_15664);
or U19862 (N_19862,N_18658,N_13087);
and U19863 (N_19863,N_13499,N_17504);
and U19864 (N_19864,N_18009,N_13390);
nor U19865 (N_19865,N_17321,N_13436);
xor U19866 (N_19866,N_15092,N_15828);
and U19867 (N_19867,N_13648,N_16814);
nor U19868 (N_19868,N_13919,N_13497);
nand U19869 (N_19869,N_17545,N_17703);
or U19870 (N_19870,N_16264,N_16165);
nand U19871 (N_19871,N_13956,N_16129);
nand U19872 (N_19872,N_16160,N_13773);
xor U19873 (N_19873,N_16824,N_17439);
or U19874 (N_19874,N_16302,N_12965);
or U19875 (N_19875,N_17122,N_15145);
and U19876 (N_19876,N_16953,N_17001);
or U19877 (N_19877,N_15495,N_15770);
nor U19878 (N_19878,N_18215,N_16206);
or U19879 (N_19879,N_12638,N_15954);
or U19880 (N_19880,N_13354,N_17409);
nor U19881 (N_19881,N_13213,N_13612);
and U19882 (N_19882,N_17908,N_15613);
nor U19883 (N_19883,N_16438,N_16831);
xnor U19884 (N_19884,N_16749,N_18618);
nand U19885 (N_19885,N_12748,N_16904);
xnor U19886 (N_19886,N_17660,N_12860);
nand U19887 (N_19887,N_18217,N_14218);
and U19888 (N_19888,N_18632,N_14263);
and U19889 (N_19889,N_12791,N_14103);
xor U19890 (N_19890,N_16424,N_17357);
xnor U19891 (N_19891,N_15348,N_16839);
nor U19892 (N_19892,N_14299,N_18028);
nor U19893 (N_19893,N_17023,N_14179);
and U19894 (N_19894,N_16187,N_15813);
nand U19895 (N_19895,N_17597,N_14657);
nand U19896 (N_19896,N_17653,N_14293);
nand U19897 (N_19897,N_17701,N_17477);
nand U19898 (N_19898,N_16829,N_14018);
nand U19899 (N_19899,N_13089,N_15716);
and U19900 (N_19900,N_12870,N_14353);
nor U19901 (N_19901,N_18119,N_18711);
nor U19902 (N_19902,N_14317,N_16477);
or U19903 (N_19903,N_12897,N_17170);
nand U19904 (N_19904,N_17556,N_15273);
nand U19905 (N_19905,N_14800,N_16420);
nand U19906 (N_19906,N_18707,N_17857);
nor U19907 (N_19907,N_17180,N_17652);
nand U19908 (N_19908,N_12705,N_14652);
xnor U19909 (N_19909,N_14232,N_12733);
and U19910 (N_19910,N_15347,N_16430);
xor U19911 (N_19911,N_14164,N_13739);
xnor U19912 (N_19912,N_18354,N_14170);
xnor U19913 (N_19913,N_15515,N_16970);
nand U19914 (N_19914,N_17394,N_15182);
and U19915 (N_19915,N_14327,N_17578);
or U19916 (N_19916,N_14373,N_16185);
and U19917 (N_19917,N_15703,N_16097);
xnor U19918 (N_19918,N_13841,N_12729);
or U19919 (N_19919,N_15661,N_16748);
and U19920 (N_19920,N_16152,N_18610);
or U19921 (N_19921,N_17743,N_18461);
and U19922 (N_19922,N_17797,N_16051);
xnor U19923 (N_19923,N_18686,N_17913);
or U19924 (N_19924,N_13798,N_13760);
xnor U19925 (N_19925,N_12611,N_16579);
or U19926 (N_19926,N_17644,N_18004);
nand U19927 (N_19927,N_16673,N_14546);
or U19928 (N_19928,N_18044,N_16396);
and U19929 (N_19929,N_15537,N_13072);
nor U19930 (N_19930,N_18125,N_16140);
or U19931 (N_19931,N_15216,N_17617);
xor U19932 (N_19932,N_16305,N_12687);
nor U19933 (N_19933,N_14110,N_12521);
nor U19934 (N_19934,N_17173,N_15652);
or U19935 (N_19935,N_16750,N_12502);
xnor U19936 (N_19936,N_17088,N_12636);
xnor U19937 (N_19937,N_17348,N_16214);
xnor U19938 (N_19938,N_13531,N_14836);
or U19939 (N_19939,N_17757,N_14390);
xor U19940 (N_19940,N_12901,N_13246);
and U19941 (N_19941,N_17770,N_13535);
and U19942 (N_19942,N_16173,N_16428);
or U19943 (N_19943,N_15518,N_18376);
or U19944 (N_19944,N_13772,N_13545);
nor U19945 (N_19945,N_16842,N_16406);
nor U19946 (N_19946,N_13762,N_14050);
nor U19947 (N_19947,N_13392,N_13091);
or U19948 (N_19948,N_17037,N_15853);
or U19949 (N_19949,N_17605,N_12829);
and U19950 (N_19950,N_14056,N_16364);
xnor U19951 (N_19951,N_16576,N_17144);
or U19952 (N_19952,N_16773,N_17376);
nand U19953 (N_19953,N_14205,N_18136);
or U19954 (N_19954,N_13584,N_16990);
nand U19955 (N_19955,N_15178,N_15670);
xnor U19956 (N_19956,N_14810,N_18147);
nand U19957 (N_19957,N_16566,N_17449);
or U19958 (N_19958,N_13661,N_13172);
nand U19959 (N_19959,N_16348,N_13634);
or U19960 (N_19960,N_18740,N_15321);
and U19961 (N_19961,N_14134,N_15194);
or U19962 (N_19962,N_13724,N_12995);
nand U19963 (N_19963,N_15748,N_17419);
xor U19964 (N_19964,N_17879,N_14347);
or U19965 (N_19965,N_14278,N_18175);
nor U19966 (N_19966,N_18717,N_16327);
or U19967 (N_19967,N_17553,N_14495);
nor U19968 (N_19968,N_18394,N_14644);
and U19969 (N_19969,N_18328,N_14280);
xnor U19970 (N_19970,N_14118,N_16913);
nand U19971 (N_19971,N_15516,N_14303);
or U19972 (N_19972,N_14900,N_12666);
xnor U19973 (N_19973,N_14279,N_15740);
nor U19974 (N_19974,N_15960,N_12982);
or U19975 (N_19975,N_17452,N_15746);
or U19976 (N_19976,N_15634,N_15367);
or U19977 (N_19977,N_12751,N_14242);
nor U19978 (N_19978,N_14534,N_15256);
and U19979 (N_19979,N_16725,N_14937);
xnor U19980 (N_19980,N_12685,N_14498);
and U19981 (N_19981,N_17071,N_15977);
and U19982 (N_19982,N_17092,N_14229);
nor U19983 (N_19983,N_12501,N_14383);
nor U19984 (N_19984,N_17711,N_16463);
nand U19985 (N_19985,N_13017,N_18302);
or U19986 (N_19986,N_13366,N_14367);
nand U19987 (N_19987,N_14842,N_17665);
xnor U19988 (N_19988,N_16412,N_12971);
or U19989 (N_19989,N_13923,N_12558);
nor U19990 (N_19990,N_16620,N_13852);
nand U19991 (N_19991,N_16825,N_13058);
or U19992 (N_19992,N_15865,N_13635);
nand U19993 (N_19993,N_14224,N_12508);
nor U19994 (N_19994,N_16701,N_17164);
xnor U19995 (N_19995,N_15160,N_18630);
xnor U19996 (N_19996,N_18392,N_18395);
and U19997 (N_19997,N_15743,N_16423);
nor U19998 (N_19998,N_18022,N_17397);
nor U19999 (N_19999,N_14677,N_14913);
nor U20000 (N_20000,N_16612,N_13260);
nor U20001 (N_20001,N_17502,N_16293);
and U20002 (N_20002,N_14806,N_14562);
nand U20003 (N_20003,N_14751,N_13543);
and U20004 (N_20004,N_15118,N_15100);
and U20005 (N_20005,N_12823,N_14064);
nor U20006 (N_20006,N_12746,N_13136);
nand U20007 (N_20007,N_13646,N_13944);
and U20008 (N_20008,N_16776,N_18016);
nand U20009 (N_20009,N_14681,N_15498);
xnor U20010 (N_20010,N_13462,N_15917);
nor U20011 (N_20011,N_14624,N_12943);
or U20012 (N_20012,N_12691,N_18407);
or U20013 (N_20013,N_13571,N_13878);
xor U20014 (N_20014,N_15261,N_13890);
and U20015 (N_20015,N_14491,N_17212);
or U20016 (N_20016,N_12660,N_13195);
xor U20017 (N_20017,N_13057,N_14375);
nor U20018 (N_20018,N_13716,N_15837);
nand U20019 (N_20019,N_13978,N_17719);
or U20020 (N_20020,N_14791,N_18104);
or U20021 (N_20021,N_17621,N_15259);
nor U20022 (N_20022,N_15390,N_15433);
xor U20023 (N_20023,N_17837,N_12538);
xor U20024 (N_20024,N_14090,N_13065);
xnor U20025 (N_20025,N_15507,N_14304);
and U20026 (N_20026,N_14324,N_18361);
or U20027 (N_20027,N_15036,N_17875);
or U20028 (N_20028,N_12763,N_17715);
nor U20029 (N_20029,N_14649,N_13160);
and U20030 (N_20030,N_17587,N_16273);
nand U20031 (N_20031,N_13360,N_17278);
and U20032 (N_20032,N_14211,N_15198);
nand U20033 (N_20033,N_17772,N_12506);
nand U20034 (N_20034,N_13049,N_17850);
or U20035 (N_20035,N_16113,N_15657);
nor U20036 (N_20036,N_16670,N_14014);
or U20037 (N_20037,N_13672,N_12801);
or U20038 (N_20038,N_12841,N_17700);
nand U20039 (N_20039,N_15423,N_13359);
nand U20040 (N_20040,N_17045,N_16544);
and U20041 (N_20041,N_17706,N_14407);
nand U20042 (N_20042,N_17686,N_17583);
and U20043 (N_20043,N_13517,N_15863);
or U20044 (N_20044,N_15765,N_13652);
or U20045 (N_20045,N_14371,N_16098);
or U20046 (N_20046,N_14380,N_14884);
or U20047 (N_20047,N_13361,N_17815);
nor U20048 (N_20048,N_14123,N_15750);
or U20049 (N_20049,N_14048,N_16199);
and U20050 (N_20050,N_16672,N_13340);
xnor U20051 (N_20051,N_17555,N_14287);
and U20052 (N_20052,N_18642,N_13985);
xnor U20053 (N_20053,N_15496,N_15669);
or U20054 (N_20054,N_16083,N_17113);
or U20055 (N_20055,N_16259,N_13673);
nor U20056 (N_20056,N_16746,N_17143);
and U20057 (N_20057,N_17593,N_12541);
nor U20058 (N_20058,N_13146,N_15816);
nand U20059 (N_20059,N_12504,N_18153);
or U20060 (N_20060,N_15489,N_12994);
xor U20061 (N_20061,N_16977,N_15878);
nand U20062 (N_20062,N_17109,N_16954);
and U20063 (N_20063,N_18634,N_18725);
and U20064 (N_20064,N_15199,N_12940);
and U20065 (N_20065,N_17393,N_13783);
or U20066 (N_20066,N_15754,N_13789);
nor U20067 (N_20067,N_16956,N_12551);
or U20068 (N_20068,N_14741,N_16810);
xnor U20069 (N_20069,N_14470,N_15666);
nand U20070 (N_20070,N_13200,N_18477);
nor U20071 (N_20071,N_12699,N_13435);
and U20072 (N_20072,N_17447,N_13683);
and U20073 (N_20073,N_17620,N_13082);
nand U20074 (N_20074,N_17396,N_16942);
nor U20075 (N_20075,N_13444,N_15227);
nand U20076 (N_20076,N_16380,N_15773);
or U20077 (N_20077,N_15774,N_18470);
nor U20078 (N_20078,N_13947,N_17103);
xnor U20079 (N_20079,N_13240,N_14598);
xnor U20080 (N_20080,N_13897,N_15630);
nand U20081 (N_20081,N_17862,N_16378);
or U20082 (N_20082,N_15541,N_14045);
nor U20083 (N_20083,N_17309,N_17830);
or U20084 (N_20084,N_16930,N_13924);
xor U20085 (N_20085,N_17411,N_15699);
or U20086 (N_20086,N_14490,N_16935);
nor U20087 (N_20087,N_12555,N_14770);
or U20088 (N_20088,N_16322,N_13939);
nand U20089 (N_20089,N_16549,N_13729);
xnor U20090 (N_20090,N_13719,N_14344);
or U20091 (N_20091,N_14252,N_17683);
xnor U20092 (N_20092,N_13452,N_14576);
or U20093 (N_20093,N_13750,N_14645);
nand U20094 (N_20094,N_15293,N_16248);
xor U20095 (N_20095,N_17611,N_15014);
xnor U20096 (N_20096,N_15738,N_16276);
xnor U20097 (N_20097,N_17943,N_18026);
xor U20098 (N_20098,N_17891,N_15512);
nand U20099 (N_20099,N_14409,N_18298);
nand U20100 (N_20100,N_13854,N_12693);
nand U20101 (N_20101,N_14284,N_16202);
nand U20102 (N_20102,N_17817,N_12820);
or U20103 (N_20103,N_17920,N_12572);
nand U20104 (N_20104,N_14273,N_13626);
xor U20105 (N_20105,N_15752,N_13306);
nand U20106 (N_20106,N_16459,N_15637);
or U20107 (N_20107,N_16443,N_14560);
or U20108 (N_20108,N_15477,N_13370);
nand U20109 (N_20109,N_18180,N_13487);
nor U20110 (N_20110,N_15956,N_15771);
or U20111 (N_20111,N_13965,N_16597);
or U20112 (N_20112,N_12967,N_17139);
xnor U20113 (N_20113,N_18114,N_18597);
nor U20114 (N_20114,N_15444,N_12802);
and U20115 (N_20115,N_14104,N_18013);
nand U20116 (N_20116,N_13507,N_14387);
nand U20117 (N_20117,N_16493,N_18015);
nor U20118 (N_20118,N_17625,N_16946);
nand U20119 (N_20119,N_16087,N_18374);
nor U20120 (N_20120,N_18451,N_15524);
nand U20121 (N_20121,N_16590,N_16998);
xnor U20122 (N_20122,N_16497,N_15381);
xor U20123 (N_20123,N_15545,N_15730);
xor U20124 (N_20124,N_13001,N_15826);
nor U20125 (N_20125,N_15566,N_16769);
nand U20126 (N_20126,N_18569,N_13647);
nand U20127 (N_20127,N_15369,N_16376);
nor U20128 (N_20128,N_15267,N_17563);
or U20129 (N_20129,N_12816,N_16724);
nor U20130 (N_20130,N_14907,N_15353);
or U20131 (N_20131,N_16759,N_17202);
and U20132 (N_20132,N_16377,N_12630);
nor U20133 (N_20133,N_12856,N_15365);
and U20134 (N_20134,N_14368,N_15466);
nor U20135 (N_20135,N_17462,N_18172);
nand U20136 (N_20136,N_18207,N_12862);
or U20137 (N_20137,N_16446,N_15737);
nor U20138 (N_20138,N_16890,N_18516);
and U20139 (N_20139,N_16384,N_16122);
nand U20140 (N_20140,N_12883,N_17785);
nor U20141 (N_20141,N_18293,N_14316);
and U20142 (N_20142,N_16723,N_13832);
nand U20143 (N_20143,N_14949,N_15555);
or U20144 (N_20144,N_13521,N_16661);
or U20145 (N_20145,N_12570,N_15635);
or U20146 (N_20146,N_17160,N_12898);
xor U20147 (N_20147,N_18368,N_16238);
and U20148 (N_20148,N_13066,N_15792);
xnor U20149 (N_20149,N_15470,N_17742);
nand U20150 (N_20150,N_14699,N_18692);
nand U20151 (N_20151,N_12525,N_18340);
and U20152 (N_20152,N_13286,N_15829);
or U20153 (N_20153,N_15523,N_17574);
or U20154 (N_20154,N_17842,N_18229);
nor U20155 (N_20155,N_16551,N_12750);
or U20156 (N_20156,N_13971,N_13599);
nor U20157 (N_20157,N_14306,N_13660);
and U20158 (N_20158,N_18038,N_14630);
xor U20159 (N_20159,N_17185,N_14485);
nor U20160 (N_20160,N_18174,N_12617);
nor U20161 (N_20161,N_13253,N_15225);
xor U20162 (N_20162,N_16733,N_18568);
nand U20163 (N_20163,N_14696,N_18749);
and U20164 (N_20164,N_15436,N_16713);
nand U20165 (N_20165,N_16314,N_15894);
xnor U20166 (N_20166,N_16304,N_16317);
or U20167 (N_20167,N_15217,N_15624);
or U20168 (N_20168,N_14340,N_14228);
or U20169 (N_20169,N_17725,N_15386);
nand U20170 (N_20170,N_13601,N_13817);
xor U20171 (N_20171,N_13754,N_16628);
and U20172 (N_20172,N_15410,N_18706);
xnor U20173 (N_20173,N_14146,N_18389);
nor U20174 (N_20174,N_18341,N_17833);
and U20175 (N_20175,N_14087,N_17484);
nand U20176 (N_20176,N_14329,N_18666);
xnor U20177 (N_20177,N_16240,N_18330);
and U20178 (N_20178,N_18713,N_16792);
or U20179 (N_20179,N_13530,N_14141);
and U20180 (N_20180,N_14267,N_17740);
nand U20181 (N_20181,N_18188,N_17730);
xnor U20182 (N_20182,N_17499,N_12800);
and U20183 (N_20183,N_15223,N_16887);
and U20184 (N_20184,N_15315,N_13868);
xor U20185 (N_20185,N_15078,N_17096);
xnor U20186 (N_20186,N_17166,N_14443);
nand U20187 (N_20187,N_13802,N_14678);
and U20188 (N_20188,N_15968,N_18650);
and U20189 (N_20189,N_16162,N_14625);
and U20190 (N_20190,N_16078,N_16494);
xnor U20191 (N_20191,N_17600,N_12721);
nor U20192 (N_20192,N_17073,N_15358);
and U20193 (N_20193,N_12602,N_17331);
nand U20194 (N_20194,N_16355,N_17404);
xnor U20195 (N_20195,N_17695,N_17501);
or U20196 (N_20196,N_18602,N_14320);
and U20197 (N_20197,N_17446,N_18551);
xnor U20198 (N_20198,N_14629,N_18546);
and U20199 (N_20199,N_13301,N_13167);
and U20200 (N_20200,N_16676,N_14986);
nor U20201 (N_20201,N_17036,N_18336);
or U20202 (N_20202,N_15910,N_14666);
nand U20203 (N_20203,N_18592,N_13787);
nand U20204 (N_20204,N_15676,N_15844);
or U20205 (N_20205,N_12891,N_14574);
xor U20206 (N_20206,N_17286,N_17315);
nand U20207 (N_20207,N_16923,N_13119);
or U20208 (N_20208,N_18519,N_17648);
and U20209 (N_20209,N_14393,N_12845);
xor U20210 (N_20210,N_17777,N_13972);
nor U20211 (N_20211,N_13912,N_15591);
and U20212 (N_20212,N_15207,N_18055);
nand U20213 (N_20213,N_13294,N_13537);
nor U20214 (N_20214,N_12735,N_13888);
xor U20215 (N_20215,N_15457,N_12528);
nand U20216 (N_20216,N_13680,N_12697);
nor U20217 (N_20217,N_15573,N_15169);
or U20218 (N_20218,N_14709,N_17243);
xnor U20219 (N_20219,N_17575,N_18729);
and U20220 (N_20220,N_16241,N_16541);
xor U20221 (N_20221,N_13555,N_14661);
nand U20222 (N_20222,N_15404,N_15075);
or U20223 (N_20223,N_16945,N_15408);
or U20224 (N_20224,N_15736,N_17567);
nor U20225 (N_20225,N_12513,N_17415);
xor U20226 (N_20226,N_16308,N_16253);
xnor U20227 (N_20227,N_13493,N_18066);
xor U20228 (N_20228,N_12796,N_13936);
and U20229 (N_20229,N_16256,N_14089);
xor U20230 (N_20230,N_15592,N_15467);
or U20231 (N_20231,N_14635,N_13206);
nor U20232 (N_20232,N_12848,N_15149);
nand U20233 (N_20233,N_15204,N_17265);
nor U20234 (N_20234,N_16254,N_14864);
or U20235 (N_20235,N_13928,N_16486);
or U20236 (N_20236,N_13282,N_18534);
or U20237 (N_20237,N_14959,N_14896);
nor U20238 (N_20238,N_15790,N_13700);
nor U20239 (N_20239,N_14897,N_12649);
and U20240 (N_20240,N_16483,N_15305);
or U20241 (N_20241,N_16182,N_12827);
xor U20242 (N_20242,N_12850,N_12614);
nor U20243 (N_20243,N_17915,N_17082);
xor U20244 (N_20244,N_13381,N_16057);
nand U20245 (N_20245,N_14860,N_13424);
and U20246 (N_20246,N_17159,N_14126);
xor U20247 (N_20247,N_14963,N_14017);
and U20248 (N_20248,N_16621,N_18453);
or U20249 (N_20249,N_12587,N_13161);
nand U20250 (N_20250,N_17761,N_15521);
and U20251 (N_20251,N_15316,N_16387);
and U20252 (N_20252,N_12516,N_12999);
and U20253 (N_20253,N_13860,N_13732);
xnor U20254 (N_20254,N_12774,N_15022);
nand U20255 (N_20255,N_15483,N_14622);
nand U20256 (N_20256,N_13099,N_16079);
nor U20257 (N_20257,N_16822,N_14866);
or U20258 (N_20258,N_15201,N_13491);
and U20259 (N_20259,N_14301,N_16899);
nor U20260 (N_20260,N_18235,N_14525);
xnor U20261 (N_20261,N_15662,N_13478);
and U20262 (N_20262,N_16194,N_15663);
or U20263 (N_20263,N_14827,N_16552);
nand U20264 (N_20264,N_14350,N_12923);
and U20265 (N_20265,N_14128,N_15948);
nor U20266 (N_20266,N_15057,N_13197);
xor U20267 (N_20267,N_14797,N_18092);
and U20268 (N_20268,N_17317,N_14338);
nor U20269 (N_20269,N_15918,N_18061);
xor U20270 (N_20270,N_15179,N_14790);
and U20271 (N_20271,N_12563,N_17145);
nand U20272 (N_20272,N_16949,N_13339);
nand U20273 (N_20273,N_16382,N_13470);
xor U20274 (N_20274,N_13996,N_14707);
or U20275 (N_20275,N_17453,N_16764);
nor U20276 (N_20276,N_16952,N_17466);
and U20277 (N_20277,N_17581,N_14241);
nor U20278 (N_20278,N_18474,N_13892);
or U20279 (N_20279,N_16863,N_16313);
and U20280 (N_20280,N_17983,N_13604);
and U20281 (N_20281,N_12628,N_16029);
and U20282 (N_20282,N_17052,N_17494);
or U20283 (N_20283,N_14235,N_14855);
nor U20284 (N_20284,N_16912,N_12836);
nand U20285 (N_20285,N_13135,N_12594);
nand U20286 (N_20286,N_17340,N_14972);
xnor U20287 (N_20287,N_13371,N_15868);
nor U20288 (N_20288,N_16367,N_14292);
or U20289 (N_20289,N_13304,N_15379);
or U20290 (N_20290,N_13820,N_14156);
xor U20291 (N_20291,N_13504,N_13830);
and U20292 (N_20292,N_17072,N_14750);
xor U20293 (N_20293,N_13606,N_17951);
nor U20294 (N_20294,N_13081,N_16788);
nor U20295 (N_20295,N_18452,N_13080);
or U20296 (N_20296,N_17853,N_16220);
or U20297 (N_20297,N_13367,N_17325);
nand U20298 (N_20298,N_12904,N_12770);
and U20299 (N_20299,N_15291,N_15650);
xor U20300 (N_20300,N_17163,N_17076);
xor U20301 (N_20301,N_15180,N_16485);
nand U20302 (N_20302,N_18307,N_17229);
and U20303 (N_20303,N_12605,N_18413);
nor U20304 (N_20304,N_16033,N_13034);
or U20305 (N_20305,N_18527,N_16176);
xor U20306 (N_20306,N_12633,N_17406);
nand U20307 (N_20307,N_16651,N_14508);
or U20308 (N_20308,N_16344,N_18438);
xor U20309 (N_20309,N_14755,N_15279);
nand U20310 (N_20310,N_16509,N_18456);
and U20311 (N_20311,N_14439,N_14386);
or U20312 (N_20312,N_15675,N_12745);
or U20313 (N_20313,N_12703,N_16032);
nand U20314 (N_20314,N_13158,N_14183);
and U20315 (N_20315,N_12849,N_13651);
nand U20316 (N_20316,N_16856,N_14112);
and U20317 (N_20317,N_15561,N_12753);
or U20318 (N_20318,N_15647,N_13098);
or U20319 (N_20319,N_13257,N_13993);
or U20320 (N_20320,N_14405,N_15121);
nand U20321 (N_20321,N_14381,N_15913);
nand U20322 (N_20322,N_17986,N_16442);
nor U20323 (N_20323,N_18234,N_17541);
and U20324 (N_20324,N_16532,N_13645);
and U20325 (N_20325,N_12678,N_15034);
nand U20326 (N_20326,N_14336,N_13926);
nor U20327 (N_20327,N_14933,N_18212);
nand U20328 (N_20328,N_13482,N_14227);
or U20329 (N_20329,N_17960,N_17748);
and U20330 (N_20330,N_12980,N_14691);
nor U20331 (N_20331,N_12621,N_14817);
nor U20332 (N_20332,N_14916,N_14756);
or U20333 (N_20333,N_17775,N_13728);
or U20334 (N_20334,N_13740,N_15745);
nand U20335 (N_20335,N_13094,N_16691);
nand U20336 (N_20336,N_14296,N_16786);
xor U20337 (N_20337,N_13406,N_17305);
nor U20338 (N_20338,N_18154,N_14449);
xnor U20339 (N_20339,N_15850,N_14923);
xnor U20340 (N_20340,N_16353,N_14533);
nor U20341 (N_20341,N_15403,N_18186);
and U20342 (N_20342,N_15927,N_16868);
nor U20343 (N_20343,N_15544,N_18249);
or U20344 (N_20344,N_13344,N_16698);
or U20345 (N_20345,N_14082,N_16244);
or U20346 (N_20346,N_13580,N_13831);
and U20347 (N_20347,N_16252,N_18375);
or U20348 (N_20348,N_18518,N_16472);
nor U20349 (N_20349,N_18062,N_15338);
xor U20350 (N_20350,N_14994,N_18338);
xor U20351 (N_20351,N_17614,N_13520);
and U20352 (N_20352,N_14465,N_13063);
nand U20353 (N_20353,N_17291,N_15434);
nand U20354 (N_20354,N_16128,N_16632);
and U20355 (N_20355,N_17431,N_14807);
xor U20356 (N_20356,N_12552,N_12945);
or U20357 (N_20357,N_14244,N_18540);
and U20358 (N_20358,N_13825,N_14114);
and U20359 (N_20359,N_18146,N_15583);
nor U20360 (N_20360,N_15761,N_16615);
and U20361 (N_20361,N_12842,N_17368);
or U20362 (N_20362,N_18620,N_18355);
xor U20363 (N_20363,N_15415,N_15162);
nand U20364 (N_20364,N_15425,N_14745);
xnor U20365 (N_20365,N_13386,N_14762);
nand U20366 (N_20366,N_15001,N_17663);
or U20367 (N_20367,N_15290,N_18272);
nor U20368 (N_20368,N_17724,N_18469);
nand U20369 (N_20369,N_16840,N_13312);
and U20370 (N_20370,N_12744,N_17284);
nor U20371 (N_20371,N_15157,N_12826);
or U20372 (N_20372,N_14838,N_17391);
nor U20373 (N_20373,N_18744,N_15366);
or U20374 (N_20374,N_15644,N_14867);
or U20375 (N_20375,N_15362,N_13273);
or U20376 (N_20376,N_14735,N_12664);
or U20377 (N_20377,N_18128,N_18531);
nor U20378 (N_20378,N_18296,N_16657);
nand U20379 (N_20379,N_15260,N_14138);
or U20380 (N_20380,N_13264,N_16561);
and U20381 (N_20381,N_16170,N_13280);
or U20382 (N_20382,N_14074,N_18492);
nor U20383 (N_20383,N_17038,N_17268);
xnor U20384 (N_20384,N_13804,N_12920);
xnor U20385 (N_20385,N_15312,N_18541);
xor U20386 (N_20386,N_15719,N_13654);
or U20387 (N_20387,N_16524,N_18619);
xnor U20388 (N_20388,N_13357,N_12970);
nand U20389 (N_20389,N_14073,N_16263);
nor U20390 (N_20390,N_17508,N_15177);
nand U20391 (N_20391,N_16605,N_15510);
nand U20392 (N_20392,N_18219,N_16702);
xnor U20393 (N_20393,N_13100,N_16523);
and U20394 (N_20394,N_13012,N_14979);
nand U20395 (N_20395,N_16224,N_15645);
nor U20396 (N_20396,N_16816,N_15674);
or U20397 (N_20397,N_17010,N_18572);
and U20398 (N_20398,N_17040,N_17147);
and U20399 (N_20399,N_17829,N_16565);
xor U20400 (N_20400,N_18476,N_14516);
nand U20401 (N_20401,N_18047,N_17874);
nor U20402 (N_20402,N_13145,N_17343);
xor U20403 (N_20403,N_16236,N_18253);
nor U20404 (N_20404,N_18032,N_14403);
and U20405 (N_20405,N_13627,N_16011);
nand U20406 (N_20406,N_16476,N_13277);
nand U20407 (N_20407,N_17000,N_17110);
and U20408 (N_20408,N_16151,N_16465);
nand U20409 (N_20409,N_18636,N_14047);
or U20410 (N_20410,N_17689,N_13613);
xor U20411 (N_20411,N_16851,N_17474);
nand U20412 (N_20412,N_16992,N_15127);
nand U20413 (N_20413,N_16100,N_13021);
nand U20414 (N_20414,N_12686,N_16562);
xor U20415 (N_20415,N_14489,N_13463);
nor U20416 (N_20416,N_16471,N_16648);
nand U20417 (N_20417,N_17256,N_13668);
and U20418 (N_20418,N_14366,N_16050);
xor U20419 (N_20419,N_18327,N_16867);
nand U20420 (N_20420,N_18322,N_17399);
xnor U20421 (N_20421,N_13421,N_16365);
nand U20422 (N_20422,N_12880,N_18239);
xor U20423 (N_20423,N_12518,N_12709);
nand U20424 (N_20424,N_14157,N_18510);
nor U20425 (N_20425,N_13641,N_13033);
nand U20426 (N_20426,N_14476,N_15627);
xor U20427 (N_20427,N_13123,N_14219);
or U20428 (N_20428,N_16613,N_18576);
xor U20429 (N_20429,N_17647,N_14378);
xnor U20430 (N_20430,N_15882,N_13433);
nand U20431 (N_20431,N_13083,N_17055);
and U20432 (N_20432,N_18384,N_16167);
nor U20433 (N_20433,N_12854,N_13075);
nand U20434 (N_20434,N_18566,N_17793);
nand U20435 (N_20435,N_18349,N_15025);
nand U20436 (N_20436,N_15317,N_17985);
nor U20437 (N_20437,N_14962,N_15926);
nor U20438 (N_20438,N_15887,N_18507);
nor U20439 (N_20439,N_15526,N_17804);
and U20440 (N_20440,N_14207,N_16278);
xnor U20441 (N_20441,N_18615,N_16560);
nor U20442 (N_20442,N_15230,N_13250);
xnor U20443 (N_20443,N_14246,N_14789);
or U20444 (N_20444,N_15582,N_14010);
nor U20445 (N_20445,N_13391,N_13170);
xnor U20446 (N_20446,N_18670,N_16475);
xnor U20447 (N_20447,N_15804,N_15147);
and U20448 (N_20448,N_18383,N_15568);
or U20449 (N_20449,N_14522,N_15808);
or U20450 (N_20450,N_17522,N_14209);
and U20451 (N_20451,N_12648,N_16844);
or U20452 (N_20452,N_17277,N_17639);
nor U20453 (N_20453,N_13102,N_13864);
nor U20454 (N_20454,N_13245,N_14659);
nand U20455 (N_20455,N_16556,N_15469);
xor U20456 (N_20456,N_18557,N_18672);
xnor U20457 (N_20457,N_13758,N_15244);
or U20458 (N_20458,N_14318,N_13505);
nor U20459 (N_20459,N_15378,N_16320);
nand U20460 (N_20460,N_16538,N_14849);
xor U20461 (N_20461,N_15058,N_12992);
nor U20462 (N_20462,N_15938,N_13749);
and U20463 (N_20463,N_12588,N_16196);
or U20464 (N_20464,N_17168,N_17254);
and U20465 (N_20465,N_17982,N_17723);
or U20466 (N_20466,N_14452,N_16722);
nand U20467 (N_20467,N_14738,N_15643);
or U20468 (N_20468,N_13713,N_14798);
nor U20469 (N_20469,N_13855,N_17007);
nor U20470 (N_20470,N_16940,N_14415);
or U20471 (N_20471,N_14300,N_16489);
nand U20472 (N_20472,N_14783,N_14515);
and U20473 (N_20473,N_16989,N_13768);
nand U20474 (N_20474,N_14130,N_18625);
nand U20475 (N_20475,N_14102,N_13844);
xor U20476 (N_20476,N_17818,N_16794);
nand U20477 (N_20477,N_18073,N_13352);
nand U20478 (N_20478,N_18623,N_15821);
or U20479 (N_20479,N_17852,N_14839);
nor U20480 (N_20480,N_13202,N_17807);
and U20481 (N_20481,N_15109,N_17802);
or U20482 (N_20482,N_15696,N_14982);
nand U20483 (N_20483,N_17709,N_14722);
and U20484 (N_20484,N_18570,N_16369);
or U20485 (N_20485,N_16864,N_16704);
xor U20486 (N_20486,N_14151,N_17627);
or U20487 (N_20487,N_14256,N_15139);
nand U20488 (N_20488,N_15116,N_13054);
and U20489 (N_20489,N_13801,N_14204);
xnor U20490 (N_20490,N_16272,N_15375);
nand U20491 (N_20491,N_12832,N_17707);
nand U20492 (N_20492,N_16800,N_16640);
and U20493 (N_20493,N_14078,N_13108);
nand U20494 (N_20494,N_16994,N_14459);
nor U20495 (N_20495,N_13010,N_15155);
and U20496 (N_20496,N_18508,N_14966);
nand U20497 (N_20497,N_17204,N_13995);
xnor U20498 (N_20498,N_18315,N_15084);
and U20499 (N_20499,N_13586,N_16653);
nor U20500 (N_20500,N_17954,N_16580);
nor U20501 (N_20501,N_12679,N_14127);
or U20502 (N_20502,N_17618,N_13380);
xnor U20503 (N_20503,N_18121,N_15920);
or U20504 (N_20504,N_12626,N_13847);
nor U20505 (N_20505,N_18425,N_16474);
xnor U20506 (N_20506,N_15909,N_18279);
xor U20507 (N_20507,N_16095,N_18521);
or U20508 (N_20508,N_17264,N_15597);
or U20509 (N_20509,N_18702,N_15095);
xnor U20510 (N_20510,N_12629,N_17914);
or U20511 (N_20511,N_13488,N_17455);
or U20512 (N_20512,N_15398,N_13742);
nor U20513 (N_20513,N_14984,N_13055);
or U20514 (N_20514,N_14308,N_12938);
xnor U20515 (N_20515,N_17381,N_15485);
xnor U20516 (N_20516,N_15851,N_17538);
nand U20517 (N_20517,N_16039,N_14796);
nor U20518 (N_20518,N_16111,N_17894);
and U20519 (N_20519,N_13101,N_14194);
nand U20520 (N_20520,N_18222,N_13998);
nor U20521 (N_20521,N_17554,N_16603);
nand U20522 (N_20522,N_16070,N_16246);
nor U20523 (N_20523,N_15272,N_18052);
nand U20524 (N_20524,N_17844,N_18701);
xor U20525 (N_20525,N_17942,N_16692);
nand U20526 (N_20526,N_14603,N_14191);
nand U20527 (N_20527,N_14596,N_18611);
nor U20528 (N_20528,N_18471,N_14537);
and U20529 (N_20529,N_17342,N_14731);
or U20530 (N_20530,N_18639,N_17058);
and U20531 (N_20531,N_13934,N_16126);
nor U20532 (N_20532,N_15550,N_14440);
or U20533 (N_20533,N_15168,N_18665);
xnor U20534 (N_20534,N_13800,N_18669);
and U20535 (N_20535,N_14752,N_18137);
and U20536 (N_20536,N_14702,N_17795);
xor U20537 (N_20537,N_13032,N_18727);
and U20538 (N_20538,N_16703,N_15864);
nor U20539 (N_20539,N_12808,N_16085);
or U20540 (N_20540,N_17086,N_12553);
or U20541 (N_20541,N_16850,N_17320);
or U20542 (N_20542,N_12987,N_18068);
and U20543 (N_20543,N_14469,N_17903);
nor U20544 (N_20544,N_17974,N_14395);
nor U20545 (N_20545,N_18218,N_13449);
and U20546 (N_20546,N_17372,N_16914);
nand U20547 (N_20547,N_13808,N_15006);
and U20548 (N_20548,N_16569,N_13982);
nor U20549 (N_20549,N_16383,N_15090);
or U20550 (N_20550,N_15679,N_14605);
nand U20551 (N_20551,N_16801,N_17435);
nand U20552 (N_20552,N_16416,N_13829);
nor U20553 (N_20553,N_15601,N_17104);
or U20554 (N_20554,N_17056,N_13207);
nor U20555 (N_20555,N_14788,N_15146);
and U20556 (N_20556,N_13308,N_17704);
and U20557 (N_20557,N_15480,N_13043);
nand U20558 (N_20558,N_16363,N_18679);
nand U20559 (N_20559,N_12997,N_13369);
and U20560 (N_20560,N_14057,N_17004);
and U20561 (N_20561,N_16901,N_15233);
nor U20562 (N_20562,N_14076,N_18455);
nand U20563 (N_20563,N_15859,N_16859);
nor U20564 (N_20564,N_12741,N_16526);
or U20565 (N_20565,N_18732,N_13885);
xnor U20566 (N_20566,N_17382,N_15694);
xor U20567 (N_20567,N_15187,N_14258);
nor U20568 (N_20568,N_17308,N_15577);
nor U20569 (N_20569,N_16116,N_16881);
xnor U20570 (N_20570,N_14182,N_16084);
nor U20571 (N_20571,N_14297,N_16296);
and U20572 (N_20572,N_13182,N_17978);
xor U20573 (N_20573,N_17642,N_16920);
and U20574 (N_20574,N_18360,N_16142);
xor U20575 (N_20575,N_12941,N_16403);
nor U20576 (N_20576,N_16845,N_14046);
nand U20577 (N_20577,N_14901,N_16622);
nor U20578 (N_20578,N_13726,N_16758);
and U20579 (N_20579,N_12984,N_18437);
xor U20580 (N_20580,N_17994,N_12917);
nor U20581 (N_20581,N_14729,N_15331);
or U20582 (N_20582,N_16351,N_18031);
nand U20583 (N_20583,N_17218,N_12650);
xor U20584 (N_20584,N_14610,N_17585);
or U20585 (N_20585,N_14411,N_17020);
nand U20586 (N_20586,N_16213,N_16135);
nor U20587 (N_20587,N_17872,N_13481);
xnor U20588 (N_20588,N_14091,N_15206);
and U20589 (N_20589,N_17705,N_15020);
nand U20590 (N_20590,N_17781,N_17386);
nand U20591 (N_20591,N_14268,N_13711);
or U20592 (N_20592,N_18090,N_14724);
xor U20593 (N_20593,N_18011,N_17046);
and U20594 (N_20594,N_13331,N_18364);
and U20595 (N_20595,N_17398,N_16086);
xnor U20596 (N_20596,N_14512,N_15814);
or U20597 (N_20597,N_14086,N_14558);
and U20598 (N_20598,N_14416,N_16742);
or U20599 (N_20599,N_18687,N_13975);
xnor U20600 (N_20600,N_15210,N_17763);
and U20601 (N_20601,N_15460,N_14749);
nand U20602 (N_20602,N_15004,N_18088);
and U20603 (N_20603,N_15595,N_14730);
or U20604 (N_20604,N_17824,N_18544);
and U20605 (N_20605,N_16721,N_16231);
nor U20606 (N_20606,N_14700,N_16461);
nor U20607 (N_20607,N_15080,N_18187);
and U20608 (N_20608,N_12855,N_15830);
or U20609 (N_20609,N_12724,N_14564);
nor U20610 (N_20610,N_18274,N_18562);
or U20611 (N_20611,N_15822,N_14069);
xor U20612 (N_20612,N_12989,N_14129);
xor U20613 (N_20613,N_18609,N_16250);
or U20614 (N_20614,N_15077,N_14068);
nor U20615 (N_20615,N_12527,N_17864);
nor U20616 (N_20616,N_16121,N_18730);
nor U20617 (N_20617,N_13445,N_16123);
nand U20618 (N_20618,N_17290,N_15452);
or U20619 (N_20619,N_15086,N_14794);
and U20620 (N_20620,N_17223,N_13528);
xnor U20621 (N_20621,N_18351,N_14446);
or U20622 (N_20622,N_12704,N_14540);
and U20623 (N_20623,N_16980,N_16262);
xor U20624 (N_20624,N_15240,N_12512);
and U20625 (N_20625,N_14955,N_16311);
nand U20626 (N_20626,N_18096,N_12962);
xnor U20627 (N_20627,N_15040,N_12582);
nand U20628 (N_20628,N_15936,N_14438);
xor U20629 (N_20629,N_18748,N_15356);
nor U20630 (N_20630,N_14264,N_15332);
nand U20631 (N_20631,N_13512,N_12544);
nor U20632 (N_20632,N_18123,N_17063);
nand U20633 (N_20633,N_17289,N_15847);
nand U20634 (N_20634,N_15693,N_17799);
xnor U20635 (N_20635,N_16564,N_13828);
or U20636 (N_20636,N_17897,N_13394);
xor U20637 (N_20637,N_15039,N_14051);
or U20638 (N_20638,N_13674,N_12927);
and U20639 (N_20639,N_14106,N_16944);
or U20640 (N_20640,N_15277,N_13723);
nor U20641 (N_20641,N_14999,N_14764);
and U20642 (N_20642,N_12752,N_14025);
and U20643 (N_20643,N_17591,N_14276);
and U20644 (N_20644,N_14253,N_14417);
nor U20645 (N_20645,N_13173,N_17099);
or U20646 (N_20646,N_13579,N_16671);
and U20647 (N_20647,N_17059,N_12759);
nand U20648 (N_20648,N_14400,N_15340);
nand U20649 (N_20649,N_16739,N_15059);
nand U20650 (N_20650,N_14309,N_13650);
or U20651 (N_20651,N_15432,N_15374);
or U20652 (N_20652,N_16611,N_13480);
nor U20653 (N_20653,N_12990,N_15973);
nor U20654 (N_20654,N_17302,N_14689);
nor U20655 (N_20655,N_13942,N_16925);
or U20656 (N_20656,N_13016,N_17975);
nor U20657 (N_20657,N_17674,N_12556);
and U20658 (N_20658,N_18024,N_17745);
xnor U20659 (N_20659,N_13590,N_13776);
nand U20660 (N_20660,N_13251,N_15678);
and U20661 (N_20661,N_16891,N_17573);
nand U20662 (N_20662,N_18158,N_15534);
and U20663 (N_20663,N_15019,N_18657);
and U20664 (N_20664,N_18622,N_17428);
or U20665 (N_20665,N_15141,N_18001);
or U20666 (N_20666,N_18745,N_16770);
and U20667 (N_20667,N_15055,N_18499);
and U20668 (N_20668,N_17509,N_18594);
nand U20669 (N_20669,N_16235,N_16699);
nand U20670 (N_20670,N_17834,N_14844);
or U20671 (N_20671,N_13883,N_15522);
or U20672 (N_20672,N_17867,N_17114);
and U20673 (N_20673,N_13228,N_13318);
and U20674 (N_20674,N_16089,N_12725);
and U20675 (N_20675,N_16107,N_17987);
nand U20676 (N_20676,N_18166,N_17426);
and U20677 (N_20677,N_12635,N_16542);
and U20678 (N_20678,N_15782,N_13666);
or U20679 (N_20679,N_17936,N_16310);
nand U20680 (N_20680,N_16117,N_15506);
or U20681 (N_20681,N_16338,N_18152);
and U20682 (N_20682,N_16760,N_15958);
and U20683 (N_20683,N_16715,N_15231);
nand U20684 (N_20684,N_15363,N_17313);
or U20685 (N_20685,N_14184,N_18415);
xnor U20686 (N_20686,N_17796,N_17138);
nor U20687 (N_20687,N_13899,N_14918);
and U20688 (N_20688,N_13039,N_16309);
or U20689 (N_20689,N_17425,N_18718);
xnor U20690 (N_20690,N_16216,N_14613);
nand U20691 (N_20691,N_13208,N_18367);
nand U20692 (N_20692,N_17950,N_17329);
or U20693 (N_20693,N_16402,N_15170);
nor U20694 (N_20694,N_13385,N_16880);
nand U20695 (N_20695,N_16247,N_17461);
nand U20696 (N_20696,N_14518,N_18352);
or U20697 (N_20697,N_16044,N_12536);
nor U20698 (N_20698,N_17923,N_13974);
or U20699 (N_20699,N_13247,N_13585);
xnor U20700 (N_20700,N_14530,N_13887);
xnor U20701 (N_20701,N_18236,N_12732);
or U20702 (N_20702,N_15586,N_18191);
or U20703 (N_20703,N_17939,N_14898);
xor U20704 (N_20704,N_16203,N_15490);
xnor U20705 (N_20705,N_12786,N_16843);
nor U20706 (N_20706,N_16455,N_14402);
xor U20707 (N_20707,N_15838,N_12825);
xnor U20708 (N_20708,N_15417,N_18348);
xnor U20709 (N_20709,N_13902,N_14572);
or U20710 (N_20710,N_15689,N_13792);
xor U20711 (N_20711,N_13256,N_14914);
nor U20712 (N_20712,N_15245,N_15482);
nor U20713 (N_20713,N_14940,N_15779);
or U20714 (N_20714,N_17196,N_18746);
xor U20715 (N_20715,N_13422,N_17750);
and U20716 (N_20716,N_16063,N_17497);
and U20717 (N_20717,N_13176,N_13440);
xor U20718 (N_20718,N_17498,N_18112);
nor U20719 (N_20719,N_12988,N_14389);
nand U20720 (N_20720,N_17132,N_18190);
or U20721 (N_20721,N_15446,N_18660);
xor U20722 (N_20722,N_13640,N_14845);
or U20723 (N_20723,N_17536,N_15896);
nor U20724 (N_20724,N_14165,N_14926);
nand U20725 (N_20725,N_12838,N_16753);
or U20726 (N_20726,N_16315,N_18366);
nand U20727 (N_20727,N_17333,N_12931);
nand U20728 (N_20728,N_18164,N_14753);
and U20729 (N_20729,N_16826,N_17595);
nand U20730 (N_20730,N_13879,N_14711);
and U20731 (N_20731,N_16802,N_18457);
xnor U20732 (N_20732,N_18195,N_18614);
and U20733 (N_20733,N_13093,N_16834);
nand U20734 (N_20734,N_15136,N_16058);
or U20735 (N_20735,N_14606,N_16092);
and U20736 (N_20736,N_16630,N_13898);
nor U20737 (N_20737,N_17165,N_17931);
nand U20738 (N_20738,N_18629,N_16427);
xnor U20739 (N_20739,N_12717,N_13297);
or U20740 (N_20740,N_14758,N_14175);
nor U20741 (N_20741,N_18058,N_15192);
xnor U20742 (N_20742,N_15108,N_18183);
and U20743 (N_20743,N_12958,N_16232);
nand U20744 (N_20744,N_13721,N_15701);
and U20745 (N_20745,N_17791,N_18533);
nor U20746 (N_20746,N_16333,N_13871);
xnor U20747 (N_20747,N_12533,N_18286);
and U20748 (N_20748,N_13329,N_18419);
nand U20749 (N_20749,N_16554,N_14307);
nand U20750 (N_20750,N_15329,N_13194);
nand U20751 (N_20751,N_18503,N_13338);
nand U20752 (N_20752,N_16207,N_18712);
and U20753 (N_20753,N_17771,N_17964);
xnor U20754 (N_20754,N_12577,N_12593);
nand U20755 (N_20755,N_12991,N_18640);
nand U20756 (N_20756,N_13925,N_14216);
nand U20757 (N_20757,N_16849,N_12833);
or U20758 (N_20758,N_16606,N_13785);
nor U20759 (N_20759,N_13159,N_18265);
nor U20760 (N_20760,N_13757,N_18439);
xor U20761 (N_20761,N_17596,N_12574);
nor U20762 (N_20762,N_14643,N_15142);
or U20763 (N_20763,N_18662,N_16799);
nor U20764 (N_20764,N_18003,N_18346);
nand U20765 (N_20765,N_13187,N_17480);
nand U20766 (N_20766,N_12865,N_14351);
xor U20767 (N_20767,N_15682,N_17367);
nand U20768 (N_20768,N_13376,N_14251);
and U20769 (N_20769,N_18142,N_13415);
and U20770 (N_20770,N_14614,N_18025);
nor U20771 (N_20771,N_13741,N_14815);
nor U20772 (N_20772,N_14359,N_17064);
nor U20773 (N_20773,N_15735,N_18449);
nor U20774 (N_20774,N_16584,N_14523);
and U20775 (N_20775,N_12919,N_17868);
nand U20776 (N_20776,N_16986,N_16510);
xor U20777 (N_20777,N_16106,N_15453);
nand U20778 (N_20778,N_13418,N_13794);
and U20779 (N_20779,N_16765,N_18230);
and U20780 (N_20780,N_16848,N_13429);
and U20781 (N_20781,N_17266,N_14821);
xnor U20782 (N_20782,N_13805,N_14628);
xnor U20783 (N_20783,N_14941,N_14163);
and U20784 (N_20784,N_17549,N_16481);
xor U20785 (N_20785,N_14220,N_17017);
and U20786 (N_20786,N_13275,N_16821);
nor U20787 (N_20787,N_18046,N_18299);
or U20788 (N_20788,N_12701,N_16060);
and U20789 (N_20789,N_14043,N_14247);
nand U20790 (N_20790,N_15685,N_12663);
xnor U20791 (N_20791,N_16180,N_15755);
and U20792 (N_20792,N_13546,N_15382);
nand U20793 (N_20793,N_13954,N_13180);
and U20794 (N_20794,N_12581,N_12985);
nor U20795 (N_20795,N_13217,N_17335);
and U20796 (N_20796,N_16346,N_12643);
or U20797 (N_20797,N_13731,N_12546);
xnor U20798 (N_20798,N_16146,N_18377);
nand U20799 (N_20799,N_16762,N_17637);
xnor U20800 (N_20800,N_17026,N_18323);
nor U20801 (N_20801,N_17779,N_13402);
xor U20802 (N_20802,N_14852,N_18196);
or U20803 (N_20803,N_14527,N_12731);
or U20804 (N_20804,N_13703,N_13314);
nand U20805 (N_20805,N_14703,N_13014);
xnor U20806 (N_20806,N_18412,N_16506);
nand U20807 (N_20807,N_14563,N_15609);
or U20808 (N_20808,N_14612,N_16299);
or U20809 (N_20809,N_17568,N_18565);
nor U20810 (N_20810,N_14948,N_12631);
nand U20811 (N_20811,N_16968,N_14149);
nand U20812 (N_20812,N_18373,N_17029);
nor U20813 (N_20813,N_17323,N_15990);
xnor U20814 (N_20814,N_18520,N_17699);
xnor U20815 (N_20815,N_14079,N_14499);
xnor U20816 (N_20816,N_14768,N_14650);
nor U20817 (N_20817,N_18206,N_13086);
or U20818 (N_20818,N_15313,N_15400);
nand U20819 (N_20819,N_13210,N_14887);
and U20820 (N_20820,N_18582,N_17021);
and U20821 (N_20821,N_16449,N_13427);
and U20822 (N_20822,N_14036,N_18685);
and U20823 (N_20823,N_12529,N_16181);
nor U20824 (N_20824,N_14044,N_13659);
nand U20825 (N_20825,N_18094,N_14553);
xnor U20826 (N_20826,N_15575,N_17615);
or U20827 (N_20827,N_14397,N_18432);
nor U20828 (N_20828,N_15441,N_13810);
nor U20829 (N_20829,N_14784,N_15801);
xnor U20830 (N_20830,N_14782,N_13676);
or U20831 (N_20831,N_12568,N_18316);
nor U20832 (N_20832,N_13812,N_14767);
nor U20833 (N_20833,N_13229,N_18287);
xor U20834 (N_20834,N_17537,N_16239);
nor U20835 (N_20835,N_15048,N_13632);
nor U20836 (N_20836,N_13688,N_17146);
xor U20837 (N_20837,N_16023,N_13193);
xnor U20838 (N_20838,N_17814,N_16303);
xnor U20839 (N_20839,N_17609,N_15037);
nand U20840 (N_20840,N_13305,N_13296);
nand U20841 (N_20841,N_17336,N_14326);
or U20842 (N_20842,N_17456,N_14740);
or U20843 (N_20843,N_13946,N_13443);
nor U20844 (N_20844,N_17008,N_15764);
or U20845 (N_20845,N_17624,N_17227);
xor U20846 (N_20846,N_18514,N_16270);
nor U20847 (N_20847,N_17334,N_16119);
and U20848 (N_20848,N_15458,N_15611);
nand U20849 (N_20849,N_14977,N_13383);
xnor U20850 (N_20850,N_14862,N_12963);
and U20851 (N_20851,N_15257,N_16462);
nor U20852 (N_20852,N_15209,N_12713);
or U20853 (N_20853,N_15690,N_15942);
xor U20854 (N_20854,N_17200,N_18721);
or U20855 (N_20855,N_12547,N_14226);
and U20856 (N_20856,N_16115,N_12953);
xnor U20857 (N_20857,N_17945,N_15337);
and U20858 (N_20858,N_18226,N_18242);
and U20859 (N_20859,N_16362,N_16933);
nor U20860 (N_20860,N_13447,N_17389);
xor U20861 (N_20861,N_13687,N_15253);
xor U20862 (N_20862,N_12622,N_12712);
or U20863 (N_20863,N_14514,N_16922);
xor U20864 (N_20864,N_14608,N_14723);
and U20865 (N_20865,N_13496,N_17992);
or U20866 (N_20866,N_13458,N_14358);
xor U20867 (N_20867,N_17009,N_17319);
and U20868 (N_20868,N_14180,N_18282);
nor U20869 (N_20869,N_18487,N_13874);
xnor U20870 (N_20870,N_15673,N_18194);
nand U20871 (N_20871,N_15268,N_13563);
xor U20872 (N_20872,N_15914,N_18682);
nand U20873 (N_20873,N_15965,N_17192);
and U20874 (N_20874,N_14176,N_16728);
or U20875 (N_20875,N_14477,N_16277);
or U20876 (N_20876,N_14410,N_13070);
xor U20877 (N_20877,N_18017,N_12726);
or U20878 (N_20878,N_16072,N_17442);
and U20879 (N_20879,N_16394,N_13292);
xor U20880 (N_20880,N_12604,N_14531);
and U20881 (N_20881,N_13456,N_15481);
nor U20882 (N_20882,N_12942,N_15989);
xor U20883 (N_20883,N_13375,N_17925);
or U20884 (N_20884,N_13026,N_12738);
nor U20885 (N_20885,N_13211,N_16938);
and U20886 (N_20886,N_17937,N_17013);
or U20887 (N_20887,N_17529,N_14777);
nor U20888 (N_20888,N_14221,N_16193);
and U20889 (N_20889,N_18051,N_13503);
and U20890 (N_20890,N_12716,N_12809);
or U20891 (N_20891,N_17470,N_16507);
nand U20892 (N_20892,N_14878,N_16179);
xnor U20893 (N_20893,N_17094,N_13790);
nor U20894 (N_20894,N_16861,N_15947);
or U20895 (N_20895,N_14312,N_13882);
nand U20896 (N_20896,N_13025,N_18035);
xnor U20897 (N_20897,N_16806,N_18408);
and U20898 (N_20898,N_17755,N_17407);
or U20899 (N_20899,N_15810,N_15600);
or U20900 (N_20900,N_12728,N_13060);
nor U20901 (N_20901,N_17905,N_17906);
nor U20902 (N_20902,N_14419,N_16932);
or U20903 (N_20903,N_17322,N_17024);
or U20904 (N_20904,N_12866,N_15427);
nand U20905 (N_20905,N_18555,N_13088);
xor U20906 (N_20906,N_16103,N_14077);
nand U20907 (N_20907,N_16756,N_18549);
xor U20908 (N_20908,N_15747,N_17053);
nand U20909 (N_20909,N_12843,N_12589);
and U20910 (N_20910,N_16408,N_17851);
nand U20911 (N_20911,N_15276,N_14535);
xor U20912 (N_20912,N_14187,N_16066);
and U20913 (N_20913,N_14814,N_15812);
xnor U20914 (N_20914,N_14517,N_16726);
and U20915 (N_20915,N_14277,N_17669);
nand U20916 (N_20916,N_13141,N_17812);
nand U20917 (N_20917,N_17631,N_13506);
xor U20918 (N_20918,N_16166,N_15120);
and U20919 (N_20919,N_18664,N_17786);
or U20920 (N_20920,N_13678,N_13466);
or U20921 (N_20921,N_17640,N_18593);
xor U20922 (N_20922,N_18150,N_17846);
nor U20923 (N_20923,N_16808,N_14448);
or U20924 (N_20924,N_13348,N_15935);
xnor U20925 (N_20925,N_13524,N_18118);
nand U20926 (N_20926,N_13547,N_16451);
and U20927 (N_20927,N_13453,N_14248);
and U20928 (N_20928,N_14924,N_16793);
xor U20929 (N_20929,N_16138,N_15151);
nor U20930 (N_20930,N_17294,N_15262);
nor U20931 (N_20931,N_13763,N_13147);
nand U20932 (N_20932,N_14936,N_12620);
nor U20933 (N_20933,N_18441,N_16540);
and U20934 (N_20934,N_13915,N_17967);
nor U20935 (N_20935,N_12612,N_15598);
nand U20936 (N_20936,N_18700,N_18472);
or U20937 (N_20937,N_16678,N_15945);
nand U20938 (N_20938,N_17219,N_17438);
xor U20939 (N_20939,N_15692,N_17900);
xnor U20940 (N_20940,N_12578,N_17838);
xor U20941 (N_20941,N_16388,N_16582);
or U20942 (N_20942,N_17434,N_14245);
nor U20943 (N_20943,N_15546,N_17490);
nand U20944 (N_20944,N_16139,N_14957);
nor U20945 (N_20945,N_13551,N_16984);
or U20946 (N_20946,N_16772,N_17606);
and U20947 (N_20947,N_13144,N_15163);
nand U20948 (N_20948,N_16885,N_16820);
nand U20949 (N_20949,N_17712,N_15823);
xor U20950 (N_20950,N_13983,N_18529);
or U20951 (N_20951,N_12531,N_15842);
and U20952 (N_20952,N_18628,N_17821);
nand U20953 (N_20953,N_16587,N_12627);
nand U20954 (N_20954,N_18185,N_14906);
xnor U20955 (N_20955,N_15402,N_13061);
nand U20956 (N_20956,N_16433,N_17338);
or U20957 (N_20957,N_16133,N_15574);
nand U20958 (N_20958,N_15005,N_18532);
and U20959 (N_20959,N_12932,N_15835);
xor U20960 (N_20960,N_14586,N_16626);
nor U20961 (N_20961,N_12535,N_16048);
or U20962 (N_20962,N_18070,N_18617);
or U20963 (N_20963,N_16168,N_12928);
or U20964 (N_20964,N_17083,N_14829);
nor U20965 (N_20965,N_15553,N_18447);
or U20966 (N_20966,N_15472,N_17002);
and U20967 (N_20967,N_18165,N_13205);
xor U20968 (N_20968,N_13234,N_15478);
xnor U20969 (N_20969,N_15035,N_16735);
and U20970 (N_20970,N_16832,N_14374);
nand U20971 (N_20971,N_13921,N_17310);
xnor U20972 (N_20972,N_13920,N_17118);
nor U20973 (N_20973,N_15102,N_18674);
nor U20974 (N_20974,N_14019,N_18405);
and U20975 (N_20975,N_17766,N_12642);
nor U20976 (N_20976,N_15302,N_14274);
and U20977 (N_20977,N_16024,N_17789);
nand U20978 (N_20978,N_15174,N_14903);
nand U20979 (N_20979,N_16732,N_13414);
nor U20980 (N_20980,N_16685,N_15010);
nor U20981 (N_20981,N_16379,N_18645);
or U20982 (N_20982,N_12688,N_14993);
nand U20983 (N_20983,N_14494,N_15978);
xnor U20984 (N_20984,N_17731,N_17141);
nor U20985 (N_20985,N_15951,N_15171);
nand U20986 (N_20986,N_15183,N_16521);
or U20987 (N_20987,N_13589,N_17883);
xnor U20988 (N_20988,N_14431,N_17390);
and U20989 (N_20989,N_17457,N_17780);
nor U20990 (N_20990,N_17893,N_13046);
or U20991 (N_20991,N_18120,N_13020);
and U20992 (N_20992,N_17613,N_14561);
and U20993 (N_20993,N_14915,N_15508);
or U20994 (N_20994,N_13353,N_13288);
nor U20995 (N_20995,N_17809,N_12844);
nand U20996 (N_20996,N_14988,N_14208);
xnor U20997 (N_20997,N_17130,N_15165);
and U20998 (N_20998,N_18053,N_17603);
and U20999 (N_20999,N_13819,N_18605);
or U21000 (N_21000,N_15373,N_17003);
nand U21001 (N_21001,N_18661,N_14812);
and U21002 (N_21002,N_13695,N_15984);
or U21003 (N_21003,N_14352,N_17778);
and U21004 (N_21004,N_17101,N_13358);
and U21005 (N_21005,N_17495,N_12852);
or U21006 (N_21006,N_12875,N_14550);
or U21007 (N_21007,N_17861,N_16155);
xnor U21008 (N_21008,N_17855,N_17019);
nand U21009 (N_21009,N_15959,N_16150);
nor U21010 (N_21010,N_12766,N_17245);
or U21011 (N_21011,N_12514,N_16343);
nand U21012 (N_21012,N_18122,N_17318);
and U21013 (N_21013,N_12944,N_15641);
nor U21014 (N_21014,N_15051,N_16547);
nor U21015 (N_21015,N_13365,N_13044);
or U21016 (N_21016,N_12922,N_15412);
nor U21017 (N_21017,N_14616,N_16395);
or U21018 (N_21018,N_14085,N_13935);
xor U21019 (N_21019,N_14889,N_15345);
and U21020 (N_21020,N_15228,N_17561);
nor U21021 (N_21021,N_17178,N_15819);
or U21022 (N_21022,N_18649,N_14328);
nor U21023 (N_21023,N_13894,N_15769);
xnor U21024 (N_21024,N_15535,N_14778);
nor U21025 (N_21025,N_14442,N_17360);
or U21026 (N_21026,N_15869,N_16695);
xor U21027 (N_21027,N_18045,N_13519);
or U21028 (N_21028,N_16610,N_18110);
or U21029 (N_21029,N_18607,N_15361);
and U21030 (N_21030,N_15191,N_17876);
xnor U21031 (N_21031,N_14369,N_17854);
nor U21032 (N_21032,N_13549,N_15323);
nand U21033 (N_21033,N_18406,N_13833);
and U21034 (N_21034,N_15263,N_13347);
or U21035 (N_21035,N_13811,N_17066);
nor U21036 (N_21036,N_18445,N_16041);
xnor U21037 (N_21037,N_14881,N_15069);
nand U21038 (N_21038,N_13191,N_18143);
nor U21039 (N_21039,N_18372,N_15306);
or U21040 (N_21040,N_18381,N_14364);
and U21041 (N_21041,N_15392,N_15520);
nor U21042 (N_21042,N_13966,N_17074);
or U21043 (N_21043,N_15659,N_15907);
and U21044 (N_21044,N_17882,N_15360);
or U21045 (N_21045,N_13751,N_17123);
or U21046 (N_21046,N_14028,N_13056);
and U21047 (N_21047,N_16487,N_13637);
nand U21048 (N_21048,N_17570,N_13403);
nand U21049 (N_21049,N_15599,N_14566);
nand U21050 (N_21050,N_14254,N_15684);
or U21051 (N_21051,N_13121,N_13166);
and U21052 (N_21052,N_14732,N_15011);
xnor U21053 (N_21053,N_17831,N_13765);
or U21054 (N_21054,N_16971,N_13162);
or U21055 (N_21055,N_13069,N_16637);
and U21056 (N_21056,N_18435,N_13022);
xor U21057 (N_21057,N_13753,N_15128);
xor U21058 (N_21058,N_14456,N_14973);
or U21059 (N_21059,N_17142,N_13077);
and U21060 (N_21060,N_17297,N_12756);
or U21061 (N_21061,N_15213,N_13408);
xnor U21062 (N_21062,N_16504,N_16407);
or U21063 (N_21063,N_18344,N_18436);
nand U21064 (N_21064,N_17378,N_13509);
xor U21065 (N_21065,N_16192,N_18086);
xnor U21066 (N_21066,N_13714,N_13281);
and U21067 (N_21067,N_14567,N_13209);
nor U21068 (N_21068,N_15855,N_16910);
nand U21069 (N_21069,N_13441,N_14161);
nand U21070 (N_21070,N_14119,N_16836);
xnor U21071 (N_21071,N_18574,N_13598);
xnor U21072 (N_21072,N_16539,N_14831);
nor U21073 (N_21073,N_13454,N_15854);
nand U21074 (N_21074,N_12760,N_14012);
and U21075 (N_21075,N_13224,N_13168);
or U21076 (N_21076,N_14931,N_15529);
nor U21077 (N_21077,N_14444,N_16761);
xor U21078 (N_21078,N_18281,N_15656);
nor U21079 (N_21079,N_13686,N_12926);
xnor U21080 (N_21080,N_16002,N_13393);
or U21081 (N_21081,N_15704,N_17832);
or U21082 (N_21082,N_14910,N_16911);
nand U21083 (N_21083,N_15161,N_13186);
nand U21084 (N_21084,N_16937,N_13857);
or U21085 (N_21085,N_16666,N_18254);
nor U21086 (N_21086,N_12906,N_13685);
and U21087 (N_21087,N_15632,N_14437);
xnor U21088 (N_21088,N_13600,N_13671);
or U21089 (N_21089,N_14976,N_16297);
or U21090 (N_21090,N_14747,N_15372);
xnor U21091 (N_21091,N_17988,N_15021);
nand U21092 (N_21092,N_13542,N_16124);
xnor U21093 (N_21093,N_18681,N_13048);
xor U21094 (N_21094,N_16289,N_14813);
xor U21095 (N_21095,N_18379,N_14133);
xor U21096 (N_21096,N_13821,N_12907);
and U21097 (N_21097,N_14833,N_13152);
xnor U21098 (N_21098,N_12952,N_16370);
and U21099 (N_21099,N_16368,N_13143);
nor U21100 (N_21100,N_17237,N_12885);
or U21101 (N_21101,N_14511,N_15158);
nor U21102 (N_21102,N_15416,N_15314);
nor U21103 (N_21103,N_18198,N_18131);
nand U21104 (N_21104,N_17678,N_18552);
or U21105 (N_21105,N_12585,N_12798);
xor U21106 (N_21106,N_12564,N_13198);
and U21107 (N_21107,N_16001,N_17205);
or U21108 (N_21108,N_18513,N_16511);
or U21109 (N_21109,N_16936,N_13968);
and U21110 (N_21110,N_12519,N_13489);
nand U21111 (N_21111,N_13124,N_13396);
nor U21112 (N_21112,N_14322,N_14555);
nand U21113 (N_21113,N_17767,N_17933);
nand U21114 (N_21114,N_15930,N_14426);
nor U21115 (N_21115,N_18356,N_12757);
and U21116 (N_21116,N_16009,N_17233);
nand U21117 (N_21117,N_17283,N_13872);
nor U21118 (N_21118,N_15621,N_17493);
nor U21119 (N_21119,N_15786,N_12754);
or U21120 (N_21120,N_12730,N_16005);
and U21121 (N_21121,N_15607,N_14663);
and U21122 (N_21122,N_12851,N_13941);
or U21123 (N_21123,N_15640,N_13518);
and U21124 (N_21124,N_12706,N_13346);
and U21125 (N_21125,N_16318,N_15012);
or U21126 (N_21126,N_13845,N_15780);
or U21127 (N_21127,N_14763,N_15406);
nand U21128 (N_21128,N_12708,N_16469);
and U21129 (N_21129,N_14890,N_14097);
and U21130 (N_21130,N_15387,N_13137);
nand U21131 (N_21131,N_17491,N_17330);
nand U21132 (N_21132,N_18560,N_16853);
nand U21133 (N_21133,N_16548,N_16965);
and U21134 (N_21134,N_16917,N_13132);
nor U21135 (N_21135,N_16458,N_17926);
nor U21136 (N_21136,N_16013,N_15820);
nor U21137 (N_21137,N_13566,N_14458);
xor U21138 (N_21138,N_16281,N_18161);
xnor U21139 (N_21139,N_18689,N_17102);
nand U21140 (N_21140,N_18189,N_17298);
xor U21141 (N_21141,N_14513,N_16434);
nand U21142 (N_21142,N_13665,N_17400);
nand U21143 (N_21143,N_12918,N_14200);
nand U21144 (N_21144,N_14919,N_18486);
nand U21145 (N_21145,N_16878,N_17582);
nand U21146 (N_21146,N_16948,N_13837);
nor U21147 (N_21147,N_12702,N_16818);
nand U21148 (N_21148,N_15326,N_17250);
nor U21149 (N_21149,N_13336,N_18201);
xor U21150 (N_21150,N_12523,N_18410);
or U21151 (N_21151,N_18291,N_13963);
xor U21152 (N_21152,N_13560,N_13973);
xor U21153 (N_21153,N_16222,N_12879);
or U21154 (N_21154,N_17337,N_13556);
xor U21155 (N_21155,N_18741,N_13780);
xor U21156 (N_21156,N_18502,N_13118);
nor U21157 (N_21157,N_12839,N_15479);
and U21158 (N_21158,N_16419,N_18723);
and U21159 (N_21159,N_16674,N_16334);
or U21160 (N_21160,N_15426,N_13388);
nor U21161 (N_21161,N_14342,N_13962);
nand U21162 (N_21162,N_18668,N_16398);
nand U21163 (N_21163,N_17714,N_14551);
nand U21164 (N_21164,N_17835,N_15639);
xor U21165 (N_21165,N_18097,N_18006);
xnor U21166 (N_21166,N_13483,N_13826);
and U21167 (N_21167,N_14793,N_15029);
and U21168 (N_21168,N_16655,N_13558);
or U21169 (N_21169,N_16325,N_18126);
nand U21170 (N_21170,N_17421,N_14868);
or U21171 (N_21171,N_13448,N_15793);
nor U21172 (N_21172,N_14980,N_16638);
xnor U21173 (N_21173,N_15873,N_13856);
and U21174 (N_21174,N_12955,N_16267);
nand U21175 (N_21175,N_17762,N_17352);
xor U21176 (N_21176,N_13085,N_16218);
xor U21177 (N_21177,N_14288,N_14640);
nand U21178 (N_21178,N_15980,N_13002);
nand U21179 (N_21179,N_17681,N_16838);
nand U21180 (N_21180,N_13992,N_17211);
and U21181 (N_21181,N_16957,N_12505);
or U21182 (N_21182,N_13525,N_16586);
or U21183 (N_21183,N_17225,N_17199);
xnor U21184 (N_21184,N_18526,N_18033);
nor U21185 (N_21185,N_14799,N_13007);
nor U21186 (N_21186,N_12889,N_16341);
nand U21187 (N_21187,N_16889,N_18698);
or U21188 (N_21188,N_12810,N_14105);
xor U21189 (N_21189,N_12710,N_14243);
xor U21190 (N_21190,N_15596,N_14436);
or U21191 (N_21191,N_15106,N_16571);
nand U21192 (N_21192,N_17717,N_18303);
and U21193 (N_21193,N_12768,N_14168);
nand U21194 (N_21194,N_16215,N_14588);
xor U21195 (N_21195,N_18391,N_15330);
nand U21196 (N_21196,N_13775,N_18671);
nand U21197 (N_21197,N_13644,N_16410);
or U21198 (N_21198,N_13177,N_17207);
xor U21199 (N_21199,N_12803,N_13319);
and U21200 (N_21200,N_15110,N_17288);
xor U21201 (N_21201,N_15465,N_14372);
or U21202 (N_21202,N_15563,N_15923);
xnor U21203 (N_21203,N_14819,N_15557);
or U21204 (N_21204,N_17458,N_17823);
or U21205 (N_21205,N_13682,N_15255);
xor U21206 (N_21206,N_12974,N_14070);
or U21207 (N_21207,N_12968,N_12899);
or U21208 (N_21208,N_16719,N_15341);
and U21209 (N_21209,N_12824,N_16429);
nand U21210 (N_21210,N_14120,N_15648);
xnor U21211 (N_21211,N_14370,N_17783);
nor U21212 (N_21212,N_13110,N_14002);
or U21213 (N_21213,N_15885,N_17949);
nand U21214 (N_21214,N_13045,N_14255);
nand U21215 (N_21215,N_12669,N_14647);
nand U21216 (N_21216,N_14225,N_12711);
nor U21217 (N_21217,N_17759,N_14332);
nand U21218 (N_21218,N_16601,N_14600);
nor U21219 (N_21219,N_12861,N_15584);
nor U21220 (N_21220,N_13911,N_16006);
and U21221 (N_21221,N_15649,N_13300);
nand U21222 (N_21222,N_17280,N_16360);
nor U21223 (N_21223,N_13262,N_18091);
nand U21224 (N_21224,N_13510,N_14325);
nor U21225 (N_21225,N_16675,N_15122);
nor U21226 (N_21226,N_16959,N_13188);
nand U21227 (N_21227,N_14020,N_14547);
xor U21228 (N_21228,N_16230,N_14391);
nor U21229 (N_21229,N_15397,N_15785);
xnor U21230 (N_21230,N_16027,N_13859);
or U21231 (N_21231,N_16641,N_17299);
xnor U21232 (N_21232,N_17355,N_17576);
nor U21233 (N_21233,N_13623,N_16137);
nand U21234 (N_21234,N_15971,N_13952);
nand U21235 (N_21235,N_17922,N_14840);
nand U21236 (N_21236,N_17758,N_16633);
nor U21237 (N_21237,N_13709,N_13309);
and U21238 (N_21238,N_16927,N_17577);
or U21239 (N_21239,N_18332,N_12797);
xor U21240 (N_21240,N_12787,N_14759);
xnor U21241 (N_21241,N_14593,N_15103);
and U21242 (N_21242,N_14694,N_12765);
xor U21243 (N_21243,N_16358,N_14049);
or U21244 (N_21244,N_14147,N_16280);
nand U21245 (N_21245,N_14385,N_12668);
or U21246 (N_21246,N_17031,N_13950);
nor U21247 (N_21247,N_15552,N_12576);
or U21248 (N_21248,N_17248,N_14824);
nand U21249 (N_21249,N_17944,N_15044);
xnor U21250 (N_21250,N_18295,N_15421);
and U21251 (N_21251,N_15530,N_13858);
and U21252 (N_21252,N_17629,N_18333);
and U21253 (N_21253,N_15698,N_16283);
xor U21254 (N_21254,N_18228,N_14427);
xnor U21255 (N_21255,N_14084,N_15234);
nand U21256 (N_21256,N_15628,N_18100);
or U21257 (N_21257,N_16080,N_14769);
nor U21258 (N_21258,N_17413,N_14971);
or U21259 (N_21259,N_17471,N_12978);
or U21260 (N_21260,N_14792,N_15671);
or U21261 (N_21261,N_14345,N_18388);
xor U21262 (N_21262,N_14802,N_16512);
xor U21263 (N_21263,N_16751,N_18450);
nor U21264 (N_21264,N_14856,N_13853);
xor U21265 (N_21265,N_15531,N_16285);
and U21266 (N_21266,N_18448,N_18528);
or U21267 (N_21267,N_18564,N_12624);
or U21268 (N_21268,N_16012,N_14376);
or U21269 (N_21269,N_13559,N_14261);
nor U21270 (N_21270,N_18240,N_13541);
nand U21271 (N_21271,N_13249,N_18506);
or U21272 (N_21272,N_18589,N_14686);
nor U21273 (N_21273,N_15430,N_15451);
or U21274 (N_21274,N_16047,N_16169);
nor U21275 (N_21275,N_17363,N_12530);
nor U21276 (N_21276,N_13778,N_17210);
and U21277 (N_21277,N_14496,N_14706);
or U21278 (N_21278,N_16682,N_15564);
and U21279 (N_21279,N_15473,N_16664);
and U21280 (N_21280,N_15249,N_14420);
nor U21281 (N_21281,N_12616,N_15658);
or U21282 (N_21282,N_15998,N_17039);
nand U21283 (N_21283,N_16677,N_16782);
nand U21284 (N_21284,N_18691,N_16976);
nor U21285 (N_21285,N_15903,N_16684);
or U21286 (N_21286,N_16156,N_17911);
xor U21287 (N_21287,N_17927,N_16950);
nand U21288 (N_21288,N_12534,N_15807);
nor U21289 (N_21289,N_18504,N_14787);
xor U21290 (N_21290,N_14765,N_12559);
or U21291 (N_21291,N_18109,N_16488);
xor U21292 (N_21292,N_18380,N_15089);
and U21293 (N_21293,N_13107,N_17516);
xnor U21294 (N_21294,N_12503,N_14497);
nand U21295 (N_21295,N_18276,N_14132);
or U21296 (N_21296,N_12881,N_13467);
nor U21297 (N_21297,N_17760,N_14414);
or U21298 (N_21298,N_18371,N_18246);
nand U21299 (N_21299,N_18396,N_17645);
nand U21300 (N_21300,N_13922,N_13550);
and U21301 (N_21301,N_15395,N_13534);
nand U21302 (N_21302,N_12937,N_17690);
and U21303 (N_21303,N_16817,N_18378);
xor U21304 (N_21304,N_15912,N_17917);
nand U21305 (N_21305,N_15503,N_17353);
nand U21306 (N_21306,N_17068,N_17995);
and U21307 (N_21307,N_13004,N_18084);
nor U21308 (N_21308,N_17087,N_15440);
and U21309 (N_21309,N_16328,N_13327);
nor U21310 (N_21310,N_13036,N_16031);
or U21311 (N_21311,N_13587,N_16397);
or U21312 (N_21312,N_14843,N_12761);
or U21313 (N_21313,N_16689,N_12586);
xor U21314 (N_21314,N_16337,N_17890);
and U21315 (N_21315,N_13128,N_17344);
or U21316 (N_21316,N_15712,N_12583);
xor U21317 (N_21317,N_12619,N_12657);
xor U21318 (N_21318,N_18243,N_16260);
xnor U21319 (N_21319,N_16809,N_17506);
nor U21320 (N_21320,N_14023,N_14029);
nor U21321 (N_21321,N_13799,N_14305);
or U21322 (N_21322,N_15845,N_15653);
or U21323 (N_21323,N_13807,N_14524);
nand U21324 (N_21324,N_13782,N_18019);
or U21325 (N_21325,N_17708,N_13265);
and U21326 (N_21326,N_17437,N_17959);
xnor U21327 (N_21327,N_18641,N_14725);
xor U21328 (N_21328,N_13508,N_17149);
xnor U21329 (N_21329,N_18266,N_17963);
xnor U21330 (N_21330,N_16335,N_18598);
xor U21331 (N_21331,N_16876,N_15638);
nand U21332 (N_21332,N_15104,N_12807);
or U21333 (N_21333,N_14093,N_15884);
xnor U21334 (N_21334,N_14330,N_17514);
or U21335 (N_21335,N_16807,N_18320);
or U21336 (N_21336,N_12979,N_15940);
nor U21337 (N_21337,N_14178,N_13786);
nand U21338 (N_21338,N_17235,N_14580);
xor U21339 (N_21339,N_13322,N_17107);
or U21340 (N_21340,N_13477,N_13142);
or U21341 (N_21341,N_15983,N_13532);
xnor U21342 (N_21342,N_17078,N_14237);
nor U21343 (N_21343,N_15056,N_17079);
nand U21344 (N_21344,N_12830,N_14283);
nand U21345 (N_21345,N_13189,N_15218);
xnor U21346 (N_21346,N_18495,N_17940);
xor U21347 (N_21347,N_17912,N_16108);
xor U21348 (N_21348,N_14294,N_16091);
or U21349 (N_21349,N_12662,N_15082);
nor U21350 (N_21350,N_16609,N_12900);
and U21351 (N_21351,N_13267,N_17246);
and U21352 (N_21352,N_15519,N_16588);
or U21353 (N_21353,N_15411,N_14592);
and U21354 (N_21354,N_18599,N_13349);
nor U21355 (N_21355,N_17756,N_17722);
xnor U21356 (N_21356,N_14021,N_16964);
nand U21357 (N_21357,N_13285,N_16258);
nor U21358 (N_21358,N_16174,N_15933);
nor U21359 (N_21359,N_15401,N_12795);
nand U21360 (N_21360,N_13702,N_12771);
nor U21361 (N_21361,N_12590,N_16287);
or U21362 (N_21362,N_13886,N_13105);
and U21363 (N_21363,N_13324,N_17300);
nor U21364 (N_21364,N_13788,N_18735);
and U21365 (N_21365,N_16754,N_13522);
and U21366 (N_21366,N_14529,N_14545);
nand U21367 (N_21367,N_15827,N_13748);
xnor U21368 (N_21368,N_17301,N_12618);
xor U21369 (N_21369,N_16186,N_16708);
or U21370 (N_21370,N_17451,N_12884);
xor U21371 (N_21371,N_17041,N_12893);
xor U21372 (N_21372,N_14272,N_18350);
nand U21373 (N_21373,N_16374,N_12625);
and U21374 (N_21374,N_14142,N_14604);
nor U21375 (N_21375,N_14618,N_13933);
or U21376 (N_21376,N_16294,N_13227);
or U21377 (N_21377,N_17405,N_13103);
nor U21378 (N_21378,N_15322,N_17726);
nor U21379 (N_21379,N_15429,N_17720);
and U21380 (N_21380,N_14148,N_13174);
xor U21381 (N_21381,N_13697,N_16903);
nand U21382 (N_21382,N_14169,N_17359);
nand U21383 (N_21383,N_16208,N_16731);
and U21384 (N_21384,N_13698,N_14921);
and U21385 (N_21385,N_13106,N_17295);
and U21386 (N_21386,N_12764,N_17193);
or U21387 (N_21387,N_14257,N_18144);
nand U21388 (N_21388,N_14445,N_16161);
xnor U21389 (N_21389,N_12543,N_12998);
xnor U21390 (N_21390,N_14360,N_14185);
nor U21391 (N_21391,N_16245,N_18382);
and U21392 (N_21392,N_17747,N_15538);
nor U21393 (N_21393,N_17980,N_18397);
xor U21394 (N_21394,N_16456,N_15214);
and U21395 (N_21395,N_14693,N_13957);
and U21396 (N_21396,N_18192,N_13148);
nor U21397 (N_21397,N_13827,N_15399);
nor U21398 (N_21398,N_17189,N_18525);
xnor U21399 (N_21399,N_16967,N_12613);
nor U21400 (N_21400,N_17650,N_18027);
nand U21401 (N_21401,N_17241,N_18454);
nand U21402 (N_21402,N_18573,N_18176);
nand U21403 (N_21403,N_17580,N_17673);
or U21404 (N_21404,N_16600,N_16447);
and U21405 (N_21405,N_18479,N_15509);
nand U21406 (N_21406,N_13984,N_12665);
nor U21407 (N_21407,N_15744,N_17152);
or U21408 (N_21408,N_16872,N_17311);
nand U21409 (N_21409,N_15560,N_16559);
nand U21410 (N_21410,N_14683,N_14861);
and U21411 (N_21411,N_15063,N_18359);
or U21412 (N_21412,N_16714,N_15105);
nand U21413 (N_21413,N_14651,N_17749);
nor U21414 (N_21414,N_13084,N_15633);
and U21415 (N_21415,N_13255,N_13591);
and U21416 (N_21416,N_12873,N_14189);
nor U21417 (N_21417,N_13492,N_14339);
xor U21418 (N_21418,N_14398,N_14581);
nand U21419 (N_21419,N_16572,N_16931);
nor U21420 (N_21420,N_17221,N_13031);
nand U21421 (N_21421,N_17746,N_18595);
or U21422 (N_21422,N_17124,N_17424);
or U21423 (N_21423,N_17881,N_13236);
nand U21424 (N_21424,N_15967,N_15618);
nand U21425 (N_21425,N_17025,N_14131);
or U21426 (N_21426,N_13592,N_12654);
xnor U21427 (N_21427,N_17548,N_16918);
xnor U21428 (N_21428,N_18558,N_13823);
nand U21429 (N_21429,N_18257,N_13900);
and U21430 (N_21430,N_16375,N_15113);
nand U21431 (N_21431,N_17095,N_13694);
nand U21432 (N_21432,N_17356,N_16599);
nor U21433 (N_21433,N_13907,N_13959);
nor U21434 (N_21434,N_17362,N_17526);
and U21435 (N_21435,N_17443,N_15298);
or U21436 (N_21436,N_16421,N_15241);
and U21437 (N_21437,N_15117,N_17887);
or U21438 (N_21438,N_18167,N_13062);
nand U21439 (N_21439,N_14672,N_15893);
nand U21440 (N_21440,N_12692,N_18041);
xor U21441 (N_21441,N_18127,N_18043);
nor U21442 (N_21442,N_14958,N_18133);
nand U21443 (N_21443,N_17551,N_15015);
and U21444 (N_21444,N_17958,N_16088);
nor U21445 (N_21445,N_15687,N_14239);
nand U21446 (N_21446,N_12500,N_13115);
and U21447 (N_21447,N_14233,N_13880);
nor U21448 (N_21448,N_15219,N_15085);
or U21449 (N_21449,N_16884,N_16191);
and U21450 (N_21450,N_15540,N_14236);
nand U21451 (N_21451,N_18251,N_15710);
xnor U21452 (N_21452,N_14583,N_13342);
or U21453 (N_21453,N_14905,N_17564);
or U21454 (N_21454,N_16894,N_14040);
and U21455 (N_21455,N_15195,N_17140);
or U21456 (N_21456,N_15076,N_18462);
nor U21457 (N_21457,N_14075,N_13578);
nand U21458 (N_21458,N_17126,N_14685);
nand U21459 (N_21459,N_17429,N_13215);
xor U21460 (N_21460,N_15758,N_18223);
or U21461 (N_21461,N_15612,N_17546);
nor U21462 (N_21462,N_14520,N_13516);
and U21463 (N_21463,N_16073,N_14117);
xor U21464 (N_21464,N_13271,N_14549);
xor U21465 (N_21465,N_16625,N_13064);
nand U21466 (N_21466,N_16190,N_15994);
xnor U21467 (N_21467,N_18357,N_13355);
and U21468 (N_21468,N_13006,N_13628);
nand U21469 (N_21469,N_14775,N_17148);
nand U21470 (N_21470,N_15603,N_17979);
nor U21471 (N_21471,N_16219,N_14455);
nor U21472 (N_21472,N_14795,N_14144);
or U21473 (N_21473,N_17197,N_14421);
nand U21474 (N_21474,N_17513,N_18021);
nor U21475 (N_21475,N_17792,N_13430);
nand U21476 (N_21476,N_18034,N_17242);
and U21477 (N_21477,N_13781,N_15093);
xnor U21478 (N_21478,N_14809,N_15722);
xnor U21479 (N_21479,N_17260,N_14461);
xor U21480 (N_21480,N_16399,N_14430);
nor U21481 (N_21481,N_13472,N_15919);
xor U21482 (N_21482,N_18501,N_12672);
or U21483 (N_21483,N_17505,N_13473);
and U21484 (N_21484,N_14928,N_14394);
and U21485 (N_21485,N_12682,N_15499);
nor U21486 (N_21486,N_15925,N_14698);
nand U21487 (N_21487,N_14987,N_16659);
nand U21488 (N_21488,N_13218,N_17408);
or U21489 (N_21489,N_15824,N_17608);
nand U21490 (N_21490,N_15924,N_15054);
xor U21491 (N_21491,N_14847,N_18401);
and U21492 (N_21492,N_16067,N_18319);
nor U21493 (N_21493,N_14418,N_14960);
nand U21494 (N_21494,N_14594,N_14121);
or U21495 (N_21495,N_14676,N_13639);
or U21496 (N_21496,N_14473,N_17234);
nand U21497 (N_21497,N_14985,N_15517);
nor U21498 (N_21498,N_13471,N_12864);
and U21499 (N_21499,N_16237,N_13904);
or U21500 (N_21500,N_18141,N_13469);
nor U21501 (N_21501,N_15175,N_14811);
nor U21502 (N_21502,N_15946,N_14095);
or U21503 (N_21503,N_17932,N_16171);
and U21504 (N_21504,N_13474,N_15585);
nand U21505 (N_21505,N_15098,N_16882);
nand U21506 (N_21506,N_18647,N_13814);
nor U21507 (N_21507,N_13374,N_14670);
nor U21508 (N_21508,N_16372,N_16035);
nand U21509 (N_21509,N_13708,N_17475);
nand U21510 (N_21510,N_17880,N_15438);
xnor U21511 (N_21511,N_14071,N_16454);
and U21512 (N_21512,N_15672,N_18646);
xnor U21513 (N_21513,N_15811,N_18489);
or U21514 (N_21514,N_14846,N_15777);
or U21515 (N_21515,N_13552,N_18363);
or U21516 (N_21516,N_16154,N_14323);
nand U21517 (N_21517,N_14942,N_14922);
nor U21518 (N_21518,N_15708,N_14462);
nand U21519 (N_21519,N_13727,N_13455);
xor U21520 (N_21520,N_15486,N_14266);
nand U21521 (N_21521,N_17238,N_14026);
nor U21522 (N_21522,N_16865,N_18314);
or U21523 (N_21523,N_16929,N_14429);
or U21524 (N_21524,N_18429,N_13730);
or U21525 (N_21525,N_14668,N_17069);
xor U21526 (N_21526,N_13842,N_18404);
and U21527 (N_21527,N_15172,N_15532);
or U21528 (N_21528,N_15222,N_13241);
xor U21529 (N_21529,N_16339,N_14761);
nand U21530 (N_21530,N_18157,N_17247);
and U21531 (N_21531,N_15324,N_13777);
nor U21532 (N_21532,N_12888,N_16900);
or U21533 (N_21533,N_16757,N_13870);
nor U21534 (N_21534,N_17935,N_16869);
or U21535 (N_21535,N_13834,N_18715);
nor U21536 (N_21536,N_17281,N_13574);
or U21537 (N_21537,N_16740,N_15969);
nor U21538 (N_21538,N_17542,N_17859);
or U21539 (N_21539,N_15768,N_14737);
xnor U21540 (N_21540,N_13774,N_14413);
nor U21541 (N_21541,N_13439,N_17478);
or U21542 (N_21542,N_16404,N_18078);
and U21543 (N_21543,N_18204,N_17392);
nand U21544 (N_21544,N_13013,N_18612);
xnor U21545 (N_21545,N_14981,N_13513);
nor U21546 (N_21546,N_13127,N_17826);
nor U21547 (N_21547,N_15594,N_17784);
nand U21548 (N_21548,N_14363,N_16736);
and U21549 (N_21549,N_14714,N_16717);
nor U21550 (N_21550,N_16973,N_14983);
nand U21551 (N_21551,N_15463,N_16624);
or U21552 (N_21552,N_18267,N_12524);
and U21553 (N_21553,N_13410,N_13185);
and U21554 (N_21554,N_14285,N_15094);
nor U21555 (N_21555,N_17157,N_13003);
xor U21556 (N_21556,N_13583,N_12632);
xnor U21557 (N_21557,N_14480,N_18699);
nor U21558 (N_21558,N_16647,N_17738);
and U21559 (N_21559,N_12794,N_12916);
or U21560 (N_21560,N_17370,N_13029);
and U21561 (N_21561,N_13840,N_15629);
xor U21562 (N_21562,N_15742,N_16385);
nor U21563 (N_21563,N_12634,N_17684);
and U21564 (N_21564,N_17928,N_13216);
nor U21565 (N_21565,N_15798,N_17528);
xor U21566 (N_21566,N_12846,N_14153);
and U21567 (N_21567,N_18280,N_12913);
nor U21568 (N_21568,N_14230,N_17910);
nand U21569 (N_21569,N_12947,N_18580);
and U21570 (N_21570,N_17685,N_14701);
xor U21571 (N_21571,N_17739,N_14565);
xnor U21572 (N_21572,N_18065,N_18292);
or U21573 (N_21573,N_13958,N_17351);
nor U21574 (N_21574,N_17559,N_18159);
nor U21575 (N_21575,N_15131,N_12743);
xor U21576 (N_21576,N_18273,N_18149);
xnor U21577 (N_21577,N_16643,N_14970);
nand U21578 (N_21578,N_15542,N_14475);
nand U21579 (N_21579,N_15431,N_12641);
nand U21580 (N_21580,N_15714,N_14092);
xnor U21581 (N_21581,N_14399,N_16777);
xnor U21582 (N_21582,N_16893,N_16916);
nor U21583 (N_21583,N_18554,N_15944);
nor U21584 (N_21584,N_17345,N_17531);
and U21585 (N_21585,N_14482,N_17811);
nand U21586 (N_21586,N_17224,N_17034);
xor U21587 (N_21587,N_17869,N_15852);
nor U21588 (N_21588,N_14642,N_13231);
xnor U21589 (N_21589,N_13917,N_15939);
and U21590 (N_21590,N_14519,N_17646);
xnor U21591 (N_21591,N_12606,N_14944);
nand U21592 (N_21592,N_17090,N_16716);
and U21593 (N_21593,N_13692,N_16787);
xnor U21594 (N_21594,N_14990,N_14382);
xor U21595 (N_21595,N_17934,N_16282);
nor U21596 (N_21596,N_18490,N_18498);
xor U21597 (N_21597,N_18559,N_14150);
nand U21598 (N_21598,N_14083,N_13214);
and U21599 (N_21599,N_16470,N_14573);
or U21600 (N_21600,N_17432,N_15189);
nor U21601 (N_21601,N_18339,N_18591);
nand U21602 (N_21602,N_13450,N_12515);
nor U21603 (N_21603,N_16515,N_16960);
nor U21604 (N_21604,N_15435,N_17287);
nor U21605 (N_21605,N_13252,N_16969);
xor U21606 (N_21606,N_18252,N_16906);
nor U21607 (N_21607,N_13746,N_12775);
and U21608 (N_21608,N_14027,N_16688);
nand U21609 (N_21609,N_17973,N_12661);
or U21610 (N_21610,N_15941,N_17808);
nand U21611 (N_21611,N_18480,N_18680);
or U21612 (N_21612,N_16457,N_12573);
nand U21613 (N_21613,N_16951,N_13690);
xnor U21614 (N_21614,N_18736,N_18162);
nor U21615 (N_21615,N_12951,N_16342);
nand U21616 (N_21616,N_13298,N_18345);
nand U21617 (N_21617,N_17307,N_15154);
and U21618 (N_21618,N_15475,N_17188);
nor U21619 (N_21619,N_15185,N_14952);
nand U21620 (N_21620,N_18603,N_13913);
nor U21621 (N_21621,N_17517,N_18567);
nor U21622 (N_21622,N_14996,N_18317);
nor U21623 (N_21623,N_16707,N_12935);
xor U21624 (N_21624,N_17636,N_13625);
xnor U21625 (N_21625,N_14822,N_13171);
and U21626 (N_21626,N_12598,N_16340);
and U21627 (N_21627,N_17420,N_13684);
xor U21628 (N_21628,N_13420,N_16392);
nor U21629 (N_21629,N_13953,N_13254);
or U21630 (N_21630,N_17938,N_15763);
nand U21631 (N_21631,N_17121,N_12804);
and U21632 (N_21632,N_18627,N_14569);
and U21633 (N_21633,N_15502,N_16819);
nor U21634 (N_21634,N_15981,N_15424);
and U21635 (N_21635,N_16614,N_14038);
xor U21636 (N_21636,N_13332,N_15961);
nor U21637 (N_21637,N_13400,N_15578);
and U21638 (N_21638,N_12948,N_17473);
or U21639 (N_21639,N_12921,N_14388);
or U21640 (N_21640,N_17680,N_16987);
xor U21641 (N_21641,N_17892,N_15992);
nand U21642 (N_21642,N_13643,N_15150);
nor U21643 (N_21643,N_12782,N_14055);
and U21644 (N_21644,N_14450,N_12857);
or U21645 (N_21645,N_17688,N_12539);
nand U21646 (N_21646,N_14447,N_16531);
xor U21647 (N_21647,N_14478,N_16996);
xor U21648 (N_21648,N_18054,N_14932);
xor U21649 (N_21649,N_15547,N_18057);
nor U21650 (N_21650,N_16527,N_18434);
or U21651 (N_21651,N_13875,N_18210);
nand U21652 (N_21652,N_14188,N_15848);
nor U21653 (N_21653,N_15514,N_18139);
nand U21654 (N_21654,N_16411,N_17533);
and U21655 (N_21655,N_16790,N_17825);
xnor U21656 (N_21656,N_15733,N_16132);
nor U21657 (N_21657,N_18285,N_14501);
or U21658 (N_21658,N_14096,N_14721);
xor U21659 (N_21659,N_14249,N_16593);
xor U21660 (N_21660,N_17981,N_17489);
nand U21661 (N_21661,N_13350,N_16479);
nor U21662 (N_21662,N_14509,N_17612);
xor U21663 (N_21663,N_18297,N_16665);
nor U21664 (N_21664,N_16781,N_16700);
nand U21665 (N_21665,N_12831,N_18517);
nand U21666 (N_21666,N_17519,N_16686);
and U21667 (N_21667,N_14667,N_16043);
nor U21668 (N_21668,N_18284,N_18205);
xnor U21669 (N_21669,N_18049,N_16061);
nor U21670 (N_21670,N_13116,N_13270);
xor U21671 (N_21671,N_13630,N_17787);
and U21672 (N_21672,N_17423,N_17198);
or U21673 (N_21673,N_16823,N_14585);
or U21674 (N_21674,N_12975,N_18311);
or U21675 (N_21675,N_18326,N_16153);
nor U21676 (N_21676,N_17865,N_17091);
and U21677 (N_21677,N_14830,N_17512);
and U21678 (N_21678,N_13502,N_14460);
xnor U21679 (N_21679,N_18659,N_17153);
or U21680 (N_21680,N_18737,N_17511);
xor U21681 (N_21681,N_12977,N_12847);
nand U21682 (N_21682,N_14196,N_12835);
or U21683 (N_21683,N_15266,N_18613);
and U21684 (N_21684,N_17801,N_12908);
xnor U21685 (N_21685,N_18310,N_17520);
and U21686 (N_21686,N_18409,N_14088);
xor U21687 (N_21687,N_12758,N_15371);
xnor U21688 (N_21688,N_15527,N_14041);
nor U21689 (N_21689,N_15414,N_15471);
or U21690 (N_21690,N_15756,N_16743);
or U21691 (N_21691,N_13226,N_14679);
nor U21692 (N_21692,N_15265,N_16496);
nor U21693 (N_21693,N_17990,N_14713);
nand U21694 (N_21694,N_18601,N_18703);
and U21695 (N_21695,N_17380,N_13609);
nand U21696 (N_21696,N_15439,N_15533);
nand U21697 (N_21697,N_17602,N_17154);
nand U21698 (N_21698,N_16019,N_14823);
nand U21699 (N_21699,N_16435,N_17220);
xnor U21700 (N_21700,N_17769,N_18182);
nor U21701 (N_21701,N_13047,N_15389);
xor U21702 (N_21702,N_15788,N_12790);
nand U21703 (N_21703,N_17293,N_14260);
nand U21704 (N_21704,N_15999,N_15897);
and U21705 (N_21705,N_16284,N_17946);
or U21706 (N_21706,N_18347,N_18064);
xor U21707 (N_21707,N_14422,N_16631);
xor U21708 (N_21708,N_17610,N_15726);
nand U21709 (N_21709,N_15380,N_15915);
and U21710 (N_21710,N_12723,N_14974);
and U21711 (N_21711,N_14152,N_12677);
and U21712 (N_21712,N_15073,N_16164);
nand U21713 (N_21713,N_13283,N_14726);
nand U21714 (N_21714,N_15459,N_12714);
nand U21715 (N_21715,N_17952,N_16038);
or U21716 (N_21716,N_14712,N_15576);
or U21717 (N_21717,N_15695,N_17116);
nand U21718 (N_21718,N_17186,N_14880);
xnor U21719 (N_21719,N_13412,N_14633);
or U21720 (N_21720,N_18695,N_16943);
nor U21721 (N_21721,N_15247,N_13515);
or U21722 (N_21722,N_13035,N_18290);
or U21723 (N_21723,N_18585,N_14828);
or U21724 (N_21724,N_16437,N_15815);
xnor U21725 (N_21725,N_13813,N_14950);
or U21726 (N_21726,N_17081,N_16003);
xnor U21727 (N_21727,N_17171,N_15834);
and U21728 (N_21728,N_15061,N_14556);
nand U21729 (N_21729,N_12966,N_13459);
or U21730 (N_21730,N_15536,N_17097);
and U21731 (N_21731,N_13738,N_14171);
nand U21732 (N_21732,N_13766,N_13446);
nor U21733 (N_21733,N_13707,N_14158);
nor U21734 (N_21734,N_13743,N_14978);
xnor U21735 (N_21735,N_15350,N_17375);
and U21736 (N_21736,N_12776,N_15060);
or U21737 (N_21737,N_12644,N_12983);
or U21738 (N_21738,N_15364,N_17292);
or U21739 (N_21739,N_15861,N_18225);
and U21740 (N_21740,N_16645,N_17174);
nand U21741 (N_21741,N_14463,N_17217);
or U21742 (N_21742,N_14602,N_13906);
nor U21743 (N_21743,N_16909,N_17601);
nor U21744 (N_21744,N_13024,N_13011);
xor U21745 (N_21745,N_14240,N_14015);
nor U21746 (N_21746,N_14190,N_15226);
and U21747 (N_21747,N_16490,N_13313);
xor U21748 (N_21748,N_16874,N_12610);
xnor U21749 (N_21749,N_18459,N_17361);
or U21750 (N_21750,N_14871,N_18241);
or U21751 (N_21751,N_16102,N_13356);
or U21752 (N_21752,N_15236,N_17997);
nor U21753 (N_21753,N_18427,N_18621);
or U21754 (N_21754,N_17216,N_14584);
and U21755 (N_21755,N_15979,N_13027);
or U21756 (N_21756,N_17948,N_14673);
and U21757 (N_21757,N_12645,N_13839);
nor U21758 (N_21758,N_17070,N_14739);
or U21759 (N_21759,N_16581,N_17651);
nand U21760 (N_21760,N_14464,N_18370);
nor U21761 (N_21761,N_16629,N_14007);
xnor U21762 (N_21762,N_17377,N_14536);
or U21763 (N_21763,N_14930,N_14834);
and U21764 (N_21764,N_15101,N_14311);
or U21765 (N_21765,N_16780,N_15660);
nand U21766 (N_21766,N_17098,N_16663);
nor U21767 (N_21767,N_18575,N_14675);
and U21768 (N_21768,N_17468,N_17006);
xor U21769 (N_21769,N_14454,N_16738);
nor U21770 (N_21770,N_14206,N_17177);
nor U21771 (N_21771,N_16888,N_14776);
nor U21772 (N_21772,N_16795,N_18156);
and U21773 (N_21773,N_17279,N_17956);
nand U21774 (N_21774,N_18608,N_14636);
or U21775 (N_21775,N_15357,N_16828);
and U21776 (N_21776,N_13154,N_12600);
nand U21777 (N_21777,N_18386,N_17877);
xor U21778 (N_21778,N_17599,N_17158);
and U21779 (N_21779,N_15299,N_17049);
and U21780 (N_21780,N_16503,N_17849);
xor U21781 (N_21781,N_13008,N_17727);
and U21782 (N_21782,N_12934,N_18522);
nor U21783 (N_21783,N_17764,N_14052);
nand U21784 (N_21784,N_13199,N_18023);
nand U21785 (N_21785,N_17898,N_16436);
nor U21786 (N_21786,N_13770,N_16589);
xor U21787 (N_21787,N_16158,N_15264);
nand U21788 (N_21788,N_13042,N_12575);
nor U21789 (N_21789,N_18655,N_15753);
and U21790 (N_21790,N_17848,N_13990);
or U21791 (N_21791,N_12896,N_13622);
and U21792 (N_21792,N_17607,N_13514);
nand U21793 (N_21793,N_17788,N_14660);
or U21794 (N_21794,N_15697,N_16752);
nor U21795 (N_21795,N_14909,N_13988);
and U21796 (N_21796,N_16720,N_15982);
xor U21797 (N_21797,N_18385,N_13867);
nand U21798 (N_21798,N_15759,N_14934);
or U21799 (N_21799,N_18203,N_14492);
xor U21800 (N_21800,N_13940,N_15405);
nand U21801 (N_21801,N_17800,N_17492);
nor U21802 (N_21802,N_17679,N_13596);
xnor U21803 (N_21803,N_16662,N_13326);
nor U21804 (N_21804,N_13619,N_14032);
nor U21805 (N_21805,N_18171,N_12887);
nor U21806 (N_21806,N_18000,N_15270);
and U21807 (N_21807,N_16775,N_15497);
xnor U21808 (N_21808,N_13756,N_16619);
xor U21809 (N_21809,N_13387,N_13153);
nand U21810 (N_21810,N_16400,N_15043);
or U21811 (N_21811,N_15024,N_15208);
nor U21812 (N_21812,N_14486,N_14377);
and U21813 (N_21813,N_14992,N_17051);
nor U21814 (N_21814,N_15651,N_14259);
or U21815 (N_21815,N_16741,N_17535);
and U21816 (N_21816,N_17030,N_18077);
xor U21817 (N_21817,N_17628,N_18491);
or U21818 (N_21818,N_16112,N_15731);
xnor U21819 (N_21819,N_17208,N_17203);
or U21820 (N_21820,N_16409,N_13431);
and U21821 (N_21821,N_17255,N_17655);
nand U21822 (N_21822,N_12698,N_12895);
nor U21823 (N_21823,N_17454,N_13221);
and U21824 (N_21824,N_16595,N_16567);
nand U21825 (N_21825,N_17521,N_13561);
nor U21826 (N_21826,N_17998,N_16251);
xnor U21827 (N_21827,N_13235,N_18581);
nor U21828 (N_21828,N_18387,N_14250);
or U21829 (N_21829,N_17507,N_13901);
xnor U21830 (N_21830,N_15246,N_14404);
or U21831 (N_21831,N_18693,N_14757);
and U21832 (N_21832,N_12579,N_13964);
xor U21833 (N_21833,N_12912,N_13848);
nand U21834 (N_21834,N_16130,N_12969);
nand U21835 (N_21835,N_18115,N_17167);
or U21836 (N_21836,N_13238,N_16209);
and U21837 (N_21837,N_17445,N_15065);
or U21838 (N_21838,N_13291,N_16074);
and U21839 (N_21839,N_13611,N_13689);
nor U21840 (N_21840,N_12747,N_15455);
and U21841 (N_21841,N_15018,N_17901);
xor U21842 (N_21842,N_17916,N_16766);
nand U21843 (N_21843,N_13351,N_18111);
xor U21844 (N_21844,N_12783,N_13564);
xnor U21845 (N_21845,N_15447,N_18334);
xnor U21846 (N_21846,N_16618,N_18072);
xnor U21847 (N_21847,N_15825,N_14493);
or U21848 (N_21848,N_16955,N_17228);
nor U21849 (N_21849,N_15409,N_18277);
xnor U21850 (N_21850,N_17016,N_15505);
xor U21851 (N_21851,N_16718,N_15383);
nand U21852 (N_21852,N_12740,N_16811);
nand U21853 (N_21853,N_18708,N_16269);
or U21854 (N_21854,N_16516,N_13861);
nand U21855 (N_21855,N_13610,N_14995);
and U21856 (N_21856,N_14601,N_17966);
or U21857 (N_21857,N_13850,N_16895);
nand U21858 (N_21858,N_14680,N_13529);
nand U21859 (N_21859,N_16681,N_17267);
xnor U21860 (N_21860,N_16862,N_18129);
nor U21861 (N_21861,N_15344,N_18588);
and U21862 (N_21862,N_14968,N_17332);
nand U21863 (N_21863,N_16147,N_18135);
nor U21864 (N_21864,N_15283,N_14004);
nand U21865 (N_21865,N_17422,N_17060);
and U21866 (N_21866,N_13745,N_16330);
nor U21867 (N_21867,N_14883,N_18523);
xnor U21868 (N_21868,N_15030,N_18288);
xor U21869 (N_21869,N_14506,N_14331);
or U21870 (N_21870,N_15278,N_12607);
and U21871 (N_21871,N_17534,N_17214);
nand U21872 (N_21872,N_14054,N_16227);
and U21873 (N_21873,N_16870,N_13248);
or U21874 (N_21874,N_14893,N_14781);
nand U21875 (N_21875,N_16157,N_16048);
nand U21876 (N_21876,N_13299,N_12802);
or U21877 (N_21877,N_14173,N_16594);
xor U21878 (N_21878,N_14096,N_13669);
xnor U21879 (N_21879,N_15265,N_15511);
nor U21880 (N_21880,N_15459,N_18100);
nand U21881 (N_21881,N_13255,N_17884);
and U21882 (N_21882,N_17768,N_15449);
nand U21883 (N_21883,N_13764,N_12864);
nor U21884 (N_21884,N_14911,N_16932);
xor U21885 (N_21885,N_14121,N_18185);
and U21886 (N_21886,N_13501,N_17311);
nand U21887 (N_21887,N_14793,N_13131);
nand U21888 (N_21888,N_15768,N_15487);
nand U21889 (N_21889,N_17263,N_16170);
nand U21890 (N_21890,N_17879,N_16506);
and U21891 (N_21891,N_13320,N_14346);
nor U21892 (N_21892,N_17188,N_15133);
nor U21893 (N_21893,N_15620,N_18670);
and U21894 (N_21894,N_17085,N_16435);
and U21895 (N_21895,N_16755,N_16658);
nor U21896 (N_21896,N_18548,N_16119);
xor U21897 (N_21897,N_16194,N_15661);
nand U21898 (N_21898,N_12520,N_17544);
or U21899 (N_21899,N_17553,N_18673);
nor U21900 (N_21900,N_14788,N_18141);
or U21901 (N_21901,N_14035,N_15254);
xnor U21902 (N_21902,N_17099,N_18729);
nand U21903 (N_21903,N_12716,N_15267);
or U21904 (N_21904,N_13232,N_13480);
and U21905 (N_21905,N_18544,N_13859);
nand U21906 (N_21906,N_13952,N_12594);
xnor U21907 (N_21907,N_12858,N_15273);
nand U21908 (N_21908,N_14542,N_16145);
nand U21909 (N_21909,N_15437,N_15315);
and U21910 (N_21910,N_15911,N_17853);
xor U21911 (N_21911,N_18001,N_17768);
and U21912 (N_21912,N_14794,N_16173);
or U21913 (N_21913,N_13255,N_17204);
xor U21914 (N_21914,N_13055,N_16923);
and U21915 (N_21915,N_13804,N_13289);
nand U21916 (N_21916,N_13762,N_13564);
and U21917 (N_21917,N_14645,N_16395);
or U21918 (N_21918,N_14408,N_16090);
nand U21919 (N_21919,N_12525,N_17982);
or U21920 (N_21920,N_16839,N_12626);
or U21921 (N_21921,N_17082,N_16070);
nor U21922 (N_21922,N_16109,N_15291);
nand U21923 (N_21923,N_18409,N_14510);
nand U21924 (N_21924,N_13347,N_18471);
nand U21925 (N_21925,N_17839,N_14516);
xnor U21926 (N_21926,N_13087,N_18267);
or U21927 (N_21927,N_18061,N_16230);
xnor U21928 (N_21928,N_18577,N_16301);
nand U21929 (N_21929,N_12978,N_14651);
nor U21930 (N_21930,N_13021,N_18124);
nor U21931 (N_21931,N_14754,N_15725);
or U21932 (N_21932,N_18139,N_16300);
or U21933 (N_21933,N_17435,N_17886);
nor U21934 (N_21934,N_18080,N_15552);
or U21935 (N_21935,N_13642,N_13427);
xor U21936 (N_21936,N_18553,N_17996);
nand U21937 (N_21937,N_16257,N_13007);
and U21938 (N_21938,N_16553,N_16983);
and U21939 (N_21939,N_16337,N_16100);
nand U21940 (N_21940,N_16679,N_13874);
nand U21941 (N_21941,N_15725,N_13487);
nand U21942 (N_21942,N_15099,N_18315);
and U21943 (N_21943,N_18092,N_13620);
or U21944 (N_21944,N_17156,N_12955);
or U21945 (N_21945,N_18723,N_13494);
nand U21946 (N_21946,N_17362,N_18509);
nand U21947 (N_21947,N_17466,N_14852);
nand U21948 (N_21948,N_17410,N_12711);
nand U21949 (N_21949,N_14366,N_16118);
nor U21950 (N_21950,N_16255,N_15687);
or U21951 (N_21951,N_16849,N_14467);
xor U21952 (N_21952,N_18663,N_13598);
nor U21953 (N_21953,N_13695,N_16635);
or U21954 (N_21954,N_13318,N_18130);
and U21955 (N_21955,N_14192,N_18125);
and U21956 (N_21956,N_15310,N_16566);
xor U21957 (N_21957,N_14301,N_16488);
nor U21958 (N_21958,N_18419,N_13752);
nor U21959 (N_21959,N_13085,N_13791);
nand U21960 (N_21960,N_15459,N_17251);
xnor U21961 (N_21961,N_14031,N_16621);
xor U21962 (N_21962,N_17532,N_15469);
nor U21963 (N_21963,N_13988,N_12935);
xor U21964 (N_21964,N_17213,N_12951);
and U21965 (N_21965,N_15617,N_14485);
and U21966 (N_21966,N_13340,N_16233);
or U21967 (N_21967,N_12586,N_16007);
or U21968 (N_21968,N_14415,N_14994);
nor U21969 (N_21969,N_15499,N_17501);
and U21970 (N_21970,N_14299,N_13007);
and U21971 (N_21971,N_16315,N_15830);
or U21972 (N_21972,N_17963,N_17489);
and U21973 (N_21973,N_17669,N_14072);
xor U21974 (N_21974,N_15409,N_16213);
or U21975 (N_21975,N_12767,N_17527);
xnor U21976 (N_21976,N_17038,N_16223);
nand U21977 (N_21977,N_17186,N_15201);
xor U21978 (N_21978,N_17633,N_16277);
or U21979 (N_21979,N_14256,N_15004);
and U21980 (N_21980,N_13479,N_16622);
nor U21981 (N_21981,N_15211,N_15494);
or U21982 (N_21982,N_14764,N_14129);
xnor U21983 (N_21983,N_14815,N_18204);
nor U21984 (N_21984,N_14948,N_12591);
nand U21985 (N_21985,N_17954,N_14453);
xnor U21986 (N_21986,N_12568,N_13194);
nor U21987 (N_21987,N_15080,N_14364);
and U21988 (N_21988,N_15546,N_13253);
or U21989 (N_21989,N_14361,N_12935);
xor U21990 (N_21990,N_18014,N_14893);
xnor U21991 (N_21991,N_18161,N_14537);
and U21992 (N_21992,N_13444,N_18152);
nor U21993 (N_21993,N_17041,N_14670);
nand U21994 (N_21994,N_15099,N_15854);
or U21995 (N_21995,N_15825,N_15736);
or U21996 (N_21996,N_17142,N_12995);
xor U21997 (N_21997,N_17378,N_17548);
nand U21998 (N_21998,N_13305,N_12528);
and U21999 (N_21999,N_16887,N_16435);
and U22000 (N_22000,N_13495,N_13930);
nor U22001 (N_22001,N_15649,N_14008);
nand U22002 (N_22002,N_16368,N_16799);
and U22003 (N_22003,N_16075,N_18145);
nor U22004 (N_22004,N_17760,N_17865);
and U22005 (N_22005,N_13376,N_14274);
nand U22006 (N_22006,N_15771,N_17301);
xor U22007 (N_22007,N_17399,N_17971);
or U22008 (N_22008,N_17564,N_13398);
or U22009 (N_22009,N_13102,N_18741);
or U22010 (N_22010,N_16748,N_14889);
nand U22011 (N_22011,N_14151,N_15199);
nor U22012 (N_22012,N_18456,N_12675);
nand U22013 (N_22013,N_17827,N_15125);
xor U22014 (N_22014,N_12567,N_16804);
nor U22015 (N_22015,N_18049,N_13628);
or U22016 (N_22016,N_18709,N_18139);
nor U22017 (N_22017,N_18252,N_13054);
xor U22018 (N_22018,N_16675,N_17379);
and U22019 (N_22019,N_12811,N_14508);
and U22020 (N_22020,N_15835,N_15946);
and U22021 (N_22021,N_17413,N_17326);
or U22022 (N_22022,N_15332,N_16280);
or U22023 (N_22023,N_15545,N_14198);
and U22024 (N_22024,N_14183,N_16248);
or U22025 (N_22025,N_14392,N_18594);
and U22026 (N_22026,N_13732,N_12936);
nand U22027 (N_22027,N_12871,N_16165);
xnor U22028 (N_22028,N_13163,N_12955);
and U22029 (N_22029,N_17025,N_17001);
or U22030 (N_22030,N_13688,N_14069);
xnor U22031 (N_22031,N_16449,N_14748);
or U22032 (N_22032,N_17169,N_12987);
nor U22033 (N_22033,N_14742,N_15971);
nor U22034 (N_22034,N_17588,N_14451);
nand U22035 (N_22035,N_14205,N_17942);
and U22036 (N_22036,N_17389,N_12921);
nand U22037 (N_22037,N_15741,N_16057);
nor U22038 (N_22038,N_15554,N_18016);
nand U22039 (N_22039,N_14621,N_14100);
nor U22040 (N_22040,N_13662,N_15409);
nand U22041 (N_22041,N_15667,N_13425);
nand U22042 (N_22042,N_13728,N_14142);
nand U22043 (N_22043,N_17689,N_16547);
nor U22044 (N_22044,N_18256,N_13078);
or U22045 (N_22045,N_17708,N_18110);
xnor U22046 (N_22046,N_16338,N_13207);
and U22047 (N_22047,N_13943,N_16981);
nor U22048 (N_22048,N_12717,N_12946);
xnor U22049 (N_22049,N_14830,N_17521);
and U22050 (N_22050,N_14022,N_18478);
or U22051 (N_22051,N_15061,N_12987);
nand U22052 (N_22052,N_13765,N_16784);
and U22053 (N_22053,N_14398,N_18061);
nor U22054 (N_22054,N_15875,N_18265);
xor U22055 (N_22055,N_17097,N_13701);
nor U22056 (N_22056,N_15195,N_14831);
xor U22057 (N_22057,N_18227,N_12730);
nand U22058 (N_22058,N_15623,N_14966);
xor U22059 (N_22059,N_14561,N_12570);
nor U22060 (N_22060,N_15032,N_17470);
and U22061 (N_22061,N_18360,N_15258);
and U22062 (N_22062,N_15452,N_13919);
xor U22063 (N_22063,N_14902,N_14051);
nor U22064 (N_22064,N_15550,N_16258);
nand U22065 (N_22065,N_18174,N_18095);
and U22066 (N_22066,N_14121,N_14378);
xor U22067 (N_22067,N_15881,N_12877);
xnor U22068 (N_22068,N_18054,N_15224);
nand U22069 (N_22069,N_15632,N_12634);
nor U22070 (N_22070,N_15649,N_12502);
or U22071 (N_22071,N_16000,N_14525);
xor U22072 (N_22072,N_14436,N_15350);
nor U22073 (N_22073,N_14717,N_17507);
and U22074 (N_22074,N_15176,N_18576);
xor U22075 (N_22075,N_14233,N_13405);
nand U22076 (N_22076,N_14881,N_17497);
or U22077 (N_22077,N_18056,N_18290);
nor U22078 (N_22078,N_13961,N_18505);
or U22079 (N_22079,N_17922,N_16376);
nor U22080 (N_22080,N_15008,N_12521);
nand U22081 (N_22081,N_15466,N_15564);
or U22082 (N_22082,N_13053,N_13848);
nor U22083 (N_22083,N_14454,N_16576);
nand U22084 (N_22084,N_14948,N_15997);
nor U22085 (N_22085,N_16641,N_13498);
nand U22086 (N_22086,N_16824,N_15224);
nor U22087 (N_22087,N_13763,N_15485);
nor U22088 (N_22088,N_15816,N_14885);
nor U22089 (N_22089,N_18039,N_17823);
nand U22090 (N_22090,N_13123,N_15611);
nor U22091 (N_22091,N_14515,N_15617);
nor U22092 (N_22092,N_14533,N_13087);
nand U22093 (N_22093,N_14711,N_15459);
xnor U22094 (N_22094,N_14372,N_16948);
and U22095 (N_22095,N_15196,N_16614);
or U22096 (N_22096,N_18530,N_17868);
and U22097 (N_22097,N_18553,N_13475);
and U22098 (N_22098,N_15326,N_13887);
nand U22099 (N_22099,N_12660,N_14469);
nand U22100 (N_22100,N_12726,N_12853);
and U22101 (N_22101,N_14322,N_15248);
or U22102 (N_22102,N_12699,N_14859);
nand U22103 (N_22103,N_13251,N_12888);
xor U22104 (N_22104,N_17910,N_15196);
xor U22105 (N_22105,N_15269,N_13312);
nor U22106 (N_22106,N_14309,N_16556);
xnor U22107 (N_22107,N_14107,N_15452);
and U22108 (N_22108,N_17620,N_14256);
xnor U22109 (N_22109,N_17327,N_18587);
nor U22110 (N_22110,N_17331,N_13246);
nor U22111 (N_22111,N_12730,N_14479);
nor U22112 (N_22112,N_17895,N_15427);
nand U22113 (N_22113,N_15698,N_17925);
xnor U22114 (N_22114,N_13649,N_16633);
xor U22115 (N_22115,N_18233,N_16484);
or U22116 (N_22116,N_17666,N_17862);
and U22117 (N_22117,N_13344,N_16362);
xnor U22118 (N_22118,N_14250,N_17474);
or U22119 (N_22119,N_13450,N_14875);
and U22120 (N_22120,N_18357,N_14362);
xnor U22121 (N_22121,N_16607,N_14696);
or U22122 (N_22122,N_14059,N_15791);
or U22123 (N_22123,N_13547,N_13495);
and U22124 (N_22124,N_17422,N_13819);
or U22125 (N_22125,N_14492,N_15692);
nand U22126 (N_22126,N_14051,N_13612);
or U22127 (N_22127,N_17125,N_12662);
nand U22128 (N_22128,N_17568,N_15560);
and U22129 (N_22129,N_16125,N_16419);
nand U22130 (N_22130,N_18476,N_18543);
xor U22131 (N_22131,N_16765,N_12664);
nand U22132 (N_22132,N_13074,N_16689);
nor U22133 (N_22133,N_16410,N_12679);
nor U22134 (N_22134,N_15936,N_16609);
nand U22135 (N_22135,N_16881,N_15153);
nor U22136 (N_22136,N_17427,N_16129);
nor U22137 (N_22137,N_13994,N_15914);
xnor U22138 (N_22138,N_18156,N_16030);
nor U22139 (N_22139,N_13683,N_16284);
and U22140 (N_22140,N_16926,N_18053);
nand U22141 (N_22141,N_12990,N_18343);
and U22142 (N_22142,N_16166,N_15747);
xnor U22143 (N_22143,N_16679,N_15206);
or U22144 (N_22144,N_15858,N_14149);
nand U22145 (N_22145,N_16097,N_14916);
or U22146 (N_22146,N_12824,N_14597);
or U22147 (N_22147,N_18008,N_15144);
nand U22148 (N_22148,N_18050,N_14561);
and U22149 (N_22149,N_12579,N_12620);
and U22150 (N_22150,N_13021,N_16430);
xor U22151 (N_22151,N_14145,N_15717);
xnor U22152 (N_22152,N_15857,N_17533);
nor U22153 (N_22153,N_18050,N_18027);
and U22154 (N_22154,N_17963,N_12804);
and U22155 (N_22155,N_16448,N_18073);
nand U22156 (N_22156,N_14248,N_12788);
nor U22157 (N_22157,N_18632,N_15142);
nand U22158 (N_22158,N_18195,N_17143);
and U22159 (N_22159,N_15832,N_12683);
nand U22160 (N_22160,N_16460,N_13130);
nand U22161 (N_22161,N_13706,N_18608);
and U22162 (N_22162,N_17633,N_15357);
nor U22163 (N_22163,N_13899,N_15821);
nor U22164 (N_22164,N_16046,N_12759);
nor U22165 (N_22165,N_18077,N_17097);
nor U22166 (N_22166,N_13596,N_18083);
xor U22167 (N_22167,N_15243,N_16416);
or U22168 (N_22168,N_16628,N_17017);
nor U22169 (N_22169,N_16575,N_14954);
and U22170 (N_22170,N_15180,N_17362);
nor U22171 (N_22171,N_18311,N_14646);
nor U22172 (N_22172,N_17563,N_14053);
or U22173 (N_22173,N_14714,N_12606);
xnor U22174 (N_22174,N_18288,N_17614);
nand U22175 (N_22175,N_16011,N_18328);
nand U22176 (N_22176,N_13348,N_13742);
nand U22177 (N_22177,N_17938,N_13560);
and U22178 (N_22178,N_17098,N_18155);
and U22179 (N_22179,N_13690,N_16958);
and U22180 (N_22180,N_17896,N_15941);
nor U22181 (N_22181,N_15888,N_17543);
or U22182 (N_22182,N_15006,N_14966);
and U22183 (N_22183,N_14131,N_14628);
xnor U22184 (N_22184,N_18283,N_16658);
nand U22185 (N_22185,N_18438,N_17436);
nand U22186 (N_22186,N_17317,N_14182);
and U22187 (N_22187,N_16102,N_16457);
nand U22188 (N_22188,N_13205,N_18008);
or U22189 (N_22189,N_13342,N_16713);
or U22190 (N_22190,N_18280,N_17718);
and U22191 (N_22191,N_18318,N_15330);
or U22192 (N_22192,N_12813,N_13502);
nand U22193 (N_22193,N_16106,N_12840);
and U22194 (N_22194,N_13186,N_16969);
or U22195 (N_22195,N_12899,N_18601);
and U22196 (N_22196,N_12669,N_16777);
nor U22197 (N_22197,N_14499,N_17330);
and U22198 (N_22198,N_14792,N_18328);
nand U22199 (N_22199,N_13778,N_16440);
nor U22200 (N_22200,N_14649,N_14969);
and U22201 (N_22201,N_14074,N_13734);
or U22202 (N_22202,N_14148,N_16076);
and U22203 (N_22203,N_15595,N_17666);
or U22204 (N_22204,N_16875,N_17461);
xnor U22205 (N_22205,N_16212,N_17193);
nand U22206 (N_22206,N_16078,N_14371);
nor U22207 (N_22207,N_14510,N_16138);
xor U22208 (N_22208,N_16728,N_13065);
nor U22209 (N_22209,N_17096,N_18121);
or U22210 (N_22210,N_13269,N_18046);
nand U22211 (N_22211,N_13077,N_14699);
xor U22212 (N_22212,N_14079,N_15313);
nor U22213 (N_22213,N_17924,N_17262);
or U22214 (N_22214,N_13261,N_16266);
nor U22215 (N_22215,N_15003,N_15433);
and U22216 (N_22216,N_15291,N_14851);
nand U22217 (N_22217,N_14636,N_15736);
nor U22218 (N_22218,N_14642,N_15851);
and U22219 (N_22219,N_15349,N_17062);
nor U22220 (N_22220,N_14542,N_12739);
nand U22221 (N_22221,N_15277,N_17684);
nand U22222 (N_22222,N_13883,N_12862);
nand U22223 (N_22223,N_14287,N_15313);
or U22224 (N_22224,N_17165,N_17182);
nand U22225 (N_22225,N_13971,N_18724);
nor U22226 (N_22226,N_13067,N_14489);
and U22227 (N_22227,N_17160,N_16936);
nand U22228 (N_22228,N_18077,N_15796);
and U22229 (N_22229,N_16099,N_18329);
nor U22230 (N_22230,N_17302,N_14029);
and U22231 (N_22231,N_14109,N_15169);
or U22232 (N_22232,N_13289,N_17204);
and U22233 (N_22233,N_18123,N_14978);
and U22234 (N_22234,N_18746,N_14647);
or U22235 (N_22235,N_15438,N_16772);
xnor U22236 (N_22236,N_14354,N_13738);
nand U22237 (N_22237,N_13532,N_17619);
xnor U22238 (N_22238,N_15183,N_17120);
or U22239 (N_22239,N_15321,N_13373);
or U22240 (N_22240,N_17450,N_17070);
nor U22241 (N_22241,N_13806,N_17219);
nand U22242 (N_22242,N_12753,N_15781);
nor U22243 (N_22243,N_16650,N_14769);
or U22244 (N_22244,N_14827,N_16274);
nand U22245 (N_22245,N_17071,N_13768);
nand U22246 (N_22246,N_15568,N_13302);
and U22247 (N_22247,N_13250,N_16581);
nor U22248 (N_22248,N_17966,N_15594);
or U22249 (N_22249,N_15855,N_16122);
or U22250 (N_22250,N_17309,N_18064);
xnor U22251 (N_22251,N_14400,N_15370);
or U22252 (N_22252,N_16229,N_14165);
or U22253 (N_22253,N_15843,N_18301);
nand U22254 (N_22254,N_15120,N_13017);
or U22255 (N_22255,N_14895,N_15353);
xnor U22256 (N_22256,N_14004,N_15008);
or U22257 (N_22257,N_18573,N_18109);
and U22258 (N_22258,N_15247,N_16263);
or U22259 (N_22259,N_14410,N_15967);
xnor U22260 (N_22260,N_16418,N_14034);
xor U22261 (N_22261,N_14124,N_16608);
or U22262 (N_22262,N_17757,N_17699);
xnor U22263 (N_22263,N_14565,N_16205);
or U22264 (N_22264,N_14034,N_12996);
nand U22265 (N_22265,N_16245,N_14862);
xnor U22266 (N_22266,N_17400,N_17448);
or U22267 (N_22267,N_15894,N_16305);
nor U22268 (N_22268,N_14679,N_18656);
and U22269 (N_22269,N_13286,N_14923);
or U22270 (N_22270,N_14662,N_18522);
or U22271 (N_22271,N_18561,N_18424);
nor U22272 (N_22272,N_12945,N_17229);
nand U22273 (N_22273,N_14183,N_18558);
nand U22274 (N_22274,N_18317,N_17185);
xnor U22275 (N_22275,N_12864,N_14327);
nor U22276 (N_22276,N_17467,N_14334);
or U22277 (N_22277,N_17902,N_16502);
nor U22278 (N_22278,N_16551,N_15792);
or U22279 (N_22279,N_13010,N_15173);
nand U22280 (N_22280,N_16788,N_17054);
nor U22281 (N_22281,N_15167,N_13185);
and U22282 (N_22282,N_18333,N_13428);
nand U22283 (N_22283,N_15012,N_13752);
or U22284 (N_22284,N_17967,N_13163);
or U22285 (N_22285,N_13120,N_17037);
and U22286 (N_22286,N_16581,N_13519);
nand U22287 (N_22287,N_17218,N_12901);
xnor U22288 (N_22288,N_18122,N_13327);
nand U22289 (N_22289,N_15876,N_13285);
xor U22290 (N_22290,N_14210,N_15759);
and U22291 (N_22291,N_13612,N_18074);
nand U22292 (N_22292,N_16926,N_13301);
nor U22293 (N_22293,N_13986,N_17503);
or U22294 (N_22294,N_16273,N_17939);
or U22295 (N_22295,N_13635,N_16322);
and U22296 (N_22296,N_13517,N_18480);
nand U22297 (N_22297,N_13047,N_16176);
nand U22298 (N_22298,N_18690,N_16496);
or U22299 (N_22299,N_13580,N_15409);
or U22300 (N_22300,N_17631,N_17137);
xnor U22301 (N_22301,N_13067,N_12681);
nor U22302 (N_22302,N_17303,N_13580);
xor U22303 (N_22303,N_17797,N_17440);
xnor U22304 (N_22304,N_13560,N_14750);
and U22305 (N_22305,N_14706,N_16178);
xnor U22306 (N_22306,N_17437,N_15510);
nand U22307 (N_22307,N_14632,N_15251);
xnor U22308 (N_22308,N_17901,N_16884);
xor U22309 (N_22309,N_13405,N_14494);
nand U22310 (N_22310,N_17655,N_14688);
and U22311 (N_22311,N_17752,N_16378);
nand U22312 (N_22312,N_18419,N_13635);
nand U22313 (N_22313,N_12626,N_18652);
and U22314 (N_22314,N_13239,N_12569);
nor U22315 (N_22315,N_16989,N_15418);
nand U22316 (N_22316,N_14313,N_13696);
and U22317 (N_22317,N_17170,N_14038);
or U22318 (N_22318,N_13354,N_18040);
or U22319 (N_22319,N_16877,N_16454);
nand U22320 (N_22320,N_13253,N_16158);
or U22321 (N_22321,N_18389,N_14634);
or U22322 (N_22322,N_15685,N_16303);
nor U22323 (N_22323,N_17516,N_18475);
or U22324 (N_22324,N_12980,N_18531);
and U22325 (N_22325,N_17592,N_13553);
and U22326 (N_22326,N_18213,N_13604);
xnor U22327 (N_22327,N_13720,N_16208);
or U22328 (N_22328,N_16228,N_17432);
nor U22329 (N_22329,N_18667,N_17525);
nor U22330 (N_22330,N_13767,N_17050);
xor U22331 (N_22331,N_18282,N_12640);
xor U22332 (N_22332,N_16438,N_12721);
xor U22333 (N_22333,N_15156,N_13470);
or U22334 (N_22334,N_17143,N_17792);
nor U22335 (N_22335,N_14428,N_14408);
and U22336 (N_22336,N_15862,N_16686);
and U22337 (N_22337,N_14047,N_14889);
nand U22338 (N_22338,N_14392,N_13209);
xnor U22339 (N_22339,N_16237,N_13642);
and U22340 (N_22340,N_16375,N_15581);
or U22341 (N_22341,N_16519,N_17815);
and U22342 (N_22342,N_16353,N_17412);
and U22343 (N_22343,N_18483,N_16679);
xnor U22344 (N_22344,N_12646,N_12701);
xnor U22345 (N_22345,N_15913,N_16946);
and U22346 (N_22346,N_17902,N_16151);
and U22347 (N_22347,N_17897,N_14914);
nor U22348 (N_22348,N_15185,N_14030);
nor U22349 (N_22349,N_14998,N_13136);
or U22350 (N_22350,N_18617,N_16757);
or U22351 (N_22351,N_15008,N_18140);
xnor U22352 (N_22352,N_13205,N_13773);
xor U22353 (N_22353,N_13063,N_13361);
xnor U22354 (N_22354,N_17394,N_15556);
xor U22355 (N_22355,N_14020,N_18276);
or U22356 (N_22356,N_15861,N_18578);
nand U22357 (N_22357,N_16699,N_14312);
nand U22358 (N_22358,N_16774,N_18128);
nor U22359 (N_22359,N_14793,N_17723);
xor U22360 (N_22360,N_14492,N_18097);
and U22361 (N_22361,N_14653,N_12730);
or U22362 (N_22362,N_17141,N_18208);
nor U22363 (N_22363,N_15112,N_16467);
or U22364 (N_22364,N_14123,N_16283);
xor U22365 (N_22365,N_12800,N_14309);
nand U22366 (N_22366,N_12770,N_12948);
nand U22367 (N_22367,N_14675,N_13880);
nand U22368 (N_22368,N_15505,N_14342);
nand U22369 (N_22369,N_12549,N_14764);
xor U22370 (N_22370,N_17051,N_14410);
nand U22371 (N_22371,N_13520,N_12563);
nand U22372 (N_22372,N_13795,N_18285);
nor U22373 (N_22373,N_14605,N_18260);
nor U22374 (N_22374,N_16072,N_18416);
nor U22375 (N_22375,N_17489,N_17888);
and U22376 (N_22376,N_14473,N_13246);
and U22377 (N_22377,N_14085,N_18203);
nor U22378 (N_22378,N_15472,N_18511);
nor U22379 (N_22379,N_17242,N_13057);
nand U22380 (N_22380,N_12707,N_15816);
nand U22381 (N_22381,N_15164,N_15406);
xor U22382 (N_22382,N_17072,N_16801);
xor U22383 (N_22383,N_18273,N_17972);
nor U22384 (N_22384,N_18267,N_15539);
nor U22385 (N_22385,N_16377,N_12965);
nand U22386 (N_22386,N_15044,N_18656);
or U22387 (N_22387,N_17947,N_13115);
or U22388 (N_22388,N_15964,N_16608);
or U22389 (N_22389,N_17054,N_17766);
nand U22390 (N_22390,N_16616,N_18533);
and U22391 (N_22391,N_17591,N_15610);
xnor U22392 (N_22392,N_16512,N_17262);
or U22393 (N_22393,N_17461,N_14267);
or U22394 (N_22394,N_15835,N_12656);
nand U22395 (N_22395,N_16533,N_13446);
or U22396 (N_22396,N_17173,N_18243);
or U22397 (N_22397,N_16208,N_13341);
or U22398 (N_22398,N_14887,N_17770);
and U22399 (N_22399,N_17465,N_14366);
nand U22400 (N_22400,N_14976,N_15752);
or U22401 (N_22401,N_16505,N_14088);
and U22402 (N_22402,N_17729,N_13365);
nor U22403 (N_22403,N_13577,N_16986);
and U22404 (N_22404,N_17176,N_17860);
xor U22405 (N_22405,N_16006,N_16619);
xnor U22406 (N_22406,N_17660,N_16744);
or U22407 (N_22407,N_13871,N_17118);
and U22408 (N_22408,N_15313,N_13020);
xor U22409 (N_22409,N_15099,N_16211);
xnor U22410 (N_22410,N_15923,N_17289);
nand U22411 (N_22411,N_15340,N_17350);
and U22412 (N_22412,N_16605,N_13605);
nor U22413 (N_22413,N_13786,N_14775);
or U22414 (N_22414,N_17227,N_18038);
xor U22415 (N_22415,N_13852,N_17710);
and U22416 (N_22416,N_17985,N_12593);
and U22417 (N_22417,N_15124,N_14692);
or U22418 (N_22418,N_17615,N_15356);
and U22419 (N_22419,N_17593,N_18241);
nand U22420 (N_22420,N_16033,N_16752);
nor U22421 (N_22421,N_13135,N_13985);
nand U22422 (N_22422,N_16027,N_16660);
and U22423 (N_22423,N_13138,N_18234);
xor U22424 (N_22424,N_12900,N_15823);
xor U22425 (N_22425,N_13933,N_12512);
xor U22426 (N_22426,N_14233,N_15058);
nor U22427 (N_22427,N_12539,N_13308);
nand U22428 (N_22428,N_16284,N_13095);
and U22429 (N_22429,N_17558,N_17272);
and U22430 (N_22430,N_14067,N_18014);
nand U22431 (N_22431,N_13800,N_15792);
and U22432 (N_22432,N_13680,N_16675);
xnor U22433 (N_22433,N_18274,N_13066);
and U22434 (N_22434,N_13360,N_14900);
or U22435 (N_22435,N_16629,N_14335);
and U22436 (N_22436,N_17703,N_16768);
nand U22437 (N_22437,N_16062,N_13878);
nand U22438 (N_22438,N_18308,N_17368);
or U22439 (N_22439,N_15928,N_16745);
xor U22440 (N_22440,N_13771,N_16305);
nand U22441 (N_22441,N_14802,N_16097);
xnor U22442 (N_22442,N_15747,N_13631);
and U22443 (N_22443,N_14926,N_15490);
nor U22444 (N_22444,N_16502,N_14647);
xnor U22445 (N_22445,N_15965,N_14460);
xor U22446 (N_22446,N_16419,N_16849);
or U22447 (N_22447,N_17186,N_13558);
nand U22448 (N_22448,N_16549,N_17334);
or U22449 (N_22449,N_14331,N_14522);
xor U22450 (N_22450,N_13831,N_14440);
xnor U22451 (N_22451,N_17817,N_12786);
nand U22452 (N_22452,N_16997,N_16786);
nor U22453 (N_22453,N_14668,N_16555);
nor U22454 (N_22454,N_13204,N_18535);
and U22455 (N_22455,N_18620,N_17445);
nor U22456 (N_22456,N_17501,N_13993);
or U22457 (N_22457,N_17130,N_16273);
and U22458 (N_22458,N_15702,N_18265);
xor U22459 (N_22459,N_16947,N_17188);
xnor U22460 (N_22460,N_13393,N_16843);
or U22461 (N_22461,N_13702,N_13760);
nor U22462 (N_22462,N_16337,N_16408);
or U22463 (N_22463,N_14870,N_18348);
nor U22464 (N_22464,N_13350,N_17419);
nor U22465 (N_22465,N_18243,N_17863);
and U22466 (N_22466,N_13652,N_14843);
xor U22467 (N_22467,N_15755,N_13884);
nand U22468 (N_22468,N_14690,N_13026);
xor U22469 (N_22469,N_16503,N_14128);
nand U22470 (N_22470,N_15255,N_13075);
xor U22471 (N_22471,N_17495,N_13075);
nand U22472 (N_22472,N_12574,N_16801);
and U22473 (N_22473,N_15266,N_17324);
xnor U22474 (N_22474,N_16854,N_15789);
nand U22475 (N_22475,N_17552,N_18369);
and U22476 (N_22476,N_16774,N_15254);
xnor U22477 (N_22477,N_18028,N_15587);
nor U22478 (N_22478,N_18720,N_17384);
nand U22479 (N_22479,N_16165,N_18370);
or U22480 (N_22480,N_18706,N_17977);
or U22481 (N_22481,N_18340,N_16816);
xnor U22482 (N_22482,N_12666,N_15734);
and U22483 (N_22483,N_17492,N_16350);
xnor U22484 (N_22484,N_14884,N_16380);
and U22485 (N_22485,N_15144,N_14448);
xor U22486 (N_22486,N_17543,N_13397);
xor U22487 (N_22487,N_14687,N_17913);
nand U22488 (N_22488,N_14311,N_14773);
nand U22489 (N_22489,N_17844,N_12780);
nand U22490 (N_22490,N_16294,N_16237);
nor U22491 (N_22491,N_14186,N_17489);
and U22492 (N_22492,N_16115,N_13888);
or U22493 (N_22493,N_18567,N_15013);
nand U22494 (N_22494,N_15306,N_16398);
nor U22495 (N_22495,N_15639,N_14069);
xnor U22496 (N_22496,N_18088,N_16091);
nor U22497 (N_22497,N_15590,N_16047);
and U22498 (N_22498,N_13183,N_16513);
and U22499 (N_22499,N_13746,N_16053);
xnor U22500 (N_22500,N_17073,N_17795);
nor U22501 (N_22501,N_14372,N_13703);
nand U22502 (N_22502,N_16460,N_15480);
nand U22503 (N_22503,N_16282,N_16449);
nand U22504 (N_22504,N_14819,N_13798);
or U22505 (N_22505,N_17567,N_17607);
nand U22506 (N_22506,N_18076,N_12816);
nor U22507 (N_22507,N_16289,N_18691);
xor U22508 (N_22508,N_14918,N_14423);
xnor U22509 (N_22509,N_18387,N_15068);
nor U22510 (N_22510,N_17867,N_15270);
and U22511 (N_22511,N_16752,N_16616);
nand U22512 (N_22512,N_13018,N_18621);
or U22513 (N_22513,N_15858,N_13549);
nand U22514 (N_22514,N_14180,N_15840);
xnor U22515 (N_22515,N_12934,N_13662);
or U22516 (N_22516,N_13336,N_15416);
or U22517 (N_22517,N_15453,N_17211);
or U22518 (N_22518,N_18211,N_16165);
nor U22519 (N_22519,N_16605,N_18058);
or U22520 (N_22520,N_16953,N_15279);
nand U22521 (N_22521,N_17787,N_18646);
nor U22522 (N_22522,N_14045,N_12663);
nor U22523 (N_22523,N_18604,N_16580);
nor U22524 (N_22524,N_13147,N_16107);
nor U22525 (N_22525,N_17615,N_18255);
and U22526 (N_22526,N_15673,N_17582);
nand U22527 (N_22527,N_13423,N_14339);
nor U22528 (N_22528,N_17770,N_18101);
nand U22529 (N_22529,N_16199,N_14597);
and U22530 (N_22530,N_15777,N_17619);
or U22531 (N_22531,N_17707,N_15450);
nor U22532 (N_22532,N_17083,N_15392);
or U22533 (N_22533,N_13494,N_13462);
and U22534 (N_22534,N_15131,N_17727);
xnor U22535 (N_22535,N_16914,N_18128);
nand U22536 (N_22536,N_14091,N_15695);
nand U22537 (N_22537,N_17637,N_15459);
xnor U22538 (N_22538,N_17457,N_13096);
nand U22539 (N_22539,N_15622,N_15985);
and U22540 (N_22540,N_18144,N_18165);
and U22541 (N_22541,N_18009,N_14123);
nand U22542 (N_22542,N_12964,N_13890);
and U22543 (N_22543,N_17919,N_17090);
xnor U22544 (N_22544,N_17228,N_17605);
xor U22545 (N_22545,N_15474,N_16465);
nand U22546 (N_22546,N_14196,N_18309);
and U22547 (N_22547,N_16180,N_14247);
or U22548 (N_22548,N_16454,N_12522);
xnor U22549 (N_22549,N_12845,N_18429);
xnor U22550 (N_22550,N_15869,N_15013);
and U22551 (N_22551,N_14195,N_16204);
xor U22552 (N_22552,N_14029,N_17442);
or U22553 (N_22553,N_15389,N_14829);
nand U22554 (N_22554,N_16039,N_16528);
and U22555 (N_22555,N_13713,N_16322);
and U22556 (N_22556,N_15350,N_17462);
or U22557 (N_22557,N_14489,N_14573);
and U22558 (N_22558,N_17631,N_16695);
xnor U22559 (N_22559,N_15102,N_14096);
and U22560 (N_22560,N_13421,N_14502);
and U22561 (N_22561,N_14668,N_15454);
nor U22562 (N_22562,N_17892,N_15214);
or U22563 (N_22563,N_13592,N_15723);
nor U22564 (N_22564,N_14675,N_17133);
or U22565 (N_22565,N_14823,N_17020);
nand U22566 (N_22566,N_15359,N_18344);
nor U22567 (N_22567,N_16486,N_15239);
xor U22568 (N_22568,N_16301,N_12747);
nor U22569 (N_22569,N_14010,N_13070);
xor U22570 (N_22570,N_14845,N_13677);
nand U22571 (N_22571,N_13528,N_14381);
or U22572 (N_22572,N_15637,N_14046);
nor U22573 (N_22573,N_16697,N_14992);
and U22574 (N_22574,N_14143,N_15829);
and U22575 (N_22575,N_14658,N_12989);
xor U22576 (N_22576,N_17789,N_13793);
xnor U22577 (N_22577,N_14441,N_13131);
nand U22578 (N_22578,N_17622,N_14614);
xor U22579 (N_22579,N_13180,N_13840);
nor U22580 (N_22580,N_15414,N_15831);
or U22581 (N_22581,N_13193,N_16368);
nand U22582 (N_22582,N_17462,N_16682);
and U22583 (N_22583,N_14182,N_13962);
xor U22584 (N_22584,N_15533,N_13985);
nand U22585 (N_22585,N_17165,N_17895);
nor U22586 (N_22586,N_12919,N_14942);
and U22587 (N_22587,N_12504,N_18667);
nor U22588 (N_22588,N_14413,N_16806);
nor U22589 (N_22589,N_13132,N_13305);
xor U22590 (N_22590,N_16488,N_16545);
or U22591 (N_22591,N_14959,N_15690);
and U22592 (N_22592,N_15566,N_15042);
and U22593 (N_22593,N_16233,N_17135);
nand U22594 (N_22594,N_17522,N_15600);
nor U22595 (N_22595,N_14037,N_15877);
and U22596 (N_22596,N_17381,N_14913);
nor U22597 (N_22597,N_13117,N_12511);
xnor U22598 (N_22598,N_16442,N_13883);
and U22599 (N_22599,N_15115,N_16906);
and U22600 (N_22600,N_14937,N_14524);
and U22601 (N_22601,N_13495,N_17596);
and U22602 (N_22602,N_13319,N_13672);
nand U22603 (N_22603,N_16848,N_18654);
nor U22604 (N_22604,N_15594,N_12828);
and U22605 (N_22605,N_14991,N_17511);
xor U22606 (N_22606,N_14206,N_16016);
nor U22607 (N_22607,N_14586,N_16575);
nor U22608 (N_22608,N_13971,N_17883);
and U22609 (N_22609,N_13514,N_16623);
and U22610 (N_22610,N_13268,N_17926);
and U22611 (N_22611,N_15700,N_15001);
or U22612 (N_22612,N_16081,N_15193);
nor U22613 (N_22613,N_17270,N_13926);
or U22614 (N_22614,N_15877,N_15439);
nor U22615 (N_22615,N_14548,N_15360);
or U22616 (N_22616,N_16062,N_12755);
and U22617 (N_22617,N_18190,N_18731);
and U22618 (N_22618,N_17213,N_17785);
nor U22619 (N_22619,N_14379,N_18058);
nand U22620 (N_22620,N_17706,N_17321);
or U22621 (N_22621,N_12804,N_13360);
nand U22622 (N_22622,N_12869,N_17381);
and U22623 (N_22623,N_17116,N_16204);
or U22624 (N_22624,N_17591,N_16728);
nand U22625 (N_22625,N_13325,N_12548);
or U22626 (N_22626,N_17520,N_17112);
nor U22627 (N_22627,N_17694,N_13511);
nor U22628 (N_22628,N_16537,N_18693);
nand U22629 (N_22629,N_16793,N_15596);
xor U22630 (N_22630,N_18427,N_17587);
nand U22631 (N_22631,N_13951,N_14886);
xor U22632 (N_22632,N_12701,N_15578);
xnor U22633 (N_22633,N_13987,N_16897);
or U22634 (N_22634,N_16503,N_13828);
nand U22635 (N_22635,N_15615,N_16776);
or U22636 (N_22636,N_17460,N_17382);
nand U22637 (N_22637,N_16781,N_15959);
or U22638 (N_22638,N_18343,N_16487);
nor U22639 (N_22639,N_15829,N_17232);
or U22640 (N_22640,N_18748,N_13300);
and U22641 (N_22641,N_17260,N_12684);
nor U22642 (N_22642,N_14898,N_14060);
or U22643 (N_22643,N_13948,N_18297);
nor U22644 (N_22644,N_15405,N_18465);
nor U22645 (N_22645,N_18160,N_18003);
xor U22646 (N_22646,N_13135,N_16753);
nand U22647 (N_22647,N_13530,N_14501);
nor U22648 (N_22648,N_15634,N_14927);
xnor U22649 (N_22649,N_12857,N_17430);
nor U22650 (N_22650,N_18563,N_16082);
and U22651 (N_22651,N_14658,N_16810);
and U22652 (N_22652,N_13146,N_13046);
or U22653 (N_22653,N_16343,N_14811);
nor U22654 (N_22654,N_15671,N_17959);
nor U22655 (N_22655,N_14390,N_14300);
nor U22656 (N_22656,N_17209,N_12536);
and U22657 (N_22657,N_14634,N_15015);
nand U22658 (N_22658,N_12911,N_16083);
or U22659 (N_22659,N_12624,N_14745);
xnor U22660 (N_22660,N_13341,N_14892);
xnor U22661 (N_22661,N_15083,N_17491);
xor U22662 (N_22662,N_14461,N_16132);
nand U22663 (N_22663,N_13342,N_13892);
and U22664 (N_22664,N_12719,N_14238);
xor U22665 (N_22665,N_14184,N_18683);
or U22666 (N_22666,N_18201,N_18051);
xnor U22667 (N_22667,N_13531,N_13657);
nand U22668 (N_22668,N_16862,N_17698);
nand U22669 (N_22669,N_13191,N_18641);
and U22670 (N_22670,N_17849,N_17843);
or U22671 (N_22671,N_13059,N_13748);
xnor U22672 (N_22672,N_14932,N_15102);
nand U22673 (N_22673,N_16897,N_16159);
nand U22674 (N_22674,N_13377,N_14781);
and U22675 (N_22675,N_16247,N_16776);
nand U22676 (N_22676,N_12529,N_12795);
xor U22677 (N_22677,N_18642,N_17683);
xor U22678 (N_22678,N_14029,N_18665);
nand U22679 (N_22679,N_18095,N_17305);
nor U22680 (N_22680,N_16917,N_18609);
or U22681 (N_22681,N_13732,N_14537);
nand U22682 (N_22682,N_14443,N_13028);
nand U22683 (N_22683,N_13135,N_13213);
xnor U22684 (N_22684,N_13053,N_17254);
xnor U22685 (N_22685,N_18192,N_15560);
or U22686 (N_22686,N_13766,N_16521);
and U22687 (N_22687,N_16001,N_16020);
and U22688 (N_22688,N_17480,N_15088);
and U22689 (N_22689,N_15362,N_16649);
or U22690 (N_22690,N_15707,N_15491);
or U22691 (N_22691,N_14444,N_17094);
and U22692 (N_22692,N_13341,N_13579);
xnor U22693 (N_22693,N_14867,N_12712);
and U22694 (N_22694,N_16546,N_17519);
and U22695 (N_22695,N_18638,N_17713);
and U22696 (N_22696,N_13477,N_17775);
nor U22697 (N_22697,N_14241,N_17162);
and U22698 (N_22698,N_17438,N_13900);
xnor U22699 (N_22699,N_16618,N_12980);
or U22700 (N_22700,N_14777,N_16369);
or U22701 (N_22701,N_13550,N_14905);
and U22702 (N_22702,N_15127,N_15349);
nor U22703 (N_22703,N_17790,N_15793);
or U22704 (N_22704,N_18357,N_18228);
nand U22705 (N_22705,N_16105,N_15478);
nor U22706 (N_22706,N_17238,N_13885);
nand U22707 (N_22707,N_17267,N_15730);
nor U22708 (N_22708,N_13655,N_13164);
or U22709 (N_22709,N_14504,N_14633);
and U22710 (N_22710,N_17872,N_13384);
nor U22711 (N_22711,N_17286,N_18611);
xor U22712 (N_22712,N_18171,N_17363);
nor U22713 (N_22713,N_14347,N_15063);
xnor U22714 (N_22714,N_14656,N_18257);
and U22715 (N_22715,N_15636,N_17714);
and U22716 (N_22716,N_15181,N_16248);
xnor U22717 (N_22717,N_16820,N_16530);
nand U22718 (N_22718,N_13258,N_17292);
and U22719 (N_22719,N_16609,N_12839);
and U22720 (N_22720,N_17975,N_13507);
nor U22721 (N_22721,N_14701,N_15968);
nor U22722 (N_22722,N_17355,N_14768);
nand U22723 (N_22723,N_12732,N_15504);
and U22724 (N_22724,N_13318,N_13758);
or U22725 (N_22725,N_15171,N_18435);
or U22726 (N_22726,N_15324,N_15291);
and U22727 (N_22727,N_15112,N_15346);
nor U22728 (N_22728,N_13308,N_17548);
or U22729 (N_22729,N_18143,N_15114);
nor U22730 (N_22730,N_14334,N_16363);
or U22731 (N_22731,N_15433,N_12645);
xor U22732 (N_22732,N_17442,N_17055);
nor U22733 (N_22733,N_17563,N_14888);
or U22734 (N_22734,N_17428,N_18482);
nand U22735 (N_22735,N_15006,N_13239);
or U22736 (N_22736,N_18605,N_15666);
or U22737 (N_22737,N_18535,N_13474);
and U22738 (N_22738,N_15910,N_12566);
and U22739 (N_22739,N_17326,N_15080);
and U22740 (N_22740,N_16716,N_14735);
and U22741 (N_22741,N_18250,N_16007);
nand U22742 (N_22742,N_13724,N_16793);
xnor U22743 (N_22743,N_15221,N_12593);
nand U22744 (N_22744,N_17387,N_15425);
nor U22745 (N_22745,N_18275,N_16978);
xnor U22746 (N_22746,N_17551,N_13840);
nor U22747 (N_22747,N_15237,N_14016);
xor U22748 (N_22748,N_16001,N_15274);
xor U22749 (N_22749,N_16264,N_12889);
xnor U22750 (N_22750,N_13989,N_12839);
nand U22751 (N_22751,N_13436,N_14310);
nand U22752 (N_22752,N_15150,N_17291);
nand U22753 (N_22753,N_16490,N_14639);
nand U22754 (N_22754,N_12535,N_13117);
or U22755 (N_22755,N_14588,N_14058);
xor U22756 (N_22756,N_14762,N_17510);
or U22757 (N_22757,N_12970,N_13362);
nand U22758 (N_22758,N_16283,N_16750);
and U22759 (N_22759,N_16600,N_12786);
nand U22760 (N_22760,N_18193,N_16987);
xor U22761 (N_22761,N_14735,N_17041);
or U22762 (N_22762,N_18208,N_18059);
nand U22763 (N_22763,N_16365,N_14316);
or U22764 (N_22764,N_12909,N_18238);
and U22765 (N_22765,N_14503,N_15575);
and U22766 (N_22766,N_18353,N_13849);
nor U22767 (N_22767,N_13267,N_16604);
nor U22768 (N_22768,N_14914,N_17151);
or U22769 (N_22769,N_17034,N_15505);
xnor U22770 (N_22770,N_18610,N_18023);
nor U22771 (N_22771,N_16270,N_16855);
nor U22772 (N_22772,N_13557,N_13834);
nor U22773 (N_22773,N_12888,N_14038);
or U22774 (N_22774,N_14997,N_16489);
nand U22775 (N_22775,N_17883,N_16371);
xor U22776 (N_22776,N_18463,N_17029);
or U22777 (N_22777,N_12584,N_12817);
nor U22778 (N_22778,N_14523,N_17758);
and U22779 (N_22779,N_18464,N_15973);
and U22780 (N_22780,N_12619,N_17309);
xor U22781 (N_22781,N_18195,N_14332);
or U22782 (N_22782,N_17183,N_13697);
and U22783 (N_22783,N_16195,N_16372);
or U22784 (N_22784,N_15756,N_17060);
nand U22785 (N_22785,N_13482,N_14084);
nor U22786 (N_22786,N_18479,N_15518);
nor U22787 (N_22787,N_14762,N_17042);
or U22788 (N_22788,N_14596,N_17875);
xnor U22789 (N_22789,N_14674,N_13668);
nand U22790 (N_22790,N_14833,N_15769);
xor U22791 (N_22791,N_17948,N_16765);
nand U22792 (N_22792,N_15999,N_16048);
xnor U22793 (N_22793,N_13163,N_17247);
or U22794 (N_22794,N_13743,N_14713);
xor U22795 (N_22795,N_14675,N_15989);
nand U22796 (N_22796,N_17639,N_13210);
and U22797 (N_22797,N_17503,N_14133);
or U22798 (N_22798,N_14863,N_16817);
nor U22799 (N_22799,N_17561,N_18377);
xnor U22800 (N_22800,N_15789,N_16733);
nand U22801 (N_22801,N_14329,N_18306);
and U22802 (N_22802,N_18307,N_16103);
and U22803 (N_22803,N_16784,N_18156);
and U22804 (N_22804,N_18248,N_15301);
and U22805 (N_22805,N_14171,N_14848);
or U22806 (N_22806,N_18273,N_15434);
and U22807 (N_22807,N_13134,N_15465);
nor U22808 (N_22808,N_15812,N_14615);
and U22809 (N_22809,N_13215,N_13810);
nor U22810 (N_22810,N_17444,N_18009);
nor U22811 (N_22811,N_17620,N_14850);
or U22812 (N_22812,N_12761,N_14857);
nor U22813 (N_22813,N_17607,N_14813);
nor U22814 (N_22814,N_13111,N_13541);
or U22815 (N_22815,N_18144,N_15931);
xnor U22816 (N_22816,N_18146,N_17897);
or U22817 (N_22817,N_17367,N_14539);
or U22818 (N_22818,N_17220,N_18427);
xnor U22819 (N_22819,N_17681,N_16883);
nor U22820 (N_22820,N_16500,N_13202);
nand U22821 (N_22821,N_15941,N_14246);
xor U22822 (N_22822,N_17100,N_14206);
nand U22823 (N_22823,N_15925,N_15373);
or U22824 (N_22824,N_13305,N_17757);
and U22825 (N_22825,N_17499,N_17896);
nor U22826 (N_22826,N_18514,N_14214);
or U22827 (N_22827,N_14361,N_17939);
and U22828 (N_22828,N_16388,N_16418);
or U22829 (N_22829,N_13114,N_18601);
nand U22830 (N_22830,N_16403,N_18505);
and U22831 (N_22831,N_16480,N_15205);
nand U22832 (N_22832,N_17962,N_14847);
and U22833 (N_22833,N_12692,N_13829);
nand U22834 (N_22834,N_14950,N_13691);
nand U22835 (N_22835,N_14959,N_15801);
nor U22836 (N_22836,N_14940,N_17721);
nor U22837 (N_22837,N_17312,N_15969);
or U22838 (N_22838,N_15972,N_15781);
nand U22839 (N_22839,N_15903,N_13220);
nor U22840 (N_22840,N_15030,N_16452);
nand U22841 (N_22841,N_18582,N_17414);
nand U22842 (N_22842,N_14245,N_18321);
nand U22843 (N_22843,N_16700,N_14844);
nand U22844 (N_22844,N_12773,N_18324);
nor U22845 (N_22845,N_15643,N_18301);
or U22846 (N_22846,N_14944,N_13046);
or U22847 (N_22847,N_14527,N_16419);
nand U22848 (N_22848,N_17170,N_17716);
nand U22849 (N_22849,N_16166,N_16415);
xnor U22850 (N_22850,N_16754,N_16154);
nand U22851 (N_22851,N_17480,N_12794);
or U22852 (N_22852,N_17066,N_12884);
nand U22853 (N_22853,N_18704,N_18730);
or U22854 (N_22854,N_13817,N_15518);
nand U22855 (N_22855,N_15238,N_14984);
or U22856 (N_22856,N_18724,N_15183);
or U22857 (N_22857,N_12919,N_16031);
nand U22858 (N_22858,N_14630,N_15529);
nand U22859 (N_22859,N_14398,N_18709);
xnor U22860 (N_22860,N_17579,N_17442);
nor U22861 (N_22861,N_17310,N_14054);
nand U22862 (N_22862,N_17650,N_13509);
nor U22863 (N_22863,N_13936,N_17413);
nand U22864 (N_22864,N_15507,N_16105);
or U22865 (N_22865,N_13245,N_14334);
xnor U22866 (N_22866,N_17184,N_15280);
or U22867 (N_22867,N_16022,N_17667);
nand U22868 (N_22868,N_13202,N_12951);
and U22869 (N_22869,N_16449,N_14380);
and U22870 (N_22870,N_14607,N_15746);
xnor U22871 (N_22871,N_16197,N_15940);
xnor U22872 (N_22872,N_14766,N_12739);
xor U22873 (N_22873,N_13296,N_17215);
or U22874 (N_22874,N_17601,N_13822);
nor U22875 (N_22875,N_16262,N_18091);
nand U22876 (N_22876,N_14109,N_15221);
xnor U22877 (N_22877,N_18294,N_14509);
xor U22878 (N_22878,N_17570,N_13330);
xor U22879 (N_22879,N_13599,N_14898);
and U22880 (N_22880,N_17582,N_13162);
and U22881 (N_22881,N_15095,N_16709);
or U22882 (N_22882,N_17728,N_13308);
and U22883 (N_22883,N_13013,N_13529);
or U22884 (N_22884,N_16035,N_18364);
nor U22885 (N_22885,N_18398,N_15500);
nand U22886 (N_22886,N_16436,N_13946);
and U22887 (N_22887,N_17650,N_16586);
and U22888 (N_22888,N_18395,N_15020);
nor U22889 (N_22889,N_12903,N_18018);
xnor U22890 (N_22890,N_17834,N_17417);
and U22891 (N_22891,N_13584,N_15959);
nor U22892 (N_22892,N_16586,N_12758);
or U22893 (N_22893,N_13310,N_18045);
or U22894 (N_22894,N_14554,N_17707);
and U22895 (N_22895,N_15495,N_16007);
nor U22896 (N_22896,N_17580,N_17303);
xnor U22897 (N_22897,N_18528,N_13392);
xor U22898 (N_22898,N_16983,N_13315);
or U22899 (N_22899,N_17533,N_18690);
or U22900 (N_22900,N_14504,N_13018);
and U22901 (N_22901,N_16342,N_15518);
xnor U22902 (N_22902,N_16234,N_13217);
and U22903 (N_22903,N_13607,N_15678);
nor U22904 (N_22904,N_14913,N_14014);
or U22905 (N_22905,N_18356,N_16153);
xnor U22906 (N_22906,N_17177,N_16139);
nor U22907 (N_22907,N_12508,N_14315);
or U22908 (N_22908,N_16220,N_15948);
and U22909 (N_22909,N_15017,N_15561);
or U22910 (N_22910,N_17211,N_17321);
nor U22911 (N_22911,N_13378,N_14962);
and U22912 (N_22912,N_13584,N_15426);
nand U22913 (N_22913,N_14897,N_13188);
xnor U22914 (N_22914,N_17488,N_13504);
xnor U22915 (N_22915,N_15740,N_15643);
nor U22916 (N_22916,N_17451,N_12939);
nor U22917 (N_22917,N_16734,N_14305);
nand U22918 (N_22918,N_16024,N_16397);
nor U22919 (N_22919,N_17705,N_12722);
or U22920 (N_22920,N_14216,N_15258);
nand U22921 (N_22921,N_18640,N_12925);
xor U22922 (N_22922,N_12509,N_14360);
nor U22923 (N_22923,N_16686,N_17672);
or U22924 (N_22924,N_16475,N_14240);
and U22925 (N_22925,N_14883,N_16803);
or U22926 (N_22926,N_13273,N_16026);
nand U22927 (N_22927,N_17001,N_16603);
xor U22928 (N_22928,N_12950,N_14379);
and U22929 (N_22929,N_16925,N_12658);
and U22930 (N_22930,N_15271,N_16399);
nand U22931 (N_22931,N_13919,N_17315);
nor U22932 (N_22932,N_18512,N_16118);
nand U22933 (N_22933,N_16514,N_16815);
or U22934 (N_22934,N_13463,N_16617);
xor U22935 (N_22935,N_18378,N_17248);
xor U22936 (N_22936,N_13326,N_14155);
or U22937 (N_22937,N_17145,N_16756);
nand U22938 (N_22938,N_14567,N_15061);
nor U22939 (N_22939,N_17506,N_13655);
and U22940 (N_22940,N_16455,N_13409);
xnor U22941 (N_22941,N_12560,N_13391);
xnor U22942 (N_22942,N_13487,N_15548);
nand U22943 (N_22943,N_17225,N_15863);
nor U22944 (N_22944,N_12997,N_17392);
and U22945 (N_22945,N_13563,N_14185);
nor U22946 (N_22946,N_15567,N_14347);
nor U22947 (N_22947,N_13246,N_12912);
or U22948 (N_22948,N_15196,N_17480);
xnor U22949 (N_22949,N_14811,N_18510);
and U22950 (N_22950,N_16268,N_16353);
or U22951 (N_22951,N_18355,N_14141);
or U22952 (N_22952,N_13248,N_16960);
or U22953 (N_22953,N_15309,N_12811);
and U22954 (N_22954,N_15257,N_17298);
nor U22955 (N_22955,N_14037,N_13748);
and U22956 (N_22956,N_14361,N_16434);
and U22957 (N_22957,N_14102,N_17586);
nand U22958 (N_22958,N_18311,N_14386);
xnor U22959 (N_22959,N_18308,N_16368);
nand U22960 (N_22960,N_17729,N_18138);
nor U22961 (N_22961,N_18673,N_16848);
and U22962 (N_22962,N_14176,N_18513);
xor U22963 (N_22963,N_17684,N_17398);
and U22964 (N_22964,N_16852,N_17449);
nand U22965 (N_22965,N_17643,N_16241);
nand U22966 (N_22966,N_13553,N_16656);
nor U22967 (N_22967,N_18230,N_14831);
or U22968 (N_22968,N_18496,N_16409);
or U22969 (N_22969,N_14248,N_15545);
or U22970 (N_22970,N_18138,N_12528);
and U22971 (N_22971,N_16993,N_17970);
xnor U22972 (N_22972,N_14326,N_17088);
nand U22973 (N_22973,N_18220,N_15484);
xnor U22974 (N_22974,N_12580,N_18160);
xnor U22975 (N_22975,N_15456,N_16995);
nand U22976 (N_22976,N_12886,N_13776);
or U22977 (N_22977,N_14101,N_13324);
or U22978 (N_22978,N_17720,N_16801);
or U22979 (N_22979,N_18406,N_13420);
nand U22980 (N_22980,N_14503,N_15987);
or U22981 (N_22981,N_12637,N_17376);
and U22982 (N_22982,N_17770,N_14706);
and U22983 (N_22983,N_17458,N_17537);
and U22984 (N_22984,N_13173,N_12598);
and U22985 (N_22985,N_18547,N_17263);
nand U22986 (N_22986,N_16152,N_15195);
nor U22987 (N_22987,N_18377,N_13614);
and U22988 (N_22988,N_12868,N_12601);
and U22989 (N_22989,N_18587,N_15712);
or U22990 (N_22990,N_12599,N_16435);
nand U22991 (N_22991,N_17951,N_18209);
nor U22992 (N_22992,N_18395,N_18316);
and U22993 (N_22993,N_13870,N_14862);
xor U22994 (N_22994,N_16078,N_13259);
or U22995 (N_22995,N_17389,N_12540);
xor U22996 (N_22996,N_12655,N_15785);
or U22997 (N_22997,N_16246,N_12652);
nand U22998 (N_22998,N_14049,N_15733);
nor U22999 (N_22999,N_14811,N_18085);
and U23000 (N_23000,N_18077,N_13998);
and U23001 (N_23001,N_15949,N_15436);
xor U23002 (N_23002,N_14178,N_14456);
nor U23003 (N_23003,N_12532,N_13318);
and U23004 (N_23004,N_15227,N_15730);
and U23005 (N_23005,N_13115,N_17687);
nor U23006 (N_23006,N_17999,N_15269);
or U23007 (N_23007,N_18233,N_17669);
xor U23008 (N_23008,N_13713,N_14835);
nand U23009 (N_23009,N_15594,N_13257);
or U23010 (N_23010,N_14193,N_14661);
and U23011 (N_23011,N_17352,N_17470);
nand U23012 (N_23012,N_14927,N_15624);
or U23013 (N_23013,N_18410,N_14902);
and U23014 (N_23014,N_17335,N_17167);
or U23015 (N_23015,N_16897,N_15598);
nor U23016 (N_23016,N_16286,N_17213);
nand U23017 (N_23017,N_18106,N_18211);
or U23018 (N_23018,N_13926,N_12508);
xnor U23019 (N_23019,N_17055,N_15829);
xor U23020 (N_23020,N_13101,N_14113);
or U23021 (N_23021,N_18134,N_17309);
nor U23022 (N_23022,N_13899,N_16427);
xnor U23023 (N_23023,N_13046,N_16120);
nor U23024 (N_23024,N_17435,N_17330);
or U23025 (N_23025,N_14072,N_15703);
nand U23026 (N_23026,N_13887,N_16397);
or U23027 (N_23027,N_17591,N_14759);
nand U23028 (N_23028,N_13295,N_15369);
nand U23029 (N_23029,N_17520,N_16345);
nor U23030 (N_23030,N_12837,N_18440);
xor U23031 (N_23031,N_12916,N_16317);
xnor U23032 (N_23032,N_14717,N_13925);
or U23033 (N_23033,N_14532,N_17772);
and U23034 (N_23034,N_14823,N_12538);
and U23035 (N_23035,N_15749,N_17533);
and U23036 (N_23036,N_17401,N_14638);
nand U23037 (N_23037,N_12847,N_18709);
or U23038 (N_23038,N_16160,N_15864);
and U23039 (N_23039,N_14192,N_13593);
or U23040 (N_23040,N_18585,N_15596);
or U23041 (N_23041,N_15886,N_16976);
nand U23042 (N_23042,N_15096,N_16195);
and U23043 (N_23043,N_14040,N_14037);
nor U23044 (N_23044,N_18202,N_15220);
xor U23045 (N_23045,N_14809,N_14237);
nand U23046 (N_23046,N_13585,N_15044);
or U23047 (N_23047,N_14884,N_17470);
xor U23048 (N_23048,N_14029,N_15380);
xnor U23049 (N_23049,N_14459,N_13144);
nand U23050 (N_23050,N_13364,N_12986);
or U23051 (N_23051,N_15107,N_12747);
and U23052 (N_23052,N_17762,N_12751);
nor U23053 (N_23053,N_16747,N_12971);
or U23054 (N_23054,N_15277,N_12703);
and U23055 (N_23055,N_18267,N_16732);
or U23056 (N_23056,N_15633,N_17971);
nor U23057 (N_23057,N_18605,N_18041);
or U23058 (N_23058,N_18740,N_18205);
nor U23059 (N_23059,N_16099,N_16894);
or U23060 (N_23060,N_17590,N_13543);
nand U23061 (N_23061,N_16305,N_14080);
or U23062 (N_23062,N_14407,N_17834);
or U23063 (N_23063,N_18481,N_16545);
and U23064 (N_23064,N_17172,N_16166);
xor U23065 (N_23065,N_13063,N_18598);
and U23066 (N_23066,N_13356,N_14349);
xnor U23067 (N_23067,N_15461,N_12938);
xor U23068 (N_23068,N_14434,N_14997);
xnor U23069 (N_23069,N_16349,N_14270);
and U23070 (N_23070,N_13038,N_18663);
or U23071 (N_23071,N_12651,N_14490);
nor U23072 (N_23072,N_17962,N_16233);
or U23073 (N_23073,N_13418,N_16206);
and U23074 (N_23074,N_16660,N_17955);
xor U23075 (N_23075,N_17569,N_18543);
xor U23076 (N_23076,N_14116,N_16320);
nand U23077 (N_23077,N_18193,N_12867);
nor U23078 (N_23078,N_12851,N_14898);
or U23079 (N_23079,N_14882,N_14263);
or U23080 (N_23080,N_17190,N_13412);
or U23081 (N_23081,N_12715,N_18405);
and U23082 (N_23082,N_12705,N_14047);
and U23083 (N_23083,N_18480,N_16011);
nand U23084 (N_23084,N_14679,N_13961);
nor U23085 (N_23085,N_17962,N_16833);
nor U23086 (N_23086,N_15531,N_13281);
and U23087 (N_23087,N_16031,N_14438);
or U23088 (N_23088,N_15814,N_14018);
and U23089 (N_23089,N_17155,N_13514);
or U23090 (N_23090,N_14788,N_17688);
or U23091 (N_23091,N_13265,N_16512);
and U23092 (N_23092,N_17322,N_13608);
and U23093 (N_23093,N_17486,N_18374);
nor U23094 (N_23094,N_15700,N_14002);
xor U23095 (N_23095,N_17705,N_15027);
or U23096 (N_23096,N_18620,N_14461);
or U23097 (N_23097,N_15725,N_17678);
xor U23098 (N_23098,N_18465,N_18357);
nor U23099 (N_23099,N_14367,N_12523);
nor U23100 (N_23100,N_16119,N_18341);
xor U23101 (N_23101,N_15947,N_14339);
nand U23102 (N_23102,N_14133,N_13545);
xnor U23103 (N_23103,N_18509,N_16445);
or U23104 (N_23104,N_17598,N_12563);
or U23105 (N_23105,N_17490,N_12894);
xor U23106 (N_23106,N_14296,N_15358);
nand U23107 (N_23107,N_16950,N_17589);
xnor U23108 (N_23108,N_17340,N_18516);
nor U23109 (N_23109,N_14503,N_12777);
or U23110 (N_23110,N_14793,N_14046);
nand U23111 (N_23111,N_13428,N_13794);
nand U23112 (N_23112,N_16187,N_15890);
and U23113 (N_23113,N_16963,N_17050);
and U23114 (N_23114,N_17452,N_15597);
or U23115 (N_23115,N_17270,N_18479);
or U23116 (N_23116,N_12535,N_17792);
and U23117 (N_23117,N_17760,N_14664);
nand U23118 (N_23118,N_17377,N_14031);
xnor U23119 (N_23119,N_13340,N_13331);
and U23120 (N_23120,N_13321,N_17814);
xnor U23121 (N_23121,N_18569,N_18731);
xor U23122 (N_23122,N_17451,N_15021);
or U23123 (N_23123,N_18557,N_14223);
xor U23124 (N_23124,N_13939,N_13197);
xor U23125 (N_23125,N_17091,N_18560);
or U23126 (N_23126,N_18409,N_13827);
nor U23127 (N_23127,N_17616,N_16778);
and U23128 (N_23128,N_14706,N_17189);
nor U23129 (N_23129,N_13214,N_13014);
nor U23130 (N_23130,N_13501,N_12822);
nor U23131 (N_23131,N_17843,N_12648);
and U23132 (N_23132,N_16330,N_14604);
nor U23133 (N_23133,N_17613,N_17630);
nor U23134 (N_23134,N_15300,N_16728);
and U23135 (N_23135,N_17190,N_13665);
nand U23136 (N_23136,N_13405,N_18119);
or U23137 (N_23137,N_15769,N_16662);
or U23138 (N_23138,N_13839,N_13918);
nor U23139 (N_23139,N_17572,N_13837);
xor U23140 (N_23140,N_14382,N_16762);
nand U23141 (N_23141,N_16142,N_18689);
or U23142 (N_23142,N_16433,N_17848);
and U23143 (N_23143,N_13881,N_15763);
nor U23144 (N_23144,N_15026,N_15917);
xnor U23145 (N_23145,N_14434,N_14210);
nand U23146 (N_23146,N_12977,N_16477);
nor U23147 (N_23147,N_15089,N_14820);
nor U23148 (N_23148,N_16072,N_14795);
xor U23149 (N_23149,N_15035,N_18480);
xor U23150 (N_23150,N_13750,N_17972);
xor U23151 (N_23151,N_16956,N_17077);
nand U23152 (N_23152,N_14758,N_15754);
and U23153 (N_23153,N_16611,N_18731);
nand U23154 (N_23154,N_13661,N_14408);
xnor U23155 (N_23155,N_17474,N_15188);
nor U23156 (N_23156,N_17095,N_17249);
xnor U23157 (N_23157,N_13372,N_17350);
xor U23158 (N_23158,N_17654,N_16024);
nor U23159 (N_23159,N_17816,N_13587);
or U23160 (N_23160,N_13446,N_18291);
nand U23161 (N_23161,N_14989,N_16456);
xnor U23162 (N_23162,N_13569,N_13667);
xnor U23163 (N_23163,N_14172,N_16327);
xnor U23164 (N_23164,N_13400,N_14036);
nor U23165 (N_23165,N_15721,N_16253);
nand U23166 (N_23166,N_16365,N_16470);
nor U23167 (N_23167,N_16689,N_17378);
nor U23168 (N_23168,N_13807,N_13543);
or U23169 (N_23169,N_17552,N_15442);
nor U23170 (N_23170,N_15856,N_13470);
or U23171 (N_23171,N_15167,N_14911);
nand U23172 (N_23172,N_15471,N_16327);
or U23173 (N_23173,N_14063,N_14803);
or U23174 (N_23174,N_16551,N_16445);
nand U23175 (N_23175,N_17712,N_13413);
or U23176 (N_23176,N_12964,N_14240);
or U23177 (N_23177,N_14349,N_17277);
nand U23178 (N_23178,N_15241,N_14116);
nor U23179 (N_23179,N_14012,N_16366);
nand U23180 (N_23180,N_13292,N_16339);
and U23181 (N_23181,N_14270,N_17697);
xor U23182 (N_23182,N_18269,N_13029);
nand U23183 (N_23183,N_15817,N_16737);
nand U23184 (N_23184,N_17222,N_15998);
and U23185 (N_23185,N_15905,N_12964);
nor U23186 (N_23186,N_16786,N_15824);
and U23187 (N_23187,N_17917,N_17530);
nand U23188 (N_23188,N_18286,N_16099);
or U23189 (N_23189,N_14133,N_12602);
or U23190 (N_23190,N_17119,N_18025);
xnor U23191 (N_23191,N_14872,N_17175);
nor U23192 (N_23192,N_18730,N_14345);
nor U23193 (N_23193,N_12538,N_15934);
xnor U23194 (N_23194,N_15357,N_16468);
nor U23195 (N_23195,N_18080,N_14747);
and U23196 (N_23196,N_15802,N_14523);
and U23197 (N_23197,N_17132,N_13830);
and U23198 (N_23198,N_15976,N_18583);
xor U23199 (N_23199,N_12778,N_15135);
nor U23200 (N_23200,N_14928,N_16086);
xnor U23201 (N_23201,N_12713,N_12592);
and U23202 (N_23202,N_14373,N_12504);
nand U23203 (N_23203,N_13607,N_17081);
xor U23204 (N_23204,N_16228,N_18498);
nor U23205 (N_23205,N_12631,N_13948);
nand U23206 (N_23206,N_17841,N_12597);
or U23207 (N_23207,N_15961,N_15945);
nand U23208 (N_23208,N_15936,N_12898);
or U23209 (N_23209,N_17681,N_17209);
and U23210 (N_23210,N_16630,N_14066);
nand U23211 (N_23211,N_15667,N_16684);
xnor U23212 (N_23212,N_17647,N_15206);
or U23213 (N_23213,N_18687,N_16808);
and U23214 (N_23214,N_14913,N_12612);
and U23215 (N_23215,N_15148,N_14491);
xnor U23216 (N_23216,N_16712,N_14310);
and U23217 (N_23217,N_18301,N_13985);
nand U23218 (N_23218,N_16730,N_17632);
or U23219 (N_23219,N_17782,N_18611);
nand U23220 (N_23220,N_18014,N_12821);
and U23221 (N_23221,N_12850,N_16190);
or U23222 (N_23222,N_17741,N_14574);
xnor U23223 (N_23223,N_13353,N_17917);
and U23224 (N_23224,N_14464,N_17536);
xnor U23225 (N_23225,N_16613,N_15083);
or U23226 (N_23226,N_15068,N_14334);
xnor U23227 (N_23227,N_15448,N_14601);
nand U23228 (N_23228,N_15608,N_18238);
nand U23229 (N_23229,N_13965,N_14506);
nand U23230 (N_23230,N_18159,N_15342);
nand U23231 (N_23231,N_15052,N_16790);
xor U23232 (N_23232,N_14347,N_17299);
and U23233 (N_23233,N_13884,N_14407);
and U23234 (N_23234,N_13025,N_14649);
and U23235 (N_23235,N_18565,N_12962);
and U23236 (N_23236,N_14642,N_15222);
or U23237 (N_23237,N_13364,N_14130);
xor U23238 (N_23238,N_15763,N_17330);
and U23239 (N_23239,N_17008,N_17471);
or U23240 (N_23240,N_16326,N_17080);
and U23241 (N_23241,N_18403,N_12934);
nor U23242 (N_23242,N_15032,N_17664);
xnor U23243 (N_23243,N_16187,N_13031);
nand U23244 (N_23244,N_16037,N_13292);
or U23245 (N_23245,N_16123,N_16750);
xnor U23246 (N_23246,N_17308,N_18095);
and U23247 (N_23247,N_16559,N_13585);
nand U23248 (N_23248,N_12755,N_17782);
and U23249 (N_23249,N_14695,N_16333);
xnor U23250 (N_23250,N_16438,N_17371);
and U23251 (N_23251,N_18335,N_15756);
nor U23252 (N_23252,N_16605,N_13347);
or U23253 (N_23253,N_14486,N_12615);
and U23254 (N_23254,N_15899,N_12770);
nor U23255 (N_23255,N_14915,N_15073);
or U23256 (N_23256,N_18562,N_12702);
xnor U23257 (N_23257,N_17883,N_16385);
xor U23258 (N_23258,N_18015,N_16074);
nand U23259 (N_23259,N_17871,N_17948);
and U23260 (N_23260,N_13107,N_17570);
nor U23261 (N_23261,N_16081,N_17675);
and U23262 (N_23262,N_12551,N_17194);
nand U23263 (N_23263,N_15864,N_18725);
nor U23264 (N_23264,N_14520,N_15251);
or U23265 (N_23265,N_16694,N_14269);
nor U23266 (N_23266,N_13351,N_17346);
or U23267 (N_23267,N_13579,N_16700);
xor U23268 (N_23268,N_12647,N_15399);
nand U23269 (N_23269,N_13182,N_12950);
and U23270 (N_23270,N_14790,N_13551);
nor U23271 (N_23271,N_18557,N_13054);
nand U23272 (N_23272,N_13084,N_17680);
and U23273 (N_23273,N_13470,N_18711);
and U23274 (N_23274,N_14811,N_18714);
nand U23275 (N_23275,N_12847,N_13664);
nor U23276 (N_23276,N_17332,N_15782);
xor U23277 (N_23277,N_14104,N_14278);
nand U23278 (N_23278,N_16760,N_13621);
and U23279 (N_23279,N_16086,N_15439);
and U23280 (N_23280,N_16410,N_18391);
nor U23281 (N_23281,N_13313,N_15074);
or U23282 (N_23282,N_13843,N_16336);
nor U23283 (N_23283,N_16640,N_13004);
nor U23284 (N_23284,N_16417,N_16939);
or U23285 (N_23285,N_13874,N_16818);
or U23286 (N_23286,N_15724,N_17490);
or U23287 (N_23287,N_18353,N_12689);
or U23288 (N_23288,N_13319,N_16433);
nor U23289 (N_23289,N_14870,N_12937);
xnor U23290 (N_23290,N_14184,N_12607);
and U23291 (N_23291,N_15980,N_15686);
or U23292 (N_23292,N_16902,N_18544);
xnor U23293 (N_23293,N_16672,N_13698);
nor U23294 (N_23294,N_17256,N_17924);
or U23295 (N_23295,N_16783,N_15566);
or U23296 (N_23296,N_16386,N_17858);
nand U23297 (N_23297,N_14738,N_17000);
nand U23298 (N_23298,N_18216,N_16450);
and U23299 (N_23299,N_15405,N_18236);
and U23300 (N_23300,N_16263,N_13031);
nor U23301 (N_23301,N_14141,N_13845);
nor U23302 (N_23302,N_16293,N_16741);
or U23303 (N_23303,N_18383,N_15813);
or U23304 (N_23304,N_17642,N_13677);
nor U23305 (N_23305,N_15536,N_16289);
xor U23306 (N_23306,N_12865,N_14756);
nor U23307 (N_23307,N_12998,N_15262);
and U23308 (N_23308,N_16545,N_14241);
or U23309 (N_23309,N_16838,N_14789);
or U23310 (N_23310,N_15130,N_13448);
or U23311 (N_23311,N_18435,N_12570);
or U23312 (N_23312,N_18280,N_17511);
nand U23313 (N_23313,N_18022,N_18723);
or U23314 (N_23314,N_14019,N_14653);
nor U23315 (N_23315,N_17207,N_18413);
nor U23316 (N_23316,N_17759,N_14920);
xnor U23317 (N_23317,N_15887,N_14564);
nor U23318 (N_23318,N_15981,N_13753);
nor U23319 (N_23319,N_13203,N_14742);
xor U23320 (N_23320,N_15301,N_14639);
and U23321 (N_23321,N_14988,N_18244);
or U23322 (N_23322,N_17962,N_16751);
and U23323 (N_23323,N_16686,N_12987);
xor U23324 (N_23324,N_15568,N_18235);
xor U23325 (N_23325,N_13715,N_16385);
nand U23326 (N_23326,N_14219,N_12688);
nor U23327 (N_23327,N_18297,N_13087);
xor U23328 (N_23328,N_16731,N_13492);
and U23329 (N_23329,N_13612,N_15074);
xor U23330 (N_23330,N_16170,N_14880);
and U23331 (N_23331,N_17002,N_16676);
or U23332 (N_23332,N_17935,N_15245);
or U23333 (N_23333,N_16471,N_14457);
or U23334 (N_23334,N_13437,N_18467);
and U23335 (N_23335,N_16726,N_17282);
and U23336 (N_23336,N_16318,N_15598);
nor U23337 (N_23337,N_16862,N_16816);
xnor U23338 (N_23338,N_16140,N_16222);
or U23339 (N_23339,N_16383,N_15165);
nor U23340 (N_23340,N_17590,N_15610);
xor U23341 (N_23341,N_18145,N_12850);
xor U23342 (N_23342,N_14407,N_13642);
xnor U23343 (N_23343,N_15379,N_16404);
or U23344 (N_23344,N_13969,N_12953);
nor U23345 (N_23345,N_14598,N_13879);
and U23346 (N_23346,N_16850,N_15265);
or U23347 (N_23347,N_13740,N_13961);
and U23348 (N_23348,N_15100,N_17090);
nor U23349 (N_23349,N_13003,N_14699);
and U23350 (N_23350,N_18371,N_13288);
nand U23351 (N_23351,N_18386,N_15623);
xnor U23352 (N_23352,N_12552,N_15294);
nor U23353 (N_23353,N_17115,N_13816);
and U23354 (N_23354,N_17776,N_13640);
xnor U23355 (N_23355,N_18483,N_13352);
or U23356 (N_23356,N_16355,N_16653);
or U23357 (N_23357,N_17068,N_12729);
nand U23358 (N_23358,N_12933,N_13168);
nand U23359 (N_23359,N_15012,N_17822);
xnor U23360 (N_23360,N_16926,N_15420);
nand U23361 (N_23361,N_17776,N_15583);
xnor U23362 (N_23362,N_13398,N_16272);
xor U23363 (N_23363,N_16167,N_13642);
and U23364 (N_23364,N_14564,N_17587);
nor U23365 (N_23365,N_12912,N_13588);
and U23366 (N_23366,N_14507,N_15581);
or U23367 (N_23367,N_13490,N_17899);
xnor U23368 (N_23368,N_13159,N_16750);
xor U23369 (N_23369,N_15896,N_18192);
or U23370 (N_23370,N_18684,N_12775);
nand U23371 (N_23371,N_16437,N_18319);
or U23372 (N_23372,N_14601,N_13624);
xnor U23373 (N_23373,N_12532,N_12909);
and U23374 (N_23374,N_14971,N_17744);
or U23375 (N_23375,N_16525,N_16759);
or U23376 (N_23376,N_13105,N_18459);
and U23377 (N_23377,N_14361,N_12641);
or U23378 (N_23378,N_13647,N_12708);
nor U23379 (N_23379,N_13137,N_16523);
nand U23380 (N_23380,N_17351,N_14327);
xnor U23381 (N_23381,N_17923,N_12736);
xnor U23382 (N_23382,N_12581,N_18061);
xor U23383 (N_23383,N_13587,N_13401);
or U23384 (N_23384,N_17743,N_17798);
nor U23385 (N_23385,N_13750,N_18423);
nand U23386 (N_23386,N_12749,N_16222);
nor U23387 (N_23387,N_18225,N_17146);
nor U23388 (N_23388,N_16933,N_14444);
or U23389 (N_23389,N_14672,N_14578);
nor U23390 (N_23390,N_12961,N_17079);
or U23391 (N_23391,N_12507,N_18638);
and U23392 (N_23392,N_13372,N_17049);
and U23393 (N_23393,N_18369,N_17206);
and U23394 (N_23394,N_18616,N_14011);
or U23395 (N_23395,N_14379,N_12510);
nor U23396 (N_23396,N_14052,N_18387);
xnor U23397 (N_23397,N_15397,N_17915);
nand U23398 (N_23398,N_12558,N_12999);
xnor U23399 (N_23399,N_17663,N_12847);
or U23400 (N_23400,N_16468,N_12933);
and U23401 (N_23401,N_12896,N_15123);
or U23402 (N_23402,N_12969,N_14147);
nand U23403 (N_23403,N_14801,N_18647);
xor U23404 (N_23404,N_13184,N_16778);
nand U23405 (N_23405,N_17502,N_17038);
and U23406 (N_23406,N_15853,N_16024);
nor U23407 (N_23407,N_16922,N_15458);
or U23408 (N_23408,N_14647,N_17025);
and U23409 (N_23409,N_16277,N_13028);
and U23410 (N_23410,N_15428,N_16343);
xnor U23411 (N_23411,N_16870,N_15810);
xnor U23412 (N_23412,N_13306,N_17401);
nand U23413 (N_23413,N_16229,N_13514);
nor U23414 (N_23414,N_12738,N_17391);
or U23415 (N_23415,N_14804,N_15667);
nor U23416 (N_23416,N_14437,N_13952);
xnor U23417 (N_23417,N_13726,N_14812);
nand U23418 (N_23418,N_18540,N_15291);
and U23419 (N_23419,N_12816,N_14524);
nor U23420 (N_23420,N_15008,N_14469);
and U23421 (N_23421,N_18712,N_17463);
and U23422 (N_23422,N_18297,N_17256);
and U23423 (N_23423,N_14326,N_16821);
nand U23424 (N_23424,N_13995,N_17461);
or U23425 (N_23425,N_15816,N_17932);
or U23426 (N_23426,N_13583,N_18302);
or U23427 (N_23427,N_17658,N_16743);
nor U23428 (N_23428,N_14391,N_15370);
nor U23429 (N_23429,N_16457,N_15748);
nand U23430 (N_23430,N_15199,N_17743);
or U23431 (N_23431,N_18321,N_17874);
nor U23432 (N_23432,N_16424,N_16576);
and U23433 (N_23433,N_15903,N_15344);
nand U23434 (N_23434,N_14504,N_13973);
xor U23435 (N_23435,N_17610,N_14419);
xnor U23436 (N_23436,N_18717,N_12634);
and U23437 (N_23437,N_17643,N_15296);
or U23438 (N_23438,N_14296,N_13681);
xnor U23439 (N_23439,N_16510,N_13689);
nand U23440 (N_23440,N_15955,N_16704);
nand U23441 (N_23441,N_14583,N_17584);
nor U23442 (N_23442,N_12721,N_14987);
nand U23443 (N_23443,N_14061,N_14528);
xnor U23444 (N_23444,N_14997,N_13142);
or U23445 (N_23445,N_18087,N_15272);
nand U23446 (N_23446,N_14708,N_15257);
xor U23447 (N_23447,N_12917,N_15343);
xnor U23448 (N_23448,N_13641,N_13285);
nand U23449 (N_23449,N_17215,N_16577);
nand U23450 (N_23450,N_14847,N_18328);
nor U23451 (N_23451,N_16802,N_18449);
nand U23452 (N_23452,N_18268,N_13440);
or U23453 (N_23453,N_12764,N_12908);
nand U23454 (N_23454,N_17238,N_12797);
or U23455 (N_23455,N_13667,N_14510);
xor U23456 (N_23456,N_16337,N_17244);
and U23457 (N_23457,N_15346,N_13160);
nand U23458 (N_23458,N_13643,N_13199);
nand U23459 (N_23459,N_17611,N_15961);
nor U23460 (N_23460,N_18290,N_15697);
nand U23461 (N_23461,N_15804,N_18559);
xor U23462 (N_23462,N_17207,N_15324);
or U23463 (N_23463,N_13553,N_13249);
nor U23464 (N_23464,N_13573,N_17171);
and U23465 (N_23465,N_13013,N_15242);
or U23466 (N_23466,N_17832,N_13043);
nor U23467 (N_23467,N_15769,N_15502);
and U23468 (N_23468,N_17022,N_13437);
and U23469 (N_23469,N_15908,N_13430);
nand U23470 (N_23470,N_18366,N_15144);
or U23471 (N_23471,N_17371,N_17484);
nand U23472 (N_23472,N_14684,N_16430);
nand U23473 (N_23473,N_17886,N_15521);
or U23474 (N_23474,N_17604,N_12716);
xnor U23475 (N_23475,N_16703,N_13378);
nor U23476 (N_23476,N_16307,N_12794);
and U23477 (N_23477,N_14753,N_14323);
nor U23478 (N_23478,N_16496,N_15774);
or U23479 (N_23479,N_18385,N_16301);
nand U23480 (N_23480,N_17232,N_15708);
nand U23481 (N_23481,N_16178,N_17263);
nor U23482 (N_23482,N_14682,N_15564);
xor U23483 (N_23483,N_17876,N_14085);
and U23484 (N_23484,N_15439,N_16145);
or U23485 (N_23485,N_13994,N_16412);
xor U23486 (N_23486,N_16879,N_15588);
or U23487 (N_23487,N_13538,N_15094);
xnor U23488 (N_23488,N_14630,N_14262);
nor U23489 (N_23489,N_18079,N_16669);
and U23490 (N_23490,N_13717,N_17422);
and U23491 (N_23491,N_16616,N_17959);
or U23492 (N_23492,N_16894,N_16025);
xor U23493 (N_23493,N_17667,N_16673);
or U23494 (N_23494,N_13858,N_14156);
xor U23495 (N_23495,N_16204,N_15663);
or U23496 (N_23496,N_18263,N_13209);
or U23497 (N_23497,N_18414,N_16518);
nor U23498 (N_23498,N_15252,N_17929);
and U23499 (N_23499,N_18481,N_16721);
and U23500 (N_23500,N_12928,N_16389);
and U23501 (N_23501,N_16912,N_13280);
xnor U23502 (N_23502,N_17212,N_17080);
and U23503 (N_23503,N_12938,N_16033);
nand U23504 (N_23504,N_18052,N_15680);
nand U23505 (N_23505,N_16991,N_17087);
nor U23506 (N_23506,N_16755,N_16109);
xnor U23507 (N_23507,N_17612,N_15251);
and U23508 (N_23508,N_17709,N_18147);
and U23509 (N_23509,N_14328,N_16750);
and U23510 (N_23510,N_14931,N_12811);
nor U23511 (N_23511,N_12902,N_16127);
nor U23512 (N_23512,N_12591,N_18177);
nand U23513 (N_23513,N_12889,N_13246);
xor U23514 (N_23514,N_13844,N_18050);
and U23515 (N_23515,N_18446,N_16251);
nor U23516 (N_23516,N_16795,N_18126);
and U23517 (N_23517,N_13108,N_12999);
nand U23518 (N_23518,N_17621,N_13531);
or U23519 (N_23519,N_18686,N_14672);
or U23520 (N_23520,N_12750,N_15469);
and U23521 (N_23521,N_14263,N_13243);
xor U23522 (N_23522,N_12989,N_18369);
nor U23523 (N_23523,N_14329,N_14938);
xor U23524 (N_23524,N_15452,N_16088);
or U23525 (N_23525,N_15640,N_15052);
xnor U23526 (N_23526,N_12854,N_15503);
or U23527 (N_23527,N_17390,N_15917);
xnor U23528 (N_23528,N_13324,N_14486);
or U23529 (N_23529,N_17428,N_16447);
xor U23530 (N_23530,N_17753,N_14952);
xnor U23531 (N_23531,N_13107,N_17062);
nor U23532 (N_23532,N_18101,N_17200);
xor U23533 (N_23533,N_17388,N_13668);
nand U23534 (N_23534,N_13560,N_16563);
or U23535 (N_23535,N_14621,N_12865);
or U23536 (N_23536,N_17743,N_14661);
nand U23537 (N_23537,N_18452,N_18736);
nor U23538 (N_23538,N_15783,N_12846);
nor U23539 (N_23539,N_15343,N_14596);
nand U23540 (N_23540,N_12859,N_18474);
nand U23541 (N_23541,N_13076,N_17832);
nor U23542 (N_23542,N_14061,N_15241);
or U23543 (N_23543,N_15589,N_16712);
and U23544 (N_23544,N_12552,N_13563);
nand U23545 (N_23545,N_18118,N_14691);
and U23546 (N_23546,N_14014,N_15268);
nand U23547 (N_23547,N_12939,N_13347);
nand U23548 (N_23548,N_12954,N_14936);
or U23549 (N_23549,N_18420,N_16161);
nand U23550 (N_23550,N_17439,N_14652);
and U23551 (N_23551,N_15637,N_14687);
nor U23552 (N_23552,N_17084,N_14238);
and U23553 (N_23553,N_14985,N_13031);
nor U23554 (N_23554,N_15090,N_16173);
xor U23555 (N_23555,N_14966,N_18292);
nand U23556 (N_23556,N_16300,N_17440);
or U23557 (N_23557,N_13333,N_17144);
and U23558 (N_23558,N_17038,N_13155);
xor U23559 (N_23559,N_17748,N_15996);
nand U23560 (N_23560,N_14532,N_13420);
nor U23561 (N_23561,N_17738,N_14766);
and U23562 (N_23562,N_12515,N_15136);
nand U23563 (N_23563,N_15818,N_14753);
and U23564 (N_23564,N_16880,N_18041);
nand U23565 (N_23565,N_14611,N_17167);
nand U23566 (N_23566,N_17867,N_14686);
and U23567 (N_23567,N_16581,N_12647);
xor U23568 (N_23568,N_13683,N_14275);
nand U23569 (N_23569,N_13442,N_15969);
nor U23570 (N_23570,N_16998,N_17499);
xnor U23571 (N_23571,N_13988,N_17236);
nand U23572 (N_23572,N_17001,N_15399);
nor U23573 (N_23573,N_15766,N_14041);
and U23574 (N_23574,N_16807,N_17907);
nand U23575 (N_23575,N_15819,N_14381);
nand U23576 (N_23576,N_17900,N_17978);
or U23577 (N_23577,N_16733,N_17382);
nand U23578 (N_23578,N_17397,N_17985);
xor U23579 (N_23579,N_15228,N_16688);
nor U23580 (N_23580,N_18223,N_18393);
nor U23581 (N_23581,N_14121,N_12901);
nand U23582 (N_23582,N_17865,N_14374);
xnor U23583 (N_23583,N_13562,N_14776);
nor U23584 (N_23584,N_17590,N_14577);
nor U23585 (N_23585,N_18378,N_15609);
and U23586 (N_23586,N_14140,N_15897);
xor U23587 (N_23587,N_15602,N_15046);
and U23588 (N_23588,N_18667,N_12509);
nor U23589 (N_23589,N_13804,N_17983);
xnor U23590 (N_23590,N_15286,N_18056);
and U23591 (N_23591,N_18053,N_18461);
xor U23592 (N_23592,N_16577,N_18508);
nor U23593 (N_23593,N_16867,N_17661);
xor U23594 (N_23594,N_18140,N_16001);
nand U23595 (N_23595,N_18153,N_13994);
nor U23596 (N_23596,N_13942,N_16757);
or U23597 (N_23597,N_17082,N_16076);
nor U23598 (N_23598,N_17251,N_15691);
xor U23599 (N_23599,N_15524,N_15903);
nor U23600 (N_23600,N_14233,N_15089);
and U23601 (N_23601,N_15303,N_14363);
nor U23602 (N_23602,N_15226,N_14363);
or U23603 (N_23603,N_18179,N_14234);
nor U23604 (N_23604,N_14009,N_13966);
and U23605 (N_23605,N_12704,N_15558);
or U23606 (N_23606,N_15107,N_12578);
or U23607 (N_23607,N_14595,N_17599);
nand U23608 (N_23608,N_18520,N_13559);
and U23609 (N_23609,N_16507,N_17108);
nor U23610 (N_23610,N_17740,N_16632);
nand U23611 (N_23611,N_16659,N_16896);
nand U23612 (N_23612,N_16684,N_16931);
nor U23613 (N_23613,N_13394,N_18336);
or U23614 (N_23614,N_12979,N_17624);
xnor U23615 (N_23615,N_13407,N_13564);
xnor U23616 (N_23616,N_15277,N_16827);
and U23617 (N_23617,N_13172,N_13975);
or U23618 (N_23618,N_16183,N_12649);
xnor U23619 (N_23619,N_13987,N_15641);
or U23620 (N_23620,N_12793,N_17405);
and U23621 (N_23621,N_18687,N_17143);
xor U23622 (N_23622,N_13490,N_16050);
xnor U23623 (N_23623,N_17304,N_13053);
or U23624 (N_23624,N_15654,N_12779);
xnor U23625 (N_23625,N_15132,N_16864);
nor U23626 (N_23626,N_12662,N_18582);
or U23627 (N_23627,N_17751,N_16292);
xnor U23628 (N_23628,N_17021,N_13308);
or U23629 (N_23629,N_16023,N_13849);
nor U23630 (N_23630,N_14972,N_18352);
nor U23631 (N_23631,N_15491,N_14295);
nand U23632 (N_23632,N_13076,N_13582);
or U23633 (N_23633,N_13965,N_12815);
nor U23634 (N_23634,N_16638,N_17348);
or U23635 (N_23635,N_14112,N_18126);
nand U23636 (N_23636,N_18431,N_16301);
xnor U23637 (N_23637,N_16299,N_13782);
xor U23638 (N_23638,N_14904,N_13848);
or U23639 (N_23639,N_12672,N_13388);
xor U23640 (N_23640,N_15083,N_15169);
nor U23641 (N_23641,N_16300,N_13091);
or U23642 (N_23642,N_16627,N_13584);
or U23643 (N_23643,N_14185,N_13909);
nor U23644 (N_23644,N_15695,N_15247);
nor U23645 (N_23645,N_14158,N_15006);
xor U23646 (N_23646,N_13689,N_17192);
xor U23647 (N_23647,N_16689,N_14191);
nor U23648 (N_23648,N_14603,N_17219);
nor U23649 (N_23649,N_13980,N_18678);
nand U23650 (N_23650,N_16685,N_13407);
and U23651 (N_23651,N_18244,N_13297);
nand U23652 (N_23652,N_13975,N_17802);
or U23653 (N_23653,N_14756,N_12574);
xor U23654 (N_23654,N_14481,N_16681);
and U23655 (N_23655,N_13326,N_17780);
xnor U23656 (N_23656,N_12752,N_15872);
and U23657 (N_23657,N_15643,N_13435);
nand U23658 (N_23658,N_14926,N_15394);
xor U23659 (N_23659,N_14770,N_14514);
nor U23660 (N_23660,N_15216,N_18528);
xor U23661 (N_23661,N_17411,N_13011);
or U23662 (N_23662,N_12649,N_12622);
and U23663 (N_23663,N_17731,N_17567);
and U23664 (N_23664,N_15324,N_17336);
xor U23665 (N_23665,N_16601,N_13021);
nor U23666 (N_23666,N_14874,N_15880);
nor U23667 (N_23667,N_18425,N_18365);
nor U23668 (N_23668,N_16343,N_16518);
and U23669 (N_23669,N_15231,N_17611);
nand U23670 (N_23670,N_16584,N_15728);
nor U23671 (N_23671,N_17903,N_15157);
nand U23672 (N_23672,N_17226,N_13393);
xnor U23673 (N_23673,N_14045,N_15657);
or U23674 (N_23674,N_14749,N_13360);
xor U23675 (N_23675,N_15388,N_17824);
xnor U23676 (N_23676,N_13680,N_15825);
nand U23677 (N_23677,N_15501,N_14025);
nor U23678 (N_23678,N_13649,N_13758);
and U23679 (N_23679,N_17321,N_16652);
xnor U23680 (N_23680,N_17067,N_17888);
nor U23681 (N_23681,N_17895,N_15760);
nand U23682 (N_23682,N_14994,N_14869);
xnor U23683 (N_23683,N_17013,N_13605);
and U23684 (N_23684,N_13591,N_16213);
xnor U23685 (N_23685,N_16152,N_13355);
and U23686 (N_23686,N_17881,N_16496);
nand U23687 (N_23687,N_17659,N_16524);
nor U23688 (N_23688,N_17138,N_14416);
nor U23689 (N_23689,N_15136,N_17438);
xnor U23690 (N_23690,N_14373,N_14119);
xnor U23691 (N_23691,N_16759,N_18478);
xor U23692 (N_23692,N_17767,N_15160);
nand U23693 (N_23693,N_12827,N_14670);
xor U23694 (N_23694,N_14771,N_18348);
nor U23695 (N_23695,N_15682,N_14522);
or U23696 (N_23696,N_13796,N_14805);
or U23697 (N_23697,N_15176,N_12555);
nand U23698 (N_23698,N_15022,N_14852);
nor U23699 (N_23699,N_16303,N_16551);
and U23700 (N_23700,N_14879,N_18220);
xor U23701 (N_23701,N_15807,N_12686);
or U23702 (N_23702,N_16029,N_16445);
xnor U23703 (N_23703,N_12865,N_16392);
nand U23704 (N_23704,N_14409,N_13180);
nor U23705 (N_23705,N_15602,N_12735);
and U23706 (N_23706,N_16329,N_16835);
or U23707 (N_23707,N_14594,N_15749);
xor U23708 (N_23708,N_14677,N_12740);
or U23709 (N_23709,N_13906,N_17482);
and U23710 (N_23710,N_14438,N_17694);
or U23711 (N_23711,N_13836,N_12702);
or U23712 (N_23712,N_13801,N_15136);
or U23713 (N_23713,N_14739,N_15056);
nor U23714 (N_23714,N_18457,N_14113);
xnor U23715 (N_23715,N_18272,N_15493);
xnor U23716 (N_23716,N_12701,N_15255);
and U23717 (N_23717,N_18283,N_12980);
nand U23718 (N_23718,N_18209,N_18614);
xor U23719 (N_23719,N_13921,N_17013);
or U23720 (N_23720,N_15745,N_16888);
nor U23721 (N_23721,N_14308,N_12546);
or U23722 (N_23722,N_18280,N_14790);
or U23723 (N_23723,N_16491,N_16414);
or U23724 (N_23724,N_18588,N_18360);
or U23725 (N_23725,N_18617,N_17438);
xor U23726 (N_23726,N_16043,N_17337);
and U23727 (N_23727,N_12555,N_18652);
xnor U23728 (N_23728,N_15460,N_17414);
and U23729 (N_23729,N_17042,N_17201);
or U23730 (N_23730,N_14017,N_12775);
nand U23731 (N_23731,N_17624,N_13818);
xor U23732 (N_23732,N_14793,N_17293);
nand U23733 (N_23733,N_15759,N_17968);
or U23734 (N_23734,N_14980,N_15180);
and U23735 (N_23735,N_16680,N_18011);
or U23736 (N_23736,N_14034,N_15560);
nand U23737 (N_23737,N_13364,N_14376);
or U23738 (N_23738,N_17345,N_16159);
or U23739 (N_23739,N_14276,N_14582);
nand U23740 (N_23740,N_13156,N_17482);
and U23741 (N_23741,N_17888,N_12889);
xnor U23742 (N_23742,N_16436,N_18331);
or U23743 (N_23743,N_13103,N_18305);
nand U23744 (N_23744,N_18071,N_15686);
nor U23745 (N_23745,N_14757,N_16608);
and U23746 (N_23746,N_14454,N_12699);
or U23747 (N_23747,N_15928,N_18461);
nand U23748 (N_23748,N_14691,N_13930);
or U23749 (N_23749,N_13100,N_15112);
xor U23750 (N_23750,N_12907,N_15438);
nor U23751 (N_23751,N_15382,N_14458);
nand U23752 (N_23752,N_17262,N_17038);
xnor U23753 (N_23753,N_16757,N_16498);
nor U23754 (N_23754,N_18081,N_14865);
nor U23755 (N_23755,N_13712,N_13760);
nand U23756 (N_23756,N_14906,N_18428);
or U23757 (N_23757,N_12639,N_14087);
and U23758 (N_23758,N_15226,N_12585);
nor U23759 (N_23759,N_18065,N_12823);
and U23760 (N_23760,N_17370,N_14192);
nor U23761 (N_23761,N_17813,N_16450);
xnor U23762 (N_23762,N_17324,N_15901);
nor U23763 (N_23763,N_13866,N_14449);
or U23764 (N_23764,N_14200,N_16549);
or U23765 (N_23765,N_12537,N_16674);
nor U23766 (N_23766,N_14411,N_16783);
nand U23767 (N_23767,N_18414,N_16175);
and U23768 (N_23768,N_18498,N_15092);
nand U23769 (N_23769,N_12550,N_14085);
or U23770 (N_23770,N_13263,N_17116);
and U23771 (N_23771,N_18656,N_18528);
or U23772 (N_23772,N_18202,N_16990);
nor U23773 (N_23773,N_15292,N_14743);
xor U23774 (N_23774,N_12975,N_18359);
xnor U23775 (N_23775,N_14315,N_16190);
xnor U23776 (N_23776,N_14780,N_18539);
nor U23777 (N_23777,N_16360,N_15329);
xor U23778 (N_23778,N_13738,N_16438);
nor U23779 (N_23779,N_14806,N_16791);
nor U23780 (N_23780,N_12914,N_15561);
and U23781 (N_23781,N_14458,N_14873);
and U23782 (N_23782,N_12613,N_13307);
xnor U23783 (N_23783,N_13123,N_18584);
xor U23784 (N_23784,N_17187,N_13182);
and U23785 (N_23785,N_16992,N_14725);
or U23786 (N_23786,N_18483,N_17683);
or U23787 (N_23787,N_18482,N_14158);
xor U23788 (N_23788,N_16179,N_14220);
xor U23789 (N_23789,N_18654,N_13825);
nor U23790 (N_23790,N_18534,N_16311);
xnor U23791 (N_23791,N_13770,N_16916);
nor U23792 (N_23792,N_16065,N_13889);
or U23793 (N_23793,N_16821,N_12595);
and U23794 (N_23794,N_12756,N_17760);
nand U23795 (N_23795,N_16314,N_16217);
or U23796 (N_23796,N_12813,N_12583);
nand U23797 (N_23797,N_15829,N_16877);
xor U23798 (N_23798,N_17407,N_16488);
and U23799 (N_23799,N_18641,N_16442);
or U23800 (N_23800,N_17875,N_17516);
nand U23801 (N_23801,N_16880,N_17293);
nand U23802 (N_23802,N_12663,N_18216);
nand U23803 (N_23803,N_15931,N_15527);
nor U23804 (N_23804,N_15945,N_17433);
and U23805 (N_23805,N_14855,N_15744);
and U23806 (N_23806,N_13637,N_13615);
and U23807 (N_23807,N_14525,N_12652);
and U23808 (N_23808,N_14855,N_18457);
or U23809 (N_23809,N_18169,N_14609);
xnor U23810 (N_23810,N_16846,N_16941);
or U23811 (N_23811,N_16221,N_15472);
or U23812 (N_23812,N_18743,N_12643);
xnor U23813 (N_23813,N_17115,N_14974);
nor U23814 (N_23814,N_13542,N_17748);
nor U23815 (N_23815,N_14717,N_15236);
or U23816 (N_23816,N_16259,N_16198);
nor U23817 (N_23817,N_13124,N_13714);
and U23818 (N_23818,N_14770,N_13856);
and U23819 (N_23819,N_13231,N_16098);
xor U23820 (N_23820,N_14848,N_18587);
xnor U23821 (N_23821,N_16261,N_14782);
nand U23822 (N_23822,N_16353,N_17219);
nor U23823 (N_23823,N_16851,N_13590);
nor U23824 (N_23824,N_16906,N_17451);
xnor U23825 (N_23825,N_18081,N_16202);
nand U23826 (N_23826,N_17575,N_16539);
nand U23827 (N_23827,N_14772,N_17263);
nor U23828 (N_23828,N_14566,N_13917);
xnor U23829 (N_23829,N_15728,N_18523);
nor U23830 (N_23830,N_15612,N_16305);
and U23831 (N_23831,N_16702,N_13473);
and U23832 (N_23832,N_13713,N_13967);
nand U23833 (N_23833,N_16341,N_12617);
and U23834 (N_23834,N_14515,N_16181);
nor U23835 (N_23835,N_16511,N_14727);
xor U23836 (N_23836,N_14614,N_18069);
nor U23837 (N_23837,N_13652,N_13095);
xor U23838 (N_23838,N_17745,N_18193);
xnor U23839 (N_23839,N_17857,N_18078);
nand U23840 (N_23840,N_17676,N_16438);
or U23841 (N_23841,N_13368,N_18713);
or U23842 (N_23842,N_15117,N_17722);
and U23843 (N_23843,N_15253,N_12912);
and U23844 (N_23844,N_12699,N_17934);
xor U23845 (N_23845,N_12561,N_15096);
and U23846 (N_23846,N_13891,N_13700);
nor U23847 (N_23847,N_18359,N_17666);
xor U23848 (N_23848,N_18213,N_16616);
and U23849 (N_23849,N_16535,N_15969);
or U23850 (N_23850,N_15163,N_14107);
and U23851 (N_23851,N_16768,N_18555);
and U23852 (N_23852,N_17382,N_18367);
nor U23853 (N_23853,N_14084,N_17527);
xnor U23854 (N_23854,N_16398,N_15863);
nor U23855 (N_23855,N_16821,N_16324);
xnor U23856 (N_23856,N_12698,N_14285);
or U23857 (N_23857,N_18332,N_15223);
nand U23858 (N_23858,N_12792,N_13004);
nor U23859 (N_23859,N_16381,N_14438);
xnor U23860 (N_23860,N_16344,N_16740);
or U23861 (N_23861,N_12604,N_16275);
nor U23862 (N_23862,N_16831,N_17779);
xnor U23863 (N_23863,N_16694,N_18172);
or U23864 (N_23864,N_13933,N_15086);
and U23865 (N_23865,N_17472,N_14589);
nand U23866 (N_23866,N_17033,N_16197);
xnor U23867 (N_23867,N_18034,N_16102);
xor U23868 (N_23868,N_17310,N_17977);
and U23869 (N_23869,N_12961,N_13511);
nor U23870 (N_23870,N_15630,N_14725);
or U23871 (N_23871,N_14326,N_13402);
nor U23872 (N_23872,N_12601,N_13726);
and U23873 (N_23873,N_14456,N_14213);
nor U23874 (N_23874,N_16823,N_17566);
nor U23875 (N_23875,N_16641,N_13698);
xnor U23876 (N_23876,N_17509,N_13000);
nor U23877 (N_23877,N_15079,N_14618);
xor U23878 (N_23878,N_14694,N_12990);
xor U23879 (N_23879,N_17566,N_14380);
xnor U23880 (N_23880,N_15996,N_13534);
and U23881 (N_23881,N_17997,N_15050);
nor U23882 (N_23882,N_14598,N_17183);
and U23883 (N_23883,N_13335,N_17648);
nor U23884 (N_23884,N_17253,N_16888);
xor U23885 (N_23885,N_15002,N_15457);
xnor U23886 (N_23886,N_15563,N_13150);
and U23887 (N_23887,N_16669,N_13714);
xor U23888 (N_23888,N_17714,N_16339);
and U23889 (N_23889,N_13788,N_15173);
xnor U23890 (N_23890,N_12751,N_16379);
nor U23891 (N_23891,N_17786,N_15726);
and U23892 (N_23892,N_16443,N_15974);
nor U23893 (N_23893,N_14088,N_13095);
xor U23894 (N_23894,N_13783,N_17097);
nor U23895 (N_23895,N_13893,N_15986);
nand U23896 (N_23896,N_16330,N_17203);
nor U23897 (N_23897,N_13932,N_13561);
nor U23898 (N_23898,N_12595,N_13628);
nor U23899 (N_23899,N_16265,N_18073);
and U23900 (N_23900,N_17433,N_13572);
nand U23901 (N_23901,N_17138,N_15142);
or U23902 (N_23902,N_18587,N_17832);
and U23903 (N_23903,N_17078,N_14292);
or U23904 (N_23904,N_14536,N_15509);
nand U23905 (N_23905,N_13652,N_13138);
or U23906 (N_23906,N_17669,N_18074);
xor U23907 (N_23907,N_18302,N_15944);
nor U23908 (N_23908,N_12918,N_17001);
nor U23909 (N_23909,N_15429,N_13751);
or U23910 (N_23910,N_14854,N_16741);
and U23911 (N_23911,N_13162,N_18677);
xnor U23912 (N_23912,N_13116,N_13386);
or U23913 (N_23913,N_16860,N_16131);
and U23914 (N_23914,N_12734,N_15182);
and U23915 (N_23915,N_16807,N_15157);
or U23916 (N_23916,N_18479,N_17492);
and U23917 (N_23917,N_16568,N_17796);
nand U23918 (N_23918,N_16510,N_18108);
nor U23919 (N_23919,N_13025,N_17198);
nand U23920 (N_23920,N_13893,N_12909);
xnor U23921 (N_23921,N_16424,N_13962);
and U23922 (N_23922,N_18679,N_17169);
xor U23923 (N_23923,N_14857,N_14986);
or U23924 (N_23924,N_13375,N_16556);
nand U23925 (N_23925,N_13533,N_18675);
nor U23926 (N_23926,N_14665,N_14508);
nor U23927 (N_23927,N_12903,N_16770);
xnor U23928 (N_23928,N_18321,N_17707);
nor U23929 (N_23929,N_14514,N_13458);
xor U23930 (N_23930,N_13753,N_12527);
xnor U23931 (N_23931,N_12860,N_13321);
and U23932 (N_23932,N_16171,N_18601);
nand U23933 (N_23933,N_15527,N_17554);
nand U23934 (N_23934,N_16701,N_15056);
nor U23935 (N_23935,N_16079,N_13112);
nand U23936 (N_23936,N_14097,N_16207);
nor U23937 (N_23937,N_16114,N_15092);
nand U23938 (N_23938,N_13044,N_17497);
nand U23939 (N_23939,N_14329,N_16178);
nand U23940 (N_23940,N_13594,N_14364);
nand U23941 (N_23941,N_16202,N_17373);
and U23942 (N_23942,N_18718,N_14456);
nor U23943 (N_23943,N_17005,N_13149);
or U23944 (N_23944,N_13181,N_16137);
xor U23945 (N_23945,N_12636,N_13053);
or U23946 (N_23946,N_15859,N_16479);
and U23947 (N_23947,N_14647,N_13871);
or U23948 (N_23948,N_14545,N_16515);
nor U23949 (N_23949,N_16729,N_17473);
nand U23950 (N_23950,N_14917,N_18018);
and U23951 (N_23951,N_13059,N_18424);
xor U23952 (N_23952,N_18317,N_16047);
xnor U23953 (N_23953,N_15620,N_14079);
nand U23954 (N_23954,N_16663,N_15220);
xor U23955 (N_23955,N_16337,N_17131);
xor U23956 (N_23956,N_18608,N_16018);
or U23957 (N_23957,N_14814,N_15217);
nand U23958 (N_23958,N_14696,N_15392);
nand U23959 (N_23959,N_16974,N_13838);
nand U23960 (N_23960,N_12739,N_18008);
nand U23961 (N_23961,N_14738,N_17950);
or U23962 (N_23962,N_15005,N_13140);
and U23963 (N_23963,N_16554,N_18177);
nand U23964 (N_23964,N_17820,N_17282);
and U23965 (N_23965,N_14129,N_15475);
or U23966 (N_23966,N_17286,N_14916);
or U23967 (N_23967,N_13659,N_17112);
nand U23968 (N_23968,N_14054,N_17906);
and U23969 (N_23969,N_15811,N_16707);
nor U23970 (N_23970,N_14312,N_18148);
nand U23971 (N_23971,N_17898,N_16066);
xnor U23972 (N_23972,N_15239,N_16235);
nand U23973 (N_23973,N_15752,N_13462);
nand U23974 (N_23974,N_15599,N_18719);
or U23975 (N_23975,N_13657,N_17760);
nor U23976 (N_23976,N_14419,N_15057);
and U23977 (N_23977,N_18184,N_16318);
xor U23978 (N_23978,N_18618,N_13558);
xnor U23979 (N_23979,N_18101,N_14108);
xor U23980 (N_23980,N_18611,N_12710);
xnor U23981 (N_23981,N_17360,N_17060);
nor U23982 (N_23982,N_14658,N_17334);
nor U23983 (N_23983,N_15149,N_16149);
nor U23984 (N_23984,N_15397,N_13630);
or U23985 (N_23985,N_16699,N_14409);
nand U23986 (N_23986,N_16526,N_17112);
nor U23987 (N_23987,N_18522,N_16419);
nand U23988 (N_23988,N_15827,N_16486);
nand U23989 (N_23989,N_14896,N_16904);
or U23990 (N_23990,N_15375,N_14480);
nor U23991 (N_23991,N_16188,N_15680);
nor U23992 (N_23992,N_17651,N_13880);
nor U23993 (N_23993,N_15501,N_12796);
xnor U23994 (N_23994,N_15077,N_12986);
nand U23995 (N_23995,N_13720,N_16448);
or U23996 (N_23996,N_15640,N_16432);
or U23997 (N_23997,N_17964,N_16010);
xor U23998 (N_23998,N_13600,N_16562);
nor U23999 (N_23999,N_13376,N_15767);
and U24000 (N_24000,N_17039,N_12795);
or U24001 (N_24001,N_14504,N_16227);
or U24002 (N_24002,N_14257,N_17023);
nand U24003 (N_24003,N_18254,N_16180);
nand U24004 (N_24004,N_12865,N_16851);
and U24005 (N_24005,N_17156,N_18464);
xnor U24006 (N_24006,N_18474,N_15692);
nand U24007 (N_24007,N_12588,N_14955);
nand U24008 (N_24008,N_18725,N_13545);
nor U24009 (N_24009,N_14045,N_12724);
nor U24010 (N_24010,N_12661,N_15458);
nand U24011 (N_24011,N_18126,N_14190);
xnor U24012 (N_24012,N_16160,N_16021);
or U24013 (N_24013,N_17536,N_18727);
and U24014 (N_24014,N_17950,N_15983);
xor U24015 (N_24015,N_14672,N_17811);
nand U24016 (N_24016,N_16043,N_14047);
nand U24017 (N_24017,N_13787,N_18345);
xnor U24018 (N_24018,N_18655,N_12534);
xnor U24019 (N_24019,N_15420,N_15116);
and U24020 (N_24020,N_16140,N_18368);
and U24021 (N_24021,N_17098,N_12871);
nand U24022 (N_24022,N_16618,N_18103);
or U24023 (N_24023,N_18325,N_17474);
and U24024 (N_24024,N_12811,N_13178);
and U24025 (N_24025,N_16174,N_14235);
xor U24026 (N_24026,N_13520,N_14970);
nor U24027 (N_24027,N_15560,N_18402);
xor U24028 (N_24028,N_13031,N_14188);
nor U24029 (N_24029,N_14136,N_13263);
or U24030 (N_24030,N_17115,N_14153);
xor U24031 (N_24031,N_15980,N_16471);
or U24032 (N_24032,N_14284,N_14493);
and U24033 (N_24033,N_16328,N_13154);
or U24034 (N_24034,N_16177,N_13268);
or U24035 (N_24035,N_13412,N_14752);
xor U24036 (N_24036,N_17512,N_15087);
nor U24037 (N_24037,N_17902,N_18538);
or U24038 (N_24038,N_15729,N_16177);
or U24039 (N_24039,N_17380,N_13202);
nand U24040 (N_24040,N_17806,N_16194);
xor U24041 (N_24041,N_14486,N_14215);
xnor U24042 (N_24042,N_15723,N_14818);
xnor U24043 (N_24043,N_14951,N_14268);
nand U24044 (N_24044,N_13821,N_17029);
nor U24045 (N_24045,N_13538,N_14419);
and U24046 (N_24046,N_16966,N_18039);
nand U24047 (N_24047,N_18396,N_14032);
xnor U24048 (N_24048,N_13076,N_15972);
nor U24049 (N_24049,N_14711,N_13640);
nor U24050 (N_24050,N_18059,N_12838);
or U24051 (N_24051,N_14094,N_13151);
nor U24052 (N_24052,N_17035,N_14972);
nor U24053 (N_24053,N_14144,N_14396);
xnor U24054 (N_24054,N_14098,N_14613);
nand U24055 (N_24055,N_14996,N_14298);
xnor U24056 (N_24056,N_13466,N_17145);
nand U24057 (N_24057,N_15872,N_13895);
nor U24058 (N_24058,N_12634,N_14898);
and U24059 (N_24059,N_12896,N_12774);
nor U24060 (N_24060,N_15715,N_16693);
nor U24061 (N_24061,N_15980,N_17000);
nor U24062 (N_24062,N_17803,N_16150);
nand U24063 (N_24063,N_14760,N_17310);
xnor U24064 (N_24064,N_16415,N_14306);
and U24065 (N_24065,N_12559,N_12813);
and U24066 (N_24066,N_18381,N_18166);
nor U24067 (N_24067,N_13130,N_14487);
nand U24068 (N_24068,N_15620,N_13256);
xnor U24069 (N_24069,N_14712,N_15956);
or U24070 (N_24070,N_16636,N_14797);
nand U24071 (N_24071,N_12928,N_17510);
or U24072 (N_24072,N_18591,N_17849);
xor U24073 (N_24073,N_13120,N_18593);
xnor U24074 (N_24074,N_17369,N_12560);
nand U24075 (N_24075,N_14277,N_12806);
or U24076 (N_24076,N_13569,N_18074);
xnor U24077 (N_24077,N_15156,N_15327);
nor U24078 (N_24078,N_15767,N_14720);
nand U24079 (N_24079,N_18065,N_16708);
xnor U24080 (N_24080,N_17827,N_18184);
xnor U24081 (N_24081,N_17026,N_14516);
or U24082 (N_24082,N_14841,N_14355);
or U24083 (N_24083,N_15930,N_16945);
xor U24084 (N_24084,N_18739,N_18126);
or U24085 (N_24085,N_16230,N_12584);
and U24086 (N_24086,N_13941,N_16229);
and U24087 (N_24087,N_13752,N_15047);
and U24088 (N_24088,N_18323,N_16245);
and U24089 (N_24089,N_17046,N_14153);
xnor U24090 (N_24090,N_13460,N_13225);
or U24091 (N_24091,N_17930,N_17277);
or U24092 (N_24092,N_12634,N_14345);
or U24093 (N_24093,N_18423,N_15796);
nand U24094 (N_24094,N_13559,N_13741);
and U24095 (N_24095,N_13961,N_18346);
nand U24096 (N_24096,N_16944,N_17061);
xor U24097 (N_24097,N_16152,N_13104);
nand U24098 (N_24098,N_17558,N_18088);
nand U24099 (N_24099,N_16541,N_16846);
xnor U24100 (N_24100,N_14153,N_15318);
and U24101 (N_24101,N_16217,N_15252);
nor U24102 (N_24102,N_12770,N_12551);
nor U24103 (N_24103,N_17663,N_17993);
and U24104 (N_24104,N_17898,N_17085);
and U24105 (N_24105,N_13258,N_15161);
xor U24106 (N_24106,N_17856,N_18314);
xor U24107 (N_24107,N_13432,N_13216);
nand U24108 (N_24108,N_17484,N_18665);
xor U24109 (N_24109,N_15944,N_16710);
or U24110 (N_24110,N_14811,N_18423);
xor U24111 (N_24111,N_17891,N_13491);
nor U24112 (N_24112,N_12774,N_16579);
nor U24113 (N_24113,N_18077,N_18071);
nor U24114 (N_24114,N_15673,N_17654);
xor U24115 (N_24115,N_17661,N_16979);
or U24116 (N_24116,N_14101,N_15026);
xor U24117 (N_24117,N_18246,N_14898);
nor U24118 (N_24118,N_12552,N_12943);
or U24119 (N_24119,N_17667,N_14158);
and U24120 (N_24120,N_18672,N_17449);
and U24121 (N_24121,N_16393,N_16361);
nor U24122 (N_24122,N_14617,N_15722);
xnor U24123 (N_24123,N_13805,N_13643);
or U24124 (N_24124,N_17610,N_18267);
xnor U24125 (N_24125,N_18679,N_12918);
xor U24126 (N_24126,N_18197,N_14299);
or U24127 (N_24127,N_16763,N_15869);
xor U24128 (N_24128,N_14091,N_12767);
or U24129 (N_24129,N_15586,N_14372);
or U24130 (N_24130,N_14267,N_13801);
or U24131 (N_24131,N_18333,N_15066);
or U24132 (N_24132,N_18020,N_17013);
and U24133 (N_24133,N_15998,N_16845);
nor U24134 (N_24134,N_14963,N_13218);
nor U24135 (N_24135,N_12609,N_16041);
xor U24136 (N_24136,N_13077,N_17799);
or U24137 (N_24137,N_16072,N_12555);
nand U24138 (N_24138,N_16947,N_17924);
or U24139 (N_24139,N_15699,N_17803);
nand U24140 (N_24140,N_16401,N_12534);
and U24141 (N_24141,N_16066,N_13732);
xnor U24142 (N_24142,N_12961,N_14991);
xor U24143 (N_24143,N_13373,N_16567);
xor U24144 (N_24144,N_16294,N_14861);
nand U24145 (N_24145,N_18181,N_15775);
nand U24146 (N_24146,N_14705,N_13261);
xor U24147 (N_24147,N_14688,N_15726);
and U24148 (N_24148,N_18192,N_14010);
and U24149 (N_24149,N_15538,N_13059);
nand U24150 (N_24150,N_12675,N_12833);
xnor U24151 (N_24151,N_15760,N_12814);
or U24152 (N_24152,N_14623,N_12929);
xnor U24153 (N_24153,N_18061,N_16608);
nor U24154 (N_24154,N_12799,N_13155);
nor U24155 (N_24155,N_14223,N_15596);
or U24156 (N_24156,N_14318,N_17019);
xor U24157 (N_24157,N_16119,N_14085);
or U24158 (N_24158,N_15566,N_15602);
nand U24159 (N_24159,N_17257,N_17219);
and U24160 (N_24160,N_16370,N_12676);
nand U24161 (N_24161,N_14310,N_15748);
nand U24162 (N_24162,N_15538,N_18345);
and U24163 (N_24163,N_15885,N_14952);
nand U24164 (N_24164,N_14091,N_18277);
and U24165 (N_24165,N_18531,N_15383);
or U24166 (N_24166,N_16008,N_18501);
or U24167 (N_24167,N_14913,N_16936);
or U24168 (N_24168,N_18267,N_15461);
xnor U24169 (N_24169,N_17828,N_16730);
xor U24170 (N_24170,N_12757,N_17814);
and U24171 (N_24171,N_12869,N_14747);
nor U24172 (N_24172,N_15962,N_14390);
xnor U24173 (N_24173,N_14678,N_14109);
nor U24174 (N_24174,N_15451,N_13251);
and U24175 (N_24175,N_16197,N_13919);
and U24176 (N_24176,N_18472,N_14028);
nand U24177 (N_24177,N_16540,N_18493);
or U24178 (N_24178,N_15131,N_15944);
and U24179 (N_24179,N_17588,N_18051);
and U24180 (N_24180,N_14248,N_18470);
nor U24181 (N_24181,N_16136,N_15418);
nor U24182 (N_24182,N_14505,N_16596);
or U24183 (N_24183,N_15982,N_15194);
nand U24184 (N_24184,N_14828,N_12786);
nand U24185 (N_24185,N_14255,N_14700);
nand U24186 (N_24186,N_16412,N_15714);
or U24187 (N_24187,N_13908,N_15080);
nor U24188 (N_24188,N_15757,N_14974);
xor U24189 (N_24189,N_15276,N_13659);
nor U24190 (N_24190,N_13926,N_17886);
or U24191 (N_24191,N_13351,N_12523);
nand U24192 (N_24192,N_15464,N_17477);
nand U24193 (N_24193,N_17068,N_18263);
nor U24194 (N_24194,N_14880,N_15644);
and U24195 (N_24195,N_13259,N_12663);
nor U24196 (N_24196,N_15314,N_12877);
or U24197 (N_24197,N_16489,N_15392);
and U24198 (N_24198,N_18478,N_14985);
nor U24199 (N_24199,N_13973,N_17620);
nand U24200 (N_24200,N_12864,N_14993);
or U24201 (N_24201,N_14110,N_15900);
and U24202 (N_24202,N_18290,N_12894);
nand U24203 (N_24203,N_18382,N_13364);
xnor U24204 (N_24204,N_17609,N_17355);
and U24205 (N_24205,N_12874,N_14314);
nor U24206 (N_24206,N_13292,N_15225);
or U24207 (N_24207,N_13284,N_17808);
xor U24208 (N_24208,N_18235,N_17185);
or U24209 (N_24209,N_14886,N_15511);
and U24210 (N_24210,N_12519,N_13063);
or U24211 (N_24211,N_16986,N_15504);
xor U24212 (N_24212,N_17699,N_15070);
xor U24213 (N_24213,N_12514,N_14004);
nand U24214 (N_24214,N_12836,N_17746);
or U24215 (N_24215,N_16095,N_13322);
nand U24216 (N_24216,N_14048,N_14157);
xor U24217 (N_24217,N_12528,N_13693);
nor U24218 (N_24218,N_17499,N_17999);
or U24219 (N_24219,N_16863,N_12914);
and U24220 (N_24220,N_14360,N_15904);
or U24221 (N_24221,N_18016,N_16422);
and U24222 (N_24222,N_17671,N_13636);
or U24223 (N_24223,N_15945,N_13252);
xor U24224 (N_24224,N_17484,N_15963);
and U24225 (N_24225,N_15335,N_16937);
and U24226 (N_24226,N_13564,N_14146);
or U24227 (N_24227,N_16492,N_17270);
nor U24228 (N_24228,N_15897,N_12781);
nand U24229 (N_24229,N_17804,N_14997);
nand U24230 (N_24230,N_16419,N_18547);
nand U24231 (N_24231,N_16050,N_13774);
and U24232 (N_24232,N_14109,N_13702);
and U24233 (N_24233,N_17739,N_13102);
nand U24234 (N_24234,N_16582,N_17792);
xor U24235 (N_24235,N_13797,N_15092);
and U24236 (N_24236,N_13608,N_17314);
and U24237 (N_24237,N_18554,N_13287);
nand U24238 (N_24238,N_13918,N_18036);
nand U24239 (N_24239,N_15531,N_15949);
nand U24240 (N_24240,N_17071,N_16097);
and U24241 (N_24241,N_16891,N_13117);
xor U24242 (N_24242,N_15926,N_13247);
or U24243 (N_24243,N_13012,N_13741);
xnor U24244 (N_24244,N_16375,N_13261);
nor U24245 (N_24245,N_14282,N_13884);
and U24246 (N_24246,N_13930,N_18004);
xnor U24247 (N_24247,N_12544,N_13268);
and U24248 (N_24248,N_14460,N_17078);
and U24249 (N_24249,N_16310,N_12856);
nor U24250 (N_24250,N_17486,N_18658);
xor U24251 (N_24251,N_17940,N_16482);
xnor U24252 (N_24252,N_15668,N_13325);
nand U24253 (N_24253,N_13997,N_17812);
and U24254 (N_24254,N_17737,N_17406);
nand U24255 (N_24255,N_14939,N_13646);
xor U24256 (N_24256,N_13629,N_17704);
or U24257 (N_24257,N_17355,N_12843);
and U24258 (N_24258,N_13143,N_15505);
nand U24259 (N_24259,N_16896,N_16995);
nand U24260 (N_24260,N_14438,N_16646);
nand U24261 (N_24261,N_16974,N_17759);
nand U24262 (N_24262,N_18633,N_16390);
xnor U24263 (N_24263,N_17248,N_18655);
or U24264 (N_24264,N_12762,N_15645);
nand U24265 (N_24265,N_17212,N_18133);
nand U24266 (N_24266,N_15425,N_16972);
xnor U24267 (N_24267,N_13068,N_18295);
nor U24268 (N_24268,N_15265,N_16620);
xnor U24269 (N_24269,N_14470,N_15901);
nand U24270 (N_24270,N_15521,N_15478);
nand U24271 (N_24271,N_18312,N_17634);
nor U24272 (N_24272,N_16321,N_17523);
nor U24273 (N_24273,N_18529,N_13536);
or U24274 (N_24274,N_18065,N_17937);
nand U24275 (N_24275,N_18514,N_15983);
xor U24276 (N_24276,N_16487,N_17942);
nand U24277 (N_24277,N_16943,N_17130);
and U24278 (N_24278,N_17741,N_15113);
nor U24279 (N_24279,N_12528,N_17714);
nor U24280 (N_24280,N_14331,N_14175);
and U24281 (N_24281,N_16987,N_13088);
xor U24282 (N_24282,N_18521,N_14378);
nor U24283 (N_24283,N_12754,N_12881);
xnor U24284 (N_24284,N_17357,N_17686);
xor U24285 (N_24285,N_14636,N_16442);
or U24286 (N_24286,N_18503,N_14088);
nand U24287 (N_24287,N_16384,N_15104);
or U24288 (N_24288,N_13478,N_15211);
nand U24289 (N_24289,N_12535,N_17071);
xor U24290 (N_24290,N_13411,N_16966);
or U24291 (N_24291,N_17125,N_14251);
xnor U24292 (N_24292,N_15089,N_16307);
xnor U24293 (N_24293,N_14428,N_16782);
and U24294 (N_24294,N_17863,N_14636);
and U24295 (N_24295,N_16144,N_17948);
or U24296 (N_24296,N_14804,N_16955);
nor U24297 (N_24297,N_18156,N_14290);
nor U24298 (N_24298,N_18160,N_17282);
and U24299 (N_24299,N_18605,N_12774);
or U24300 (N_24300,N_13780,N_15360);
and U24301 (N_24301,N_12865,N_14806);
and U24302 (N_24302,N_15334,N_13725);
xnor U24303 (N_24303,N_14590,N_14076);
or U24304 (N_24304,N_15204,N_18521);
or U24305 (N_24305,N_15863,N_13887);
or U24306 (N_24306,N_12649,N_15737);
or U24307 (N_24307,N_16473,N_16933);
nand U24308 (N_24308,N_17651,N_17151);
xnor U24309 (N_24309,N_17032,N_14067);
nand U24310 (N_24310,N_14205,N_14494);
nor U24311 (N_24311,N_16311,N_13517);
nor U24312 (N_24312,N_16177,N_15635);
and U24313 (N_24313,N_12707,N_13501);
or U24314 (N_24314,N_14427,N_15938);
nand U24315 (N_24315,N_16088,N_17973);
nor U24316 (N_24316,N_18747,N_15579);
or U24317 (N_24317,N_16561,N_15773);
xor U24318 (N_24318,N_15618,N_13800);
nand U24319 (N_24319,N_13295,N_17267);
xnor U24320 (N_24320,N_14406,N_14974);
and U24321 (N_24321,N_17330,N_16964);
nor U24322 (N_24322,N_16790,N_13502);
nand U24323 (N_24323,N_13618,N_17416);
nand U24324 (N_24324,N_16414,N_15003);
nor U24325 (N_24325,N_15449,N_18141);
and U24326 (N_24326,N_15242,N_16262);
nand U24327 (N_24327,N_15176,N_14216);
nand U24328 (N_24328,N_14174,N_16454);
xnor U24329 (N_24329,N_17266,N_14649);
nor U24330 (N_24330,N_16267,N_12878);
xnor U24331 (N_24331,N_15696,N_12827);
nand U24332 (N_24332,N_13397,N_14945);
and U24333 (N_24333,N_14220,N_17611);
nand U24334 (N_24334,N_18416,N_13443);
nand U24335 (N_24335,N_13668,N_18736);
nand U24336 (N_24336,N_16812,N_15334);
nand U24337 (N_24337,N_14675,N_13001);
nor U24338 (N_24338,N_13183,N_14245);
xor U24339 (N_24339,N_17157,N_14899);
nand U24340 (N_24340,N_13789,N_17504);
or U24341 (N_24341,N_14863,N_17403);
xnor U24342 (N_24342,N_18008,N_13990);
or U24343 (N_24343,N_17211,N_17823);
or U24344 (N_24344,N_14160,N_16336);
and U24345 (N_24345,N_18157,N_17540);
xor U24346 (N_24346,N_16112,N_18245);
xnor U24347 (N_24347,N_13414,N_15930);
and U24348 (N_24348,N_14987,N_15941);
nand U24349 (N_24349,N_18382,N_13799);
or U24350 (N_24350,N_14923,N_13245);
nor U24351 (N_24351,N_12800,N_13521);
xor U24352 (N_24352,N_15538,N_16675);
or U24353 (N_24353,N_17777,N_13022);
or U24354 (N_24354,N_16951,N_14093);
xor U24355 (N_24355,N_14077,N_16662);
and U24356 (N_24356,N_13113,N_13272);
or U24357 (N_24357,N_16917,N_15260);
nor U24358 (N_24358,N_16753,N_17102);
xor U24359 (N_24359,N_14961,N_18233);
or U24360 (N_24360,N_15251,N_14507);
xnor U24361 (N_24361,N_18741,N_13733);
or U24362 (N_24362,N_16214,N_14679);
nand U24363 (N_24363,N_17062,N_15817);
nand U24364 (N_24364,N_12761,N_14212);
xnor U24365 (N_24365,N_18286,N_13194);
nor U24366 (N_24366,N_15223,N_14810);
xor U24367 (N_24367,N_14074,N_15269);
xnor U24368 (N_24368,N_15515,N_13436);
and U24369 (N_24369,N_18677,N_13020);
and U24370 (N_24370,N_12580,N_14906);
nor U24371 (N_24371,N_15093,N_13760);
nand U24372 (N_24372,N_12854,N_13790);
and U24373 (N_24373,N_15202,N_13343);
xnor U24374 (N_24374,N_15680,N_14354);
nor U24375 (N_24375,N_16280,N_16194);
and U24376 (N_24376,N_17380,N_15610);
or U24377 (N_24377,N_13082,N_17800);
xor U24378 (N_24378,N_17187,N_16910);
and U24379 (N_24379,N_13081,N_13916);
nand U24380 (N_24380,N_16053,N_16462);
or U24381 (N_24381,N_18499,N_14528);
and U24382 (N_24382,N_14270,N_14024);
and U24383 (N_24383,N_13703,N_14305);
nor U24384 (N_24384,N_18074,N_16766);
or U24385 (N_24385,N_13654,N_17828);
and U24386 (N_24386,N_15103,N_14628);
nand U24387 (N_24387,N_15803,N_13038);
xor U24388 (N_24388,N_17005,N_13628);
nand U24389 (N_24389,N_14253,N_13879);
nor U24390 (N_24390,N_15121,N_15676);
or U24391 (N_24391,N_12865,N_15154);
nand U24392 (N_24392,N_12992,N_12905);
or U24393 (N_24393,N_17066,N_17469);
nand U24394 (N_24394,N_13131,N_12829);
and U24395 (N_24395,N_14264,N_18487);
xnor U24396 (N_24396,N_14838,N_12517);
or U24397 (N_24397,N_13980,N_14757);
nand U24398 (N_24398,N_15858,N_18147);
xnor U24399 (N_24399,N_17879,N_18087);
or U24400 (N_24400,N_17148,N_17056);
or U24401 (N_24401,N_16032,N_17605);
or U24402 (N_24402,N_17761,N_17496);
xor U24403 (N_24403,N_14357,N_13319);
and U24404 (N_24404,N_18586,N_17834);
xnor U24405 (N_24405,N_14203,N_17757);
or U24406 (N_24406,N_18511,N_16797);
or U24407 (N_24407,N_14490,N_15676);
or U24408 (N_24408,N_16638,N_16148);
nand U24409 (N_24409,N_13122,N_15457);
xor U24410 (N_24410,N_16482,N_13347);
or U24411 (N_24411,N_16057,N_14592);
and U24412 (N_24412,N_13346,N_15055);
nand U24413 (N_24413,N_18704,N_17097);
or U24414 (N_24414,N_16053,N_16578);
xor U24415 (N_24415,N_12975,N_14396);
and U24416 (N_24416,N_17624,N_16015);
or U24417 (N_24417,N_15753,N_12947);
xor U24418 (N_24418,N_17773,N_16144);
xnor U24419 (N_24419,N_14167,N_17991);
nor U24420 (N_24420,N_12586,N_13418);
and U24421 (N_24421,N_17494,N_17336);
nand U24422 (N_24422,N_17243,N_15373);
nand U24423 (N_24423,N_13850,N_15551);
nand U24424 (N_24424,N_17324,N_12736);
or U24425 (N_24425,N_14254,N_15517);
xor U24426 (N_24426,N_14960,N_15364);
or U24427 (N_24427,N_14391,N_18381);
nand U24428 (N_24428,N_15255,N_15135);
and U24429 (N_24429,N_16971,N_13093);
or U24430 (N_24430,N_17997,N_17635);
xnor U24431 (N_24431,N_18147,N_18207);
nor U24432 (N_24432,N_17538,N_13033);
nor U24433 (N_24433,N_16406,N_17658);
xor U24434 (N_24434,N_14267,N_17049);
nor U24435 (N_24435,N_14160,N_13650);
or U24436 (N_24436,N_15547,N_15229);
nor U24437 (N_24437,N_16466,N_18672);
or U24438 (N_24438,N_14266,N_16528);
nor U24439 (N_24439,N_15491,N_18391);
xnor U24440 (N_24440,N_12679,N_13290);
nand U24441 (N_24441,N_14208,N_15945);
or U24442 (N_24442,N_15102,N_18715);
nor U24443 (N_24443,N_17219,N_13876);
or U24444 (N_24444,N_14594,N_15088);
or U24445 (N_24445,N_13197,N_15839);
nand U24446 (N_24446,N_15393,N_13895);
nand U24447 (N_24447,N_17711,N_13913);
and U24448 (N_24448,N_17286,N_13568);
and U24449 (N_24449,N_17648,N_14483);
nand U24450 (N_24450,N_15555,N_17267);
and U24451 (N_24451,N_16226,N_17131);
nor U24452 (N_24452,N_12895,N_13350);
xor U24453 (N_24453,N_14986,N_18534);
and U24454 (N_24454,N_18096,N_14989);
or U24455 (N_24455,N_18259,N_12931);
xor U24456 (N_24456,N_15108,N_13658);
or U24457 (N_24457,N_17116,N_17179);
nand U24458 (N_24458,N_15288,N_13547);
and U24459 (N_24459,N_17513,N_17319);
xor U24460 (N_24460,N_15208,N_13858);
or U24461 (N_24461,N_16564,N_13885);
nor U24462 (N_24462,N_15659,N_18616);
and U24463 (N_24463,N_16270,N_13352);
nand U24464 (N_24464,N_15860,N_18251);
xor U24465 (N_24465,N_17641,N_16338);
nor U24466 (N_24466,N_15252,N_14150);
nor U24467 (N_24467,N_18462,N_12948);
xor U24468 (N_24468,N_15512,N_13551);
nor U24469 (N_24469,N_13470,N_17016);
nand U24470 (N_24470,N_12922,N_16179);
xor U24471 (N_24471,N_15370,N_13662);
xor U24472 (N_24472,N_16997,N_16509);
or U24473 (N_24473,N_17316,N_12973);
nor U24474 (N_24474,N_16009,N_12563);
nor U24475 (N_24475,N_18508,N_12901);
or U24476 (N_24476,N_15316,N_17976);
nor U24477 (N_24477,N_18717,N_17827);
and U24478 (N_24478,N_13804,N_18384);
or U24479 (N_24479,N_18425,N_15625);
xor U24480 (N_24480,N_13794,N_14327);
xnor U24481 (N_24481,N_18742,N_15180);
and U24482 (N_24482,N_18128,N_13236);
xnor U24483 (N_24483,N_16494,N_15164);
nand U24484 (N_24484,N_14368,N_16335);
or U24485 (N_24485,N_14791,N_13194);
or U24486 (N_24486,N_14268,N_12593);
nor U24487 (N_24487,N_12921,N_15388);
and U24488 (N_24488,N_16004,N_17638);
nor U24489 (N_24489,N_12789,N_16502);
or U24490 (N_24490,N_17247,N_17942);
nor U24491 (N_24491,N_13292,N_15296);
nand U24492 (N_24492,N_14892,N_13678);
nand U24493 (N_24493,N_16836,N_17624);
nor U24494 (N_24494,N_17541,N_17689);
nor U24495 (N_24495,N_15612,N_16245);
xnor U24496 (N_24496,N_13983,N_12613);
nand U24497 (N_24497,N_15713,N_18638);
or U24498 (N_24498,N_14073,N_12589);
and U24499 (N_24499,N_15046,N_15356);
or U24500 (N_24500,N_17796,N_14245);
and U24501 (N_24501,N_12745,N_13226);
nand U24502 (N_24502,N_18152,N_16795);
nor U24503 (N_24503,N_16515,N_12616);
xor U24504 (N_24504,N_15109,N_17750);
nor U24505 (N_24505,N_16570,N_16154);
nor U24506 (N_24506,N_12626,N_14655);
xor U24507 (N_24507,N_17106,N_14287);
nand U24508 (N_24508,N_17749,N_16002);
and U24509 (N_24509,N_17470,N_15455);
or U24510 (N_24510,N_13412,N_12569);
nor U24511 (N_24511,N_18405,N_18486);
nand U24512 (N_24512,N_16093,N_13324);
or U24513 (N_24513,N_16057,N_12619);
xnor U24514 (N_24514,N_13793,N_18378);
or U24515 (N_24515,N_18208,N_18369);
nand U24516 (N_24516,N_14226,N_17922);
nor U24517 (N_24517,N_15242,N_13739);
and U24518 (N_24518,N_15991,N_14895);
nor U24519 (N_24519,N_17979,N_17325);
nand U24520 (N_24520,N_13627,N_13263);
and U24521 (N_24521,N_18161,N_17732);
and U24522 (N_24522,N_18147,N_14847);
and U24523 (N_24523,N_16517,N_16281);
nand U24524 (N_24524,N_15096,N_13880);
nor U24525 (N_24525,N_17215,N_15914);
xor U24526 (N_24526,N_16429,N_17883);
nand U24527 (N_24527,N_16637,N_18138);
and U24528 (N_24528,N_14818,N_13669);
nor U24529 (N_24529,N_12928,N_15805);
or U24530 (N_24530,N_13617,N_16013);
xor U24531 (N_24531,N_13326,N_17262);
nand U24532 (N_24532,N_12661,N_17798);
nand U24533 (N_24533,N_14113,N_18506);
nand U24534 (N_24534,N_17077,N_17848);
xnor U24535 (N_24535,N_14426,N_17972);
xnor U24536 (N_24536,N_16999,N_14795);
or U24537 (N_24537,N_18234,N_16863);
nand U24538 (N_24538,N_12948,N_15015);
nor U24539 (N_24539,N_16852,N_17655);
or U24540 (N_24540,N_17102,N_16462);
or U24541 (N_24541,N_15719,N_15450);
nand U24542 (N_24542,N_13710,N_14559);
nand U24543 (N_24543,N_16598,N_14145);
nor U24544 (N_24544,N_16516,N_16736);
and U24545 (N_24545,N_13251,N_13603);
nor U24546 (N_24546,N_14658,N_13214);
nor U24547 (N_24547,N_14682,N_13824);
nor U24548 (N_24548,N_16627,N_15436);
nor U24549 (N_24549,N_17729,N_15166);
nor U24550 (N_24550,N_18381,N_13578);
nor U24551 (N_24551,N_15533,N_12754);
nor U24552 (N_24552,N_16352,N_13470);
nor U24553 (N_24553,N_15777,N_15968);
and U24554 (N_24554,N_14459,N_12875);
and U24555 (N_24555,N_13846,N_18021);
xor U24556 (N_24556,N_17797,N_12758);
nand U24557 (N_24557,N_17543,N_17480);
nand U24558 (N_24558,N_12954,N_12838);
nor U24559 (N_24559,N_16340,N_15762);
nor U24560 (N_24560,N_13465,N_13371);
nor U24561 (N_24561,N_16996,N_13337);
xnor U24562 (N_24562,N_18130,N_16526);
xnor U24563 (N_24563,N_13603,N_14042);
nand U24564 (N_24564,N_18483,N_13000);
nor U24565 (N_24565,N_12677,N_17272);
and U24566 (N_24566,N_13513,N_14489);
xnor U24567 (N_24567,N_13290,N_15975);
and U24568 (N_24568,N_15385,N_14910);
nor U24569 (N_24569,N_15220,N_14234);
and U24570 (N_24570,N_14965,N_12892);
nor U24571 (N_24571,N_16396,N_12913);
or U24572 (N_24572,N_17267,N_15294);
or U24573 (N_24573,N_13742,N_14121);
or U24574 (N_24574,N_14714,N_17127);
or U24575 (N_24575,N_17590,N_18355);
xor U24576 (N_24576,N_17370,N_13475);
nor U24577 (N_24577,N_13772,N_17437);
and U24578 (N_24578,N_13854,N_12779);
nand U24579 (N_24579,N_13445,N_18678);
or U24580 (N_24580,N_14699,N_15894);
or U24581 (N_24581,N_15851,N_18375);
xor U24582 (N_24582,N_17867,N_18539);
nand U24583 (N_24583,N_15899,N_16895);
or U24584 (N_24584,N_15525,N_14613);
xor U24585 (N_24585,N_13162,N_14961);
or U24586 (N_24586,N_12780,N_16361);
xor U24587 (N_24587,N_12909,N_16626);
xor U24588 (N_24588,N_13577,N_16419);
xor U24589 (N_24589,N_16556,N_17728);
xnor U24590 (N_24590,N_14142,N_16838);
and U24591 (N_24591,N_13882,N_18692);
nand U24592 (N_24592,N_17122,N_16786);
or U24593 (N_24593,N_14315,N_17587);
nand U24594 (N_24594,N_18082,N_16535);
xnor U24595 (N_24595,N_15791,N_17305);
nand U24596 (N_24596,N_17078,N_13522);
and U24597 (N_24597,N_17697,N_15233);
nand U24598 (N_24598,N_15641,N_16960);
nand U24599 (N_24599,N_13038,N_14856);
or U24600 (N_24600,N_12706,N_16792);
xnor U24601 (N_24601,N_16892,N_14006);
and U24602 (N_24602,N_13718,N_18714);
and U24603 (N_24603,N_18625,N_18287);
or U24604 (N_24604,N_12598,N_18005);
xnor U24605 (N_24605,N_13774,N_17376);
xor U24606 (N_24606,N_16372,N_17547);
xnor U24607 (N_24607,N_13899,N_16776);
nor U24608 (N_24608,N_16508,N_14863);
nand U24609 (N_24609,N_16620,N_17055);
xor U24610 (N_24610,N_14778,N_17988);
xor U24611 (N_24611,N_14054,N_17051);
nand U24612 (N_24612,N_16305,N_17676);
xnor U24613 (N_24613,N_16608,N_14740);
and U24614 (N_24614,N_16768,N_15098);
nor U24615 (N_24615,N_15705,N_16441);
xnor U24616 (N_24616,N_14614,N_16600);
and U24617 (N_24617,N_17404,N_16684);
xor U24618 (N_24618,N_18696,N_13966);
xnor U24619 (N_24619,N_12809,N_12526);
and U24620 (N_24620,N_12650,N_18500);
nand U24621 (N_24621,N_18267,N_17727);
nor U24622 (N_24622,N_17962,N_18433);
nor U24623 (N_24623,N_15010,N_16603);
or U24624 (N_24624,N_15601,N_13494);
or U24625 (N_24625,N_16230,N_18488);
or U24626 (N_24626,N_13997,N_13085);
and U24627 (N_24627,N_17850,N_14847);
nor U24628 (N_24628,N_14426,N_14116);
nor U24629 (N_24629,N_17784,N_15015);
and U24630 (N_24630,N_14132,N_18022);
nand U24631 (N_24631,N_18184,N_14142);
nand U24632 (N_24632,N_17836,N_17379);
and U24633 (N_24633,N_14344,N_14114);
or U24634 (N_24634,N_14871,N_15604);
nand U24635 (N_24635,N_15225,N_17345);
or U24636 (N_24636,N_12502,N_17893);
or U24637 (N_24637,N_15244,N_17033);
and U24638 (N_24638,N_18607,N_16112);
nor U24639 (N_24639,N_13658,N_12654);
or U24640 (N_24640,N_17344,N_17024);
and U24641 (N_24641,N_13021,N_17455);
or U24642 (N_24642,N_12514,N_18021);
or U24643 (N_24643,N_13730,N_12816);
and U24644 (N_24644,N_13742,N_16094);
or U24645 (N_24645,N_14077,N_17532);
xnor U24646 (N_24646,N_16553,N_16434);
xor U24647 (N_24647,N_14617,N_13747);
nor U24648 (N_24648,N_13451,N_13965);
xor U24649 (N_24649,N_13628,N_14810);
nor U24650 (N_24650,N_15994,N_16072);
nor U24651 (N_24651,N_13533,N_14309);
nor U24652 (N_24652,N_18172,N_17620);
or U24653 (N_24653,N_16556,N_15283);
xor U24654 (N_24654,N_13863,N_15516);
and U24655 (N_24655,N_14991,N_15585);
nor U24656 (N_24656,N_18128,N_16639);
nor U24657 (N_24657,N_13231,N_13573);
nand U24658 (N_24658,N_15024,N_16677);
nand U24659 (N_24659,N_14874,N_14982);
nand U24660 (N_24660,N_13335,N_12811);
and U24661 (N_24661,N_17769,N_18071);
nor U24662 (N_24662,N_16051,N_13224);
and U24663 (N_24663,N_16582,N_18120);
nand U24664 (N_24664,N_16487,N_15526);
or U24665 (N_24665,N_14931,N_14348);
and U24666 (N_24666,N_14052,N_15994);
nand U24667 (N_24667,N_18306,N_13402);
nand U24668 (N_24668,N_15633,N_17302);
or U24669 (N_24669,N_13190,N_16430);
and U24670 (N_24670,N_15435,N_16938);
or U24671 (N_24671,N_14007,N_13599);
and U24672 (N_24672,N_15299,N_18546);
nor U24673 (N_24673,N_15338,N_13391);
nor U24674 (N_24674,N_13371,N_14354);
nand U24675 (N_24675,N_13882,N_13175);
or U24676 (N_24676,N_12874,N_18304);
or U24677 (N_24677,N_15863,N_14087);
nand U24678 (N_24678,N_14921,N_15071);
or U24679 (N_24679,N_18012,N_14696);
or U24680 (N_24680,N_17281,N_17294);
xnor U24681 (N_24681,N_13862,N_15980);
nand U24682 (N_24682,N_13267,N_18018);
xor U24683 (N_24683,N_18078,N_15343);
and U24684 (N_24684,N_17571,N_17226);
xor U24685 (N_24685,N_17233,N_17437);
nor U24686 (N_24686,N_16545,N_13325);
or U24687 (N_24687,N_18663,N_16852);
or U24688 (N_24688,N_14297,N_18277);
or U24689 (N_24689,N_13970,N_15200);
and U24690 (N_24690,N_17009,N_14593);
nor U24691 (N_24691,N_15976,N_18068);
nor U24692 (N_24692,N_18568,N_16431);
nand U24693 (N_24693,N_17365,N_13865);
nor U24694 (N_24694,N_14363,N_12874);
or U24695 (N_24695,N_15185,N_17026);
or U24696 (N_24696,N_16542,N_13035);
nand U24697 (N_24697,N_18737,N_16800);
or U24698 (N_24698,N_16728,N_18597);
nand U24699 (N_24699,N_17892,N_13140);
or U24700 (N_24700,N_12918,N_18678);
or U24701 (N_24701,N_14009,N_14830);
nor U24702 (N_24702,N_13772,N_17467);
and U24703 (N_24703,N_14586,N_12501);
nor U24704 (N_24704,N_13380,N_16730);
or U24705 (N_24705,N_18167,N_17654);
nor U24706 (N_24706,N_17964,N_18685);
nor U24707 (N_24707,N_14437,N_17053);
and U24708 (N_24708,N_17965,N_17340);
and U24709 (N_24709,N_13617,N_14328);
and U24710 (N_24710,N_15098,N_12776);
nand U24711 (N_24711,N_15894,N_17751);
and U24712 (N_24712,N_16297,N_12648);
nand U24713 (N_24713,N_18212,N_15547);
xor U24714 (N_24714,N_13272,N_14127);
nor U24715 (N_24715,N_12833,N_16918);
nor U24716 (N_24716,N_15794,N_16582);
xnor U24717 (N_24717,N_18352,N_13647);
and U24718 (N_24718,N_15157,N_15985);
and U24719 (N_24719,N_17086,N_15125);
or U24720 (N_24720,N_17578,N_16262);
nor U24721 (N_24721,N_14520,N_17826);
and U24722 (N_24722,N_16083,N_14156);
xor U24723 (N_24723,N_18418,N_13212);
nor U24724 (N_24724,N_15163,N_14445);
nor U24725 (N_24725,N_15826,N_12600);
nand U24726 (N_24726,N_12914,N_12663);
nand U24727 (N_24727,N_16386,N_16650);
nor U24728 (N_24728,N_16027,N_13311);
and U24729 (N_24729,N_13818,N_14112);
nand U24730 (N_24730,N_15884,N_16039);
xor U24731 (N_24731,N_14367,N_14480);
or U24732 (N_24732,N_13353,N_17488);
nand U24733 (N_24733,N_12953,N_17098);
nor U24734 (N_24734,N_17828,N_17587);
nor U24735 (N_24735,N_14722,N_18635);
and U24736 (N_24736,N_15668,N_17890);
and U24737 (N_24737,N_17407,N_17806);
nand U24738 (N_24738,N_13214,N_16885);
nand U24739 (N_24739,N_16146,N_13369);
nor U24740 (N_24740,N_15606,N_14230);
or U24741 (N_24741,N_15350,N_18718);
and U24742 (N_24742,N_14187,N_12757);
and U24743 (N_24743,N_17965,N_14767);
xnor U24744 (N_24744,N_15705,N_14913);
xor U24745 (N_24745,N_15490,N_17660);
or U24746 (N_24746,N_16904,N_17080);
and U24747 (N_24747,N_13935,N_14476);
or U24748 (N_24748,N_16317,N_13330);
xor U24749 (N_24749,N_13872,N_16397);
xor U24750 (N_24750,N_17070,N_14223);
nor U24751 (N_24751,N_14037,N_14251);
nand U24752 (N_24752,N_18452,N_15387);
nand U24753 (N_24753,N_15712,N_17471);
nand U24754 (N_24754,N_16232,N_16536);
xor U24755 (N_24755,N_15426,N_14783);
or U24756 (N_24756,N_18723,N_13931);
nand U24757 (N_24757,N_15015,N_15481);
nand U24758 (N_24758,N_15953,N_13150);
xor U24759 (N_24759,N_18472,N_13010);
or U24760 (N_24760,N_15503,N_18034);
or U24761 (N_24761,N_16254,N_17436);
nor U24762 (N_24762,N_13008,N_15136);
or U24763 (N_24763,N_13915,N_16728);
xnor U24764 (N_24764,N_12940,N_18077);
or U24765 (N_24765,N_16332,N_16026);
and U24766 (N_24766,N_15287,N_17257);
nor U24767 (N_24767,N_15720,N_14837);
nand U24768 (N_24768,N_13164,N_16064);
or U24769 (N_24769,N_16713,N_17233);
and U24770 (N_24770,N_13640,N_14452);
nor U24771 (N_24771,N_17221,N_18644);
nand U24772 (N_24772,N_18640,N_16120);
nor U24773 (N_24773,N_18250,N_17957);
nor U24774 (N_24774,N_13498,N_14768);
and U24775 (N_24775,N_15384,N_16597);
nand U24776 (N_24776,N_16047,N_15636);
xnor U24777 (N_24777,N_17963,N_13921);
xnor U24778 (N_24778,N_15078,N_16216);
nand U24779 (N_24779,N_18028,N_14217);
xnor U24780 (N_24780,N_18045,N_16097);
or U24781 (N_24781,N_12549,N_16087);
and U24782 (N_24782,N_15388,N_16956);
xnor U24783 (N_24783,N_16174,N_14523);
xnor U24784 (N_24784,N_13052,N_12665);
or U24785 (N_24785,N_14232,N_13994);
nand U24786 (N_24786,N_12964,N_14099);
and U24787 (N_24787,N_17928,N_14388);
nand U24788 (N_24788,N_16331,N_15464);
nor U24789 (N_24789,N_12917,N_13741);
or U24790 (N_24790,N_14605,N_18003);
xor U24791 (N_24791,N_12945,N_14917);
nor U24792 (N_24792,N_14606,N_15577);
and U24793 (N_24793,N_14306,N_16020);
nor U24794 (N_24794,N_14967,N_12714);
xnor U24795 (N_24795,N_16241,N_13942);
nor U24796 (N_24796,N_17008,N_16061);
nor U24797 (N_24797,N_14823,N_12623);
nand U24798 (N_24798,N_14956,N_15332);
or U24799 (N_24799,N_14559,N_15676);
nor U24800 (N_24800,N_15449,N_18740);
xor U24801 (N_24801,N_16857,N_12659);
or U24802 (N_24802,N_16343,N_12557);
nor U24803 (N_24803,N_14428,N_14404);
xnor U24804 (N_24804,N_16274,N_12764);
and U24805 (N_24805,N_13089,N_17886);
nand U24806 (N_24806,N_16925,N_13910);
nor U24807 (N_24807,N_12786,N_18258);
nor U24808 (N_24808,N_14127,N_13841);
or U24809 (N_24809,N_17158,N_14116);
or U24810 (N_24810,N_16235,N_18154);
and U24811 (N_24811,N_16702,N_17790);
xor U24812 (N_24812,N_17780,N_14737);
or U24813 (N_24813,N_13869,N_15583);
nand U24814 (N_24814,N_18056,N_14256);
xnor U24815 (N_24815,N_16532,N_18204);
xor U24816 (N_24816,N_13298,N_16104);
and U24817 (N_24817,N_16770,N_14979);
nor U24818 (N_24818,N_13072,N_13186);
nor U24819 (N_24819,N_15025,N_16790);
nand U24820 (N_24820,N_14145,N_12976);
and U24821 (N_24821,N_17580,N_13208);
xnor U24822 (N_24822,N_16240,N_13297);
or U24823 (N_24823,N_18696,N_17794);
nor U24824 (N_24824,N_13999,N_14531);
nand U24825 (N_24825,N_15832,N_17051);
nand U24826 (N_24826,N_18745,N_16192);
nand U24827 (N_24827,N_14292,N_14320);
or U24828 (N_24828,N_15269,N_16293);
xnor U24829 (N_24829,N_16464,N_16349);
nand U24830 (N_24830,N_15677,N_16942);
nand U24831 (N_24831,N_16527,N_18038);
nor U24832 (N_24832,N_14086,N_15420);
nor U24833 (N_24833,N_13682,N_17127);
nor U24834 (N_24834,N_13987,N_17211);
nor U24835 (N_24835,N_15074,N_16668);
xor U24836 (N_24836,N_12855,N_12873);
xor U24837 (N_24837,N_16684,N_17944);
and U24838 (N_24838,N_18210,N_15523);
nor U24839 (N_24839,N_18021,N_12639);
and U24840 (N_24840,N_18209,N_15143);
xor U24841 (N_24841,N_15777,N_17541);
nor U24842 (N_24842,N_12943,N_18494);
xnor U24843 (N_24843,N_14149,N_18168);
nor U24844 (N_24844,N_15158,N_13985);
nor U24845 (N_24845,N_17365,N_17808);
nor U24846 (N_24846,N_14672,N_18610);
nand U24847 (N_24847,N_12615,N_16643);
and U24848 (N_24848,N_18205,N_17397);
and U24849 (N_24849,N_17366,N_16058);
nor U24850 (N_24850,N_18327,N_15332);
nor U24851 (N_24851,N_16120,N_17101);
nor U24852 (N_24852,N_17383,N_13932);
xnor U24853 (N_24853,N_17058,N_16003);
xor U24854 (N_24854,N_15099,N_13002);
and U24855 (N_24855,N_16359,N_17663);
and U24856 (N_24856,N_17313,N_18377);
xor U24857 (N_24857,N_13881,N_13878);
xor U24858 (N_24858,N_14113,N_14784);
or U24859 (N_24859,N_12963,N_16675);
nor U24860 (N_24860,N_16195,N_17844);
and U24861 (N_24861,N_14072,N_13329);
and U24862 (N_24862,N_14574,N_16608);
nor U24863 (N_24863,N_18183,N_13606);
nand U24864 (N_24864,N_14823,N_16619);
nand U24865 (N_24865,N_15417,N_16744);
and U24866 (N_24866,N_17268,N_18614);
nor U24867 (N_24867,N_16683,N_16075);
nand U24868 (N_24868,N_18183,N_18728);
or U24869 (N_24869,N_14064,N_13233);
nor U24870 (N_24870,N_13647,N_16193);
nand U24871 (N_24871,N_16808,N_15522);
or U24872 (N_24872,N_17728,N_18123);
nand U24873 (N_24873,N_18692,N_16680);
xor U24874 (N_24874,N_15342,N_17359);
xor U24875 (N_24875,N_14825,N_17036);
or U24876 (N_24876,N_15788,N_16955);
or U24877 (N_24877,N_15645,N_14959);
nand U24878 (N_24878,N_13387,N_17732);
or U24879 (N_24879,N_17357,N_14086);
nand U24880 (N_24880,N_15320,N_16832);
xor U24881 (N_24881,N_17368,N_18044);
nand U24882 (N_24882,N_16130,N_13621);
or U24883 (N_24883,N_12802,N_18249);
xnor U24884 (N_24884,N_18354,N_16876);
xor U24885 (N_24885,N_14556,N_18207);
and U24886 (N_24886,N_17269,N_15657);
or U24887 (N_24887,N_17328,N_13796);
nor U24888 (N_24888,N_13665,N_17604);
or U24889 (N_24889,N_13974,N_14292);
and U24890 (N_24890,N_17625,N_17352);
nor U24891 (N_24891,N_15807,N_15908);
or U24892 (N_24892,N_16331,N_13389);
nor U24893 (N_24893,N_18387,N_17584);
nor U24894 (N_24894,N_13364,N_15893);
nor U24895 (N_24895,N_18291,N_16322);
xnor U24896 (N_24896,N_17663,N_17925);
and U24897 (N_24897,N_14104,N_16931);
nand U24898 (N_24898,N_17094,N_18646);
and U24899 (N_24899,N_14455,N_14810);
xor U24900 (N_24900,N_16385,N_17283);
and U24901 (N_24901,N_17661,N_17410);
nand U24902 (N_24902,N_14966,N_15883);
nor U24903 (N_24903,N_17806,N_15537);
nand U24904 (N_24904,N_13932,N_18334);
and U24905 (N_24905,N_16015,N_15306);
and U24906 (N_24906,N_16259,N_18452);
or U24907 (N_24907,N_16700,N_15704);
and U24908 (N_24908,N_14624,N_14753);
and U24909 (N_24909,N_13907,N_16550);
nor U24910 (N_24910,N_15683,N_13886);
and U24911 (N_24911,N_14186,N_17862);
or U24912 (N_24912,N_16154,N_17204);
or U24913 (N_24913,N_17168,N_14460);
nand U24914 (N_24914,N_16291,N_15284);
nor U24915 (N_24915,N_17915,N_14470);
or U24916 (N_24916,N_16656,N_13144);
xnor U24917 (N_24917,N_13469,N_17092);
or U24918 (N_24918,N_13311,N_15711);
and U24919 (N_24919,N_14525,N_16653);
and U24920 (N_24920,N_18746,N_16573);
nand U24921 (N_24921,N_12992,N_17494);
or U24922 (N_24922,N_18695,N_15771);
or U24923 (N_24923,N_15455,N_13967);
xor U24924 (N_24924,N_13867,N_17167);
nand U24925 (N_24925,N_16415,N_13244);
and U24926 (N_24926,N_17797,N_15024);
nor U24927 (N_24927,N_12586,N_17147);
and U24928 (N_24928,N_14751,N_14312);
nand U24929 (N_24929,N_16965,N_12768);
nand U24930 (N_24930,N_13469,N_14657);
and U24931 (N_24931,N_17945,N_12921);
nor U24932 (N_24932,N_14497,N_13692);
nor U24933 (N_24933,N_15018,N_16156);
or U24934 (N_24934,N_14611,N_14182);
and U24935 (N_24935,N_15348,N_12910);
and U24936 (N_24936,N_13039,N_18490);
or U24937 (N_24937,N_16961,N_14721);
nand U24938 (N_24938,N_13117,N_14571);
nand U24939 (N_24939,N_17030,N_17325);
and U24940 (N_24940,N_18564,N_15410);
and U24941 (N_24941,N_13209,N_13158);
or U24942 (N_24942,N_18650,N_16669);
and U24943 (N_24943,N_14343,N_14871);
nand U24944 (N_24944,N_17933,N_18557);
nand U24945 (N_24945,N_18267,N_12568);
and U24946 (N_24946,N_14198,N_15969);
nor U24947 (N_24947,N_15543,N_13035);
and U24948 (N_24948,N_17356,N_16050);
and U24949 (N_24949,N_18657,N_13657);
or U24950 (N_24950,N_12686,N_13024);
and U24951 (N_24951,N_16267,N_16284);
or U24952 (N_24952,N_13184,N_15724);
nand U24953 (N_24953,N_17133,N_15945);
nand U24954 (N_24954,N_17270,N_13633);
and U24955 (N_24955,N_13357,N_16703);
nor U24956 (N_24956,N_12576,N_17127);
and U24957 (N_24957,N_15174,N_15554);
nand U24958 (N_24958,N_16739,N_17436);
nand U24959 (N_24959,N_14741,N_18049);
xnor U24960 (N_24960,N_16083,N_14619);
or U24961 (N_24961,N_16157,N_13519);
nor U24962 (N_24962,N_13992,N_16525);
and U24963 (N_24963,N_17285,N_18084);
nand U24964 (N_24964,N_14001,N_13960);
nor U24965 (N_24965,N_14556,N_18467);
and U24966 (N_24966,N_17188,N_16833);
nor U24967 (N_24967,N_18033,N_13193);
and U24968 (N_24968,N_17141,N_17587);
nand U24969 (N_24969,N_13992,N_18287);
and U24970 (N_24970,N_16347,N_15254);
or U24971 (N_24971,N_14114,N_16249);
or U24972 (N_24972,N_14382,N_16346);
nor U24973 (N_24973,N_12837,N_18298);
nor U24974 (N_24974,N_16027,N_18095);
nand U24975 (N_24975,N_18190,N_14436);
nor U24976 (N_24976,N_13782,N_14899);
nor U24977 (N_24977,N_16882,N_17650);
xnor U24978 (N_24978,N_13966,N_17307);
xnor U24979 (N_24979,N_16552,N_13788);
nor U24980 (N_24980,N_16911,N_14169);
xor U24981 (N_24981,N_16833,N_16628);
nand U24982 (N_24982,N_13539,N_15394);
and U24983 (N_24983,N_18436,N_15983);
nand U24984 (N_24984,N_16845,N_14963);
or U24985 (N_24985,N_13103,N_12913);
or U24986 (N_24986,N_14005,N_15056);
nand U24987 (N_24987,N_18205,N_13780);
or U24988 (N_24988,N_13378,N_14184);
or U24989 (N_24989,N_15637,N_17807);
nand U24990 (N_24990,N_17420,N_14243);
or U24991 (N_24991,N_18471,N_14362);
nand U24992 (N_24992,N_15791,N_13055);
or U24993 (N_24993,N_13541,N_15947);
or U24994 (N_24994,N_13696,N_15897);
xor U24995 (N_24995,N_17609,N_14703);
nand U24996 (N_24996,N_14742,N_16665);
or U24997 (N_24997,N_14242,N_17842);
xnor U24998 (N_24998,N_17645,N_14364);
nand U24999 (N_24999,N_17095,N_14150);
and UO_0 (O_0,N_19476,N_20603);
nand UO_1 (O_1,N_22433,N_21286);
xnor UO_2 (O_2,N_24606,N_23250);
nand UO_3 (O_3,N_23410,N_22284);
nand UO_4 (O_4,N_24584,N_23003);
or UO_5 (O_5,N_22193,N_24973);
nor UO_6 (O_6,N_19137,N_21641);
nor UO_7 (O_7,N_22832,N_20228);
nand UO_8 (O_8,N_18995,N_22196);
and UO_9 (O_9,N_21432,N_21183);
or UO_10 (O_10,N_20252,N_21667);
or UO_11 (O_11,N_21004,N_21738);
and UO_12 (O_12,N_22904,N_24580);
and UO_13 (O_13,N_24978,N_21799);
and UO_14 (O_14,N_24175,N_23112);
nand UO_15 (O_15,N_24850,N_22113);
and UO_16 (O_16,N_20501,N_20073);
and UO_17 (O_17,N_19768,N_21867);
nand UO_18 (O_18,N_21508,N_20506);
or UO_19 (O_19,N_24768,N_20816);
nand UO_20 (O_20,N_19592,N_23154);
nand UO_21 (O_21,N_19717,N_24953);
and UO_22 (O_22,N_23006,N_24569);
nand UO_23 (O_23,N_19651,N_20849);
nand UO_24 (O_24,N_19020,N_19293);
nor UO_25 (O_25,N_19231,N_19048);
nand UO_26 (O_26,N_22243,N_20237);
nor UO_27 (O_27,N_21801,N_22941);
and UO_28 (O_28,N_24017,N_20780);
nor UO_29 (O_29,N_23636,N_20767);
nand UO_30 (O_30,N_19492,N_21790);
and UO_31 (O_31,N_21614,N_21953);
and UO_32 (O_32,N_21418,N_24706);
nor UO_33 (O_33,N_23982,N_24397);
nor UO_34 (O_34,N_24105,N_19914);
and UO_35 (O_35,N_20362,N_20659);
nor UO_36 (O_36,N_23035,N_19736);
nor UO_37 (O_37,N_21864,N_23625);
and UO_38 (O_38,N_20021,N_19983);
nor UO_39 (O_39,N_20456,N_21431);
or UO_40 (O_40,N_23283,N_19694);
and UO_41 (O_41,N_20467,N_24027);
nand UO_42 (O_42,N_24415,N_19656);
nor UO_43 (O_43,N_23858,N_19999);
and UO_44 (O_44,N_24049,N_22963);
and UO_45 (O_45,N_20848,N_23307);
nand UO_46 (O_46,N_20739,N_24000);
or UO_47 (O_47,N_22856,N_20498);
nand UO_48 (O_48,N_21853,N_18907);
or UO_49 (O_49,N_21701,N_22507);
nor UO_50 (O_50,N_21501,N_22150);
xnor UO_51 (O_51,N_18785,N_24742);
nand UO_52 (O_52,N_24680,N_24724);
nand UO_53 (O_53,N_24373,N_24298);
or UO_54 (O_54,N_21369,N_21902);
or UO_55 (O_55,N_21816,N_21274);
or UO_56 (O_56,N_20920,N_18841);
nor UO_57 (O_57,N_19980,N_24575);
xor UO_58 (O_58,N_20496,N_22700);
nor UO_59 (O_59,N_19838,N_21765);
nand UO_60 (O_60,N_21281,N_22945);
and UO_61 (O_61,N_21015,N_22631);
xnor UO_62 (O_62,N_22979,N_21311);
or UO_63 (O_63,N_20083,N_24735);
nand UO_64 (O_64,N_22007,N_20040);
or UO_65 (O_65,N_22137,N_24755);
and UO_66 (O_66,N_20323,N_19728);
and UO_67 (O_67,N_20941,N_19082);
and UO_68 (O_68,N_23058,N_19818);
or UO_69 (O_69,N_21118,N_18777);
xor UO_70 (O_70,N_24754,N_19077);
xnor UO_71 (O_71,N_21607,N_21065);
or UO_72 (O_72,N_20262,N_24380);
nor UO_73 (O_73,N_21206,N_19128);
nor UO_74 (O_74,N_19991,N_23381);
or UO_75 (O_75,N_18831,N_24544);
nand UO_76 (O_76,N_19166,N_23439);
nor UO_77 (O_77,N_20829,N_24582);
xnor UO_78 (O_78,N_22417,N_20776);
nor UO_79 (O_79,N_18924,N_24124);
nand UO_80 (O_80,N_22850,N_20759);
and UO_81 (O_81,N_20598,N_23957);
nand UO_82 (O_82,N_22056,N_23737);
nor UO_83 (O_83,N_19262,N_21037);
nand UO_84 (O_84,N_22048,N_21958);
nand UO_85 (O_85,N_23918,N_20960);
or UO_86 (O_86,N_20278,N_23649);
nand UO_87 (O_87,N_18860,N_21456);
nand UO_88 (O_88,N_19148,N_22237);
nand UO_89 (O_89,N_18973,N_19690);
nand UO_90 (O_90,N_23643,N_22896);
xnor UO_91 (O_91,N_21944,N_19979);
nor UO_92 (O_92,N_20214,N_24103);
and UO_93 (O_93,N_24834,N_19844);
and UO_94 (O_94,N_22613,N_19143);
or UO_95 (O_95,N_21376,N_24288);
nand UO_96 (O_96,N_20076,N_21811);
xnor UO_97 (O_97,N_18882,N_24360);
and UO_98 (O_98,N_24263,N_19475);
and UO_99 (O_99,N_19035,N_23683);
and UO_100 (O_100,N_24371,N_20585);
or UO_101 (O_101,N_22512,N_21074);
xnor UO_102 (O_102,N_23747,N_22790);
xnor UO_103 (O_103,N_20288,N_23458);
or UO_104 (O_104,N_22277,N_22639);
or UO_105 (O_105,N_21740,N_20538);
nand UO_106 (O_106,N_23533,N_19207);
nor UO_107 (O_107,N_24980,N_22972);
or UO_108 (O_108,N_18898,N_19296);
or UO_109 (O_109,N_18974,N_19874);
or UO_110 (O_110,N_21457,N_18796);
and UO_111 (O_111,N_19100,N_23952);
nand UO_112 (O_112,N_21787,N_24656);
and UO_113 (O_113,N_20365,N_19558);
nand UO_114 (O_114,N_23243,N_22106);
nand UO_115 (O_115,N_22651,N_24223);
and UO_116 (O_116,N_20921,N_20660);
or UO_117 (O_117,N_23367,N_21886);
or UO_118 (O_118,N_22879,N_19674);
nand UO_119 (O_119,N_20572,N_24699);
xnor UO_120 (O_120,N_23732,N_21935);
or UO_121 (O_121,N_21513,N_22042);
nand UO_122 (O_122,N_23323,N_22374);
or UO_123 (O_123,N_20063,N_19418);
nand UO_124 (O_124,N_22161,N_20976);
or UO_125 (O_125,N_24076,N_24142);
nor UO_126 (O_126,N_21692,N_21574);
and UO_127 (O_127,N_24244,N_23133);
and UO_128 (O_128,N_20211,N_23720);
or UO_129 (O_129,N_21039,N_23885);
nor UO_130 (O_130,N_24395,N_24410);
xor UO_131 (O_131,N_22623,N_22802);
or UO_132 (O_132,N_22021,N_21377);
xor UO_133 (O_133,N_19198,N_24739);
nand UO_134 (O_134,N_23221,N_23734);
or UO_135 (O_135,N_22707,N_23779);
xor UO_136 (O_136,N_21444,N_21287);
and UO_137 (O_137,N_18789,N_19356);
xor UO_138 (O_138,N_20452,N_24287);
xnor UO_139 (O_139,N_24711,N_23024);
xnor UO_140 (O_140,N_24871,N_19856);
and UO_141 (O_141,N_19222,N_24198);
nor UO_142 (O_142,N_21411,N_22934);
xnor UO_143 (O_143,N_24452,N_21256);
or UO_144 (O_144,N_23363,N_21949);
nand UO_145 (O_145,N_22951,N_20200);
or UO_146 (O_146,N_19494,N_21794);
or UO_147 (O_147,N_24473,N_22662);
or UO_148 (O_148,N_20640,N_21477);
xnor UO_149 (O_149,N_22486,N_21537);
nor UO_150 (O_150,N_20355,N_22404);
xnor UO_151 (O_151,N_23531,N_22083);
or UO_152 (O_152,N_19902,N_22275);
nand UO_153 (O_153,N_22684,N_19240);
and UO_154 (O_154,N_18851,N_20050);
nand UO_155 (O_155,N_20238,N_20706);
nand UO_156 (O_156,N_19320,N_23043);
and UO_157 (O_157,N_21270,N_20689);
nor UO_158 (O_158,N_23429,N_21919);
nor UO_159 (O_159,N_24228,N_21463);
and UO_160 (O_160,N_23695,N_22897);
or UO_161 (O_161,N_23705,N_23856);
nor UO_162 (O_162,N_20004,N_23749);
or UO_163 (O_163,N_19400,N_23633);
or UO_164 (O_164,N_20353,N_19517);
and UO_165 (O_165,N_24719,N_23394);
and UO_166 (O_166,N_22840,N_19364);
nand UO_167 (O_167,N_20663,N_24885);
nand UO_168 (O_168,N_19556,N_23128);
xnor UO_169 (O_169,N_23741,N_22779);
and UO_170 (O_170,N_19923,N_18773);
xor UO_171 (O_171,N_22207,N_23699);
or UO_172 (O_172,N_23645,N_24418);
xor UO_173 (O_173,N_24422,N_23159);
nand UO_174 (O_174,N_20242,N_22589);
and UO_175 (O_175,N_20629,N_21649);
or UO_176 (O_176,N_20779,N_21521);
or UO_177 (O_177,N_20518,N_21770);
and UO_178 (O_178,N_21086,N_20898);
nor UO_179 (O_179,N_23377,N_19875);
and UO_180 (O_180,N_20328,N_20126);
xor UO_181 (O_181,N_24894,N_19942);
nand UO_182 (O_182,N_19948,N_20109);
or UO_183 (O_183,N_24374,N_19336);
nor UO_184 (O_184,N_21713,N_19568);
nand UO_185 (O_185,N_20606,N_21581);
nor UO_186 (O_186,N_19343,N_19646);
and UO_187 (O_187,N_24110,N_23914);
xnor UO_188 (O_188,N_22049,N_22645);
nor UO_189 (O_189,N_19686,N_23913);
and UO_190 (O_190,N_21893,N_23748);
and UO_191 (O_191,N_23021,N_21878);
xnor UO_192 (O_192,N_21851,N_22480);
and UO_193 (O_193,N_23138,N_21977);
or UO_194 (O_194,N_23151,N_21450);
xor UO_195 (O_195,N_19798,N_23566);
nand UO_196 (O_196,N_23286,N_23099);
and UO_197 (O_197,N_19287,N_23718);
xor UO_198 (O_198,N_24698,N_23074);
xnor UO_199 (O_199,N_21361,N_24929);
xor UO_200 (O_200,N_22523,N_21900);
nor UO_201 (O_201,N_21197,N_24831);
xor UO_202 (O_202,N_23976,N_23130);
xor UO_203 (O_203,N_21626,N_22233);
nor UO_204 (O_204,N_24348,N_19537);
xor UO_205 (O_205,N_19088,N_18966);
nand UO_206 (O_206,N_20623,N_24256);
xor UO_207 (O_207,N_20907,N_20914);
nand UO_208 (O_208,N_21401,N_20236);
nand UO_209 (O_209,N_21446,N_19775);
nand UO_210 (O_210,N_20951,N_24773);
nor UO_211 (O_211,N_24559,N_20903);
or UO_212 (O_212,N_23326,N_23218);
and UO_213 (O_213,N_21407,N_19858);
and UO_214 (O_214,N_23481,N_20010);
nand UO_215 (O_215,N_19031,N_19519);
and UO_216 (O_216,N_22408,N_23382);
or UO_217 (O_217,N_19053,N_18854);
and UO_218 (O_218,N_19586,N_24196);
nor UO_219 (O_219,N_18969,N_19976);
nor UO_220 (O_220,N_21233,N_23254);
xor UO_221 (O_221,N_24682,N_20985);
and UO_222 (O_222,N_21166,N_19968);
nand UO_223 (O_223,N_24787,N_22105);
xnor UO_224 (O_224,N_23091,N_20442);
and UO_225 (O_225,N_20166,N_22381);
nand UO_226 (O_226,N_19094,N_19459);
nor UO_227 (O_227,N_23215,N_24435);
and UO_228 (O_228,N_20547,N_23269);
xor UO_229 (O_229,N_22723,N_23068);
nor UO_230 (O_230,N_22013,N_19414);
or UO_231 (O_231,N_22428,N_23543);
xor UO_232 (O_232,N_24121,N_21227);
nor UO_233 (O_233,N_23846,N_24138);
or UO_234 (O_234,N_20979,N_20641);
nor UO_235 (O_235,N_24558,N_23251);
nor UO_236 (O_236,N_23805,N_24084);
and UO_237 (O_237,N_24922,N_24383);
xnor UO_238 (O_238,N_22079,N_19486);
or UO_239 (O_239,N_24564,N_24357);
nor UO_240 (O_240,N_20874,N_21198);
nor UO_241 (O_241,N_20709,N_24734);
or UO_242 (O_242,N_21800,N_21204);
nor UO_243 (O_243,N_22311,N_24858);
xor UO_244 (O_244,N_24339,N_24997);
or UO_245 (O_245,N_20583,N_21621);
nand UO_246 (O_246,N_21035,N_20644);
and UO_247 (O_247,N_21689,N_21364);
nor UO_248 (O_248,N_22906,N_19830);
xor UO_249 (O_249,N_19572,N_23238);
nand UO_250 (O_250,N_19273,N_19557);
or UO_251 (O_251,N_19878,N_19772);
xor UO_252 (O_252,N_22654,N_22778);
nor UO_253 (O_253,N_19750,N_22045);
or UO_254 (O_254,N_24286,N_24468);
nor UO_255 (O_255,N_22306,N_22289);
nand UO_256 (O_256,N_19480,N_23796);
xor UO_257 (O_257,N_21484,N_19407);
or UO_258 (O_258,N_22175,N_24501);
and UO_259 (O_259,N_24224,N_19609);
nor UO_260 (O_260,N_20826,N_23514);
xor UO_261 (O_261,N_19988,N_22482);
or UO_262 (O_262,N_18862,N_20906);
nand UO_263 (O_263,N_21041,N_21474);
xnor UO_264 (O_264,N_21234,N_22808);
or UO_265 (O_265,N_20910,N_24630);
nor UO_266 (O_266,N_24006,N_21303);
nor UO_267 (O_267,N_24405,N_24292);
or UO_268 (O_268,N_23657,N_22057);
nand UO_269 (O_269,N_19934,N_21638);
or UO_270 (O_270,N_24060,N_24269);
and UO_271 (O_271,N_20795,N_24639);
xnor UO_272 (O_272,N_19006,N_23665);
or UO_273 (O_273,N_19041,N_21615);
or UO_274 (O_274,N_20661,N_22354);
or UO_275 (O_275,N_24800,N_24191);
and UO_276 (O_276,N_21176,N_18858);
nor UO_277 (O_277,N_18988,N_20299);
nand UO_278 (O_278,N_20343,N_22873);
and UO_279 (O_279,N_22719,N_23430);
nor UO_280 (O_280,N_24647,N_19249);
nor UO_281 (O_281,N_23380,N_18847);
xnor UO_282 (O_282,N_22813,N_19477);
xor UO_283 (O_283,N_22564,N_21647);
nand UO_284 (O_284,N_19420,N_21622);
nand UO_285 (O_285,N_24577,N_22276);
and UO_286 (O_286,N_20577,N_23950);
or UO_287 (O_287,N_21138,N_21100);
nand UO_288 (O_288,N_24497,N_19941);
or UO_289 (O_289,N_20463,N_23886);
nor UO_290 (O_290,N_18934,N_23685);
and UO_291 (O_291,N_19561,N_24109);
or UO_292 (O_292,N_19472,N_24107);
nand UO_293 (O_293,N_19510,N_20449);
xnor UO_294 (O_294,N_23833,N_19160);
and UO_295 (O_295,N_21729,N_19051);
or UO_296 (O_296,N_19354,N_20808);
xnor UO_297 (O_297,N_22741,N_21993);
xnor UO_298 (O_298,N_22722,N_20727);
or UO_299 (O_299,N_19629,N_22219);
xnor UO_300 (O_300,N_24725,N_20206);
or UO_301 (O_301,N_21651,N_20479);
or UO_302 (O_302,N_23217,N_21006);
nor UO_303 (O_303,N_24021,N_23968);
nor UO_304 (O_304,N_23418,N_24805);
xor UO_305 (O_305,N_21273,N_22477);
nand UO_306 (O_306,N_19398,N_19920);
nor UO_307 (O_307,N_20049,N_22823);
or UO_308 (O_308,N_22641,N_22916);
nor UO_309 (O_309,N_20873,N_21742);
and UO_310 (O_310,N_19797,N_23707);
nor UO_311 (O_311,N_21684,N_20665);
nand UO_312 (O_312,N_20305,N_18819);
xnor UO_313 (O_313,N_22035,N_21490);
or UO_314 (O_314,N_23146,N_19023);
nor UO_315 (O_315,N_19086,N_23455);
xnor UO_316 (O_316,N_23437,N_19089);
xnor UO_317 (O_317,N_21072,N_22212);
or UO_318 (O_318,N_20711,N_21170);
nand UO_319 (O_319,N_23010,N_23270);
xnor UO_320 (O_320,N_22368,N_22747);
and UO_321 (O_321,N_24576,N_23922);
and UO_322 (O_322,N_23216,N_19816);
nand UO_323 (O_323,N_21955,N_21105);
nand UO_324 (O_324,N_21603,N_21119);
nor UO_325 (O_325,N_19248,N_23352);
or UO_326 (O_326,N_24972,N_19227);
xnor UO_327 (O_327,N_20033,N_24516);
nor UO_328 (O_328,N_21524,N_19072);
and UO_329 (O_329,N_23386,N_21384);
xnor UO_330 (O_330,N_18903,N_22253);
nor UO_331 (O_331,N_20740,N_24909);
xor UO_332 (O_332,N_24048,N_22385);
xnor UO_333 (O_333,N_22740,N_22658);
nor UO_334 (O_334,N_21033,N_21016);
and UO_335 (O_335,N_23702,N_22209);
xor UO_336 (O_336,N_21871,N_19066);
and UO_337 (O_337,N_23731,N_24458);
and UO_338 (O_338,N_21036,N_18997);
and UO_339 (O_339,N_19260,N_23174);
nand UO_340 (O_340,N_19058,N_24425);
or UO_341 (O_341,N_23529,N_23780);
nand UO_342 (O_342,N_22165,N_18991);
xnor UO_343 (O_343,N_21317,N_21720);
or UO_344 (O_344,N_19478,N_20578);
and UO_345 (O_345,N_21698,N_23763);
nand UO_346 (O_346,N_21116,N_24090);
or UO_347 (O_347,N_20959,N_20485);
or UO_348 (O_348,N_19842,N_22214);
and UO_349 (O_349,N_20142,N_19623);
nand UO_350 (O_350,N_23654,N_20386);
and UO_351 (O_351,N_23750,N_19577);
nand UO_352 (O_352,N_21366,N_24556);
or UO_353 (O_353,N_22070,N_24152);
and UO_354 (O_354,N_19621,N_19784);
nor UO_355 (O_355,N_22052,N_20643);
nand UO_356 (O_356,N_23434,N_21946);
xor UO_357 (O_357,N_23231,N_24163);
nor UO_358 (O_358,N_22016,N_22821);
nand UO_359 (O_359,N_19799,N_19722);
nand UO_360 (O_360,N_23427,N_21012);
nor UO_361 (O_361,N_20195,N_19812);
xnor UO_362 (O_362,N_19678,N_20617);
nand UO_363 (O_363,N_21329,N_23304);
xnor UO_364 (O_364,N_21080,N_19275);
or UO_365 (O_365,N_20805,N_24471);
or UO_366 (O_366,N_20302,N_22975);
nor UO_367 (O_367,N_20034,N_20190);
or UO_368 (O_368,N_22678,N_18993);
or UO_369 (O_369,N_23414,N_20441);
nor UO_370 (O_370,N_23915,N_19453);
nand UO_371 (O_371,N_23884,N_24283);
nor UO_372 (O_372,N_24161,N_21824);
or UO_373 (O_373,N_24687,N_21964);
or UO_374 (O_374,N_20859,N_23896);
and UO_375 (O_375,N_20523,N_20513);
nor UO_376 (O_376,N_22012,N_23296);
xnor UO_377 (O_377,N_23357,N_20886);
nor UO_378 (O_378,N_19068,N_23605);
nor UO_379 (O_379,N_21391,N_24986);
nor UO_380 (O_380,N_21127,N_24939);
xnor UO_381 (O_381,N_22483,N_20847);
or UO_382 (O_382,N_20146,N_22504);
nor UO_383 (O_383,N_23416,N_22915);
or UO_384 (O_384,N_20042,N_22818);
nor UO_385 (O_385,N_22458,N_23632);
nor UO_386 (O_386,N_24085,N_22123);
nor UO_387 (O_387,N_22340,N_20789);
and UO_388 (O_388,N_20838,N_24883);
and UO_389 (O_389,N_19987,N_22810);
nand UO_390 (O_390,N_20308,N_23348);
xnor UO_391 (O_391,N_24015,N_19712);
nor UO_392 (O_392,N_23530,N_21817);
nor UO_393 (O_393,N_23839,N_24485);
xor UO_394 (O_394,N_22498,N_21454);
nor UO_395 (O_395,N_20932,N_24213);
nand UO_396 (O_396,N_22545,N_19887);
xnor UO_397 (O_397,N_23358,N_20948);
nand UO_398 (O_398,N_23421,N_23892);
or UO_399 (O_399,N_19584,N_24819);
nand UO_400 (O_400,N_18765,N_20212);
nand UO_401 (O_401,N_22539,N_20690);
xnor UO_402 (O_402,N_22101,N_23509);
nand UO_403 (O_403,N_19447,N_19916);
nor UO_404 (O_404,N_24779,N_24284);
and UO_405 (O_405,N_20990,N_20209);
and UO_406 (O_406,N_22612,N_21929);
xnor UO_407 (O_407,N_19854,N_24583);
nand UO_408 (O_408,N_21514,N_21048);
xor UO_409 (O_409,N_24472,N_20973);
or UO_410 (O_410,N_21066,N_21843);
and UO_411 (O_411,N_21756,N_20336);
or UO_412 (O_412,N_22258,N_20310);
nand UO_413 (O_413,N_23178,N_20373);
nand UO_414 (O_414,N_22771,N_23958);
or UO_415 (O_415,N_21439,N_20356);
xnor UO_416 (O_416,N_24036,N_20187);
nor UO_417 (O_417,N_21712,N_21814);
and UO_418 (O_418,N_21153,N_22592);
and UO_419 (O_419,N_23369,N_20000);
nor UO_420 (O_420,N_23308,N_20558);
xnor UO_421 (O_421,N_22770,N_19698);
nor UO_422 (O_422,N_24310,N_24300);
and UO_423 (O_423,N_24892,N_18880);
and UO_424 (O_424,N_21754,N_21310);
or UO_425 (O_425,N_20773,N_21763);
nor UO_426 (O_426,N_21840,N_22097);
and UO_427 (O_427,N_24114,N_19993);
nor UO_428 (O_428,N_24753,N_22093);
or UO_429 (O_429,N_24747,N_24836);
xor UO_430 (O_430,N_22877,N_20991);
nor UO_431 (O_431,N_21970,N_22050);
xor UO_432 (O_432,N_19140,N_23453);
and UO_433 (O_433,N_24775,N_23592);
xor UO_434 (O_434,N_18939,N_23587);
nand UO_435 (O_435,N_19938,N_24227);
xnor UO_436 (O_436,N_22824,N_23753);
and UO_437 (O_437,N_19202,N_21648);
xnor UO_438 (O_438,N_21263,N_21355);
or UO_439 (O_439,N_24302,N_23825);
nand UO_440 (O_440,N_24597,N_19669);
nand UO_441 (O_441,N_21275,N_24345);
xnor UO_442 (O_442,N_22577,N_24180);
and UO_443 (O_443,N_22980,N_19831);
xnor UO_444 (O_444,N_20604,N_19042);
or UO_445 (O_445,N_19789,N_21239);
nand UO_446 (O_446,N_22073,N_20550);
and UO_447 (O_447,N_23199,N_23635);
nor UO_448 (O_448,N_22878,N_24062);
xnor UO_449 (O_449,N_24572,N_22343);
xnor UO_450 (O_450,N_23200,N_24545);
xor UO_451 (O_451,N_21768,N_18908);
xor UO_452 (O_452,N_24679,N_19982);
and UO_453 (O_453,N_22336,N_22495);
or UO_454 (O_454,N_24306,N_23696);
nand UO_455 (O_455,N_24989,N_22845);
and UO_456 (O_456,N_21566,N_21264);
or UO_457 (O_457,N_21038,N_20793);
or UO_458 (O_458,N_23502,N_23474);
nor UO_459 (O_459,N_21818,N_18822);
nor UO_460 (O_460,N_24511,N_21018);
nor UO_461 (O_461,N_20009,N_21736);
and UO_462 (O_462,N_20056,N_22520);
nand UO_463 (O_463,N_21382,N_24063);
nor UO_464 (O_464,N_24955,N_23090);
and UO_465 (O_465,N_21157,N_22299);
nor UO_466 (O_466,N_19157,N_19467);
nand UO_467 (O_467,N_24586,N_21297);
xor UO_468 (O_468,N_21640,N_23208);
xnor UO_469 (O_469,N_22830,N_23594);
or UO_470 (O_470,N_20435,N_22034);
nand UO_471 (O_471,N_21344,N_24377);
or UO_472 (O_472,N_21905,N_22127);
or UO_473 (O_473,N_21847,N_19161);
or UO_474 (O_474,N_20279,N_24562);
or UO_475 (O_475,N_24305,N_21858);
nor UO_476 (O_476,N_23375,N_23114);
nor UO_477 (O_477,N_20173,N_23582);
or UO_478 (O_478,N_22862,N_21936);
or UO_479 (O_479,N_24866,N_22349);
nand UO_480 (O_480,N_20224,N_20207);
nand UO_481 (O_481,N_22999,N_22278);
or UO_482 (O_482,N_23309,N_23565);
nor UO_483 (O_483,N_24795,N_20667);
nor UO_484 (O_484,N_19965,N_19841);
nor UO_485 (O_485,N_21509,N_21831);
nor UO_486 (O_486,N_19975,N_22466);
or UO_487 (O_487,N_22438,N_23120);
or UO_488 (O_488,N_20183,N_22393);
or UO_489 (O_489,N_20400,N_23807);
or UO_490 (O_490,N_20700,N_20069);
or UO_491 (O_491,N_24813,N_23642);
nand UO_492 (O_492,N_22230,N_24113);
nand UO_493 (O_493,N_23033,N_20445);
nand UO_494 (O_494,N_20717,N_23712);
and UO_495 (O_495,N_18982,N_20845);
and UO_496 (O_496,N_21282,N_22600);
nand UO_497 (O_497,N_24384,N_24675);
or UO_498 (O_498,N_22331,N_22389);
xor UO_499 (O_499,N_19259,N_22554);
nand UO_500 (O_500,N_24399,N_22659);
or UO_501 (O_501,N_21587,N_21396);
or UO_502 (O_502,N_19479,N_20102);
nand UO_503 (O_503,N_20961,N_24760);
and UO_504 (O_504,N_22925,N_20648);
and UO_505 (O_505,N_21142,N_21702);
xnor UO_506 (O_506,N_20148,N_23588);
xnor UO_507 (O_507,N_22478,N_24788);
and UO_508 (O_508,N_20251,N_20239);
nor UO_509 (O_509,N_23867,N_21228);
xor UO_510 (O_510,N_19907,N_20204);
and UO_511 (O_511,N_20947,N_20208);
nor UO_512 (O_512,N_22792,N_21942);
or UO_513 (O_513,N_22936,N_23770);
nor UO_514 (O_514,N_21972,N_19636);
nand UO_515 (O_515,N_23752,N_19021);
and UO_516 (O_516,N_23658,N_24259);
and UO_517 (O_517,N_22383,N_22245);
or UO_518 (O_518,N_21512,N_19996);
and UO_519 (O_519,N_21541,N_24316);
xor UO_520 (O_520,N_19576,N_22051);
and UO_521 (O_521,N_21194,N_23225);
or UO_522 (O_522,N_21250,N_20919);
or UO_523 (O_523,N_23697,N_24661);
or UO_524 (O_524,N_21681,N_23371);
xor UO_525 (O_525,N_19951,N_20374);
nand UO_526 (O_526,N_21351,N_22114);
xnor UO_527 (O_527,N_21440,N_20059);
nand UO_528 (O_528,N_22714,N_22942);
nor UO_529 (O_529,N_19375,N_21455);
nor UO_530 (O_530,N_23239,N_20199);
or UO_531 (O_531,N_22536,N_23639);
nand UO_532 (O_532,N_21110,N_20213);
and UO_533 (O_533,N_20217,N_24478);
and UO_534 (O_534,N_19639,N_21745);
nand UO_535 (O_535,N_24212,N_22914);
and UO_536 (O_536,N_22055,N_21055);
and UO_537 (O_537,N_20790,N_19550);
nor UO_538 (O_538,N_23791,N_20320);
and UO_539 (O_539,N_24931,N_22729);
nor UO_540 (O_540,N_20646,N_20702);
nand UO_541 (O_541,N_21123,N_24416);
or UO_542 (O_542,N_19186,N_22305);
nand UO_543 (O_543,N_19239,N_21318);
nand UO_544 (O_544,N_21887,N_24434);
nand UO_545 (O_545,N_19670,N_22390);
nand UO_546 (O_546,N_24177,N_23282);
xnor UO_547 (O_547,N_22735,N_22529);
or UO_548 (O_548,N_20472,N_21832);
and UO_549 (O_549,N_24047,N_23105);
and UO_550 (O_550,N_23379,N_23841);
or UO_551 (O_551,N_23262,N_21926);
nand UO_552 (O_552,N_22198,N_23845);
xor UO_553 (O_553,N_23498,N_22889);
nand UO_554 (O_554,N_20058,N_18837);
and UO_555 (O_555,N_18820,N_20607);
nand UO_556 (O_556,N_23946,N_19582);
or UO_557 (O_557,N_19062,N_20258);
and UO_558 (O_558,N_24925,N_22699);
and UO_559 (O_559,N_21109,N_21673);
and UO_560 (O_560,N_21555,N_22227);
and UO_561 (O_561,N_22399,N_19108);
and UO_562 (O_562,N_19268,N_23370);
nand UO_563 (O_563,N_20488,N_23118);
xnor UO_564 (O_564,N_19960,N_21325);
nand UO_565 (O_565,N_19450,N_19465);
xnor UO_566 (O_566,N_20115,N_21011);
nor UO_567 (O_567,N_24536,N_19085);
or UO_568 (O_568,N_21114,N_22638);
xnor UO_569 (O_569,N_19740,N_23002);
nand UO_570 (O_570,N_21082,N_18770);
or UO_571 (O_571,N_24426,N_24309);
nand UO_572 (O_572,N_20852,N_22852);
nand UO_573 (O_573,N_23803,N_21497);
xnor UO_574 (O_574,N_22382,N_22679);
nor UO_575 (O_575,N_22582,N_22876);
nor UO_576 (O_576,N_24143,N_19595);
xor UO_577 (O_577,N_21106,N_22672);
or UO_578 (O_578,N_20119,N_19536);
or UO_579 (O_579,N_19012,N_18918);
nor UO_580 (O_580,N_19419,N_22344);
or UO_581 (O_581,N_22894,N_24176);
and UO_582 (O_582,N_23129,N_24253);
nand UO_583 (O_583,N_23924,N_20651);
and UO_584 (O_584,N_20107,N_21288);
xor UO_585 (O_585,N_24921,N_23467);
nor UO_586 (O_586,N_22882,N_23951);
xor UO_587 (O_587,N_20269,N_20232);
nor UO_588 (O_588,N_21945,N_23402);
xor UO_589 (O_589,N_23905,N_20731);
nor UO_590 (O_590,N_24367,N_21600);
or UO_591 (O_591,N_21582,N_22670);
xor UO_592 (O_592,N_24341,N_23517);
nand UO_593 (O_593,N_22886,N_21852);
xnor UO_594 (O_594,N_18792,N_24590);
or UO_595 (O_595,N_24835,N_20930);
nand UO_596 (O_596,N_24064,N_20297);
xor UO_597 (O_597,N_20231,N_18876);
nor UO_598 (O_598,N_24072,N_22801);
or UO_599 (O_599,N_19504,N_22259);
and UO_600 (O_600,N_24878,N_23818);
or UO_601 (O_601,N_20439,N_19511);
nor UO_602 (O_602,N_18965,N_24517);
nor UO_603 (O_603,N_19624,N_22216);
nand UO_604 (O_604,N_22831,N_18829);
or UO_605 (O_605,N_20283,N_19913);
nor UO_606 (O_606,N_19119,N_18865);
and UO_607 (O_607,N_21252,N_23488);
xor UO_608 (O_608,N_22162,N_24344);
nor UO_609 (O_609,N_19280,N_18774);
nand UO_610 (O_610,N_22286,N_19985);
xnor UO_611 (O_611,N_24400,N_23134);
and UO_612 (O_612,N_22296,N_20516);
nor UO_613 (O_613,N_20715,N_24585);
xor UO_614 (O_614,N_19508,N_19331);
nand UO_615 (O_615,N_22966,N_22601);
xor UO_616 (O_616,N_23465,N_18897);
nor UO_617 (O_617,N_19645,N_19491);
and UO_618 (O_618,N_24902,N_24442);
or UO_619 (O_619,N_20595,N_24453);
or UO_620 (O_620,N_24127,N_21976);
or UO_621 (O_621,N_20517,N_18845);
or UO_622 (O_622,N_20270,N_21149);
xnor UO_623 (O_623,N_23906,N_22372);
xor UO_624 (O_624,N_24183,N_20575);
and UO_625 (O_625,N_24940,N_23048);
nand UO_626 (O_626,N_20628,N_23290);
or UO_627 (O_627,N_19429,N_24557);
or UO_628 (O_628,N_19081,N_20394);
xnor UO_629 (O_629,N_20605,N_23921);
xor UO_630 (O_630,N_20304,N_24145);
nand UO_631 (O_631,N_24201,N_24466);
nor UO_632 (O_632,N_19738,N_19279);
nor UO_633 (O_633,N_23113,N_20108);
xor UO_634 (O_634,N_20413,N_23015);
xnor UO_635 (O_635,N_23733,N_20163);
xnor UO_636 (O_636,N_22716,N_23062);
or UO_637 (O_637,N_23482,N_20936);
and UO_638 (O_638,N_21480,N_19215);
nor UO_639 (O_639,N_23077,N_22964);
or UO_640 (O_640,N_22283,N_22842);
xor UO_641 (O_641,N_24243,N_24745);
nand UO_642 (O_642,N_19358,N_20543);
or UO_643 (O_643,N_19229,N_23201);
nor UO_644 (O_644,N_24261,N_22224);
nand UO_645 (O_645,N_24718,N_24678);
nand UO_646 (O_646,N_23965,N_23081);
or UO_647 (O_647,N_19329,N_24636);
or UO_648 (O_648,N_21385,N_22782);
and UO_649 (O_649,N_23548,N_24769);
or UO_650 (O_650,N_21573,N_21388);
and UO_651 (O_651,N_20088,N_18817);
nor UO_652 (O_652,N_19243,N_21219);
nor UO_653 (O_653,N_21182,N_22712);
nor UO_654 (O_654,N_20783,N_21894);
nand UO_655 (O_655,N_19446,N_19926);
xnor UO_656 (O_656,N_19885,N_20272);
xnor UO_657 (O_657,N_21722,N_22334);
xor UO_658 (O_658,N_22402,N_23859);
or UO_659 (O_659,N_24948,N_20477);
or UO_660 (O_660,N_20367,N_20784);
or UO_661 (O_661,N_21855,N_19442);
and UO_662 (O_662,N_20937,N_22310);
nand UO_663 (O_663,N_23994,N_23738);
and UO_664 (O_664,N_24165,N_24462);
nor UO_665 (O_665,N_22036,N_24538);
nor UO_666 (O_666,N_23878,N_24221);
nand UO_667 (O_667,N_23891,N_22037);
and UO_668 (O_668,N_19495,N_21184);
nand UO_669 (O_669,N_22351,N_21828);
or UO_670 (O_670,N_22616,N_21044);
and UO_671 (O_671,N_24663,N_22606);
xnor UO_672 (O_672,N_24872,N_20129);
or UO_673 (O_673,N_23802,N_24061);
nor UO_674 (O_674,N_20155,N_23664);
nor UO_675 (O_675,N_20289,N_24907);
nand UO_676 (O_676,N_24886,N_18866);
or UO_677 (O_677,N_20913,N_19218);
nand UO_678 (O_678,N_20635,N_21335);
or UO_679 (O_679,N_19244,N_19748);
or UO_680 (O_680,N_24120,N_23131);
xor UO_681 (O_681,N_19696,N_19648);
or UO_682 (O_682,N_23451,N_21637);
nor UO_683 (O_683,N_23932,N_23678);
or UO_684 (O_684,N_23709,N_22125);
and UO_685 (O_685,N_20478,N_20799);
xnor UO_686 (O_686,N_20306,N_19406);
or UO_687 (O_687,N_23089,N_18842);
nand UO_688 (O_688,N_20410,N_19766);
xor UO_689 (O_689,N_21591,N_19405);
nor UO_690 (O_690,N_23558,N_21950);
or UO_691 (O_691,N_24660,N_24713);
and UO_692 (O_692,N_23338,N_23778);
nor UO_693 (O_693,N_21269,N_24710);
xnor UO_694 (O_694,N_19840,N_22210);
and UO_695 (O_695,N_24086,N_24607);
nand UO_696 (O_696,N_18852,N_21795);
nor UO_697 (O_697,N_20624,N_21496);
and UO_698 (O_698,N_22611,N_19337);
nand UO_699 (O_699,N_21934,N_20876);
nor UO_700 (O_700,N_23190,N_20725);
nand UO_701 (O_701,N_19109,N_21160);
or UO_702 (O_702,N_19889,N_20520);
xor UO_703 (O_703,N_19791,N_24281);
nor UO_704 (O_704,N_21328,N_19300);
nor UO_705 (O_705,N_19971,N_21980);
nor UO_706 (O_706,N_22077,N_23316);
xnor UO_707 (O_707,N_21984,N_19488);
nand UO_708 (O_708,N_22475,N_21101);
and UO_709 (O_709,N_22459,N_21180);
nand UO_710 (O_710,N_23220,N_19369);
and UO_711 (O_711,N_19434,N_19566);
nor UO_712 (O_712,N_23536,N_23223);
or UO_713 (O_713,N_21342,N_23599);
nor UO_714 (O_714,N_21247,N_22596);
nand UO_715 (O_715,N_21813,N_22192);
or UO_716 (O_716,N_20530,N_21459);
nand UO_717 (O_717,N_22176,N_24185);
xor UO_718 (O_718,N_23330,N_24822);
nor UO_719 (O_719,N_20011,N_21836);
xnor UO_720 (O_720,N_24840,N_22609);
nand UO_721 (O_721,N_22129,N_19654);
nor UO_722 (O_722,N_20411,N_21136);
and UO_723 (O_723,N_19116,N_23469);
nand UO_724 (O_724,N_23507,N_23782);
nand UO_725 (O_725,N_19252,N_22285);
nand UO_726 (O_726,N_19129,N_20596);
nand UO_727 (O_727,N_20012,N_21410);
nor UO_728 (O_728,N_22809,N_21974);
and UO_729 (O_729,N_19444,N_20327);
nand UO_730 (O_730,N_19899,N_24635);
or UO_731 (O_731,N_23389,N_22517);
or UO_732 (O_732,N_24295,N_22450);
and UO_733 (O_733,N_19028,N_23652);
nand UO_734 (O_734,N_19050,N_21062);
or UO_735 (O_735,N_19173,N_20926);
nor UO_736 (O_736,N_21542,N_23562);
nor UO_737 (O_737,N_23095,N_22030);
nand UO_738 (O_738,N_21236,N_23318);
and UO_739 (O_739,N_24817,N_22282);
nor UO_740 (O_740,N_20864,N_24731);
or UO_741 (O_741,N_20203,N_20175);
or UO_742 (O_742,N_21833,N_20461);
nand UO_743 (O_743,N_18931,N_24133);
nand UO_744 (O_744,N_21462,N_23942);
nor UO_745 (O_745,N_21820,N_24868);
nor UO_746 (O_746,N_24708,N_20775);
nand UO_747 (O_747,N_24406,N_22086);
xnor UO_748 (O_748,N_24247,N_22836);
nor UO_749 (O_749,N_23539,N_20354);
nor UO_750 (O_750,N_20966,N_20832);
or UO_751 (O_751,N_22429,N_18869);
and UO_752 (O_752,N_24318,N_23277);
xor UO_753 (O_753,N_19721,N_22624);
nor UO_754 (O_754,N_22593,N_24644);
nand UO_755 (O_755,N_22061,N_24023);
and UO_756 (O_756,N_20223,N_23816);
or UO_757 (O_757,N_23065,N_22186);
nor UO_758 (O_758,N_21954,N_22533);
or UO_759 (O_759,N_21966,N_19203);
or UO_760 (O_760,N_22693,N_18871);
and UO_761 (O_761,N_21597,N_24393);
xor UO_762 (O_762,N_20614,N_21280);
xor UO_763 (O_763,N_23917,N_22320);
nand UO_764 (O_764,N_21741,N_23609);
xor UO_765 (O_765,N_21313,N_20404);
nor UO_766 (O_766,N_18815,N_19135);
nand UO_767 (O_767,N_21715,N_24388);
and UO_768 (O_768,N_23561,N_22548);
nand UO_769 (O_769,N_21265,N_23291);
and UO_770 (O_770,N_19211,N_24368);
nor UO_771 (O_771,N_24005,N_24381);
xor UO_772 (O_772,N_19790,N_23079);
nor UO_773 (O_773,N_22315,N_18953);
or UO_774 (O_774,N_20032,N_20573);
nand UO_775 (O_775,N_19762,N_23758);
or UO_776 (O_776,N_21730,N_19056);
and UO_777 (O_777,N_22487,N_20749);
nand UO_778 (O_778,N_22029,N_19029);
nor UO_779 (O_779,N_24920,N_23975);
and UO_780 (O_780,N_24464,N_23172);
nor UO_781 (O_781,N_24066,N_24242);
or UO_782 (O_782,N_24225,N_20368);
xnor UO_783 (O_783,N_21343,N_20721);
xor UO_784 (O_784,N_21546,N_20745);
xor UO_785 (O_785,N_19505,N_23191);
and UO_786 (O_786,N_21639,N_22905);
and UO_787 (O_787,N_23462,N_20811);
xnor UO_788 (O_788,N_19597,N_19397);
xnor UO_789 (O_789,N_19005,N_24617);
nor UO_790 (O_790,N_19107,N_18848);
or UO_791 (O_791,N_19298,N_20935);
nand UO_792 (O_792,N_23014,N_24231);
nand UO_793 (O_793,N_22146,N_22255);
or UO_794 (O_794,N_24520,N_19445);
nor UO_795 (O_795,N_20726,N_23849);
and UO_796 (O_796,N_20293,N_20286);
nor UO_797 (O_797,N_23009,N_19683);
or UO_798 (O_798,N_19808,N_23668);
nand UO_799 (O_799,N_20544,N_19664);
and UO_800 (O_800,N_19745,N_23960);
and UO_801 (O_801,N_24645,N_23904);
and UO_802 (O_802,N_23938,N_19921);
and UO_803 (O_803,N_20567,N_23510);
nand UO_804 (O_804,N_22290,N_20339);
or UO_805 (O_805,N_19800,N_21710);
or UO_806 (O_806,N_24293,N_19316);
nor UO_807 (O_807,N_21084,N_19346);
or UO_808 (O_808,N_20249,N_23771);
or UO_809 (O_809,N_23117,N_23933);
xor UO_810 (O_810,N_19424,N_19185);
nand UO_811 (O_811,N_24716,N_21545);
nand UO_812 (O_812,N_18833,N_20405);
xnor UO_813 (O_813,N_20121,N_19742);
xnor UO_814 (O_814,N_23263,N_23675);
nor UO_815 (O_815,N_21827,N_19873);
xor UO_816 (O_816,N_18956,N_20495);
nor UO_817 (O_817,N_19134,N_20671);
or UO_818 (O_818,N_20754,N_23192);
xnor UO_819 (O_819,N_22804,N_22484);
and UO_820 (O_820,N_19112,N_19813);
nand UO_821 (O_821,N_23673,N_21620);
or UO_822 (O_822,N_20683,N_22166);
xnor UO_823 (O_823,N_20118,N_21644);
and UO_824 (O_824,N_24039,N_24874);
and UO_825 (O_825,N_21911,N_21341);
or UO_826 (O_826,N_23978,N_19111);
or UO_827 (O_827,N_23969,N_24741);
nand UO_828 (O_828,N_20197,N_22316);
and UO_829 (O_829,N_22521,N_20803);
or UO_830 (O_830,N_19655,N_19820);
nand UO_831 (O_831,N_22525,N_20574);
nand UO_832 (O_832,N_22121,N_22668);
xor UO_833 (O_833,N_24097,N_23491);
and UO_834 (O_834,N_20219,N_23017);
or UO_835 (O_835,N_20184,N_19538);
xor UO_836 (O_836,N_20549,N_22452);
nand UO_837 (O_837,N_22135,N_23110);
nor UO_838 (O_838,N_22562,N_23124);
xnor UO_839 (O_839,N_23676,N_21262);
nor UO_840 (O_840,N_18758,N_24136);
nor UO_841 (O_841,N_22503,N_23992);
xnor UO_842 (O_842,N_21428,N_24265);
xnor UO_843 (O_843,N_24571,N_20888);
or UO_844 (O_844,N_23836,N_24843);
and UO_845 (O_845,N_21586,N_20235);
nand UO_846 (O_846,N_24943,N_19126);
nand UO_847 (O_847,N_19493,N_19904);
and UO_848 (O_848,N_21889,N_23927);
and UO_849 (O_849,N_24214,N_22501);
nor UO_850 (O_850,N_20916,N_19046);
and UO_851 (O_851,N_20186,N_18994);
nand UO_852 (O_852,N_24928,N_20134);
xor UO_853 (O_853,N_19033,N_20772);
and UO_854 (O_854,N_20758,N_20608);
and UO_855 (O_855,N_19804,N_22401);
xor UO_856 (O_856,N_19247,N_18755);
nor UO_857 (O_857,N_22437,N_21706);
nor UO_858 (O_858,N_21956,N_23173);
and UO_859 (O_859,N_22989,N_23293);
nor UO_860 (O_860,N_20182,N_19385);
and UO_861 (O_861,N_19605,N_20466);
nor UO_862 (O_862,N_24683,N_24324);
or UO_863 (O_863,N_23563,N_24671);
and UO_864 (O_864,N_20557,N_24375);
xnor UO_865 (O_865,N_21453,N_18838);
nor UO_866 (O_866,N_20664,N_23919);
and UO_867 (O_867,N_21482,N_22665);
xnor UO_868 (O_868,N_21753,N_20931);
nand UO_869 (O_869,N_23405,N_20553);
or UO_870 (O_870,N_24119,N_23495);
nand UO_871 (O_871,N_19732,N_23353);
nor UO_872 (O_872,N_20020,N_24618);
nand UO_873 (O_873,N_20100,N_22576);
and UO_874 (O_874,N_19313,N_19821);
and UO_875 (O_875,N_24503,N_24791);
or UO_876 (O_876,N_19835,N_20141);
nor UO_877 (O_877,N_19589,N_24568);
or UO_878 (O_878,N_20075,N_22683);
and UO_879 (O_879,N_21169,N_23339);
nand UO_880 (O_880,N_24901,N_20494);
xnor UO_881 (O_881,N_22954,N_19502);
nor UO_882 (O_882,N_24189,N_22869);
or UO_883 (O_883,N_20342,N_22983);
xnor UO_884 (O_884,N_22169,N_23332);
nor UO_885 (O_885,N_22203,N_19915);
nand UO_886 (O_886,N_20999,N_21449);
nor UO_887 (O_887,N_19071,N_18870);
xor UO_888 (O_888,N_22561,N_21635);
nand UO_889 (O_889,N_24869,N_19853);
nand UO_890 (O_890,N_23819,N_24848);
nand UO_891 (O_891,N_19049,N_24749);
nand UO_892 (O_892,N_23039,N_21279);
and UO_893 (O_893,N_22527,N_19897);
or UO_894 (O_894,N_19318,N_19383);
and UO_895 (O_895,N_19253,N_21024);
and UO_896 (O_896,N_19426,N_22329);
nand UO_897 (O_897,N_21943,N_23998);
nand UO_898 (O_898,N_23163,N_23944);
or UO_899 (O_899,N_18763,N_21760);
nand UO_900 (O_900,N_23496,N_19679);
nand UO_901 (O_901,N_18946,N_19896);
nor UO_902 (O_902,N_22570,N_21856);
xnor UO_903 (O_903,N_23947,N_20712);
nand UO_904 (O_904,N_21705,N_24167);
xor UO_905 (O_905,N_20409,N_23787);
nor UO_906 (O_906,N_19396,N_20865);
nand UO_907 (O_907,N_21301,N_20720);
xnor UO_908 (O_908,N_19214,N_22038);
nand UO_909 (O_909,N_23519,N_19715);
xor UO_910 (O_910,N_20432,N_18874);
xnor UO_911 (O_911,N_21337,N_19890);
and UO_912 (O_912,N_21804,N_20233);
nor UO_913 (O_913,N_22540,N_20958);
and UO_914 (O_914,N_19839,N_22435);
and UO_915 (O_915,N_18928,N_23037);
nand UO_916 (O_916,N_23031,N_22544);
and UO_917 (O_917,N_23973,N_21679);
or UO_918 (O_918,N_23941,N_21195);
nor UO_919 (O_919,N_22455,N_23762);
nor UO_920 (O_920,N_20275,N_22660);
or UO_921 (O_921,N_22817,N_23559);
nor UO_922 (O_922,N_21315,N_20398);
and UO_923 (O_923,N_19395,N_20751);
xnor UO_924 (O_924,N_23127,N_21520);
and UO_925 (O_925,N_20743,N_20055);
or UO_926 (O_926,N_21773,N_24830);
or UO_927 (O_927,N_23436,N_21718);
nand UO_928 (O_928,N_19756,N_19966);
and UO_929 (O_929,N_22849,N_24513);
nor UO_930 (O_930,N_21229,N_21158);
and UO_931 (O_931,N_20078,N_22446);
or UO_932 (O_932,N_22522,N_22298);
nor UO_933 (O_933,N_20770,N_22784);
nor UO_934 (O_934,N_24796,N_22257);
or UO_935 (O_935,N_23494,N_24949);
xor UO_936 (O_936,N_19681,N_21690);
nor UO_937 (O_937,N_24624,N_21090);
nand UO_938 (O_938,N_22221,N_22040);
or UO_939 (O_939,N_21748,N_24430);
or UO_940 (O_940,N_19224,N_21350);
nand UO_941 (O_941,N_20422,N_21533);
or UO_942 (O_942,N_24864,N_23240);
nand UO_943 (O_943,N_19413,N_18884);
or UO_944 (O_944,N_19295,N_24440);
xor UO_945 (O_945,N_22065,N_20956);
nor UO_946 (O_946,N_20072,N_23207);
or UO_947 (O_947,N_20450,N_20470);
nor UO_948 (O_948,N_19314,N_23092);
nand UO_949 (O_949,N_21162,N_24524);
nor UO_950 (O_950,N_24327,N_23152);
or UO_951 (O_951,N_19267,N_23050);
and UO_952 (O_952,N_23794,N_22348);
nor UO_953 (O_953,N_22022,N_20315);
nor UO_954 (O_954,N_24825,N_22149);
and UO_955 (O_955,N_19559,N_24320);
nand UO_956 (O_956,N_20732,N_18873);
or UO_957 (O_957,N_24154,N_19008);
xnor UO_958 (O_958,N_24625,N_23314);
nor UO_959 (O_959,N_19781,N_22604);
or UO_960 (O_960,N_24134,N_19630);
nand UO_961 (O_961,N_19855,N_24044);
xnor UO_962 (O_962,N_20137,N_19608);
and UO_963 (O_963,N_19565,N_21782);
nand UO_964 (O_964,N_20023,N_24257);
nand UO_965 (O_965,N_24677,N_21458);
and UO_966 (O_966,N_24402,N_22469);
nor UO_967 (O_967,N_24354,N_22001);
xnor UO_968 (O_968,N_23863,N_24827);
nand UO_969 (O_969,N_24685,N_21316);
nand UO_970 (O_970,N_20649,N_20526);
nand UO_971 (O_971,N_20147,N_22420);
nand UO_972 (O_972,N_22443,N_24890);
xor UO_973 (O_973,N_20734,N_23419);
and UO_974 (O_974,N_21857,N_19440);
or UO_975 (O_975,N_20802,N_22271);
xor UO_976 (O_976,N_24463,N_21370);
xor UO_977 (O_977,N_19093,N_23612);
xor UO_978 (O_978,N_19770,N_23567);
or UO_979 (O_979,N_20539,N_23929);
or UO_980 (O_980,N_22694,N_22984);
and UO_981 (O_981,N_21527,N_20817);
nand UO_982 (O_982,N_19641,N_23988);
and UO_983 (O_983,N_21551,N_20340);
or UO_984 (O_984,N_22157,N_24633);
nand UO_985 (O_985,N_21590,N_21327);
nand UO_986 (O_986,N_18960,N_20503);
and UO_987 (O_987,N_22547,N_22669);
nand UO_988 (O_988,N_19374,N_22920);
nor UO_989 (O_989,N_19532,N_24923);
nand UO_990 (O_990,N_23333,N_21465);
nand UO_991 (O_991,N_19862,N_21220);
xnor UO_992 (O_992,N_23898,N_20540);
nand UO_993 (O_993,N_24414,N_23417);
nor UO_994 (O_994,N_19523,N_21983);
or UO_995 (O_995,N_23742,N_22431);
or UO_996 (O_996,N_22573,N_24996);
and UO_997 (O_997,N_22552,N_22362);
nor UO_998 (O_998,N_23055,N_22046);
or UO_999 (O_999,N_19113,N_19925);
and UO_1000 (O_1000,N_19102,N_20152);
xnor UO_1001 (O_1001,N_20457,N_22430);
xor UO_1002 (O_1002,N_19361,N_22974);
nand UO_1003 (O_1003,N_20612,N_21320);
nor UO_1004 (O_1004,N_18868,N_20730);
nor UO_1005 (O_1005,N_21881,N_24303);
and UO_1006 (O_1006,N_21134,N_24338);
nand UO_1007 (O_1007,N_24301,N_18791);
xnor UO_1008 (O_1008,N_23493,N_22120);
nand UO_1009 (O_1009,N_24346,N_22599);
or UO_1010 (O_1010,N_22309,N_23313);
nand UO_1011 (O_1011,N_22650,N_19013);
nor UO_1012 (O_1012,N_23209,N_23404);
nor UO_1013 (O_1013,N_19002,N_24555);
nand UO_1014 (O_1014,N_20169,N_18967);
and UO_1015 (O_1015,N_24820,N_23568);
or UO_1016 (O_1016,N_22776,N_19195);
nor UO_1017 (O_1017,N_23011,N_23399);
or UO_1018 (O_1018,N_23088,N_24140);
nor UO_1019 (O_1019,N_24111,N_24985);
nand UO_1020 (O_1020,N_19574,N_20243);
nor UO_1021 (O_1021,N_21693,N_21908);
nand UO_1022 (O_1022,N_19543,N_21994);
nand UO_1023 (O_1023,N_22893,N_18900);
nor UO_1024 (O_1024,N_22549,N_21668);
or UO_1025 (O_1025,N_19317,N_24613);
and UO_1026 (O_1026,N_23844,N_20508);
and UO_1027 (O_1027,N_21716,N_23689);
or UO_1028 (O_1028,N_24358,N_23751);
and UO_1029 (O_1029,N_19365,N_22783);
or UO_1030 (O_1030,N_21152,N_24249);
nor UO_1031 (O_1031,N_19264,N_20346);
xor UO_1032 (O_1032,N_23962,N_24855);
nand UO_1033 (O_1033,N_21967,N_21145);
nor UO_1034 (O_1034,N_19435,N_19045);
or UO_1035 (O_1035,N_21746,N_20925);
or UO_1036 (O_1036,N_21243,N_20273);
xnor UO_1037 (O_1037,N_20338,N_20091);
xor UO_1038 (O_1038,N_20431,N_22407);
xor UO_1039 (O_1039,N_18761,N_19170);
xor UO_1040 (O_1040,N_24905,N_19774);
nor UO_1041 (O_1041,N_19431,N_24347);
nor UO_1042 (O_1042,N_21526,N_21205);
xor UO_1043 (O_1043,N_19828,N_19888);
nor UO_1044 (O_1044,N_19955,N_21245);
nand UO_1045 (O_1045,N_20002,N_20418);
xor UO_1046 (O_1046,N_20752,N_20066);
xnor UO_1047 (O_1047,N_23554,N_20892);
or UO_1048 (O_1048,N_21099,N_22014);
xnor UO_1049 (O_1049,N_22854,N_24184);
xor UO_1050 (O_1050,N_20158,N_19297);
xnor UO_1051 (O_1051,N_22163,N_19438);
nor UO_1052 (O_1052,N_19631,N_23835);
or UO_1053 (O_1053,N_20890,N_23428);
nor UO_1054 (O_1054,N_20933,N_19087);
xor UO_1055 (O_1055,N_24726,N_24043);
nor UO_1056 (O_1056,N_22642,N_23555);
xnor UO_1057 (O_1057,N_21659,N_22326);
nor UO_1058 (O_1058,N_23362,N_21631);
or UO_1059 (O_1059,N_20427,N_24482);
nand UO_1060 (O_1060,N_21251,N_23986);
nand UO_1061 (O_1061,N_24029,N_24457);
nor UO_1062 (O_1062,N_22991,N_19776);
nand UO_1063 (O_1063,N_20533,N_24802);
xnor UO_1064 (O_1064,N_19404,N_23572);
or UO_1065 (O_1065,N_21481,N_24646);
and UO_1066 (O_1066,N_24723,N_20918);
and UO_1067 (O_1067,N_22598,N_22910);
nand UO_1068 (O_1068,N_20176,N_20560);
xnor UO_1069 (O_1069,N_18828,N_22933);
xor UO_1070 (O_1070,N_22993,N_20962);
xor UO_1071 (O_1071,N_22909,N_23630);
nand UO_1072 (O_1072,N_24946,N_19079);
and UO_1073 (O_1073,N_21387,N_18768);
nor UO_1074 (O_1074,N_22943,N_21133);
and UO_1075 (O_1075,N_21171,N_21352);
or UO_1076 (O_1076,N_24417,N_22369);
and UO_1077 (O_1077,N_23627,N_24326);
nor UO_1078 (O_1078,N_24828,N_18947);
nor UO_1079 (O_1079,N_20757,N_19196);
nand UO_1080 (O_1080,N_19294,N_22519);
or UO_1081 (O_1081,N_23744,N_20881);
or UO_1082 (O_1082,N_23104,N_23060);
nand UO_1083 (O_1083,N_22144,N_21751);
xor UO_1084 (O_1084,N_19663,N_24207);
and UO_1085 (O_1085,N_20419,N_21529);
and UO_1086 (O_1086,N_19534,N_20672);
nor UO_1087 (O_1087,N_23786,N_23045);
and UO_1088 (O_1088,N_20866,N_23257);
xor UO_1089 (O_1089,N_22386,N_21225);
nor UO_1090 (O_1090,N_19011,N_19388);
nor UO_1091 (O_1091,N_21025,N_22104);
and UO_1092 (O_1092,N_20376,N_22448);
xor UO_1093 (O_1093,N_23287,N_20682);
or UO_1094 (O_1094,N_23925,N_20654);
or UO_1095 (O_1095,N_22841,N_22535);
or UO_1096 (O_1096,N_19281,N_24546);
and UO_1097 (O_1097,N_22375,N_19507);
nor UO_1098 (O_1098,N_19846,N_20412);
nor UO_1099 (O_1099,N_20633,N_21185);
or UO_1100 (O_1100,N_19719,N_21755);
and UO_1101 (O_1101,N_20216,N_20564);
nand UO_1102 (O_1102,N_22099,N_23187);
or UO_1103 (O_1103,N_23618,N_21001);
or UO_1104 (O_1104,N_21425,N_21416);
or UO_1105 (O_1105,N_19210,N_19947);
or UO_1106 (O_1106,N_18922,N_23194);
and UO_1107 (O_1107,N_21218,N_23390);
and UO_1108 (O_1108,N_18818,N_19578);
xnor UO_1109 (O_1109,N_20536,N_22288);
nand UO_1110 (O_1110,N_20534,N_20658);
nor UO_1111 (O_1111,N_23783,N_24891);
xor UO_1112 (O_1112,N_24752,N_22743);
nand UO_1113 (O_1113,N_21298,N_20112);
or UO_1114 (O_1114,N_20038,N_23590);
nor UO_1115 (O_1115,N_21875,N_20359);
xnor UO_1116 (O_1116,N_20008,N_24459);
or UO_1117 (O_1117,N_24480,N_24229);
and UO_1118 (O_1118,N_23985,N_19325);
nor UO_1119 (O_1119,N_21051,N_24115);
nand UO_1120 (O_1120,N_23391,N_23032);
nor UO_1121 (O_1121,N_23882,N_18913);
or UO_1122 (O_1122,N_21761,N_23746);
nand UO_1123 (O_1123,N_22218,N_22768);
and UO_1124 (O_1124,N_21222,N_23224);
xor UO_1125 (O_1125,N_22332,N_24236);
and UO_1126 (O_1126,N_20750,N_20117);
nand UO_1127 (O_1127,N_23500,N_24548);
and UO_1128 (O_1128,N_21061,N_20965);
nand UO_1129 (O_1129,N_24032,N_22960);
or UO_1130 (O_1130,N_20205,N_20981);
xnor UO_1131 (O_1131,N_19454,N_20330);
xnor UO_1132 (O_1132,N_22424,N_20970);
and UO_1133 (O_1133,N_19969,N_23228);
or UO_1134 (O_1134,N_24778,N_22913);
nand UO_1135 (O_1135,N_18804,N_21210);
xnor UO_1136 (O_1136,N_23023,N_19266);
or UO_1137 (O_1137,N_23445,N_20652);
nor UO_1138 (O_1138,N_19090,N_24232);
and UO_1139 (O_1139,N_20934,N_23503);
and UO_1140 (O_1140,N_21201,N_23971);
nand UO_1141 (O_1141,N_24009,N_23573);
xor UO_1142 (O_1142,N_21070,N_23424);
nor UO_1143 (O_1143,N_22620,N_19958);
or UO_1144 (O_1144,N_20819,N_21774);
nor UO_1145 (O_1145,N_19305,N_20215);
xor UO_1146 (O_1146,N_22509,N_20103);
or UO_1147 (O_1147,N_22213,N_19908);
xor UO_1148 (O_1148,N_24512,N_20133);
or UO_1149 (O_1149,N_22748,N_23182);
xnor UO_1150 (O_1150,N_24190,N_21933);
xor UO_1151 (O_1151,N_21083,N_20764);
xnor UO_1152 (O_1152,N_19199,N_23834);
xor UO_1153 (O_1153,N_21922,N_22177);
nand UO_1154 (O_1154,N_24436,N_24372);
nand UO_1155 (O_1155,N_24861,N_19122);
xnor UO_1156 (O_1156,N_24523,N_20125);
or UO_1157 (O_1157,N_19911,N_24439);
or UO_1158 (O_1158,N_24250,N_18933);
nand UO_1159 (O_1159,N_24994,N_23659);
nor UO_1160 (O_1160,N_21606,N_21657);
nand UO_1161 (O_1161,N_19449,N_24233);
or UO_1162 (O_1162,N_22308,N_21495);
nand UO_1163 (O_1163,N_22396,N_21688);
xnor UO_1164 (O_1164,N_20546,N_23219);
nor UO_1165 (O_1165,N_22787,N_21075);
nor UO_1166 (O_1166,N_21576,N_20019);
and UO_1167 (O_1167,N_22168,N_23604);
and UO_1168 (O_1168,N_21986,N_23213);
or UO_1169 (O_1169,N_21565,N_23497);
and UO_1170 (O_1170,N_21548,N_22937);
nor UO_1171 (O_1171,N_24851,N_21098);
and UO_1172 (O_1172,N_21650,N_24712);
nand UO_1173 (O_1173,N_20744,N_23259);
xor UO_1174 (O_1174,N_24627,N_21177);
nand UO_1175 (O_1175,N_21839,N_18888);
xor UO_1176 (O_1176,N_23713,N_21199);
nor UO_1177 (O_1177,N_21299,N_22202);
nor UO_1178 (O_1178,N_23275,N_24908);
nand UO_1179 (O_1179,N_22610,N_18809);
or UO_1180 (O_1180,N_19289,N_22366);
and UO_1181 (O_1181,N_23866,N_19497);
and UO_1182 (O_1182,N_19487,N_19972);
nand UO_1183 (O_1183,N_19973,N_20505);
xnor UO_1184 (O_1184,N_22058,N_20030);
nor UO_1185 (O_1185,N_21487,N_23144);
and UO_1186 (O_1186,N_23183,N_23102);
or UO_1187 (O_1187,N_20781,N_23479);
and UO_1188 (O_1188,N_24240,N_22805);
and UO_1189 (O_1189,N_24481,N_22957);
nor UO_1190 (O_1190,N_19865,N_22087);
nand UO_1191 (O_1191,N_22608,N_19585);
nand UO_1192 (O_1192,N_24467,N_19251);
xnor UO_1193 (O_1193,N_22363,N_18893);
nor UO_1194 (O_1194,N_22337,N_22339);
nor UO_1195 (O_1195,N_21079,N_19163);
xnor UO_1196 (O_1196,N_23547,N_23279);
nand UO_1197 (O_1197,N_23000,N_24128);
or UO_1198 (O_1198,N_21321,N_23595);
nor UO_1199 (O_1199,N_20392,N_21677);
nand UO_1200 (O_1200,N_23476,N_22844);
or UO_1201 (O_1201,N_20185,N_21558);
nor UO_1202 (O_1202,N_20588,N_19524);
nand UO_1203 (O_1203,N_23756,N_23505);
or UO_1204 (O_1204,N_24199,N_20532);
nand UO_1205 (O_1205,N_21081,N_24343);
xnor UO_1206 (O_1206,N_24722,N_23054);
nor UO_1207 (O_1207,N_21009,N_22017);
nor UO_1208 (O_1208,N_19682,N_24220);
or UO_1209 (O_1209,N_23669,N_22733);
xnor UO_1210 (O_1210,N_22868,N_23407);
or UO_1211 (O_1211,N_24941,N_22307);
and UO_1212 (O_1212,N_20762,N_19703);
xor UO_1213 (O_1213,N_22807,N_18886);
nor UO_1214 (O_1214,N_21947,N_20138);
or UO_1215 (O_1215,N_24770,N_20068);
nand UO_1216 (O_1216,N_22786,N_22231);
and UO_1217 (O_1217,N_21414,N_19022);
nand UO_1218 (O_1218,N_23520,N_23278);
xor UO_1219 (O_1219,N_20676,N_20841);
and UO_1220 (O_1220,N_20590,N_24510);
nor UO_1221 (O_1221,N_20917,N_21348);
or UO_1222 (O_1222,N_22262,N_21992);
and UO_1223 (O_1223,N_22189,N_23361);
nand UO_1224 (O_1224,N_23140,N_19986);
nand UO_1225 (O_1225,N_24409,N_20669);
and UO_1226 (O_1226,N_22273,N_22185);
nor UO_1227 (O_1227,N_22081,N_20940);
nor UO_1228 (O_1228,N_19792,N_19927);
nand UO_1229 (O_1229,N_19386,N_21890);
and UO_1230 (O_1230,N_19705,N_24042);
nand UO_1231 (O_1231,N_19114,N_23959);
nor UO_1232 (O_1232,N_19531,N_23608);
and UO_1233 (O_1233,N_24215,N_22471);
nand UO_1234 (O_1234,N_20454,N_22474);
nor UO_1235 (O_1235,N_19024,N_21294);
xor UO_1236 (O_1236,N_22414,N_20257);
and UO_1237 (O_1237,N_18771,N_20379);
nand UO_1238 (O_1238,N_24331,N_22646);
nor UO_1239 (O_1239,N_22524,N_19443);
nand UO_1240 (O_1240,N_20696,N_20510);
nand UO_1241 (O_1241,N_23295,N_21429);
nand UO_1242 (O_1242,N_22398,N_23266);
nand UO_1243 (O_1243,N_20015,N_22075);
xnor UO_1244 (O_1244,N_21122,N_23574);
xnor UO_1245 (O_1245,N_21598,N_20329);
or UO_1246 (O_1246,N_22067,N_20527);
nor UO_1247 (O_1247,N_20455,N_21502);
or UO_1248 (O_1248,N_24291,N_23879);
xnor UO_1249 (O_1249,N_19489,N_22138);
xor UO_1250 (O_1250,N_19220,N_19945);
xnor UO_1251 (O_1251,N_22518,N_23760);
nor UO_1252 (O_1252,N_21290,N_22447);
or UO_1253 (O_1253,N_21579,N_20110);
or UO_1254 (O_1254,N_21941,N_23426);
nor UO_1255 (O_1255,N_24093,N_24470);
xnor UO_1256 (O_1256,N_21903,N_22098);
nor UO_1257 (O_1257,N_22775,N_19653);
nor UO_1258 (O_1258,N_21059,N_21556);
xor UO_1259 (O_1259,N_22785,N_21877);
nand UO_1260 (O_1260,N_24013,N_22280);
or UO_1261 (O_1261,N_20381,N_19803);
nand UO_1262 (O_1262,N_20842,N_19255);
or UO_1263 (O_1263,N_20978,N_20469);
or UO_1264 (O_1264,N_19165,N_21493);
nor UO_1265 (O_1265,N_22403,N_19702);
or UO_1266 (O_1266,N_19164,N_21865);
xor UO_1267 (O_1267,N_24998,N_24028);
or UO_1268 (O_1268,N_23466,N_20625);
or UO_1269 (O_1269,N_19917,N_19864);
and UO_1270 (O_1270,N_22342,N_19044);
or UO_1271 (O_1271,N_21850,N_22201);
nand UO_1272 (O_1272,N_20407,N_22681);
nor UO_1273 (O_1273,N_20480,N_20597);
xnor UO_1274 (O_1274,N_24081,N_19096);
and UO_1275 (O_1275,N_21135,N_20514);
or UO_1276 (O_1276,N_20096,N_24122);
and UO_1277 (O_1277,N_21058,N_21471);
nand UO_1278 (O_1278,N_20621,N_19380);
nand UO_1279 (O_1279,N_20253,N_19462);
and UO_1280 (O_1280,N_20736,N_19003);
nor UO_1281 (O_1281,N_23185,N_22159);
nor UO_1282 (O_1282,N_22615,N_22133);
or UO_1283 (O_1283,N_19937,N_19261);
nand UO_1284 (O_1284,N_21190,N_21293);
nand UO_1285 (O_1285,N_22513,N_22449);
nor UO_1286 (O_1286,N_22268,N_24541);
xnor UO_1287 (O_1287,N_21815,N_22982);
or UO_1288 (O_1288,N_24823,N_23687);
and UO_1289 (O_1289,N_24812,N_18834);
nor UO_1290 (O_1290,N_23934,N_24008);
and UO_1291 (O_1291,N_20382,N_18912);
nor UO_1292 (O_1292,N_20521,N_20611);
nor UO_1293 (O_1293,N_23535,N_19879);
xor UO_1294 (O_1294,N_21998,N_22923);
xor UO_1295 (O_1295,N_21981,N_21226);
xnor UO_1296 (O_1296,N_24667,N_21863);
or UO_1297 (O_1297,N_19007,N_18823);
nand UO_1298 (O_1298,N_22208,N_21113);
and UO_1299 (O_1299,N_24151,N_21435);
xnor UO_1300 (O_1300,N_19901,N_23222);
xor UO_1301 (O_1301,N_22627,N_24807);
nor UO_1302 (O_1302,N_23853,N_23877);
nand UO_1303 (O_1303,N_22861,N_19309);
and UO_1304 (O_1304,N_23432,N_19188);
or UO_1305 (O_1305,N_21221,N_22955);
nor UO_1306 (O_1306,N_24915,N_22758);
nand UO_1307 (O_1307,N_24490,N_19570);
xor UO_1308 (O_1308,N_19437,N_22745);
or UO_1309 (O_1309,N_21672,N_23912);
and UO_1310 (O_1310,N_18901,N_20255);
and UO_1311 (O_1311,N_23499,N_21124);
xor UO_1312 (O_1312,N_19644,N_23276);
or UO_1313 (O_1313,N_22109,N_23492);
or UO_1314 (O_1314,N_20963,N_24987);
nand UO_1315 (O_1315,N_20177,N_23663);
and UO_1316 (O_1316,N_24737,N_21687);
nor UO_1317 (O_1317,N_24153,N_21924);
or UO_1318 (O_1318,N_24961,N_21503);
and UO_1319 (O_1319,N_23977,N_24361);
or UO_1320 (O_1320,N_23025,N_20402);
nand UO_1321 (O_1321,N_21951,N_21492);
nand UO_1322 (O_1322,N_23790,N_24809);
nor UO_1323 (O_1323,N_22234,N_23103);
or UO_1324 (O_1324,N_19749,N_24967);
nor UO_1325 (O_1325,N_19692,N_23894);
or UO_1326 (O_1326,N_19819,N_21583);
nand UO_1327 (O_1327,N_22009,N_22986);
nand UO_1328 (O_1328,N_19836,N_23211);
nor UO_1329 (O_1329,N_21664,N_23292);
nand UO_1330 (O_1330,N_19015,N_23871);
or UO_1331 (O_1331,N_21717,N_24728);
or UO_1332 (O_1332,N_21792,N_22152);
nand UO_1333 (O_1333,N_22917,N_19647);
and UO_1334 (O_1334,N_22080,N_22174);
and UO_1335 (O_1335,N_22929,N_24799);
nand UO_1336 (O_1336,N_24587,N_23403);
nand UO_1337 (O_1337,N_21478,N_20742);
nor UO_1338 (O_1338,N_18836,N_24889);
or UO_1339 (O_1339,N_21821,N_24157);
nor UO_1340 (O_1340,N_19714,N_19642);
and UO_1341 (O_1341,N_19171,N_24614);
and UO_1342 (O_1342,N_20295,N_19886);
or UO_1343 (O_1343,N_22820,N_23920);
nor UO_1344 (O_1344,N_21517,N_21948);
xor UO_1345 (O_1345,N_22248,N_23984);
xor UO_1346 (O_1346,N_24727,N_18951);
or UO_1347 (O_1347,N_23340,N_21888);
and UO_1348 (O_1348,N_19893,N_21213);
nor UO_1349 (O_1349,N_21010,N_20296);
xnor UO_1350 (O_1350,N_18786,N_23026);
and UO_1351 (O_1351,N_19837,N_20748);
nand UO_1352 (O_1352,N_22359,N_21961);
nand UO_1353 (O_1353,N_20569,N_23071);
nor UO_1354 (O_1354,N_22460,N_22578);
nand UO_1355 (O_1355,N_24290,N_23901);
and UO_1356 (O_1356,N_18830,N_23804);
or UO_1357 (O_1357,N_19054,N_20474);
nor UO_1358 (O_1358,N_24325,N_20371);
or UO_1359 (O_1359,N_21783,N_18810);
nor UO_1360 (O_1360,N_24304,N_20620);
nor UO_1361 (O_1361,N_22708,N_21346);
nor UO_1362 (O_1362,N_23989,N_23372);
nand UO_1363 (O_1363,N_20397,N_23703);
nor UO_1364 (O_1364,N_19697,N_22136);
xor UO_1365 (O_1365,N_19861,N_20481);
or UO_1366 (O_1366,N_18896,N_21952);
nand UO_1367 (O_1367,N_20144,N_19127);
nand UO_1368 (O_1368,N_20244,N_24068);
and UO_1369 (O_1369,N_20375,N_23598);
or UO_1370 (O_1370,N_24927,N_19509);
or UO_1371 (O_1371,N_22619,N_19739);
nand UO_1372 (O_1372,N_24323,N_24887);
and UO_1373 (O_1373,N_22411,N_22085);
nor UO_1374 (O_1374,N_21358,N_22709);
xor UO_1375 (O_1375,N_22996,N_22235);
nor UO_1376 (O_1376,N_19688,N_24648);
xor UO_1377 (O_1377,N_21187,N_21735);
or UO_1378 (O_1378,N_23769,N_23648);
nand UO_1379 (O_1379,N_18972,N_23354);
nor UO_1380 (O_1380,N_21539,N_24391);
xnor UO_1381 (O_1381,N_19602,N_19226);
nand UO_1382 (O_1382,N_23463,N_24170);
nor UO_1383 (O_1383,N_23073,N_24879);
and UO_1384 (O_1384,N_23446,N_20191);
nand UO_1385 (O_1385,N_19436,N_19097);
nor UO_1386 (O_1386,N_23822,N_20274);
nand UO_1387 (O_1387,N_24308,N_22445);
nor UO_1388 (O_1388,N_20818,N_19120);
or UO_1389 (O_1389,N_23013,N_21163);
and UO_1390 (O_1390,N_21613,N_24130);
nor UO_1391 (O_1391,N_21663,N_18855);
nand UO_1392 (O_1392,N_20902,N_22618);
nand UO_1393 (O_1393,N_23123,N_20350);
xor UO_1394 (O_1394,N_21053,N_23489);
and UO_1395 (O_1395,N_19620,N_20263);
and UO_1396 (O_1396,N_21897,N_21434);
nand UO_1397 (O_1397,N_20154,N_23289);
xor UO_1398 (O_1398,N_21628,N_24312);
or UO_1399 (O_1399,N_21326,N_22655);
nor UO_1400 (O_1400,N_20026,N_20352);
and UO_1401 (O_1401,N_24602,N_18861);
and UO_1402 (O_1402,N_22183,N_19628);
or UO_1403 (O_1403,N_19661,N_20995);
xor UO_1404 (O_1404,N_20728,N_20280);
nor UO_1405 (O_1405,N_20846,N_24814);
nand UO_1406 (O_1406,N_20984,N_20632);
and UO_1407 (O_1407,N_22674,N_21808);
xnor UO_1408 (O_1408,N_21780,N_18802);
xnor UO_1409 (O_1409,N_21000,N_21835);
and UO_1410 (O_1410,N_23051,N_24270);
or UO_1411 (O_1411,N_18784,N_24376);
or UO_1412 (O_1412,N_20554,N_20704);
nand UO_1413 (O_1413,N_23701,N_20486);
nor UO_1414 (O_1414,N_24763,N_19427);
nor UO_1415 (O_1415,N_22944,N_19660);
nand UO_1416 (O_1416,N_21181,N_23781);
nand UO_1417 (O_1417,N_20908,N_22444);
or UO_1418 (O_1418,N_23601,N_21580);
or UO_1419 (O_1419,N_22595,N_19744);
nor UO_1420 (O_1420,N_20674,N_21826);
and UO_1421 (O_1421,N_23583,N_24947);
or UO_1422 (O_1422,N_23828,N_23317);
or UO_1423 (O_1423,N_22270,N_19225);
nand UO_1424 (O_1424,N_23589,N_24046);
nand UO_1425 (O_1425,N_22685,N_22442);
or UO_1426 (O_1426,N_20344,N_18799);
nand UO_1427 (O_1427,N_22892,N_22543);
nand UO_1428 (O_1428,N_24824,N_23761);
and UO_1429 (O_1429,N_24688,N_20193);
or UO_1430 (O_1430,N_24001,N_20492);
nand UO_1431 (O_1431,N_24897,N_21880);
and UO_1432 (O_1432,N_24020,N_24867);
xor UO_1433 (O_1433,N_20071,N_23272);
nor UO_1434 (O_1434,N_19709,N_22293);
and UO_1435 (O_1435,N_20321,N_19763);
nor UO_1436 (O_1436,N_19393,N_21017);
xor UO_1437 (O_1437,N_24098,N_19055);
nand UO_1438 (O_1438,N_19235,N_20265);
nand UO_1439 (O_1439,N_19514,N_23776);
nand UO_1440 (O_1440,N_20081,N_20681);
nor UO_1441 (O_1441,N_20586,N_19254);
and UO_1442 (O_1442,N_20824,N_24896);
or UO_1443 (O_1443,N_22190,N_24786);
and UO_1444 (O_1444,N_20957,N_22353);
nor UO_1445 (O_1445,N_21610,N_24704);
nand UO_1446 (O_1446,N_22319,N_21665);
or UO_1447 (O_1447,N_21271,N_18976);
xor UO_1448 (O_1448,N_23591,N_22632);
and UO_1449 (O_1449,N_20156,N_18989);
nand UO_1450 (O_1450,N_24274,N_23234);
nor UO_1451 (O_1451,N_20879,N_22406);
or UO_1452 (O_1452,N_22751,N_22314);
nor UO_1453 (O_1453,N_19657,N_20980);
nand UO_1454 (O_1454,N_20844,N_21834);
nor UO_1455 (O_1455,N_23109,N_23461);
xor UO_1456 (O_1456,N_22220,N_20311);
nor UO_1457 (O_1457,N_24437,N_21491);
xnor UO_1458 (O_1458,N_20230,N_24403);
nor UO_1459 (O_1459,N_19326,N_24052);
xnor UO_1460 (O_1460,N_22799,N_24294);
and UO_1461 (O_1461,N_19614,N_19713);
nand UO_1462 (O_1462,N_18979,N_21757);
or UO_1463 (O_1463,N_24099,N_24700);
and UO_1464 (O_1464,N_20347,N_19562);
nand UO_1465 (O_1465,N_19579,N_22742);
or UO_1466 (O_1466,N_21676,N_23693);
and UO_1467 (O_1467,N_21126,N_18978);
nand UO_1468 (O_1468,N_19954,N_23579);
xnor UO_1469 (O_1469,N_24783,N_19984);
and UO_1470 (O_1470,N_22387,N_20345);
nor UO_1471 (O_1471,N_24601,N_24487);
nand UO_1472 (O_1472,N_23557,N_20854);
xnor UO_1473 (O_1473,N_21324,N_24280);
xnor UO_1474 (O_1474,N_23955,N_23454);
or UO_1475 (O_1475,N_23087,N_24522);
or UO_1476 (O_1476,N_18943,N_21461);
and UO_1477 (O_1477,N_22588,N_23022);
nand UO_1478 (O_1478,N_24447,N_19256);
nand UO_1479 (O_1479,N_22968,N_22806);
and UO_1480 (O_1480,N_21844,N_22200);
nor UO_1481 (O_1481,N_19174,N_20897);
and UO_1482 (O_1482,N_24488,N_22647);
or UO_1483 (O_1483,N_23928,N_19615);
xor UO_1484 (O_1484,N_23680,N_23343);
xnor UO_1485 (O_1485,N_23135,N_20738);
nand UO_1486 (O_1486,N_22170,N_19685);
and UO_1487 (O_1487,N_21419,N_24811);
xnor UO_1488 (O_1488,N_22292,N_22206);
nor UO_1489 (O_1489,N_22978,N_19662);
nor UO_1490 (O_1490,N_20086,N_19939);
or UO_1491 (O_1491,N_22857,N_19708);
and UO_1492 (O_1492,N_21588,N_23937);
nand UO_1493 (O_1493,N_21916,N_19898);
and UO_1494 (O_1494,N_21468,N_20131);
xor UO_1495 (O_1495,N_24095,N_18754);
and UO_1496 (O_1496,N_20438,N_19957);
or UO_1497 (O_1497,N_21148,N_23153);
and UO_1498 (O_1498,N_20093,N_22269);
nor UO_1499 (O_1499,N_23611,N_23739);
nor UO_1500 (O_1500,N_24200,N_22365);
and UO_1501 (O_1501,N_23126,N_18780);
xnor UO_1502 (O_1502,N_22397,N_23086);
nor UO_1503 (O_1503,N_23049,N_23047);
nand UO_1504 (O_1504,N_21363,N_23028);
nor UO_1505 (O_1505,N_21322,N_23083);
or UO_1506 (O_1506,N_24144,N_20284);
or UO_1507 (O_1507,N_24150,N_21276);
or UO_1508 (O_1508,N_24053,N_20525);
nor UO_1509 (O_1509,N_23096,N_23861);
nor UO_1510 (O_1510,N_23736,N_21914);
and UO_1511 (O_1511,N_20801,N_22361);
nand UO_1512 (O_1512,N_19500,N_20077);
nor UO_1513 (O_1513,N_19430,N_22958);
nand UO_1514 (O_1514,N_20835,N_23616);
or UO_1515 (O_1515,N_23132,N_20140);
or UO_1516 (O_1516,N_22252,N_24689);
xnor UO_1517 (O_1517,N_20955,N_24701);
and UO_1518 (O_1518,N_18766,N_20915);
and UO_1519 (O_1519,N_22851,N_22666);
nor UO_1520 (O_1520,N_24952,N_20904);
xnor UO_1521 (O_1521,N_21069,N_20880);
or UO_1522 (O_1522,N_18843,N_22664);
or UO_1523 (O_1523,N_22692,N_20064);
nand UO_1524 (O_1524,N_23890,N_24491);
xnor UO_1525 (O_1525,N_23468,N_23483);
xor UO_1526 (O_1526,N_19675,N_20130);
xor UO_1527 (O_1527,N_22931,N_24534);
or UO_1528 (O_1528,N_21530,N_19099);
or UO_1529 (O_1529,N_23460,N_23522);
xor UO_1530 (O_1530,N_22470,N_23242);
nor UO_1531 (O_1531,N_24499,N_19801);
and UO_1532 (O_1532,N_19162,N_20796);
nand UO_1533 (O_1533,N_22204,N_21131);
and UO_1534 (O_1534,N_24938,N_22141);
or UO_1535 (O_1535,N_21253,N_19213);
xor UO_1536 (O_1536,N_22797,N_21255);
or UO_1537 (O_1537,N_23930,N_20602);
and UO_1538 (O_1538,N_21413,N_21732);
nand UO_1539 (O_1539,N_21057,N_19704);
or UO_1540 (O_1540,N_24445,N_22583);
or UO_1541 (O_1541,N_20647,N_20031);
nand UO_1542 (O_1542,N_21519,N_19687);
nor UO_1543 (O_1543,N_22705,N_23100);
xor UO_1544 (O_1544,N_24884,N_24502);
and UO_1545 (O_1545,N_20292,N_21211);
nand UO_1546 (O_1546,N_24238,N_21304);
or UO_1547 (O_1547,N_22321,N_22497);
xnor UO_1548 (O_1548,N_20459,N_23473);
xnor UO_1549 (O_1549,N_20024,N_24797);
nand UO_1550 (O_1550,N_24852,N_20971);
nand UO_1551 (O_1551,N_19598,N_19460);
and UO_1552 (O_1552,N_18856,N_23939);
xor UO_1553 (O_1553,N_23670,N_18987);
xor UO_1554 (O_1554,N_24082,N_21091);
xnor UO_1555 (O_1555,N_24738,N_24455);
xnor UO_1556 (O_1556,N_21354,N_24771);
or UO_1557 (O_1557,N_19377,N_24588);
nor UO_1558 (O_1558,N_22246,N_18875);
nand UO_1559 (O_1559,N_21200,N_24854);
or UO_1560 (O_1560,N_19718,N_22033);
nand UO_1561 (O_1561,N_21023,N_19060);
nor UO_1562 (O_1562,N_21087,N_22391);
and UO_1563 (O_1563,N_22531,N_23184);
nand UO_1564 (O_1564,N_19516,N_23544);
xnor UO_1565 (O_1565,N_19918,N_22328);
or UO_1566 (O_1566,N_20823,N_22405);
nand UO_1567 (O_1567,N_19115,N_20045);
nand UO_1568 (O_1568,N_22112,N_23241);
or UO_1569 (O_1569,N_21161,N_21499);
nand UO_1570 (O_1570,N_24975,N_23176);
or UO_1571 (O_1571,N_18930,N_20922);
nor UO_1572 (O_1572,N_18919,N_21784);
nor UO_1573 (O_1573,N_19723,N_22657);
nand UO_1574 (O_1574,N_24370,N_22464);
xnor UO_1575 (O_1575,N_24957,N_20178);
nand UO_1576 (O_1576,N_21686,N_23518);
or UO_1577 (O_1577,N_23288,N_19847);
and UO_1578 (O_1578,N_22215,N_24681);
and UO_1579 (O_1579,N_22574,N_24709);
nor UO_1580 (O_1580,N_23899,N_23027);
or UO_1581 (O_1581,N_23578,N_21985);
nand UO_1582 (O_1582,N_24252,N_23335);
nand UO_1583 (O_1583,N_20953,N_21424);
xor UO_1584 (O_1584,N_20281,N_19811);
nand UO_1585 (O_1585,N_20153,N_22226);
nand UO_1586 (O_1586,N_18825,N_24205);
nor UO_1587 (O_1587,N_23995,N_19146);
and UO_1588 (O_1588,N_19153,N_19368);
and UO_1589 (O_1589,N_24424,N_21540);
and UO_1590 (O_1590,N_23180,N_19832);
xor UO_1591 (O_1591,N_21268,N_22774);
xnor UO_1592 (O_1592,N_23911,N_22158);
and UO_1593 (O_1593,N_23294,N_23388);
and UO_1594 (O_1594,N_23875,N_19355);
and UO_1595 (O_1595,N_22423,N_20746);
or UO_1596 (O_1596,N_23082,N_24171);
nor UO_1597 (O_1597,N_24102,N_21666);
or UO_1598 (O_1598,N_21307,N_18879);
xnor UO_1599 (O_1599,N_22981,N_20820);
xnor UO_1600 (O_1600,N_20447,N_22110);
xnor UO_1601 (O_1601,N_21284,N_24146);
nor UO_1602 (O_1602,N_24605,N_21345);
nor UO_1603 (O_1603,N_22881,N_23797);
xnor UO_1604 (O_1604,N_20541,N_20443);
or UO_1605 (O_1605,N_21532,N_18964);
and UO_1606 (O_1606,N_23842,N_23170);
nor UO_1607 (O_1607,N_24330,N_20694);
nand UO_1608 (O_1608,N_19833,N_18921);
xor UO_1609 (O_1609,N_23256,N_22091);
or UO_1610 (O_1610,N_24518,N_22261);
or UO_1611 (O_1611,N_22173,N_24443);
nor UO_1612 (O_1612,N_23070,N_21825);
nand UO_1613 (O_1613,N_24780,N_23981);
or UO_1614 (O_1614,N_24806,N_20771);
and UO_1615 (O_1615,N_23936,N_24641);
nand UO_1616 (O_1616,N_22928,N_24958);
or UO_1617 (O_1617,N_24758,N_23961);
or UO_1618 (O_1618,N_21802,N_23281);
nand UO_1619 (O_1619,N_23171,N_22511);
and UO_1620 (O_1620,N_24248,N_19324);
or UO_1621 (O_1621,N_21978,N_20714);
nor UO_1622 (O_1622,N_24413,N_18881);
nor UO_1623 (O_1623,N_19333,N_20946);
nor UO_1624 (O_1624,N_23725,N_20701);
nand UO_1625 (O_1625,N_24993,N_18812);
xor UO_1626 (O_1626,N_22781,N_19805);
nor UO_1627 (O_1627,N_19546,N_24561);
nand UO_1628 (O_1628,N_23634,N_20451);
xor UO_1629 (O_1629,N_22499,N_20318);
nand UO_1630 (O_1630,N_22451,N_20885);
xnor UO_1631 (O_1631,N_19542,N_21323);
nor UO_1632 (O_1632,N_24147,N_22415);
nor UO_1633 (O_1633,N_20484,N_23870);
or UO_1634 (O_1634,N_24337,N_20769);
nor UO_1635 (O_1635,N_23448,N_23993);
and UO_1636 (O_1636,N_19506,N_19014);
and UO_1637 (O_1637,N_24307,N_23724);
nand UO_1638 (O_1638,N_22710,N_24010);
nand UO_1639 (O_1639,N_24565,N_19826);
or UO_1640 (O_1640,N_21612,N_24552);
xnor UO_1641 (O_1641,N_23740,N_19618);
or UO_1642 (O_1642,N_20634,N_21494);
nand UO_1643 (O_1643,N_24219,N_19753);
nor UO_1644 (O_1644,N_19930,N_21714);
nor UO_1645 (O_1645,N_24649,N_24362);
or UO_1646 (O_1646,N_22260,N_21031);
nor UO_1647 (O_1647,N_21417,N_20319);
nand UO_1648 (O_1648,N_18788,N_19074);
or UO_1649 (O_1649,N_20562,N_18940);
or UO_1650 (O_1650,N_23830,N_19677);
and UO_1651 (O_1651,N_21128,N_19802);
and UO_1652 (O_1652,N_24600,N_21873);
nor UO_1653 (O_1653,N_23076,N_19635);
or UO_1654 (O_1654,N_23004,N_21412);
and UO_1655 (O_1655,N_22766,N_19882);
nor UO_1656 (O_1656,N_22094,N_24784);
or UO_1657 (O_1657,N_21132,N_22191);
or UO_1658 (O_1658,N_24255,N_21423);
and UO_1659 (O_1659,N_20448,N_20170);
or UO_1660 (O_1660,N_24964,N_21562);
nand UO_1661 (O_1661,N_19411,N_23773);
or UO_1662 (O_1662,N_24666,N_24960);
and UO_1663 (O_1663,N_22142,N_24531);
nor UO_1664 (O_1664,N_19348,N_24349);
and UO_1665 (O_1665,N_21309,N_24208);
xor UO_1666 (O_1666,N_21296,N_23264);
and UO_1667 (O_1667,N_19469,N_24016);
xor UO_1668 (O_1668,N_22843,N_20460);
or UO_1669 (O_1669,N_23232,N_21694);
or UO_1670 (O_1670,N_20830,N_24088);
nand UO_1671 (O_1671,N_24695,N_20092);
nand UO_1672 (O_1672,N_21725,N_23711);
and UO_1673 (O_1673,N_18935,N_21518);
and UO_1674 (O_1674,N_19883,N_20462);
xnor UO_1675 (O_1675,N_21772,N_21584);
and UO_1676 (O_1676,N_24966,N_24363);
and UO_1677 (O_1677,N_21671,N_22116);
and UO_1678 (O_1678,N_24913,N_18958);
or UO_1679 (O_1679,N_22323,N_21241);
nor UO_1680 (O_1680,N_19498,N_21314);
and UO_1681 (O_1681,N_20165,N_23312);
and UO_1682 (O_1682,N_23412,N_22027);
nor UO_1683 (O_1683,N_21957,N_18814);
and UO_1684 (O_1684,N_24432,N_23210);
or UO_1685 (O_1685,N_22322,N_23324);
and UO_1686 (O_1686,N_24392,N_19238);
nor UO_1687 (O_1687,N_21096,N_22063);
nand UO_1688 (O_1688,N_20048,N_24732);
or UO_1689 (O_1689,N_22002,N_24847);
and UO_1690 (O_1690,N_24087,N_23189);
nor UO_1691 (O_1691,N_18807,N_24765);
nand UO_1692 (O_1692,N_19149,N_24222);
or UO_1693 (O_1693,N_21658,N_19040);
xor UO_1694 (O_1694,N_21721,N_19755);
nand UO_1695 (O_1695,N_22251,N_21822);
and UO_1696 (O_1696,N_23328,N_23692);
or UO_1697 (O_1697,N_22720,N_23620);
or UO_1698 (O_1698,N_21785,N_21806);
nor UO_1699 (O_1699,N_21020,N_21884);
nand UO_1700 (O_1700,N_23764,N_23811);
nand UO_1701 (O_1701,N_24720,N_18996);
nand UO_1702 (O_1702,N_22355,N_22870);
nand UO_1703 (O_1703,N_19389,N_23881);
nor UO_1704 (O_1704,N_21289,N_21737);
or UO_1705 (O_1705,N_19136,N_23143);
nand UO_1706 (O_1706,N_18941,N_19649);
nand UO_1707 (O_1707,N_23655,N_20939);
and UO_1708 (O_1708,N_20196,N_22603);
xnor UO_1709 (O_1709,N_23052,N_19706);
nor UO_1710 (O_1710,N_19323,N_22345);
or UO_1711 (O_1711,N_22379,N_22690);
xnor UO_1712 (O_1712,N_23571,N_21704);
xnor UO_1713 (O_1713,N_22294,N_19197);
nor UO_1714 (O_1714,N_23366,N_22256);
nor UO_1715 (O_1715,N_24540,N_19328);
xor UO_1716 (O_1716,N_23158,N_23477);
nor UO_1717 (O_1717,N_22563,N_21823);
or UO_1718 (O_1718,N_21629,N_22467);
xnor UO_1719 (O_1719,N_19026,N_22118);
xnor UO_1720 (O_1720,N_19378,N_20763);
nand UO_1721 (O_1721,N_23470,N_22302);
or UO_1722 (O_1722,N_20434,N_22026);
and UO_1723 (O_1723,N_21214,N_23435);
nand UO_1724 (O_1724,N_23007,N_20982);
and UO_1725 (O_1725,N_24460,N_18977);
or UO_1726 (O_1726,N_21238,N_22515);
xor UO_1727 (O_1727,N_23686,N_24669);
nand UO_1728 (O_1728,N_21572,N_22488);
nand UO_1729 (O_1729,N_21593,N_19263);
or UO_1730 (O_1730,N_20062,N_22932);
and UO_1731 (O_1731,N_24024,N_20894);
or UO_1732 (O_1732,N_19470,N_21758);
nor UO_1733 (O_1733,N_22325,N_19701);
xnor UO_1734 (O_1734,N_24045,N_24126);
nor UO_1735 (O_1735,N_22689,N_20326);
or UO_1736 (O_1736,N_19850,N_23829);
or UO_1737 (O_1737,N_22875,N_21633);
and UO_1738 (O_1738,N_21338,N_24818);
or UO_1739 (O_1739,N_24169,N_18760);
or UO_1740 (O_1740,N_20420,N_21266);
and UO_1741 (O_1741,N_23840,N_23360);
nand UO_1742 (O_1742,N_21267,N_20591);
nor UO_1743 (O_1743,N_24599,N_21486);
xnor UO_1744 (O_1744,N_20804,N_24604);
nand UO_1745 (O_1745,N_24059,N_20151);
or UO_1746 (O_1746,N_24692,N_23832);
nand UO_1747 (O_1747,N_18895,N_22479);
nand UO_1748 (O_1748,N_21167,N_19018);
and UO_1749 (O_1749,N_22962,N_22263);
and UO_1750 (O_1750,N_20609,N_24750);
or UO_1751 (O_1751,N_20565,N_24652);
and UO_1752 (O_1752,N_19959,N_19872);
xor UO_1753 (O_1753,N_20688,N_24446);
xnor UO_1754 (O_1754,N_24461,N_19069);
xor UO_1755 (O_1755,N_20766,N_23197);
nand UO_1756 (O_1756,N_24782,N_21191);
or UO_1757 (O_1757,N_24816,N_20098);
xnor UO_1758 (O_1758,N_24733,N_22895);
nand UO_1759 (O_1759,N_21634,N_22041);
and UO_1760 (O_1760,N_21332,N_23838);
nand UO_1761 (O_1761,N_19387,N_23864);
nor UO_1762 (O_1762,N_21917,N_24125);
and UO_1763 (O_1763,N_23681,N_24285);
or UO_1764 (O_1764,N_23945,N_24321);
or UO_1765 (O_1765,N_19417,N_24543);
and UO_1766 (O_1766,N_20774,N_22031);
nand UO_1767 (O_1767,N_24408,N_19525);
xor UO_1768 (O_1768,N_19552,N_19627);
xnor UO_1769 (O_1769,N_23963,N_22147);
xor UO_1770 (O_1770,N_24849,N_19743);
and UO_1771 (O_1771,N_20401,N_20998);
nand UO_1772 (O_1772,N_22179,N_20399);
or UO_1773 (O_1773,N_23056,N_21433);
nand UO_1774 (O_1774,N_21969,N_19352);
nand UO_1775 (O_1775,N_24366,N_20483);
xor UO_1776 (O_1776,N_19919,N_23280);
xnor UO_1777 (O_1777,N_19665,N_21125);
xnor UO_1778 (O_1778,N_22250,N_20615);
xor UO_1779 (O_1779,N_20765,N_22066);
and UO_1780 (O_1780,N_21089,N_19587);
xnor UO_1781 (O_1781,N_23359,N_19590);
and UO_1782 (O_1782,N_22053,N_19793);
nor UO_1783 (O_1783,N_23285,N_24970);
and UO_1784 (O_1784,N_22921,N_21932);
nand UO_1785 (O_1785,N_20785,N_20593);
nand UO_1786 (O_1786,N_20225,N_21691);
nor UO_1787 (O_1787,N_22155,N_20566);
or UO_1788 (O_1788,N_20723,N_23305);
nand UO_1789 (O_1789,N_24950,N_19130);
or UO_1790 (O_1790,N_24535,N_20065);
and UO_1791 (O_1791,N_24856,N_19990);
xnor UO_1792 (O_1792,N_21003,N_21536);
or UO_1793 (O_1793,N_21776,N_19940);
nor UO_1794 (O_1794,N_19372,N_23273);
nand UO_1795 (O_1795,N_23167,N_19580);
xor UO_1796 (O_1796,N_18839,N_22926);
or UO_1797 (O_1797,N_21791,N_19154);
and UO_1798 (O_1798,N_22737,N_18803);
and UO_1799 (O_1799,N_20160,N_20834);
nor UO_1800 (O_1800,N_22502,N_21415);
nand UO_1801 (O_1801,N_20425,N_21030);
nand UO_1802 (O_1802,N_20545,N_21460);
or UO_1803 (O_1803,N_24549,N_21139);
nand UO_1804 (O_1804,N_19291,N_21235);
nor UO_1805 (O_1805,N_24116,N_20446);
nor UO_1806 (O_1806,N_20695,N_19204);
or UO_1807 (O_1807,N_23115,N_22567);
and UO_1808 (O_1808,N_20599,N_21421);
or UO_1809 (O_1809,N_19234,N_22384);
nand UO_1810 (O_1810,N_24289,N_22371);
and UO_1811 (O_1811,N_19880,N_23910);
nand UO_1812 (O_1812,N_19924,N_21347);
nor UO_1813 (O_1813,N_18827,N_22626);
and UO_1814 (O_1814,N_18906,N_20627);
and UO_1815 (O_1815,N_20905,N_22829);
xnor UO_1816 (O_1816,N_20325,N_20568);
nand UO_1817 (O_1817,N_23524,N_18911);
xor UO_1818 (O_1818,N_24040,N_19468);
nor UO_1819 (O_1819,N_19415,N_22082);
nor UO_1820 (O_1820,N_21739,N_20909);
or UO_1821 (O_1821,N_19528,N_24429);
xnor UO_1822 (O_1822,N_24862,N_24135);
nand UO_1823 (O_1823,N_22976,N_21601);
and UO_1824 (O_1824,N_18775,N_23431);
and UO_1825 (O_1825,N_22542,N_20143);
xnor UO_1826 (O_1826,N_22364,N_23629);
or UO_1827 (O_1827,N_21915,N_24743);
or UO_1828 (O_1828,N_21819,N_21809);
or UO_1829 (O_1829,N_23413,N_20895);
xnor UO_1830 (O_1830,N_22291,N_19037);
nor UO_1831 (O_1831,N_19065,N_21467);
xor UO_1832 (O_1832,N_22848,N_20822);
or UO_1833 (O_1833,N_22217,N_19809);
nor UO_1834 (O_1834,N_18999,N_22935);
nor UO_1835 (O_1835,N_23327,N_23869);
or UO_1836 (O_1836,N_22148,N_22633);
nor UO_1837 (O_1837,N_20017,N_22566);
and UO_1838 (O_1838,N_19527,N_20708);
nand UO_1839 (O_1839,N_23674,N_19964);
xor UO_1840 (O_1840,N_20761,N_21837);
xor UO_1841 (O_1841,N_21427,N_20331);
and UO_1842 (O_1842,N_21360,N_22847);
nor UO_1843 (O_1843,N_18894,N_19206);
and UO_1844 (O_1844,N_21305,N_21538);
nor UO_1845 (O_1845,N_22281,N_23815);
nand UO_1846 (O_1846,N_19895,N_21525);
and UO_1847 (O_1847,N_20384,N_21695);
nand UO_1848 (O_1848,N_24521,N_23459);
or UO_1849 (O_1849,N_24311,N_21240);
or UO_1850 (O_1850,N_19603,N_18915);
or UO_1851 (O_1851,N_20855,N_24945);
or UO_1852 (O_1852,N_18923,N_24139);
xor UO_1853 (O_1853,N_24969,N_23798);
or UO_1854 (O_1854,N_22228,N_24860);
and UO_1855 (O_1855,N_18849,N_23698);
and UO_1856 (O_1856,N_23053,N_19638);
or UO_1857 (O_1857,N_23145,N_22028);
and UO_1858 (O_1858,N_20097,N_19133);
and UO_1859 (O_1859,N_23195,N_24873);
xnor UO_1860 (O_1860,N_23647,N_20631);
nand UO_1861 (O_1861,N_22195,N_22744);
nor UO_1862 (O_1862,N_18872,N_18917);
xor UO_1863 (O_1863,N_22607,N_21404);
or UO_1864 (O_1864,N_18968,N_20489);
and UO_1865 (O_1865,N_22911,N_22456);
xnor UO_1866 (O_1866,N_22172,N_22765);
nand UO_1867 (O_1867,N_21193,N_19869);
xor UO_1868 (O_1868,N_19522,N_24498);
xnor UO_1869 (O_1869,N_24514,N_24756);
and UO_1870 (O_1870,N_22653,N_20120);
or UO_1871 (O_1871,N_20307,N_23722);
nor UO_1872 (O_1872,N_21308,N_21373);
nand UO_1873 (O_1873,N_24026,N_22788);
xnor UO_1874 (O_1874,N_24266,N_20650);
or UO_1875 (O_1875,N_24638,N_19141);
or UO_1876 (O_1876,N_21097,N_23226);
xnor UO_1877 (O_1877,N_22863,N_22054);
nand UO_1878 (O_1878,N_24593,N_20074);
xor UO_1879 (O_1879,N_23916,N_23600);
nor UO_1880 (O_1880,N_24254,N_24598);
nand UO_1881 (O_1881,N_20060,N_22827);
and UO_1882 (O_1882,N_22295,N_22553);
nand UO_1883 (O_1883,N_22985,N_21381);
and UO_1884 (O_1884,N_21047,N_24707);
nor UO_1885 (O_1885,N_19778,N_21405);
nor UO_1886 (O_1886,N_22023,N_23443);
nand UO_1887 (O_1887,N_20786,N_19067);
and UO_1888 (O_1888,N_22100,N_19707);
or UO_1889 (O_1889,N_23166,N_23660);
and UO_1890 (O_1890,N_23441,N_19274);
nand UO_1891 (O_1891,N_18942,N_23044);
and UO_1892 (O_1892,N_24494,N_22432);
nand UO_1893 (O_1893,N_20316,N_18892);
nor UO_1894 (O_1894,N_24983,N_21752);
nand UO_1895 (O_1895,N_19695,N_21406);
or UO_1896 (O_1896,N_22673,N_20563);
nand UO_1897 (O_1897,N_21560,N_24197);
and UO_1898 (O_1898,N_24456,N_21609);
xnor UO_1899 (O_1899,N_21845,N_24533);
nand UO_1900 (O_1900,N_21155,N_22558);
and UO_1901 (O_1901,N_19807,N_23908);
nor UO_1902 (O_1902,N_24857,N_20132);
nand UO_1903 (O_1903,N_18826,N_24173);
nor UO_1904 (O_1904,N_20301,N_23406);
nor UO_1905 (O_1905,N_22095,N_22130);
nor UO_1906 (O_1906,N_21990,N_21378);
xor UO_1907 (O_1907,N_22630,N_20515);
nand UO_1908 (O_1908,N_24500,N_21646);
nor UO_1909 (O_1909,N_24643,N_20499);
or UO_1910 (O_1910,N_24553,N_24640);
or UO_1911 (O_1911,N_20524,N_21940);
nand UO_1912 (O_1912,N_19667,N_24182);
nor UO_1913 (O_1913,N_20884,N_24881);
nand UO_1914 (O_1914,N_21618,N_19138);
and UO_1915 (O_1915,N_21632,N_24610);
or UO_1916 (O_1916,N_23956,N_22825);
nor UO_1917 (O_1917,N_22115,N_22011);
or UO_1918 (O_1918,N_23193,N_22378);
or UO_1919 (O_1919,N_24299,N_21728);
or UO_1920 (O_1920,N_24296,N_20095);
and UO_1921 (O_1921,N_19423,N_22671);
nand UO_1922 (O_1922,N_24022,N_24092);
xnor UO_1923 (O_1923,N_21043,N_21796);
and UO_1924 (O_1924,N_22151,N_20188);
nor UO_1925 (O_1925,N_18787,N_23409);
nand UO_1926 (O_1926,N_19175,N_20430);
xor UO_1927 (O_1927,N_23581,N_24623);
nor UO_1928 (O_1928,N_23814,N_20964);
or UO_1929 (O_1929,N_24519,N_20977);
nand UO_1930 (O_1930,N_20417,N_24959);
or UO_1931 (O_1931,N_18783,N_20393);
nor UO_1932 (O_1932,N_23252,N_24067);
nand UO_1933 (O_1933,N_20592,N_21868);
and UO_1934 (O_1934,N_20377,N_20171);
nand UO_1935 (O_1935,N_19339,N_24875);
and UO_1936 (O_1936,N_22494,N_24479);
or UO_1937 (O_1937,N_24012,N_22092);
nand UO_1938 (O_1938,N_21567,N_19616);
xor UO_1939 (O_1939,N_21653,N_19903);
nand UO_1940 (O_1940,N_23157,N_22131);
nor UO_1941 (O_1941,N_22084,N_18959);
or UO_1942 (O_1942,N_21571,N_19036);
nand UO_1943 (O_1943,N_20172,N_23179);
nand UO_1944 (O_1944,N_21531,N_24329);
or UO_1945 (O_1945,N_21202,N_19025);
nor UO_1946 (O_1946,N_21005,N_19132);
nand UO_1947 (O_1947,N_21168,N_20760);
nor UO_1948 (O_1948,N_20264,N_24801);
nand UO_1949 (O_1949,N_19884,N_18998);
and UO_1950 (O_1950,N_23631,N_23996);
or UO_1951 (O_1951,N_24465,N_19250);
nand UO_1952 (O_1952,N_19172,N_19892);
xor UO_1953 (O_1953,N_20261,N_18778);
xnor UO_1954 (O_1954,N_21511,N_20969);
nand UO_1955 (O_1955,N_24620,N_23656);
and UO_1956 (O_1956,N_22132,N_24730);
and UO_1957 (O_1957,N_21696,N_21535);
and UO_1958 (O_1958,N_24837,N_19953);
or UO_1959 (O_1959,N_19271,N_24251);
nand UO_1960 (O_1960,N_21892,N_20869);
xor UO_1961 (O_1961,N_21544,N_22594);
xor UO_1962 (O_1962,N_23868,N_23880);
xnor UO_1963 (O_1963,N_23255,N_21217);
xnor UO_1964 (O_1964,N_23766,N_22476);
xnor UO_1965 (O_1965,N_19795,N_23628);
nor UO_1966 (O_1966,N_20210,N_24844);
xnor UO_1967 (O_1967,N_18961,N_24258);
nand UO_1968 (O_1968,N_24942,N_23464);
xor UO_1969 (O_1969,N_22649,N_23235);
or UO_1970 (O_1970,N_23641,N_19699);
nand UO_1971 (O_1971,N_22313,N_22967);
nor UO_1972 (O_1972,N_23012,N_22556);
or UO_1973 (O_1973,N_20054,N_24203);
nand UO_1974 (O_1974,N_24484,N_21674);
xnor UO_1975 (O_1975,N_21988,N_19765);
and UO_1976 (O_1976,N_20250,N_22532);
nand UO_1977 (O_1977,N_21029,N_24662);
and UO_1978 (O_1978,N_20810,N_23034);
nand UO_1979 (O_1979,N_24276,N_19283);
or UO_1980 (O_1980,N_19184,N_21861);
xor UO_1981 (O_1981,N_21682,N_21027);
nand UO_1982 (O_1982,N_18904,N_23397);
nand UO_1983 (O_1983,N_22264,N_21359);
or UO_1984 (O_1984,N_23850,N_19787);
or UO_1985 (O_1985,N_23821,N_22625);
or UO_1986 (O_1986,N_20619,N_24762);
nor UO_1987 (O_1987,N_19786,N_19852);
or UO_1988 (O_1988,N_19142,N_20006);
nor UO_1989 (O_1989,N_23854,N_20370);
nand UO_1990 (O_1990,N_22757,N_18779);
and UO_1991 (O_1991,N_20677,N_22900);
xor UO_1992 (O_1992,N_20348,N_19433);
nor UO_1993 (O_1993,N_21733,N_19201);
or UO_1994 (O_1994,N_19092,N_23661);
nand UO_1995 (O_1995,N_24785,N_21150);
or UO_1996 (O_1996,N_19691,N_18936);
nand UO_1997 (O_1997,N_19515,N_24355);
nand UO_1998 (O_1998,N_21426,N_22419);
nor UO_1999 (O_1999,N_20929,N_21285);
and UO_2000 (O_2000,N_23999,N_19741);
nor UO_2001 (O_2001,N_21272,N_23093);
or UO_2002 (O_2002,N_20519,N_20287);
or UO_2003 (O_2003,N_19017,N_22973);
xor UO_2004 (O_2004,N_22803,N_23974);
nor UO_2005 (O_2005,N_19684,N_23449);
and UO_2006 (O_2006,N_21578,N_20104);
nand UO_2007 (O_2007,N_23373,N_23420);
and UO_2008 (O_2008,N_24065,N_21534);
nor UO_2009 (O_2009,N_24078,N_23057);
nand UO_2010 (O_2010,N_22780,N_20579);
nor UO_2011 (O_2011,N_20622,N_19301);
or UO_2012 (O_2012,N_21394,N_20853);
and UO_2013 (O_2013,N_23873,N_21021);
and UO_2014 (O_2014,N_22791,N_24073);
xnor UO_2015 (O_2015,N_24241,N_24160);
and UO_2016 (O_2016,N_22279,N_24477);
xor UO_2017 (O_2017,N_21930,N_23303);
and UO_2018 (O_2018,N_20509,N_22853);
nand UO_2019 (O_2019,N_24815,N_18863);
nand UO_2020 (O_2020,N_20875,N_24239);
nand UO_2021 (O_2021,N_23161,N_21724);
and UO_2022 (O_2022,N_20241,N_21968);
or UO_2023 (O_2023,N_18805,N_19302);
nor UO_2024 (O_2024,N_22726,N_22652);
and UO_2025 (O_2025,N_20013,N_21882);
nand UO_2026 (O_2026,N_22508,N_23585);
or UO_2027 (O_2027,N_24774,N_20882);
and UO_2028 (O_2028,N_22648,N_19518);
xor UO_2029 (O_2029,N_24761,N_24527);
and UO_2030 (O_2030,N_19867,N_21778);
nor UO_2031 (O_2031,N_21973,N_23119);
and UO_2032 (O_2032,N_20294,N_20860);
nand UO_2033 (O_2033,N_19070,N_24665);
or UO_2034 (O_2034,N_19894,N_19321);
nand UO_2035 (O_2035,N_24589,N_24933);
and UO_2036 (O_2036,N_24579,N_22903);
nand UO_2037 (O_2037,N_19794,N_24839);
nand UO_2038 (O_2038,N_21357,N_23852);
nand UO_2039 (O_2039,N_19593,N_24619);
nor UO_2040 (O_2040,N_19512,N_23788);
and UO_2041 (O_2041,N_20685,N_23036);
xnor UO_2042 (O_2042,N_20675,N_24275);
and UO_2043 (O_2043,N_21034,N_19633);
and UO_2044 (O_2044,N_21838,N_19084);
nand UO_2045 (O_2045,N_24314,N_23299);
nand UO_2046 (O_2046,N_23553,N_22346);
nor UO_2047 (O_2047,N_22724,N_24313);
and UO_2048 (O_2048,N_22422,N_24932);
xor UO_2049 (O_2049,N_20248,N_22119);
and UO_2050 (O_2050,N_20831,N_21727);
nor UO_2051 (O_2051,N_22338,N_23810);
or UO_2052 (O_2052,N_21995,N_24826);
nor UO_2053 (O_2053,N_18905,N_24703);
nor UO_2054 (O_2054,N_21088,N_24789);
xnor UO_2055 (O_2055,N_23395,N_21767);
and UO_2056 (O_2056,N_20893,N_21437);
and UO_2057 (O_2057,N_18949,N_20737);
or UO_2058 (O_2058,N_19541,N_23244);
and UO_2059 (O_2059,N_22239,N_23619);
xor UO_2060 (O_2060,N_19970,N_20986);
nand UO_2061 (O_2061,N_20529,N_23142);
nand UO_2062 (O_2062,N_20551,N_22006);
or UO_2063 (O_2063,N_19183,N_22481);
and UO_2064 (O_2064,N_20724,N_20465);
and UO_2065 (O_2065,N_24668,N_23378);
or UO_2066 (O_2066,N_21208,N_22327);
nand UO_2067 (O_2067,N_23268,N_19560);
xor UO_2068 (O_2068,N_24919,N_23075);
and UO_2069 (O_2069,N_24664,N_19746);
xor UO_2070 (O_2070,N_22153,N_21617);
nor UO_2071 (O_2071,N_24267,N_20582);
nand UO_2072 (O_2072,N_24650,N_18801);
and UO_2073 (O_2073,N_22199,N_19613);
or UO_2074 (O_2074,N_19310,N_24096);
xor UO_2075 (O_2075,N_20395,N_22614);
or UO_2076 (O_2076,N_19061,N_22000);
nor UO_2077 (O_2077,N_22560,N_22715);
and UO_2078 (O_2078,N_18885,N_23708);
xnor UO_2079 (O_2079,N_19382,N_24632);
nand UO_2080 (O_2080,N_23851,N_20391);
nor UO_2081 (O_2081,N_21067,N_20403);
and UO_2082 (O_2082,N_20366,N_20872);
nand UO_2083 (O_2083,N_24427,N_21390);
and UO_2084 (O_2084,N_22102,N_24777);
xnor UO_2085 (O_2085,N_20924,N_23644);
nand UO_2086 (O_2086,N_19650,N_18962);
and UO_2087 (O_2087,N_23767,N_24264);
nand UO_2088 (O_2088,N_22232,N_22546);
and UO_2089 (O_2089,N_20735,N_22472);
and UO_2090 (O_2090,N_23719,N_19817);
and UO_2091 (O_2091,N_21594,N_21073);
xor UO_2092 (O_2092,N_21371,N_20707);
nor UO_2093 (O_2093,N_23727,N_23926);
and UO_2094 (O_2094,N_20522,N_24670);
or UO_2095 (O_2095,N_22434,N_19950);
nand UO_2096 (O_2096,N_21498,N_23301);
nand UO_2097 (O_2097,N_23808,N_20576);
or UO_2098 (O_2098,N_20341,N_19600);
or UO_2099 (O_2099,N_23258,N_20179);
and UO_2100 (O_2100,N_24912,N_22505);
xor UO_2101 (O_2101,N_21261,N_24530);
and UO_2102 (O_2102,N_21918,N_21237);
nor UO_2103 (O_2103,N_19783,N_24578);
and UO_2104 (O_2104,N_23490,N_19553);
and UO_2105 (O_2105,N_19501,N_22695);
or UO_2106 (O_2106,N_20792,N_21259);
nand UO_2107 (O_2107,N_20535,N_22871);
or UO_2108 (O_2108,N_23320,N_21592);
nor UO_2109 (O_2109,N_23480,N_23615);
xor UO_2110 (O_2110,N_24030,N_23827);
nand UO_2111 (O_2111,N_22457,N_22767);
or UO_2112 (O_2112,N_19181,N_22590);
nand UO_2113 (O_2113,N_19551,N_20135);
or UO_2114 (O_2114,N_19073,N_20733);
or UO_2115 (O_2115,N_22047,N_24279);
or UO_2116 (O_2116,N_19860,N_22946);
nand UO_2117 (O_2117,N_19700,N_23487);
nor UO_2118 (O_2118,N_19464,N_21485);
nand UO_2119 (O_2119,N_23768,N_22772);
nor UO_2120 (O_2120,N_21032,N_22814);
and UO_2121 (O_2121,N_19177,N_18821);
xnor UO_2122 (O_2122,N_19583,N_21192);
or UO_2123 (O_2123,N_21726,N_23136);
nand UO_2124 (O_2124,N_19180,N_21353);
nor UO_2125 (O_2125,N_24038,N_19912);
nand UO_2126 (O_2126,N_21846,N_21807);
nor UO_2127 (O_2127,N_20988,N_21340);
or UO_2128 (O_2128,N_24210,N_24149);
xnor UO_2129 (O_2129,N_24603,N_19731);
nor UO_2130 (O_2130,N_20070,N_24104);
nor UO_2131 (O_2131,N_22761,N_23584);
or UO_2132 (O_2132,N_21938,N_20202);
nor UO_2133 (O_2133,N_20084,N_23640);
xor UO_2134 (O_2134,N_19269,N_20945);
or UO_2135 (O_2135,N_22812,N_24492);
nor UO_2136 (O_2136,N_23478,N_20309);
and UO_2137 (O_2137,N_21052,N_18824);
nand UO_2138 (O_2138,N_24245,N_19659);
nor UO_2139 (O_2139,N_19039,N_18980);
xor UO_2140 (O_2140,N_22676,N_19503);
nand UO_2141 (O_2141,N_18927,N_19103);
xnor UO_2142 (O_2142,N_23186,N_19121);
or UO_2143 (O_2143,N_19209,N_24419);
xor UO_2144 (O_2144,N_22575,N_19946);
and UO_2145 (O_2145,N_19340,N_21625);
or UO_2146 (O_2146,N_22025,N_20180);
nor UO_2147 (O_2147,N_24378,N_21448);
xor UO_2148 (O_2148,N_21488,N_19409);
xor UO_2149 (O_2149,N_24690,N_23513);
or UO_2150 (O_2150,N_19236,N_21655);
and UO_2151 (O_2151,N_21330,N_18808);
xor UO_2152 (O_2152,N_21254,N_20390);
xnor UO_2153 (O_2153,N_19725,N_22970);
or UO_2154 (O_2154,N_22948,N_21140);
nor UO_2155 (O_2155,N_20868,N_21093);
xor UO_2156 (O_2156,N_19242,N_24202);
nand UO_2157 (O_2157,N_18798,N_21685);
nand UO_2158 (O_2158,N_21928,N_24352);
and UO_2159 (O_2159,N_20221,N_22822);
nor UO_2160 (O_2160,N_20067,N_19332);
and UO_2161 (O_2161,N_20018,N_24991);
nor UO_2162 (O_2162,N_23063,N_19995);
and UO_2163 (O_2163,N_24792,N_21231);
xnor UO_2164 (O_2164,N_22819,N_22043);
nor UO_2165 (O_2165,N_21711,N_21660);
xor UO_2166 (O_2166,N_20277,N_19422);
nand UO_2167 (O_2167,N_21076,N_23066);
xor UO_2168 (O_2168,N_19059,N_24567);
or UO_2169 (O_2169,N_21764,N_19857);
xor UO_2170 (O_2170,N_19104,N_20974);
nor UO_2171 (O_2171,N_24018,N_24694);
or UO_2172 (O_2172,N_24002,N_24772);
or UO_2173 (O_2173,N_19758,N_23415);
and UO_2174 (O_2174,N_24390,N_21899);
and UO_2175 (O_2175,N_24192,N_22333);
and UO_2176 (O_2176,N_24537,N_19286);
nor UO_2177 (O_2177,N_23368,N_22069);
or UO_2178 (O_2178,N_24396,N_24721);
nor UO_2179 (O_2179,N_20159,N_20645);
nand UO_2180 (O_2180,N_24365,N_19485);
xor UO_2181 (O_2181,N_21789,N_21400);
nand UO_2182 (O_2182,N_22591,N_24566);
nor UO_2183 (O_2183,N_19223,N_19402);
nor UO_2184 (O_2184,N_19312,N_21207);
and UO_2185 (O_2185,N_22661,N_19131);
and UO_2186 (O_2186,N_21697,N_20161);
or UO_2187 (O_2187,N_21862,N_22688);
nand UO_2188 (O_2188,N_20372,N_21937);
and UO_2189 (O_2189,N_20406,N_24684);
nor UO_2190 (O_2190,N_23637,N_23196);
and UO_2191 (O_2191,N_20993,N_20697);
nor UO_2192 (O_2192,N_23204,N_20777);
nand UO_2193 (O_2193,N_20722,N_23321);
nor UO_2194 (O_2194,N_22833,N_21619);
xor UO_2195 (O_2195,N_18764,N_20437);
nand UO_2196 (O_2196,N_24893,N_21750);
nand UO_2197 (O_2197,N_21172,N_21895);
and UO_2198 (O_2198,N_19771,N_22763);
nor UO_2199 (O_2199,N_20581,N_20164);
nor UO_2200 (O_2200,N_20870,N_23569);
nand UO_2201 (O_2201,N_19591,N_19232);
and UO_2202 (O_2202,N_19931,N_22538);
or UO_2203 (O_2203,N_23857,N_23789);
or UO_2204 (O_2204,N_22891,N_22858);
or UO_2205 (O_2205,N_21398,N_24336);
or UO_2206 (O_2206,N_24273,N_19216);
and UO_2207 (O_2207,N_20476,N_22752);
and UO_2208 (O_2208,N_24094,N_20303);
and UO_2209 (O_2209,N_23755,N_20181);
or UO_2210 (O_2210,N_22461,N_18952);
or UO_2211 (O_2211,N_22489,N_20878);
nand UO_2212 (O_2212,N_23329,N_24421);
nand UO_2213 (O_2213,N_23214,N_22160);
and UO_2214 (O_2214,N_21669,N_19521);
and UO_2215 (O_2215,N_20337,N_20827);
nor UO_2216 (O_2216,N_19159,N_22068);
xor UO_2217 (O_2217,N_21451,N_20943);
or UO_2218 (O_2218,N_24611,N_22629);
xnor UO_2219 (O_2219,N_22605,N_22901);
and UO_2220 (O_2220,N_22759,N_22864);
and UO_2221 (O_2221,N_24158,N_19619);
and UO_2222 (O_2222,N_24616,N_22427);
nor UO_2223 (O_2223,N_19724,N_20680);
or UO_2224 (O_2224,N_22409,N_24767);
nor UO_2225 (O_2225,N_20507,N_23759);
or UO_2226 (O_2226,N_20912,N_22352);
or UO_2227 (O_2227,N_23526,N_24340);
xor UO_2228 (O_2228,N_20429,N_23551);
nand UO_2229 (O_2229,N_23800,N_24174);
or UO_2230 (O_2230,N_22004,N_21906);
nand UO_2231 (O_2231,N_24846,N_18984);
nor UO_2232 (O_2232,N_22711,N_19626);
nor UO_2233 (O_2233,N_24496,N_24055);
and UO_2234 (O_2234,N_22773,N_23606);
nand UO_2235 (O_2235,N_24282,N_24334);
or UO_2236 (O_2236,N_21143,N_20482);
xnor UO_2237 (O_2237,N_20189,N_19625);
nor UO_2238 (O_2238,N_20385,N_19734);
or UO_2239 (O_2239,N_21146,N_24914);
xor UO_2240 (O_2240,N_24117,N_20911);
and UO_2241 (O_2241,N_22182,N_24845);
nor UO_2242 (O_2242,N_21554,N_20987);
nor UO_2243 (O_2243,N_20014,N_19150);
or UO_2244 (O_2244,N_21550,N_19391);
xnor UO_2245 (O_2245,N_23817,N_18981);
xor UO_2246 (O_2246,N_20247,N_20788);
nand UO_2247 (O_2247,N_19526,N_20692);
nand UO_2248 (O_2248,N_20388,N_19547);
xor UO_2249 (O_2249,N_19228,N_21362);
and UO_2250 (O_2250,N_21196,N_22580);
nand UO_2251 (O_2251,N_21645,N_20007);
nand UO_2252 (O_2252,N_21212,N_24156);
or UO_2253 (O_2253,N_23876,N_19549);
xor UO_2254 (O_2254,N_21771,N_21793);
or UO_2255 (O_2255,N_19217,N_20149);
and UO_2256 (O_2256,N_21408,N_24382);
xnor UO_2257 (O_2257,N_22643,N_20415);
nand UO_2258 (O_2258,N_19827,N_19484);
and UO_2259 (O_2259,N_21050,N_20349);
nand UO_2260 (O_2260,N_24148,N_20162);
nor UO_2261 (O_2261,N_22020,N_24178);
nor UO_2262 (O_2262,N_20174,N_19900);
xnor UO_2263 (O_2263,N_22890,N_19473);
and UO_2264 (O_2264,N_24803,N_24211);
and UO_2265 (O_2265,N_22728,N_19110);
xnor UO_2266 (O_2266,N_22111,N_23575);
and UO_2267 (O_2267,N_21111,N_19760);
nor UO_2268 (O_2268,N_20113,N_24776);
and UO_2269 (O_2269,N_20453,N_19567);
or UO_2270 (O_2270,N_19278,N_23646);
or UO_2271 (O_2271,N_19773,N_19637);
or UO_2272 (O_2272,N_23909,N_20871);
xor UO_2273 (O_2273,N_23576,N_23577);
nor UO_2274 (O_2274,N_19607,N_24899);
xor UO_2275 (O_2275,N_21910,N_21608);
and UO_2276 (O_2276,N_18954,N_24080);
nand UO_2277 (O_2277,N_23137,N_22394);
nor UO_2278 (O_2278,N_21319,N_21829);
and UO_2279 (O_2279,N_22559,N_22528);
nor UO_2280 (O_2280,N_20741,N_22956);
xnor UO_2281 (O_2281,N_18756,N_23300);
nand UO_2282 (O_2282,N_24034,N_21179);
and UO_2283 (O_2283,N_19064,N_23546);
or UO_2284 (O_2284,N_21008,N_20046);
nor UO_2285 (O_2285,N_23349,N_20079);
and UO_2286 (O_2286,N_21505,N_21178);
or UO_2287 (O_2287,N_22634,N_20039);
or UO_2288 (O_2288,N_20035,N_23016);
and UO_2289 (O_2289,N_20900,N_19727);
and UO_2290 (O_2290,N_22834,N_21489);
nor UO_2291 (O_2291,N_22995,N_20718);
or UO_2292 (O_2292,N_19359,N_24560);
and UO_2293 (O_2293,N_21045,N_22950);
and UO_2294 (O_2294,N_18990,N_20245);
xor UO_2295 (O_2295,N_22541,N_22789);
or UO_2296 (O_2296,N_23198,N_22510);
xor UO_2297 (O_2297,N_23160,N_23704);
xor UO_2298 (O_2298,N_18948,N_18853);
nand UO_2299 (O_2299,N_19963,N_20271);
or UO_2300 (O_2300,N_23347,N_20996);
nand UO_2301 (O_2301,N_21379,N_20052);
nor UO_2302 (O_2302,N_21349,N_19513);
or UO_2303 (O_2303,N_21662,N_21283);
and UO_2304 (O_2304,N_23983,N_23650);
nand UO_2305 (O_2305,N_21749,N_20005);
nand UO_2306 (O_2306,N_23792,N_23621);
xor UO_2307 (O_2307,N_23820,N_21805);
xnor UO_2308 (O_2308,N_19720,N_23297);
nor UO_2309 (O_2309,N_23966,N_22107);
and UO_2310 (O_2310,N_24906,N_21189);
xor UO_2311 (O_2311,N_20490,N_22526);
nor UO_2312 (O_2312,N_21068,N_22764);
nor UO_2313 (O_2313,N_21115,N_21549);
xor UO_2314 (O_2314,N_21430,N_20378);
and UO_2315 (O_2315,N_22421,N_21971);
nand UO_2316 (O_2316,N_22413,N_19237);
and UO_2317 (O_2317,N_20994,N_20380);
xnor UO_2318 (O_2318,N_24350,N_24451);
nand UO_2319 (O_2319,N_20440,N_20600);
and UO_2320 (O_2320,N_24859,N_21523);
nor UO_2321 (O_2321,N_19668,N_21723);
nor UO_2322 (O_2322,N_18955,N_23626);
nor UO_2323 (O_2323,N_21397,N_22117);
and UO_2324 (O_2324,N_21438,N_19906);
nand UO_2325 (O_2325,N_18864,N_23342);
xor UO_2326 (O_2326,N_23267,N_23230);
xor UO_2327 (O_2327,N_22756,N_22373);
xnor UO_2328 (O_2328,N_21516,N_22865);
xnor UO_2329 (O_2329,N_20260,N_19009);
nand UO_2330 (O_2330,N_23485,N_19306);
nor UO_2331 (O_2331,N_23653,N_23248);
nand UO_2332 (O_2332,N_22838,N_20851);
nand UO_2333 (O_2333,N_21506,N_19520);
and UO_2334 (O_2334,N_18800,N_22621);
or UO_2335 (O_2335,N_19233,N_24898);
or UO_2336 (O_2336,N_23080,N_24444);
nand UO_2337 (O_2337,N_24995,N_22637);
nor UO_2338 (O_2338,N_21049,N_24118);
and UO_2339 (O_2339,N_23512,N_23785);
and UO_2340 (O_2340,N_23721,N_21028);
or UO_2341 (O_2341,N_23772,N_19710);
and UO_2342 (O_2342,N_24079,N_20369);
nand UO_2343 (O_2343,N_20332,N_20699);
or UO_2344 (O_2344,N_18750,N_24335);
xnor UO_2345 (O_2345,N_24963,N_22912);
or UO_2346 (O_2346,N_21872,N_21991);
xor UO_2347 (O_2347,N_23613,N_23364);
and UO_2348 (O_2348,N_22872,N_23355);
nand UO_2349 (O_2349,N_24821,N_23175);
or UO_2350 (O_2350,N_19845,N_21627);
or UO_2351 (O_2351,N_21744,N_24493);
nor UO_2352 (O_2352,N_20436,N_24277);
or UO_2353 (O_2353,N_22335,N_19456);
or UO_2354 (O_2354,N_20234,N_23521);
and UO_2355 (O_2355,N_21186,N_24164);
nor UO_2356 (O_2356,N_22837,N_24057);
nor UO_2357 (O_2357,N_21874,N_22032);
and UO_2358 (O_2358,N_24041,N_20383);
or UO_2359 (O_2359,N_21830,N_21393);
xnor UO_2360 (O_2360,N_23691,N_20089);
and UO_2361 (O_2361,N_19594,N_23560);
nand UO_2362 (O_2362,N_20357,N_19192);
nor UO_2363 (O_2363,N_23597,N_22018);
and UO_2364 (O_2364,N_18925,N_19357);
nor UO_2365 (O_2365,N_21137,N_19075);
xnor UO_2366 (O_2366,N_24736,N_22225);
and UO_2367 (O_2367,N_19276,N_23274);
and UO_2368 (O_2368,N_24658,N_21445);
xnor UO_2369 (O_2369,N_19258,N_20719);
and UO_2370 (O_2370,N_24804,N_24615);
and UO_2371 (O_2371,N_24642,N_18772);
nor UO_2372 (O_2372,N_21661,N_24595);
or UO_2373 (O_2373,N_23812,N_21879);
and UO_2374 (O_2374,N_19780,N_18932);
and UO_2375 (O_2375,N_19711,N_23148);
nor UO_2376 (O_2376,N_23765,N_19047);
and UO_2377 (O_2377,N_21708,N_19806);
or UO_2378 (O_2378,N_22725,N_19178);
xor UO_2379 (O_2379,N_21442,N_19981);
nor UO_2380 (O_2380,N_20891,N_24956);
nand UO_2381 (O_2381,N_19933,N_23715);
and UO_2382 (O_2382,N_22436,N_21144);
and UO_2383 (O_2383,N_23564,N_22240);
or UO_2384 (O_2384,N_22143,N_20335);
nor UO_2385 (O_2385,N_21564,N_20791);
nand UO_2386 (O_2386,N_24106,N_23029);
xor UO_2387 (O_2387,N_22395,N_22178);
nor UO_2388 (O_2388,N_24676,N_24900);
nor UO_2389 (O_2389,N_18781,N_22254);
or UO_2390 (O_2390,N_21883,N_21939);
or UO_2391 (O_2391,N_19001,N_21466);
nand UO_2392 (O_2392,N_23948,N_19754);
or UO_2393 (O_2393,N_21151,N_20363);
or UO_2394 (O_2394,N_24204,N_24798);
nand UO_2395 (O_2395,N_19371,N_24162);
and UO_2396 (O_2396,N_21904,N_19829);
and UO_2397 (O_2397,N_20282,N_24992);
and UO_2398 (O_2398,N_21339,N_24581);
nand UO_2399 (O_2399,N_19158,N_20246);
or UO_2400 (O_2400,N_22367,N_23106);
nor UO_2401 (O_2401,N_21258,N_22303);
nand UO_2402 (O_2402,N_24781,N_18910);
and UO_2403 (O_2403,N_23425,N_20594);
xor UO_2404 (O_2404,N_21876,N_21470);
nand UO_2405 (O_2405,N_22537,N_23122);
xor UO_2406 (O_2406,N_19304,N_23775);
and UO_2407 (O_2407,N_20423,N_23393);
nor UO_2408 (O_2408,N_20500,N_22272);
and UO_2409 (O_2409,N_19246,N_21165);
or UO_2410 (O_2410,N_21812,N_24917);
or UO_2411 (O_2411,N_24014,N_21367);
nand UO_2412 (O_2412,N_22746,N_19977);
nor UO_2413 (O_2413,N_22994,N_21108);
xor UO_2414 (O_2414,N_23730,N_23020);
nand UO_2415 (O_2415,N_23793,N_19843);
xnor UO_2416 (O_2416,N_20201,N_21356);
nor UO_2417 (O_2417,N_20468,N_23714);
nand UO_2418 (O_2418,N_20798,N_23038);
nor UO_2419 (O_2419,N_24937,N_18887);
nor UO_2420 (O_2420,N_19612,N_21788);
or UO_2421 (O_2421,N_23954,N_18926);
or UO_2422 (O_2422,N_20814,N_20601);
and UO_2423 (O_2423,N_22360,N_23422);
xor UO_2424 (O_2424,N_21103,N_20414);
and UO_2425 (O_2425,N_23344,N_18950);
and UO_2426 (O_2426,N_23700,N_23346);
nor UO_2427 (O_2427,N_21700,N_23671);
xnor UO_2428 (O_2428,N_20753,N_23862);
nor UO_2429 (O_2429,N_23990,N_21848);
or UO_2430 (O_2430,N_24924,N_24971);
nand UO_2431 (O_2431,N_22579,N_21300);
xor UO_2432 (O_2432,N_24977,N_23061);
nand UO_2433 (O_2433,N_24657,N_18795);
xor UO_2434 (O_2434,N_24328,N_20713);
nor UO_2435 (O_2435,N_24508,N_24895);
or UO_2436 (O_2436,N_23723,N_20082);
or UO_2437 (O_2437,N_20043,N_23310);
and UO_2438 (O_2438,N_20313,N_20812);
or UO_2439 (O_2439,N_19277,N_24322);
or UO_2440 (O_2440,N_23247,N_19194);
nand UO_2441 (O_2441,N_20618,N_22357);
nand UO_2442 (O_2442,N_22440,N_24075);
nand UO_2443 (O_2443,N_22584,N_23125);
nand UO_2444 (O_2444,N_19401,N_22754);
and UO_2445 (O_2445,N_20027,N_20768);
and UO_2446 (O_2446,N_24528,N_21248);
and UO_2447 (O_2447,N_23447,N_19125);
nand UO_2448 (O_2448,N_20259,N_20139);
xor UO_2449 (O_2449,N_19030,N_22952);
nor UO_2450 (O_2450,N_22324,N_21779);
nor UO_2451 (O_2451,N_19782,N_23341);
xnor UO_2452 (O_2452,N_22180,N_20360);
xor UO_2453 (O_2453,N_19208,N_23233);
nand UO_2454 (O_2454,N_22039,N_19151);
nand UO_2455 (O_2455,N_23964,N_20528);
and UO_2456 (O_2456,N_21443,N_20150);
and UO_2457 (O_2457,N_19338,N_23337);
nor UO_2458 (O_2458,N_21589,N_22721);
or UO_2459 (O_2459,N_18850,N_24353);
and UO_2460 (O_2460,N_21507,N_22701);
xor UO_2461 (O_2461,N_21577,N_23902);
xnor UO_2462 (O_2462,N_20361,N_24999);
and UO_2463 (O_2463,N_23108,N_24386);
xor UO_2464 (O_2464,N_20610,N_19080);
nor UO_2465 (O_2465,N_22636,N_23903);
nor UO_2466 (O_2466,N_19730,N_20747);
xor UO_2467 (O_2467,N_22988,N_23334);
xnor UO_2468 (O_2468,N_24007,N_22426);
xor UO_2469 (O_2469,N_24751,N_22738);
nor UO_2470 (O_2470,N_23907,N_20475);
xor UO_2471 (O_2471,N_20105,N_21999);
xor UO_2472 (O_2472,N_22500,N_22874);
xnor UO_2473 (O_2473,N_19272,N_19871);
xnor UO_2474 (O_2474,N_23141,N_20047);
xnor UO_2475 (O_2475,N_21154,N_19666);
xnor UO_2476 (O_2476,N_18846,N_20531);
and UO_2477 (O_2477,N_19245,N_18793);
nand UO_2478 (O_2478,N_21675,N_24934);
nand UO_2479 (O_2479,N_22370,N_24364);
nand UO_2480 (O_2480,N_19533,N_24412);
nor UO_2481 (O_2481,N_19548,N_24218);
nor UO_2482 (O_2482,N_20312,N_22581);
xor UO_2483 (O_2483,N_22205,N_22706);
nor UO_2484 (O_2484,N_24877,N_22491);
or UO_2485 (O_2485,N_20276,N_23188);
xnor UO_2486 (O_2486,N_21117,N_24693);
nand UO_2487 (O_2487,N_19632,N_21570);
and UO_2488 (O_2488,N_19673,N_21071);
nand UO_2489 (O_2489,N_23872,N_19205);
nand UO_2490 (O_2490,N_21368,N_24863);
nand UO_2491 (O_2491,N_23501,N_23943);
nor UO_2492 (O_2492,N_19379,N_22796);
or UO_2493 (O_2493,N_23511,N_22969);
xor UO_2494 (O_2494,N_22247,N_19564);
xnor UO_2495 (O_2495,N_23979,N_19010);
nand UO_2496 (O_2496,N_19078,N_21306);
or UO_2497 (O_2497,N_24278,N_24132);
nor UO_2498 (O_2498,N_22656,N_22949);
xnor UO_2499 (O_2499,N_22750,N_24351);
and UO_2500 (O_2500,N_22555,N_24209);
xor UO_2501 (O_2501,N_19038,N_18816);
nor UO_2502 (O_2502,N_23809,N_21797);
xnor UO_2503 (O_2503,N_20416,N_19330);
xor UO_2504 (O_2504,N_22587,N_21841);
nand UO_2505 (O_2505,N_24705,N_21054);
nand UO_2506 (O_2506,N_19952,N_20800);
and UO_2507 (O_2507,N_20106,N_21515);
xnor UO_2508 (O_2508,N_20136,N_21064);
xor UO_2509 (O_2509,N_19588,N_21173);
nor UO_2510 (O_2510,N_19956,N_20268);
nor UO_2511 (O_2511,N_20497,N_22739);
xnor UO_2512 (O_2512,N_21602,N_21436);
nand UO_2513 (O_2513,N_20928,N_21479);
xnor UO_2514 (O_2514,N_19425,N_23757);
and UO_2515 (O_2515,N_20220,N_19032);
or UO_2516 (O_2516,N_23411,N_23813);
and UO_2517 (O_2517,N_21224,N_20087);
xnor UO_2518 (O_2518,N_23408,N_23622);
xnor UO_2519 (O_2519,N_20858,N_23059);
nand UO_2520 (O_2520,N_19441,N_21923);
and UO_2521 (O_2521,N_21257,N_21775);
xor UO_2522 (O_2522,N_19563,N_20041);
or UO_2523 (O_2523,N_21920,N_19000);
nor UO_2524 (O_2524,N_22187,N_21680);
nand UO_2525 (O_2525,N_23365,N_23019);
nand UO_2526 (O_2526,N_20222,N_20655);
xor UO_2527 (O_2527,N_20950,N_20589);
or UO_2528 (O_2528,N_22749,N_22698);
and UO_2529 (O_2529,N_20094,N_21085);
nand UO_2530 (O_2530,N_23302,N_24268);
or UO_2531 (O_2531,N_22939,N_24495);
and UO_2532 (O_2532,N_23111,N_21223);
or UO_2533 (O_2533,N_19432,N_24542);
and UO_2534 (O_2534,N_21709,N_23253);
xnor UO_2535 (O_2535,N_19671,N_20333);
xnor UO_2536 (O_2536,N_19643,N_19106);
or UO_2537 (O_2537,N_19241,N_22793);
nand UO_2538 (O_2538,N_23593,N_19155);
xnor UO_2539 (O_2539,N_20053,N_23078);
nor UO_2540 (O_2540,N_20797,N_19935);
xor UO_2541 (O_2541,N_20051,N_18757);
or UO_2542 (O_2542,N_24515,N_23164);
and UO_2543 (O_2543,N_18867,N_19169);
or UO_2544 (O_2544,N_20856,N_20833);
xor UO_2545 (O_2545,N_20755,N_24469);
nand UO_2546 (O_2546,N_19168,N_19870);
nand UO_2547 (O_2547,N_23607,N_24654);
nand UO_2548 (O_2548,N_19998,N_21302);
nand UO_2549 (O_2549,N_19751,N_19416);
nand UO_2550 (O_2550,N_23001,N_24271);
or UO_2551 (O_2551,N_21372,N_21611);
and UO_2552 (O_2552,N_19815,N_19189);
xor UO_2553 (O_2553,N_21026,N_21652);
and UO_2554 (O_2554,N_24031,N_23350);
and UO_2555 (O_2555,N_24506,N_22828);
xor UO_2556 (O_2556,N_24547,N_20691);
or UO_2557 (O_2557,N_19027,N_22317);
or UO_2558 (O_2558,N_22691,N_21781);
nand UO_2559 (O_2559,N_20025,N_24794);
nor UO_2560 (O_2560,N_22867,N_18759);
and UO_2561 (O_2561,N_21810,N_21561);
nor UO_2562 (O_2562,N_19322,N_19752);
and UO_2563 (O_2563,N_20314,N_23084);
nor UO_2564 (O_2564,N_24757,N_24910);
nand UO_2565 (O_2565,N_20587,N_22400);
and UO_2566 (O_2566,N_23735,N_22410);
and UO_2567 (O_2567,N_24790,N_23325);
nand UO_2568 (O_2568,N_21759,N_20290);
xor UO_2569 (O_2569,N_24962,N_19098);
xor UO_2570 (O_2570,N_24984,N_19824);
nand UO_2571 (O_2571,N_22551,N_23538);
or UO_2572 (O_2572,N_20099,N_20322);
xor UO_2573 (O_2573,N_24011,N_24672);
nor UO_2574 (O_2574,N_20678,N_24759);
and UO_2575 (O_2575,N_23710,N_23743);
and UO_2576 (O_2576,N_19362,N_19265);
xor UO_2577 (O_2577,N_21585,N_18753);
and UO_2578 (O_2578,N_22961,N_19676);
and UO_2579 (O_2579,N_18970,N_23537);
nand UO_2580 (O_2580,N_23552,N_20613);
and UO_2581 (O_2581,N_20036,N_23442);
and UO_2582 (O_2582,N_20387,N_24853);
or UO_2583 (O_2583,N_24089,N_19530);
nor UO_2584 (O_2584,N_21022,N_22687);
and UO_2585 (O_2585,N_21719,N_21769);
xnor UO_2586 (O_2586,N_21092,N_23392);
nor UO_2587 (O_2587,N_21656,N_18971);
and UO_2588 (O_2588,N_20389,N_18767);
and UO_2589 (O_2589,N_20124,N_23101);
and UO_2590 (O_2590,N_20807,N_23261);
and UO_2591 (O_2591,N_20975,N_21854);
xnor UO_2592 (O_2592,N_22924,N_22884);
nand UO_2593 (O_2593,N_20639,N_24389);
and UO_2594 (O_2594,N_22571,N_19535);
nand UO_2595 (O_2595,N_20828,N_22734);
and UO_2596 (O_2596,N_20861,N_18920);
and UO_2597 (O_2597,N_22971,N_20580);
nor UO_2598 (O_2598,N_24193,N_24123);
or UO_2599 (O_2599,N_19016,N_23717);
nand UO_2600 (O_2600,N_22907,N_19545);
and UO_2601 (O_2601,N_23991,N_19606);
and UO_2602 (O_2602,N_24965,N_22898);
xor UO_2603 (O_2603,N_23322,N_23716);
or UO_2604 (O_2604,N_19471,N_23484);
and UO_2605 (O_2605,N_23064,N_19452);
nor UO_2606 (O_2606,N_20983,N_20630);
or UO_2607 (O_2607,N_19876,N_20825);
or UO_2608 (O_2608,N_20487,N_22727);
nor UO_2609 (O_2609,N_21129,N_22585);
xor UO_2610 (O_2610,N_22940,N_21102);
and UO_2611 (O_2611,N_19672,N_19823);
nand UO_2612 (O_2612,N_22492,N_21522);
and UO_2613 (O_2613,N_20954,N_22376);
nand UO_2614 (O_2614,N_22059,N_24691);
or UO_2615 (O_2615,N_19658,N_23315);
or UO_2616 (O_2616,N_22463,N_21623);
nor UO_2617 (O_2617,N_21007,N_24262);
nor UO_2618 (O_2618,N_22938,N_18877);
and UO_2619 (O_2619,N_21063,N_23319);
xnor UO_2620 (O_2620,N_23205,N_21249);
nor UO_2621 (O_2621,N_22418,N_19777);
nor UO_2622 (O_2622,N_24217,N_22794);
nor UO_2623 (O_2623,N_20666,N_22485);
nand UO_2624 (O_2624,N_18857,N_19193);
or UO_2625 (O_2625,N_22015,N_23883);
nor UO_2626 (O_2626,N_22060,N_21331);
nand UO_2627 (O_2627,N_23165,N_24622);
and UO_2628 (O_2628,N_21743,N_20809);
and UO_2629 (O_2629,N_24058,N_20638);
xor UO_2630 (O_2630,N_18891,N_22635);
xnor UO_2631 (O_2631,N_19118,N_23438);
and UO_2632 (O_2632,N_23801,N_19290);
and UO_2633 (O_2633,N_24168,N_20899);
nand UO_2634 (O_2634,N_24591,N_19575);
and UO_2635 (O_2635,N_19726,N_24918);
xnor UO_2636 (O_2636,N_24083,N_22194);
nor UO_2637 (O_2637,N_20883,N_24379);
xnor UO_2638 (O_2638,N_24673,N_19344);
and UO_2639 (O_2639,N_24431,N_20167);
xnor UO_2640 (O_2640,N_24407,N_20684);
or UO_2641 (O_2641,N_19167,N_24438);
nor UO_2642 (O_2642,N_22347,N_22223);
and UO_2643 (O_2643,N_24216,N_19943);
nand UO_2644 (O_2644,N_24071,N_22128);
nor UO_2645 (O_2645,N_20111,N_22730);
nor UO_2646 (O_2646,N_24951,N_20657);
and UO_2647 (O_2647,N_23311,N_19994);
and UO_2648 (O_2648,N_24505,N_19421);
nor UO_2649 (O_2649,N_23586,N_21295);
nand UO_2650 (O_2650,N_22008,N_19571);
nor UO_2651 (O_2651,N_20555,N_20813);
and UO_2652 (O_2652,N_21596,N_22188);
or UO_2653 (O_2653,N_20128,N_23679);
or UO_2654 (O_2654,N_22078,N_24903);
xor UO_2655 (O_2655,N_24186,N_24108);
and UO_2656 (O_2656,N_19366,N_24880);
and UO_2657 (O_2657,N_24077,N_21605);
and UO_2658 (O_2658,N_19936,N_19403);
or UO_2659 (O_2659,N_22557,N_23336);
nor UO_2660 (O_2660,N_21703,N_20218);
xnor UO_2661 (O_2661,N_23967,N_22908);
nand UO_2662 (O_2662,N_22468,N_20949);
and UO_2663 (O_2663,N_23900,N_21147);
nor UO_2664 (O_2664,N_20458,N_19961);
xor UO_2665 (O_2665,N_19451,N_21292);
xor UO_2666 (O_2666,N_22266,N_24904);
nor UO_2667 (O_2667,N_19997,N_23610);
or UO_2668 (O_2668,N_22732,N_19152);
nor UO_2669 (O_2669,N_20502,N_21599);
nand UO_2670 (O_2670,N_19063,N_19043);
xnor UO_2671 (O_2671,N_21859,N_24686);
and UO_2672 (O_2672,N_19187,N_21921);
or UO_2673 (O_2673,N_19345,N_21630);
or UO_2674 (O_2674,N_20548,N_21107);
nor UO_2675 (O_2675,N_24342,N_19810);
nand UO_2676 (O_2676,N_22181,N_22572);
xor UO_2677 (O_2677,N_22380,N_22953);
nand UO_2678 (O_2678,N_24297,N_23682);
nand UO_2679 (O_2679,N_23331,N_22859);
nor UO_2680 (O_2680,N_24486,N_21215);
nand UO_2681 (O_2681,N_23690,N_21242);
nand UO_2682 (O_2682,N_19299,N_24091);
or UO_2683 (O_2683,N_18811,N_22702);
or UO_2684 (O_2684,N_20729,N_21909);
and UO_2685 (O_2685,N_24474,N_21447);
nand UO_2686 (O_2686,N_23953,N_20285);
nand UO_2687 (O_2687,N_24976,N_22330);
nor UO_2688 (O_2688,N_22493,N_24968);
or UO_2689 (O_2689,N_23940,N_21989);
nor UO_2690 (O_2690,N_19144,N_19341);
xor UO_2691 (O_2691,N_21164,N_18751);
and UO_2692 (O_2692,N_22003,N_22211);
and UO_2693 (O_2693,N_21901,N_18835);
and UO_2694 (O_2694,N_18813,N_23284);
and UO_2695 (O_2695,N_20656,N_19796);
nand UO_2696 (O_2696,N_23515,N_24865);
nand UO_2697 (O_2697,N_19145,N_23433);
nand UO_2698 (O_2698,N_20942,N_21504);
xor UO_2699 (O_2699,N_23206,N_20194);
xnor UO_2700 (O_2700,N_22755,N_20815);
or UO_2701 (O_2701,N_20351,N_22156);
and UO_2702 (O_2702,N_23887,N_19891);
and UO_2703 (O_2703,N_21569,N_23545);
and UO_2704 (O_2704,N_23306,N_21975);
xnor UO_2705 (O_2705,N_18899,N_19928);
or UO_2706 (O_2706,N_23972,N_22139);
nor UO_2707 (O_2707,N_23596,N_20863);
xor UO_2708 (O_2708,N_19759,N_23745);
nor UO_2709 (O_2709,N_21786,N_22769);
or UO_2710 (O_2710,N_21654,N_21156);
nand UO_2711 (O_2711,N_20266,N_20687);
or UO_2712 (O_2712,N_23067,N_24069);
xor UO_2713 (O_2713,N_19539,N_24729);
xnor UO_2714 (O_2714,N_23072,N_24195);
nand UO_2715 (O_2715,N_23486,N_20227);
and UO_2716 (O_2716,N_23107,N_23824);
or UO_2717 (O_2717,N_24235,N_21475);
and UO_2718 (O_2718,N_21230,N_19334);
nand UO_2719 (O_2719,N_21624,N_21392);
nand UO_2720 (O_2720,N_21246,N_21731);
nand UO_2721 (O_2721,N_23570,N_21464);
or UO_2722 (O_2722,N_24246,N_22197);
and UO_2723 (O_2723,N_19461,N_23398);
nand UO_2724 (O_2724,N_20653,N_24833);
nor UO_2725 (O_2725,N_23260,N_22718);
and UO_2726 (O_2726,N_24433,N_22777);
or UO_2727 (O_2727,N_20512,N_20424);
or UO_2728 (O_2728,N_23504,N_19176);
and UO_2729 (O_2729,N_19689,N_22569);
or UO_2730 (O_2730,N_23549,N_20364);
nand UO_2731 (O_2731,N_21907,N_20022);
and UO_2732 (O_2732,N_19866,N_24930);
nand UO_2733 (O_2733,N_24573,N_23728);
xor UO_2734 (O_2734,N_19581,N_23706);
and UO_2735 (O_2735,N_21927,N_20408);
nand UO_2736 (O_2736,N_20122,N_22899);
xnor UO_2737 (O_2737,N_24882,N_22318);
xnor UO_2738 (O_2738,N_18938,N_23847);
or UO_2739 (O_2739,N_23249,N_18929);
nor UO_2740 (O_2740,N_20756,N_21040);
nor UO_2741 (O_2741,N_23777,N_21209);
xor UO_2742 (O_2742,N_23169,N_24628);
nor UO_2743 (O_2743,N_18914,N_24155);
and UO_2744 (O_2744,N_22462,N_19399);
and UO_2745 (O_2745,N_24037,N_23889);
and UO_2746 (O_2746,N_19034,N_19095);
or UO_2747 (O_2747,N_19761,N_22167);
or UO_2748 (O_2748,N_21979,N_23688);
and UO_2749 (O_2749,N_23452,N_23997);
or UO_2750 (O_2750,N_22795,N_18782);
or UO_2751 (O_2751,N_23345,N_23236);
nand UO_2752 (O_2752,N_22762,N_24394);
xnor UO_2753 (O_2753,N_24428,N_19769);
or UO_2754 (O_2754,N_20867,N_20298);
xor UO_2755 (O_2755,N_23843,N_21636);
nor UO_2756 (O_2756,N_20123,N_19466);
or UO_2757 (O_2757,N_23097,N_24655);
or UO_2758 (O_2758,N_19601,N_22550);
nor UO_2759 (O_2759,N_19191,N_19311);
or UO_2760 (O_2760,N_21734,N_19910);
nand UO_2761 (O_2761,N_22134,N_19257);
and UO_2762 (O_2762,N_21094,N_19779);
xor UO_2763 (O_2763,N_18890,N_21965);
or UO_2764 (O_2764,N_20433,N_20561);
xnor UO_2765 (O_2765,N_20542,N_21842);
nor UO_2766 (O_2766,N_24981,N_20157);
or UO_2767 (O_2767,N_24539,N_19392);
or UO_2768 (O_2768,N_22184,N_18844);
and UO_2769 (O_2769,N_24056,N_23893);
or UO_2770 (O_2770,N_23085,N_21766);
nor UO_2771 (O_2771,N_20240,N_22122);
nor UO_2772 (O_2772,N_22990,N_22568);
nand UO_2773 (O_2773,N_23471,N_21365);
or UO_2774 (O_2774,N_24166,N_22304);
or UO_2775 (O_2775,N_22108,N_24319);
nor UO_2776 (O_2776,N_24074,N_19922);
or UO_2777 (O_2777,N_24916,N_23806);
and UO_2778 (O_2778,N_20116,N_21441);
and UO_2779 (O_2779,N_21121,N_21960);
xor UO_2780 (O_2780,N_21528,N_19978);
nand UO_2781 (O_2781,N_22089,N_21141);
nor UO_2782 (O_2782,N_19474,N_24926);
and UO_2783 (O_2783,N_21866,N_24748);
or UO_2784 (O_2784,N_20491,N_21963);
nand UO_2785 (O_2785,N_21277,N_20428);
or UO_2786 (O_2786,N_20806,N_22736);
and UO_2787 (O_2787,N_22640,N_24766);
xor UO_2788 (O_2788,N_19859,N_19825);
nor UO_2789 (O_2789,N_22145,N_20559);
and UO_2790 (O_2790,N_20029,N_18986);
xnor UO_2791 (O_2791,N_23684,N_22506);
xor UO_2792 (O_2792,N_21925,N_22287);
nand UO_2793 (O_2793,N_19285,N_21707);
xnor UO_2794 (O_2794,N_18832,N_23666);
and UO_2795 (O_2795,N_24715,N_22644);
and UO_2796 (O_2796,N_24315,N_23672);
or UO_2797 (O_2797,N_22696,N_21278);
nor UO_2798 (O_2798,N_21216,N_20080);
nand UO_2799 (O_2799,N_22238,N_21798);
and UO_2800 (O_2800,N_22753,N_22998);
or UO_2801 (O_2801,N_24717,N_20003);
xnor UO_2802 (O_2802,N_19367,N_23638);
nor UO_2803 (O_2803,N_21996,N_24141);
and UO_2804 (O_2804,N_21104,N_23534);
nand UO_2805 (O_2805,N_18983,N_24050);
xnor UO_2806 (O_2806,N_21013,N_22731);
and UO_2807 (O_2807,N_19596,N_18806);
xor UO_2808 (O_2808,N_22880,N_18859);
nor UO_2809 (O_2809,N_24181,N_21553);
nor UO_2810 (O_2810,N_21174,N_24051);
or UO_2811 (O_2811,N_23970,N_19640);
and UO_2812 (O_2812,N_22597,N_24033);
xor UO_2813 (O_2813,N_24112,N_22815);
and UO_2814 (O_2814,N_19147,N_20896);
or UO_2815 (O_2815,N_20673,N_18963);
and UO_2816 (O_2816,N_19381,N_22534);
xnor UO_2817 (O_2817,N_22164,N_19851);
nor UO_2818 (O_2818,N_24187,N_19052);
nor UO_2819 (O_2819,N_24003,N_22855);
and UO_2820 (O_2820,N_23229,N_20837);
xor UO_2821 (O_2821,N_21402,N_22453);
or UO_2822 (O_2822,N_19622,N_19308);
nor UO_2823 (O_2823,N_18916,N_23624);
nand UO_2824 (O_2824,N_22126,N_21112);
nor UO_2825 (O_2825,N_21120,N_21891);
and UO_2826 (O_2826,N_21747,N_23602);
nor UO_2827 (O_2827,N_24131,N_22617);
or UO_2828 (O_2828,N_20989,N_24746);
or UO_2829 (O_2829,N_22439,N_21380);
nor UO_2830 (O_2830,N_21559,N_20877);
or UO_2831 (O_2831,N_21869,N_20923);
xor UO_2832 (O_2832,N_21849,N_22816);
or UO_2833 (O_2833,N_23617,N_23651);
xor UO_2834 (O_2834,N_24420,N_19716);
nor UO_2835 (O_2835,N_19909,N_22088);
nand UO_2836 (O_2836,N_22019,N_20396);
xnor UO_2837 (O_2837,N_23865,N_19499);
xnor UO_2838 (O_2838,N_23121,N_21203);
xor UO_2839 (O_2839,N_22171,N_22922);
and UO_2840 (O_2840,N_24841,N_21552);
or UO_2841 (O_2841,N_24659,N_23040);
nand UO_2842 (O_2842,N_24526,N_23116);
or UO_2843 (O_2843,N_19212,N_21002);
nand UO_2844 (O_2844,N_21896,N_22044);
nor UO_2845 (O_2845,N_22300,N_24489);
nor UO_2846 (O_2846,N_20857,N_19351);
xor UO_2847 (O_2847,N_20421,N_22965);
and UO_2848 (O_2848,N_18883,N_23888);
nand UO_2849 (O_2849,N_23356,N_20668);
xnor UO_2850 (O_2850,N_20334,N_20267);
and UO_2851 (O_2851,N_20636,N_19373);
or UO_2852 (O_2852,N_19967,N_24592);
or UO_2853 (O_2853,N_19303,N_24637);
xor UO_2854 (O_2854,N_23444,N_23376);
nor UO_2855 (O_2855,N_22675,N_19376);
nand UO_2856 (O_2856,N_22663,N_20028);
xor UO_2857 (O_2857,N_20044,N_20662);
nand UO_2858 (O_2858,N_23246,N_19814);
xor UO_2859 (O_2859,N_22565,N_20698);
and UO_2860 (O_2860,N_24764,N_19490);
and UO_2861 (O_2861,N_24982,N_22677);
nand UO_2862 (O_2862,N_20787,N_24179);
nand UO_2863 (O_2863,N_24974,N_20291);
nor UO_2864 (O_2864,N_20968,N_24838);
or UO_2865 (O_2865,N_23540,N_20693);
and UO_2866 (O_2866,N_20992,N_23542);
xor UO_2867 (O_2867,N_19868,N_23837);
xor UO_2868 (O_2868,N_22154,N_22465);
and UO_2869 (O_2869,N_24936,N_21409);
and UO_2870 (O_2870,N_19117,N_24237);
or UO_2871 (O_2871,N_22682,N_19483);
xor UO_2872 (O_2872,N_23623,N_22071);
nor UO_2873 (O_2873,N_23826,N_21913);
xnor UO_2874 (O_2874,N_24570,N_18769);
and UO_2875 (O_2875,N_24450,N_18762);
xnor UO_2876 (O_2876,N_22249,N_24317);
and UO_2877 (O_2877,N_19540,N_23265);
xnor UO_2878 (O_2878,N_23525,N_23855);
xnor UO_2879 (O_2879,N_21670,N_19390);
and UO_2880 (O_2880,N_23874,N_22927);
nand UO_2881 (O_2881,N_21399,N_21383);
nor UO_2882 (O_2882,N_24532,N_24944);
xnor UO_2883 (O_2883,N_19292,N_20952);
xor UO_2884 (O_2884,N_21982,N_20556);
nor UO_2885 (O_2885,N_22717,N_19004);
xor UO_2886 (O_2886,N_24504,N_18985);
nor UO_2887 (O_2887,N_22835,N_19179);
xnor UO_2888 (O_2888,N_23550,N_23506);
and UO_2889 (O_2889,N_20927,N_21260);
nand UO_2890 (O_2890,N_24401,N_19156);
and UO_2891 (O_2891,N_24714,N_21557);
nor UO_2892 (O_2892,N_21046,N_19735);
or UO_2893 (O_2893,N_20889,N_24448);
nor UO_2894 (O_2894,N_19905,N_24100);
and UO_2895 (O_2895,N_24702,N_20493);
and UO_2896 (O_2896,N_22312,N_20843);
or UO_2897 (O_2897,N_23041,N_22703);
and UO_2898 (O_2898,N_22416,N_21563);
or UO_2899 (O_2899,N_21188,N_19481);
xor UO_2900 (O_2900,N_21547,N_24423);
or UO_2901 (O_2901,N_24385,N_20778);
xnor UO_2902 (O_2902,N_24651,N_21312);
and UO_2903 (O_2903,N_19634,N_20840);
nand UO_2904 (O_2904,N_23980,N_23069);
or UO_2905 (O_2905,N_18957,N_21699);
or UO_2906 (O_2906,N_20057,N_21042);
or UO_2907 (O_2907,N_22826,N_21159);
nand UO_2908 (O_2908,N_19083,N_19288);
xnor UO_2909 (O_2909,N_23580,N_20037);
xnor UO_2910 (O_2910,N_18889,N_19439);
nor UO_2911 (O_2911,N_19482,N_23694);
nor UO_2912 (O_2912,N_21643,N_21395);
and UO_2913 (O_2913,N_23516,N_23603);
nand UO_2914 (O_2914,N_19555,N_23831);
xnor UO_2915 (O_2915,N_21014,N_23423);
nand UO_2916 (O_2916,N_22236,N_23754);
or UO_2917 (O_2917,N_19929,N_19091);
or UO_2918 (O_2918,N_22096,N_21678);
nand UO_2919 (O_2919,N_24876,N_23018);
and UO_2920 (O_2920,N_22010,N_19284);
xor UO_2921 (O_2921,N_24574,N_23384);
nand UO_2922 (O_2922,N_20114,N_23271);
nor UO_2923 (O_2923,N_20850,N_24035);
nand UO_2924 (O_2924,N_18909,N_24674);
nor UO_2925 (O_2925,N_18840,N_19747);
or UO_2926 (O_2926,N_21568,N_23729);
xnor UO_2927 (O_2927,N_18902,N_21510);
nor UO_2928 (O_2928,N_24509,N_19788);
and UO_2929 (O_2929,N_21333,N_24653);
nor UO_2930 (O_2930,N_20997,N_21962);
or UO_2931 (O_2931,N_23931,N_23472);
or UO_2932 (O_2932,N_20226,N_19319);
or UO_2933 (O_2933,N_19327,N_22839);
or UO_2934 (O_2934,N_21389,N_23351);
nand UO_2935 (O_2935,N_22516,N_23237);
nand UO_2936 (O_2936,N_19363,N_22930);
nor UO_2937 (O_2937,N_22602,N_19863);
and UO_2938 (O_2938,N_22992,N_20537);
xnor UO_2939 (O_2939,N_24629,N_20145);
and UO_2940 (O_2940,N_19076,N_24634);
nand UO_2941 (O_2941,N_21543,N_24954);
and UO_2942 (O_2942,N_23008,N_22392);
nor UO_2943 (O_2943,N_24554,N_23799);
xor UO_2944 (O_2944,N_19057,N_20198);
and UO_2945 (O_2945,N_21469,N_24025);
nand UO_2946 (O_2946,N_24612,N_22866);
nor UO_2947 (O_2947,N_23030,N_24359);
nand UO_2948 (O_2948,N_19737,N_20473);
nand UO_2949 (O_2949,N_21870,N_23374);
and UO_2950 (O_2950,N_23895,N_23860);
nor UO_2951 (O_2951,N_20679,N_23005);
xor UO_2952 (O_2952,N_24990,N_21604);
or UO_2953 (O_2953,N_24206,N_20862);
nor UO_2954 (O_2954,N_21777,N_21885);
or UO_2955 (O_2955,N_20670,N_21473);
nand UO_2956 (O_2956,N_20085,N_24631);
nand UO_2957 (O_2957,N_19350,N_23139);
nor UO_2958 (O_2958,N_20616,N_21060);
or UO_2959 (O_2959,N_21336,N_24563);
or UO_2960 (O_2960,N_19733,N_19604);
nor UO_2961 (O_2961,N_23203,N_20001);
nand UO_2962 (O_2962,N_24808,N_21422);
nand UO_2963 (O_2963,N_24697,N_23508);
nor UO_2964 (O_2964,N_23147,N_22622);
or UO_2965 (O_2965,N_23042,N_22241);
or UO_2966 (O_2966,N_21931,N_22490);
or UO_2967 (O_2967,N_18878,N_22860);
nand UO_2968 (O_2968,N_19610,N_19360);
or UO_2969 (O_2969,N_19219,N_23245);
and UO_2970 (O_2970,N_24626,N_23556);
xnor UO_2971 (O_2971,N_22024,N_24551);
and UO_2972 (O_2972,N_22425,N_24740);
xor UO_2973 (O_2973,N_23046,N_19949);
xor UO_2974 (O_2974,N_19307,N_21476);
and UO_2975 (O_2975,N_23541,N_22229);
xor UO_2976 (O_2976,N_20710,N_22977);
and UO_2977 (O_2977,N_23156,N_22947);
nor UO_2978 (O_2978,N_21912,N_22713);
and UO_2979 (O_2979,N_24159,N_24744);
and UO_2980 (O_2980,N_22005,N_23098);
nand UO_2981 (O_2981,N_19200,N_20464);
xor UO_2982 (O_2982,N_23949,N_19458);
and UO_2983 (O_2983,N_19190,N_22680);
and UO_2984 (O_2984,N_22800,N_21575);
or UO_2985 (O_2985,N_18975,N_23177);
and UO_2986 (O_2986,N_19105,N_20887);
or UO_2987 (O_2987,N_24404,N_22902);
nor UO_2988 (O_2988,N_22846,N_24842);
xor UO_2989 (O_2989,N_24475,N_20471);
or UO_2990 (O_2990,N_18752,N_19757);
xnor UO_2991 (O_2991,N_23475,N_23383);
xnor UO_2992 (O_2992,N_22301,N_19370);
or UO_2993 (O_2993,N_22103,N_20504);
nor UO_2994 (O_2994,N_19680,N_24369);
xnor UO_2995 (O_2995,N_21403,N_20716);
nand UO_2996 (O_2996,N_22356,N_20782);
and UO_2997 (O_2997,N_20821,N_24810);
or UO_2998 (O_2998,N_22064,N_19342);
nand UO_2999 (O_2999,N_19412,N_19282);
endmodule