module basic_1500_15000_2000_10_levels_1xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
nor U0 (N_0,In_370,In_16);
nor U1 (N_1,In_215,In_1135);
and U2 (N_2,In_188,In_106);
or U3 (N_3,In_194,In_250);
and U4 (N_4,In_805,In_1121);
or U5 (N_5,In_1114,In_131);
and U6 (N_6,In_921,In_1013);
and U7 (N_7,In_1085,In_1434);
nand U8 (N_8,In_1494,In_950);
or U9 (N_9,In_368,In_135);
nor U10 (N_10,In_967,In_1314);
or U11 (N_11,In_915,In_1134);
nor U12 (N_12,In_1398,In_560);
nand U13 (N_13,In_1413,In_882);
and U14 (N_14,In_886,In_1111);
and U15 (N_15,In_260,In_1054);
or U16 (N_16,In_437,In_226);
or U17 (N_17,In_781,In_1029);
or U18 (N_18,In_552,In_1160);
or U19 (N_19,In_1427,In_382);
nand U20 (N_20,In_1337,In_182);
or U21 (N_21,In_551,In_42);
nand U22 (N_22,In_797,In_1390);
or U23 (N_23,In_76,In_729);
nor U24 (N_24,In_414,In_1419);
and U25 (N_25,In_1373,In_528);
nor U26 (N_26,In_707,In_851);
nand U27 (N_27,In_201,In_1051);
nand U28 (N_28,In_1275,In_1458);
nand U29 (N_29,In_933,In_1002);
nor U30 (N_30,In_1197,In_564);
and U31 (N_31,In_1243,In_218);
nand U32 (N_32,In_635,In_542);
and U33 (N_33,In_648,In_1222);
or U34 (N_34,In_259,In_1081);
nor U35 (N_35,In_1195,In_67);
nor U36 (N_36,In_1225,In_265);
nand U37 (N_37,In_189,In_1187);
and U38 (N_38,In_477,In_231);
nor U39 (N_39,In_1168,In_1167);
nor U40 (N_40,In_748,In_190);
nor U41 (N_41,In_789,In_1097);
or U42 (N_42,In_270,In_45);
nand U43 (N_43,In_823,In_1253);
nand U44 (N_44,In_868,In_756);
or U45 (N_45,In_483,In_1368);
nor U46 (N_46,In_644,In_329);
nor U47 (N_47,In_1402,In_827);
or U48 (N_48,In_1035,In_152);
or U49 (N_49,In_1291,In_565);
and U50 (N_50,In_1481,In_1150);
or U51 (N_51,In_98,In_213);
nand U52 (N_52,In_25,In_52);
and U53 (N_53,In_1418,In_350);
and U54 (N_54,In_1037,In_714);
or U55 (N_55,In_222,In_1162);
or U56 (N_56,In_148,In_1038);
or U57 (N_57,In_62,In_824);
or U58 (N_58,In_296,In_500);
nor U59 (N_59,In_88,In_1175);
nand U60 (N_60,In_604,In_818);
and U61 (N_61,In_280,In_1347);
nand U62 (N_62,In_1020,In_1351);
nand U63 (N_63,In_1272,In_765);
and U64 (N_64,In_1247,In_115);
nand U65 (N_65,In_1157,In_1058);
and U66 (N_66,In_848,In_864);
or U67 (N_67,In_833,In_1193);
nand U68 (N_68,In_924,In_1386);
and U69 (N_69,In_1204,In_576);
or U70 (N_70,In_123,In_1077);
or U71 (N_71,In_675,In_1228);
nand U72 (N_72,In_743,In_1389);
nor U73 (N_73,In_429,In_1305);
xnor U74 (N_74,In_220,In_898);
or U75 (N_75,In_285,In_703);
and U76 (N_76,In_1101,In_327);
and U77 (N_77,In_757,In_1053);
or U78 (N_78,In_232,In_255);
nor U79 (N_79,In_1493,In_1444);
nor U80 (N_80,In_1060,In_341);
or U81 (N_81,In_1359,In_1001);
nor U82 (N_82,In_464,In_186);
and U83 (N_83,In_1469,In_300);
and U84 (N_84,In_1268,In_172);
or U85 (N_85,In_205,In_1461);
or U86 (N_86,In_1464,In_1353);
nand U87 (N_87,In_1235,In_1179);
and U88 (N_88,In_1178,In_585);
nand U89 (N_89,In_1124,In_1487);
and U90 (N_90,In_466,In_1426);
nand U91 (N_91,In_816,In_455);
and U92 (N_92,In_1151,In_333);
or U93 (N_93,In_17,In_573);
or U94 (N_94,In_400,In_0);
and U95 (N_95,In_1290,In_1218);
and U96 (N_96,In_180,In_1457);
or U97 (N_97,In_277,In_490);
and U98 (N_98,In_209,In_849);
and U99 (N_99,In_1468,In_86);
or U100 (N_100,In_650,In_751);
or U101 (N_101,In_301,In_968);
nand U102 (N_102,In_1030,In_607);
or U103 (N_103,In_1176,In_1416);
or U104 (N_104,In_14,In_1063);
and U105 (N_105,In_484,In_264);
nor U106 (N_106,In_1489,In_695);
nand U107 (N_107,In_592,In_1278);
or U108 (N_108,In_705,In_151);
nand U109 (N_109,In_90,In_93);
nor U110 (N_110,In_363,In_931);
and U111 (N_111,In_1399,In_195);
nand U112 (N_112,In_1472,In_319);
nor U113 (N_113,In_836,In_1246);
or U114 (N_114,In_1266,In_872);
and U115 (N_115,In_601,In_562);
or U116 (N_116,In_38,In_1344);
and U117 (N_117,In_1092,In_1408);
or U118 (N_118,In_632,In_393);
nor U119 (N_119,In_309,In_909);
nand U120 (N_120,In_1448,In_223);
nand U121 (N_121,In_1201,In_1138);
nand U122 (N_122,In_352,In_411);
or U123 (N_123,In_124,In_1083);
and U124 (N_124,In_404,In_196);
nor U125 (N_125,In_877,In_728);
nand U126 (N_126,In_237,In_690);
and U127 (N_127,In_631,In_41);
nor U128 (N_128,In_853,In_206);
nor U129 (N_129,In_651,In_846);
nor U130 (N_130,In_896,In_621);
or U131 (N_131,In_951,In_646);
and U132 (N_132,In_1375,In_252);
and U133 (N_133,In_396,In_1057);
and U134 (N_134,In_1161,In_1379);
nor U135 (N_135,In_842,In_624);
and U136 (N_136,In_626,In_859);
nor U137 (N_137,In_1106,In_672);
nand U138 (N_138,In_12,In_181);
or U139 (N_139,In_699,In_200);
nor U140 (N_140,In_494,In_73);
and U141 (N_141,In_378,In_1123);
nor U142 (N_142,In_480,In_608);
nand U143 (N_143,In_1285,In_142);
nor U144 (N_144,In_1358,In_376);
nor U145 (N_145,In_1429,In_917);
and U146 (N_146,In_869,In_609);
nand U147 (N_147,In_1364,In_262);
nand U148 (N_148,In_902,In_517);
nor U149 (N_149,In_901,In_278);
nand U150 (N_150,In_1442,In_279);
and U151 (N_151,In_457,In_734);
nor U152 (N_152,In_1237,In_927);
or U153 (N_153,In_1384,In_778);
nand U154 (N_154,In_318,In_612);
or U155 (N_155,In_1192,In_111);
and U156 (N_156,In_183,In_1455);
and U157 (N_157,In_932,In_1211);
and U158 (N_158,In_597,In_1282);
nand U159 (N_159,In_1251,In_1074);
xor U160 (N_160,In_1028,In_671);
nor U161 (N_161,In_865,In_1424);
or U162 (N_162,In_143,In_923);
or U163 (N_163,In_101,In_605);
nor U164 (N_164,In_548,In_1329);
nor U165 (N_165,In_1104,In_1226);
and U166 (N_166,In_170,In_380);
nor U167 (N_167,In_1198,In_449);
or U168 (N_168,In_419,In_364);
and U169 (N_169,In_460,In_486);
or U170 (N_170,In_303,In_1477);
and U171 (N_171,In_964,In_345);
nand U172 (N_172,In_10,In_74);
nor U173 (N_173,In_1324,In_1169);
and U174 (N_174,In_595,In_990);
nor U175 (N_175,In_759,In_39);
nor U176 (N_176,In_779,In_563);
xnor U177 (N_177,In_239,In_764);
nand U178 (N_178,In_619,In_1122);
nor U179 (N_179,In_815,In_822);
nand U180 (N_180,In_735,In_1450);
nand U181 (N_181,In_787,In_89);
nor U182 (N_182,In_1465,In_745);
nor U183 (N_183,In_1079,In_792);
nand U184 (N_184,In_784,In_769);
or U185 (N_185,In_543,In_701);
nor U186 (N_186,In_1017,In_852);
or U187 (N_187,In_850,In_1146);
nand U188 (N_188,In_503,In_193);
and U189 (N_189,In_825,In_510);
and U190 (N_190,In_1100,In_991);
nor U191 (N_191,In_776,In_808);
nand U192 (N_192,In_1338,In_398);
nor U193 (N_193,In_969,In_2);
and U194 (N_194,In_294,In_240);
or U195 (N_195,In_1470,In_929);
or U196 (N_196,In_68,In_351);
nand U197 (N_197,In_938,In_254);
or U198 (N_198,In_1491,In_1127);
nand U199 (N_199,In_844,In_275);
and U200 (N_200,In_1260,In_1440);
nand U201 (N_201,In_811,In_1473);
or U202 (N_202,In_652,In_744);
or U203 (N_203,In_1062,In_912);
or U204 (N_204,In_1087,In_117);
nand U205 (N_205,In_356,In_439);
and U206 (N_206,In_31,In_1366);
or U207 (N_207,In_365,In_611);
nand U208 (N_208,In_717,In_770);
nand U209 (N_209,In_1476,In_1367);
and U210 (N_210,In_478,In_810);
nand U211 (N_211,In_1056,In_801);
nand U212 (N_212,In_282,In_112);
nor U213 (N_213,In_791,In_761);
and U214 (N_214,In_8,In_955);
and U215 (N_215,In_120,In_187);
or U216 (N_216,In_654,In_375);
nor U217 (N_217,In_1288,In_475);
or U218 (N_218,In_1327,In_1447);
and U219 (N_219,In_108,In_3);
nor U220 (N_220,In_557,In_1446);
and U221 (N_221,In_1279,In_965);
nor U222 (N_222,In_1380,In_758);
and U223 (N_223,In_267,In_890);
and U224 (N_224,In_1080,In_1300);
nand U225 (N_225,In_408,In_273);
or U226 (N_226,In_405,In_613);
and U227 (N_227,In_249,In_1262);
or U228 (N_228,In_1423,In_775);
nor U229 (N_229,In_1003,In_1016);
and U230 (N_230,In_698,In_1234);
or U231 (N_231,In_48,In_1188);
or U232 (N_232,In_907,In_246);
or U233 (N_233,In_772,In_1224);
xor U234 (N_234,In_403,In_317);
nor U235 (N_235,In_1349,In_313);
or U236 (N_236,In_184,In_1012);
nor U237 (N_237,In_905,In_311);
and U238 (N_238,In_1208,In_456);
or U239 (N_239,In_589,In_1027);
nor U240 (N_240,In_1065,In_293);
or U241 (N_241,In_1158,In_212);
or U242 (N_242,In_686,In_1021);
nand U243 (N_243,In_1374,In_953);
and U244 (N_244,In_963,In_786);
nand U245 (N_245,In_308,In_50);
nor U246 (N_246,In_1009,In_1369);
and U247 (N_247,In_1112,In_578);
nor U248 (N_248,In_133,In_526);
nor U249 (N_249,In_628,In_1050);
nor U250 (N_250,In_795,In_540);
nor U251 (N_251,In_855,In_1490);
nand U252 (N_252,In_230,In_536);
and U253 (N_253,In_625,In_803);
or U254 (N_254,In_569,In_620);
and U255 (N_255,In_243,In_474);
and U256 (N_256,In_1292,In_1041);
nand U257 (N_257,In_730,In_660);
nor U258 (N_258,In_1189,In_322);
nor U259 (N_259,In_434,In_1287);
nand U260 (N_260,In_344,In_1073);
nand U261 (N_261,In_1277,In_109);
nor U262 (N_262,In_1397,In_1276);
nor U263 (N_263,In_1335,In_1330);
nor U264 (N_264,In_1245,In_1174);
nand U265 (N_265,In_11,In_332);
or U266 (N_266,In_535,In_489);
nor U267 (N_267,In_753,In_347);
and U268 (N_268,In_1432,In_1042);
nand U269 (N_269,In_683,In_71);
and U270 (N_270,In_538,In_1181);
or U271 (N_271,In_369,In_1166);
nand U272 (N_272,In_1115,In_661);
nand U273 (N_273,In_331,In_998);
nor U274 (N_274,In_383,In_879);
nor U275 (N_275,In_1372,In_723);
nor U276 (N_276,In_337,In_740);
and U277 (N_277,In_1164,In_166);
and U278 (N_278,In_706,In_271);
nand U279 (N_279,In_981,In_72);
nor U280 (N_280,In_718,In_867);
nand U281 (N_281,In_961,In_330);
and U282 (N_282,In_338,In_391);
and U283 (N_283,In_502,In_247);
or U284 (N_284,In_420,In_627);
or U285 (N_285,In_568,In_992);
nand U286 (N_286,In_1240,In_559);
or U287 (N_287,In_372,In_83);
nand U288 (N_288,In_197,In_986);
and U289 (N_289,In_81,In_1154);
nand U290 (N_290,In_524,In_688);
nand U291 (N_291,In_424,In_684);
or U292 (N_292,In_1485,In_43);
nand U293 (N_293,In_141,In_549);
nor U294 (N_294,In_919,In_92);
and U295 (N_295,In_302,In_377);
nand U296 (N_296,In_722,In_1019);
nand U297 (N_297,In_689,In_579);
and U298 (N_298,In_1371,In_60);
nor U299 (N_299,In_739,In_451);
nor U300 (N_300,In_556,In_659);
and U301 (N_301,In_284,In_59);
nor U302 (N_302,In_1196,In_1126);
or U303 (N_303,In_614,In_208);
and U304 (N_304,In_422,In_574);
or U305 (N_305,In_1322,In_937);
or U306 (N_306,In_162,In_288);
and U307 (N_307,In_870,In_1496);
and U308 (N_308,In_1309,In_51);
nor U309 (N_309,In_27,In_1411);
or U310 (N_310,In_482,In_922);
or U311 (N_311,In_977,In_492);
nand U312 (N_312,In_1071,In_894);
and U313 (N_313,In_445,In_1387);
nand U314 (N_314,In_335,In_738);
and U315 (N_315,In_1325,In_866);
or U316 (N_316,In_219,In_1216);
nor U317 (N_317,In_415,In_407);
or U318 (N_318,In_397,In_643);
and U319 (N_319,In_518,In_1421);
nand U320 (N_320,In_34,In_1203);
nor U321 (N_321,In_721,In_885);
and U322 (N_322,In_947,In_447);
or U323 (N_323,In_1125,In_655);
and U324 (N_324,In_532,In_980);
nand U325 (N_325,In_908,In_1233);
nand U326 (N_326,In_1190,In_1241);
and U327 (N_327,In_725,In_719);
or U328 (N_328,In_204,In_1248);
or U329 (N_329,In_1069,In_916);
and U330 (N_330,In_28,In_583);
nand U331 (N_331,In_506,In_340);
nor U332 (N_332,In_1381,In_450);
or U333 (N_333,In_315,In_346);
nand U334 (N_334,In_1010,In_541);
xnor U335 (N_335,In_203,In_23);
and U336 (N_336,In_5,In_1334);
nand U337 (N_337,In_1348,In_920);
nand U338 (N_338,In_995,In_496);
and U339 (N_339,In_697,In_873);
nand U340 (N_340,In_153,In_895);
nand U341 (N_341,In_458,In_513);
and U342 (N_342,In_1156,In_834);
nand U343 (N_343,In_724,In_1215);
and U344 (N_344,In_1116,In_666);
or U345 (N_345,In_736,In_392);
or U346 (N_346,In_668,In_47);
nor U347 (N_347,In_1205,In_670);
and U348 (N_348,In_945,In_1438);
or U349 (N_349,In_600,In_1008);
or U350 (N_350,In_1018,In_1183);
or U351 (N_351,In_1346,In_566);
nor U352 (N_352,In_286,In_793);
nor U353 (N_353,In_1295,In_155);
or U354 (N_354,In_942,In_1425);
or U355 (N_355,In_432,In_1091);
xnor U356 (N_356,In_53,In_1257);
nand U357 (N_357,In_860,In_1378);
or U358 (N_358,In_747,In_1383);
and U359 (N_359,In_910,In_547);
nand U360 (N_360,In_463,In_80);
nor U361 (N_361,In_354,In_639);
or U362 (N_362,In_1441,In_617);
or U363 (N_363,In_1370,In_662);
or U364 (N_364,In_469,In_289);
nand U365 (N_365,In_537,In_946);
nand U366 (N_366,In_534,In_591);
nand U367 (N_367,In_202,In_87);
and U368 (N_368,In_1401,In_1113);
nor U369 (N_369,In_107,In_687);
nand U370 (N_370,In_948,In_305);
nand U371 (N_371,In_716,In_1043);
nand U372 (N_372,In_358,In_105);
nand U373 (N_373,In_394,In_1171);
nor U374 (N_374,In_826,In_857);
nand U375 (N_375,In_348,In_462);
and U376 (N_376,In_1177,In_641);
xnor U377 (N_377,In_1143,In_1297);
nor U378 (N_378,In_390,In_1170);
nor U379 (N_379,In_130,In_571);
and U380 (N_380,In_731,In_1471);
nor U381 (N_381,In_1492,In_838);
or U382 (N_382,In_134,In_245);
and U383 (N_383,In_1064,In_384);
nand U384 (N_384,In_1172,In_732);
nor U385 (N_385,In_975,In_427);
nand U386 (N_386,In_993,In_1213);
and U387 (N_387,In_610,In_712);
or U388 (N_388,In_49,In_978);
or U389 (N_389,In_516,In_957);
nor U390 (N_390,In_1086,In_1137);
or U391 (N_391,In_395,In_1267);
or U392 (N_392,In_1395,In_314);
or U393 (N_393,In_26,In_1439);
nor U394 (N_394,In_1155,In_830);
nand U395 (N_395,In_1252,In_622);
nand U396 (N_396,In_499,In_737);
nand U397 (N_397,In_653,In_935);
nand U398 (N_398,In_649,In_29);
nand U399 (N_399,In_173,In_299);
or U400 (N_400,In_742,In_1463);
nor U401 (N_401,In_1236,In_1130);
or U402 (N_402,In_914,In_799);
nor U403 (N_403,In_1453,In_679);
nor U404 (N_404,In_1159,In_276);
nor U405 (N_405,In_856,In_1049);
and U406 (N_406,In_244,In_523);
or U407 (N_407,In_362,In_216);
or U408 (N_408,In_1406,In_715);
and U409 (N_409,In_1034,In_623);
nor U410 (N_410,In_567,In_269);
or U411 (N_411,In_304,In_958);
nand U412 (N_412,In_310,In_1342);
and U413 (N_413,In_75,In_323);
or U414 (N_414,In_199,In_785);
or U415 (N_415,In_1403,In_1396);
nand U416 (N_416,In_884,In_1318);
and U417 (N_417,In_553,In_939);
or U418 (N_418,In_1452,In_307);
and U419 (N_419,In_291,In_1321);
and U420 (N_420,In_1117,In_144);
or U421 (N_421,In_1149,In_99);
or U422 (N_422,In_1298,In_1223);
and U423 (N_423,In_436,In_1283);
nand U424 (N_424,In_361,In_353);
and U425 (N_425,In_966,In_95);
or U426 (N_426,In_1294,In_656);
nand U427 (N_427,In_806,In_1296);
and U428 (N_428,In_1007,In_527);
nand U429 (N_429,In_667,In_1102);
or U430 (N_430,In_1333,In_821);
or U431 (N_431,In_292,In_1238);
nor U432 (N_432,In_1023,In_261);
nand U433 (N_433,In_1466,In_1120);
and U434 (N_434,In_1084,In_430);
nand U435 (N_435,In_1207,In_709);
or U436 (N_436,In_804,In_171);
nand U437 (N_437,In_749,In_515);
nand U438 (N_438,In_1200,In_248);
or U439 (N_439,In_1214,In_1362);
nand U440 (N_440,In_373,In_1180);
nor U441 (N_441,In_211,In_587);
nand U442 (N_442,In_1316,In_520);
nor U443 (N_443,In_642,In_1404);
nor U444 (N_444,In_533,In_572);
nor U445 (N_445,In_227,In_1147);
or U446 (N_446,In_943,In_371);
and U447 (N_447,In_174,In_1133);
or U448 (N_448,In_1109,In_633);
and U449 (N_449,In_191,In_835);
nor U450 (N_450,In_91,In_1339);
nand U451 (N_451,In_678,In_674);
nand U452 (N_452,In_1265,In_1099);
nand U453 (N_453,In_295,In_682);
nand U454 (N_454,In_77,In_1352);
and U455 (N_455,In_402,In_987);
and U456 (N_456,In_754,In_645);
nor U457 (N_457,In_343,In_1128);
or U458 (N_458,In_426,In_416);
nand U459 (N_459,In_1250,In_1264);
nand U460 (N_460,In_1345,In_97);
nand U461 (N_461,In_1317,In_1459);
nor U462 (N_462,In_956,In_36);
nor U463 (N_463,In_521,In_1036);
nor U464 (N_464,In_467,In_752);
xor U465 (N_465,In_802,In_593);
nor U466 (N_466,In_1420,In_994);
or U467 (N_467,In_167,In_545);
nor U468 (N_468,In_618,In_1249);
nand U469 (N_469,In_1412,In_94);
or U470 (N_470,In_606,In_433);
or U471 (N_471,In_1495,In_1497);
nand U472 (N_472,In_630,In_1061);
or U473 (N_473,In_1328,In_883);
or U474 (N_474,In_1132,In_70);
nand U475 (N_475,In_798,In_893);
or U476 (N_476,In_1385,In_1289);
nand U477 (N_477,In_949,In_511);
and U478 (N_478,In_580,In_127);
or U479 (N_479,In_125,In_1340);
nand U480 (N_480,In_741,In_1382);
and U481 (N_481,In_1070,In_1141);
nand U482 (N_482,In_268,In_1341);
and U483 (N_483,In_558,In_339);
or U484 (N_484,In_746,In_228);
or U485 (N_485,In_221,In_1059);
or U486 (N_486,In_1139,In_140);
nor U487 (N_487,In_1005,In_185);
and U488 (N_488,In_1273,In_509);
and U489 (N_489,In_479,In_1319);
nor U490 (N_490,In_122,In_970);
and U491 (N_491,In_1221,In_1410);
or U492 (N_492,In_888,In_839);
nor U493 (N_493,In_812,In_236);
and U494 (N_494,In_636,In_473);
nand U495 (N_495,In_767,In_1148);
or U496 (N_496,In_974,In_733);
nor U497 (N_497,In_198,In_952);
xnor U498 (N_498,In_904,In_512);
nor U499 (N_499,In_399,In_1436);
or U500 (N_500,In_1405,In_96);
nor U501 (N_501,In_570,In_615);
or U502 (N_502,In_1428,In_444);
or U503 (N_503,In_150,In_603);
nor U504 (N_504,In_78,In_582);
nand U505 (N_505,In_629,In_704);
and U506 (N_506,In_529,In_1271);
or U507 (N_507,In_1145,In_22);
or U508 (N_508,In_1015,In_104);
or U509 (N_509,In_1119,In_1355);
or U510 (N_510,In_35,In_750);
or U511 (N_511,In_1323,In_1217);
nand U512 (N_512,In_15,In_638);
or U513 (N_513,In_1365,In_1022);
nor U514 (N_514,In_1032,In_766);
nor U515 (N_515,In_413,In_283);
nor U516 (N_516,In_1098,In_409);
nor U517 (N_517,In_324,In_522);
nor U518 (N_518,In_1025,In_1094);
or U519 (N_519,In_428,In_1004);
nand U520 (N_520,In_913,In_366);
nor U521 (N_521,In_57,In_207);
nor U522 (N_522,In_177,In_481);
and U523 (N_523,In_1284,In_476);
xor U524 (N_524,In_1129,In_979);
nand U525 (N_525,In_1310,In_114);
or U526 (N_526,In_960,In_681);
nor U527 (N_527,In_326,In_6);
nand U528 (N_528,In_1072,In_491);
nor U529 (N_529,In_918,In_1407);
nand U530 (N_530,In_1093,In_814);
or U531 (N_531,In_768,In_982);
or U532 (N_532,In_1286,In_858);
nor U533 (N_533,In_1308,In_944);
nor U534 (N_534,In_1078,In_472);
and U535 (N_535,In_164,In_941);
or U536 (N_536,In_1209,In_1307);
nor U537 (N_537,In_325,In_316);
nand U538 (N_538,In_158,In_33);
nor U539 (N_539,In_1443,In_720);
and U540 (N_540,In_891,In_861);
and U541 (N_541,In_1082,In_1131);
nand U542 (N_542,In_1299,In_1409);
nor U543 (N_543,In_771,In_577);
or U544 (N_544,In_1363,In_1144);
nor U545 (N_545,In_774,In_539);
nand U546 (N_546,In_381,In_498);
or U547 (N_547,In_1075,In_1388);
or U548 (N_548,In_930,In_711);
or U549 (N_549,In_440,In_132);
nor U550 (N_550,In_387,In_983);
or U551 (N_551,In_1194,In_1173);
nand U552 (N_552,In_694,In_82);
and U553 (N_553,In_819,In_1088);
or U554 (N_554,In_755,In_514);
nor U555 (N_555,In_334,In_900);
or U556 (N_556,In_1392,In_320);
or U557 (N_557,In_1486,In_897);
and U558 (N_558,In_796,In_926);
and U559 (N_559,In_290,In_1430);
and U560 (N_560,In_1313,In_1445);
nor U561 (N_561,In_899,In_258);
nand U562 (N_562,In_224,In_163);
and U563 (N_563,In_1259,In_24);
and U564 (N_564,In_40,In_1263);
or U565 (N_565,In_119,In_1024);
nor U566 (N_566,In_1391,In_61);
or U567 (N_567,In_1244,In_1484);
or U568 (N_568,In_418,In_487);
nor U569 (N_569,In_546,In_875);
and U570 (N_570,In_84,In_453);
nor U571 (N_571,In_410,In_807);
nor U572 (N_572,In_417,In_599);
nor U573 (N_573,In_69,In_156);
nor U574 (N_574,In_845,In_306);
and U575 (N_575,In_575,In_336);
nor U576 (N_576,In_590,In_880);
and U577 (N_577,In_298,In_702);
or U578 (N_578,In_1256,In_1229);
nand U579 (N_579,In_680,In_1000);
or U580 (N_580,In_145,In_762);
xnor U581 (N_581,In_878,In_1255);
nand U582 (N_582,In_708,In_235);
or U583 (N_583,In_1498,In_452);
xor U584 (N_584,In_438,In_1011);
or U585 (N_585,In_137,In_726);
or U586 (N_586,In_1274,In_263);
and U587 (N_587,In_147,In_1231);
or U588 (N_588,In_1354,In_1046);
nand U589 (N_589,In_973,In_501);
nand U590 (N_590,In_525,In_1356);
or U591 (N_591,In_146,In_1033);
and U592 (N_592,In_954,In_1261);
or U593 (N_593,In_103,In_56);
and U594 (N_594,In_1,In_234);
and U595 (N_595,In_1067,In_1006);
or U596 (N_596,In_1361,In_443);
nand U597 (N_597,In_1343,In_1206);
nand U598 (N_598,In_210,In_256);
nor U599 (N_599,In_700,In_817);
nor U600 (N_600,In_66,In_959);
nand U601 (N_601,In_1040,In_178);
and U602 (N_602,In_554,In_459);
nand U603 (N_603,In_266,In_862);
nor U604 (N_604,In_657,In_1417);
nor U605 (N_605,In_1220,In_505);
nand U606 (N_606,In_1331,In_1230);
nand U607 (N_607,In_386,In_1210);
or U608 (N_608,In_7,In_116);
nor U609 (N_609,In_647,In_1332);
nor U610 (N_610,In_389,In_1449);
or U611 (N_611,In_54,In_713);
nand U612 (N_612,In_1431,In_829);
or U613 (N_613,In_677,In_832);
or U614 (N_614,In_1303,In_727);
and U615 (N_615,In_843,In_1191);
or U616 (N_616,In_1451,In_21);
and U617 (N_617,In_691,In_663);
nor U618 (N_618,In_800,In_876);
and U619 (N_619,In_1269,In_287);
or U620 (N_620,In_128,In_379);
and U621 (N_621,In_1152,In_1219);
nand U622 (N_622,In_1281,In_471);
nor U623 (N_623,In_1422,In_328);
and U624 (N_624,In_126,In_1326);
and U625 (N_625,In_176,In_1474);
nor U626 (N_626,In_544,In_100);
and U627 (N_627,In_1095,In_1414);
or U628 (N_628,In_1096,In_175);
or U629 (N_629,In_217,In_272);
or U630 (N_630,In_1415,In_435);
and U631 (N_631,In_911,In_1433);
or U632 (N_632,In_367,In_696);
nor U633 (N_633,In_1499,In_401);
or U634 (N_634,In_1479,In_470);
nand U635 (N_635,In_1184,In_928);
nor U636 (N_636,In_692,In_1475);
nor U637 (N_637,In_1227,In_531);
nand U638 (N_638,In_1302,In_242);
nor U639 (N_639,In_813,In_1052);
nand U640 (N_640,In_976,In_1153);
or U641 (N_641,In_693,In_1315);
nor U642 (N_642,In_1182,In_504);
nand U643 (N_643,In_1435,In_446);
or U644 (N_644,In_634,In_594);
and U645 (N_645,In_1306,In_1478);
nor U646 (N_646,In_773,In_442);
or U647 (N_647,In_598,In_355);
or U648 (N_648,In_18,In_154);
nor U649 (N_649,In_55,In_790);
nand U650 (N_650,In_431,In_794);
nor U651 (N_651,In_863,In_179);
and U652 (N_652,In_1108,In_1185);
nand U653 (N_653,In_1357,In_999);
nor U654 (N_654,In_588,In_493);
or U655 (N_655,In_550,In_673);
or U656 (N_656,In_1254,In_1232);
or U657 (N_657,In_1377,In_602);
or U658 (N_658,In_1044,In_229);
nand U659 (N_659,In_871,In_1242);
nand U660 (N_660,In_1068,In_497);
nor U661 (N_661,In_903,In_925);
or U662 (N_662,In_423,In_782);
nand U663 (N_663,In_58,In_406);
or U664 (N_664,In_63,In_1107);
or U665 (N_665,In_581,In_519);
or U666 (N_666,In_312,In_1048);
or U667 (N_667,In_138,In_637);
or U668 (N_668,In_454,In_32);
nand U669 (N_669,In_640,In_65);
nor U670 (N_670,In_669,In_30);
and U671 (N_671,In_1110,In_1270);
or U672 (N_672,In_887,In_1311);
nor U673 (N_673,In_1293,In_1045);
or U674 (N_674,In_665,In_214);
nand U675 (N_675,In_360,In_1360);
nor U676 (N_676,In_831,In_788);
and U677 (N_677,In_19,In_763);
nor U678 (N_678,In_840,In_906);
or U679 (N_679,In_385,In_79);
and U680 (N_680,In_1047,In_157);
nand U681 (N_681,In_321,In_760);
or U682 (N_682,In_710,In_251);
nor U683 (N_683,In_488,In_121);
and U684 (N_684,In_837,In_616);
and U685 (N_685,In_881,In_685);
and U686 (N_686,In_1066,In_1456);
nand U687 (N_687,In_1136,In_584);
and U688 (N_688,In_1026,In_297);
and U689 (N_689,In_1031,In_1165);
or U690 (N_690,In_495,In_461);
or U691 (N_691,In_342,In_4);
or U692 (N_692,In_238,In_448);
nor U693 (N_693,In_159,In_1089);
or U694 (N_694,In_1258,In_441);
and U695 (N_695,In_874,In_257);
and U696 (N_696,In_160,In_1199);
nor U697 (N_697,In_1320,In_37);
and U698 (N_698,In_828,In_1301);
or U699 (N_699,In_854,In_149);
nand U700 (N_700,In_984,In_85);
nor U701 (N_701,In_192,In_1280);
and U702 (N_702,In_1488,In_988);
nand U703 (N_703,In_997,In_136);
and U704 (N_704,In_777,In_664);
nand U705 (N_705,In_233,In_1014);
or U706 (N_706,In_892,In_561);
or U707 (N_707,In_359,In_169);
or U708 (N_708,In_241,In_113);
or U709 (N_709,In_465,In_1350);
or U710 (N_710,In_972,In_485);
or U711 (N_711,In_1103,In_809);
nor U712 (N_712,In_962,In_161);
nor U713 (N_713,In_847,In_1090);
and U714 (N_714,In_936,In_996);
or U715 (N_715,In_9,In_13);
nor U716 (N_716,In_274,In_44);
xnor U717 (N_717,In_530,In_118);
nor U718 (N_718,In_555,In_1202);
or U719 (N_719,In_110,In_507);
and U720 (N_720,In_586,In_1312);
and U721 (N_721,In_1482,In_1118);
nor U722 (N_722,In_1467,In_820);
nor U723 (N_723,In_783,In_934);
or U724 (N_724,In_889,In_468);
or U725 (N_725,In_421,In_658);
and U726 (N_726,In_46,In_165);
and U727 (N_727,In_1393,In_596);
nand U728 (N_728,In_940,In_357);
nand U729 (N_729,In_1437,In_253);
nor U730 (N_730,In_989,In_1239);
nor U731 (N_731,In_349,In_425);
or U732 (N_732,In_1076,In_1394);
nand U733 (N_733,In_1105,In_1483);
and U734 (N_734,In_1304,In_780);
and U735 (N_735,In_1140,In_374);
nor U736 (N_736,In_1055,In_1212);
nand U737 (N_737,In_129,In_1336);
and U738 (N_738,In_20,In_281);
or U739 (N_739,In_508,In_841);
and U740 (N_740,In_1454,In_102);
or U741 (N_741,In_1462,In_1460);
nand U742 (N_742,In_139,In_971);
and U743 (N_743,In_1400,In_676);
nor U744 (N_744,In_1142,In_1186);
nor U745 (N_745,In_225,In_1163);
nor U746 (N_746,In_388,In_1039);
and U747 (N_747,In_1376,In_168);
and U748 (N_748,In_412,In_1480);
and U749 (N_749,In_64,In_985);
and U750 (N_750,In_1261,In_1267);
and U751 (N_751,In_522,In_825);
nor U752 (N_752,In_721,In_142);
or U753 (N_753,In_1477,In_1114);
and U754 (N_754,In_614,In_531);
nor U755 (N_755,In_1310,In_190);
or U756 (N_756,In_345,In_1393);
or U757 (N_757,In_1425,In_280);
nor U758 (N_758,In_533,In_619);
or U759 (N_759,In_566,In_896);
and U760 (N_760,In_1405,In_1075);
and U761 (N_761,In_303,In_1014);
and U762 (N_762,In_926,In_1269);
nor U763 (N_763,In_451,In_969);
nand U764 (N_764,In_189,In_487);
nor U765 (N_765,In_1150,In_63);
and U766 (N_766,In_1000,In_1459);
and U767 (N_767,In_163,In_546);
or U768 (N_768,In_643,In_829);
or U769 (N_769,In_610,In_595);
nor U770 (N_770,In_65,In_1058);
nand U771 (N_771,In_1071,In_1318);
nor U772 (N_772,In_311,In_13);
nor U773 (N_773,In_436,In_505);
nor U774 (N_774,In_927,In_597);
nand U775 (N_775,In_61,In_187);
and U776 (N_776,In_460,In_1423);
or U777 (N_777,In_1174,In_391);
or U778 (N_778,In_1246,In_343);
nand U779 (N_779,In_1483,In_148);
nand U780 (N_780,In_625,In_7);
nor U781 (N_781,In_1030,In_1366);
nor U782 (N_782,In_1215,In_313);
nor U783 (N_783,In_959,In_176);
and U784 (N_784,In_1433,In_1000);
and U785 (N_785,In_493,In_1187);
or U786 (N_786,In_219,In_293);
nor U787 (N_787,In_612,In_978);
nor U788 (N_788,In_791,In_236);
or U789 (N_789,In_1477,In_1257);
or U790 (N_790,In_692,In_831);
nand U791 (N_791,In_1234,In_1411);
and U792 (N_792,In_1445,In_427);
nor U793 (N_793,In_1382,In_255);
nor U794 (N_794,In_890,In_1220);
or U795 (N_795,In_1187,In_1388);
and U796 (N_796,In_655,In_1059);
or U797 (N_797,In_605,In_870);
nor U798 (N_798,In_850,In_607);
and U799 (N_799,In_249,In_1354);
nor U800 (N_800,In_962,In_512);
or U801 (N_801,In_569,In_594);
and U802 (N_802,In_540,In_190);
or U803 (N_803,In_1226,In_785);
nor U804 (N_804,In_298,In_808);
nor U805 (N_805,In_1290,In_783);
nor U806 (N_806,In_609,In_1485);
nor U807 (N_807,In_1393,In_1127);
nand U808 (N_808,In_1408,In_647);
and U809 (N_809,In_382,In_283);
nor U810 (N_810,In_19,In_1280);
and U811 (N_811,In_1477,In_1395);
nor U812 (N_812,In_532,In_667);
and U813 (N_813,In_950,In_694);
or U814 (N_814,In_264,In_335);
nand U815 (N_815,In_67,In_1294);
and U816 (N_816,In_57,In_1045);
and U817 (N_817,In_943,In_917);
nand U818 (N_818,In_335,In_187);
nand U819 (N_819,In_1406,In_264);
and U820 (N_820,In_520,In_1209);
or U821 (N_821,In_435,In_91);
nand U822 (N_822,In_337,In_1415);
or U823 (N_823,In_60,In_1440);
nand U824 (N_824,In_507,In_691);
nand U825 (N_825,In_451,In_438);
or U826 (N_826,In_1129,In_659);
and U827 (N_827,In_1000,In_1341);
nand U828 (N_828,In_762,In_1394);
nand U829 (N_829,In_1223,In_783);
or U830 (N_830,In_455,In_954);
or U831 (N_831,In_1303,In_1034);
nand U832 (N_832,In_443,In_62);
nand U833 (N_833,In_1223,In_653);
and U834 (N_834,In_155,In_1395);
nand U835 (N_835,In_1312,In_512);
or U836 (N_836,In_332,In_968);
or U837 (N_837,In_1154,In_424);
nand U838 (N_838,In_922,In_356);
nand U839 (N_839,In_624,In_1227);
and U840 (N_840,In_161,In_486);
or U841 (N_841,In_1339,In_13);
and U842 (N_842,In_468,In_1121);
or U843 (N_843,In_552,In_634);
nor U844 (N_844,In_49,In_906);
nand U845 (N_845,In_921,In_1471);
and U846 (N_846,In_918,In_1364);
nand U847 (N_847,In_745,In_442);
nor U848 (N_848,In_202,In_626);
nand U849 (N_849,In_1137,In_754);
or U850 (N_850,In_1134,In_550);
and U851 (N_851,In_299,In_328);
nand U852 (N_852,In_1477,In_1027);
and U853 (N_853,In_276,In_1448);
and U854 (N_854,In_330,In_39);
nand U855 (N_855,In_55,In_987);
and U856 (N_856,In_514,In_835);
nor U857 (N_857,In_1471,In_633);
and U858 (N_858,In_213,In_299);
nand U859 (N_859,In_923,In_1035);
or U860 (N_860,In_1092,In_775);
nand U861 (N_861,In_491,In_910);
or U862 (N_862,In_1338,In_1118);
nor U863 (N_863,In_1128,In_493);
nand U864 (N_864,In_933,In_116);
and U865 (N_865,In_753,In_905);
nor U866 (N_866,In_1091,In_1314);
nand U867 (N_867,In_1392,In_15);
nand U868 (N_868,In_805,In_1263);
and U869 (N_869,In_98,In_1398);
and U870 (N_870,In_1295,In_673);
nand U871 (N_871,In_706,In_482);
nand U872 (N_872,In_1021,In_1186);
nand U873 (N_873,In_647,In_680);
or U874 (N_874,In_550,In_1074);
or U875 (N_875,In_593,In_655);
and U876 (N_876,In_600,In_606);
and U877 (N_877,In_1400,In_373);
or U878 (N_878,In_158,In_27);
nor U879 (N_879,In_724,In_1087);
and U880 (N_880,In_479,In_151);
and U881 (N_881,In_656,In_807);
and U882 (N_882,In_546,In_946);
nor U883 (N_883,In_927,In_1172);
or U884 (N_884,In_427,In_1130);
and U885 (N_885,In_357,In_1389);
nor U886 (N_886,In_672,In_275);
nor U887 (N_887,In_652,In_1460);
and U888 (N_888,In_1268,In_192);
xnor U889 (N_889,In_734,In_545);
nor U890 (N_890,In_1464,In_757);
nor U891 (N_891,In_98,In_312);
and U892 (N_892,In_1209,In_743);
and U893 (N_893,In_65,In_1107);
and U894 (N_894,In_740,In_1001);
or U895 (N_895,In_1146,In_264);
and U896 (N_896,In_128,In_1164);
and U897 (N_897,In_1135,In_105);
nor U898 (N_898,In_880,In_828);
nor U899 (N_899,In_1354,In_1358);
or U900 (N_900,In_87,In_1219);
nor U901 (N_901,In_43,In_682);
or U902 (N_902,In_1098,In_1379);
and U903 (N_903,In_1228,In_1014);
nor U904 (N_904,In_952,In_1348);
and U905 (N_905,In_553,In_387);
nand U906 (N_906,In_1439,In_1106);
and U907 (N_907,In_1165,In_504);
and U908 (N_908,In_256,In_972);
nand U909 (N_909,In_1128,In_724);
or U910 (N_910,In_493,In_1041);
nor U911 (N_911,In_280,In_1307);
nand U912 (N_912,In_527,In_229);
xnor U913 (N_913,In_573,In_429);
nand U914 (N_914,In_36,In_852);
and U915 (N_915,In_682,In_1030);
nor U916 (N_916,In_242,In_173);
nand U917 (N_917,In_492,In_942);
nand U918 (N_918,In_831,In_1493);
nor U919 (N_919,In_449,In_847);
nor U920 (N_920,In_835,In_77);
or U921 (N_921,In_1097,In_231);
nor U922 (N_922,In_1385,In_1263);
nand U923 (N_923,In_601,In_783);
and U924 (N_924,In_526,In_1058);
and U925 (N_925,In_335,In_1458);
nor U926 (N_926,In_522,In_1129);
or U927 (N_927,In_1394,In_615);
nand U928 (N_928,In_142,In_1462);
nand U929 (N_929,In_682,In_245);
and U930 (N_930,In_1472,In_1441);
nand U931 (N_931,In_466,In_988);
or U932 (N_932,In_1000,In_593);
nor U933 (N_933,In_451,In_231);
nor U934 (N_934,In_938,In_68);
nor U935 (N_935,In_236,In_285);
nand U936 (N_936,In_1029,In_879);
nand U937 (N_937,In_37,In_1017);
and U938 (N_938,In_155,In_571);
and U939 (N_939,In_772,In_636);
nor U940 (N_940,In_1390,In_1274);
nand U941 (N_941,In_1224,In_1261);
and U942 (N_942,In_400,In_712);
nand U943 (N_943,In_1346,In_1229);
or U944 (N_944,In_1357,In_466);
and U945 (N_945,In_1096,In_126);
nor U946 (N_946,In_999,In_939);
nor U947 (N_947,In_913,In_1294);
and U948 (N_948,In_180,In_1396);
or U949 (N_949,In_780,In_1297);
nor U950 (N_950,In_797,In_1195);
nand U951 (N_951,In_466,In_529);
or U952 (N_952,In_794,In_524);
or U953 (N_953,In_974,In_570);
nand U954 (N_954,In_486,In_61);
nor U955 (N_955,In_798,In_999);
nor U956 (N_956,In_1026,In_1409);
and U957 (N_957,In_848,In_1096);
and U958 (N_958,In_1414,In_476);
or U959 (N_959,In_1033,In_1272);
nor U960 (N_960,In_1323,In_799);
or U961 (N_961,In_193,In_427);
nor U962 (N_962,In_308,In_582);
and U963 (N_963,In_864,In_931);
nor U964 (N_964,In_890,In_1356);
and U965 (N_965,In_1055,In_1190);
nand U966 (N_966,In_703,In_942);
and U967 (N_967,In_763,In_1039);
or U968 (N_968,In_581,In_1226);
nand U969 (N_969,In_1499,In_946);
nor U970 (N_970,In_385,In_756);
nand U971 (N_971,In_475,In_1193);
or U972 (N_972,In_349,In_517);
and U973 (N_973,In_1428,In_1067);
nand U974 (N_974,In_641,In_1328);
nor U975 (N_975,In_581,In_470);
and U976 (N_976,In_349,In_27);
and U977 (N_977,In_299,In_633);
or U978 (N_978,In_994,In_334);
and U979 (N_979,In_1198,In_1233);
and U980 (N_980,In_231,In_481);
nand U981 (N_981,In_1197,In_173);
or U982 (N_982,In_464,In_525);
nor U983 (N_983,In_235,In_841);
or U984 (N_984,In_600,In_368);
nand U985 (N_985,In_911,In_88);
nand U986 (N_986,In_257,In_73);
nor U987 (N_987,In_168,In_652);
nand U988 (N_988,In_361,In_750);
nor U989 (N_989,In_249,In_7);
and U990 (N_990,In_425,In_1473);
and U991 (N_991,In_41,In_1133);
nand U992 (N_992,In_435,In_296);
and U993 (N_993,In_1044,In_1439);
nor U994 (N_994,In_289,In_462);
nor U995 (N_995,In_923,In_964);
and U996 (N_996,In_1453,In_1480);
and U997 (N_997,In_289,In_598);
and U998 (N_998,In_621,In_819);
xnor U999 (N_999,In_1397,In_187);
or U1000 (N_1000,In_1081,In_312);
nor U1001 (N_1001,In_1031,In_115);
and U1002 (N_1002,In_828,In_542);
nand U1003 (N_1003,In_1212,In_299);
or U1004 (N_1004,In_1420,In_1495);
and U1005 (N_1005,In_415,In_1133);
or U1006 (N_1006,In_764,In_537);
nor U1007 (N_1007,In_822,In_744);
or U1008 (N_1008,In_1174,In_570);
nand U1009 (N_1009,In_248,In_966);
nor U1010 (N_1010,In_1255,In_402);
and U1011 (N_1011,In_73,In_1121);
nor U1012 (N_1012,In_1114,In_1177);
or U1013 (N_1013,In_288,In_531);
and U1014 (N_1014,In_527,In_1342);
or U1015 (N_1015,In_1320,In_685);
and U1016 (N_1016,In_722,In_756);
nor U1017 (N_1017,In_1333,In_732);
nand U1018 (N_1018,In_1424,In_665);
nand U1019 (N_1019,In_1077,In_419);
nand U1020 (N_1020,In_476,In_879);
or U1021 (N_1021,In_1076,In_460);
or U1022 (N_1022,In_1318,In_480);
and U1023 (N_1023,In_883,In_442);
nor U1024 (N_1024,In_74,In_517);
nand U1025 (N_1025,In_418,In_751);
or U1026 (N_1026,In_1324,In_468);
nand U1027 (N_1027,In_406,In_920);
xor U1028 (N_1028,In_956,In_1469);
nand U1029 (N_1029,In_1440,In_1392);
nand U1030 (N_1030,In_687,In_234);
nor U1031 (N_1031,In_649,In_1014);
and U1032 (N_1032,In_255,In_12);
and U1033 (N_1033,In_303,In_937);
or U1034 (N_1034,In_129,In_1043);
and U1035 (N_1035,In_725,In_467);
nor U1036 (N_1036,In_371,In_1457);
nor U1037 (N_1037,In_643,In_186);
nand U1038 (N_1038,In_1261,In_884);
and U1039 (N_1039,In_652,In_1398);
and U1040 (N_1040,In_542,In_216);
nor U1041 (N_1041,In_1130,In_424);
nor U1042 (N_1042,In_1283,In_1081);
nor U1043 (N_1043,In_970,In_824);
and U1044 (N_1044,In_692,In_11);
nand U1045 (N_1045,In_1458,In_819);
nor U1046 (N_1046,In_1262,In_33);
nand U1047 (N_1047,In_394,In_600);
and U1048 (N_1048,In_167,In_355);
nand U1049 (N_1049,In_1350,In_1014);
or U1050 (N_1050,In_1300,In_1232);
nand U1051 (N_1051,In_1420,In_1343);
nor U1052 (N_1052,In_230,In_549);
nand U1053 (N_1053,In_177,In_1023);
nor U1054 (N_1054,In_1132,In_1419);
or U1055 (N_1055,In_1047,In_1251);
nor U1056 (N_1056,In_641,In_26);
and U1057 (N_1057,In_368,In_1380);
nor U1058 (N_1058,In_1150,In_567);
and U1059 (N_1059,In_894,In_323);
and U1060 (N_1060,In_1124,In_610);
or U1061 (N_1061,In_384,In_987);
nand U1062 (N_1062,In_1409,In_942);
nor U1063 (N_1063,In_591,In_1097);
nand U1064 (N_1064,In_318,In_95);
or U1065 (N_1065,In_839,In_27);
nand U1066 (N_1066,In_1157,In_887);
nor U1067 (N_1067,In_1456,In_471);
nor U1068 (N_1068,In_1416,In_1355);
nor U1069 (N_1069,In_833,In_633);
or U1070 (N_1070,In_393,In_315);
nand U1071 (N_1071,In_594,In_1248);
or U1072 (N_1072,In_417,In_1012);
and U1073 (N_1073,In_1427,In_1195);
or U1074 (N_1074,In_1478,In_1255);
nand U1075 (N_1075,In_735,In_1430);
nor U1076 (N_1076,In_1415,In_832);
or U1077 (N_1077,In_1311,In_1155);
or U1078 (N_1078,In_820,In_1069);
nand U1079 (N_1079,In_1009,In_76);
nand U1080 (N_1080,In_976,In_1090);
and U1081 (N_1081,In_1289,In_353);
or U1082 (N_1082,In_1183,In_817);
or U1083 (N_1083,In_1205,In_1217);
and U1084 (N_1084,In_1302,In_1102);
or U1085 (N_1085,In_1364,In_855);
nor U1086 (N_1086,In_1160,In_765);
nand U1087 (N_1087,In_44,In_615);
or U1088 (N_1088,In_890,In_800);
nand U1089 (N_1089,In_450,In_635);
nor U1090 (N_1090,In_1352,In_1212);
and U1091 (N_1091,In_1348,In_325);
or U1092 (N_1092,In_81,In_579);
and U1093 (N_1093,In_633,In_933);
or U1094 (N_1094,In_190,In_755);
nand U1095 (N_1095,In_1339,In_542);
nor U1096 (N_1096,In_257,In_288);
and U1097 (N_1097,In_552,In_781);
or U1098 (N_1098,In_221,In_576);
or U1099 (N_1099,In_1388,In_1413);
or U1100 (N_1100,In_527,In_366);
nand U1101 (N_1101,In_1104,In_930);
nand U1102 (N_1102,In_1188,In_901);
nor U1103 (N_1103,In_644,In_357);
and U1104 (N_1104,In_145,In_869);
and U1105 (N_1105,In_1037,In_751);
or U1106 (N_1106,In_1086,In_1450);
nand U1107 (N_1107,In_340,In_82);
nand U1108 (N_1108,In_1234,In_1276);
and U1109 (N_1109,In_171,In_627);
nand U1110 (N_1110,In_120,In_309);
nand U1111 (N_1111,In_646,In_79);
nand U1112 (N_1112,In_34,In_94);
and U1113 (N_1113,In_1055,In_806);
and U1114 (N_1114,In_1318,In_932);
and U1115 (N_1115,In_66,In_212);
or U1116 (N_1116,In_107,In_51);
or U1117 (N_1117,In_1291,In_885);
nand U1118 (N_1118,In_119,In_909);
nor U1119 (N_1119,In_1235,In_748);
and U1120 (N_1120,In_1218,In_902);
and U1121 (N_1121,In_427,In_1143);
nand U1122 (N_1122,In_86,In_733);
or U1123 (N_1123,In_310,In_214);
and U1124 (N_1124,In_625,In_1232);
and U1125 (N_1125,In_2,In_913);
nand U1126 (N_1126,In_1120,In_438);
and U1127 (N_1127,In_1443,In_146);
and U1128 (N_1128,In_1365,In_1328);
nand U1129 (N_1129,In_301,In_753);
nand U1130 (N_1130,In_195,In_1217);
and U1131 (N_1131,In_1144,In_197);
and U1132 (N_1132,In_377,In_1475);
and U1133 (N_1133,In_755,In_281);
nand U1134 (N_1134,In_1469,In_1006);
nand U1135 (N_1135,In_155,In_1398);
and U1136 (N_1136,In_356,In_1472);
nor U1137 (N_1137,In_810,In_929);
or U1138 (N_1138,In_262,In_763);
nor U1139 (N_1139,In_86,In_15);
or U1140 (N_1140,In_455,In_692);
and U1141 (N_1141,In_947,In_1169);
and U1142 (N_1142,In_1475,In_462);
nand U1143 (N_1143,In_978,In_112);
xor U1144 (N_1144,In_473,In_1397);
or U1145 (N_1145,In_941,In_564);
nand U1146 (N_1146,In_396,In_1347);
nor U1147 (N_1147,In_772,In_1377);
and U1148 (N_1148,In_1332,In_639);
nor U1149 (N_1149,In_1387,In_782);
or U1150 (N_1150,In_995,In_1430);
nor U1151 (N_1151,In_1298,In_900);
nor U1152 (N_1152,In_802,In_759);
nor U1153 (N_1153,In_498,In_198);
or U1154 (N_1154,In_202,In_442);
nor U1155 (N_1155,In_1490,In_1268);
nand U1156 (N_1156,In_448,In_119);
nor U1157 (N_1157,In_453,In_1072);
or U1158 (N_1158,In_854,In_1420);
nor U1159 (N_1159,In_98,In_10);
nor U1160 (N_1160,In_399,In_1295);
and U1161 (N_1161,In_548,In_352);
or U1162 (N_1162,In_271,In_777);
or U1163 (N_1163,In_1242,In_67);
or U1164 (N_1164,In_940,In_517);
and U1165 (N_1165,In_90,In_387);
or U1166 (N_1166,In_409,In_207);
nand U1167 (N_1167,In_1301,In_981);
nand U1168 (N_1168,In_920,In_820);
or U1169 (N_1169,In_1171,In_299);
and U1170 (N_1170,In_74,In_607);
nand U1171 (N_1171,In_611,In_1215);
and U1172 (N_1172,In_709,In_1231);
and U1173 (N_1173,In_184,In_978);
or U1174 (N_1174,In_1250,In_674);
or U1175 (N_1175,In_431,In_1125);
nor U1176 (N_1176,In_1113,In_1314);
or U1177 (N_1177,In_443,In_746);
and U1178 (N_1178,In_165,In_1076);
nand U1179 (N_1179,In_1129,In_771);
or U1180 (N_1180,In_266,In_1084);
nor U1181 (N_1181,In_747,In_524);
and U1182 (N_1182,In_839,In_801);
nand U1183 (N_1183,In_294,In_1159);
nor U1184 (N_1184,In_625,In_80);
or U1185 (N_1185,In_843,In_1278);
nand U1186 (N_1186,In_323,In_655);
nand U1187 (N_1187,In_1414,In_708);
and U1188 (N_1188,In_946,In_963);
nor U1189 (N_1189,In_519,In_454);
nor U1190 (N_1190,In_1353,In_728);
nand U1191 (N_1191,In_286,In_1444);
or U1192 (N_1192,In_1318,In_1428);
or U1193 (N_1193,In_810,In_2);
and U1194 (N_1194,In_1253,In_613);
nand U1195 (N_1195,In_1094,In_15);
nor U1196 (N_1196,In_1442,In_1302);
or U1197 (N_1197,In_921,In_967);
nand U1198 (N_1198,In_766,In_315);
or U1199 (N_1199,In_795,In_1012);
and U1200 (N_1200,In_771,In_582);
and U1201 (N_1201,In_337,In_968);
nor U1202 (N_1202,In_506,In_586);
or U1203 (N_1203,In_1198,In_148);
and U1204 (N_1204,In_1179,In_567);
nor U1205 (N_1205,In_948,In_1471);
nand U1206 (N_1206,In_55,In_111);
nand U1207 (N_1207,In_181,In_1408);
nor U1208 (N_1208,In_488,In_1156);
nand U1209 (N_1209,In_860,In_416);
nand U1210 (N_1210,In_1008,In_850);
and U1211 (N_1211,In_1462,In_1237);
and U1212 (N_1212,In_1484,In_1238);
nor U1213 (N_1213,In_1351,In_521);
or U1214 (N_1214,In_1018,In_628);
nand U1215 (N_1215,In_54,In_987);
nor U1216 (N_1216,In_1449,In_614);
nand U1217 (N_1217,In_1414,In_374);
nor U1218 (N_1218,In_176,In_1187);
or U1219 (N_1219,In_437,In_352);
nand U1220 (N_1220,In_484,In_665);
nor U1221 (N_1221,In_1205,In_208);
and U1222 (N_1222,In_15,In_585);
and U1223 (N_1223,In_733,In_1329);
nor U1224 (N_1224,In_122,In_385);
nand U1225 (N_1225,In_1016,In_173);
nor U1226 (N_1226,In_687,In_97);
or U1227 (N_1227,In_605,In_1397);
or U1228 (N_1228,In_43,In_821);
nand U1229 (N_1229,In_449,In_171);
and U1230 (N_1230,In_666,In_1316);
or U1231 (N_1231,In_10,In_654);
and U1232 (N_1232,In_1096,In_2);
or U1233 (N_1233,In_832,In_619);
nor U1234 (N_1234,In_239,In_1287);
nand U1235 (N_1235,In_934,In_37);
nor U1236 (N_1236,In_473,In_887);
nor U1237 (N_1237,In_860,In_605);
or U1238 (N_1238,In_838,In_756);
nor U1239 (N_1239,In_73,In_1450);
and U1240 (N_1240,In_645,In_36);
nand U1241 (N_1241,In_718,In_1193);
or U1242 (N_1242,In_265,In_1035);
nand U1243 (N_1243,In_194,In_1472);
nor U1244 (N_1244,In_969,In_342);
nand U1245 (N_1245,In_436,In_81);
xor U1246 (N_1246,In_357,In_1372);
or U1247 (N_1247,In_114,In_177);
or U1248 (N_1248,In_969,In_133);
or U1249 (N_1249,In_794,In_1160);
or U1250 (N_1250,In_697,In_66);
or U1251 (N_1251,In_530,In_636);
nor U1252 (N_1252,In_374,In_1098);
or U1253 (N_1253,In_485,In_1425);
nand U1254 (N_1254,In_1378,In_544);
and U1255 (N_1255,In_749,In_720);
and U1256 (N_1256,In_188,In_34);
nand U1257 (N_1257,In_329,In_918);
and U1258 (N_1258,In_1104,In_594);
nor U1259 (N_1259,In_512,In_1482);
nor U1260 (N_1260,In_1217,In_616);
or U1261 (N_1261,In_527,In_394);
or U1262 (N_1262,In_645,In_266);
xnor U1263 (N_1263,In_531,In_643);
nor U1264 (N_1264,In_1075,In_489);
or U1265 (N_1265,In_526,In_359);
and U1266 (N_1266,In_231,In_1042);
or U1267 (N_1267,In_537,In_742);
or U1268 (N_1268,In_1170,In_507);
nand U1269 (N_1269,In_280,In_1109);
nand U1270 (N_1270,In_552,In_465);
and U1271 (N_1271,In_312,In_722);
and U1272 (N_1272,In_113,In_498);
nand U1273 (N_1273,In_1455,In_309);
or U1274 (N_1274,In_1197,In_1138);
and U1275 (N_1275,In_1313,In_125);
nand U1276 (N_1276,In_1168,In_616);
nand U1277 (N_1277,In_1263,In_1074);
and U1278 (N_1278,In_747,In_450);
nor U1279 (N_1279,In_655,In_254);
nor U1280 (N_1280,In_333,In_583);
and U1281 (N_1281,In_350,In_1118);
nor U1282 (N_1282,In_338,In_1229);
nand U1283 (N_1283,In_4,In_1127);
and U1284 (N_1284,In_1147,In_276);
or U1285 (N_1285,In_1435,In_220);
nor U1286 (N_1286,In_227,In_150);
or U1287 (N_1287,In_413,In_1052);
and U1288 (N_1288,In_1238,In_1382);
or U1289 (N_1289,In_764,In_19);
or U1290 (N_1290,In_1156,In_693);
nand U1291 (N_1291,In_99,In_871);
or U1292 (N_1292,In_1068,In_1028);
nand U1293 (N_1293,In_1415,In_52);
nor U1294 (N_1294,In_428,In_121);
nand U1295 (N_1295,In_985,In_124);
nand U1296 (N_1296,In_177,In_1277);
nor U1297 (N_1297,In_1343,In_336);
or U1298 (N_1298,In_1039,In_844);
nand U1299 (N_1299,In_512,In_155);
and U1300 (N_1300,In_774,In_957);
and U1301 (N_1301,In_1406,In_1487);
nor U1302 (N_1302,In_404,In_542);
or U1303 (N_1303,In_497,In_104);
and U1304 (N_1304,In_362,In_1445);
nor U1305 (N_1305,In_942,In_1259);
nand U1306 (N_1306,In_211,In_364);
nand U1307 (N_1307,In_209,In_314);
nor U1308 (N_1308,In_1031,In_1221);
or U1309 (N_1309,In_691,In_327);
nand U1310 (N_1310,In_1061,In_1244);
nor U1311 (N_1311,In_386,In_1389);
nand U1312 (N_1312,In_343,In_123);
or U1313 (N_1313,In_392,In_176);
and U1314 (N_1314,In_257,In_1379);
and U1315 (N_1315,In_162,In_989);
and U1316 (N_1316,In_1332,In_192);
nor U1317 (N_1317,In_828,In_686);
and U1318 (N_1318,In_636,In_607);
or U1319 (N_1319,In_996,In_1274);
nor U1320 (N_1320,In_1136,In_711);
or U1321 (N_1321,In_21,In_160);
or U1322 (N_1322,In_1024,In_1389);
nor U1323 (N_1323,In_365,In_1286);
nor U1324 (N_1324,In_613,In_908);
nand U1325 (N_1325,In_1113,In_982);
nor U1326 (N_1326,In_1257,In_439);
nor U1327 (N_1327,In_1337,In_1129);
nand U1328 (N_1328,In_793,In_239);
or U1329 (N_1329,In_706,In_1006);
or U1330 (N_1330,In_807,In_1213);
nor U1331 (N_1331,In_451,In_1400);
or U1332 (N_1332,In_584,In_165);
nor U1333 (N_1333,In_559,In_142);
nand U1334 (N_1334,In_303,In_925);
or U1335 (N_1335,In_1483,In_595);
and U1336 (N_1336,In_990,In_449);
nand U1337 (N_1337,In_939,In_618);
and U1338 (N_1338,In_1073,In_1326);
nor U1339 (N_1339,In_687,In_1269);
and U1340 (N_1340,In_81,In_355);
or U1341 (N_1341,In_221,In_13);
or U1342 (N_1342,In_1013,In_215);
and U1343 (N_1343,In_211,In_612);
nand U1344 (N_1344,In_1199,In_152);
or U1345 (N_1345,In_374,In_829);
and U1346 (N_1346,In_533,In_462);
nand U1347 (N_1347,In_1220,In_1442);
nor U1348 (N_1348,In_1344,In_1062);
nand U1349 (N_1349,In_1344,In_79);
or U1350 (N_1350,In_1390,In_1186);
xnor U1351 (N_1351,In_257,In_764);
and U1352 (N_1352,In_1208,In_402);
and U1353 (N_1353,In_771,In_185);
or U1354 (N_1354,In_1407,In_1299);
or U1355 (N_1355,In_1083,In_1205);
and U1356 (N_1356,In_97,In_1215);
nor U1357 (N_1357,In_945,In_767);
and U1358 (N_1358,In_150,In_687);
nor U1359 (N_1359,In_867,In_161);
nor U1360 (N_1360,In_1114,In_979);
or U1361 (N_1361,In_523,In_209);
nand U1362 (N_1362,In_41,In_53);
nor U1363 (N_1363,In_475,In_614);
and U1364 (N_1364,In_1230,In_1138);
or U1365 (N_1365,In_831,In_204);
nor U1366 (N_1366,In_507,In_485);
nand U1367 (N_1367,In_1016,In_961);
and U1368 (N_1368,In_1485,In_1305);
xnor U1369 (N_1369,In_697,In_796);
or U1370 (N_1370,In_1132,In_660);
or U1371 (N_1371,In_26,In_67);
nand U1372 (N_1372,In_477,In_125);
nor U1373 (N_1373,In_141,In_1138);
nand U1374 (N_1374,In_320,In_297);
and U1375 (N_1375,In_1218,In_827);
nand U1376 (N_1376,In_418,In_1468);
and U1377 (N_1377,In_988,In_304);
or U1378 (N_1378,In_824,In_988);
nand U1379 (N_1379,In_780,In_420);
nor U1380 (N_1380,In_622,In_196);
nand U1381 (N_1381,In_1058,In_1162);
and U1382 (N_1382,In_257,In_1157);
nor U1383 (N_1383,In_1094,In_1268);
nor U1384 (N_1384,In_1079,In_261);
and U1385 (N_1385,In_375,In_1346);
nor U1386 (N_1386,In_59,In_901);
and U1387 (N_1387,In_180,In_710);
nand U1388 (N_1388,In_1121,In_163);
nor U1389 (N_1389,In_1445,In_639);
or U1390 (N_1390,In_719,In_598);
and U1391 (N_1391,In_295,In_116);
nand U1392 (N_1392,In_305,In_1099);
nand U1393 (N_1393,In_551,In_1245);
nand U1394 (N_1394,In_431,In_571);
nor U1395 (N_1395,In_600,In_1238);
nor U1396 (N_1396,In_671,In_823);
or U1397 (N_1397,In_1168,In_1315);
or U1398 (N_1398,In_413,In_231);
or U1399 (N_1399,In_1262,In_605);
or U1400 (N_1400,In_386,In_358);
nand U1401 (N_1401,In_427,In_62);
or U1402 (N_1402,In_1009,In_658);
and U1403 (N_1403,In_1178,In_940);
nand U1404 (N_1404,In_491,In_762);
nor U1405 (N_1405,In_1224,In_236);
nand U1406 (N_1406,In_458,In_92);
nor U1407 (N_1407,In_1341,In_1408);
nand U1408 (N_1408,In_327,In_475);
or U1409 (N_1409,In_1096,In_668);
nand U1410 (N_1410,In_1253,In_291);
nor U1411 (N_1411,In_348,In_899);
or U1412 (N_1412,In_543,In_682);
and U1413 (N_1413,In_400,In_966);
nor U1414 (N_1414,In_1145,In_173);
or U1415 (N_1415,In_1258,In_84);
nor U1416 (N_1416,In_304,In_809);
nor U1417 (N_1417,In_60,In_1139);
nand U1418 (N_1418,In_578,In_1462);
or U1419 (N_1419,In_971,In_748);
nor U1420 (N_1420,In_914,In_257);
nand U1421 (N_1421,In_174,In_202);
nand U1422 (N_1422,In_1143,In_747);
or U1423 (N_1423,In_79,In_382);
or U1424 (N_1424,In_214,In_246);
xor U1425 (N_1425,In_1485,In_336);
nand U1426 (N_1426,In_507,In_1348);
nor U1427 (N_1427,In_262,In_1231);
nor U1428 (N_1428,In_736,In_1309);
nand U1429 (N_1429,In_1106,In_841);
and U1430 (N_1430,In_306,In_716);
or U1431 (N_1431,In_1372,In_99);
nand U1432 (N_1432,In_1489,In_67);
or U1433 (N_1433,In_915,In_1459);
nor U1434 (N_1434,In_1459,In_300);
and U1435 (N_1435,In_10,In_814);
nor U1436 (N_1436,In_1332,In_680);
nand U1437 (N_1437,In_353,In_1474);
and U1438 (N_1438,In_688,In_1221);
nor U1439 (N_1439,In_599,In_1191);
or U1440 (N_1440,In_247,In_281);
or U1441 (N_1441,In_900,In_351);
or U1442 (N_1442,In_1040,In_735);
or U1443 (N_1443,In_1287,In_965);
nor U1444 (N_1444,In_899,In_1336);
nand U1445 (N_1445,In_1451,In_1260);
nor U1446 (N_1446,In_1176,In_80);
nor U1447 (N_1447,In_547,In_191);
nand U1448 (N_1448,In_1418,In_1066);
nand U1449 (N_1449,In_1280,In_152);
nand U1450 (N_1450,In_46,In_906);
and U1451 (N_1451,In_1046,In_959);
nand U1452 (N_1452,In_64,In_523);
nand U1453 (N_1453,In_498,In_395);
or U1454 (N_1454,In_1140,In_854);
nand U1455 (N_1455,In_1337,In_335);
and U1456 (N_1456,In_116,In_1109);
nand U1457 (N_1457,In_1197,In_98);
nor U1458 (N_1458,In_24,In_1470);
nor U1459 (N_1459,In_971,In_104);
nor U1460 (N_1460,In_55,In_1228);
and U1461 (N_1461,In_477,In_1076);
nor U1462 (N_1462,In_1204,In_915);
or U1463 (N_1463,In_146,In_78);
nand U1464 (N_1464,In_1132,In_403);
and U1465 (N_1465,In_1236,In_1370);
and U1466 (N_1466,In_153,In_913);
nor U1467 (N_1467,In_1223,In_987);
nand U1468 (N_1468,In_642,In_425);
and U1469 (N_1469,In_401,In_57);
nand U1470 (N_1470,In_598,In_1001);
and U1471 (N_1471,In_178,In_1222);
and U1472 (N_1472,In_397,In_59);
nor U1473 (N_1473,In_566,In_1273);
nand U1474 (N_1474,In_1436,In_1296);
nor U1475 (N_1475,In_470,In_19);
or U1476 (N_1476,In_751,In_405);
or U1477 (N_1477,In_450,In_1363);
or U1478 (N_1478,In_721,In_486);
and U1479 (N_1479,In_873,In_793);
and U1480 (N_1480,In_681,In_15);
and U1481 (N_1481,In_827,In_714);
or U1482 (N_1482,In_248,In_1470);
nor U1483 (N_1483,In_1113,In_186);
or U1484 (N_1484,In_866,In_942);
and U1485 (N_1485,In_278,In_551);
nor U1486 (N_1486,In_53,In_1175);
or U1487 (N_1487,In_855,In_164);
and U1488 (N_1488,In_1091,In_1031);
and U1489 (N_1489,In_1373,In_891);
or U1490 (N_1490,In_310,In_1225);
nand U1491 (N_1491,In_874,In_527);
nand U1492 (N_1492,In_1014,In_276);
nand U1493 (N_1493,In_259,In_700);
or U1494 (N_1494,In_1274,In_1420);
or U1495 (N_1495,In_1064,In_297);
nor U1496 (N_1496,In_224,In_201);
or U1497 (N_1497,In_1115,In_1335);
and U1498 (N_1498,In_934,In_1454);
nand U1499 (N_1499,In_1420,In_1149);
and U1500 (N_1500,N_163,N_427);
nor U1501 (N_1501,N_205,N_2);
or U1502 (N_1502,N_306,N_371);
nor U1503 (N_1503,N_358,N_1424);
and U1504 (N_1504,N_588,N_361);
and U1505 (N_1505,N_193,N_5);
nand U1506 (N_1506,N_373,N_445);
nand U1507 (N_1507,N_1413,N_362);
nor U1508 (N_1508,N_913,N_58);
nand U1509 (N_1509,N_1171,N_90);
and U1510 (N_1510,N_1197,N_1081);
and U1511 (N_1511,N_679,N_111);
and U1512 (N_1512,N_1407,N_98);
or U1513 (N_1513,N_949,N_1307);
or U1514 (N_1514,N_250,N_1003);
nor U1515 (N_1515,N_484,N_165);
nor U1516 (N_1516,N_904,N_1093);
nand U1517 (N_1517,N_566,N_198);
or U1518 (N_1518,N_118,N_855);
or U1519 (N_1519,N_1417,N_1135);
and U1520 (N_1520,N_1042,N_1000);
and U1521 (N_1521,N_359,N_737);
and U1522 (N_1522,N_342,N_286);
and U1523 (N_1523,N_208,N_1066);
nor U1524 (N_1524,N_1087,N_1217);
and U1525 (N_1525,N_496,N_655);
and U1526 (N_1526,N_754,N_334);
nand U1527 (N_1527,N_89,N_1123);
nor U1528 (N_1528,N_1484,N_860);
nor U1529 (N_1529,N_460,N_1129);
or U1530 (N_1530,N_652,N_1422);
nor U1531 (N_1531,N_1305,N_764);
nor U1532 (N_1532,N_311,N_388);
or U1533 (N_1533,N_1258,N_987);
nor U1534 (N_1534,N_1026,N_1226);
and U1535 (N_1535,N_1437,N_922);
nand U1536 (N_1536,N_866,N_835);
or U1537 (N_1537,N_573,N_278);
nand U1538 (N_1538,N_1419,N_967);
nor U1539 (N_1539,N_1256,N_1368);
nor U1540 (N_1540,N_11,N_788);
nor U1541 (N_1541,N_390,N_1266);
nor U1542 (N_1542,N_554,N_37);
nor U1543 (N_1543,N_352,N_221);
or U1544 (N_1544,N_826,N_676);
or U1545 (N_1545,N_104,N_106);
or U1546 (N_1546,N_374,N_216);
nand U1547 (N_1547,N_736,N_762);
or U1548 (N_1548,N_513,N_418);
or U1549 (N_1549,N_919,N_1382);
nor U1550 (N_1550,N_1487,N_447);
nand U1551 (N_1551,N_295,N_529);
nand U1552 (N_1552,N_1240,N_551);
nand U1553 (N_1553,N_1239,N_211);
and U1554 (N_1554,N_616,N_1136);
or U1555 (N_1555,N_607,N_766);
nand U1556 (N_1556,N_844,N_91);
and U1557 (N_1557,N_1331,N_853);
nand U1558 (N_1558,N_833,N_1139);
or U1559 (N_1559,N_915,N_316);
or U1560 (N_1560,N_631,N_717);
and U1561 (N_1561,N_1015,N_82);
nor U1562 (N_1562,N_950,N_1128);
nor U1563 (N_1563,N_813,N_1109);
and U1564 (N_1564,N_333,N_173);
nand U1565 (N_1565,N_559,N_1450);
or U1566 (N_1566,N_271,N_617);
and U1567 (N_1567,N_71,N_1145);
nor U1568 (N_1568,N_688,N_1200);
or U1569 (N_1569,N_391,N_121);
and U1570 (N_1570,N_206,N_673);
and U1571 (N_1571,N_647,N_1435);
or U1572 (N_1572,N_1350,N_264);
nand U1573 (N_1573,N_642,N_629);
and U1574 (N_1574,N_1257,N_579);
xnor U1575 (N_1575,N_451,N_870);
or U1576 (N_1576,N_452,N_1065);
nand U1577 (N_1577,N_419,N_1308);
or U1578 (N_1578,N_758,N_694);
nand U1579 (N_1579,N_479,N_544);
nand U1580 (N_1580,N_1489,N_1027);
nor U1581 (N_1581,N_439,N_738);
and U1582 (N_1582,N_428,N_299);
and U1583 (N_1583,N_1159,N_882);
or U1584 (N_1584,N_847,N_492);
nor U1585 (N_1585,N_680,N_220);
or U1586 (N_1586,N_1259,N_725);
or U1587 (N_1587,N_751,N_908);
nor U1588 (N_1588,N_572,N_257);
or U1589 (N_1589,N_819,N_718);
nor U1590 (N_1590,N_901,N_1161);
or U1591 (N_1591,N_719,N_321);
or U1592 (N_1592,N_594,N_848);
nor U1593 (N_1593,N_1119,N_666);
nand U1594 (N_1594,N_1048,N_760);
nand U1595 (N_1595,N_356,N_1034);
nor U1596 (N_1596,N_809,N_574);
nand U1597 (N_1597,N_734,N_437);
nor U1598 (N_1598,N_849,N_1383);
xnor U1599 (N_1599,N_910,N_836);
or U1600 (N_1600,N_103,N_1190);
or U1601 (N_1601,N_1233,N_400);
xnor U1602 (N_1602,N_33,N_20);
and U1603 (N_1603,N_35,N_1323);
nor U1604 (N_1604,N_1432,N_255);
nand U1605 (N_1605,N_494,N_76);
and U1606 (N_1606,N_567,N_521);
nand U1607 (N_1607,N_1423,N_1284);
or U1608 (N_1608,N_1204,N_41);
nand U1609 (N_1609,N_234,N_1293);
nand U1610 (N_1610,N_1398,N_1112);
and U1611 (N_1611,N_548,N_1211);
or U1612 (N_1612,N_202,N_223);
nand U1613 (N_1613,N_183,N_55);
nand U1614 (N_1614,N_473,N_97);
or U1615 (N_1615,N_998,N_863);
and U1616 (N_1616,N_959,N_520);
nor U1617 (N_1617,N_1245,N_805);
or U1618 (N_1618,N_1189,N_335);
nor U1619 (N_1619,N_381,N_1300);
nand U1620 (N_1620,N_692,N_75);
and U1621 (N_1621,N_477,N_525);
nor U1622 (N_1622,N_269,N_1446);
and U1623 (N_1623,N_1184,N_137);
nand U1624 (N_1624,N_774,N_1374);
nor U1625 (N_1625,N_1228,N_899);
nor U1626 (N_1626,N_409,N_1409);
nor U1627 (N_1627,N_219,N_1169);
nand U1628 (N_1628,N_57,N_867);
and U1629 (N_1629,N_538,N_1277);
nor U1630 (N_1630,N_1491,N_258);
and U1631 (N_1631,N_948,N_1358);
nor U1632 (N_1632,N_1388,N_389);
and U1633 (N_1633,N_8,N_1349);
and U1634 (N_1634,N_743,N_1203);
nor U1635 (N_1635,N_136,N_1143);
nand U1636 (N_1636,N_1411,N_1131);
and U1637 (N_1637,N_620,N_667);
or U1638 (N_1638,N_968,N_589);
nor U1639 (N_1639,N_480,N_1214);
nand U1640 (N_1640,N_831,N_1219);
or U1641 (N_1641,N_348,N_285);
and U1642 (N_1642,N_615,N_1478);
or U1643 (N_1643,N_1325,N_931);
nand U1644 (N_1644,N_808,N_1166);
nor U1645 (N_1645,N_172,N_293);
or U1646 (N_1646,N_1077,N_896);
nor U1647 (N_1647,N_14,N_197);
nor U1648 (N_1648,N_1071,N_527);
and U1649 (N_1649,N_481,N_38);
and U1650 (N_1650,N_1242,N_1140);
or U1651 (N_1651,N_524,N_95);
nor U1652 (N_1652,N_1352,N_310);
nor U1653 (N_1653,N_126,N_29);
or U1654 (N_1654,N_1188,N_735);
nand U1655 (N_1655,N_545,N_1414);
and U1656 (N_1656,N_564,N_53);
nor U1657 (N_1657,N_792,N_979);
xnor U1658 (N_1658,N_128,N_99);
nor U1659 (N_1659,N_86,N_581);
nand U1660 (N_1660,N_174,N_1229);
nand U1661 (N_1661,N_937,N_537);
and U1662 (N_1662,N_1311,N_982);
nand U1663 (N_1663,N_984,N_974);
or U1664 (N_1664,N_338,N_304);
nor U1665 (N_1665,N_244,N_1223);
and U1666 (N_1666,N_1141,N_812);
and U1667 (N_1667,N_94,N_143);
and U1668 (N_1668,N_516,N_739);
or U1669 (N_1669,N_778,N_330);
or U1670 (N_1670,N_996,N_1443);
nand U1671 (N_1671,N_112,N_318);
and U1672 (N_1672,N_508,N_113);
and U1673 (N_1673,N_73,N_450);
and U1674 (N_1674,N_823,N_555);
or U1675 (N_1675,N_355,N_1336);
or U1676 (N_1676,N_145,N_252);
nand U1677 (N_1677,N_552,N_19);
nor U1678 (N_1678,N_79,N_1154);
nand U1679 (N_1679,N_324,N_156);
nor U1680 (N_1680,N_889,N_1039);
or U1681 (N_1681,N_52,N_983);
or U1682 (N_1682,N_561,N_991);
nor U1683 (N_1683,N_1436,N_1102);
nand U1684 (N_1684,N_740,N_417);
or U1685 (N_1685,N_783,N_1367);
or U1686 (N_1686,N_224,N_556);
nor U1687 (N_1687,N_1069,N_1182);
and U1688 (N_1688,N_1465,N_370);
or U1689 (N_1689,N_1442,N_468);
nand U1690 (N_1690,N_657,N_1391);
nor U1691 (N_1691,N_1355,N_1457);
or U1692 (N_1692,N_683,N_307);
nor U1693 (N_1693,N_105,N_1227);
nor U1694 (N_1694,N_265,N_852);
nand U1695 (N_1695,N_85,N_801);
nor U1696 (N_1696,N_1183,N_1453);
nor U1697 (N_1697,N_1281,N_1086);
and U1698 (N_1698,N_1279,N_1202);
nand U1699 (N_1699,N_432,N_64);
and U1700 (N_1700,N_353,N_880);
nand U1701 (N_1701,N_472,N_1199);
nor U1702 (N_1702,N_24,N_547);
nand U1703 (N_1703,N_1317,N_721);
or U1704 (N_1704,N_1180,N_421);
or U1705 (N_1705,N_789,N_1447);
or U1706 (N_1706,N_677,N_1341);
and U1707 (N_1707,N_861,N_997);
nand U1708 (N_1708,N_27,N_1137);
or U1709 (N_1709,N_971,N_435);
nand U1710 (N_1710,N_213,N_383);
nand U1711 (N_1711,N_645,N_1116);
nor U1712 (N_1712,N_3,N_412);
nor U1713 (N_1713,N_1377,N_1362);
nand U1714 (N_1714,N_1080,N_606);
nand U1715 (N_1715,N_802,N_962);
and U1716 (N_1716,N_578,N_730);
nor U1717 (N_1717,N_753,N_47);
and U1718 (N_1718,N_815,N_78);
and U1719 (N_1719,N_294,N_117);
nand U1720 (N_1720,N_366,N_595);
xor U1721 (N_1721,N_992,N_386);
nor U1722 (N_1722,N_685,N_1068);
nand U1723 (N_1723,N_716,N_1096);
nand U1724 (N_1724,N_1033,N_43);
or U1725 (N_1725,N_936,N_167);
and U1726 (N_1726,N_176,N_614);
nor U1727 (N_1727,N_748,N_981);
or U1728 (N_1728,N_1405,N_993);
nor U1729 (N_1729,N_830,N_933);
nand U1730 (N_1730,N_1264,N_712);
nor U1731 (N_1731,N_434,N_622);
or U1732 (N_1732,N_894,N_1043);
and U1733 (N_1733,N_270,N_988);
nor U1734 (N_1734,N_1243,N_907);
or U1735 (N_1735,N_251,N_1370);
nor U1736 (N_1736,N_838,N_66);
nand U1737 (N_1737,N_241,N_12);
nand U1738 (N_1738,N_953,N_1455);
nand U1739 (N_1739,N_312,N_1016);
or U1740 (N_1740,N_980,N_1270);
or U1741 (N_1741,N_61,N_1486);
and U1742 (N_1742,N_1492,N_890);
nand U1743 (N_1743,N_943,N_456);
and U1744 (N_1744,N_1208,N_536);
or U1745 (N_1745,N_775,N_232);
or U1746 (N_1746,N_429,N_724);
and U1747 (N_1747,N_501,N_807);
nor U1748 (N_1748,N_1014,N_532);
or U1749 (N_1749,N_810,N_1191);
xnor U1750 (N_1750,N_1290,N_142);
and U1751 (N_1751,N_1276,N_275);
xnor U1752 (N_1752,N_28,N_336);
or U1753 (N_1753,N_1070,N_598);
nand U1754 (N_1754,N_1364,N_1361);
nor U1755 (N_1755,N_972,N_1301);
or U1756 (N_1756,N_414,N_711);
nand U1757 (N_1757,N_1474,N_218);
nand U1758 (N_1758,N_865,N_144);
nand U1759 (N_1759,N_515,N_570);
nor U1760 (N_1760,N_509,N_332);
and U1761 (N_1761,N_850,N_770);
nand U1762 (N_1762,N_328,N_497);
nand U1763 (N_1763,N_669,N_1064);
nor U1764 (N_1764,N_927,N_1162);
nor U1765 (N_1765,N_1328,N_1386);
and U1766 (N_1766,N_969,N_96);
or U1767 (N_1767,N_609,N_888);
or U1768 (N_1768,N_522,N_1216);
and U1769 (N_1769,N_168,N_1091);
or U1770 (N_1770,N_1302,N_425);
nand U1771 (N_1771,N_776,N_408);
and U1772 (N_1772,N_16,N_272);
or U1773 (N_1773,N_0,N_671);
nand U1774 (N_1774,N_284,N_192);
or U1775 (N_1775,N_700,N_1312);
and U1776 (N_1776,N_466,N_83);
or U1777 (N_1777,N_186,N_531);
nand U1778 (N_1778,N_196,N_1092);
nand U1779 (N_1779,N_323,N_396);
or U1780 (N_1780,N_1155,N_814);
nand U1781 (N_1781,N_787,N_116);
nor U1782 (N_1782,N_841,N_832);
nand U1783 (N_1783,N_640,N_1241);
or U1784 (N_1784,N_1347,N_1175);
nor U1785 (N_1785,N_610,N_420);
or U1786 (N_1786,N_940,N_486);
and U1787 (N_1787,N_1032,N_1150);
nand U1788 (N_1788,N_237,N_1428);
nand U1789 (N_1789,N_540,N_583);
or U1790 (N_1790,N_592,N_571);
nand U1791 (N_1791,N_1339,N_1057);
and U1792 (N_1792,N_438,N_175);
or U1793 (N_1793,N_1466,N_458);
nand U1794 (N_1794,N_715,N_668);
xnor U1795 (N_1795,N_793,N_1187);
nor U1796 (N_1796,N_277,N_1329);
and U1797 (N_1797,N_932,N_13);
nand U1798 (N_1798,N_63,N_1089);
nand U1799 (N_1799,N_604,N_152);
nand U1800 (N_1800,N_781,N_897);
and U1801 (N_1801,N_1117,N_611);
nand U1802 (N_1802,N_873,N_1);
nor U1803 (N_1803,N_856,N_10);
nor U1804 (N_1804,N_1022,N_519);
and U1805 (N_1805,N_254,N_209);
nor U1806 (N_1806,N_869,N_157);
nor U1807 (N_1807,N_1469,N_1261);
or U1808 (N_1808,N_1084,N_1072);
nor U1809 (N_1809,N_1220,N_461);
nor U1810 (N_1810,N_1097,N_431);
nand U1811 (N_1811,N_874,N_1498);
nand U1812 (N_1812,N_25,N_1018);
and U1813 (N_1813,N_151,N_231);
nor U1814 (N_1814,N_875,N_1062);
or U1815 (N_1815,N_1113,N_459);
nor U1816 (N_1816,N_1130,N_489);
and U1817 (N_1817,N_1303,N_706);
and U1818 (N_1818,N_911,N_314);
nor U1819 (N_1819,N_906,N_22);
nor U1820 (N_1820,N_697,N_661);
nand U1821 (N_1821,N_1394,N_406);
nand U1822 (N_1822,N_1222,N_276);
and U1823 (N_1823,N_1295,N_273);
nor U1824 (N_1824,N_1348,N_84);
or U1825 (N_1825,N_1473,N_1292);
nor U1826 (N_1826,N_1110,N_476);
or U1827 (N_1827,N_653,N_504);
and U1828 (N_1828,N_1001,N_964);
or U1829 (N_1829,N_1025,N_1082);
and U1830 (N_1830,N_297,N_394);
nor U1831 (N_1831,N_146,N_769);
or U1832 (N_1832,N_759,N_684);
or U1833 (N_1833,N_1354,N_1058);
nor U1834 (N_1834,N_1497,N_1315);
nor U1835 (N_1835,N_124,N_1353);
and U1836 (N_1836,N_120,N_1114);
and U1837 (N_1837,N_703,N_46);
nand U1838 (N_1838,N_1250,N_1415);
or U1839 (N_1839,N_291,N_138);
or U1840 (N_1840,N_1262,N_914);
or U1841 (N_1841,N_302,N_298);
or U1842 (N_1842,N_204,N_1471);
or U1843 (N_1843,N_487,N_887);
and U1844 (N_1844,N_290,N_153);
or U1845 (N_1845,N_512,N_523);
and U1846 (N_1846,N_313,N_100);
or U1847 (N_1847,N_1299,N_1456);
or U1848 (N_1848,N_375,N_1010);
or U1849 (N_1849,N_895,N_483);
and U1850 (N_1850,N_1313,N_682);
nand U1851 (N_1851,N_811,N_627);
and U1852 (N_1852,N_1425,N_961);
nand U1853 (N_1853,N_354,N_621);
or U1854 (N_1854,N_119,N_1271);
and U1855 (N_1855,N_1366,N_893);
or U1856 (N_1856,N_966,N_1209);
nor U1857 (N_1857,N_1314,N_868);
and U1858 (N_1858,N_123,N_941);
or U1859 (N_1859,N_791,N_1318);
or U1860 (N_1860,N_1152,N_876);
or U1861 (N_1861,N_1365,N_637);
or U1862 (N_1862,N_1106,N_263);
nand U1863 (N_1863,N_18,N_1462);
nand U1864 (N_1864,N_839,N_467);
nor U1865 (N_1865,N_199,N_862);
and U1866 (N_1866,N_970,N_771);
or U1867 (N_1867,N_920,N_289);
or U1868 (N_1868,N_1378,N_1310);
nand U1869 (N_1869,N_986,N_1372);
nor U1870 (N_1870,N_619,N_1192);
and U1871 (N_1871,N_939,N_825);
xor U1872 (N_1872,N_1105,N_924);
nor U1873 (N_1873,N_816,N_827);
nand U1874 (N_1874,N_87,N_587);
or U1875 (N_1875,N_1074,N_1401);
nor U1876 (N_1876,N_1344,N_1179);
nor U1877 (N_1877,N_351,N_1439);
nor U1878 (N_1878,N_798,N_296);
nor U1879 (N_1879,N_162,N_534);
and U1880 (N_1880,N_376,N_742);
and U1881 (N_1881,N_184,N_1280);
nor U1882 (N_1882,N_773,N_1412);
nand U1883 (N_1883,N_347,N_644);
and U1884 (N_1884,N_88,N_557);
and U1885 (N_1885,N_1149,N_245);
or U1886 (N_1886,N_32,N_1104);
nor U1887 (N_1887,N_745,N_804);
or U1888 (N_1888,N_710,N_1173);
nor U1889 (N_1889,N_879,N_1458);
or U1890 (N_1890,N_928,N_1024);
nand U1891 (N_1891,N_806,N_159);
nor U1892 (N_1892,N_246,N_1063);
or U1893 (N_1893,N_1249,N_9);
nor U1894 (N_1894,N_820,N_227);
or U1895 (N_1895,N_48,N_1195);
nand U1896 (N_1896,N_634,N_475);
nand U1897 (N_1897,N_958,N_720);
or U1898 (N_1898,N_687,N_1363);
nor U1899 (N_1899,N_1075,N_1163);
nor U1900 (N_1900,N_1283,N_1434);
or U1901 (N_1901,N_169,N_31);
nand U1902 (N_1902,N_563,N_1265);
nand U1903 (N_1903,N_580,N_490);
nor U1904 (N_1904,N_1196,N_401);
or U1905 (N_1905,N_1120,N_1332);
and U1906 (N_1906,N_1146,N_1481);
and U1907 (N_1907,N_1017,N_49);
nand U1908 (N_1908,N_678,N_125);
nor U1909 (N_1909,N_372,N_584);
and U1910 (N_1910,N_883,N_149);
nand U1911 (N_1911,N_664,N_1231);
or U1912 (N_1912,N_903,N_498);
and U1913 (N_1913,N_709,N_1052);
or U1914 (N_1914,N_238,N_658);
and U1915 (N_1915,N_1406,N_1099);
nor U1916 (N_1916,N_871,N_1011);
and U1917 (N_1917,N_550,N_325);
or U1918 (N_1918,N_660,N_975);
and U1919 (N_1919,N_114,N_995);
nor U1920 (N_1920,N_287,N_1269);
nor U1921 (N_1921,N_1490,N_1403);
or U1922 (N_1922,N_42,N_575);
and U1923 (N_1923,N_261,N_398);
and U1924 (N_1924,N_1322,N_474);
nor U1925 (N_1925,N_946,N_590);
nor U1926 (N_1926,N_469,N_799);
or U1927 (N_1927,N_746,N_562);
nor U1928 (N_1928,N_568,N_80);
or U1929 (N_1929,N_708,N_796);
and U1930 (N_1930,N_643,N_340);
xnor U1931 (N_1931,N_229,N_1273);
or U1932 (N_1932,N_1285,N_59);
nand U1933 (N_1933,N_403,N_916);
nor U1934 (N_1934,N_281,N_885);
and U1935 (N_1935,N_1007,N_378);
nor U1936 (N_1936,N_1291,N_926);
nor U1937 (N_1937,N_857,N_1021);
nor U1938 (N_1938,N_385,N_898);
nand U1939 (N_1939,N_1420,N_262);
or U1940 (N_1940,N_233,N_30);
xor U1941 (N_1941,N_670,N_756);
nand U1942 (N_1942,N_1138,N_705);
nand U1943 (N_1943,N_840,N_944);
nand U1944 (N_1944,N_155,N_207);
or U1945 (N_1945,N_1047,N_1330);
nor U1946 (N_1946,N_491,N_1441);
and U1947 (N_1947,N_923,N_533);
and U1948 (N_1948,N_1267,N_1178);
and U1949 (N_1949,N_482,N_918);
nor U1950 (N_1950,N_1212,N_274);
nand U1951 (N_1951,N_1193,N_686);
or U1952 (N_1952,N_166,N_1252);
nand U1953 (N_1953,N_794,N_543);
and U1954 (N_1954,N_1198,N_957);
and U1955 (N_1955,N_488,N_1454);
or U1956 (N_1956,N_1286,N_600);
and U1957 (N_1957,N_675,N_154);
and U1958 (N_1958,N_1340,N_267);
and U1959 (N_1959,N_623,N_565);
and U1960 (N_1960,N_553,N_4);
nor U1961 (N_1961,N_605,N_413);
nor U1962 (N_1962,N_1186,N_1224);
and U1963 (N_1963,N_1356,N_194);
or U1964 (N_1964,N_1384,N_761);
and U1965 (N_1965,N_546,N_722);
or U1966 (N_1966,N_1073,N_693);
or U1967 (N_1967,N_350,N_628);
nor U1968 (N_1968,N_457,N_150);
nor U1969 (N_1969,N_1321,N_430);
nor U1970 (N_1970,N_36,N_471);
nand U1971 (N_1971,N_593,N_74);
nor U1972 (N_1972,N_747,N_750);
and U1973 (N_1973,N_1373,N_230);
or U1974 (N_1974,N_1319,N_599);
and U1975 (N_1975,N_1030,N_701);
and U1976 (N_1976,N_228,N_1004);
nor U1977 (N_1977,N_343,N_785);
nand U1978 (N_1978,N_530,N_1351);
or U1979 (N_1979,N_455,N_344);
or U1980 (N_1980,N_1181,N_1357);
or U1981 (N_1981,N_650,N_1289);
nand U1982 (N_1982,N_1444,N_341);
or U1983 (N_1983,N_161,N_626);
nand U1984 (N_1984,N_514,N_1275);
or U1985 (N_1985,N_139,N_65);
nor U1986 (N_1986,N_1438,N_842);
or U1987 (N_1987,N_1185,N_925);
nor U1988 (N_1988,N_994,N_1095);
nand U1989 (N_1989,N_665,N_1061);
nand U1990 (N_1990,N_1326,N_989);
nor U1991 (N_1991,N_635,N_360);
nand U1992 (N_1992,N_1125,N_1067);
or U1993 (N_1993,N_129,N_591);
nand U1994 (N_1994,N_34,N_1006);
or U1995 (N_1995,N_1429,N_872);
nor U1996 (N_1996,N_102,N_1133);
nand U1997 (N_1997,N_179,N_978);
nand U1998 (N_1998,N_1055,N_1038);
nor U1999 (N_1999,N_463,N_596);
and U2000 (N_2000,N_44,N_503);
and U2001 (N_2001,N_535,N_1142);
nor U2002 (N_2002,N_200,N_1393);
xnor U2003 (N_2003,N_1343,N_444);
or U2004 (N_2004,N_674,N_1260);
or U2005 (N_2005,N_1480,N_1153);
or U2006 (N_2006,N_384,N_399);
and U2007 (N_2007,N_1168,N_777);
and U2008 (N_2008,N_891,N_945);
nor U2009 (N_2009,N_107,N_843);
nor U2010 (N_2010,N_726,N_930);
nor U2011 (N_2011,N_1049,N_259);
nand U2012 (N_2012,N_1451,N_1157);
and U2013 (N_2013,N_1255,N_440);
and U2014 (N_2014,N_624,N_506);
nor U2015 (N_2015,N_542,N_1232);
nand U2016 (N_2016,N_411,N_367);
nor U2017 (N_2017,N_1205,N_1496);
and U2018 (N_2018,N_377,N_821);
nor U2019 (N_2019,N_1375,N_779);
or U2020 (N_2020,N_1333,N_1076);
and U2021 (N_2021,N_1008,N_728);
or U2022 (N_2022,N_326,N_1397);
xor U2023 (N_2023,N_786,N_260);
and U2024 (N_2024,N_952,N_188);
or U2025 (N_2025,N_1031,N_140);
and U2026 (N_2026,N_510,N_464);
or U2027 (N_2027,N_1108,N_1392);
or U2028 (N_2028,N_266,N_1100);
or U2029 (N_2029,N_443,N_1005);
nand U2030 (N_2030,N_749,N_929);
nand U2031 (N_2031,N_1399,N_1111);
and U2032 (N_2032,N_1337,N_1054);
nor U2033 (N_2033,N_1127,N_646);
nor U2034 (N_2034,N_518,N_851);
or U2035 (N_2035,N_729,N_656);
or U2036 (N_2036,N_1144,N_723);
nand U2037 (N_2037,N_1094,N_51);
and U2038 (N_2038,N_160,N_1176);
and U2039 (N_2039,N_878,N_178);
nor U2040 (N_2040,N_40,N_1488);
nor U2041 (N_2041,N_834,N_433);
and U2042 (N_2042,N_613,N_243);
nand U2043 (N_2043,N_495,N_215);
or U2044 (N_2044,N_1126,N_426);
and U2045 (N_2045,N_985,N_636);
nor U2046 (N_2046,N_1334,N_951);
and U2047 (N_2047,N_846,N_191);
or U2048 (N_2048,N_649,N_1472);
nor U2049 (N_2049,N_240,N_612);
or U2050 (N_2050,N_303,N_1020);
nand U2051 (N_2051,N_214,N_539);
nand U2052 (N_2052,N_1060,N_1013);
nor U2053 (N_2053,N_280,N_892);
or U2054 (N_2054,N_422,N_135);
nor U2055 (N_2055,N_1410,N_714);
nand U2056 (N_2056,N_81,N_387);
nor U2057 (N_2057,N_1174,N_190);
nor U2058 (N_2058,N_1402,N_226);
and U2059 (N_2059,N_639,N_392);
nor U2060 (N_2060,N_21,N_1387);
nand U2061 (N_2061,N_1177,N_1132);
nor U2062 (N_2062,N_797,N_393);
or U2063 (N_2063,N_973,N_1327);
and U2064 (N_2064,N_625,N_110);
or U2065 (N_2065,N_424,N_305);
nand U2066 (N_2066,N_1234,N_279);
and U2067 (N_2067,N_829,N_1460);
nand U2068 (N_2068,N_1371,N_999);
and U2069 (N_2069,N_757,N_1044);
nand U2070 (N_2070,N_1476,N_288);
nand U2071 (N_2071,N_45,N_337);
or U2072 (N_2072,N_180,N_1421);
nor U2073 (N_2073,N_446,N_239);
or U2074 (N_2074,N_608,N_956);
or U2075 (N_2075,N_1172,N_648);
and U2076 (N_2076,N_147,N_1040);
and U2077 (N_2077,N_1230,N_256);
nand U2078 (N_2078,N_1342,N_108);
or U2079 (N_2079,N_938,N_662);
and U2080 (N_2080,N_780,N_505);
nand U2081 (N_2081,N_618,N_511);
or U2082 (N_2082,N_15,N_1298);
and U2083 (N_2083,N_1468,N_651);
xor U2084 (N_2084,N_1467,N_1483);
nor U2085 (N_2085,N_247,N_1085);
and U2086 (N_2086,N_1029,N_1418);
or U2087 (N_2087,N_1408,N_698);
nor U2088 (N_2088,N_854,N_1461);
xnor U2089 (N_2089,N_210,N_1268);
or U2090 (N_2090,N_1288,N_507);
or U2091 (N_2091,N_248,N_1045);
or U2092 (N_2092,N_1083,N_1090);
or U2093 (N_2093,N_62,N_115);
or U2094 (N_2094,N_130,N_242);
or U2095 (N_2095,N_768,N_1236);
or U2096 (N_2096,N_23,N_942);
nand U2097 (N_2097,N_1151,N_1160);
nor U2098 (N_2098,N_225,N_141);
or U2099 (N_2099,N_1207,N_69);
and U2100 (N_2100,N_1445,N_101);
and U2101 (N_2101,N_283,N_1056);
and U2102 (N_2102,N_921,N_1335);
nor U2103 (N_2103,N_1495,N_1316);
and U2104 (N_2104,N_1272,N_465);
nand U2105 (N_2105,N_349,N_1221);
or U2106 (N_2106,N_309,N_395);
or U2107 (N_2107,N_691,N_790);
nor U2108 (N_2108,N_133,N_947);
nand U2109 (N_2109,N_441,N_803);
xor U2110 (N_2110,N_1380,N_449);
or U2111 (N_2111,N_68,N_1246);
or U2112 (N_2112,N_585,N_345);
or U2113 (N_2113,N_282,N_26);
or U2114 (N_2114,N_689,N_1009);
and U2115 (N_2115,N_39,N_502);
or U2116 (N_2116,N_603,N_763);
nor U2117 (N_2117,N_881,N_837);
and U2118 (N_2118,N_365,N_327);
nand U2119 (N_2119,N_1304,N_407);
and U2120 (N_2120,N_1244,N_1287);
and U2121 (N_2121,N_1296,N_1059);
nand U2122 (N_2122,N_576,N_1088);
and U2123 (N_2123,N_902,N_1274);
or U2124 (N_2124,N_1431,N_732);
nor U2125 (N_2125,N_1475,N_767);
nor U2126 (N_2126,N_1470,N_77);
nand U2127 (N_2127,N_132,N_182);
or U2128 (N_2128,N_1124,N_363);
or U2129 (N_2129,N_1194,N_822);
nor U2130 (N_2130,N_500,N_752);
nand U2131 (N_2131,N_1002,N_17);
or U2132 (N_2132,N_1294,N_1430);
nor U2133 (N_2133,N_1201,N_1426);
nor U2134 (N_2134,N_1134,N_1041);
nor U2135 (N_2135,N_364,N_92);
or U2136 (N_2136,N_346,N_877);
or U2137 (N_2137,N_917,N_203);
and U2138 (N_2138,N_369,N_402);
and U2139 (N_2139,N_1433,N_442);
and U2140 (N_2140,N_772,N_187);
nor U2141 (N_2141,N_659,N_217);
and U2142 (N_2142,N_379,N_1482);
or U2143 (N_2143,N_470,N_1381);
nand U2144 (N_2144,N_1448,N_1251);
or U2145 (N_2145,N_301,N_148);
nor U2146 (N_2146,N_253,N_558);
nor U2147 (N_2147,N_602,N_1396);
and U2148 (N_2148,N_1165,N_690);
nor U2149 (N_2149,N_1463,N_268);
or U2150 (N_2150,N_1115,N_517);
nor U2151 (N_2151,N_597,N_1037);
nor U2152 (N_2152,N_884,N_50);
nand U2153 (N_2153,N_733,N_485);
nor U2154 (N_2154,N_1449,N_977);
nand U2155 (N_2155,N_1452,N_60);
nand U2156 (N_2156,N_380,N_1379);
nor U2157 (N_2157,N_1101,N_909);
nor U2158 (N_2158,N_824,N_744);
nand U2159 (N_2159,N_1051,N_795);
or U2160 (N_2160,N_454,N_436);
and U2161 (N_2161,N_67,N_1385);
nand U2162 (N_2162,N_1404,N_638);
and U2163 (N_2163,N_322,N_493);
nand U2164 (N_2164,N_1247,N_331);
and U2165 (N_2165,N_1218,N_630);
and U2166 (N_2166,N_1036,N_1464);
nand U2167 (N_2167,N_633,N_1346);
or U2168 (N_2168,N_577,N_672);
or U2169 (N_2169,N_308,N_189);
or U2170 (N_2170,N_1248,N_696);
or U2171 (N_2171,N_905,N_1485);
nor U2172 (N_2172,N_6,N_1156);
nor U2173 (N_2173,N_319,N_317);
or U2174 (N_2174,N_755,N_586);
or U2175 (N_2175,N_1306,N_478);
nor U2176 (N_2176,N_1053,N_1098);
nor U2177 (N_2177,N_158,N_410);
nor U2178 (N_2178,N_1170,N_397);
and U2179 (N_2179,N_963,N_1237);
or U2180 (N_2180,N_70,N_1324);
and U2181 (N_2181,N_912,N_1359);
nand U2182 (N_2182,N_955,N_1148);
and U2183 (N_2183,N_181,N_741);
nand U2184 (N_2184,N_818,N_702);
xor U2185 (N_2185,N_731,N_800);
nor U2186 (N_2186,N_1282,N_954);
nor U2187 (N_2187,N_828,N_1499);
nand U2188 (N_2188,N_1278,N_1238);
or U2189 (N_2189,N_784,N_1477);
nor U2190 (N_2190,N_934,N_699);
and U2191 (N_2191,N_1254,N_935);
nor U2192 (N_2192,N_900,N_526);
nand U2193 (N_2193,N_632,N_177);
nand U2194 (N_2194,N_765,N_864);
or U2195 (N_2195,N_1078,N_453);
nor U2196 (N_2196,N_654,N_1103);
and U2197 (N_2197,N_171,N_1147);
nor U2198 (N_2198,N_195,N_164);
xor U2199 (N_2199,N_1206,N_1012);
nand U2200 (N_2200,N_1479,N_859);
and U2201 (N_2201,N_56,N_134);
or U2202 (N_2202,N_329,N_1400);
nand U2203 (N_2203,N_990,N_1210);
and U2204 (N_2204,N_1369,N_1376);
nor U2205 (N_2205,N_817,N_1493);
or U2206 (N_2206,N_292,N_528);
and U2207 (N_2207,N_704,N_1427);
nand U2208 (N_2208,N_415,N_7);
or U2209 (N_2209,N_1167,N_499);
nor U2210 (N_2210,N_416,N_601);
or U2211 (N_2211,N_727,N_170);
nand U2212 (N_2212,N_127,N_1440);
or U2213 (N_2213,N_1118,N_1320);
nor U2214 (N_2214,N_1459,N_462);
nand U2215 (N_2215,N_222,N_109);
and U2216 (N_2216,N_560,N_1028);
and U2217 (N_2217,N_965,N_1164);
and U2218 (N_2218,N_1046,N_300);
or U2219 (N_2219,N_54,N_1253);
nand U2220 (N_2220,N_357,N_1395);
or U2221 (N_2221,N_212,N_713);
nor U2222 (N_2222,N_1035,N_1360);
or U2223 (N_2223,N_315,N_1019);
and U2224 (N_2224,N_1079,N_1158);
nand U2225 (N_2225,N_1225,N_1215);
and U2226 (N_2226,N_1107,N_886);
and U2227 (N_2227,N_368,N_582);
nor U2228 (N_2228,N_549,N_641);
nand U2229 (N_2229,N_1263,N_72);
and U2230 (N_2230,N_681,N_131);
nand U2231 (N_2231,N_1416,N_782);
nand U2232 (N_2232,N_201,N_122);
nor U2233 (N_2233,N_1235,N_845);
nor U2234 (N_2234,N_569,N_1121);
or U2235 (N_2235,N_1023,N_1345);
and U2236 (N_2236,N_707,N_960);
and U2237 (N_2237,N_1122,N_423);
nand U2238 (N_2238,N_320,N_382);
and U2239 (N_2239,N_93,N_858);
xor U2240 (N_2240,N_404,N_1338);
and U2241 (N_2241,N_1050,N_1494);
and U2242 (N_2242,N_1390,N_235);
or U2243 (N_2243,N_339,N_663);
or U2244 (N_2244,N_1309,N_185);
and U2245 (N_2245,N_236,N_448);
or U2246 (N_2246,N_695,N_1389);
or U2247 (N_2247,N_249,N_1213);
or U2248 (N_2248,N_541,N_976);
or U2249 (N_2249,N_405,N_1297);
nand U2250 (N_2250,N_696,N_581);
nor U2251 (N_2251,N_1125,N_1073);
or U2252 (N_2252,N_1160,N_1003);
and U2253 (N_2253,N_208,N_1022);
nand U2254 (N_2254,N_1377,N_84);
nor U2255 (N_2255,N_320,N_285);
nor U2256 (N_2256,N_1126,N_996);
or U2257 (N_2257,N_892,N_793);
and U2258 (N_2258,N_1127,N_1272);
nor U2259 (N_2259,N_1157,N_1035);
nand U2260 (N_2260,N_1048,N_285);
nand U2261 (N_2261,N_851,N_1417);
nor U2262 (N_2262,N_1494,N_856);
and U2263 (N_2263,N_1313,N_350);
and U2264 (N_2264,N_979,N_1056);
and U2265 (N_2265,N_453,N_118);
nor U2266 (N_2266,N_679,N_186);
nor U2267 (N_2267,N_21,N_180);
xnor U2268 (N_2268,N_1427,N_773);
and U2269 (N_2269,N_1075,N_588);
and U2270 (N_2270,N_255,N_609);
or U2271 (N_2271,N_166,N_1320);
nand U2272 (N_2272,N_744,N_569);
or U2273 (N_2273,N_1368,N_74);
nand U2274 (N_2274,N_460,N_34);
nor U2275 (N_2275,N_822,N_498);
or U2276 (N_2276,N_646,N_38);
and U2277 (N_2277,N_796,N_223);
nand U2278 (N_2278,N_483,N_519);
nand U2279 (N_2279,N_1027,N_1308);
and U2280 (N_2280,N_966,N_1073);
and U2281 (N_2281,N_1016,N_820);
or U2282 (N_2282,N_1124,N_1458);
or U2283 (N_2283,N_1469,N_754);
nor U2284 (N_2284,N_819,N_1470);
or U2285 (N_2285,N_704,N_794);
nor U2286 (N_2286,N_47,N_554);
and U2287 (N_2287,N_895,N_1064);
and U2288 (N_2288,N_396,N_553);
nor U2289 (N_2289,N_655,N_95);
and U2290 (N_2290,N_1291,N_23);
nand U2291 (N_2291,N_1442,N_1329);
or U2292 (N_2292,N_907,N_1270);
nand U2293 (N_2293,N_386,N_836);
or U2294 (N_2294,N_847,N_65);
nor U2295 (N_2295,N_1393,N_1053);
nand U2296 (N_2296,N_486,N_1363);
nand U2297 (N_2297,N_591,N_233);
or U2298 (N_2298,N_341,N_652);
nor U2299 (N_2299,N_1491,N_474);
nand U2300 (N_2300,N_843,N_680);
and U2301 (N_2301,N_84,N_83);
nor U2302 (N_2302,N_470,N_620);
nand U2303 (N_2303,N_537,N_533);
nor U2304 (N_2304,N_758,N_672);
and U2305 (N_2305,N_406,N_403);
nor U2306 (N_2306,N_673,N_1337);
nor U2307 (N_2307,N_1065,N_1062);
and U2308 (N_2308,N_1156,N_1137);
or U2309 (N_2309,N_1395,N_1166);
nor U2310 (N_2310,N_159,N_912);
or U2311 (N_2311,N_992,N_1306);
or U2312 (N_2312,N_1237,N_1252);
nand U2313 (N_2313,N_878,N_458);
and U2314 (N_2314,N_1078,N_846);
and U2315 (N_2315,N_822,N_1472);
or U2316 (N_2316,N_561,N_341);
and U2317 (N_2317,N_792,N_144);
or U2318 (N_2318,N_323,N_583);
or U2319 (N_2319,N_2,N_1153);
nand U2320 (N_2320,N_828,N_894);
and U2321 (N_2321,N_1334,N_1319);
nor U2322 (N_2322,N_1298,N_1382);
nor U2323 (N_2323,N_480,N_1147);
nand U2324 (N_2324,N_936,N_1208);
nor U2325 (N_2325,N_1362,N_25);
nand U2326 (N_2326,N_690,N_852);
or U2327 (N_2327,N_22,N_778);
or U2328 (N_2328,N_1159,N_304);
nor U2329 (N_2329,N_784,N_837);
and U2330 (N_2330,N_118,N_355);
nor U2331 (N_2331,N_1200,N_995);
nand U2332 (N_2332,N_1223,N_44);
nand U2333 (N_2333,N_1290,N_472);
nand U2334 (N_2334,N_1145,N_1142);
nand U2335 (N_2335,N_555,N_1246);
nand U2336 (N_2336,N_960,N_1301);
or U2337 (N_2337,N_952,N_1123);
or U2338 (N_2338,N_743,N_710);
nor U2339 (N_2339,N_73,N_852);
and U2340 (N_2340,N_125,N_165);
nor U2341 (N_2341,N_567,N_994);
nor U2342 (N_2342,N_1040,N_729);
nand U2343 (N_2343,N_579,N_1040);
nor U2344 (N_2344,N_267,N_1296);
or U2345 (N_2345,N_719,N_600);
or U2346 (N_2346,N_707,N_664);
or U2347 (N_2347,N_1330,N_141);
and U2348 (N_2348,N_815,N_814);
nand U2349 (N_2349,N_1403,N_551);
nor U2350 (N_2350,N_573,N_465);
or U2351 (N_2351,N_1372,N_863);
nor U2352 (N_2352,N_364,N_367);
nand U2353 (N_2353,N_1,N_314);
nand U2354 (N_2354,N_1080,N_870);
nand U2355 (N_2355,N_56,N_1248);
or U2356 (N_2356,N_1157,N_1011);
nor U2357 (N_2357,N_1203,N_404);
or U2358 (N_2358,N_166,N_269);
nor U2359 (N_2359,N_1296,N_1078);
nor U2360 (N_2360,N_548,N_652);
nor U2361 (N_2361,N_1383,N_742);
nor U2362 (N_2362,N_1456,N_741);
or U2363 (N_2363,N_672,N_1017);
or U2364 (N_2364,N_138,N_1348);
and U2365 (N_2365,N_913,N_498);
and U2366 (N_2366,N_634,N_117);
nor U2367 (N_2367,N_120,N_330);
and U2368 (N_2368,N_203,N_12);
or U2369 (N_2369,N_427,N_282);
and U2370 (N_2370,N_1457,N_1026);
or U2371 (N_2371,N_952,N_1061);
nand U2372 (N_2372,N_1267,N_363);
and U2373 (N_2373,N_1353,N_643);
nand U2374 (N_2374,N_1423,N_949);
nand U2375 (N_2375,N_1100,N_982);
nor U2376 (N_2376,N_736,N_605);
or U2377 (N_2377,N_224,N_429);
nand U2378 (N_2378,N_1427,N_486);
and U2379 (N_2379,N_86,N_721);
and U2380 (N_2380,N_975,N_1465);
or U2381 (N_2381,N_1131,N_29);
and U2382 (N_2382,N_154,N_1356);
nand U2383 (N_2383,N_616,N_1095);
and U2384 (N_2384,N_413,N_356);
nand U2385 (N_2385,N_625,N_1183);
and U2386 (N_2386,N_1018,N_505);
or U2387 (N_2387,N_1227,N_383);
nor U2388 (N_2388,N_512,N_1481);
nor U2389 (N_2389,N_808,N_1379);
and U2390 (N_2390,N_1146,N_1483);
nor U2391 (N_2391,N_768,N_1070);
or U2392 (N_2392,N_428,N_1253);
and U2393 (N_2393,N_1400,N_526);
or U2394 (N_2394,N_557,N_732);
nand U2395 (N_2395,N_1258,N_1166);
nand U2396 (N_2396,N_991,N_604);
nand U2397 (N_2397,N_105,N_534);
and U2398 (N_2398,N_532,N_739);
and U2399 (N_2399,N_1203,N_1347);
nor U2400 (N_2400,N_1011,N_260);
or U2401 (N_2401,N_2,N_1087);
and U2402 (N_2402,N_899,N_338);
or U2403 (N_2403,N_150,N_1178);
or U2404 (N_2404,N_1290,N_167);
or U2405 (N_2405,N_475,N_1097);
nand U2406 (N_2406,N_24,N_235);
nor U2407 (N_2407,N_1111,N_962);
nor U2408 (N_2408,N_1151,N_1489);
and U2409 (N_2409,N_340,N_480);
nand U2410 (N_2410,N_1168,N_778);
nor U2411 (N_2411,N_798,N_126);
and U2412 (N_2412,N_1181,N_952);
nor U2413 (N_2413,N_640,N_519);
nand U2414 (N_2414,N_1248,N_136);
or U2415 (N_2415,N_1471,N_298);
nor U2416 (N_2416,N_283,N_181);
nand U2417 (N_2417,N_1352,N_767);
or U2418 (N_2418,N_83,N_1177);
nand U2419 (N_2419,N_1268,N_485);
and U2420 (N_2420,N_1394,N_708);
or U2421 (N_2421,N_901,N_707);
nor U2422 (N_2422,N_1,N_1080);
xnor U2423 (N_2423,N_1434,N_228);
or U2424 (N_2424,N_25,N_1495);
and U2425 (N_2425,N_269,N_263);
nor U2426 (N_2426,N_1030,N_1284);
or U2427 (N_2427,N_1395,N_1319);
xor U2428 (N_2428,N_1348,N_265);
and U2429 (N_2429,N_616,N_1444);
nor U2430 (N_2430,N_1456,N_1367);
nand U2431 (N_2431,N_1485,N_1490);
or U2432 (N_2432,N_1196,N_444);
and U2433 (N_2433,N_776,N_505);
nor U2434 (N_2434,N_151,N_641);
nor U2435 (N_2435,N_621,N_1410);
and U2436 (N_2436,N_420,N_283);
nor U2437 (N_2437,N_158,N_1156);
nor U2438 (N_2438,N_670,N_416);
nor U2439 (N_2439,N_1298,N_788);
nor U2440 (N_2440,N_1318,N_952);
nor U2441 (N_2441,N_1080,N_553);
nor U2442 (N_2442,N_322,N_1055);
nor U2443 (N_2443,N_568,N_330);
or U2444 (N_2444,N_509,N_1301);
nor U2445 (N_2445,N_570,N_622);
and U2446 (N_2446,N_928,N_789);
nand U2447 (N_2447,N_143,N_494);
or U2448 (N_2448,N_1414,N_44);
or U2449 (N_2449,N_1418,N_1376);
nand U2450 (N_2450,N_328,N_909);
nor U2451 (N_2451,N_201,N_1148);
nand U2452 (N_2452,N_1426,N_311);
nor U2453 (N_2453,N_764,N_788);
nand U2454 (N_2454,N_988,N_1414);
or U2455 (N_2455,N_189,N_1141);
or U2456 (N_2456,N_647,N_1385);
and U2457 (N_2457,N_761,N_506);
or U2458 (N_2458,N_1112,N_848);
nor U2459 (N_2459,N_1152,N_1088);
nand U2460 (N_2460,N_408,N_407);
and U2461 (N_2461,N_411,N_124);
and U2462 (N_2462,N_809,N_1099);
nor U2463 (N_2463,N_967,N_1009);
and U2464 (N_2464,N_101,N_875);
and U2465 (N_2465,N_334,N_675);
and U2466 (N_2466,N_1042,N_178);
nor U2467 (N_2467,N_1036,N_45);
and U2468 (N_2468,N_1372,N_883);
and U2469 (N_2469,N_187,N_1220);
and U2470 (N_2470,N_1091,N_1071);
or U2471 (N_2471,N_127,N_823);
nor U2472 (N_2472,N_1319,N_866);
nor U2473 (N_2473,N_121,N_1138);
and U2474 (N_2474,N_1409,N_189);
and U2475 (N_2475,N_1379,N_1002);
nand U2476 (N_2476,N_321,N_655);
nor U2477 (N_2477,N_1316,N_174);
or U2478 (N_2478,N_1355,N_584);
nand U2479 (N_2479,N_838,N_810);
and U2480 (N_2480,N_1487,N_1173);
or U2481 (N_2481,N_573,N_467);
nand U2482 (N_2482,N_1296,N_1377);
nand U2483 (N_2483,N_1307,N_1172);
nand U2484 (N_2484,N_341,N_1113);
xnor U2485 (N_2485,N_236,N_1106);
nand U2486 (N_2486,N_312,N_474);
nor U2487 (N_2487,N_1176,N_691);
and U2488 (N_2488,N_817,N_346);
or U2489 (N_2489,N_264,N_293);
nand U2490 (N_2490,N_1452,N_474);
and U2491 (N_2491,N_1160,N_1433);
or U2492 (N_2492,N_223,N_180);
nor U2493 (N_2493,N_600,N_451);
or U2494 (N_2494,N_1037,N_110);
and U2495 (N_2495,N_867,N_1271);
nor U2496 (N_2496,N_726,N_331);
or U2497 (N_2497,N_1144,N_220);
and U2498 (N_2498,N_175,N_1457);
nand U2499 (N_2499,N_86,N_872);
or U2500 (N_2500,N_994,N_127);
and U2501 (N_2501,N_730,N_625);
and U2502 (N_2502,N_930,N_1485);
and U2503 (N_2503,N_1248,N_401);
or U2504 (N_2504,N_892,N_858);
or U2505 (N_2505,N_1478,N_1169);
and U2506 (N_2506,N_205,N_1136);
or U2507 (N_2507,N_770,N_627);
or U2508 (N_2508,N_1228,N_829);
nand U2509 (N_2509,N_574,N_1411);
nand U2510 (N_2510,N_44,N_822);
and U2511 (N_2511,N_26,N_580);
nand U2512 (N_2512,N_901,N_499);
and U2513 (N_2513,N_1092,N_1196);
and U2514 (N_2514,N_244,N_1281);
or U2515 (N_2515,N_214,N_592);
nand U2516 (N_2516,N_948,N_156);
and U2517 (N_2517,N_483,N_687);
nand U2518 (N_2518,N_261,N_1269);
nor U2519 (N_2519,N_2,N_1204);
nand U2520 (N_2520,N_491,N_1234);
or U2521 (N_2521,N_1388,N_1468);
or U2522 (N_2522,N_1044,N_275);
or U2523 (N_2523,N_1334,N_773);
and U2524 (N_2524,N_323,N_60);
nor U2525 (N_2525,N_854,N_554);
and U2526 (N_2526,N_862,N_153);
or U2527 (N_2527,N_149,N_393);
nand U2528 (N_2528,N_90,N_69);
nand U2529 (N_2529,N_364,N_1130);
or U2530 (N_2530,N_1217,N_194);
nand U2531 (N_2531,N_27,N_230);
nor U2532 (N_2532,N_1202,N_946);
nand U2533 (N_2533,N_380,N_1366);
nand U2534 (N_2534,N_327,N_1023);
or U2535 (N_2535,N_293,N_272);
nand U2536 (N_2536,N_481,N_1303);
nor U2537 (N_2537,N_1141,N_1067);
or U2538 (N_2538,N_84,N_1283);
nor U2539 (N_2539,N_32,N_65);
or U2540 (N_2540,N_294,N_1331);
nand U2541 (N_2541,N_1367,N_366);
nor U2542 (N_2542,N_518,N_1091);
or U2543 (N_2543,N_1449,N_530);
nor U2544 (N_2544,N_1143,N_671);
nand U2545 (N_2545,N_1177,N_1032);
nand U2546 (N_2546,N_515,N_1080);
and U2547 (N_2547,N_1046,N_337);
nor U2548 (N_2548,N_1440,N_9);
or U2549 (N_2549,N_123,N_839);
or U2550 (N_2550,N_1352,N_948);
or U2551 (N_2551,N_1349,N_660);
and U2552 (N_2552,N_42,N_547);
or U2553 (N_2553,N_523,N_7);
nand U2554 (N_2554,N_883,N_619);
nand U2555 (N_2555,N_677,N_437);
or U2556 (N_2556,N_10,N_203);
nand U2557 (N_2557,N_1089,N_105);
and U2558 (N_2558,N_794,N_743);
nand U2559 (N_2559,N_166,N_790);
and U2560 (N_2560,N_884,N_1294);
and U2561 (N_2561,N_227,N_271);
nor U2562 (N_2562,N_1268,N_1445);
nor U2563 (N_2563,N_259,N_1231);
and U2564 (N_2564,N_1468,N_918);
or U2565 (N_2565,N_1290,N_492);
nor U2566 (N_2566,N_1408,N_811);
nand U2567 (N_2567,N_927,N_1337);
nor U2568 (N_2568,N_317,N_1495);
nand U2569 (N_2569,N_1079,N_454);
and U2570 (N_2570,N_1257,N_228);
nand U2571 (N_2571,N_1247,N_1283);
nor U2572 (N_2572,N_419,N_438);
nand U2573 (N_2573,N_1106,N_279);
or U2574 (N_2574,N_289,N_906);
and U2575 (N_2575,N_1205,N_643);
nand U2576 (N_2576,N_1025,N_441);
nor U2577 (N_2577,N_1278,N_509);
or U2578 (N_2578,N_1498,N_101);
and U2579 (N_2579,N_363,N_422);
nand U2580 (N_2580,N_1420,N_131);
or U2581 (N_2581,N_1114,N_515);
and U2582 (N_2582,N_825,N_1377);
nor U2583 (N_2583,N_60,N_1298);
nor U2584 (N_2584,N_1255,N_307);
or U2585 (N_2585,N_170,N_237);
nor U2586 (N_2586,N_967,N_88);
nand U2587 (N_2587,N_864,N_1337);
and U2588 (N_2588,N_647,N_904);
or U2589 (N_2589,N_49,N_628);
and U2590 (N_2590,N_581,N_1136);
nand U2591 (N_2591,N_1420,N_43);
or U2592 (N_2592,N_969,N_630);
or U2593 (N_2593,N_424,N_94);
or U2594 (N_2594,N_1179,N_1319);
nor U2595 (N_2595,N_1232,N_688);
and U2596 (N_2596,N_99,N_202);
nand U2597 (N_2597,N_302,N_1462);
or U2598 (N_2598,N_1234,N_1211);
nand U2599 (N_2599,N_545,N_873);
nor U2600 (N_2600,N_1173,N_1021);
nor U2601 (N_2601,N_8,N_1354);
and U2602 (N_2602,N_587,N_896);
and U2603 (N_2603,N_1380,N_278);
or U2604 (N_2604,N_1090,N_1238);
or U2605 (N_2605,N_1375,N_830);
nand U2606 (N_2606,N_681,N_474);
nor U2607 (N_2607,N_130,N_75);
and U2608 (N_2608,N_762,N_913);
nor U2609 (N_2609,N_963,N_547);
or U2610 (N_2610,N_349,N_710);
nor U2611 (N_2611,N_1432,N_785);
nor U2612 (N_2612,N_1287,N_357);
and U2613 (N_2613,N_1157,N_564);
xor U2614 (N_2614,N_548,N_1188);
nor U2615 (N_2615,N_999,N_961);
nor U2616 (N_2616,N_1239,N_451);
and U2617 (N_2617,N_87,N_1113);
nor U2618 (N_2618,N_827,N_1461);
nor U2619 (N_2619,N_501,N_84);
and U2620 (N_2620,N_361,N_481);
or U2621 (N_2621,N_1194,N_201);
nor U2622 (N_2622,N_417,N_1492);
or U2623 (N_2623,N_1329,N_1494);
and U2624 (N_2624,N_1163,N_1030);
and U2625 (N_2625,N_788,N_22);
and U2626 (N_2626,N_39,N_1378);
nor U2627 (N_2627,N_925,N_404);
and U2628 (N_2628,N_249,N_411);
nor U2629 (N_2629,N_1275,N_587);
or U2630 (N_2630,N_880,N_150);
nor U2631 (N_2631,N_590,N_93);
nor U2632 (N_2632,N_1018,N_345);
and U2633 (N_2633,N_300,N_1270);
and U2634 (N_2634,N_1484,N_938);
nor U2635 (N_2635,N_1471,N_997);
nand U2636 (N_2636,N_510,N_1344);
nor U2637 (N_2637,N_1415,N_1247);
nand U2638 (N_2638,N_919,N_1291);
nor U2639 (N_2639,N_1158,N_476);
nor U2640 (N_2640,N_4,N_634);
and U2641 (N_2641,N_436,N_887);
and U2642 (N_2642,N_187,N_192);
nor U2643 (N_2643,N_470,N_736);
nand U2644 (N_2644,N_1389,N_111);
or U2645 (N_2645,N_803,N_615);
or U2646 (N_2646,N_1081,N_959);
nor U2647 (N_2647,N_957,N_288);
nor U2648 (N_2648,N_970,N_334);
nor U2649 (N_2649,N_886,N_884);
or U2650 (N_2650,N_457,N_1375);
or U2651 (N_2651,N_819,N_929);
nor U2652 (N_2652,N_1270,N_551);
nand U2653 (N_2653,N_543,N_564);
nor U2654 (N_2654,N_718,N_1292);
or U2655 (N_2655,N_1406,N_1261);
or U2656 (N_2656,N_1318,N_383);
and U2657 (N_2657,N_1388,N_176);
nor U2658 (N_2658,N_177,N_1492);
nor U2659 (N_2659,N_1295,N_572);
nand U2660 (N_2660,N_1233,N_567);
and U2661 (N_2661,N_683,N_534);
and U2662 (N_2662,N_248,N_514);
or U2663 (N_2663,N_151,N_97);
and U2664 (N_2664,N_1318,N_481);
nor U2665 (N_2665,N_1185,N_1043);
or U2666 (N_2666,N_1294,N_1375);
or U2667 (N_2667,N_91,N_281);
nor U2668 (N_2668,N_1237,N_791);
nor U2669 (N_2669,N_1175,N_940);
or U2670 (N_2670,N_583,N_1092);
and U2671 (N_2671,N_1200,N_586);
and U2672 (N_2672,N_92,N_471);
nand U2673 (N_2673,N_448,N_452);
nand U2674 (N_2674,N_414,N_598);
and U2675 (N_2675,N_622,N_935);
nand U2676 (N_2676,N_618,N_1376);
nand U2677 (N_2677,N_136,N_216);
or U2678 (N_2678,N_411,N_219);
nor U2679 (N_2679,N_32,N_119);
or U2680 (N_2680,N_753,N_1141);
nand U2681 (N_2681,N_458,N_1467);
nor U2682 (N_2682,N_61,N_752);
or U2683 (N_2683,N_778,N_1046);
nand U2684 (N_2684,N_388,N_1079);
and U2685 (N_2685,N_494,N_315);
and U2686 (N_2686,N_590,N_699);
and U2687 (N_2687,N_75,N_544);
or U2688 (N_2688,N_498,N_552);
or U2689 (N_2689,N_1156,N_1403);
and U2690 (N_2690,N_548,N_464);
nand U2691 (N_2691,N_1289,N_439);
and U2692 (N_2692,N_680,N_826);
nand U2693 (N_2693,N_668,N_318);
nand U2694 (N_2694,N_558,N_86);
nand U2695 (N_2695,N_435,N_86);
or U2696 (N_2696,N_859,N_629);
or U2697 (N_2697,N_568,N_222);
or U2698 (N_2698,N_1187,N_1358);
nor U2699 (N_2699,N_684,N_633);
and U2700 (N_2700,N_583,N_1004);
nand U2701 (N_2701,N_1492,N_1240);
nor U2702 (N_2702,N_1354,N_1113);
and U2703 (N_2703,N_1157,N_800);
and U2704 (N_2704,N_325,N_779);
nor U2705 (N_2705,N_913,N_301);
nand U2706 (N_2706,N_1058,N_787);
or U2707 (N_2707,N_565,N_567);
and U2708 (N_2708,N_711,N_1400);
nand U2709 (N_2709,N_1107,N_373);
and U2710 (N_2710,N_1001,N_1435);
nand U2711 (N_2711,N_757,N_1305);
nor U2712 (N_2712,N_195,N_98);
and U2713 (N_2713,N_590,N_1290);
nand U2714 (N_2714,N_1064,N_953);
nor U2715 (N_2715,N_1053,N_539);
and U2716 (N_2716,N_806,N_811);
nor U2717 (N_2717,N_1071,N_281);
and U2718 (N_2718,N_1066,N_253);
and U2719 (N_2719,N_1100,N_764);
nor U2720 (N_2720,N_363,N_1397);
nor U2721 (N_2721,N_1294,N_18);
or U2722 (N_2722,N_305,N_804);
or U2723 (N_2723,N_367,N_77);
and U2724 (N_2724,N_1189,N_1485);
nor U2725 (N_2725,N_1254,N_1019);
nor U2726 (N_2726,N_1296,N_1430);
nor U2727 (N_2727,N_1200,N_102);
or U2728 (N_2728,N_815,N_288);
nand U2729 (N_2729,N_1281,N_346);
nand U2730 (N_2730,N_1320,N_611);
nor U2731 (N_2731,N_709,N_180);
or U2732 (N_2732,N_1131,N_1417);
or U2733 (N_2733,N_1465,N_652);
and U2734 (N_2734,N_1187,N_874);
or U2735 (N_2735,N_1313,N_633);
nor U2736 (N_2736,N_1314,N_60);
nand U2737 (N_2737,N_1148,N_874);
nand U2738 (N_2738,N_1379,N_970);
nor U2739 (N_2739,N_1143,N_435);
nor U2740 (N_2740,N_266,N_776);
nor U2741 (N_2741,N_1256,N_1217);
and U2742 (N_2742,N_1158,N_883);
nor U2743 (N_2743,N_538,N_784);
and U2744 (N_2744,N_814,N_1499);
nor U2745 (N_2745,N_801,N_637);
nand U2746 (N_2746,N_884,N_725);
or U2747 (N_2747,N_155,N_759);
nor U2748 (N_2748,N_800,N_644);
nand U2749 (N_2749,N_473,N_607);
nand U2750 (N_2750,N_749,N_33);
nor U2751 (N_2751,N_1234,N_678);
nand U2752 (N_2752,N_396,N_1475);
nor U2753 (N_2753,N_866,N_1226);
nand U2754 (N_2754,N_1447,N_951);
and U2755 (N_2755,N_1471,N_1141);
and U2756 (N_2756,N_5,N_626);
and U2757 (N_2757,N_1487,N_400);
or U2758 (N_2758,N_375,N_624);
nand U2759 (N_2759,N_706,N_1120);
or U2760 (N_2760,N_1358,N_1019);
nand U2761 (N_2761,N_1199,N_568);
nor U2762 (N_2762,N_694,N_836);
or U2763 (N_2763,N_571,N_610);
xnor U2764 (N_2764,N_882,N_264);
nand U2765 (N_2765,N_1378,N_933);
or U2766 (N_2766,N_622,N_1451);
nand U2767 (N_2767,N_686,N_92);
nand U2768 (N_2768,N_1120,N_206);
nand U2769 (N_2769,N_240,N_1062);
nand U2770 (N_2770,N_915,N_416);
nor U2771 (N_2771,N_1382,N_220);
nor U2772 (N_2772,N_612,N_337);
or U2773 (N_2773,N_1357,N_226);
nand U2774 (N_2774,N_1114,N_376);
or U2775 (N_2775,N_481,N_678);
nor U2776 (N_2776,N_632,N_293);
and U2777 (N_2777,N_356,N_399);
or U2778 (N_2778,N_744,N_1410);
or U2779 (N_2779,N_159,N_1449);
or U2780 (N_2780,N_205,N_1186);
nor U2781 (N_2781,N_144,N_1337);
or U2782 (N_2782,N_855,N_369);
or U2783 (N_2783,N_375,N_931);
and U2784 (N_2784,N_1016,N_365);
or U2785 (N_2785,N_1260,N_67);
and U2786 (N_2786,N_1342,N_1086);
nor U2787 (N_2787,N_605,N_1457);
or U2788 (N_2788,N_1020,N_563);
or U2789 (N_2789,N_43,N_1070);
or U2790 (N_2790,N_1157,N_1400);
and U2791 (N_2791,N_4,N_276);
and U2792 (N_2792,N_807,N_1480);
nor U2793 (N_2793,N_1040,N_698);
nand U2794 (N_2794,N_440,N_553);
or U2795 (N_2795,N_52,N_830);
nand U2796 (N_2796,N_352,N_974);
and U2797 (N_2797,N_225,N_928);
or U2798 (N_2798,N_1311,N_573);
nand U2799 (N_2799,N_868,N_778);
nor U2800 (N_2800,N_645,N_1192);
nor U2801 (N_2801,N_1470,N_1357);
nor U2802 (N_2802,N_32,N_99);
and U2803 (N_2803,N_1146,N_1055);
nand U2804 (N_2804,N_318,N_1279);
and U2805 (N_2805,N_134,N_114);
or U2806 (N_2806,N_891,N_631);
nand U2807 (N_2807,N_700,N_265);
nand U2808 (N_2808,N_1065,N_801);
nand U2809 (N_2809,N_85,N_968);
nor U2810 (N_2810,N_438,N_268);
nor U2811 (N_2811,N_1266,N_1267);
or U2812 (N_2812,N_130,N_795);
nand U2813 (N_2813,N_67,N_899);
and U2814 (N_2814,N_1458,N_425);
or U2815 (N_2815,N_141,N_1407);
and U2816 (N_2816,N_214,N_429);
or U2817 (N_2817,N_0,N_902);
nor U2818 (N_2818,N_677,N_368);
xnor U2819 (N_2819,N_1033,N_1208);
nand U2820 (N_2820,N_570,N_1497);
or U2821 (N_2821,N_879,N_13);
nand U2822 (N_2822,N_1259,N_1427);
or U2823 (N_2823,N_347,N_231);
nand U2824 (N_2824,N_1193,N_87);
nand U2825 (N_2825,N_915,N_370);
or U2826 (N_2826,N_15,N_63);
nand U2827 (N_2827,N_767,N_275);
nand U2828 (N_2828,N_813,N_1087);
or U2829 (N_2829,N_1000,N_1497);
nand U2830 (N_2830,N_1343,N_561);
and U2831 (N_2831,N_1382,N_1328);
nand U2832 (N_2832,N_1490,N_632);
nand U2833 (N_2833,N_1252,N_915);
nand U2834 (N_2834,N_1263,N_14);
xor U2835 (N_2835,N_1401,N_473);
or U2836 (N_2836,N_1093,N_1465);
and U2837 (N_2837,N_679,N_769);
or U2838 (N_2838,N_976,N_695);
nand U2839 (N_2839,N_492,N_1062);
nor U2840 (N_2840,N_268,N_920);
or U2841 (N_2841,N_812,N_93);
nand U2842 (N_2842,N_1126,N_403);
or U2843 (N_2843,N_333,N_194);
or U2844 (N_2844,N_295,N_246);
or U2845 (N_2845,N_875,N_118);
nand U2846 (N_2846,N_476,N_467);
and U2847 (N_2847,N_730,N_1353);
and U2848 (N_2848,N_545,N_1183);
and U2849 (N_2849,N_102,N_1218);
and U2850 (N_2850,N_1313,N_806);
and U2851 (N_2851,N_652,N_1393);
and U2852 (N_2852,N_309,N_886);
nand U2853 (N_2853,N_1045,N_477);
or U2854 (N_2854,N_1220,N_190);
and U2855 (N_2855,N_625,N_1371);
or U2856 (N_2856,N_559,N_786);
or U2857 (N_2857,N_922,N_751);
or U2858 (N_2858,N_848,N_402);
or U2859 (N_2859,N_1313,N_466);
nand U2860 (N_2860,N_587,N_318);
nand U2861 (N_2861,N_533,N_1153);
and U2862 (N_2862,N_436,N_1226);
or U2863 (N_2863,N_904,N_1436);
or U2864 (N_2864,N_819,N_730);
nand U2865 (N_2865,N_487,N_841);
or U2866 (N_2866,N_490,N_1318);
or U2867 (N_2867,N_319,N_312);
nor U2868 (N_2868,N_965,N_1347);
nand U2869 (N_2869,N_1092,N_1466);
nor U2870 (N_2870,N_808,N_819);
or U2871 (N_2871,N_434,N_992);
xor U2872 (N_2872,N_267,N_1292);
or U2873 (N_2873,N_1408,N_330);
nor U2874 (N_2874,N_853,N_1469);
nor U2875 (N_2875,N_1088,N_21);
nand U2876 (N_2876,N_1405,N_931);
nand U2877 (N_2877,N_971,N_1265);
and U2878 (N_2878,N_647,N_173);
or U2879 (N_2879,N_1476,N_725);
or U2880 (N_2880,N_945,N_391);
nor U2881 (N_2881,N_594,N_260);
and U2882 (N_2882,N_121,N_1119);
nand U2883 (N_2883,N_420,N_533);
and U2884 (N_2884,N_277,N_1496);
and U2885 (N_2885,N_650,N_0);
or U2886 (N_2886,N_576,N_32);
nand U2887 (N_2887,N_565,N_554);
or U2888 (N_2888,N_242,N_1176);
or U2889 (N_2889,N_1477,N_730);
and U2890 (N_2890,N_1403,N_578);
or U2891 (N_2891,N_143,N_1477);
nor U2892 (N_2892,N_1344,N_1277);
nor U2893 (N_2893,N_464,N_1356);
nand U2894 (N_2894,N_1433,N_126);
nor U2895 (N_2895,N_77,N_1133);
nor U2896 (N_2896,N_1023,N_234);
and U2897 (N_2897,N_795,N_256);
nand U2898 (N_2898,N_393,N_869);
or U2899 (N_2899,N_213,N_370);
nand U2900 (N_2900,N_78,N_106);
and U2901 (N_2901,N_1339,N_13);
nor U2902 (N_2902,N_698,N_152);
or U2903 (N_2903,N_613,N_542);
nand U2904 (N_2904,N_1262,N_1484);
and U2905 (N_2905,N_1465,N_1308);
nand U2906 (N_2906,N_675,N_1322);
or U2907 (N_2907,N_68,N_1440);
nand U2908 (N_2908,N_796,N_705);
nand U2909 (N_2909,N_111,N_1136);
and U2910 (N_2910,N_485,N_254);
nor U2911 (N_2911,N_1318,N_613);
nor U2912 (N_2912,N_960,N_936);
or U2913 (N_2913,N_13,N_708);
or U2914 (N_2914,N_619,N_1432);
nand U2915 (N_2915,N_905,N_652);
or U2916 (N_2916,N_412,N_1022);
or U2917 (N_2917,N_644,N_556);
nand U2918 (N_2918,N_1404,N_1249);
and U2919 (N_2919,N_280,N_834);
nand U2920 (N_2920,N_704,N_430);
nand U2921 (N_2921,N_1254,N_21);
nand U2922 (N_2922,N_927,N_723);
or U2923 (N_2923,N_1432,N_811);
nand U2924 (N_2924,N_560,N_1215);
or U2925 (N_2925,N_415,N_337);
or U2926 (N_2926,N_823,N_664);
and U2927 (N_2927,N_233,N_56);
nor U2928 (N_2928,N_1249,N_177);
nor U2929 (N_2929,N_156,N_1111);
and U2930 (N_2930,N_712,N_1231);
nor U2931 (N_2931,N_779,N_1439);
nand U2932 (N_2932,N_1292,N_738);
and U2933 (N_2933,N_1032,N_1456);
nor U2934 (N_2934,N_1240,N_680);
nand U2935 (N_2935,N_1338,N_172);
or U2936 (N_2936,N_1274,N_760);
nor U2937 (N_2937,N_725,N_518);
nor U2938 (N_2938,N_946,N_933);
or U2939 (N_2939,N_1342,N_313);
nor U2940 (N_2940,N_1123,N_1179);
and U2941 (N_2941,N_1238,N_411);
nand U2942 (N_2942,N_1017,N_1172);
nor U2943 (N_2943,N_1024,N_22);
and U2944 (N_2944,N_644,N_684);
or U2945 (N_2945,N_1434,N_448);
nor U2946 (N_2946,N_645,N_995);
nand U2947 (N_2947,N_753,N_1086);
nand U2948 (N_2948,N_299,N_1296);
nand U2949 (N_2949,N_904,N_596);
and U2950 (N_2950,N_2,N_1011);
and U2951 (N_2951,N_160,N_1266);
xor U2952 (N_2952,N_68,N_34);
nor U2953 (N_2953,N_624,N_1420);
or U2954 (N_2954,N_1201,N_668);
nor U2955 (N_2955,N_1049,N_1487);
nor U2956 (N_2956,N_1336,N_233);
nand U2957 (N_2957,N_1053,N_1001);
or U2958 (N_2958,N_1432,N_1266);
and U2959 (N_2959,N_320,N_214);
and U2960 (N_2960,N_1432,N_1421);
nand U2961 (N_2961,N_914,N_1492);
and U2962 (N_2962,N_606,N_422);
and U2963 (N_2963,N_1026,N_83);
nand U2964 (N_2964,N_1283,N_370);
and U2965 (N_2965,N_110,N_1167);
or U2966 (N_2966,N_199,N_1475);
or U2967 (N_2967,N_175,N_450);
nand U2968 (N_2968,N_1348,N_978);
or U2969 (N_2969,N_1005,N_1491);
or U2970 (N_2970,N_494,N_793);
and U2971 (N_2971,N_1006,N_37);
or U2972 (N_2972,N_1488,N_811);
nor U2973 (N_2973,N_722,N_597);
nand U2974 (N_2974,N_1196,N_486);
or U2975 (N_2975,N_1418,N_1183);
and U2976 (N_2976,N_501,N_1393);
or U2977 (N_2977,N_694,N_852);
and U2978 (N_2978,N_847,N_473);
xnor U2979 (N_2979,N_1014,N_702);
nand U2980 (N_2980,N_87,N_89);
or U2981 (N_2981,N_1484,N_1073);
nor U2982 (N_2982,N_676,N_324);
or U2983 (N_2983,N_912,N_186);
nand U2984 (N_2984,N_1289,N_1338);
and U2985 (N_2985,N_683,N_782);
and U2986 (N_2986,N_869,N_494);
nand U2987 (N_2987,N_1009,N_395);
or U2988 (N_2988,N_1231,N_292);
nor U2989 (N_2989,N_297,N_467);
and U2990 (N_2990,N_1363,N_222);
nor U2991 (N_2991,N_1273,N_1405);
nor U2992 (N_2992,N_1313,N_1010);
or U2993 (N_2993,N_1384,N_1108);
and U2994 (N_2994,N_628,N_1005);
nor U2995 (N_2995,N_1473,N_1409);
nor U2996 (N_2996,N_1414,N_1262);
and U2997 (N_2997,N_1416,N_162);
nand U2998 (N_2998,N_715,N_120);
or U2999 (N_2999,N_1380,N_1114);
nand U3000 (N_3000,N_2448,N_1671);
or U3001 (N_3001,N_1619,N_1872);
and U3002 (N_3002,N_2926,N_2664);
nand U3003 (N_3003,N_1588,N_2820);
and U3004 (N_3004,N_1895,N_1755);
nand U3005 (N_3005,N_2047,N_2779);
or U3006 (N_3006,N_1553,N_2328);
or U3007 (N_3007,N_2471,N_1552);
nor U3008 (N_3008,N_1854,N_2075);
nor U3009 (N_3009,N_1633,N_2059);
nor U3010 (N_3010,N_1740,N_1695);
and U3011 (N_3011,N_2366,N_1710);
nor U3012 (N_3012,N_2964,N_2032);
or U3013 (N_3013,N_1601,N_1592);
nand U3014 (N_3014,N_2469,N_1545);
and U3015 (N_3015,N_1738,N_1911);
nand U3016 (N_3016,N_1668,N_2860);
xor U3017 (N_3017,N_2805,N_2135);
nor U3018 (N_3018,N_1519,N_2463);
or U3019 (N_3019,N_2988,N_1834);
and U3020 (N_3020,N_2058,N_1946);
nand U3021 (N_3021,N_2434,N_2036);
or U3022 (N_3022,N_2626,N_2644);
xor U3023 (N_3023,N_1739,N_1888);
and U3024 (N_3024,N_2281,N_2423);
or U3025 (N_3025,N_2505,N_1696);
or U3026 (N_3026,N_1896,N_2690);
nor U3027 (N_3027,N_1792,N_1930);
and U3028 (N_3028,N_2193,N_2192);
nand U3029 (N_3029,N_1628,N_2236);
nor U3030 (N_3030,N_1608,N_2148);
nand U3031 (N_3031,N_1977,N_2649);
nand U3032 (N_3032,N_1921,N_2057);
nor U3033 (N_3033,N_2859,N_1874);
nor U3034 (N_3034,N_1630,N_2747);
and U3035 (N_3035,N_2283,N_1865);
and U3036 (N_3036,N_2321,N_1817);
nor U3037 (N_3037,N_2014,N_1596);
or U3038 (N_3038,N_2580,N_2556);
nand U3039 (N_3039,N_2396,N_2169);
and U3040 (N_3040,N_1652,N_2352);
and U3041 (N_3041,N_2833,N_2545);
or U3042 (N_3042,N_2204,N_2008);
or U3043 (N_3043,N_2186,N_1751);
and U3044 (N_3044,N_2137,N_2245);
nor U3045 (N_3045,N_2957,N_1893);
nor U3046 (N_3046,N_1706,N_1867);
and U3047 (N_3047,N_2220,N_2373);
nand U3048 (N_3048,N_2242,N_2459);
nor U3049 (N_3049,N_1535,N_1793);
or U3050 (N_3050,N_2677,N_2643);
or U3051 (N_3051,N_2138,N_1501);
nand U3052 (N_3052,N_1569,N_2409);
and U3053 (N_3053,N_1610,N_1606);
or U3054 (N_3054,N_2495,N_1522);
and U3055 (N_3055,N_1530,N_2349);
or U3056 (N_3056,N_2771,N_1791);
nand U3057 (N_3057,N_2415,N_2101);
nor U3058 (N_3058,N_2397,N_1678);
or U3059 (N_3059,N_2737,N_1887);
nor U3060 (N_3060,N_1944,N_2249);
nand U3061 (N_3061,N_2708,N_1635);
or U3062 (N_3062,N_1987,N_2834);
and U3063 (N_3063,N_2878,N_1853);
or U3064 (N_3064,N_2441,N_2661);
and U3065 (N_3065,N_2067,N_2322);
xnor U3066 (N_3066,N_2082,N_2061);
nor U3067 (N_3067,N_1849,N_1932);
nand U3068 (N_3068,N_1866,N_1900);
nor U3069 (N_3069,N_1638,N_2854);
and U3070 (N_3070,N_2460,N_2103);
or U3071 (N_3071,N_2385,N_2935);
nor U3072 (N_3072,N_1787,N_2778);
or U3073 (N_3073,N_1960,N_2080);
and U3074 (N_3074,N_2210,N_1705);
nand U3075 (N_3075,N_2143,N_2149);
nor U3076 (N_3076,N_1937,N_2630);
or U3077 (N_3077,N_2458,N_2631);
or U3078 (N_3078,N_1770,N_2377);
or U3079 (N_3079,N_2917,N_1514);
and U3080 (N_3080,N_1841,N_2002);
or U3081 (N_3081,N_2313,N_2368);
or U3082 (N_3082,N_2425,N_1744);
nor U3083 (N_3083,N_1945,N_1894);
and U3084 (N_3084,N_2121,N_2503);
or U3085 (N_3085,N_2274,N_2674);
and U3086 (N_3086,N_1838,N_1684);
or U3087 (N_3087,N_2601,N_1627);
nor U3088 (N_3088,N_1617,N_2217);
nand U3089 (N_3089,N_2003,N_2983);
nand U3090 (N_3090,N_1513,N_2603);
or U3091 (N_3091,N_2299,N_1728);
or U3092 (N_3092,N_1529,N_2710);
and U3093 (N_3093,N_2861,N_2476);
and U3094 (N_3094,N_1917,N_1583);
nor U3095 (N_3095,N_2892,N_2826);
nor U3096 (N_3096,N_2740,N_1547);
or U3097 (N_3097,N_2683,N_2344);
nand U3098 (N_3098,N_2413,N_1616);
and U3099 (N_3099,N_1557,N_2178);
or U3100 (N_3100,N_1796,N_1861);
or U3101 (N_3101,N_2386,N_2694);
or U3102 (N_3102,N_2657,N_1839);
and U3103 (N_3103,N_2345,N_1526);
or U3104 (N_3104,N_2177,N_1971);
and U3105 (N_3105,N_2754,N_2623);
or U3106 (N_3106,N_2009,N_2327);
nand U3107 (N_3107,N_1570,N_1748);
nor U3108 (N_3108,N_2931,N_1644);
or U3109 (N_3109,N_2675,N_2351);
or U3110 (N_3110,N_2090,N_2842);
or U3111 (N_3111,N_2488,N_1912);
nand U3112 (N_3112,N_2403,N_2532);
or U3113 (N_3113,N_2087,N_2038);
or U3114 (N_3114,N_2071,N_2222);
or U3115 (N_3115,N_1844,N_2006);
or U3116 (N_3116,N_1502,N_2714);
and U3117 (N_3117,N_2929,N_1711);
or U3118 (N_3118,N_2165,N_2611);
or U3119 (N_3119,N_1624,N_2232);
nor U3120 (N_3120,N_2589,N_2891);
nor U3121 (N_3121,N_2678,N_2994);
nor U3122 (N_3122,N_1807,N_2915);
nor U3123 (N_3123,N_2456,N_2965);
nor U3124 (N_3124,N_1587,N_2384);
nor U3125 (N_3125,N_2855,N_2371);
and U3126 (N_3126,N_2906,N_2596);
nor U3127 (N_3127,N_1979,N_2703);
and U3128 (N_3128,N_2319,N_1753);
or U3129 (N_3129,N_2510,N_2147);
or U3130 (N_3130,N_1717,N_2506);
nand U3131 (N_3131,N_1762,N_1618);
or U3132 (N_3132,N_2619,N_2836);
and U3133 (N_3133,N_1585,N_2986);
or U3134 (N_3134,N_2326,N_2173);
or U3135 (N_3135,N_2880,N_2231);
and U3136 (N_3136,N_1731,N_2077);
nor U3137 (N_3137,N_1968,N_2467);
and U3138 (N_3138,N_2314,N_2582);
and U3139 (N_3139,N_2911,N_2879);
nor U3140 (N_3140,N_2332,N_1732);
nor U3141 (N_3141,N_2205,N_2837);
and U3142 (N_3142,N_2337,N_2557);
nand U3143 (N_3143,N_2392,N_2381);
or U3144 (N_3144,N_2307,N_1508);
or U3145 (N_3145,N_2017,N_2435);
nand U3146 (N_3146,N_1603,N_1609);
nand U3147 (N_3147,N_2498,N_2168);
or U3148 (N_3148,N_1634,N_1850);
nor U3149 (N_3149,N_2849,N_2194);
and U3150 (N_3150,N_2440,N_2172);
or U3151 (N_3151,N_1701,N_2133);
or U3152 (N_3152,N_1563,N_1537);
nand U3153 (N_3153,N_2844,N_2374);
or U3154 (N_3154,N_2908,N_1795);
nor U3155 (N_3155,N_1540,N_2685);
nor U3156 (N_3156,N_2745,N_2115);
nand U3157 (N_3157,N_1599,N_1969);
nand U3158 (N_3158,N_2539,N_2436);
nand U3159 (N_3159,N_2579,N_2478);
nor U3160 (N_3160,N_2821,N_1980);
nand U3161 (N_3161,N_2259,N_1590);
and U3162 (N_3162,N_2789,N_1524);
and U3163 (N_3163,N_2241,N_2527);
nand U3164 (N_3164,N_2890,N_1646);
nand U3165 (N_3165,N_1811,N_2127);
or U3166 (N_3166,N_2011,N_2760);
or U3167 (N_3167,N_2991,N_1669);
and U3168 (N_3168,N_2798,N_2612);
or U3169 (N_3169,N_2736,N_2095);
and U3170 (N_3170,N_2227,N_2128);
nor U3171 (N_3171,N_1859,N_2540);
and U3172 (N_3172,N_2741,N_2054);
and U3173 (N_3173,N_2066,N_2682);
nand U3174 (N_3174,N_1639,N_1936);
nor U3175 (N_3175,N_1822,N_1768);
nor U3176 (N_3176,N_2752,N_2156);
nand U3177 (N_3177,N_1851,N_2049);
or U3178 (N_3178,N_2786,N_1730);
and U3179 (N_3179,N_1923,N_1614);
nand U3180 (N_3180,N_1901,N_2144);
and U3181 (N_3181,N_1658,N_2230);
nor U3182 (N_3182,N_1902,N_2790);
or U3183 (N_3183,N_1809,N_1892);
or U3184 (N_3184,N_1546,N_2555);
or U3185 (N_3185,N_2429,N_2875);
nor U3186 (N_3186,N_2781,N_2372);
nand U3187 (N_3187,N_2564,N_2375);
or U3188 (N_3188,N_2487,N_2370);
nand U3189 (N_3189,N_2602,N_1682);
and U3190 (N_3190,N_2079,N_1500);
nor U3191 (N_3191,N_2431,N_1881);
and U3192 (N_3192,N_2735,N_2852);
and U3193 (N_3193,N_2667,N_2722);
nand U3194 (N_3194,N_1516,N_1565);
nand U3195 (N_3195,N_1788,N_2533);
nand U3196 (N_3196,N_2195,N_2438);
or U3197 (N_3197,N_1813,N_2828);
nor U3198 (N_3198,N_2970,N_2251);
or U3199 (N_3199,N_2235,N_2025);
or U3200 (N_3200,N_1725,N_1784);
nand U3201 (N_3201,N_2605,N_1871);
and U3202 (N_3202,N_2998,N_2560);
nand U3203 (N_3203,N_2401,N_2762);
or U3204 (N_3204,N_2767,N_2997);
or U3205 (N_3205,N_2806,N_2553);
nand U3206 (N_3206,N_2813,N_2807);
or U3207 (N_3207,N_2721,N_2584);
or U3208 (N_3208,N_2485,N_2260);
nand U3209 (N_3209,N_2216,N_2428);
or U3210 (N_3210,N_2289,N_2286);
nand U3211 (N_3211,N_2829,N_2823);
and U3212 (N_3212,N_1852,N_2300);
nand U3213 (N_3213,N_2543,N_2309);
and U3214 (N_3214,N_2883,N_2520);
nor U3215 (N_3215,N_2554,N_2316);
nor U3216 (N_3216,N_1727,N_2432);
nand U3217 (N_3217,N_2018,N_1612);
xnor U3218 (N_3218,N_2412,N_1840);
or U3219 (N_3219,N_2268,N_1721);
and U3220 (N_3220,N_2160,N_2347);
nor U3221 (N_3221,N_2224,N_2175);
nor U3222 (N_3222,N_1745,N_1602);
nor U3223 (N_3223,N_2483,N_2953);
nor U3224 (N_3224,N_2992,N_1995);
nor U3225 (N_3225,N_2943,N_2551);
and U3226 (N_3226,N_2726,N_2125);
nand U3227 (N_3227,N_1800,N_2910);
nand U3228 (N_3228,N_2862,N_2362);
nor U3229 (N_3229,N_2393,N_1577);
nor U3230 (N_3230,N_2581,N_2330);
nor U3231 (N_3231,N_2907,N_1607);
nand U3232 (N_3232,N_1988,N_2457);
and U3233 (N_3233,N_2023,N_1857);
or U3234 (N_3234,N_1782,N_2398);
or U3235 (N_3235,N_1690,N_1961);
or U3236 (N_3236,N_2706,N_1919);
or U3237 (N_3237,N_2831,N_2206);
nor U3238 (N_3238,N_2407,N_2124);
nand U3239 (N_3239,N_1720,N_2119);
and U3240 (N_3240,N_2013,N_1799);
or U3241 (N_3241,N_1708,N_2824);
or U3242 (N_3242,N_1642,N_2938);
nor U3243 (N_3243,N_2772,N_2261);
nand U3244 (N_3244,N_1786,N_2461);
or U3245 (N_3245,N_2376,N_2120);
nor U3246 (N_3246,N_1972,N_2639);
or U3247 (N_3247,N_1832,N_2094);
and U3248 (N_3248,N_2507,N_1512);
or U3249 (N_3249,N_1794,N_2154);
or U3250 (N_3250,N_2999,N_2499);
nand U3251 (N_3251,N_2234,N_2141);
and U3252 (N_3252,N_1962,N_2257);
nand U3253 (N_3253,N_2214,N_2621);
and U3254 (N_3254,N_2107,N_2815);
nand U3255 (N_3255,N_2780,N_2868);
nor U3256 (N_3256,N_2599,N_1655);
and U3257 (N_3257,N_2711,N_1543);
or U3258 (N_3258,N_2001,N_2944);
nand U3259 (N_3259,N_1672,N_2742);
nor U3260 (N_3260,N_1771,N_2808);
or U3261 (N_3261,N_1951,N_1976);
or U3262 (N_3262,N_1935,N_2404);
nor U3263 (N_3263,N_1981,N_1802);
nand U3264 (N_3264,N_2524,N_2963);
nand U3265 (N_3265,N_2616,N_2816);
nand U3266 (N_3266,N_1582,N_2272);
nor U3267 (N_3267,N_1518,N_2296);
nor U3268 (N_3268,N_2365,N_2538);
or U3269 (N_3269,N_1940,N_1525);
and U3270 (N_3270,N_2768,N_2208);
and U3271 (N_3271,N_2052,N_1670);
nor U3272 (N_3272,N_1846,N_2288);
nor U3273 (N_3273,N_1922,N_1580);
xnor U3274 (N_3274,N_1949,N_2455);
nor U3275 (N_3275,N_2550,N_2652);
or U3276 (N_3276,N_1589,N_2695);
xnor U3277 (N_3277,N_1566,N_1918);
and U3278 (N_3278,N_1600,N_2012);
and U3279 (N_3279,N_2764,N_2010);
nand U3280 (N_3280,N_2114,N_1831);
and U3281 (N_3281,N_2343,N_2660);
and U3282 (N_3282,N_1562,N_1803);
or U3283 (N_3283,N_1964,N_1629);
nand U3284 (N_3284,N_2750,N_2294);
and U3285 (N_3285,N_2255,N_2191);
and U3286 (N_3286,N_2131,N_1510);
and U3287 (N_3287,N_1989,N_2720);
nor U3288 (N_3288,N_2548,N_2161);
or U3289 (N_3289,N_2521,N_1576);
nand U3290 (N_3290,N_2357,N_1666);
nor U3291 (N_3291,N_2034,N_2243);
nor U3292 (N_3292,N_2229,N_1882);
or U3293 (N_3293,N_2648,N_2671);
or U3294 (N_3294,N_2250,N_2704);
and U3295 (N_3295,N_2426,N_2367);
nand U3296 (N_3296,N_2895,N_1760);
nand U3297 (N_3297,N_2788,N_1824);
and U3298 (N_3298,N_2285,N_2586);
or U3299 (N_3299,N_2884,N_2233);
or U3300 (N_3300,N_2512,N_2200);
or U3301 (N_3301,N_2350,N_2716);
nand U3302 (N_3302,N_1722,N_2867);
or U3303 (N_3303,N_2793,N_2291);
nor U3304 (N_3304,N_2201,N_2402);
nand U3305 (N_3305,N_2874,N_1827);
and U3306 (N_3306,N_2699,N_1780);
nor U3307 (N_3307,N_2015,N_2841);
nand U3308 (N_3308,N_2853,N_2091);
nand U3309 (N_3309,N_2866,N_2575);
nand U3310 (N_3310,N_1598,N_2615);
or U3311 (N_3311,N_2989,N_1908);
nand U3312 (N_3312,N_2635,N_2587);
nor U3313 (N_3313,N_2684,N_1659);
and U3314 (N_3314,N_2787,N_2723);
nor U3315 (N_3315,N_1724,N_1568);
and U3316 (N_3316,N_2045,N_2857);
or U3317 (N_3317,N_1676,N_2338);
or U3318 (N_3318,N_2387,N_2123);
nand U3319 (N_3319,N_2702,N_2016);
nor U3320 (N_3320,N_1880,N_1656);
nor U3321 (N_3321,N_2382,N_2089);
and U3322 (N_3322,N_2305,N_2048);
nand U3323 (N_3323,N_1595,N_2676);
nand U3324 (N_3324,N_2610,N_1856);
nand U3325 (N_3325,N_2600,N_2406);
nand U3326 (N_3326,N_2620,N_1926);
and U3327 (N_3327,N_2183,N_2361);
nor U3328 (N_3328,N_2159,N_2430);
and U3329 (N_3329,N_2633,N_2697);
and U3330 (N_3330,N_1574,N_1560);
xnor U3331 (N_3331,N_2056,N_1556);
and U3332 (N_3332,N_1571,N_2496);
nor U3333 (N_3333,N_2005,N_2982);
nand U3334 (N_3334,N_2670,N_2215);
and U3335 (N_3335,N_1531,N_2419);
nor U3336 (N_3336,N_2881,N_2244);
and U3337 (N_3337,N_1691,N_2271);
nor U3338 (N_3338,N_2170,N_2563);
nor U3339 (N_3339,N_2565,N_1645);
or U3340 (N_3340,N_2663,N_2253);
nand U3341 (N_3341,N_2863,N_1998);
and U3342 (N_3342,N_2707,N_1978);
nand U3343 (N_3343,N_1815,N_2207);
nor U3344 (N_3344,N_1667,N_1662);
and U3345 (N_3345,N_2689,N_2973);
and U3346 (N_3346,N_2761,N_2814);
nor U3347 (N_3347,N_2902,N_1653);
or U3348 (N_3348,N_2072,N_2606);
and U3349 (N_3349,N_1673,N_2749);
nor U3350 (N_3350,N_2925,N_2967);
nand U3351 (N_3351,N_1761,N_2899);
nor U3352 (N_3352,N_2604,N_2282);
nand U3353 (N_3353,N_1864,N_2809);
and U3354 (N_3354,N_2665,N_2559);
and U3355 (N_3355,N_2515,N_1956);
nand U3356 (N_3356,N_2427,N_2151);
nand U3357 (N_3357,N_2197,N_2358);
and U3358 (N_3358,N_2535,N_1909);
nand U3359 (N_3359,N_2093,N_2948);
or U3360 (N_3360,N_2027,N_2951);
nand U3361 (N_3361,N_1920,N_2629);
or U3362 (N_3362,N_1804,N_1506);
nand U3363 (N_3363,N_2031,N_2627);
nor U3364 (N_3364,N_1891,N_2042);
and U3365 (N_3365,N_1643,N_2035);
nor U3366 (N_3366,N_2889,N_1876);
nor U3367 (N_3367,N_1747,N_2292);
nand U3368 (N_3368,N_2391,N_2295);
or U3369 (N_3369,N_2185,N_1651);
nand U3370 (N_3370,N_2417,N_2166);
nand U3371 (N_3371,N_2418,N_2980);
and U3372 (N_3372,N_2074,N_1611);
and U3373 (N_3373,N_2645,N_1620);
and U3374 (N_3374,N_1757,N_2731);
nand U3375 (N_3375,N_2508,N_1636);
and U3376 (N_3376,N_2150,N_2848);
and U3377 (N_3377,N_2680,N_2339);
nor U3378 (N_3378,N_2996,N_1835);
nand U3379 (N_3379,N_1776,N_1613);
or U3380 (N_3380,N_2654,N_2930);
nand U3381 (N_3381,N_2795,N_2445);
or U3382 (N_3382,N_2940,N_1503);
nor U3383 (N_3383,N_2709,N_1798);
nand U3384 (N_3384,N_2298,N_1953);
and U3385 (N_3385,N_1712,N_2977);
nand U3386 (N_3386,N_1523,N_1699);
or U3387 (N_3387,N_2053,N_2571);
nor U3388 (N_3388,N_1916,N_1847);
nor U3389 (N_3389,N_2656,N_2993);
nor U3390 (N_3390,N_2024,N_2437);
and U3391 (N_3391,N_1594,N_1975);
and U3392 (N_3392,N_1713,N_1575);
and U3393 (N_3393,N_1982,N_2378);
or U3394 (N_3394,N_1879,N_2701);
nor U3395 (N_3395,N_1763,N_2987);
nor U3396 (N_3396,N_2395,N_2746);
or U3397 (N_3397,N_2822,N_1870);
nand U3398 (N_3398,N_1842,N_1848);
nor U3399 (N_3399,N_2084,N_2497);
or U3400 (N_3400,N_2753,N_2353);
nand U3401 (N_3401,N_1914,N_2717);
and U3402 (N_3402,N_1764,N_2569);
nor U3403 (N_3403,N_2939,N_2912);
or U3404 (N_3404,N_2923,N_2791);
nand U3405 (N_3405,N_2738,N_2410);
and U3406 (N_3406,N_1715,N_2482);
and U3407 (N_3407,N_2390,N_2140);
nand U3408 (N_3408,N_1735,N_2021);
nor U3409 (N_3409,N_2333,N_1505);
nor U3410 (N_3410,N_2408,N_2713);
or U3411 (N_3411,N_2162,N_1873);
nand U3412 (N_3412,N_1756,N_2287);
nand U3413 (N_3413,N_2256,N_2715);
nand U3414 (N_3414,N_1772,N_2774);
or U3415 (N_3415,N_2696,N_2466);
nand U3416 (N_3416,N_2802,N_2182);
or U3417 (N_3417,N_1928,N_2751);
nand U3418 (N_3418,N_2422,N_2803);
nor U3419 (N_3419,N_2450,N_1622);
nor U3420 (N_3420,N_2609,N_1778);
nand U3421 (N_3421,N_2625,N_2076);
or U3422 (N_3422,N_1759,N_1536);
nand U3423 (N_3423,N_1663,N_2122);
and U3424 (N_3424,N_2636,N_2226);
and U3425 (N_3425,N_2876,N_1777);
nand U3426 (N_3426,N_2946,N_2153);
and U3427 (N_3427,N_1548,N_2552);
and U3428 (N_3428,N_2439,N_2062);
nor U3429 (N_3429,N_1504,N_2509);
or U3430 (N_3430,N_1517,N_2669);
and U3431 (N_3431,N_2896,N_1752);
or U3432 (N_3432,N_2985,N_1743);
and U3433 (N_3433,N_1929,N_2254);
and U3434 (N_3434,N_2632,N_2421);
nand U3435 (N_3435,N_2484,N_2519);
or U3436 (N_3436,N_2190,N_2920);
and U3437 (N_3437,N_2356,N_2026);
or U3438 (N_3438,N_2083,N_1700);
nor U3439 (N_3439,N_2511,N_2394);
nor U3440 (N_3440,N_1604,N_2537);
or U3441 (N_3441,N_2473,N_2870);
nand U3442 (N_3442,N_2976,N_2634);
and U3443 (N_3443,N_2613,N_2102);
and U3444 (N_3444,N_2744,N_1697);
and U3445 (N_3445,N_2187,N_1555);
nand U3446 (N_3446,N_2196,N_1773);
or U3447 (N_3447,N_2624,N_1775);
nor U3448 (N_3448,N_1597,N_2755);
or U3449 (N_3449,N_2475,N_2134);
or U3450 (N_3450,N_2481,N_2566);
or U3451 (N_3451,N_2486,N_2681);
or U3452 (N_3452,N_1886,N_2562);
nand U3453 (N_3453,N_2819,N_2145);
and U3454 (N_3454,N_2040,N_1907);
and U3455 (N_3455,N_2850,N_2942);
nand U3456 (N_3456,N_2302,N_2546);
nor U3457 (N_3457,N_2974,N_2389);
nand U3458 (N_3458,N_2468,N_2284);
nor U3459 (N_3459,N_2118,N_2536);
nor U3460 (N_3460,N_2088,N_2591);
and U3461 (N_3461,N_1591,N_2462);
nand U3462 (N_3462,N_2733,N_2280);
nor U3463 (N_3463,N_2668,N_1869);
or U3464 (N_3464,N_2578,N_2959);
nor U3465 (N_3465,N_1812,N_1833);
and U3466 (N_3466,N_2223,N_2766);
and U3467 (N_3467,N_1814,N_2491);
nand U3468 (N_3468,N_2941,N_2672);
nand U3469 (N_3469,N_2894,N_1990);
nor U3470 (N_3470,N_2388,N_1890);
and U3471 (N_3471,N_2189,N_1938);
nand U3472 (N_3472,N_1750,N_2157);
nor U3473 (N_3473,N_2163,N_2638);
nand U3474 (N_3474,N_1654,N_1878);
and U3475 (N_3475,N_2492,N_2900);
and U3476 (N_3476,N_1623,N_2158);
and U3477 (N_3477,N_1781,N_1718);
nand U3478 (N_3478,N_1819,N_2927);
or U3479 (N_3479,N_1694,N_1765);
nor U3480 (N_3480,N_2096,N_2278);
nand U3481 (N_3481,N_2801,N_1943);
nor U3482 (N_3482,N_1933,N_2360);
and U3483 (N_3483,N_2293,N_2129);
nor U3484 (N_3484,N_1675,N_2990);
and U3485 (N_3485,N_2325,N_1572);
nand U3486 (N_3486,N_2732,N_2692);
or U3487 (N_3487,N_2922,N_2901);
or U3488 (N_3488,N_2060,N_2203);
nor U3489 (N_3489,N_2174,N_2264);
nor U3490 (N_3490,N_2830,N_1955);
nor U3491 (N_3491,N_2777,N_1704);
nor U3492 (N_3492,N_2529,N_2734);
nor U3493 (N_3493,N_1843,N_1805);
nand U3494 (N_3494,N_2651,N_2310);
or U3495 (N_3495,N_1970,N_1959);
or U3496 (N_3496,N_1790,N_1785);
or U3497 (N_3497,N_1736,N_1862);
and U3498 (N_3498,N_2770,N_2950);
or U3499 (N_3499,N_2958,N_2355);
nand U3500 (N_3500,N_2724,N_2642);
and U3501 (N_3501,N_2240,N_2188);
nor U3502 (N_3502,N_2981,N_2308);
nand U3503 (N_3503,N_2465,N_1942);
and U3504 (N_3504,N_1966,N_2311);
nor U3505 (N_3505,N_2501,N_1665);
nand U3506 (N_3506,N_2743,N_2739);
nand U3507 (N_3507,N_2269,N_2909);
or U3508 (N_3508,N_2653,N_2763);
nand U3509 (N_3509,N_1957,N_2655);
or U3510 (N_3510,N_2864,N_1661);
or U3511 (N_3511,N_2567,N_1741);
nand U3512 (N_3512,N_2202,N_2019);
or U3513 (N_3513,N_1649,N_2905);
nor U3514 (N_3514,N_1991,N_2033);
and U3515 (N_3515,N_2198,N_2769);
nand U3516 (N_3516,N_2303,N_1637);
nor U3517 (N_3517,N_1816,N_2975);
nand U3518 (N_3518,N_2936,N_2116);
and U3519 (N_3519,N_2811,N_1564);
nor U3520 (N_3520,N_1657,N_2446);
or U3521 (N_3521,N_2290,N_2542);
or U3522 (N_3522,N_1974,N_1579);
nor U3523 (N_3523,N_1541,N_1534);
nor U3524 (N_3524,N_1766,N_2247);
and U3525 (N_3525,N_2152,N_1883);
and U3526 (N_3526,N_1605,N_2383);
or U3527 (N_3527,N_1687,N_2794);
nand U3528 (N_3528,N_1640,N_2238);
nand U3529 (N_3529,N_2765,N_1797);
nor U3530 (N_3530,N_2776,N_2614);
xor U3531 (N_3531,N_2593,N_2030);
or U3532 (N_3532,N_1714,N_2306);
or U3533 (N_3533,N_2098,N_1931);
nor U3534 (N_3534,N_2252,N_2525);
nand U3535 (N_3535,N_2179,N_1586);
nor U3536 (N_3536,N_2934,N_2452);
nand U3537 (N_3537,N_2444,N_2420);
nor U3538 (N_3538,N_1660,N_2775);
or U3539 (N_3539,N_1996,N_2693);
or U3540 (N_3540,N_1904,N_1924);
or U3541 (N_3541,N_1550,N_2405);
nor U3542 (N_3542,N_2176,N_1573);
or U3543 (N_3543,N_2954,N_2516);
and U3544 (N_3544,N_2758,N_2592);
nor U3545 (N_3545,N_1950,N_2181);
and U3546 (N_3546,N_2691,N_1703);
or U3547 (N_3547,N_1626,N_2126);
or U3548 (N_3548,N_2514,N_2213);
nor U3549 (N_3549,N_1681,N_2199);
nand U3550 (N_3550,N_2832,N_2972);
and U3551 (N_3551,N_1947,N_1719);
and U3552 (N_3552,N_2583,N_2044);
or U3553 (N_3553,N_2504,N_2784);
nor U3554 (N_3554,N_2847,N_2335);
or U3555 (N_3555,N_2346,N_1559);
and U3556 (N_3556,N_2359,N_2329);
or U3557 (N_3557,N_2817,N_1898);
or U3558 (N_3558,N_2518,N_2212);
nand U3559 (N_3559,N_2718,N_2051);
and U3560 (N_3560,N_2962,N_1688);
nand U3561 (N_3561,N_1897,N_1542);
and U3562 (N_3562,N_2472,N_2812);
nor U3563 (N_3563,N_1963,N_2871);
nor U3564 (N_3564,N_1994,N_2865);
nand U3565 (N_3565,N_2885,N_2000);
nand U3566 (N_3566,N_2960,N_2070);
or U3567 (N_3567,N_1733,N_2728);
nand U3568 (N_3568,N_1830,N_1877);
nand U3569 (N_3569,N_1783,N_2369);
nor U3570 (N_3570,N_2748,N_2561);
or U3571 (N_3571,N_1905,N_1734);
nand U3572 (N_3572,N_2443,N_2659);
and U3573 (N_3573,N_2797,N_1915);
nor U3574 (N_3574,N_2239,N_2531);
or U3575 (N_3575,N_2493,N_2729);
or U3576 (N_3576,N_2526,N_2064);
nor U3577 (N_3577,N_2757,N_2464);
nor U3578 (N_3578,N_1631,N_2411);
and U3579 (N_3579,N_2221,N_2276);
xnor U3580 (N_3580,N_1868,N_2167);
nor U3581 (N_3581,N_1889,N_2275);
or U3582 (N_3582,N_2955,N_2588);
or U3583 (N_3583,N_1551,N_1993);
nand U3584 (N_3584,N_1967,N_2725);
and U3585 (N_3585,N_2414,N_1779);
nor U3586 (N_3586,N_2914,N_2315);
nand U3587 (N_3587,N_2340,N_2092);
and U3588 (N_3588,N_2924,N_2494);
nor U3589 (N_3589,N_2759,N_1952);
nand U3590 (N_3590,N_2111,N_1983);
and U3591 (N_3591,N_2872,N_2218);
nor U3592 (N_3592,N_2573,N_2041);
nor U3593 (N_3593,N_2918,N_2063);
nor U3594 (N_3594,N_1539,N_1702);
nor U3595 (N_3595,N_2530,N_1774);
or U3596 (N_3596,N_2105,N_1884);
nand U3597 (N_3597,N_2873,N_2142);
nand U3598 (N_3598,N_2209,N_1863);
or U3599 (N_3599,N_2617,N_1941);
nor U3600 (N_3600,N_2100,N_2037);
nand U3601 (N_3601,N_2877,N_2109);
and U3602 (N_3602,N_2528,N_1578);
or U3603 (N_3603,N_2184,N_1913);
and U3604 (N_3604,N_2698,N_1742);
and U3605 (N_3605,N_2662,N_2312);
nand U3606 (N_3606,N_1858,N_2541);
nor U3607 (N_3607,N_2773,N_2331);
and U3608 (N_3608,N_2687,N_2246);
nor U3609 (N_3609,N_2785,N_1985);
nand U3610 (N_3610,N_2585,N_2641);
and U3611 (N_3611,N_2474,N_2595);
nand U3612 (N_3612,N_2490,N_1927);
and U3613 (N_3613,N_2597,N_2354);
nand U3614 (N_3614,N_2928,N_2979);
nor U3615 (N_3615,N_2961,N_2827);
or U3616 (N_3616,N_1992,N_2065);
or U3617 (N_3617,N_2949,N_1860);
and U3618 (N_3618,N_2869,N_2887);
or U3619 (N_3619,N_1810,N_2650);
nor U3620 (N_3620,N_2640,N_1648);
or U3621 (N_3621,N_1749,N_2796);
nand U3622 (N_3622,N_2164,N_1686);
or U3623 (N_3623,N_1515,N_1693);
nand U3624 (N_3624,N_2898,N_2856);
or U3625 (N_3625,N_2673,N_1674);
nor U3626 (N_3626,N_1677,N_1954);
nand U3627 (N_3627,N_1520,N_2318);
nand U3628 (N_3628,N_2500,N_2544);
nand U3629 (N_3629,N_2085,N_2453);
and U3630 (N_3630,N_2211,N_2416);
nor U3631 (N_3631,N_2336,N_2969);
nor U3632 (N_3632,N_1647,N_1806);
nor U3633 (N_3633,N_2263,N_2888);
nand U3634 (N_3634,N_2279,N_1855);
or U3635 (N_3635,N_1558,N_2113);
and U3636 (N_3636,N_2968,N_2522);
and U3637 (N_3637,N_1826,N_1698);
or U3638 (N_3638,N_1683,N_2171);
nor U3639 (N_3639,N_2913,N_1521);
nand U3640 (N_3640,N_1934,N_2666);
nor U3641 (N_3641,N_1899,N_2029);
or U3642 (N_3642,N_2489,N_1948);
nand U3643 (N_3643,N_2228,N_1709);
or U3644 (N_3644,N_2804,N_2324);
and U3645 (N_3645,N_2598,N_1910);
or U3646 (N_3646,N_2262,N_2686);
nand U3647 (N_3647,N_2705,N_2301);
and U3648 (N_3648,N_1823,N_2248);
nand U3649 (N_3649,N_1965,N_2470);
and U3650 (N_3650,N_2451,N_1632);
and U3651 (N_3651,N_2858,N_1828);
nand U3652 (N_3652,N_2995,N_1837);
nand U3653 (N_3653,N_1789,N_1808);
or U3654 (N_3654,N_1716,N_2097);
xnor U3655 (N_3655,N_1533,N_2956);
nor U3656 (N_3656,N_2658,N_2679);
or U3657 (N_3657,N_2517,N_2782);
and U3658 (N_3658,N_1939,N_2155);
nor U3659 (N_3659,N_2117,N_2818);
nand U3660 (N_3660,N_1707,N_2933);
or U3661 (N_3661,N_2348,N_2132);
or U3662 (N_3662,N_1821,N_1554);
nand U3663 (N_3663,N_2932,N_2081);
nand U3664 (N_3664,N_2978,N_2838);
nand U3665 (N_3665,N_1615,N_2646);
or U3666 (N_3666,N_2112,N_2628);
xor U3667 (N_3667,N_1593,N_2937);
and U3668 (N_3668,N_2258,N_2480);
nand U3669 (N_3669,N_2304,N_2323);
or U3670 (N_3670,N_2572,N_1903);
nand U3671 (N_3671,N_2400,N_2558);
and U3672 (N_3672,N_1801,N_2921);
nor U3673 (N_3673,N_1845,N_1997);
nand U3674 (N_3674,N_2297,N_1561);
nand U3675 (N_3675,N_2712,N_1875);
and U3676 (N_3676,N_2104,N_1973);
or U3677 (N_3677,N_1958,N_2568);
or U3678 (N_3678,N_2513,N_2007);
or U3679 (N_3679,N_1511,N_2576);
and U3680 (N_3680,N_2945,N_2799);
and U3681 (N_3681,N_2108,N_2363);
or U3682 (N_3682,N_2379,N_2590);
nand U3683 (N_3683,N_1836,N_1758);
nand U3684 (N_3684,N_2966,N_1829);
or U3685 (N_3685,N_1986,N_2320);
or U3686 (N_3686,N_2265,N_2136);
and U3687 (N_3687,N_2039,N_2792);
nand U3688 (N_3688,N_1746,N_2433);
nand U3689 (N_3689,N_2106,N_1509);
xor U3690 (N_3690,N_2022,N_2947);
nor U3691 (N_3691,N_2594,N_2984);
nand U3692 (N_3692,N_1726,N_2479);
or U3693 (N_3693,N_2952,N_2266);
nand U3694 (N_3694,N_2477,N_2919);
xnor U3695 (N_3695,N_2399,N_2882);
nand U3696 (N_3696,N_2380,N_2904);
nand U3697 (N_3697,N_2523,N_2897);
nand U3698 (N_3698,N_2727,N_2447);
or U3699 (N_3699,N_2237,N_2618);
nand U3700 (N_3700,N_2180,N_2277);
nand U3701 (N_3701,N_1664,N_2110);
and U3702 (N_3702,N_2073,N_2099);
or U3703 (N_3703,N_2719,N_2846);
nand U3704 (N_3704,N_2971,N_2069);
nor U3705 (N_3705,N_1528,N_1769);
and U3706 (N_3706,N_2267,N_1621);
nand U3707 (N_3707,N_1906,N_2020);
nand U3708 (N_3708,N_2839,N_2574);
nand U3709 (N_3709,N_1650,N_2840);
and U3710 (N_3710,N_1581,N_2843);
nor U3711 (N_3711,N_2078,N_2637);
nand U3712 (N_3712,N_2916,N_2607);
or U3713 (N_3713,N_1754,N_1692);
nand U3714 (N_3714,N_2317,N_1685);
or U3715 (N_3715,N_2851,N_2903);
and U3716 (N_3716,N_2454,N_2146);
nand U3717 (N_3717,N_2270,N_2273);
nor U3718 (N_3718,N_2334,N_2647);
nor U3719 (N_3719,N_2219,N_2502);
and U3720 (N_3720,N_2028,N_1584);
nand U3721 (N_3721,N_1825,N_2449);
and U3722 (N_3722,N_2534,N_2730);
nand U3723 (N_3723,N_2800,N_1641);
and U3724 (N_3724,N_2700,N_2046);
and U3725 (N_3725,N_1680,N_2608);
and U3726 (N_3726,N_2622,N_1625);
and U3727 (N_3727,N_2086,N_2845);
and U3728 (N_3728,N_2139,N_2783);
or U3729 (N_3729,N_1527,N_2442);
nor U3730 (N_3730,N_2547,N_1723);
and U3731 (N_3731,N_2225,N_1984);
xnor U3732 (N_3732,N_2577,N_1820);
nand U3733 (N_3733,N_1544,N_2424);
nand U3734 (N_3734,N_1549,N_1538);
or U3735 (N_3735,N_2055,N_1689);
and U3736 (N_3736,N_2570,N_1729);
nor U3737 (N_3737,N_1532,N_1507);
nor U3738 (N_3738,N_2756,N_2810);
nand U3739 (N_3739,N_2342,N_2068);
nor U3740 (N_3740,N_2341,N_1679);
nor U3741 (N_3741,N_1999,N_1767);
nand U3742 (N_3742,N_2893,N_2886);
and U3743 (N_3743,N_2835,N_2043);
and U3744 (N_3744,N_1737,N_1567);
nor U3745 (N_3745,N_2050,N_2688);
nand U3746 (N_3746,N_2825,N_2549);
nand U3747 (N_3747,N_2004,N_2364);
nand U3748 (N_3748,N_1818,N_1885);
and U3749 (N_3749,N_2130,N_1925);
nand U3750 (N_3750,N_2096,N_2769);
or U3751 (N_3751,N_2160,N_1632);
nor U3752 (N_3752,N_2129,N_2226);
or U3753 (N_3753,N_2562,N_1964);
or U3754 (N_3754,N_2942,N_2126);
nand U3755 (N_3755,N_2790,N_1824);
or U3756 (N_3756,N_2047,N_2137);
nor U3757 (N_3757,N_1926,N_2606);
and U3758 (N_3758,N_1734,N_2074);
or U3759 (N_3759,N_2917,N_1826);
nand U3760 (N_3760,N_2297,N_2273);
or U3761 (N_3761,N_1628,N_1549);
or U3762 (N_3762,N_2252,N_2332);
nor U3763 (N_3763,N_1821,N_2754);
nand U3764 (N_3764,N_2767,N_2993);
nor U3765 (N_3765,N_1644,N_2748);
nand U3766 (N_3766,N_1762,N_2430);
nor U3767 (N_3767,N_2796,N_1535);
or U3768 (N_3768,N_2252,N_2841);
nand U3769 (N_3769,N_2577,N_1837);
nor U3770 (N_3770,N_1926,N_2052);
nand U3771 (N_3771,N_2679,N_2559);
nand U3772 (N_3772,N_1509,N_1764);
nor U3773 (N_3773,N_2415,N_2071);
nand U3774 (N_3774,N_2931,N_2073);
nand U3775 (N_3775,N_1806,N_2215);
or U3776 (N_3776,N_1767,N_2158);
and U3777 (N_3777,N_2225,N_2098);
nand U3778 (N_3778,N_2198,N_2363);
nor U3779 (N_3779,N_2602,N_1689);
and U3780 (N_3780,N_2722,N_2979);
and U3781 (N_3781,N_2074,N_2170);
or U3782 (N_3782,N_1716,N_1883);
and U3783 (N_3783,N_2955,N_1721);
nand U3784 (N_3784,N_1702,N_2422);
and U3785 (N_3785,N_2141,N_2466);
nand U3786 (N_3786,N_2380,N_2233);
nand U3787 (N_3787,N_2479,N_2905);
and U3788 (N_3788,N_1710,N_1535);
nand U3789 (N_3789,N_1720,N_1587);
and U3790 (N_3790,N_2892,N_2387);
nand U3791 (N_3791,N_1961,N_2720);
and U3792 (N_3792,N_2770,N_2788);
nor U3793 (N_3793,N_2384,N_2114);
nor U3794 (N_3794,N_1534,N_1975);
nor U3795 (N_3795,N_2134,N_2315);
and U3796 (N_3796,N_1633,N_1660);
or U3797 (N_3797,N_1790,N_1921);
and U3798 (N_3798,N_1533,N_2306);
nor U3799 (N_3799,N_1601,N_1800);
xor U3800 (N_3800,N_1914,N_2364);
or U3801 (N_3801,N_1684,N_2232);
nor U3802 (N_3802,N_1513,N_1825);
and U3803 (N_3803,N_2314,N_2766);
and U3804 (N_3804,N_1830,N_1570);
nand U3805 (N_3805,N_1640,N_2946);
nand U3806 (N_3806,N_1961,N_2129);
nand U3807 (N_3807,N_2498,N_2518);
or U3808 (N_3808,N_1671,N_1513);
and U3809 (N_3809,N_2061,N_2133);
nor U3810 (N_3810,N_2930,N_2145);
nor U3811 (N_3811,N_2619,N_2387);
or U3812 (N_3812,N_2571,N_1940);
or U3813 (N_3813,N_1974,N_1899);
nand U3814 (N_3814,N_2945,N_2994);
nand U3815 (N_3815,N_1748,N_2858);
or U3816 (N_3816,N_1507,N_2846);
or U3817 (N_3817,N_2762,N_2821);
or U3818 (N_3818,N_2316,N_2602);
and U3819 (N_3819,N_1654,N_1598);
nand U3820 (N_3820,N_2530,N_2827);
nor U3821 (N_3821,N_2733,N_2072);
or U3822 (N_3822,N_2954,N_1716);
nand U3823 (N_3823,N_2148,N_2272);
nand U3824 (N_3824,N_2340,N_2269);
nand U3825 (N_3825,N_2332,N_1878);
and U3826 (N_3826,N_2491,N_1925);
and U3827 (N_3827,N_1819,N_2376);
or U3828 (N_3828,N_1798,N_2580);
nand U3829 (N_3829,N_2820,N_1934);
or U3830 (N_3830,N_2158,N_1977);
and U3831 (N_3831,N_2218,N_1607);
nor U3832 (N_3832,N_2662,N_2934);
nand U3833 (N_3833,N_2588,N_2782);
and U3834 (N_3834,N_1995,N_1523);
and U3835 (N_3835,N_1845,N_2380);
nand U3836 (N_3836,N_2912,N_1940);
nor U3837 (N_3837,N_2496,N_2112);
or U3838 (N_3838,N_2706,N_2698);
and U3839 (N_3839,N_1787,N_2245);
and U3840 (N_3840,N_2346,N_2468);
nand U3841 (N_3841,N_1853,N_2532);
nand U3842 (N_3842,N_1836,N_2494);
and U3843 (N_3843,N_2825,N_2576);
or U3844 (N_3844,N_1914,N_2290);
or U3845 (N_3845,N_2992,N_1892);
xnor U3846 (N_3846,N_1754,N_1908);
nor U3847 (N_3847,N_1928,N_2698);
or U3848 (N_3848,N_1920,N_1785);
or U3849 (N_3849,N_2247,N_2362);
or U3850 (N_3850,N_2016,N_1547);
nand U3851 (N_3851,N_2665,N_2490);
or U3852 (N_3852,N_2464,N_2246);
and U3853 (N_3853,N_2629,N_1842);
or U3854 (N_3854,N_2520,N_1939);
xor U3855 (N_3855,N_2153,N_2686);
and U3856 (N_3856,N_1502,N_2384);
nand U3857 (N_3857,N_1839,N_2724);
nand U3858 (N_3858,N_1898,N_1627);
nor U3859 (N_3859,N_1878,N_2109);
and U3860 (N_3860,N_1759,N_2572);
nand U3861 (N_3861,N_2797,N_2065);
or U3862 (N_3862,N_2379,N_2428);
nand U3863 (N_3863,N_2910,N_2464);
or U3864 (N_3864,N_1815,N_2765);
or U3865 (N_3865,N_2077,N_2348);
and U3866 (N_3866,N_2322,N_1790);
or U3867 (N_3867,N_1569,N_2157);
or U3868 (N_3868,N_1850,N_2895);
or U3869 (N_3869,N_2406,N_1976);
or U3870 (N_3870,N_2382,N_2802);
and U3871 (N_3871,N_2704,N_2428);
nand U3872 (N_3872,N_2877,N_2046);
or U3873 (N_3873,N_2627,N_1608);
and U3874 (N_3874,N_2125,N_2054);
nand U3875 (N_3875,N_2971,N_1774);
or U3876 (N_3876,N_2772,N_2803);
nor U3877 (N_3877,N_2663,N_2769);
nand U3878 (N_3878,N_2888,N_2547);
or U3879 (N_3879,N_2658,N_2961);
and U3880 (N_3880,N_2013,N_2771);
nand U3881 (N_3881,N_2501,N_2346);
nand U3882 (N_3882,N_2550,N_2960);
or U3883 (N_3883,N_2497,N_2869);
nand U3884 (N_3884,N_2603,N_2854);
nand U3885 (N_3885,N_1807,N_1900);
or U3886 (N_3886,N_1752,N_2888);
or U3887 (N_3887,N_2030,N_2929);
and U3888 (N_3888,N_2786,N_1963);
and U3889 (N_3889,N_1713,N_2336);
and U3890 (N_3890,N_2613,N_2681);
nand U3891 (N_3891,N_2383,N_2999);
or U3892 (N_3892,N_1893,N_1841);
nand U3893 (N_3893,N_2645,N_2626);
and U3894 (N_3894,N_2218,N_2636);
nor U3895 (N_3895,N_2336,N_2420);
and U3896 (N_3896,N_1710,N_2771);
or U3897 (N_3897,N_1724,N_2436);
xnor U3898 (N_3898,N_2195,N_2500);
nor U3899 (N_3899,N_1565,N_2356);
or U3900 (N_3900,N_2910,N_2614);
or U3901 (N_3901,N_1569,N_1507);
nor U3902 (N_3902,N_2142,N_2375);
or U3903 (N_3903,N_1827,N_2242);
nand U3904 (N_3904,N_2338,N_2883);
nand U3905 (N_3905,N_1745,N_1899);
or U3906 (N_3906,N_1585,N_2694);
nor U3907 (N_3907,N_2044,N_2897);
nor U3908 (N_3908,N_2723,N_1565);
and U3909 (N_3909,N_1813,N_2737);
or U3910 (N_3910,N_2194,N_2161);
and U3911 (N_3911,N_1691,N_1823);
or U3912 (N_3912,N_1982,N_2693);
or U3913 (N_3913,N_2397,N_1519);
nand U3914 (N_3914,N_2626,N_2056);
nor U3915 (N_3915,N_2553,N_2509);
nand U3916 (N_3916,N_2200,N_1667);
nand U3917 (N_3917,N_2256,N_1649);
nand U3918 (N_3918,N_2816,N_2676);
nand U3919 (N_3919,N_1784,N_2078);
or U3920 (N_3920,N_2762,N_1740);
nor U3921 (N_3921,N_1571,N_1700);
nand U3922 (N_3922,N_2653,N_2516);
and U3923 (N_3923,N_1972,N_2466);
or U3924 (N_3924,N_2329,N_2179);
and U3925 (N_3925,N_2490,N_1661);
nor U3926 (N_3926,N_2574,N_1759);
nand U3927 (N_3927,N_2470,N_2680);
and U3928 (N_3928,N_2990,N_2918);
or U3929 (N_3929,N_1969,N_2627);
and U3930 (N_3930,N_2814,N_2939);
and U3931 (N_3931,N_2066,N_2247);
nand U3932 (N_3932,N_1925,N_2580);
and U3933 (N_3933,N_1643,N_1645);
or U3934 (N_3934,N_1932,N_2888);
or U3935 (N_3935,N_2024,N_2937);
nor U3936 (N_3936,N_1804,N_2184);
or U3937 (N_3937,N_2165,N_2205);
nand U3938 (N_3938,N_2685,N_2129);
and U3939 (N_3939,N_2704,N_1728);
nand U3940 (N_3940,N_2856,N_1898);
and U3941 (N_3941,N_2981,N_2933);
nor U3942 (N_3942,N_1650,N_2086);
nor U3943 (N_3943,N_2330,N_1605);
nand U3944 (N_3944,N_2775,N_1737);
and U3945 (N_3945,N_2783,N_2781);
and U3946 (N_3946,N_2715,N_2871);
and U3947 (N_3947,N_1905,N_1620);
and U3948 (N_3948,N_1694,N_1992);
and U3949 (N_3949,N_1730,N_2854);
or U3950 (N_3950,N_2728,N_2326);
nand U3951 (N_3951,N_2089,N_1611);
nor U3952 (N_3952,N_1815,N_2825);
nand U3953 (N_3953,N_1719,N_1893);
or U3954 (N_3954,N_2941,N_2727);
nor U3955 (N_3955,N_1866,N_2906);
or U3956 (N_3956,N_2467,N_1590);
nor U3957 (N_3957,N_2472,N_2470);
nand U3958 (N_3958,N_1754,N_2080);
nand U3959 (N_3959,N_1619,N_2084);
and U3960 (N_3960,N_2238,N_2347);
nand U3961 (N_3961,N_2025,N_1594);
and U3962 (N_3962,N_1614,N_1969);
nand U3963 (N_3963,N_1878,N_2645);
and U3964 (N_3964,N_2486,N_2979);
nand U3965 (N_3965,N_1914,N_2088);
xor U3966 (N_3966,N_1662,N_2284);
and U3967 (N_3967,N_2337,N_1676);
or U3968 (N_3968,N_1519,N_2704);
or U3969 (N_3969,N_1708,N_1903);
or U3970 (N_3970,N_1983,N_1714);
nor U3971 (N_3971,N_2763,N_1855);
or U3972 (N_3972,N_1886,N_1506);
or U3973 (N_3973,N_2516,N_2582);
and U3974 (N_3974,N_2314,N_2708);
nand U3975 (N_3975,N_1834,N_2570);
nor U3976 (N_3976,N_2296,N_2161);
nor U3977 (N_3977,N_2401,N_1875);
nor U3978 (N_3978,N_1982,N_1808);
nor U3979 (N_3979,N_2150,N_2814);
or U3980 (N_3980,N_2882,N_2951);
or U3981 (N_3981,N_2487,N_2092);
and U3982 (N_3982,N_1549,N_2751);
or U3983 (N_3983,N_1831,N_2385);
nor U3984 (N_3984,N_1714,N_1941);
and U3985 (N_3985,N_2683,N_2861);
nand U3986 (N_3986,N_2539,N_2326);
nand U3987 (N_3987,N_2901,N_2155);
or U3988 (N_3988,N_2970,N_2595);
or U3989 (N_3989,N_1906,N_2540);
nand U3990 (N_3990,N_2585,N_1951);
and U3991 (N_3991,N_1661,N_2875);
nor U3992 (N_3992,N_1658,N_2660);
nor U3993 (N_3993,N_2859,N_2562);
nand U3994 (N_3994,N_2497,N_2788);
and U3995 (N_3995,N_1772,N_1586);
nor U3996 (N_3996,N_1772,N_2197);
or U3997 (N_3997,N_2117,N_2189);
and U3998 (N_3998,N_2228,N_1648);
and U3999 (N_3999,N_1817,N_2428);
nor U4000 (N_4000,N_1773,N_1909);
and U4001 (N_4001,N_1981,N_2693);
and U4002 (N_4002,N_1620,N_1997);
nand U4003 (N_4003,N_2736,N_2214);
nand U4004 (N_4004,N_2031,N_1520);
nand U4005 (N_4005,N_2755,N_2204);
nand U4006 (N_4006,N_2694,N_2229);
or U4007 (N_4007,N_1510,N_2391);
and U4008 (N_4008,N_1896,N_2458);
nor U4009 (N_4009,N_2992,N_2918);
nand U4010 (N_4010,N_1798,N_1760);
or U4011 (N_4011,N_2831,N_1622);
and U4012 (N_4012,N_2142,N_1793);
nand U4013 (N_4013,N_2389,N_2208);
nor U4014 (N_4014,N_2437,N_2084);
nand U4015 (N_4015,N_1799,N_2562);
nor U4016 (N_4016,N_2858,N_2324);
nor U4017 (N_4017,N_2766,N_1947);
nand U4018 (N_4018,N_2995,N_2435);
nand U4019 (N_4019,N_2273,N_1573);
nor U4020 (N_4020,N_1556,N_2773);
nor U4021 (N_4021,N_2382,N_1871);
nand U4022 (N_4022,N_1986,N_1909);
and U4023 (N_4023,N_2338,N_2621);
or U4024 (N_4024,N_2938,N_1972);
and U4025 (N_4025,N_2496,N_2030);
and U4026 (N_4026,N_2770,N_2171);
nor U4027 (N_4027,N_2608,N_2297);
nand U4028 (N_4028,N_1784,N_2721);
nor U4029 (N_4029,N_2952,N_2773);
nor U4030 (N_4030,N_2908,N_2940);
and U4031 (N_4031,N_1917,N_2375);
and U4032 (N_4032,N_2980,N_2192);
or U4033 (N_4033,N_2498,N_2215);
or U4034 (N_4034,N_1736,N_2729);
or U4035 (N_4035,N_2712,N_2353);
nand U4036 (N_4036,N_1501,N_2952);
and U4037 (N_4037,N_1986,N_2789);
or U4038 (N_4038,N_2160,N_2623);
and U4039 (N_4039,N_1804,N_2665);
and U4040 (N_4040,N_2751,N_1823);
or U4041 (N_4041,N_2835,N_1540);
nand U4042 (N_4042,N_2591,N_1601);
and U4043 (N_4043,N_2238,N_2249);
nand U4044 (N_4044,N_2068,N_2442);
nor U4045 (N_4045,N_1540,N_2033);
nor U4046 (N_4046,N_1619,N_1931);
nand U4047 (N_4047,N_2177,N_1665);
nor U4048 (N_4048,N_2256,N_2459);
and U4049 (N_4049,N_2060,N_2158);
nor U4050 (N_4050,N_2481,N_2356);
nand U4051 (N_4051,N_2590,N_1516);
or U4052 (N_4052,N_2707,N_2287);
nor U4053 (N_4053,N_1656,N_1995);
and U4054 (N_4054,N_2423,N_2487);
nor U4055 (N_4055,N_2744,N_2614);
or U4056 (N_4056,N_2943,N_2778);
nand U4057 (N_4057,N_1524,N_2175);
or U4058 (N_4058,N_1896,N_2769);
and U4059 (N_4059,N_1824,N_2741);
nor U4060 (N_4060,N_2557,N_2023);
nor U4061 (N_4061,N_1524,N_1926);
or U4062 (N_4062,N_2383,N_1881);
nand U4063 (N_4063,N_2998,N_2043);
nand U4064 (N_4064,N_1923,N_2427);
nand U4065 (N_4065,N_1909,N_2134);
nor U4066 (N_4066,N_2524,N_2722);
or U4067 (N_4067,N_1700,N_1838);
and U4068 (N_4068,N_2371,N_2814);
or U4069 (N_4069,N_2929,N_1816);
nand U4070 (N_4070,N_2802,N_1533);
and U4071 (N_4071,N_2035,N_2439);
nor U4072 (N_4072,N_2944,N_2443);
or U4073 (N_4073,N_2754,N_2935);
nand U4074 (N_4074,N_1626,N_2715);
or U4075 (N_4075,N_2783,N_2061);
nand U4076 (N_4076,N_2455,N_2487);
and U4077 (N_4077,N_1616,N_1711);
and U4078 (N_4078,N_2035,N_2651);
nor U4079 (N_4079,N_1791,N_2078);
and U4080 (N_4080,N_1694,N_2156);
and U4081 (N_4081,N_2799,N_1500);
nand U4082 (N_4082,N_2689,N_2600);
and U4083 (N_4083,N_2835,N_1886);
and U4084 (N_4084,N_1586,N_1672);
and U4085 (N_4085,N_1690,N_1627);
or U4086 (N_4086,N_2004,N_2846);
and U4087 (N_4087,N_1767,N_2109);
and U4088 (N_4088,N_1778,N_2834);
and U4089 (N_4089,N_2045,N_2600);
nand U4090 (N_4090,N_2471,N_2958);
nor U4091 (N_4091,N_2445,N_1700);
nor U4092 (N_4092,N_1725,N_2145);
and U4093 (N_4093,N_2115,N_2184);
nor U4094 (N_4094,N_1528,N_1537);
or U4095 (N_4095,N_1704,N_1808);
or U4096 (N_4096,N_1791,N_1973);
and U4097 (N_4097,N_2609,N_2784);
nor U4098 (N_4098,N_1702,N_2446);
and U4099 (N_4099,N_2643,N_1767);
nand U4100 (N_4100,N_2195,N_2981);
and U4101 (N_4101,N_2490,N_2743);
nand U4102 (N_4102,N_2848,N_2532);
nand U4103 (N_4103,N_2782,N_1706);
nor U4104 (N_4104,N_2307,N_2484);
or U4105 (N_4105,N_2888,N_1567);
or U4106 (N_4106,N_2639,N_2502);
and U4107 (N_4107,N_2092,N_2544);
or U4108 (N_4108,N_2626,N_1551);
nand U4109 (N_4109,N_2292,N_2151);
or U4110 (N_4110,N_2253,N_2494);
nand U4111 (N_4111,N_2628,N_1699);
nor U4112 (N_4112,N_1832,N_1875);
nor U4113 (N_4113,N_2478,N_2395);
and U4114 (N_4114,N_2437,N_2644);
nor U4115 (N_4115,N_2327,N_2930);
nor U4116 (N_4116,N_2514,N_2038);
or U4117 (N_4117,N_1877,N_2726);
nor U4118 (N_4118,N_1562,N_1642);
and U4119 (N_4119,N_2359,N_2971);
nor U4120 (N_4120,N_1766,N_1739);
xor U4121 (N_4121,N_2850,N_2005);
or U4122 (N_4122,N_1534,N_2319);
nor U4123 (N_4123,N_2745,N_2845);
and U4124 (N_4124,N_1849,N_1546);
and U4125 (N_4125,N_1686,N_1657);
nor U4126 (N_4126,N_2792,N_2526);
nand U4127 (N_4127,N_1856,N_1727);
or U4128 (N_4128,N_1620,N_1712);
and U4129 (N_4129,N_2750,N_2829);
or U4130 (N_4130,N_2045,N_2683);
and U4131 (N_4131,N_1834,N_2573);
nand U4132 (N_4132,N_1901,N_2963);
nand U4133 (N_4133,N_2519,N_1632);
or U4134 (N_4134,N_1987,N_1745);
nor U4135 (N_4135,N_1801,N_1547);
nor U4136 (N_4136,N_1627,N_1799);
nand U4137 (N_4137,N_1541,N_1663);
nor U4138 (N_4138,N_1884,N_2774);
nor U4139 (N_4139,N_1727,N_2163);
nand U4140 (N_4140,N_1643,N_2051);
and U4141 (N_4141,N_1907,N_2487);
nand U4142 (N_4142,N_2845,N_2569);
nor U4143 (N_4143,N_2410,N_1875);
nor U4144 (N_4144,N_1790,N_2949);
and U4145 (N_4145,N_2338,N_2377);
nor U4146 (N_4146,N_2253,N_1931);
nand U4147 (N_4147,N_2964,N_2881);
nand U4148 (N_4148,N_1572,N_2917);
nor U4149 (N_4149,N_2757,N_1577);
nor U4150 (N_4150,N_2948,N_1845);
and U4151 (N_4151,N_2759,N_1696);
and U4152 (N_4152,N_2585,N_2293);
nand U4153 (N_4153,N_2294,N_1892);
nand U4154 (N_4154,N_2778,N_1998);
nand U4155 (N_4155,N_2842,N_2650);
and U4156 (N_4156,N_1558,N_1560);
or U4157 (N_4157,N_2679,N_1818);
or U4158 (N_4158,N_2106,N_2628);
xnor U4159 (N_4159,N_2314,N_2987);
or U4160 (N_4160,N_2350,N_2558);
nand U4161 (N_4161,N_1554,N_2689);
and U4162 (N_4162,N_2452,N_1767);
nand U4163 (N_4163,N_1884,N_1636);
nor U4164 (N_4164,N_2395,N_2889);
and U4165 (N_4165,N_2775,N_2193);
or U4166 (N_4166,N_2739,N_1934);
nand U4167 (N_4167,N_2074,N_2973);
or U4168 (N_4168,N_1655,N_1844);
nand U4169 (N_4169,N_2488,N_1766);
xnor U4170 (N_4170,N_2859,N_1963);
or U4171 (N_4171,N_2353,N_2976);
nand U4172 (N_4172,N_2097,N_2558);
nand U4173 (N_4173,N_1684,N_1500);
nor U4174 (N_4174,N_2601,N_2605);
nand U4175 (N_4175,N_2106,N_2154);
nand U4176 (N_4176,N_1573,N_2125);
nor U4177 (N_4177,N_2520,N_1707);
and U4178 (N_4178,N_1653,N_1560);
or U4179 (N_4179,N_2281,N_2373);
nand U4180 (N_4180,N_1837,N_1880);
and U4181 (N_4181,N_2096,N_1715);
or U4182 (N_4182,N_1847,N_2568);
and U4183 (N_4183,N_2920,N_2415);
and U4184 (N_4184,N_2626,N_1563);
and U4185 (N_4185,N_2989,N_2210);
nor U4186 (N_4186,N_2629,N_2715);
or U4187 (N_4187,N_1819,N_2698);
nor U4188 (N_4188,N_1790,N_2393);
nor U4189 (N_4189,N_1557,N_1847);
nand U4190 (N_4190,N_2784,N_2225);
nor U4191 (N_4191,N_2072,N_2530);
or U4192 (N_4192,N_1719,N_2050);
nand U4193 (N_4193,N_2437,N_2763);
or U4194 (N_4194,N_1946,N_1818);
nor U4195 (N_4195,N_1698,N_1746);
and U4196 (N_4196,N_1813,N_1665);
nor U4197 (N_4197,N_1852,N_2329);
nor U4198 (N_4198,N_1735,N_2818);
nor U4199 (N_4199,N_1942,N_1943);
and U4200 (N_4200,N_2982,N_2483);
or U4201 (N_4201,N_1533,N_2363);
nor U4202 (N_4202,N_2477,N_2456);
and U4203 (N_4203,N_1659,N_2067);
nor U4204 (N_4204,N_1926,N_1748);
nand U4205 (N_4205,N_2341,N_2448);
nor U4206 (N_4206,N_2033,N_2840);
nor U4207 (N_4207,N_2550,N_2471);
and U4208 (N_4208,N_1702,N_2477);
nand U4209 (N_4209,N_2531,N_2614);
or U4210 (N_4210,N_2137,N_1645);
or U4211 (N_4211,N_1777,N_1799);
nand U4212 (N_4212,N_2377,N_1782);
nand U4213 (N_4213,N_2480,N_2671);
and U4214 (N_4214,N_1854,N_2283);
or U4215 (N_4215,N_2894,N_2123);
nor U4216 (N_4216,N_2378,N_2257);
nor U4217 (N_4217,N_1746,N_2206);
nand U4218 (N_4218,N_2317,N_1941);
nor U4219 (N_4219,N_2815,N_2082);
and U4220 (N_4220,N_2677,N_1650);
or U4221 (N_4221,N_1645,N_2031);
nand U4222 (N_4222,N_2370,N_1915);
nor U4223 (N_4223,N_2971,N_2949);
nor U4224 (N_4224,N_2276,N_2115);
nor U4225 (N_4225,N_2552,N_2722);
nor U4226 (N_4226,N_2419,N_1664);
nor U4227 (N_4227,N_1992,N_2896);
and U4228 (N_4228,N_2966,N_2302);
nor U4229 (N_4229,N_2386,N_2774);
or U4230 (N_4230,N_2099,N_2219);
nand U4231 (N_4231,N_2829,N_2255);
and U4232 (N_4232,N_2728,N_2021);
and U4233 (N_4233,N_2110,N_2609);
and U4234 (N_4234,N_1528,N_2098);
nand U4235 (N_4235,N_1994,N_1823);
nor U4236 (N_4236,N_2906,N_1795);
nand U4237 (N_4237,N_1865,N_1947);
or U4238 (N_4238,N_2710,N_2549);
or U4239 (N_4239,N_2235,N_2930);
nor U4240 (N_4240,N_2476,N_1847);
nor U4241 (N_4241,N_2767,N_2908);
nand U4242 (N_4242,N_1769,N_2472);
nand U4243 (N_4243,N_1508,N_2311);
or U4244 (N_4244,N_2601,N_2383);
nand U4245 (N_4245,N_1742,N_1683);
and U4246 (N_4246,N_2259,N_2831);
or U4247 (N_4247,N_2924,N_2340);
or U4248 (N_4248,N_1611,N_2192);
and U4249 (N_4249,N_2821,N_2615);
nor U4250 (N_4250,N_1858,N_2786);
or U4251 (N_4251,N_2115,N_2917);
nor U4252 (N_4252,N_1711,N_1931);
or U4253 (N_4253,N_1761,N_1570);
or U4254 (N_4254,N_2867,N_2950);
or U4255 (N_4255,N_1986,N_1711);
nand U4256 (N_4256,N_1982,N_1699);
and U4257 (N_4257,N_1955,N_1867);
nor U4258 (N_4258,N_1849,N_2441);
nor U4259 (N_4259,N_2466,N_2911);
and U4260 (N_4260,N_2538,N_2600);
nor U4261 (N_4261,N_2981,N_2964);
or U4262 (N_4262,N_2470,N_2175);
nor U4263 (N_4263,N_2567,N_2102);
nor U4264 (N_4264,N_2657,N_2824);
nor U4265 (N_4265,N_1875,N_2972);
nor U4266 (N_4266,N_2495,N_2422);
and U4267 (N_4267,N_2021,N_2173);
nor U4268 (N_4268,N_1546,N_2469);
nand U4269 (N_4269,N_2798,N_2027);
nand U4270 (N_4270,N_2633,N_2092);
nor U4271 (N_4271,N_1973,N_2695);
or U4272 (N_4272,N_2053,N_1528);
nor U4273 (N_4273,N_1877,N_1564);
nor U4274 (N_4274,N_1690,N_2739);
nor U4275 (N_4275,N_2944,N_2461);
nor U4276 (N_4276,N_2685,N_2635);
or U4277 (N_4277,N_1753,N_2886);
and U4278 (N_4278,N_1593,N_1836);
and U4279 (N_4279,N_2082,N_1889);
nand U4280 (N_4280,N_2429,N_2970);
or U4281 (N_4281,N_1734,N_2169);
nand U4282 (N_4282,N_1543,N_1758);
and U4283 (N_4283,N_1623,N_2394);
nor U4284 (N_4284,N_2198,N_2396);
nand U4285 (N_4285,N_2144,N_1917);
nor U4286 (N_4286,N_2159,N_1768);
or U4287 (N_4287,N_2087,N_2966);
nor U4288 (N_4288,N_2067,N_2031);
or U4289 (N_4289,N_2256,N_1819);
nor U4290 (N_4290,N_1709,N_2987);
nor U4291 (N_4291,N_2641,N_2796);
nor U4292 (N_4292,N_2155,N_1735);
nand U4293 (N_4293,N_2795,N_2098);
xnor U4294 (N_4294,N_2383,N_1970);
nor U4295 (N_4295,N_2625,N_2436);
or U4296 (N_4296,N_2652,N_1999);
or U4297 (N_4297,N_2757,N_2326);
or U4298 (N_4298,N_2821,N_2746);
nand U4299 (N_4299,N_2477,N_2951);
or U4300 (N_4300,N_2246,N_2770);
or U4301 (N_4301,N_1861,N_2973);
and U4302 (N_4302,N_2422,N_2667);
and U4303 (N_4303,N_2559,N_2847);
or U4304 (N_4304,N_1582,N_2174);
nand U4305 (N_4305,N_2961,N_2922);
nor U4306 (N_4306,N_2690,N_1542);
or U4307 (N_4307,N_1795,N_2957);
and U4308 (N_4308,N_1875,N_1516);
and U4309 (N_4309,N_2206,N_2017);
nor U4310 (N_4310,N_1940,N_1623);
nand U4311 (N_4311,N_1516,N_2446);
nand U4312 (N_4312,N_2075,N_1635);
and U4313 (N_4313,N_2037,N_2508);
and U4314 (N_4314,N_1950,N_1790);
or U4315 (N_4315,N_2737,N_2341);
and U4316 (N_4316,N_1627,N_1805);
nand U4317 (N_4317,N_1811,N_2556);
or U4318 (N_4318,N_1574,N_1823);
nor U4319 (N_4319,N_2458,N_2028);
nor U4320 (N_4320,N_2581,N_1570);
nor U4321 (N_4321,N_2592,N_2172);
xor U4322 (N_4322,N_1539,N_2232);
or U4323 (N_4323,N_2375,N_2510);
nand U4324 (N_4324,N_2283,N_2928);
nor U4325 (N_4325,N_2585,N_2138);
and U4326 (N_4326,N_2549,N_1656);
or U4327 (N_4327,N_1961,N_2459);
or U4328 (N_4328,N_2741,N_2750);
or U4329 (N_4329,N_2300,N_2694);
and U4330 (N_4330,N_2165,N_2750);
or U4331 (N_4331,N_2250,N_2063);
or U4332 (N_4332,N_2620,N_1753);
or U4333 (N_4333,N_2760,N_1789);
nor U4334 (N_4334,N_1972,N_2965);
nand U4335 (N_4335,N_2449,N_1870);
xor U4336 (N_4336,N_2134,N_2331);
nand U4337 (N_4337,N_2010,N_2479);
and U4338 (N_4338,N_2744,N_1632);
and U4339 (N_4339,N_1718,N_2917);
or U4340 (N_4340,N_1806,N_1762);
nor U4341 (N_4341,N_2876,N_2257);
nor U4342 (N_4342,N_2525,N_2547);
or U4343 (N_4343,N_2205,N_2523);
and U4344 (N_4344,N_1597,N_2013);
and U4345 (N_4345,N_1980,N_1919);
nor U4346 (N_4346,N_2680,N_2907);
nand U4347 (N_4347,N_1933,N_2835);
and U4348 (N_4348,N_2166,N_2464);
or U4349 (N_4349,N_2994,N_2915);
nand U4350 (N_4350,N_2928,N_2611);
nor U4351 (N_4351,N_2529,N_1802);
nand U4352 (N_4352,N_2371,N_2023);
and U4353 (N_4353,N_1883,N_2035);
or U4354 (N_4354,N_1699,N_2361);
nand U4355 (N_4355,N_2643,N_2980);
nand U4356 (N_4356,N_1995,N_1824);
nor U4357 (N_4357,N_2646,N_2263);
nor U4358 (N_4358,N_1978,N_2936);
nand U4359 (N_4359,N_1919,N_1839);
or U4360 (N_4360,N_1598,N_2116);
nand U4361 (N_4361,N_2118,N_2486);
and U4362 (N_4362,N_2588,N_2546);
nand U4363 (N_4363,N_2095,N_2104);
or U4364 (N_4364,N_2134,N_2875);
or U4365 (N_4365,N_2405,N_2970);
and U4366 (N_4366,N_2419,N_2465);
or U4367 (N_4367,N_1666,N_2753);
nand U4368 (N_4368,N_2869,N_2277);
or U4369 (N_4369,N_1514,N_2767);
or U4370 (N_4370,N_2909,N_2996);
nand U4371 (N_4371,N_1697,N_2772);
and U4372 (N_4372,N_2574,N_2722);
or U4373 (N_4373,N_1836,N_2005);
or U4374 (N_4374,N_2065,N_2664);
or U4375 (N_4375,N_2776,N_1821);
or U4376 (N_4376,N_2636,N_2906);
nor U4377 (N_4377,N_2458,N_2777);
nor U4378 (N_4378,N_2373,N_2819);
or U4379 (N_4379,N_2615,N_1714);
or U4380 (N_4380,N_2490,N_2047);
and U4381 (N_4381,N_1740,N_2781);
or U4382 (N_4382,N_2137,N_2806);
or U4383 (N_4383,N_1978,N_2999);
or U4384 (N_4384,N_1777,N_2144);
and U4385 (N_4385,N_2643,N_2079);
or U4386 (N_4386,N_1957,N_2233);
nand U4387 (N_4387,N_1778,N_2966);
and U4388 (N_4388,N_2764,N_2947);
nand U4389 (N_4389,N_1948,N_2897);
or U4390 (N_4390,N_2796,N_1715);
or U4391 (N_4391,N_2837,N_2773);
nor U4392 (N_4392,N_1819,N_2764);
or U4393 (N_4393,N_2545,N_1782);
nand U4394 (N_4394,N_2903,N_2556);
nand U4395 (N_4395,N_1606,N_2053);
nor U4396 (N_4396,N_2026,N_2934);
nor U4397 (N_4397,N_1971,N_2159);
and U4398 (N_4398,N_2086,N_2363);
nor U4399 (N_4399,N_2282,N_1940);
and U4400 (N_4400,N_1761,N_2527);
or U4401 (N_4401,N_2962,N_1841);
nand U4402 (N_4402,N_2807,N_1656);
or U4403 (N_4403,N_2899,N_2684);
and U4404 (N_4404,N_2695,N_2903);
nand U4405 (N_4405,N_2566,N_2433);
nor U4406 (N_4406,N_2746,N_1723);
or U4407 (N_4407,N_1921,N_2172);
or U4408 (N_4408,N_2876,N_2849);
nand U4409 (N_4409,N_1537,N_1832);
and U4410 (N_4410,N_2370,N_1882);
or U4411 (N_4411,N_1667,N_2213);
nand U4412 (N_4412,N_1742,N_1861);
or U4413 (N_4413,N_2713,N_2602);
nor U4414 (N_4414,N_2485,N_2802);
and U4415 (N_4415,N_2907,N_2288);
and U4416 (N_4416,N_2940,N_1850);
nand U4417 (N_4417,N_2759,N_2387);
or U4418 (N_4418,N_2062,N_2869);
or U4419 (N_4419,N_2712,N_1504);
nand U4420 (N_4420,N_2730,N_1548);
nor U4421 (N_4421,N_1823,N_1762);
nand U4422 (N_4422,N_1963,N_2805);
nand U4423 (N_4423,N_2471,N_1850);
nor U4424 (N_4424,N_2794,N_2805);
or U4425 (N_4425,N_1969,N_2510);
or U4426 (N_4426,N_2140,N_2493);
and U4427 (N_4427,N_2279,N_1937);
nand U4428 (N_4428,N_2987,N_1672);
and U4429 (N_4429,N_2017,N_2863);
and U4430 (N_4430,N_2905,N_2911);
nand U4431 (N_4431,N_2168,N_2209);
nor U4432 (N_4432,N_2291,N_2138);
or U4433 (N_4433,N_2124,N_2064);
and U4434 (N_4434,N_2755,N_2265);
nor U4435 (N_4435,N_2591,N_1531);
nor U4436 (N_4436,N_2818,N_2446);
or U4437 (N_4437,N_2545,N_2504);
or U4438 (N_4438,N_2666,N_2643);
nand U4439 (N_4439,N_2213,N_2589);
and U4440 (N_4440,N_1978,N_2521);
nor U4441 (N_4441,N_2830,N_2969);
and U4442 (N_4442,N_2514,N_1647);
nor U4443 (N_4443,N_2176,N_2891);
or U4444 (N_4444,N_2833,N_2906);
and U4445 (N_4445,N_2259,N_1894);
or U4446 (N_4446,N_2000,N_2949);
nor U4447 (N_4447,N_1747,N_2021);
nor U4448 (N_4448,N_2662,N_2184);
nor U4449 (N_4449,N_1503,N_2128);
nor U4450 (N_4450,N_1865,N_1563);
nand U4451 (N_4451,N_2157,N_2014);
or U4452 (N_4452,N_1566,N_2101);
nor U4453 (N_4453,N_2597,N_2206);
nor U4454 (N_4454,N_2194,N_2286);
or U4455 (N_4455,N_1953,N_1724);
nor U4456 (N_4456,N_1670,N_2247);
nor U4457 (N_4457,N_1859,N_2752);
and U4458 (N_4458,N_2696,N_2094);
or U4459 (N_4459,N_2075,N_2398);
nand U4460 (N_4460,N_1713,N_1636);
and U4461 (N_4461,N_2059,N_2277);
and U4462 (N_4462,N_2084,N_1578);
and U4463 (N_4463,N_1551,N_2901);
nand U4464 (N_4464,N_2180,N_1774);
nand U4465 (N_4465,N_2638,N_2291);
nand U4466 (N_4466,N_2105,N_2989);
and U4467 (N_4467,N_1813,N_2673);
or U4468 (N_4468,N_2062,N_1639);
nor U4469 (N_4469,N_2345,N_2979);
or U4470 (N_4470,N_2464,N_2274);
or U4471 (N_4471,N_2561,N_2003);
and U4472 (N_4472,N_2650,N_1723);
nand U4473 (N_4473,N_2914,N_2200);
or U4474 (N_4474,N_2285,N_2011);
or U4475 (N_4475,N_2184,N_1570);
and U4476 (N_4476,N_2588,N_1657);
or U4477 (N_4477,N_1695,N_2563);
nand U4478 (N_4478,N_2240,N_2222);
nor U4479 (N_4479,N_2834,N_2697);
or U4480 (N_4480,N_2321,N_2428);
nor U4481 (N_4481,N_1636,N_2402);
and U4482 (N_4482,N_2404,N_1666);
or U4483 (N_4483,N_2001,N_1528);
or U4484 (N_4484,N_2820,N_1625);
and U4485 (N_4485,N_1870,N_2426);
and U4486 (N_4486,N_2214,N_1852);
or U4487 (N_4487,N_1695,N_2997);
or U4488 (N_4488,N_1782,N_2819);
nor U4489 (N_4489,N_2452,N_2889);
nand U4490 (N_4490,N_1897,N_2937);
and U4491 (N_4491,N_2262,N_2877);
nand U4492 (N_4492,N_2733,N_2495);
nor U4493 (N_4493,N_1509,N_2914);
nor U4494 (N_4494,N_2817,N_2091);
nor U4495 (N_4495,N_2221,N_1891);
and U4496 (N_4496,N_2408,N_1926);
nor U4497 (N_4497,N_2009,N_1930);
nor U4498 (N_4498,N_1574,N_2411);
nor U4499 (N_4499,N_2776,N_2634);
and U4500 (N_4500,N_4419,N_3132);
nor U4501 (N_4501,N_4336,N_4048);
or U4502 (N_4502,N_3846,N_4100);
nor U4503 (N_4503,N_3813,N_3504);
or U4504 (N_4504,N_4272,N_3304);
and U4505 (N_4505,N_4080,N_4201);
or U4506 (N_4506,N_4489,N_4179);
nand U4507 (N_4507,N_3855,N_3752);
and U4508 (N_4508,N_3699,N_3391);
or U4509 (N_4509,N_4408,N_3117);
nand U4510 (N_4510,N_3259,N_3448);
nand U4511 (N_4511,N_4289,N_4233);
nor U4512 (N_4512,N_4112,N_3785);
xnor U4513 (N_4513,N_4183,N_3232);
nor U4514 (N_4514,N_4440,N_3640);
and U4515 (N_4515,N_3339,N_3289);
and U4516 (N_4516,N_3500,N_3493);
nor U4517 (N_4517,N_4007,N_3853);
and U4518 (N_4518,N_3960,N_4095);
or U4519 (N_4519,N_3756,N_4089);
nor U4520 (N_4520,N_4180,N_3608);
or U4521 (N_4521,N_4137,N_3318);
nand U4522 (N_4522,N_4287,N_3422);
and U4523 (N_4523,N_3193,N_3476);
or U4524 (N_4524,N_3187,N_4451);
and U4525 (N_4525,N_3793,N_4315);
and U4526 (N_4526,N_3256,N_4471);
or U4527 (N_4527,N_4278,N_4010);
and U4528 (N_4528,N_3874,N_4204);
nand U4529 (N_4529,N_3868,N_3225);
nor U4530 (N_4530,N_4017,N_3305);
nand U4531 (N_4531,N_3989,N_3200);
or U4532 (N_4532,N_4295,N_3085);
nor U4533 (N_4533,N_3170,N_4317);
or U4534 (N_4534,N_3636,N_3769);
or U4535 (N_4535,N_3890,N_3303);
or U4536 (N_4536,N_4014,N_3114);
nor U4537 (N_4537,N_3521,N_3815);
or U4538 (N_4538,N_3691,N_3996);
or U4539 (N_4539,N_3045,N_3923);
nand U4540 (N_4540,N_4141,N_3204);
or U4541 (N_4541,N_3872,N_3933);
nor U4542 (N_4542,N_3899,N_3341);
nor U4543 (N_4543,N_3244,N_3127);
or U4544 (N_4544,N_3362,N_3760);
nor U4545 (N_4545,N_3551,N_3441);
or U4546 (N_4546,N_3430,N_3490);
or U4547 (N_4547,N_3743,N_4426);
and U4548 (N_4548,N_3198,N_3638);
or U4549 (N_4549,N_4243,N_3069);
and U4550 (N_4550,N_4125,N_3345);
or U4551 (N_4551,N_4105,N_4199);
nand U4552 (N_4552,N_3633,N_3028);
and U4553 (N_4553,N_3566,N_4165);
nand U4554 (N_4554,N_4396,N_4088);
and U4555 (N_4555,N_3434,N_4118);
and U4556 (N_4556,N_4351,N_3829);
nor U4557 (N_4557,N_3029,N_4312);
nor U4558 (N_4558,N_3964,N_3724);
and U4559 (N_4559,N_4005,N_4032);
and U4560 (N_4560,N_3316,N_3147);
xnor U4561 (N_4561,N_3860,N_4044);
nand U4562 (N_4562,N_3040,N_3678);
nand U4563 (N_4563,N_3781,N_3352);
nand U4564 (N_4564,N_4457,N_3650);
nand U4565 (N_4565,N_4172,N_3817);
nand U4566 (N_4566,N_3308,N_4239);
and U4567 (N_4567,N_4423,N_3035);
or U4568 (N_4568,N_3292,N_3767);
or U4569 (N_4569,N_3115,N_3419);
nor U4570 (N_4570,N_3892,N_4358);
or U4571 (N_4571,N_4027,N_4302);
nand U4572 (N_4572,N_4355,N_3988);
and U4573 (N_4573,N_3524,N_4499);
nor U4574 (N_4574,N_4217,N_3651);
nor U4575 (N_4575,N_4194,N_4380);
or U4576 (N_4576,N_3424,N_4225);
xnor U4577 (N_4577,N_3428,N_3830);
or U4578 (N_4578,N_3930,N_4365);
nand U4579 (N_4579,N_3264,N_3841);
or U4580 (N_4580,N_3639,N_4131);
nand U4581 (N_4581,N_3677,N_4348);
xor U4582 (N_4582,N_3795,N_3119);
nand U4583 (N_4583,N_3942,N_4122);
or U4584 (N_4584,N_4349,N_3983);
nor U4585 (N_4585,N_3060,N_3062);
or U4586 (N_4586,N_3263,N_4364);
and U4587 (N_4587,N_3528,N_3843);
or U4588 (N_4588,N_3690,N_4393);
or U4589 (N_4589,N_3751,N_4218);
nor U4590 (N_4590,N_4448,N_3408);
and U4591 (N_4591,N_3873,N_3245);
and U4592 (N_4592,N_3274,N_3826);
or U4593 (N_4593,N_3291,N_4447);
nand U4594 (N_4594,N_3050,N_4421);
and U4595 (N_4595,N_3759,N_3597);
and U4596 (N_4596,N_4142,N_4258);
or U4597 (N_4597,N_3734,N_3038);
nand U4598 (N_4598,N_3722,N_3552);
or U4599 (N_4599,N_3842,N_3859);
and U4600 (N_4600,N_3057,N_3265);
or U4601 (N_4601,N_3415,N_3661);
nand U4602 (N_4602,N_3918,N_3295);
nor U4603 (N_4603,N_4437,N_3164);
nor U4604 (N_4604,N_4110,N_3852);
nand U4605 (N_4605,N_4203,N_4427);
nor U4606 (N_4606,N_4024,N_3664);
nand U4607 (N_4607,N_3380,N_3461);
nor U4608 (N_4608,N_3113,N_3189);
or U4609 (N_4609,N_3014,N_3705);
or U4610 (N_4610,N_3741,N_3203);
nand U4611 (N_4611,N_3550,N_3511);
and U4612 (N_4612,N_3103,N_4164);
nand U4613 (N_4613,N_3272,N_4022);
nand U4614 (N_4614,N_4046,N_3703);
nand U4615 (N_4615,N_3354,N_3966);
or U4616 (N_4616,N_3994,N_3465);
nand U4617 (N_4617,N_4316,N_3788);
or U4618 (N_4618,N_3590,N_3235);
or U4619 (N_4619,N_3181,N_3747);
nand U4620 (N_4620,N_3655,N_4453);
or U4621 (N_4621,N_4397,N_3510);
and U4622 (N_4622,N_3483,N_3279);
or U4623 (N_4623,N_3680,N_3701);
nor U4624 (N_4624,N_3665,N_4309);
or U4625 (N_4625,N_3484,N_4151);
nor U4626 (N_4626,N_4280,N_4401);
nand U4627 (N_4627,N_4111,N_3594);
nand U4628 (N_4628,N_3471,N_3418);
nor U4629 (N_4629,N_3220,N_3142);
nand U4630 (N_4630,N_3513,N_4033);
nand U4631 (N_4631,N_4381,N_4439);
and U4632 (N_4632,N_4049,N_3248);
or U4633 (N_4633,N_3392,N_3820);
nor U4634 (N_4634,N_3451,N_3086);
nand U4635 (N_4635,N_3152,N_3499);
nand U4636 (N_4636,N_3887,N_3586);
nand U4637 (N_4637,N_3439,N_3588);
nand U4638 (N_4638,N_3692,N_4284);
and U4639 (N_4639,N_4023,N_3658);
nor U4640 (N_4640,N_4050,N_4353);
and U4641 (N_4641,N_4256,N_4410);
nand U4642 (N_4642,N_3782,N_3911);
and U4643 (N_4643,N_3628,N_4436);
nand U4644 (N_4644,N_4238,N_4124);
nand U4645 (N_4645,N_3541,N_3267);
or U4646 (N_4646,N_3812,N_3847);
nand U4647 (N_4647,N_4188,N_3076);
nand U4648 (N_4648,N_4488,N_4308);
and U4649 (N_4649,N_3575,N_4159);
or U4650 (N_4650,N_3877,N_3459);
or U4651 (N_4651,N_3669,N_4412);
nand U4652 (N_4652,N_3672,N_4175);
or U4653 (N_4653,N_4301,N_4113);
and U4654 (N_4654,N_3311,N_3634);
or U4655 (N_4655,N_3931,N_3378);
nor U4656 (N_4656,N_3704,N_4285);
nand U4657 (N_4657,N_3631,N_3044);
nor U4658 (N_4658,N_3831,N_3643);
nor U4659 (N_4659,N_4341,N_3405);
nor U4660 (N_4660,N_3112,N_3998);
and U4661 (N_4661,N_4246,N_4433);
nor U4662 (N_4662,N_4260,N_4297);
or U4663 (N_4663,N_3713,N_3188);
or U4664 (N_4664,N_4407,N_4347);
or U4665 (N_4665,N_4454,N_4094);
or U4666 (N_4666,N_3410,N_3218);
nor U4667 (N_4667,N_3178,N_4461);
nand U4668 (N_4668,N_4445,N_3675);
and U4669 (N_4669,N_3128,N_3130);
or U4670 (N_4670,N_4187,N_4229);
and U4671 (N_4671,N_3558,N_3236);
or U4672 (N_4672,N_3824,N_3294);
nand U4673 (N_4673,N_3938,N_3034);
and U4674 (N_4674,N_3126,N_3070);
nor U4675 (N_4675,N_3231,N_3221);
xor U4676 (N_4676,N_4378,N_3241);
nor U4677 (N_4677,N_3089,N_3963);
nor U4678 (N_4678,N_4098,N_4102);
or U4679 (N_4679,N_3977,N_3753);
nor U4680 (N_4680,N_4265,N_4126);
or U4681 (N_4681,N_3290,N_4495);
nor U4682 (N_4682,N_3326,N_3275);
nor U4683 (N_4683,N_4452,N_3102);
nor U4684 (N_4684,N_4372,N_3041);
and U4685 (N_4685,N_3526,N_3239);
or U4686 (N_4686,N_3803,N_3323);
nor U4687 (N_4687,N_3001,N_4063);
or U4688 (N_4688,N_3844,N_3058);
nor U4689 (N_4689,N_4011,N_3023);
or U4690 (N_4690,N_3601,N_4376);
and U4691 (N_4691,N_3965,N_3440);
nand U4692 (N_4692,N_4300,N_4228);
nor U4693 (N_4693,N_3652,N_4162);
xnor U4694 (N_4694,N_3973,N_3331);
and U4695 (N_4695,N_3093,N_3412);
and U4696 (N_4696,N_3561,N_3100);
or U4697 (N_4697,N_3488,N_3941);
or U4698 (N_4698,N_3794,N_3920);
or U4699 (N_4699,N_3425,N_3662);
or U4700 (N_4700,N_4181,N_4266);
nand U4701 (N_4701,N_3017,N_3547);
and U4702 (N_4702,N_4039,N_3576);
nand U4703 (N_4703,N_3962,N_3924);
nand U4704 (N_4704,N_3463,N_3689);
nor U4705 (N_4705,N_4000,N_3879);
or U4706 (N_4706,N_3196,N_3968);
and U4707 (N_4707,N_4076,N_3325);
nand U4708 (N_4708,N_4134,N_3446);
nand U4709 (N_4709,N_3007,N_3288);
nor U4710 (N_4710,N_4171,N_3162);
nand U4711 (N_4711,N_3123,N_3447);
or U4712 (N_4712,N_3061,N_4288);
nor U4713 (N_4713,N_3516,N_3230);
nand U4714 (N_4714,N_4192,N_3522);
or U4715 (N_4715,N_3632,N_3255);
and U4716 (N_4716,N_3525,N_4320);
nand U4717 (N_4717,N_3388,N_3568);
and U4718 (N_4718,N_3377,N_4087);
nand U4719 (N_4719,N_3287,N_3833);
or U4720 (N_4720,N_4209,N_3875);
or U4721 (N_4721,N_3736,N_3997);
and U4722 (N_4722,N_4160,N_4486);
nand U4723 (N_4723,N_4369,N_3611);
and U4724 (N_4724,N_3771,N_3224);
xor U4725 (N_4725,N_3674,N_3067);
and U4726 (N_4726,N_4374,N_3420);
and U4727 (N_4727,N_3937,N_3957);
nand U4728 (N_4728,N_4082,N_3613);
or U4729 (N_4729,N_3618,N_3984);
or U4730 (N_4730,N_4247,N_3624);
nor U4731 (N_4731,N_3240,N_4186);
or U4732 (N_4732,N_3811,N_4252);
or U4733 (N_4733,N_3138,N_3518);
and U4734 (N_4734,N_3124,N_4475);
nor U4735 (N_4735,N_3464,N_4020);
or U4736 (N_4736,N_4059,N_3022);
nor U4737 (N_4737,N_4425,N_4335);
nand U4738 (N_4738,N_3864,N_3312);
or U4739 (N_4739,N_4222,N_4117);
and U4740 (N_4740,N_3506,N_3012);
nor U4741 (N_4741,N_4240,N_3083);
or U4742 (N_4742,N_4104,N_3533);
nor U4743 (N_4743,N_3851,N_4158);
and U4744 (N_4744,N_3592,N_3357);
nand U4745 (N_4745,N_3133,N_3940);
nand U4746 (N_4746,N_3945,N_3545);
and U4747 (N_4747,N_3072,N_3489);
and U4748 (N_4748,N_4148,N_4323);
or U4749 (N_4749,N_3258,N_4399);
or U4750 (N_4750,N_4479,N_3438);
nor U4751 (N_4751,N_3000,N_3149);
or U4752 (N_4752,N_3066,N_4206);
nor U4753 (N_4753,N_4394,N_3542);
or U4754 (N_4754,N_3252,N_4176);
nand U4755 (N_4755,N_3399,N_3637);
nand U4756 (N_4756,N_3707,N_3314);
and U4757 (N_4757,N_3109,N_3695);
nand U4758 (N_4758,N_4443,N_3137);
nand U4759 (N_4759,N_3955,N_3792);
nand U4760 (N_4760,N_3554,N_4115);
nor U4761 (N_4761,N_4208,N_3881);
nand U4762 (N_4762,N_3144,N_3726);
nand U4763 (N_4763,N_3698,N_3626);
or U4764 (N_4764,N_4235,N_3498);
or U4765 (N_4765,N_4119,N_3182);
and U4766 (N_4766,N_4325,N_4262);
nand U4767 (N_4767,N_4200,N_4168);
nand U4768 (N_4768,N_3171,N_3049);
nor U4769 (N_4769,N_3177,N_4483);
nor U4770 (N_4770,N_4371,N_3298);
and U4771 (N_4771,N_3565,N_3789);
nand U4772 (N_4772,N_3927,N_3816);
and U4773 (N_4773,N_3729,N_3219);
nor U4774 (N_4774,N_4136,N_3491);
nor U4775 (N_4775,N_3578,N_4268);
and U4776 (N_4776,N_3612,N_3514);
nor U4777 (N_4777,N_3379,N_3043);
nor U4778 (N_4778,N_4304,N_4129);
and U4779 (N_4779,N_3208,N_4339);
and U4780 (N_4780,N_3926,N_3384);
or U4781 (N_4781,N_3074,N_4485);
and U4782 (N_4782,N_3416,N_4491);
and U4783 (N_4783,N_3591,N_3835);
or U4784 (N_4784,N_4001,N_4153);
or U4785 (N_4785,N_3358,N_3990);
nand U4786 (N_4786,N_3361,N_3175);
nor U4787 (N_4787,N_3770,N_3478);
and U4788 (N_4788,N_3981,N_3906);
nor U4789 (N_4789,N_3088,N_4496);
nor U4790 (N_4790,N_3281,N_4074);
xnor U4791 (N_4791,N_3078,N_4191);
xor U4792 (N_4792,N_3260,N_3596);
or U4793 (N_4793,N_3229,N_4460);
and U4794 (N_4794,N_3082,N_3912);
nand U4795 (N_4795,N_4382,N_3394);
nor U4796 (N_4796,N_4464,N_3807);
nor U4797 (N_4797,N_4038,N_3036);
and U4798 (N_4798,N_4404,N_3199);
nor U4799 (N_4799,N_4429,N_4071);
and U4800 (N_4800,N_4478,N_3914);
nor U4801 (N_4801,N_3237,N_3913);
and U4802 (N_4802,N_3950,N_3366);
and U4803 (N_4803,N_3810,N_4361);
and U4804 (N_4804,N_3808,N_4254);
or U4805 (N_4805,N_4259,N_3494);
or U4806 (N_4806,N_4362,N_3694);
and U4807 (N_4807,N_3156,N_4455);
or U4808 (N_4808,N_4169,N_3742);
nor U4809 (N_4809,N_3008,N_3856);
or U4810 (N_4810,N_3242,N_3444);
and U4811 (N_4811,N_4498,N_3186);
nand U4812 (N_4812,N_3897,N_3839);
nand U4813 (N_4813,N_3857,N_4146);
nand U4814 (N_4814,N_3978,N_4279);
or U4815 (N_4815,N_3627,N_4242);
and U4816 (N_4816,N_3185,N_3688);
and U4817 (N_4817,N_3143,N_4065);
or U4818 (N_4818,N_3935,N_3139);
nor U4819 (N_4819,N_3540,N_3850);
and U4820 (N_4820,N_3276,N_3939);
nand U4821 (N_4821,N_3584,N_3991);
or U4822 (N_4822,N_3861,N_4356);
and U4823 (N_4823,N_3470,N_3167);
xnor U4824 (N_4824,N_3140,N_4311);
xor U4825 (N_4825,N_3387,N_4008);
nor U4826 (N_4826,N_3324,N_4043);
or U4827 (N_4827,N_3902,N_4350);
or U4828 (N_4828,N_4400,N_3891);
or U4829 (N_4829,N_3414,N_3825);
or U4830 (N_4830,N_3687,N_3865);
and U4831 (N_4831,N_3556,N_3667);
and U4832 (N_4832,N_3262,N_3779);
or U4833 (N_4833,N_3383,N_3548);
nor U4834 (N_4834,N_3567,N_3423);
nand U4835 (N_4835,N_3953,N_4154);
nand U4836 (N_4836,N_3025,N_4366);
or U4837 (N_4837,N_3297,N_3075);
or U4838 (N_4838,N_3740,N_4092);
and U4839 (N_4839,N_3016,N_3363);
nor U4840 (N_4840,N_4469,N_3602);
nor U4841 (N_4841,N_3531,N_4294);
nand U4842 (N_4842,N_4013,N_4422);
nor U4843 (N_4843,N_3786,N_3959);
or U4844 (N_4844,N_4081,N_4281);
and U4845 (N_4845,N_4167,N_4255);
nor U4846 (N_4846,N_4178,N_3762);
and U4847 (N_4847,N_4054,N_3046);
nand U4848 (N_4848,N_3212,N_3348);
nand U4849 (N_4849,N_4249,N_3917);
and U4850 (N_4850,N_4428,N_4416);
nand U4851 (N_4851,N_3335,N_3595);
and U4852 (N_4852,N_4047,N_3227);
nor U4853 (N_4853,N_4058,N_3557);
or U4854 (N_4854,N_3581,N_4096);
nor U4855 (N_4855,N_3614,N_3630);
or U4856 (N_4856,N_3954,N_3365);
and U4857 (N_4857,N_3179,N_4147);
and U4858 (N_4858,N_4352,N_3150);
nand U4859 (N_4859,N_3328,N_3319);
nand U4860 (N_4860,N_4232,N_3195);
or U4861 (N_4861,N_4324,N_3870);
and U4862 (N_4862,N_3160,N_4389);
or U4863 (N_4863,N_4212,N_3355);
or U4864 (N_4864,N_3059,N_4403);
and U4865 (N_4865,N_3985,N_4140);
nor U4866 (N_4866,N_3758,N_3359);
or U4867 (N_4867,N_3697,N_3895);
nand U4868 (N_4868,N_3822,N_4097);
nor U4869 (N_4869,N_3725,N_3166);
nor U4870 (N_4870,N_4431,N_4414);
nand U4871 (N_4871,N_4387,N_3976);
or U4872 (N_4872,N_3159,N_3055);
and U4873 (N_4873,N_3190,N_4484);
nor U4874 (N_4874,N_4251,N_3503);
nand U4875 (N_4875,N_4045,N_3460);
xor U4876 (N_4876,N_4286,N_4012);
or U4877 (N_4877,N_3334,N_4318);
or U4878 (N_4878,N_3944,N_4036);
or U4879 (N_4879,N_3313,N_4342);
nand U4880 (N_4880,N_3153,N_3572);
or U4881 (N_4881,N_3909,N_4101);
or U4882 (N_4882,N_3684,N_3700);
nor U4883 (N_4883,N_3823,N_3322);
and U4884 (N_4884,N_3623,N_3535);
nor U4885 (N_4885,N_3589,N_4090);
nand U4886 (N_4886,N_3080,N_3834);
nor U4887 (N_4887,N_3037,N_3712);
and U4888 (N_4888,N_4133,N_3982);
or U4889 (N_4889,N_4120,N_3949);
nand U4890 (N_4890,N_4482,N_4003);
and U4891 (N_4891,N_3191,N_3342);
nor U4892 (N_4892,N_3723,N_4337);
nor U4893 (N_4893,N_3520,N_4213);
nand U4894 (N_4894,N_3819,N_4185);
nor U4895 (N_4895,N_3610,N_4220);
and U4896 (N_4896,N_4073,N_3641);
nor U4897 (N_4897,N_4373,N_3709);
nor U4898 (N_4898,N_3946,N_3411);
nor U4899 (N_4899,N_3071,N_4487);
nor U4900 (N_4900,N_3407,N_3105);
and U4901 (N_4901,N_3893,N_3745);
nand U4902 (N_4902,N_3336,N_3719);
and U4903 (N_4903,N_3475,N_4306);
xor U4904 (N_4904,N_3226,N_4329);
or U4905 (N_4905,N_3249,N_3009);
nor U4906 (N_4906,N_4490,N_4215);
nand U4907 (N_4907,N_3508,N_3748);
and U4908 (N_4908,N_3099,N_4170);
nor U4909 (N_4909,N_3356,N_3901);
or U4910 (N_4910,N_4221,N_3398);
nand U4911 (N_4911,N_4025,N_3457);
and U4912 (N_4912,N_3777,N_3993);
and U4913 (N_4913,N_4377,N_3282);
or U4914 (N_4914,N_3992,N_4331);
nand U4915 (N_4915,N_3527,N_4424);
and U4916 (N_4916,N_3517,N_3869);
and U4917 (N_4917,N_4420,N_3098);
and U4918 (N_4918,N_3970,N_3395);
nor U4919 (N_4919,N_3453,N_4405);
or U4920 (N_4920,N_3858,N_3546);
and U4921 (N_4921,N_4360,N_3791);
xnor U4922 (N_4922,N_3209,N_4211);
nand U4923 (N_4923,N_3286,N_3136);
nor U4924 (N_4924,N_4042,N_3376);
nor U4925 (N_4925,N_3573,N_3577);
and U4926 (N_4926,N_3878,N_3215);
nor U4927 (N_4927,N_4357,N_3797);
and U4928 (N_4928,N_3727,N_3400);
and U4929 (N_4929,N_3593,N_4277);
nor U4930 (N_4930,N_4273,N_4132);
nand U4931 (N_4931,N_3337,N_3660);
nor U4932 (N_4932,N_3176,N_3682);
nor U4933 (N_4933,N_3763,N_4413);
nor U4934 (N_4934,N_3888,N_3784);
nand U4935 (N_4935,N_3375,N_4383);
nand U4936 (N_4936,N_4450,N_4015);
nand U4937 (N_4937,N_3733,N_3169);
nor U4938 (N_4938,N_4345,N_3327);
or U4939 (N_4939,N_3766,N_3299);
nand U4940 (N_4940,N_4415,N_3481);
and U4941 (N_4941,N_4016,N_3452);
and U4942 (N_4942,N_4468,N_3466);
nand U4943 (N_4943,N_3668,N_3644);
nand U4944 (N_4944,N_4114,N_4283);
or U4945 (N_4945,N_4072,N_3011);
nand U4946 (N_4946,N_3539,N_3894);
or U4947 (N_4947,N_3673,N_4236);
or U4948 (N_4948,N_4152,N_3523);
or U4949 (N_4949,N_4034,N_3353);
nor U4950 (N_4950,N_4079,N_3403);
and U4951 (N_4951,N_3192,N_3987);
or U4952 (N_4952,N_3961,N_3333);
and U4953 (N_4953,N_3670,N_3505);
and U4954 (N_4954,N_3800,N_3307);
or U4955 (N_4955,N_3486,N_3302);
or U4956 (N_4956,N_3211,N_3848);
nor U4957 (N_4957,N_3537,N_3549);
or U4958 (N_4958,N_3617,N_4121);
nor U4959 (N_4959,N_3467,N_4106);
or U4960 (N_4960,N_3271,N_3721);
nand U4961 (N_4961,N_3530,N_3479);
and U4962 (N_4962,N_3402,N_3431);
and U4963 (N_4963,N_3735,N_4275);
nor U4964 (N_4964,N_4150,N_3880);
nand U4965 (N_4965,N_3714,N_4476);
or U4966 (N_4966,N_3110,N_3645);
nand U4967 (N_4967,N_4149,N_4248);
or U4968 (N_4968,N_3396,N_3730);
and U4969 (N_4969,N_3801,N_4019);
nor U4970 (N_4970,N_3210,N_4354);
and U4971 (N_4971,N_4313,N_3340);
nor U4972 (N_4972,N_3296,N_4481);
or U4973 (N_4973,N_3223,N_3051);
or U4974 (N_4974,N_3562,N_3228);
or U4975 (N_4975,N_3889,N_4333);
or U4976 (N_4976,N_3158,N_3417);
nand U4977 (N_4977,N_3474,N_3019);
and U4978 (N_4978,N_3429,N_3956);
nand U4979 (N_4979,N_4363,N_3473);
nand U4980 (N_4980,N_4182,N_4321);
nand U4981 (N_4981,N_4002,N_4472);
nand U4982 (N_4982,N_3936,N_4359);
nand U4983 (N_4983,N_3197,N_3389);
nand U4984 (N_4984,N_3183,N_4161);
or U4985 (N_4985,N_3129,N_3174);
and U4986 (N_4986,N_3948,N_4305);
xnor U4987 (N_4987,N_4230,N_3246);
and U4988 (N_4988,N_3269,N_3635);
nand U4989 (N_4989,N_4497,N_3625);
nor U4990 (N_4990,N_3585,N_3980);
or U4991 (N_4991,N_4298,N_3092);
and U4992 (N_4992,N_3739,N_4270);
and U4993 (N_4993,N_4474,N_3656);
nand U4994 (N_4994,N_3148,N_3773);
and U4995 (N_4995,N_3679,N_3497);
or U4996 (N_4996,N_4040,N_3253);
nand U4997 (N_4997,N_3696,N_3409);
nor U4998 (N_4998,N_4292,N_3172);
or U4999 (N_4999,N_4030,N_3047);
nand U5000 (N_5000,N_3350,N_3373);
nand U5001 (N_5001,N_3905,N_4234);
nor U5002 (N_5002,N_3718,N_4216);
and U5003 (N_5003,N_3986,N_3943);
or U5004 (N_5004,N_4282,N_3922);
and U5005 (N_5005,N_3809,N_3681);
or U5006 (N_5006,N_3840,N_3828);
and U5007 (N_5007,N_4057,N_4332);
or U5008 (N_5008,N_4367,N_3107);
nor U5009 (N_5009,N_4322,N_3238);
or U5010 (N_5010,N_3344,N_3659);
nand U5011 (N_5011,N_3202,N_3031);
or U5012 (N_5012,N_3455,N_3543);
or U5013 (N_5013,N_4099,N_3580);
nor U5014 (N_5014,N_3437,N_4330);
nand U5015 (N_5015,N_3744,N_3571);
nand U5016 (N_5016,N_4402,N_3343);
and U5017 (N_5017,N_4271,N_4031);
nand U5018 (N_5018,N_4174,N_4069);
and U5019 (N_5019,N_3649,N_3056);
nor U5020 (N_5020,N_4386,N_3884);
nand U5021 (N_5021,N_3754,N_4205);
nand U5022 (N_5022,N_3780,N_4346);
or U5023 (N_5023,N_4430,N_4061);
nor U5024 (N_5024,N_3151,N_4466);
nor U5025 (N_5025,N_4409,N_4214);
and U5026 (N_5026,N_3154,N_3774);
or U5027 (N_5027,N_4257,N_3555);
and U5028 (N_5028,N_3432,N_3406);
or U5029 (N_5029,N_3134,N_4173);
and U5030 (N_5030,N_3710,N_3932);
nor U5031 (N_5031,N_4210,N_3761);
or U5032 (N_5032,N_4319,N_3720);
or U5033 (N_5033,N_3755,N_3073);
xor U5034 (N_5034,N_4261,N_3910);
nand U5035 (N_5035,N_3600,N_4128);
nor U5036 (N_5036,N_3765,N_3250);
nand U5037 (N_5037,N_3146,N_3832);
nor U5038 (N_5038,N_3663,N_3283);
or U5039 (N_5039,N_3097,N_4223);
and U5040 (N_5040,N_3728,N_4145);
and U5041 (N_5041,N_3449,N_3605);
and U5042 (N_5042,N_3386,N_4029);
and U5043 (N_5043,N_3750,N_4276);
and U5044 (N_5044,N_3309,N_4290);
and U5045 (N_5045,N_3079,N_4411);
nor U5046 (N_5046,N_4156,N_4467);
nor U5047 (N_5047,N_3671,N_3374);
or U5048 (N_5048,N_3629,N_3908);
nor U5049 (N_5049,N_4130,N_4052);
nor U5050 (N_5050,N_3849,N_3268);
nand U5051 (N_5051,N_3234,N_3118);
and U5052 (N_5052,N_3032,N_3024);
and U5053 (N_5053,N_4006,N_3347);
or U5054 (N_5054,N_3442,N_3896);
and U5055 (N_5055,N_3737,N_4463);
or U5056 (N_5056,N_3921,N_3827);
and U5057 (N_5057,N_3974,N_3845);
and U5058 (N_5058,N_4334,N_4338);
or U5059 (N_5059,N_3496,N_3052);
or U5060 (N_5060,N_3141,N_3426);
or U5061 (N_5061,N_3207,N_4068);
and U5062 (N_5062,N_3999,N_4028);
nand U5063 (N_5063,N_4231,N_3574);
nor U5064 (N_5064,N_3806,N_3004);
nor U5065 (N_5065,N_3278,N_3653);
and U5066 (N_5066,N_3157,N_3609);
and U5067 (N_5067,N_4135,N_4103);
and U5068 (N_5068,N_4462,N_3958);
and U5069 (N_5069,N_4108,N_3135);
and U5070 (N_5070,N_3603,N_3018);
nand U5071 (N_5071,N_3213,N_4473);
nand U5072 (N_5072,N_3915,N_3900);
or U5073 (N_5073,N_4055,N_3091);
or U5074 (N_5074,N_3607,N_3757);
nor U5075 (N_5075,N_4184,N_4458);
or U5076 (N_5076,N_4237,N_3201);
nor U5077 (N_5077,N_3952,N_3972);
nor U5078 (N_5078,N_3615,N_3427);
and U5079 (N_5079,N_3372,N_3370);
xnor U5080 (N_5080,N_4195,N_3616);
and U5081 (N_5081,N_3005,N_3120);
nor U5082 (N_5082,N_3064,N_3553);
nand U5083 (N_5083,N_4143,N_3717);
and U5084 (N_5084,N_3106,N_4303);
nand U5085 (N_5085,N_3686,N_3838);
nand U5086 (N_5086,N_4018,N_4144);
nand U5087 (N_5087,N_3338,N_3155);
nand U5088 (N_5088,N_4465,N_3096);
nor U5089 (N_5089,N_3243,N_3646);
nand U5090 (N_5090,N_3764,N_3364);
and U5091 (N_5091,N_3205,N_3746);
or U5092 (N_5092,N_3020,N_3916);
and U5093 (N_5093,N_3802,N_3251);
nor U5094 (N_5094,N_3560,N_3310);
nor U5095 (N_5095,N_3544,N_3015);
nor U5096 (N_5096,N_3598,N_3648);
nor U5097 (N_5097,N_3951,N_3413);
or U5098 (N_5098,N_3676,N_4456);
xnor U5099 (N_5099,N_4196,N_4435);
nand U5100 (N_5100,N_3480,N_3329);
xor U5101 (N_5101,N_4398,N_4327);
or U5102 (N_5102,N_3502,N_3622);
nand U5103 (N_5103,N_3928,N_3804);
and U5104 (N_5104,N_3693,N_3620);
or U5105 (N_5105,N_4091,N_3979);
and U5106 (N_5106,N_3975,N_3796);
and U5107 (N_5107,N_4340,N_3222);
nand U5108 (N_5108,N_3163,N_3854);
or U5109 (N_5109,N_3898,N_3529);
and U5110 (N_5110,N_4064,N_4343);
nor U5111 (N_5111,N_3995,N_3711);
or U5112 (N_5112,N_3772,N_3495);
and U5113 (N_5113,N_4155,N_3382);
nor U5114 (N_5114,N_3125,N_4449);
or U5115 (N_5115,N_4245,N_3450);
and U5116 (N_5116,N_4391,N_3006);
nor U5117 (N_5117,N_4224,N_3090);
and U5118 (N_5118,N_4470,N_4078);
nand U5119 (N_5119,N_3487,N_3716);
nand U5120 (N_5120,N_3749,N_4241);
nand U5121 (N_5121,N_4384,N_3882);
and U5122 (N_5122,N_4189,N_3485);
nand U5123 (N_5123,N_3161,N_4441);
nor U5124 (N_5124,N_3702,N_3512);
nand U5125 (N_5125,N_3919,N_4227);
or U5126 (N_5126,N_3084,N_4392);
and U5127 (N_5127,N_3469,N_4190);
and U5128 (N_5128,N_4314,N_3371);
and U5129 (N_5129,N_4444,N_3346);
or U5130 (N_5130,N_3715,N_3101);
and U5131 (N_5131,N_3277,N_3925);
and U5132 (N_5132,N_3805,N_3534);
nor U5133 (N_5133,N_3087,N_4056);
and U5134 (N_5134,N_3194,N_3837);
nor U5135 (N_5135,N_4062,N_4123);
or U5136 (N_5136,N_4026,N_4084);
and U5137 (N_5137,N_3708,N_3436);
nand U5138 (N_5138,N_3116,N_3732);
or U5139 (N_5139,N_3042,N_3217);
and U5140 (N_5140,N_3731,N_3818);
nand U5141 (N_5141,N_3472,N_3569);
or U5142 (N_5142,N_4035,N_4274);
or U5143 (N_5143,N_3907,N_3317);
nand U5144 (N_5144,N_3002,N_3257);
nand U5145 (N_5145,N_4163,N_4067);
and U5146 (N_5146,N_4197,N_3969);
nand U5147 (N_5147,N_3783,N_3738);
or U5148 (N_5148,N_3033,N_3583);
and U5149 (N_5149,N_4093,N_3108);
and U5150 (N_5150,N_4202,N_3081);
or U5151 (N_5151,N_3273,N_3515);
and U5152 (N_5152,N_3104,N_3180);
and U5153 (N_5153,N_3862,N_3967);
nand U5154 (N_5154,N_4244,N_4066);
and U5155 (N_5155,N_3404,N_4418);
nor U5156 (N_5156,N_4219,N_3619);
and U5157 (N_5157,N_3330,N_3393);
and U5158 (N_5158,N_3706,N_4021);
or U5159 (N_5159,N_4139,N_4494);
and U5160 (N_5160,N_4253,N_3492);
nand U5161 (N_5161,N_4492,N_3360);
and U5162 (N_5162,N_3443,N_3564);
nand U5163 (N_5163,N_3368,N_3165);
and U5164 (N_5164,N_3145,N_3863);
or U5165 (N_5165,N_3814,N_4432);
nor U5166 (N_5166,N_4390,N_4075);
nor U5167 (N_5167,N_3095,N_4070);
and U5168 (N_5168,N_3883,N_3871);
and U5169 (N_5169,N_3509,N_3519);
and U5170 (N_5170,N_3604,N_3021);
nand U5171 (N_5171,N_4388,N_3886);
or U5172 (N_5172,N_3349,N_3876);
and U5173 (N_5173,N_4085,N_4060);
or U5174 (N_5174,N_3435,N_3285);
and U5175 (N_5175,N_4310,N_3013);
or U5176 (N_5176,N_3501,N_3027);
nor U5177 (N_5177,N_3657,N_3026);
and U5178 (N_5178,N_3903,N_3599);
nor U5179 (N_5179,N_4138,N_4299);
nand U5180 (N_5180,N_3666,N_4477);
and U5181 (N_5181,N_3261,N_3321);
nor U5182 (N_5182,N_4379,N_4041);
or U5183 (N_5183,N_4250,N_3454);
nor U5184 (N_5184,N_4291,N_4083);
and U5185 (N_5185,N_3683,N_3111);
or U5186 (N_5186,N_3790,N_4385);
nor U5187 (N_5187,N_4177,N_3184);
or U5188 (N_5188,N_4004,N_4263);
nor U5189 (N_5189,N_4434,N_3206);
nor U5190 (N_5190,N_4264,N_3233);
or U5191 (N_5191,N_3532,N_3214);
nand U5192 (N_5192,N_4480,N_4493);
nor U5193 (N_5193,N_3866,N_3971);
or U5194 (N_5194,N_4375,N_3867);
nor U5195 (N_5195,N_3775,N_3536);
or U5196 (N_5196,N_4370,N_3768);
and U5197 (N_5197,N_3010,N_3003);
nand U5198 (N_5198,N_3482,N_4127);
and U5199 (N_5199,N_4326,N_4198);
nor U5200 (N_5200,N_4107,N_3885);
nor U5201 (N_5201,N_3929,N_3385);
and U5202 (N_5202,N_3094,N_3122);
and U5203 (N_5203,N_4307,N_3381);
and U5204 (N_5204,N_3433,N_3685);
and U5205 (N_5205,N_4053,N_3173);
or U5206 (N_5206,N_3445,N_3401);
nand U5207 (N_5207,N_4269,N_4368);
and U5208 (N_5208,N_3284,N_3077);
and U5209 (N_5209,N_3647,N_3934);
or U5210 (N_5210,N_3270,N_3559);
or U5211 (N_5211,N_3247,N_3216);
nand U5212 (N_5212,N_3563,N_3642);
nor U5213 (N_5213,N_3351,N_3587);
and U5214 (N_5214,N_4051,N_3280);
xor U5215 (N_5215,N_3367,N_3538);
and U5216 (N_5216,N_3048,N_3121);
nand U5217 (N_5217,N_3332,N_3320);
and U5218 (N_5218,N_4109,N_4077);
nand U5219 (N_5219,N_3582,N_3606);
and U5220 (N_5220,N_4438,N_3168);
and U5221 (N_5221,N_3306,N_3579);
nand U5222 (N_5222,N_3131,N_4406);
and U5223 (N_5223,N_3477,N_4207);
nor U5224 (N_5224,N_4459,N_4037);
or U5225 (N_5225,N_3798,N_4226);
or U5226 (N_5226,N_3301,N_3507);
nand U5227 (N_5227,N_3293,N_3054);
and U5228 (N_5228,N_3787,N_3621);
or U5229 (N_5229,N_4417,N_3570);
nor U5230 (N_5230,N_3458,N_3369);
nor U5231 (N_5231,N_4395,N_3821);
or U5232 (N_5232,N_4446,N_4086);
or U5233 (N_5233,N_3776,N_4328);
and U5234 (N_5234,N_3254,N_4267);
and U5235 (N_5235,N_4116,N_3421);
nand U5236 (N_5236,N_3315,N_3654);
and U5237 (N_5237,N_4442,N_4293);
or U5238 (N_5238,N_3065,N_3068);
and U5239 (N_5239,N_3456,N_3063);
and U5240 (N_5240,N_3462,N_3397);
nand U5241 (N_5241,N_4166,N_3300);
nor U5242 (N_5242,N_3947,N_3266);
nand U5243 (N_5243,N_3030,N_4009);
nor U5244 (N_5244,N_3904,N_4296);
and U5245 (N_5245,N_3053,N_4344);
nor U5246 (N_5246,N_3778,N_4157);
nor U5247 (N_5247,N_3468,N_3799);
nor U5248 (N_5248,N_3836,N_3039);
nor U5249 (N_5249,N_3390,N_4193);
and U5250 (N_5250,N_4020,N_3363);
nand U5251 (N_5251,N_3949,N_4363);
nand U5252 (N_5252,N_3728,N_3847);
or U5253 (N_5253,N_3893,N_4440);
nand U5254 (N_5254,N_3903,N_3896);
nand U5255 (N_5255,N_4422,N_4100);
nor U5256 (N_5256,N_3765,N_3598);
nand U5257 (N_5257,N_3391,N_3964);
nand U5258 (N_5258,N_4253,N_3328);
nor U5259 (N_5259,N_4151,N_3103);
and U5260 (N_5260,N_3637,N_4094);
and U5261 (N_5261,N_4299,N_4239);
and U5262 (N_5262,N_3024,N_3453);
xnor U5263 (N_5263,N_3769,N_3522);
and U5264 (N_5264,N_3282,N_3868);
nand U5265 (N_5265,N_4140,N_3057);
nor U5266 (N_5266,N_3142,N_4164);
or U5267 (N_5267,N_3466,N_4448);
and U5268 (N_5268,N_4280,N_3184);
nand U5269 (N_5269,N_3421,N_4309);
and U5270 (N_5270,N_4229,N_3078);
nor U5271 (N_5271,N_3132,N_3426);
or U5272 (N_5272,N_4148,N_3550);
nand U5273 (N_5273,N_3946,N_3068);
or U5274 (N_5274,N_4481,N_3810);
nand U5275 (N_5275,N_3006,N_4067);
and U5276 (N_5276,N_4368,N_3163);
nor U5277 (N_5277,N_3292,N_3654);
or U5278 (N_5278,N_3249,N_3304);
and U5279 (N_5279,N_4129,N_3042);
nor U5280 (N_5280,N_4345,N_3902);
or U5281 (N_5281,N_3453,N_3059);
and U5282 (N_5282,N_3464,N_3428);
nor U5283 (N_5283,N_3807,N_3165);
nor U5284 (N_5284,N_4083,N_3100);
nand U5285 (N_5285,N_3820,N_3067);
nor U5286 (N_5286,N_4062,N_3522);
nor U5287 (N_5287,N_3837,N_3726);
or U5288 (N_5288,N_3967,N_3310);
nor U5289 (N_5289,N_3522,N_4021);
xor U5290 (N_5290,N_3259,N_3220);
or U5291 (N_5291,N_3072,N_3106);
nor U5292 (N_5292,N_3079,N_4112);
and U5293 (N_5293,N_3873,N_4207);
and U5294 (N_5294,N_3513,N_3930);
xnor U5295 (N_5295,N_4202,N_3144);
nor U5296 (N_5296,N_3691,N_3582);
nand U5297 (N_5297,N_3093,N_3474);
and U5298 (N_5298,N_4357,N_3960);
nand U5299 (N_5299,N_4395,N_3616);
and U5300 (N_5300,N_3981,N_3038);
or U5301 (N_5301,N_3883,N_3703);
nor U5302 (N_5302,N_3390,N_3010);
nor U5303 (N_5303,N_3728,N_3621);
nand U5304 (N_5304,N_3472,N_3387);
xor U5305 (N_5305,N_4414,N_4179);
and U5306 (N_5306,N_4004,N_3236);
or U5307 (N_5307,N_3298,N_3905);
nor U5308 (N_5308,N_4472,N_3720);
and U5309 (N_5309,N_4298,N_3556);
or U5310 (N_5310,N_3093,N_4336);
or U5311 (N_5311,N_3383,N_3883);
or U5312 (N_5312,N_4118,N_4246);
and U5313 (N_5313,N_4213,N_4438);
and U5314 (N_5314,N_4016,N_3333);
and U5315 (N_5315,N_4154,N_3364);
nor U5316 (N_5316,N_3943,N_3405);
nand U5317 (N_5317,N_4476,N_3293);
or U5318 (N_5318,N_3429,N_3271);
nand U5319 (N_5319,N_3253,N_3403);
and U5320 (N_5320,N_3766,N_3078);
and U5321 (N_5321,N_3136,N_4440);
or U5322 (N_5322,N_3558,N_4061);
or U5323 (N_5323,N_4238,N_3838);
nor U5324 (N_5324,N_3453,N_3738);
nand U5325 (N_5325,N_4056,N_3625);
nor U5326 (N_5326,N_4414,N_4186);
nor U5327 (N_5327,N_4488,N_3168);
nand U5328 (N_5328,N_3984,N_4293);
or U5329 (N_5329,N_3767,N_3725);
or U5330 (N_5330,N_4169,N_3639);
and U5331 (N_5331,N_3390,N_3645);
and U5332 (N_5332,N_3392,N_3344);
and U5333 (N_5333,N_3666,N_3579);
nor U5334 (N_5334,N_4284,N_3000);
nor U5335 (N_5335,N_4196,N_3407);
or U5336 (N_5336,N_3464,N_3936);
nand U5337 (N_5337,N_3901,N_3237);
or U5338 (N_5338,N_4478,N_3724);
and U5339 (N_5339,N_4146,N_4133);
and U5340 (N_5340,N_3439,N_4202);
nand U5341 (N_5341,N_3063,N_3962);
and U5342 (N_5342,N_3088,N_3040);
nor U5343 (N_5343,N_3666,N_4220);
or U5344 (N_5344,N_4058,N_3045);
nor U5345 (N_5345,N_4290,N_3289);
nand U5346 (N_5346,N_4328,N_4071);
or U5347 (N_5347,N_3274,N_3877);
nand U5348 (N_5348,N_3751,N_4204);
and U5349 (N_5349,N_4090,N_3059);
or U5350 (N_5350,N_3122,N_3688);
nor U5351 (N_5351,N_3625,N_3017);
or U5352 (N_5352,N_4347,N_4146);
and U5353 (N_5353,N_4213,N_3084);
and U5354 (N_5354,N_3276,N_3134);
and U5355 (N_5355,N_4331,N_3550);
and U5356 (N_5356,N_3848,N_3765);
nand U5357 (N_5357,N_4111,N_4487);
or U5358 (N_5358,N_4460,N_4216);
or U5359 (N_5359,N_3925,N_4190);
nand U5360 (N_5360,N_3702,N_4473);
or U5361 (N_5361,N_3476,N_3738);
and U5362 (N_5362,N_4088,N_4107);
nand U5363 (N_5363,N_3514,N_4201);
or U5364 (N_5364,N_3246,N_4012);
and U5365 (N_5365,N_3077,N_3025);
nand U5366 (N_5366,N_3769,N_3104);
nor U5367 (N_5367,N_4135,N_3363);
and U5368 (N_5368,N_3241,N_3631);
nor U5369 (N_5369,N_4215,N_4131);
and U5370 (N_5370,N_4145,N_3851);
and U5371 (N_5371,N_3825,N_4117);
or U5372 (N_5372,N_4059,N_3942);
nor U5373 (N_5373,N_3141,N_3961);
and U5374 (N_5374,N_4482,N_4110);
nor U5375 (N_5375,N_4181,N_3151);
nand U5376 (N_5376,N_3896,N_4324);
nand U5377 (N_5377,N_3576,N_3857);
or U5378 (N_5378,N_3030,N_4324);
nand U5379 (N_5379,N_4214,N_4237);
and U5380 (N_5380,N_3131,N_3872);
nand U5381 (N_5381,N_3544,N_3745);
and U5382 (N_5382,N_3834,N_3200);
or U5383 (N_5383,N_3900,N_3466);
and U5384 (N_5384,N_3389,N_3118);
nand U5385 (N_5385,N_4258,N_4184);
nor U5386 (N_5386,N_4177,N_4320);
or U5387 (N_5387,N_3898,N_4422);
and U5388 (N_5388,N_4008,N_3149);
nor U5389 (N_5389,N_4360,N_3205);
or U5390 (N_5390,N_3667,N_4459);
nor U5391 (N_5391,N_3602,N_3353);
or U5392 (N_5392,N_3331,N_3176);
and U5393 (N_5393,N_3359,N_3570);
or U5394 (N_5394,N_3174,N_3387);
and U5395 (N_5395,N_3684,N_3198);
or U5396 (N_5396,N_3565,N_3747);
nor U5397 (N_5397,N_3869,N_3846);
nand U5398 (N_5398,N_3372,N_3363);
and U5399 (N_5399,N_3157,N_4294);
nand U5400 (N_5400,N_4053,N_4085);
nand U5401 (N_5401,N_3490,N_3386);
nor U5402 (N_5402,N_4409,N_3129);
and U5403 (N_5403,N_3142,N_3647);
nor U5404 (N_5404,N_4468,N_3535);
nand U5405 (N_5405,N_3981,N_3497);
or U5406 (N_5406,N_3638,N_4231);
nor U5407 (N_5407,N_3879,N_3251);
nor U5408 (N_5408,N_3824,N_3213);
or U5409 (N_5409,N_4143,N_3920);
or U5410 (N_5410,N_3609,N_3775);
nor U5411 (N_5411,N_4427,N_3921);
or U5412 (N_5412,N_3944,N_4120);
or U5413 (N_5413,N_3934,N_3228);
and U5414 (N_5414,N_4027,N_4409);
or U5415 (N_5415,N_3433,N_3565);
or U5416 (N_5416,N_3448,N_3033);
nor U5417 (N_5417,N_3340,N_3333);
or U5418 (N_5418,N_3721,N_3407);
or U5419 (N_5419,N_3756,N_3357);
and U5420 (N_5420,N_4041,N_3387);
nor U5421 (N_5421,N_4037,N_4187);
nand U5422 (N_5422,N_3566,N_4067);
and U5423 (N_5423,N_4190,N_3223);
or U5424 (N_5424,N_3378,N_3023);
and U5425 (N_5425,N_3133,N_3434);
nand U5426 (N_5426,N_4432,N_3807);
nand U5427 (N_5427,N_3494,N_4376);
nand U5428 (N_5428,N_3344,N_4077);
and U5429 (N_5429,N_4070,N_3695);
nand U5430 (N_5430,N_3276,N_4119);
and U5431 (N_5431,N_3542,N_3652);
nor U5432 (N_5432,N_4411,N_3252);
and U5433 (N_5433,N_3094,N_3943);
nand U5434 (N_5434,N_3880,N_3245);
nor U5435 (N_5435,N_4464,N_3762);
and U5436 (N_5436,N_3032,N_3549);
or U5437 (N_5437,N_3992,N_3763);
or U5438 (N_5438,N_3191,N_3492);
nor U5439 (N_5439,N_3631,N_4277);
and U5440 (N_5440,N_4487,N_4271);
nand U5441 (N_5441,N_4165,N_3644);
and U5442 (N_5442,N_4245,N_4477);
nor U5443 (N_5443,N_3466,N_3027);
or U5444 (N_5444,N_4463,N_4240);
and U5445 (N_5445,N_3006,N_4296);
or U5446 (N_5446,N_3174,N_4486);
nor U5447 (N_5447,N_4129,N_3406);
nor U5448 (N_5448,N_3763,N_3341);
or U5449 (N_5449,N_3396,N_3415);
nor U5450 (N_5450,N_3387,N_3858);
or U5451 (N_5451,N_3215,N_4408);
and U5452 (N_5452,N_3914,N_4466);
nor U5453 (N_5453,N_3069,N_3604);
or U5454 (N_5454,N_3893,N_3814);
and U5455 (N_5455,N_4487,N_4378);
or U5456 (N_5456,N_3454,N_4498);
nor U5457 (N_5457,N_3227,N_3976);
nor U5458 (N_5458,N_3469,N_3520);
and U5459 (N_5459,N_3649,N_4133);
or U5460 (N_5460,N_4334,N_3391);
nor U5461 (N_5461,N_3489,N_3685);
nand U5462 (N_5462,N_3000,N_3681);
or U5463 (N_5463,N_3705,N_4024);
or U5464 (N_5464,N_3899,N_3121);
and U5465 (N_5465,N_3938,N_3809);
and U5466 (N_5466,N_3051,N_4088);
nor U5467 (N_5467,N_3504,N_4058);
nand U5468 (N_5468,N_3579,N_3805);
and U5469 (N_5469,N_4289,N_3700);
or U5470 (N_5470,N_4320,N_4378);
nor U5471 (N_5471,N_3327,N_3673);
and U5472 (N_5472,N_3237,N_3069);
and U5473 (N_5473,N_3387,N_4067);
and U5474 (N_5474,N_3580,N_3001);
nor U5475 (N_5475,N_3278,N_4361);
nand U5476 (N_5476,N_3174,N_4437);
or U5477 (N_5477,N_3493,N_3040);
nand U5478 (N_5478,N_4493,N_3683);
xnor U5479 (N_5479,N_3076,N_4216);
nand U5480 (N_5480,N_3918,N_3933);
nor U5481 (N_5481,N_4414,N_3520);
or U5482 (N_5482,N_4047,N_3279);
nand U5483 (N_5483,N_3100,N_3174);
nand U5484 (N_5484,N_3448,N_3580);
and U5485 (N_5485,N_3833,N_3781);
or U5486 (N_5486,N_4163,N_3872);
nor U5487 (N_5487,N_3492,N_3522);
xor U5488 (N_5488,N_3253,N_3471);
nand U5489 (N_5489,N_3355,N_3025);
xor U5490 (N_5490,N_3114,N_4108);
xor U5491 (N_5491,N_4400,N_3288);
or U5492 (N_5492,N_3377,N_3885);
nor U5493 (N_5493,N_3356,N_3180);
nand U5494 (N_5494,N_3660,N_3691);
nor U5495 (N_5495,N_3966,N_3438);
nor U5496 (N_5496,N_3714,N_3925);
nor U5497 (N_5497,N_3166,N_3821);
or U5498 (N_5498,N_4039,N_4071);
or U5499 (N_5499,N_3480,N_3724);
nand U5500 (N_5500,N_3231,N_3555);
or U5501 (N_5501,N_3859,N_3161);
nor U5502 (N_5502,N_4395,N_4105);
nor U5503 (N_5503,N_4365,N_3649);
and U5504 (N_5504,N_3226,N_4300);
nand U5505 (N_5505,N_3441,N_4183);
nor U5506 (N_5506,N_3709,N_3784);
or U5507 (N_5507,N_4328,N_4014);
or U5508 (N_5508,N_3473,N_3874);
nor U5509 (N_5509,N_4163,N_3032);
nand U5510 (N_5510,N_3559,N_3052);
nand U5511 (N_5511,N_4040,N_3635);
nor U5512 (N_5512,N_3146,N_4129);
or U5513 (N_5513,N_4141,N_3298);
nor U5514 (N_5514,N_3537,N_3566);
nand U5515 (N_5515,N_3876,N_4370);
and U5516 (N_5516,N_4062,N_4445);
and U5517 (N_5517,N_4066,N_3057);
and U5518 (N_5518,N_3116,N_3128);
nand U5519 (N_5519,N_3654,N_3566);
nand U5520 (N_5520,N_4298,N_4244);
nand U5521 (N_5521,N_3868,N_4211);
and U5522 (N_5522,N_3137,N_4184);
nor U5523 (N_5523,N_4063,N_3808);
and U5524 (N_5524,N_3132,N_3007);
nor U5525 (N_5525,N_4080,N_3990);
or U5526 (N_5526,N_3703,N_3858);
and U5527 (N_5527,N_3654,N_4410);
nor U5528 (N_5528,N_3801,N_3877);
or U5529 (N_5529,N_3513,N_4427);
or U5530 (N_5530,N_3718,N_3707);
and U5531 (N_5531,N_3526,N_4385);
and U5532 (N_5532,N_3860,N_3168);
nor U5533 (N_5533,N_3180,N_3476);
nor U5534 (N_5534,N_4244,N_3517);
nor U5535 (N_5535,N_4256,N_4040);
nor U5536 (N_5536,N_3977,N_3673);
and U5537 (N_5537,N_4063,N_4300);
and U5538 (N_5538,N_3027,N_4110);
and U5539 (N_5539,N_3154,N_3276);
or U5540 (N_5540,N_3593,N_4004);
and U5541 (N_5541,N_3929,N_4270);
nand U5542 (N_5542,N_3034,N_3192);
nor U5543 (N_5543,N_3006,N_4410);
nand U5544 (N_5544,N_3635,N_4439);
nand U5545 (N_5545,N_3398,N_3578);
and U5546 (N_5546,N_3420,N_3878);
nand U5547 (N_5547,N_3007,N_4141);
and U5548 (N_5548,N_3689,N_3973);
nand U5549 (N_5549,N_3352,N_3570);
nand U5550 (N_5550,N_4107,N_4217);
nand U5551 (N_5551,N_3255,N_3062);
nor U5552 (N_5552,N_3651,N_3621);
nand U5553 (N_5553,N_4071,N_3888);
or U5554 (N_5554,N_4047,N_4358);
nor U5555 (N_5555,N_4183,N_4043);
nor U5556 (N_5556,N_4081,N_4446);
or U5557 (N_5557,N_4271,N_3842);
and U5558 (N_5558,N_4291,N_3271);
and U5559 (N_5559,N_3740,N_3215);
or U5560 (N_5560,N_3136,N_3303);
nor U5561 (N_5561,N_3970,N_4353);
and U5562 (N_5562,N_3230,N_3537);
or U5563 (N_5563,N_3794,N_3191);
and U5564 (N_5564,N_3678,N_4118);
or U5565 (N_5565,N_4010,N_4213);
or U5566 (N_5566,N_4026,N_3937);
nand U5567 (N_5567,N_4088,N_3226);
or U5568 (N_5568,N_3400,N_4239);
and U5569 (N_5569,N_4078,N_4213);
nor U5570 (N_5570,N_3372,N_3933);
nand U5571 (N_5571,N_4244,N_3054);
nor U5572 (N_5572,N_4071,N_3838);
and U5573 (N_5573,N_4384,N_3718);
nand U5574 (N_5574,N_3794,N_4164);
and U5575 (N_5575,N_4137,N_3268);
nor U5576 (N_5576,N_3690,N_3025);
and U5577 (N_5577,N_4049,N_4425);
nand U5578 (N_5578,N_4328,N_4253);
and U5579 (N_5579,N_4493,N_3058);
nor U5580 (N_5580,N_3832,N_3293);
and U5581 (N_5581,N_4485,N_4332);
and U5582 (N_5582,N_3577,N_3435);
nand U5583 (N_5583,N_3551,N_3236);
and U5584 (N_5584,N_3043,N_4003);
nor U5585 (N_5585,N_3959,N_4045);
and U5586 (N_5586,N_4158,N_4056);
nand U5587 (N_5587,N_3188,N_3603);
and U5588 (N_5588,N_3197,N_3596);
nand U5589 (N_5589,N_4160,N_3896);
nor U5590 (N_5590,N_3114,N_4242);
or U5591 (N_5591,N_4090,N_4403);
nand U5592 (N_5592,N_3962,N_3660);
or U5593 (N_5593,N_4382,N_3189);
or U5594 (N_5594,N_3103,N_3974);
or U5595 (N_5595,N_4217,N_3623);
or U5596 (N_5596,N_3324,N_4456);
nand U5597 (N_5597,N_3395,N_3619);
or U5598 (N_5598,N_3222,N_3206);
nand U5599 (N_5599,N_3567,N_3024);
nand U5600 (N_5600,N_4283,N_3907);
and U5601 (N_5601,N_4298,N_4335);
nor U5602 (N_5602,N_3711,N_4482);
and U5603 (N_5603,N_3297,N_3475);
nand U5604 (N_5604,N_4316,N_3905);
nand U5605 (N_5605,N_3062,N_3357);
nor U5606 (N_5606,N_3579,N_3791);
and U5607 (N_5607,N_3214,N_3466);
and U5608 (N_5608,N_4240,N_4256);
or U5609 (N_5609,N_3676,N_4299);
nor U5610 (N_5610,N_3099,N_3967);
and U5611 (N_5611,N_3116,N_3301);
or U5612 (N_5612,N_4247,N_4006);
and U5613 (N_5613,N_3068,N_3041);
nor U5614 (N_5614,N_4046,N_3747);
nand U5615 (N_5615,N_3380,N_3297);
and U5616 (N_5616,N_3191,N_4011);
and U5617 (N_5617,N_3494,N_4340);
nand U5618 (N_5618,N_3298,N_3034);
and U5619 (N_5619,N_4264,N_4376);
nor U5620 (N_5620,N_4453,N_3977);
and U5621 (N_5621,N_3397,N_3617);
nor U5622 (N_5622,N_3659,N_3300);
or U5623 (N_5623,N_3688,N_3210);
nor U5624 (N_5624,N_3910,N_4216);
or U5625 (N_5625,N_4127,N_4348);
nor U5626 (N_5626,N_4222,N_3065);
nand U5627 (N_5627,N_3328,N_4173);
nor U5628 (N_5628,N_3995,N_3715);
or U5629 (N_5629,N_3500,N_4482);
nand U5630 (N_5630,N_3842,N_3181);
nand U5631 (N_5631,N_4339,N_3768);
nand U5632 (N_5632,N_3639,N_4098);
nor U5633 (N_5633,N_3110,N_4079);
nor U5634 (N_5634,N_3296,N_4266);
nand U5635 (N_5635,N_3787,N_3080);
nand U5636 (N_5636,N_3404,N_4137);
or U5637 (N_5637,N_3340,N_4432);
or U5638 (N_5638,N_4428,N_3563);
nand U5639 (N_5639,N_4124,N_3697);
nand U5640 (N_5640,N_3759,N_3177);
nor U5641 (N_5641,N_3131,N_3734);
or U5642 (N_5642,N_3268,N_3175);
nand U5643 (N_5643,N_4143,N_4236);
nor U5644 (N_5644,N_4079,N_4157);
or U5645 (N_5645,N_3922,N_3102);
nand U5646 (N_5646,N_4207,N_3891);
nor U5647 (N_5647,N_3472,N_3955);
and U5648 (N_5648,N_4136,N_3609);
nor U5649 (N_5649,N_3525,N_4006);
and U5650 (N_5650,N_3080,N_3322);
nand U5651 (N_5651,N_3112,N_3409);
and U5652 (N_5652,N_3919,N_4206);
or U5653 (N_5653,N_4093,N_3843);
nand U5654 (N_5654,N_4270,N_3246);
nor U5655 (N_5655,N_3223,N_3897);
or U5656 (N_5656,N_4151,N_4431);
nand U5657 (N_5657,N_3885,N_3834);
or U5658 (N_5658,N_3794,N_4188);
nor U5659 (N_5659,N_4457,N_3664);
nand U5660 (N_5660,N_3112,N_4369);
and U5661 (N_5661,N_3825,N_3539);
and U5662 (N_5662,N_3847,N_3385);
and U5663 (N_5663,N_4229,N_3819);
nand U5664 (N_5664,N_3411,N_3464);
and U5665 (N_5665,N_3518,N_3020);
or U5666 (N_5666,N_3609,N_4290);
nor U5667 (N_5667,N_4060,N_3843);
or U5668 (N_5668,N_3301,N_3593);
nand U5669 (N_5669,N_4230,N_3853);
and U5670 (N_5670,N_3197,N_3425);
nor U5671 (N_5671,N_3871,N_3753);
or U5672 (N_5672,N_3182,N_4344);
or U5673 (N_5673,N_3513,N_3726);
or U5674 (N_5674,N_3962,N_3646);
or U5675 (N_5675,N_3870,N_4031);
or U5676 (N_5676,N_3934,N_3095);
nand U5677 (N_5677,N_4409,N_3349);
nand U5678 (N_5678,N_4052,N_3879);
or U5679 (N_5679,N_4233,N_3530);
nand U5680 (N_5680,N_3090,N_4276);
or U5681 (N_5681,N_3958,N_3432);
or U5682 (N_5682,N_4243,N_4314);
or U5683 (N_5683,N_3354,N_3425);
nand U5684 (N_5684,N_4241,N_4396);
nor U5685 (N_5685,N_4328,N_3151);
nand U5686 (N_5686,N_3329,N_3611);
nor U5687 (N_5687,N_3987,N_3246);
or U5688 (N_5688,N_3804,N_4350);
nor U5689 (N_5689,N_3289,N_3724);
nor U5690 (N_5690,N_3491,N_3840);
and U5691 (N_5691,N_4141,N_4000);
nand U5692 (N_5692,N_4229,N_4455);
or U5693 (N_5693,N_3192,N_3317);
nand U5694 (N_5694,N_4274,N_3483);
nor U5695 (N_5695,N_3403,N_3831);
nor U5696 (N_5696,N_3079,N_3193);
nor U5697 (N_5697,N_3093,N_3348);
nand U5698 (N_5698,N_3658,N_3467);
and U5699 (N_5699,N_3539,N_3708);
or U5700 (N_5700,N_3908,N_3389);
and U5701 (N_5701,N_3609,N_3386);
nand U5702 (N_5702,N_3775,N_3186);
nor U5703 (N_5703,N_4058,N_4292);
nor U5704 (N_5704,N_3582,N_4325);
nand U5705 (N_5705,N_3006,N_3226);
and U5706 (N_5706,N_3260,N_3400);
and U5707 (N_5707,N_3525,N_4237);
or U5708 (N_5708,N_4078,N_4042);
or U5709 (N_5709,N_4134,N_4445);
or U5710 (N_5710,N_4083,N_4328);
and U5711 (N_5711,N_3612,N_4015);
and U5712 (N_5712,N_3656,N_3283);
nand U5713 (N_5713,N_3352,N_3343);
and U5714 (N_5714,N_3310,N_3356);
nand U5715 (N_5715,N_3048,N_4262);
nor U5716 (N_5716,N_3115,N_3153);
xnor U5717 (N_5717,N_4054,N_3160);
or U5718 (N_5718,N_3663,N_3928);
nand U5719 (N_5719,N_3356,N_3663);
or U5720 (N_5720,N_3095,N_3154);
nand U5721 (N_5721,N_3719,N_4416);
or U5722 (N_5722,N_4443,N_3716);
xnor U5723 (N_5723,N_4210,N_3516);
or U5724 (N_5724,N_3583,N_4497);
and U5725 (N_5725,N_3225,N_3560);
nor U5726 (N_5726,N_4103,N_4302);
and U5727 (N_5727,N_3829,N_4012);
and U5728 (N_5728,N_3271,N_3463);
and U5729 (N_5729,N_3545,N_3477);
nand U5730 (N_5730,N_3190,N_3700);
and U5731 (N_5731,N_3917,N_3593);
or U5732 (N_5732,N_3143,N_3493);
or U5733 (N_5733,N_3087,N_3867);
nand U5734 (N_5734,N_3258,N_3769);
or U5735 (N_5735,N_4273,N_3625);
nand U5736 (N_5736,N_4237,N_4075);
or U5737 (N_5737,N_4050,N_4101);
nor U5738 (N_5738,N_3231,N_4239);
nand U5739 (N_5739,N_3795,N_3467);
or U5740 (N_5740,N_3579,N_3578);
and U5741 (N_5741,N_3234,N_3426);
or U5742 (N_5742,N_3925,N_4086);
and U5743 (N_5743,N_3832,N_3615);
and U5744 (N_5744,N_4333,N_3493);
and U5745 (N_5745,N_3295,N_3566);
or U5746 (N_5746,N_3726,N_3304);
and U5747 (N_5747,N_4236,N_3213);
and U5748 (N_5748,N_3761,N_4303);
and U5749 (N_5749,N_3966,N_3442);
and U5750 (N_5750,N_4051,N_3560);
nand U5751 (N_5751,N_3386,N_3099);
or U5752 (N_5752,N_3120,N_3518);
nor U5753 (N_5753,N_4128,N_4473);
and U5754 (N_5754,N_3256,N_3563);
or U5755 (N_5755,N_3442,N_4380);
and U5756 (N_5756,N_3265,N_3492);
nand U5757 (N_5757,N_3996,N_4043);
or U5758 (N_5758,N_3357,N_4442);
and U5759 (N_5759,N_3229,N_4075);
and U5760 (N_5760,N_3480,N_3638);
nand U5761 (N_5761,N_3233,N_3682);
and U5762 (N_5762,N_3153,N_3453);
or U5763 (N_5763,N_3292,N_3599);
nand U5764 (N_5764,N_3368,N_4049);
nand U5765 (N_5765,N_3625,N_4156);
nor U5766 (N_5766,N_3563,N_3340);
and U5767 (N_5767,N_3660,N_4356);
nor U5768 (N_5768,N_3921,N_3988);
nor U5769 (N_5769,N_3749,N_4231);
nor U5770 (N_5770,N_3677,N_3370);
nand U5771 (N_5771,N_3278,N_4345);
nand U5772 (N_5772,N_3751,N_3818);
and U5773 (N_5773,N_3350,N_3163);
and U5774 (N_5774,N_3369,N_3207);
nand U5775 (N_5775,N_4310,N_3237);
nor U5776 (N_5776,N_3658,N_4479);
nand U5777 (N_5777,N_3689,N_3202);
nand U5778 (N_5778,N_3245,N_3928);
nor U5779 (N_5779,N_4211,N_3884);
or U5780 (N_5780,N_3300,N_3187);
nand U5781 (N_5781,N_3321,N_4335);
or U5782 (N_5782,N_4321,N_4175);
or U5783 (N_5783,N_3939,N_3310);
and U5784 (N_5784,N_3663,N_3278);
and U5785 (N_5785,N_4376,N_4199);
nor U5786 (N_5786,N_4360,N_4138);
nor U5787 (N_5787,N_3468,N_3694);
nor U5788 (N_5788,N_3887,N_3405);
and U5789 (N_5789,N_3614,N_4199);
nor U5790 (N_5790,N_3429,N_3370);
or U5791 (N_5791,N_3269,N_3320);
and U5792 (N_5792,N_3913,N_4309);
nor U5793 (N_5793,N_3141,N_3398);
or U5794 (N_5794,N_3068,N_3376);
and U5795 (N_5795,N_3917,N_3677);
nand U5796 (N_5796,N_4228,N_3386);
or U5797 (N_5797,N_3714,N_4079);
and U5798 (N_5798,N_4196,N_3274);
and U5799 (N_5799,N_3155,N_3115);
or U5800 (N_5800,N_4150,N_3270);
xor U5801 (N_5801,N_4169,N_3965);
nor U5802 (N_5802,N_3163,N_3734);
or U5803 (N_5803,N_4200,N_3668);
nor U5804 (N_5804,N_3057,N_3617);
and U5805 (N_5805,N_4244,N_3288);
and U5806 (N_5806,N_3581,N_3353);
nand U5807 (N_5807,N_3231,N_4344);
nand U5808 (N_5808,N_4145,N_3214);
and U5809 (N_5809,N_3709,N_4494);
nor U5810 (N_5810,N_3255,N_4226);
and U5811 (N_5811,N_4387,N_4196);
nor U5812 (N_5812,N_4422,N_4256);
nand U5813 (N_5813,N_3017,N_4367);
nor U5814 (N_5814,N_3499,N_3040);
or U5815 (N_5815,N_3143,N_3006);
nand U5816 (N_5816,N_4227,N_3357);
and U5817 (N_5817,N_3409,N_4416);
nand U5818 (N_5818,N_3435,N_3833);
nor U5819 (N_5819,N_4277,N_3338);
and U5820 (N_5820,N_3950,N_3519);
or U5821 (N_5821,N_3980,N_4046);
and U5822 (N_5822,N_3780,N_3207);
or U5823 (N_5823,N_3022,N_3612);
nor U5824 (N_5824,N_3208,N_3937);
nand U5825 (N_5825,N_3867,N_4040);
xor U5826 (N_5826,N_3002,N_4386);
and U5827 (N_5827,N_3156,N_3703);
nand U5828 (N_5828,N_3747,N_3248);
nor U5829 (N_5829,N_3814,N_3302);
nor U5830 (N_5830,N_4153,N_4173);
nand U5831 (N_5831,N_3248,N_4388);
and U5832 (N_5832,N_3470,N_3022);
or U5833 (N_5833,N_4340,N_4033);
nor U5834 (N_5834,N_3908,N_3429);
nand U5835 (N_5835,N_3634,N_3254);
nand U5836 (N_5836,N_3495,N_3020);
nor U5837 (N_5837,N_3896,N_4090);
nand U5838 (N_5838,N_3042,N_3735);
nor U5839 (N_5839,N_3993,N_3810);
nand U5840 (N_5840,N_3115,N_3469);
or U5841 (N_5841,N_4158,N_4434);
nor U5842 (N_5842,N_3155,N_4058);
or U5843 (N_5843,N_3280,N_4479);
nor U5844 (N_5844,N_3645,N_4038);
or U5845 (N_5845,N_3899,N_3445);
and U5846 (N_5846,N_3170,N_3322);
or U5847 (N_5847,N_4080,N_3605);
and U5848 (N_5848,N_3643,N_3419);
nor U5849 (N_5849,N_3721,N_4009);
xnor U5850 (N_5850,N_3341,N_4403);
and U5851 (N_5851,N_3735,N_4175);
or U5852 (N_5852,N_3101,N_4497);
nor U5853 (N_5853,N_3919,N_3635);
or U5854 (N_5854,N_3191,N_4070);
or U5855 (N_5855,N_4228,N_3118);
and U5856 (N_5856,N_3524,N_4199);
nor U5857 (N_5857,N_3458,N_4075);
nand U5858 (N_5858,N_4478,N_4287);
or U5859 (N_5859,N_3503,N_4383);
nand U5860 (N_5860,N_3567,N_3154);
and U5861 (N_5861,N_3987,N_3009);
nor U5862 (N_5862,N_4271,N_3361);
nor U5863 (N_5863,N_4308,N_4201);
and U5864 (N_5864,N_4140,N_3908);
or U5865 (N_5865,N_4336,N_3914);
nand U5866 (N_5866,N_3452,N_3081);
and U5867 (N_5867,N_3327,N_3355);
nor U5868 (N_5868,N_3590,N_3027);
nand U5869 (N_5869,N_4340,N_3487);
nand U5870 (N_5870,N_4023,N_3628);
or U5871 (N_5871,N_3170,N_4387);
or U5872 (N_5872,N_3314,N_3243);
and U5873 (N_5873,N_3805,N_4125);
or U5874 (N_5874,N_4393,N_3269);
and U5875 (N_5875,N_3392,N_3951);
and U5876 (N_5876,N_4327,N_3764);
and U5877 (N_5877,N_3027,N_3968);
or U5878 (N_5878,N_3264,N_3665);
nand U5879 (N_5879,N_3227,N_4387);
nand U5880 (N_5880,N_3414,N_4344);
nor U5881 (N_5881,N_3224,N_4445);
nor U5882 (N_5882,N_4426,N_3147);
and U5883 (N_5883,N_4463,N_3031);
nor U5884 (N_5884,N_3856,N_4054);
and U5885 (N_5885,N_3544,N_3444);
xor U5886 (N_5886,N_3761,N_4151);
and U5887 (N_5887,N_3499,N_4219);
or U5888 (N_5888,N_4023,N_3757);
or U5889 (N_5889,N_4083,N_3137);
nor U5890 (N_5890,N_3883,N_3242);
and U5891 (N_5891,N_3286,N_3387);
and U5892 (N_5892,N_3377,N_3567);
nor U5893 (N_5893,N_3404,N_4388);
and U5894 (N_5894,N_3738,N_3618);
nand U5895 (N_5895,N_4243,N_4101);
nand U5896 (N_5896,N_3497,N_4316);
nand U5897 (N_5897,N_3861,N_3737);
and U5898 (N_5898,N_3783,N_3158);
nor U5899 (N_5899,N_3155,N_3976);
or U5900 (N_5900,N_3419,N_3435);
nand U5901 (N_5901,N_3927,N_3671);
nand U5902 (N_5902,N_3587,N_4198);
nor U5903 (N_5903,N_3360,N_3579);
nor U5904 (N_5904,N_3886,N_3400);
nand U5905 (N_5905,N_3594,N_3864);
or U5906 (N_5906,N_3042,N_4480);
nor U5907 (N_5907,N_3369,N_4409);
nand U5908 (N_5908,N_3170,N_3561);
nor U5909 (N_5909,N_3433,N_3868);
nand U5910 (N_5910,N_3407,N_3544);
nand U5911 (N_5911,N_3327,N_3938);
nor U5912 (N_5912,N_3506,N_3245);
nor U5913 (N_5913,N_4293,N_4077);
and U5914 (N_5914,N_3235,N_3181);
nor U5915 (N_5915,N_3028,N_3951);
nand U5916 (N_5916,N_3327,N_4466);
nor U5917 (N_5917,N_4109,N_3031);
or U5918 (N_5918,N_3337,N_3980);
and U5919 (N_5919,N_3443,N_3971);
nor U5920 (N_5920,N_3499,N_3565);
or U5921 (N_5921,N_3067,N_3872);
and U5922 (N_5922,N_4330,N_4083);
and U5923 (N_5923,N_4202,N_3215);
or U5924 (N_5924,N_3208,N_4022);
nand U5925 (N_5925,N_3829,N_3489);
or U5926 (N_5926,N_3636,N_3119);
and U5927 (N_5927,N_3602,N_3157);
or U5928 (N_5928,N_3045,N_3506);
nor U5929 (N_5929,N_4026,N_3893);
nand U5930 (N_5930,N_3704,N_4154);
nand U5931 (N_5931,N_3728,N_3251);
and U5932 (N_5932,N_3464,N_3799);
or U5933 (N_5933,N_4300,N_3380);
nor U5934 (N_5934,N_3158,N_3280);
or U5935 (N_5935,N_4105,N_3808);
nand U5936 (N_5936,N_3853,N_4295);
nor U5937 (N_5937,N_3327,N_3546);
nand U5938 (N_5938,N_3913,N_4086);
or U5939 (N_5939,N_3447,N_3813);
nor U5940 (N_5940,N_3304,N_3188);
and U5941 (N_5941,N_3017,N_4190);
nor U5942 (N_5942,N_3050,N_3610);
or U5943 (N_5943,N_3654,N_3219);
nand U5944 (N_5944,N_3545,N_3583);
nor U5945 (N_5945,N_3624,N_3625);
nor U5946 (N_5946,N_4253,N_4171);
or U5947 (N_5947,N_3022,N_4495);
or U5948 (N_5948,N_4263,N_3468);
nand U5949 (N_5949,N_3470,N_4152);
and U5950 (N_5950,N_3839,N_3986);
nor U5951 (N_5951,N_4442,N_4312);
and U5952 (N_5952,N_3726,N_3946);
xnor U5953 (N_5953,N_3331,N_4424);
nor U5954 (N_5954,N_4288,N_4087);
and U5955 (N_5955,N_3410,N_3248);
nand U5956 (N_5956,N_4083,N_3392);
nand U5957 (N_5957,N_3047,N_3232);
or U5958 (N_5958,N_3127,N_3849);
nor U5959 (N_5959,N_4370,N_4210);
nor U5960 (N_5960,N_3652,N_4099);
or U5961 (N_5961,N_3764,N_3460);
nor U5962 (N_5962,N_3196,N_4262);
nor U5963 (N_5963,N_3466,N_4445);
or U5964 (N_5964,N_4490,N_3884);
or U5965 (N_5965,N_3959,N_3478);
and U5966 (N_5966,N_3508,N_4467);
or U5967 (N_5967,N_3407,N_3973);
nor U5968 (N_5968,N_4293,N_3521);
or U5969 (N_5969,N_3174,N_4498);
nor U5970 (N_5970,N_4118,N_3539);
and U5971 (N_5971,N_3275,N_3522);
nand U5972 (N_5972,N_3608,N_3543);
or U5973 (N_5973,N_3688,N_3807);
and U5974 (N_5974,N_4386,N_3409);
and U5975 (N_5975,N_4280,N_3125);
nor U5976 (N_5976,N_3683,N_4116);
nor U5977 (N_5977,N_3907,N_3273);
nor U5978 (N_5978,N_3741,N_3398);
nor U5979 (N_5979,N_4387,N_3926);
or U5980 (N_5980,N_3557,N_3923);
or U5981 (N_5981,N_3005,N_4314);
nor U5982 (N_5982,N_3020,N_4299);
and U5983 (N_5983,N_3419,N_3857);
nand U5984 (N_5984,N_3846,N_3239);
or U5985 (N_5985,N_4165,N_4151);
or U5986 (N_5986,N_3259,N_3409);
nand U5987 (N_5987,N_3324,N_4236);
nand U5988 (N_5988,N_4479,N_3646);
nand U5989 (N_5989,N_3196,N_4496);
nand U5990 (N_5990,N_4288,N_3514);
nand U5991 (N_5991,N_3253,N_3236);
nor U5992 (N_5992,N_3119,N_3772);
nor U5993 (N_5993,N_3214,N_4075);
and U5994 (N_5994,N_3109,N_4426);
or U5995 (N_5995,N_3020,N_3006);
and U5996 (N_5996,N_4283,N_4265);
nor U5997 (N_5997,N_3065,N_3960);
nor U5998 (N_5998,N_3471,N_4023);
nand U5999 (N_5999,N_4047,N_3344);
nor U6000 (N_6000,N_4722,N_5086);
and U6001 (N_6001,N_5370,N_4619);
and U6002 (N_6002,N_5906,N_5986);
nor U6003 (N_6003,N_5314,N_4597);
and U6004 (N_6004,N_4582,N_5666);
nand U6005 (N_6005,N_4908,N_5013);
and U6006 (N_6006,N_5134,N_5369);
and U6007 (N_6007,N_5864,N_4645);
nand U6008 (N_6008,N_5233,N_4570);
or U6009 (N_6009,N_5439,N_5502);
nand U6010 (N_6010,N_4888,N_5266);
and U6011 (N_6011,N_5908,N_4896);
or U6012 (N_6012,N_5985,N_5357);
nor U6013 (N_6013,N_5801,N_5164);
or U6014 (N_6014,N_4929,N_5080);
and U6015 (N_6015,N_5259,N_5201);
nand U6016 (N_6016,N_5893,N_5088);
nor U6017 (N_6017,N_4680,N_4617);
nand U6018 (N_6018,N_4663,N_5501);
and U6019 (N_6019,N_5564,N_4938);
or U6020 (N_6020,N_4726,N_5417);
nand U6021 (N_6021,N_4798,N_5596);
nand U6022 (N_6022,N_4504,N_5308);
nand U6023 (N_6023,N_4960,N_4614);
or U6024 (N_6024,N_5144,N_5918);
or U6025 (N_6025,N_4544,N_4761);
and U6026 (N_6026,N_5447,N_4831);
nand U6027 (N_6027,N_5278,N_5847);
nand U6028 (N_6028,N_5002,N_5455);
or U6029 (N_6029,N_4751,N_5664);
or U6030 (N_6030,N_4980,N_5805);
and U6031 (N_6031,N_5896,N_5402);
nor U6032 (N_6032,N_5487,N_5273);
or U6033 (N_6033,N_5550,N_5118);
and U6034 (N_6034,N_4833,N_4507);
or U6035 (N_6035,N_5978,N_4591);
or U6036 (N_6036,N_4972,N_5970);
and U6037 (N_6037,N_5539,N_5670);
nand U6038 (N_6038,N_5915,N_5710);
nor U6039 (N_6039,N_5283,N_4709);
nand U6040 (N_6040,N_5121,N_4851);
nand U6041 (N_6041,N_4919,N_5746);
nor U6042 (N_6042,N_4599,N_5351);
and U6043 (N_6043,N_5165,N_4956);
or U6044 (N_6044,N_5195,N_4654);
nor U6045 (N_6045,N_4550,N_4703);
and U6046 (N_6046,N_5538,N_4917);
nor U6047 (N_6047,N_5738,N_5785);
nor U6048 (N_6048,N_5394,N_4937);
xnor U6049 (N_6049,N_4581,N_5781);
nor U6050 (N_6050,N_5373,N_5414);
nor U6051 (N_6051,N_5333,N_4775);
and U6052 (N_6052,N_4991,N_4575);
nand U6053 (N_6053,N_5058,N_5618);
or U6054 (N_6054,N_4732,N_5076);
nand U6055 (N_6055,N_5459,N_5728);
and U6056 (N_6056,N_5673,N_5342);
nor U6057 (N_6057,N_5755,N_5049);
and U6058 (N_6058,N_4502,N_5747);
nor U6059 (N_6059,N_5006,N_5466);
or U6060 (N_6060,N_5529,N_5602);
nand U6061 (N_6061,N_5696,N_5859);
nor U6062 (N_6062,N_5794,N_4734);
nor U6063 (N_6063,N_5226,N_4671);
or U6064 (N_6064,N_5488,N_5142);
nand U6065 (N_6065,N_5943,N_4524);
nand U6066 (N_6066,N_4670,N_5325);
nand U6067 (N_6067,N_4611,N_5196);
or U6068 (N_6068,N_5625,N_5037);
or U6069 (N_6069,N_5597,N_5018);
and U6070 (N_6070,N_5091,N_5222);
and U6071 (N_6071,N_5423,N_5850);
nand U6072 (N_6072,N_4829,N_5576);
nor U6073 (N_6073,N_5147,N_5033);
and U6074 (N_6074,N_5727,N_5900);
or U6075 (N_6075,N_4669,N_5262);
or U6076 (N_6076,N_5062,N_5969);
nor U6077 (N_6077,N_4779,N_5378);
nand U6078 (N_6078,N_4871,N_5675);
and U6079 (N_6079,N_5102,N_5247);
and U6080 (N_6080,N_5567,N_4718);
nor U6081 (N_6081,N_5729,N_5268);
or U6082 (N_6082,N_5832,N_4810);
nor U6083 (N_6083,N_5724,N_4749);
nand U6084 (N_6084,N_5234,N_4877);
nor U6085 (N_6085,N_5363,N_5108);
or U6086 (N_6086,N_5793,N_5715);
and U6087 (N_6087,N_5881,N_4790);
and U6088 (N_6088,N_5762,N_5603);
and U6089 (N_6089,N_4783,N_5372);
or U6090 (N_6090,N_5667,N_5320);
and U6091 (N_6091,N_4762,N_5679);
nor U6092 (N_6092,N_4867,N_4687);
or U6093 (N_6093,N_4700,N_5419);
or U6094 (N_6094,N_5169,N_5937);
and U6095 (N_6095,N_5189,N_5471);
nor U6096 (N_6096,N_4895,N_5537);
and U6097 (N_6097,N_4693,N_5034);
nor U6098 (N_6098,N_5964,N_5249);
or U6099 (N_6099,N_4936,N_5418);
nand U6100 (N_6100,N_5580,N_5701);
or U6101 (N_6101,N_4568,N_4714);
and U6102 (N_6102,N_5128,N_5287);
and U6103 (N_6103,N_5154,N_4786);
or U6104 (N_6104,N_4816,N_4536);
or U6105 (N_6105,N_5178,N_5512);
nor U6106 (N_6106,N_4861,N_5732);
nand U6107 (N_6107,N_5981,N_4674);
or U6108 (N_6108,N_5174,N_4750);
nor U6109 (N_6109,N_4765,N_5940);
or U6110 (N_6110,N_4975,N_4627);
nand U6111 (N_6111,N_4901,N_5607);
nor U6112 (N_6112,N_4935,N_4648);
and U6113 (N_6113,N_5548,N_4985);
nor U6114 (N_6114,N_4918,N_5008);
nand U6115 (N_6115,N_5410,N_4606);
or U6116 (N_6116,N_4845,N_4828);
or U6117 (N_6117,N_5256,N_4827);
or U6118 (N_6118,N_5484,N_5944);
or U6119 (N_6119,N_5454,N_5767);
nand U6120 (N_6120,N_5492,N_5127);
and U6121 (N_6121,N_5740,N_4961);
nand U6122 (N_6122,N_5103,N_5766);
nand U6123 (N_6123,N_4637,N_5486);
nor U6124 (N_6124,N_4883,N_5116);
and U6125 (N_6125,N_5682,N_5123);
and U6126 (N_6126,N_5185,N_4590);
and U6127 (N_6127,N_5428,N_5163);
and U6128 (N_6128,N_5568,N_5302);
nor U6129 (N_6129,N_4554,N_5431);
or U6130 (N_6130,N_4676,N_4576);
and U6131 (N_6131,N_5110,N_4994);
nor U6132 (N_6132,N_4651,N_5097);
and U6133 (N_6133,N_5555,N_5718);
or U6134 (N_6134,N_4812,N_4572);
or U6135 (N_6135,N_5072,N_5199);
or U6136 (N_6136,N_5700,N_5294);
nor U6137 (N_6137,N_5996,N_4846);
and U6138 (N_6138,N_4634,N_4657);
nand U6139 (N_6139,N_5286,N_5031);
nand U6140 (N_6140,N_4759,N_5524);
nand U6141 (N_6141,N_4552,N_5520);
nand U6142 (N_6142,N_5497,N_4844);
xnor U6143 (N_6143,N_4534,N_4787);
and U6144 (N_6144,N_5078,N_4630);
and U6145 (N_6145,N_5813,N_5546);
and U6146 (N_6146,N_5545,N_5005);
nand U6147 (N_6147,N_5400,N_5894);
nor U6148 (N_6148,N_5077,N_5133);
nand U6149 (N_6149,N_5999,N_5338);
nor U6150 (N_6150,N_5240,N_5167);
nor U6151 (N_6151,N_5748,N_5560);
xor U6152 (N_6152,N_4672,N_5723);
and U6153 (N_6153,N_5463,N_5087);
or U6154 (N_6154,N_5557,N_5769);
and U6155 (N_6155,N_5143,N_5526);
and U6156 (N_6156,N_5582,N_5117);
nor U6157 (N_6157,N_5146,N_4748);
nand U6158 (N_6158,N_5585,N_5648);
nor U6159 (N_6159,N_5562,N_4500);
and U6160 (N_6160,N_5879,N_4633);
nand U6161 (N_6161,N_5998,N_5451);
or U6162 (N_6162,N_5365,N_5802);
nand U6163 (N_6163,N_4983,N_5371);
nor U6164 (N_6164,N_5381,N_5276);
nor U6165 (N_6165,N_5329,N_5563);
nor U6166 (N_6166,N_5971,N_5092);
and U6167 (N_6167,N_5997,N_5383);
nand U6168 (N_6168,N_5022,N_4853);
nand U6169 (N_6169,N_4584,N_4602);
or U6170 (N_6170,N_5750,N_5947);
or U6171 (N_6171,N_5194,N_5852);
and U6172 (N_6172,N_4684,N_5938);
nand U6173 (N_6173,N_5623,N_4915);
nor U6174 (N_6174,N_5267,N_5742);
nor U6175 (N_6175,N_5160,N_5324);
or U6176 (N_6176,N_5404,N_4825);
or U6177 (N_6177,N_4989,N_4686);
or U6178 (N_6178,N_5109,N_5309);
nor U6179 (N_6179,N_4661,N_5967);
nor U6180 (N_6180,N_4708,N_5743);
nor U6181 (N_6181,N_5677,N_5244);
or U6182 (N_6182,N_4652,N_4868);
and U6183 (N_6183,N_5838,N_5590);
nor U6184 (N_6184,N_4885,N_5074);
and U6185 (N_6185,N_4636,N_4540);
nor U6186 (N_6186,N_5464,N_5554);
or U6187 (N_6187,N_5136,N_4737);
and U6188 (N_6188,N_4631,N_5469);
and U6189 (N_6189,N_5584,N_4515);
nand U6190 (N_6190,N_4607,N_4688);
and U6191 (N_6191,N_4594,N_4753);
nand U6192 (N_6192,N_5248,N_4859);
nor U6193 (N_6193,N_5242,N_5470);
nor U6194 (N_6194,N_5857,N_4695);
nand U6195 (N_6195,N_5835,N_5542);
and U6196 (N_6196,N_4518,N_4981);
or U6197 (N_6197,N_4875,N_5885);
nand U6198 (N_6198,N_5792,N_4589);
nor U6199 (N_6199,N_5654,N_5812);
and U6200 (N_6200,N_5699,N_5975);
or U6201 (N_6201,N_5181,N_4503);
or U6202 (N_6202,N_5780,N_5433);
or U6203 (N_6203,N_5901,N_5983);
nor U6204 (N_6204,N_4840,N_5432);
or U6205 (N_6205,N_5948,N_5961);
nor U6206 (N_6206,N_5528,N_5284);
nand U6207 (N_6207,N_4909,N_4795);
or U6208 (N_6208,N_5200,N_5485);
nor U6209 (N_6209,N_5819,N_4778);
or U6210 (N_6210,N_5071,N_4723);
and U6211 (N_6211,N_5281,N_5902);
nand U6212 (N_6212,N_5279,N_5556);
or U6213 (N_6213,N_5737,N_4966);
or U6214 (N_6214,N_4506,N_5922);
or U6215 (N_6215,N_4880,N_5422);
nand U6216 (N_6216,N_4942,N_5023);
xnor U6217 (N_6217,N_5691,N_4848);
and U6218 (N_6218,N_4921,N_5318);
and U6219 (N_6219,N_4683,N_4804);
xor U6220 (N_6220,N_5208,N_5490);
or U6221 (N_6221,N_5692,N_5095);
nor U6222 (N_6222,N_5429,N_4797);
nand U6223 (N_6223,N_4516,N_4662);
nand U6224 (N_6224,N_5703,N_5100);
nor U6225 (N_6225,N_5788,N_5571);
nand U6226 (N_6226,N_4667,N_4870);
or U6227 (N_6227,N_4934,N_5066);
and U6228 (N_6228,N_5628,N_4526);
nand U6229 (N_6229,N_4874,N_5916);
and U6230 (N_6230,N_5148,N_5229);
xnor U6231 (N_6231,N_5300,N_5060);
xnor U6232 (N_6232,N_5816,N_4558);
nand U6233 (N_6233,N_5811,N_5990);
or U6234 (N_6234,N_5213,N_5385);
nand U6235 (N_6235,N_5337,N_5375);
or U6236 (N_6236,N_5028,N_5330);
or U6237 (N_6237,N_5828,N_4603);
and U6238 (N_6238,N_4926,N_4852);
and U6239 (N_6239,N_5021,N_5430);
or U6240 (N_6240,N_5561,N_5712);
or U6241 (N_6241,N_5782,N_5877);
nand U6242 (N_6242,N_4818,N_5265);
and U6243 (N_6243,N_5068,N_4839);
and U6244 (N_6244,N_5391,N_4557);
or U6245 (N_6245,N_5674,N_5854);
nand U6246 (N_6246,N_4819,N_5652);
nor U6247 (N_6247,N_4897,N_5310);
nor U6248 (N_6248,N_5032,N_5653);
nand U6249 (N_6249,N_5587,N_4566);
nand U6250 (N_6250,N_5959,N_5549);
and U6251 (N_6251,N_5051,N_5791);
nand U6252 (N_6252,N_4701,N_5082);
nand U6253 (N_6253,N_5220,N_4613);
nor U6254 (N_6254,N_5506,N_4528);
or U6255 (N_6255,N_5861,N_4706);
nor U6256 (N_6256,N_4916,N_5680);
nand U6257 (N_6257,N_4642,N_4881);
and U6258 (N_6258,N_5536,N_4622);
and U6259 (N_6259,N_5912,N_4857);
nor U6260 (N_6260,N_4940,N_4585);
and U6261 (N_6261,N_5586,N_5368);
or U6262 (N_6262,N_5202,N_5204);
nor U6263 (N_6263,N_5209,N_4547);
nand U6264 (N_6264,N_4941,N_5296);
nand U6265 (N_6265,N_5669,N_5598);
nor U6266 (N_6266,N_5435,N_5608);
or U6267 (N_6267,N_5192,N_5166);
or U6268 (N_6268,N_5112,N_5177);
and U6269 (N_6269,N_4521,N_4612);
xnor U6270 (N_6270,N_4620,N_5437);
and U6271 (N_6271,N_4794,N_4730);
nor U6272 (N_6272,N_5408,N_5355);
and U6273 (N_6273,N_5887,N_4678);
and U6274 (N_6274,N_4979,N_5619);
or U6275 (N_6275,N_5629,N_4978);
or U6276 (N_6276,N_4533,N_5295);
nand U6277 (N_6277,N_5041,N_5016);
nor U6278 (N_6278,N_5389,N_5387);
nand U6279 (N_6279,N_4965,N_4717);
nand U6280 (N_6280,N_4922,N_5162);
and U6281 (N_6281,N_4963,N_5588);
nor U6282 (N_6282,N_5465,N_5317);
nor U6283 (N_6283,N_4580,N_5962);
nand U6284 (N_6284,N_5907,N_5786);
nand U6285 (N_6285,N_5919,N_4792);
and U6286 (N_6286,N_5480,N_5328);
nand U6287 (N_6287,N_5264,N_5450);
nor U6288 (N_6288,N_5534,N_4999);
or U6289 (N_6289,N_5662,N_5514);
nand U6290 (N_6290,N_5228,N_5952);
or U6291 (N_6291,N_5269,N_5444);
or U6292 (N_6292,N_5065,N_5245);
and U6293 (N_6293,N_5496,N_5796);
or U6294 (N_6294,N_5476,N_5739);
nand U6295 (N_6295,N_4691,N_5255);
xnor U6296 (N_6296,N_5883,N_5860);
or U6297 (N_6297,N_5804,N_4933);
or U6298 (N_6298,N_4583,N_4555);
and U6299 (N_6299,N_5218,N_4553);
nand U6300 (N_6300,N_5821,N_4729);
nand U6301 (N_6301,N_5977,N_5275);
and U6302 (N_6302,N_5698,N_5566);
nor U6303 (N_6303,N_5634,N_5868);
nand U6304 (N_6304,N_5336,N_4905);
nand U6305 (N_6305,N_5219,N_5643);
and U6306 (N_6306,N_5960,N_5137);
nand U6307 (N_6307,N_5210,N_5695);
nor U6308 (N_6308,N_5413,N_4702);
and U6309 (N_6309,N_4973,N_5053);
or U6310 (N_6310,N_5449,N_5914);
or U6311 (N_6311,N_5702,N_5246);
nor U6312 (N_6312,N_5657,N_5009);
and U6313 (N_6313,N_4882,N_5771);
or U6314 (N_6314,N_5017,N_5676);
nor U6315 (N_6315,N_5443,N_4564);
and U6316 (N_6316,N_5768,N_5182);
nor U6317 (N_6317,N_4754,N_4982);
and U6318 (N_6318,N_4559,N_4813);
or U6319 (N_6319,N_5764,N_4586);
nor U6320 (N_6320,N_5660,N_4738);
nand U6321 (N_6321,N_5614,N_5936);
and U6322 (N_6322,N_4755,N_5842);
nand U6323 (N_6323,N_5856,N_4571);
or U6324 (N_6324,N_4811,N_5579);
or U6325 (N_6325,N_5079,N_5377);
nand U6326 (N_6326,N_5522,N_5305);
nand U6327 (N_6327,N_5637,N_5610);
or U6328 (N_6328,N_5044,N_4898);
nor U6329 (N_6329,N_4742,N_5036);
or U6330 (N_6330,N_4517,N_5889);
nand U6331 (N_6331,N_5638,N_5253);
nor U6332 (N_6332,N_4739,N_5933);
or U6333 (N_6333,N_5558,N_5931);
or U6334 (N_6334,N_5353,N_4805);
nand U6335 (N_6335,N_5553,N_5083);
and U6336 (N_6336,N_5232,N_5304);
and U6337 (N_6337,N_5689,N_5453);
or U6338 (N_6338,N_5711,N_5057);
and U6339 (N_6339,N_4705,N_5913);
nor U6340 (N_6340,N_5420,N_5921);
and U6341 (N_6341,N_5697,N_5559);
or U6342 (N_6342,N_4694,N_5179);
nor U6343 (N_6343,N_5261,N_5956);
nor U6344 (N_6344,N_5014,N_5543);
and U6345 (N_6345,N_4598,N_4578);
and U6346 (N_6346,N_5401,N_5157);
and U6347 (N_6347,N_5880,N_5774);
nor U6348 (N_6348,N_5726,N_5974);
nor U6349 (N_6349,N_5161,N_5411);
and U6350 (N_6350,N_5467,N_5979);
and U6351 (N_6351,N_5968,N_4866);
and U6352 (N_6352,N_5672,N_4525);
nor U6353 (N_6353,N_5719,N_4776);
nor U6354 (N_6354,N_5849,N_4842);
nor U6355 (N_6355,N_5462,N_4713);
and U6356 (N_6356,N_4609,N_5460);
or U6357 (N_6357,N_4542,N_5285);
nand U6358 (N_6358,N_5599,N_5046);
nand U6359 (N_6359,N_5367,N_4904);
nand U6360 (N_6360,N_5833,N_5084);
nor U6361 (N_6361,N_5704,N_5225);
nor U6362 (N_6362,N_5659,N_4532);
nand U6363 (N_6363,N_5871,N_5168);
nand U6364 (N_6364,N_5911,N_5651);
nor U6365 (N_6365,N_4747,N_5869);
nand U6366 (N_6366,N_4800,N_5289);
and U6367 (N_6367,N_5254,N_5690);
or U6368 (N_6368,N_4996,N_5331);
and U6369 (N_6369,N_4699,N_5081);
and U6370 (N_6370,N_4760,N_5070);
or U6371 (N_6371,N_5839,N_5569);
and U6372 (N_6372,N_5946,N_5107);
nand U6373 (N_6373,N_4501,N_5231);
nor U6374 (N_6374,N_5733,N_5096);
nor U6375 (N_6375,N_5360,N_4696);
or U6376 (N_6376,N_4858,N_5384);
or U6377 (N_6377,N_5616,N_5935);
or U6378 (N_6378,N_5565,N_4512);
xnor U6379 (N_6379,N_5535,N_5530);
or U6380 (N_6380,N_4587,N_4505);
and U6381 (N_6381,N_5656,N_4993);
nand U6382 (N_6382,N_5848,N_5632);
nand U6383 (N_6383,N_5882,N_5544);
and U6384 (N_6384,N_4543,N_4608);
nand U6385 (N_6385,N_5438,N_5957);
nand U6386 (N_6386,N_5499,N_5841);
or U6387 (N_6387,N_4712,N_4967);
nand U6388 (N_6388,N_5809,N_4892);
and U6389 (N_6389,N_4639,N_4638);
or U6390 (N_6390,N_4588,N_4535);
or U6391 (N_6391,N_5820,N_4604);
and U6392 (N_6392,N_5577,N_4675);
nor U6393 (N_6393,N_4820,N_5518);
nand U6394 (N_6394,N_4519,N_5024);
and U6395 (N_6395,N_5217,N_4656);
nand U6396 (N_6396,N_4660,N_5658);
and U6397 (N_6397,N_4789,N_5950);
nor U6398 (N_6398,N_4899,N_5260);
nand U6399 (N_6399,N_5390,N_5193);
and U6400 (N_6400,N_5479,N_4681);
and U6401 (N_6401,N_5007,N_5405);
nor U6402 (N_6402,N_4752,N_4658);
nor U6403 (N_6403,N_5876,N_5207);
nor U6404 (N_6404,N_4809,N_4860);
and U6405 (N_6405,N_5613,N_5926);
and U6406 (N_6406,N_5714,N_5751);
nand U6407 (N_6407,N_5098,N_4796);
nand U6408 (N_6408,N_5236,N_5311);
or U6409 (N_6409,N_5844,N_4862);
and U6410 (N_6410,N_4522,N_4665);
nor U6411 (N_6411,N_5039,N_5818);
and U6412 (N_6412,N_5288,N_4682);
and U6413 (N_6413,N_5426,N_5475);
nor U6414 (N_6414,N_5446,N_4766);
nand U6415 (N_6415,N_5920,N_5966);
or U6416 (N_6416,N_5441,N_4847);
or U6417 (N_6417,N_5735,N_4957);
nor U6418 (N_6418,N_5396,N_5606);
nor U6419 (N_6419,N_4741,N_5416);
or U6420 (N_6420,N_5872,N_5516);
or U6421 (N_6421,N_5257,N_5054);
nand U6422 (N_6422,N_4984,N_5366);
and U6423 (N_6423,N_4596,N_4850);
or U6424 (N_6424,N_4689,N_4799);
nor U6425 (N_6425,N_4673,N_4595);
nand U6426 (N_6426,N_4768,N_5504);
or U6427 (N_6427,N_5251,N_5640);
nor U6428 (N_6428,N_5612,N_5620);
nor U6429 (N_6429,N_5113,N_5851);
nand U6430 (N_6430,N_5489,N_4560);
and U6431 (N_6431,N_5753,N_5930);
nor U6432 (N_6432,N_4771,N_4565);
nand U6433 (N_6433,N_5334,N_5731);
or U6434 (N_6434,N_4891,N_5326);
nand U6435 (N_6435,N_5010,N_4628);
nand U6436 (N_6436,N_4976,N_5340);
or U6437 (N_6437,N_5775,N_4530);
nand U6438 (N_6438,N_4538,N_5831);
nand U6439 (N_6439,N_5797,N_5720);
nand U6440 (N_6440,N_4869,N_5379);
or U6441 (N_6441,N_4879,N_4913);
nor U6442 (N_6442,N_5271,N_5595);
or U6443 (N_6443,N_4677,N_4577);
nor U6444 (N_6444,N_5745,N_5570);
nand U6445 (N_6445,N_5863,N_4834);
and U6446 (N_6446,N_4629,N_5823);
and U6447 (N_6447,N_5646,N_4995);
nand U6448 (N_6448,N_5583,N_4843);
or U6449 (N_6449,N_5135,N_5763);
nand U6450 (N_6450,N_4551,N_5765);
or U6451 (N_6451,N_5105,N_5075);
or U6452 (N_6452,N_5787,N_5939);
nor U6453 (N_6453,N_4600,N_4821);
and U6454 (N_6454,N_4649,N_5140);
or U6455 (N_6455,N_5349,N_5364);
nor U6456 (N_6456,N_5647,N_5635);
nor U6457 (N_6457,N_5319,N_4930);
and U6458 (N_6458,N_5929,N_5589);
nand U6459 (N_6459,N_5758,N_5293);
and U6460 (N_6460,N_5170,N_5205);
nor U6461 (N_6461,N_4626,N_4715);
nand U6462 (N_6462,N_5829,N_4894);
nor U6463 (N_6463,N_4900,N_5048);
nand U6464 (N_6464,N_4514,N_5708);
and U6465 (N_6465,N_5376,N_5198);
nand U6466 (N_6466,N_5995,N_5622);
nand U6467 (N_6467,N_5783,N_5716);
nor U6468 (N_6468,N_5734,N_5111);
nand U6469 (N_6469,N_4650,N_5779);
or U6470 (N_6470,N_5191,N_5604);
nand U6471 (N_6471,N_4711,N_5025);
or U6472 (N_6472,N_5403,N_4911);
nor U6473 (N_6473,N_5949,N_5668);
or U6474 (N_6474,N_5895,N_5397);
and U6475 (N_6475,N_5993,N_5298);
and U6476 (N_6476,N_5188,N_4807);
nand U6477 (N_6477,N_5156,N_5759);
or U6478 (N_6478,N_5029,N_5749);
and U6479 (N_6479,N_5131,N_5573);
or U6480 (N_6480,N_4666,N_5045);
and U6481 (N_6481,N_4615,N_5958);
or U6482 (N_6482,N_4986,N_4782);
nor U6483 (N_6483,N_5875,N_5197);
or U6484 (N_6484,N_5332,N_5321);
and U6485 (N_6485,N_5810,N_4757);
or U6486 (N_6486,N_5523,N_5125);
nor U6487 (N_6487,N_4948,N_5282);
nand U6488 (N_6488,N_4743,N_4889);
nor U6489 (N_6489,N_5139,N_4835);
and U6490 (N_6490,N_4610,N_5655);
and U6491 (N_6491,N_5892,N_4931);
nor U6492 (N_6492,N_5398,N_4697);
nor U6493 (N_6493,N_5019,N_4736);
nand U6494 (N_6494,N_5477,N_4832);
nor U6495 (N_6495,N_5615,N_5665);
or U6496 (N_6496,N_5509,N_4593);
or U6497 (N_6497,N_4567,N_5910);
nand U6498 (N_6498,N_5928,N_5574);
and U6499 (N_6499,N_5180,N_4510);
or U6500 (N_6500,N_5953,N_5151);
nand U6501 (N_6501,N_4971,N_4964);
or U6502 (N_6502,N_5307,N_4928);
or U6503 (N_6503,N_5322,N_5891);
and U6504 (N_6504,N_5120,N_4968);
nand U6505 (N_6505,N_5130,N_5468);
or U6506 (N_6506,N_5633,N_5059);
nand U6507 (N_6507,N_4907,N_5124);
nor U6508 (N_6508,N_5686,N_5834);
nand U6509 (N_6509,N_5104,N_5547);
or U6510 (N_6510,N_4541,N_4910);
nand U6511 (N_6511,N_5352,N_5511);
and U6512 (N_6512,N_4692,N_5661);
nor U6513 (N_6513,N_5814,N_5777);
and U6514 (N_6514,N_5153,N_4962);
or U6515 (N_6515,N_5203,N_4815);
nand U6516 (N_6516,N_5984,N_5592);
or U6517 (N_6517,N_5346,N_5313);
or U6518 (N_6518,N_4841,N_4624);
or U6519 (N_6519,N_5693,N_5495);
nand U6520 (N_6520,N_4641,N_5474);
or U6521 (N_6521,N_5027,N_5155);
nor U6522 (N_6522,N_5043,N_5644);
xnor U6523 (N_6523,N_5923,N_5684);
nand U6524 (N_6524,N_4772,N_4777);
nor U6525 (N_6525,N_5064,N_4950);
nand U6526 (N_6526,N_5532,N_5458);
nor U6527 (N_6527,N_5865,N_5374);
and U6528 (N_6528,N_4826,N_5094);
and U6529 (N_6529,N_5874,N_5899);
nand U6530 (N_6530,N_4758,N_5617);
nand U6531 (N_6531,N_4655,N_5752);
nand U6532 (N_6532,N_4764,N_5965);
nor U6533 (N_6533,N_5090,N_4621);
nor U6534 (N_6534,N_5119,N_4823);
or U6535 (N_6535,N_5846,N_4646);
and U6536 (N_6536,N_4801,N_5335);
or U6537 (N_6537,N_5808,N_5671);
nand U6538 (N_6538,N_5843,N_4569);
nor U6539 (N_6539,N_5461,N_4520);
and U6540 (N_6540,N_5837,N_5101);
or U6541 (N_6541,N_5063,N_5757);
nand U6542 (N_6542,N_4546,N_5145);
nor U6543 (N_6543,N_4720,N_4814);
nor U6544 (N_6544,N_5483,N_5223);
and U6545 (N_6545,N_4763,N_5826);
xor U6546 (N_6546,N_5224,N_5639);
nor U6547 (N_6547,N_4527,N_5085);
nor U6548 (N_6548,N_5061,N_4781);
nand U6549 (N_6549,N_4733,N_5515);
or U6550 (N_6550,N_5925,N_4927);
nor U6551 (N_6551,N_4855,N_5099);
nor U6552 (N_6552,N_5149,N_4513);
or U6553 (N_6553,N_5186,N_5982);
nor U6554 (N_6554,N_5129,N_5042);
or U6555 (N_6555,N_5442,N_5510);
and U6556 (N_6556,N_5815,N_4644);
and U6557 (N_6557,N_4865,N_5798);
nor U6558 (N_6558,N_5493,N_4988);
and U6559 (N_6559,N_4562,N_4920);
or U6560 (N_6560,N_4704,N_5056);
and U6561 (N_6561,N_4923,N_5845);
or U6562 (N_6562,N_5211,N_5406);
and U6563 (N_6563,N_5991,N_5776);
nor U6564 (N_6564,N_5945,N_4756);
or U6565 (N_6565,N_5527,N_4539);
xor U6566 (N_6566,N_5344,N_4643);
nand U6567 (N_6567,N_5361,N_5159);
nand U6568 (N_6568,N_4890,N_5992);
nand U6569 (N_6569,N_4668,N_5052);
nand U6570 (N_6570,N_5754,N_5171);
nor U6571 (N_6571,N_5237,N_4601);
nor U6572 (N_6572,N_4969,N_5932);
nor U6573 (N_6573,N_5382,N_5756);
nand U6574 (N_6574,N_4944,N_5239);
and U6575 (N_6575,N_5760,N_4902);
or U6576 (N_6576,N_5290,N_4806);
nand U6577 (N_6577,N_5362,N_5380);
nor U6578 (N_6578,N_5822,N_4716);
nand U6579 (N_6579,N_5505,N_4873);
and U6580 (N_6580,N_4808,N_4893);
and U6581 (N_6581,N_4887,N_4924);
and U6582 (N_6582,N_5212,N_4523);
or U6583 (N_6583,N_5415,N_4977);
nand U6584 (N_6584,N_4925,N_5503);
or U6585 (N_6585,N_4635,N_5761);
nor U6586 (N_6586,N_5866,N_5884);
or U6587 (N_6587,N_5855,N_4574);
or U6588 (N_6588,N_5345,N_5132);
nand U6589 (N_6589,N_5277,N_5730);
nand U6590 (N_6590,N_5508,N_5327);
nor U6591 (N_6591,N_5138,N_5853);
nor U6592 (N_6592,N_4953,N_5721);
and U6593 (N_6593,N_5354,N_5122);
or U6594 (N_6594,N_5478,N_5386);
nor U6595 (N_6595,N_5491,N_5898);
nand U6596 (N_6596,N_5440,N_5641);
or U6597 (N_6597,N_5800,N_5533);
and U6598 (N_6598,N_5250,N_5452);
and U6599 (N_6599,N_4824,N_5713);
nand U6600 (N_6600,N_4537,N_5270);
or U6601 (N_6601,N_5141,N_4549);
or U6602 (N_6602,N_5954,N_5190);
or U6603 (N_6603,N_5773,N_5227);
nand U6604 (N_6604,N_5187,N_5784);
or U6605 (N_6605,N_5878,N_4592);
and U6606 (N_6606,N_5621,N_5817);
and U6607 (N_6607,N_5531,N_5717);
nand U6608 (N_6608,N_5778,N_5770);
nor U6609 (N_6609,N_4719,N_5238);
and U6610 (N_6610,N_4659,N_4997);
or U6611 (N_6611,N_5688,N_4698);
or U6612 (N_6612,N_4949,N_5407);
nand U6613 (N_6613,N_5020,N_5393);
nand U6614 (N_6614,N_5301,N_5069);
and U6615 (N_6615,N_5280,N_5867);
nor U6616 (N_6616,N_5594,N_4746);
or U6617 (N_6617,N_5593,N_5507);
nor U6618 (N_6618,N_5649,N_5315);
and U6619 (N_6619,N_4854,N_5552);
nand U6620 (N_6620,N_4951,N_5050);
nand U6621 (N_6621,N_5303,N_4864);
or U6622 (N_6622,N_5836,N_5630);
and U6623 (N_6623,N_4573,N_5243);
nand U6624 (N_6624,N_5093,N_5631);
nor U6625 (N_6625,N_4623,N_5611);
nor U6626 (N_6626,N_5214,N_4511);
or U6627 (N_6627,N_4947,N_5886);
and U6628 (N_6628,N_4548,N_4745);
nor U6629 (N_6629,N_5252,N_4785);
nor U6630 (N_6630,N_5481,N_5241);
nor U6631 (N_6631,N_4561,N_4863);
or U6632 (N_6632,N_4653,N_5924);
nor U6633 (N_6633,N_4632,N_5980);
nand U6634 (N_6634,N_4773,N_5047);
or U6635 (N_6635,N_4943,N_5230);
or U6636 (N_6636,N_4531,N_4724);
or U6637 (N_6637,N_5955,N_5706);
nand U6638 (N_6638,N_4914,N_5681);
nor U6639 (N_6639,N_5339,N_4618);
nor U6640 (N_6640,N_5272,N_4990);
and U6641 (N_6641,N_5541,N_4770);
nand U6642 (N_6642,N_4932,N_5627);
nand U6643 (N_6643,N_5221,N_5457);
or U6644 (N_6644,N_5517,N_5888);
nand U6645 (N_6645,N_5003,N_5722);
or U6646 (N_6646,N_5636,N_5862);
or U6647 (N_6647,N_4791,N_5012);
and U6648 (N_6648,N_4987,N_4728);
or U6649 (N_6649,N_5890,N_5601);
nand U6650 (N_6650,N_5011,N_5114);
or U6651 (N_6651,N_4579,N_5513);
and U6652 (N_6652,N_5291,N_5772);
or U6653 (N_6653,N_5184,N_5274);
or U6654 (N_6654,N_4830,N_4959);
nor U6655 (N_6655,N_5525,N_4856);
and U6656 (N_6656,N_5448,N_4836);
nor U6657 (N_6657,N_4793,N_5073);
nand U6658 (N_6658,N_5359,N_5521);
or U6659 (N_6659,N_4884,N_5540);
or U6660 (N_6660,N_5663,N_5806);
nor U6661 (N_6661,N_5434,N_5347);
or U6662 (N_6662,N_4946,N_5015);
nor U6663 (N_6663,N_5741,N_4625);
nand U6664 (N_6664,N_5089,N_5989);
nand U6665 (N_6665,N_4774,N_5707);
and U6666 (N_6666,N_5412,N_5001);
or U6667 (N_6667,N_5840,N_5705);
nor U6668 (N_6668,N_5678,N_5709);
and U6669 (N_6669,N_4545,N_5498);
nand U6670 (N_6670,N_5299,N_5445);
nor U6671 (N_6671,N_4838,N_5994);
and U6672 (N_6672,N_5258,N_4556);
and U6673 (N_6673,N_5425,N_5456);
nand U6674 (N_6674,N_5951,N_4788);
or U6675 (N_6675,N_5903,N_5055);
or U6676 (N_6676,N_5427,N_5725);
and U6677 (N_6677,N_4945,N_4616);
and U6678 (N_6678,N_5235,N_5343);
nand U6679 (N_6679,N_4974,N_5038);
nand U6680 (N_6680,N_4727,N_4735);
nand U6681 (N_6681,N_4690,N_5650);
nor U6682 (N_6682,N_5988,N_4731);
and U6683 (N_6683,N_5482,N_5106);
xnor U6684 (N_6684,N_5026,N_5472);
nand U6685 (N_6685,N_4970,N_4685);
nor U6686 (N_6686,N_5827,N_5215);
and U6687 (N_6687,N_4509,N_4647);
and U6688 (N_6688,N_4906,N_5591);
nor U6689 (N_6689,N_4780,N_4784);
or U6690 (N_6690,N_5519,N_4767);
nand U6691 (N_6691,N_4955,N_4710);
or U6692 (N_6692,N_5941,N_5421);
nand U6693 (N_6693,N_5348,N_4769);
and U6694 (N_6694,N_5609,N_5292);
nand U6695 (N_6695,N_5685,N_5206);
nor U6696 (N_6696,N_4707,N_5927);
and U6697 (N_6697,N_5897,N_5917);
or U6698 (N_6698,N_4744,N_5870);
nand U6699 (N_6699,N_5581,N_5600);
nor U6700 (N_6700,N_5312,N_5972);
or U6701 (N_6701,N_5399,N_4954);
or U6702 (N_6702,N_5909,N_5316);
nand U6703 (N_6703,N_5551,N_5035);
nand U6704 (N_6704,N_5388,N_5858);
nand U6705 (N_6705,N_4803,N_5626);
or U6706 (N_6706,N_5904,N_5494);
or U6707 (N_6707,N_5799,N_4740);
xnor U6708 (N_6708,N_5830,N_5356);
or U6709 (N_6709,N_5645,N_5500);
nor U6710 (N_6710,N_5172,N_4837);
or U6711 (N_6711,N_5152,N_5173);
nor U6712 (N_6712,N_5683,N_5409);
nand U6713 (N_6713,N_4849,N_4958);
nand U6714 (N_6714,N_5790,N_4939);
and U6715 (N_6715,N_5115,N_5736);
and U6716 (N_6716,N_4817,N_5578);
and U6717 (N_6717,N_5803,N_4664);
or U6718 (N_6718,N_5642,N_5150);
or U6719 (N_6719,N_5987,N_5973);
and U6720 (N_6720,N_5873,N_4903);
nand U6721 (N_6721,N_5030,N_5216);
or U6722 (N_6722,N_5000,N_5350);
nand U6723 (N_6723,N_5263,N_5040);
and U6724 (N_6724,N_5687,N_4912);
nand U6725 (N_6725,N_5624,N_4872);
nand U6726 (N_6726,N_4878,N_5934);
nand U6727 (N_6727,N_4679,N_5395);
or U6728 (N_6728,N_5004,N_5789);
and U6729 (N_6729,N_5341,N_5323);
or U6730 (N_6730,N_5424,N_4998);
or U6731 (N_6731,N_5392,N_5825);
and U6732 (N_6732,N_5976,N_5183);
or U6733 (N_6733,N_5572,N_5158);
and U6734 (N_6734,N_4952,N_5807);
or U6735 (N_6735,N_5175,N_4563);
nand U6736 (N_6736,N_5306,N_4605);
nand U6737 (N_6737,N_5575,N_5067);
or U6738 (N_6738,N_5963,N_4640);
nor U6739 (N_6739,N_5605,N_4508);
and U6740 (N_6740,N_5942,N_5358);
or U6741 (N_6741,N_5436,N_4822);
and U6742 (N_6742,N_5297,N_4876);
and U6743 (N_6743,N_4802,N_4725);
and U6744 (N_6744,N_5126,N_5824);
nand U6745 (N_6745,N_5905,N_5795);
nand U6746 (N_6746,N_5744,N_5473);
nor U6747 (N_6747,N_4886,N_4721);
nor U6748 (N_6748,N_4992,N_5694);
nor U6749 (N_6749,N_5176,N_4529);
nor U6750 (N_6750,N_4959,N_4704);
nand U6751 (N_6751,N_5272,N_5526);
or U6752 (N_6752,N_5178,N_5405);
nor U6753 (N_6753,N_5455,N_5921);
nor U6754 (N_6754,N_5160,N_4643);
nand U6755 (N_6755,N_4771,N_4717);
or U6756 (N_6756,N_5784,N_5527);
xor U6757 (N_6757,N_5160,N_5270);
nor U6758 (N_6758,N_5097,N_4863);
and U6759 (N_6759,N_5716,N_5534);
or U6760 (N_6760,N_4745,N_5382);
or U6761 (N_6761,N_5894,N_5082);
or U6762 (N_6762,N_5841,N_5581);
nor U6763 (N_6763,N_5879,N_5280);
nand U6764 (N_6764,N_4828,N_5294);
nor U6765 (N_6765,N_5600,N_4860);
and U6766 (N_6766,N_5581,N_5874);
nand U6767 (N_6767,N_4725,N_5052);
and U6768 (N_6768,N_5842,N_5222);
nor U6769 (N_6769,N_4635,N_4984);
nor U6770 (N_6770,N_5237,N_4762);
nand U6771 (N_6771,N_4516,N_4933);
and U6772 (N_6772,N_4841,N_5926);
or U6773 (N_6773,N_5553,N_5800);
nor U6774 (N_6774,N_5252,N_5758);
and U6775 (N_6775,N_5680,N_5770);
and U6776 (N_6776,N_4505,N_5845);
nor U6777 (N_6777,N_5383,N_5169);
or U6778 (N_6778,N_5439,N_4888);
nand U6779 (N_6779,N_4941,N_5933);
and U6780 (N_6780,N_5396,N_5595);
nor U6781 (N_6781,N_5133,N_5358);
and U6782 (N_6782,N_4501,N_5051);
or U6783 (N_6783,N_5056,N_5135);
and U6784 (N_6784,N_5606,N_4920);
and U6785 (N_6785,N_4841,N_5947);
nand U6786 (N_6786,N_4981,N_5517);
nand U6787 (N_6787,N_5512,N_4810);
or U6788 (N_6788,N_5152,N_4656);
or U6789 (N_6789,N_5783,N_4721);
or U6790 (N_6790,N_5864,N_5362);
nand U6791 (N_6791,N_4697,N_4672);
nor U6792 (N_6792,N_4755,N_4538);
or U6793 (N_6793,N_4647,N_5859);
or U6794 (N_6794,N_5578,N_5194);
nand U6795 (N_6795,N_4556,N_5235);
and U6796 (N_6796,N_4823,N_5272);
or U6797 (N_6797,N_4721,N_5613);
or U6798 (N_6798,N_4815,N_5066);
and U6799 (N_6799,N_5344,N_5948);
or U6800 (N_6800,N_4533,N_5065);
nand U6801 (N_6801,N_5665,N_5655);
nor U6802 (N_6802,N_5372,N_4890);
or U6803 (N_6803,N_5685,N_5325);
nand U6804 (N_6804,N_4622,N_5569);
nor U6805 (N_6805,N_5608,N_4876);
nor U6806 (N_6806,N_5481,N_5770);
nor U6807 (N_6807,N_4907,N_5642);
nor U6808 (N_6808,N_4967,N_5447);
or U6809 (N_6809,N_5823,N_5507);
and U6810 (N_6810,N_5009,N_5533);
nand U6811 (N_6811,N_4944,N_5916);
and U6812 (N_6812,N_4812,N_5168);
and U6813 (N_6813,N_4661,N_4560);
or U6814 (N_6814,N_4846,N_5396);
and U6815 (N_6815,N_4722,N_5621);
nor U6816 (N_6816,N_5346,N_5715);
and U6817 (N_6817,N_5768,N_5455);
and U6818 (N_6818,N_4568,N_5700);
nor U6819 (N_6819,N_4980,N_5111);
or U6820 (N_6820,N_5786,N_4582);
or U6821 (N_6821,N_5357,N_5432);
or U6822 (N_6822,N_5541,N_5985);
nand U6823 (N_6823,N_5483,N_5810);
nor U6824 (N_6824,N_5003,N_4605);
or U6825 (N_6825,N_5530,N_5008);
nor U6826 (N_6826,N_4835,N_5100);
nor U6827 (N_6827,N_5831,N_5916);
and U6828 (N_6828,N_4747,N_5430);
or U6829 (N_6829,N_5031,N_5225);
or U6830 (N_6830,N_5679,N_5560);
and U6831 (N_6831,N_4572,N_5448);
and U6832 (N_6832,N_5971,N_4525);
nor U6833 (N_6833,N_4955,N_5107);
nand U6834 (N_6834,N_5345,N_4698);
nand U6835 (N_6835,N_4962,N_4820);
xnor U6836 (N_6836,N_5764,N_5485);
and U6837 (N_6837,N_5029,N_4643);
nor U6838 (N_6838,N_5246,N_4908);
and U6839 (N_6839,N_4675,N_5204);
nand U6840 (N_6840,N_5472,N_5576);
and U6841 (N_6841,N_4584,N_4589);
or U6842 (N_6842,N_5988,N_4763);
or U6843 (N_6843,N_4965,N_4616);
nor U6844 (N_6844,N_5996,N_5605);
and U6845 (N_6845,N_5126,N_5637);
nand U6846 (N_6846,N_5100,N_4554);
and U6847 (N_6847,N_4881,N_5583);
nor U6848 (N_6848,N_5385,N_5493);
or U6849 (N_6849,N_4984,N_5359);
nor U6850 (N_6850,N_4841,N_5841);
xor U6851 (N_6851,N_4521,N_5623);
nor U6852 (N_6852,N_5320,N_5089);
nor U6853 (N_6853,N_4964,N_5919);
or U6854 (N_6854,N_5310,N_5994);
nand U6855 (N_6855,N_5329,N_4683);
or U6856 (N_6856,N_5885,N_4656);
and U6857 (N_6857,N_5489,N_5969);
and U6858 (N_6858,N_5943,N_4580);
nand U6859 (N_6859,N_5521,N_4931);
or U6860 (N_6860,N_5960,N_4819);
nor U6861 (N_6861,N_4528,N_5075);
nand U6862 (N_6862,N_4938,N_5332);
and U6863 (N_6863,N_4587,N_5832);
or U6864 (N_6864,N_4695,N_5608);
nor U6865 (N_6865,N_5592,N_5844);
nor U6866 (N_6866,N_5119,N_5218);
nand U6867 (N_6867,N_5795,N_5231);
nor U6868 (N_6868,N_5475,N_5402);
and U6869 (N_6869,N_4646,N_4630);
and U6870 (N_6870,N_5244,N_5086);
and U6871 (N_6871,N_4537,N_5512);
nor U6872 (N_6872,N_5660,N_5542);
nor U6873 (N_6873,N_5649,N_4533);
or U6874 (N_6874,N_4882,N_5876);
nor U6875 (N_6875,N_5169,N_4733);
or U6876 (N_6876,N_5166,N_5353);
or U6877 (N_6877,N_4873,N_4989);
and U6878 (N_6878,N_4553,N_5331);
or U6879 (N_6879,N_4683,N_5416);
and U6880 (N_6880,N_5920,N_5571);
and U6881 (N_6881,N_5988,N_5119);
or U6882 (N_6882,N_4684,N_4748);
nor U6883 (N_6883,N_5585,N_4676);
or U6884 (N_6884,N_5573,N_5375);
nor U6885 (N_6885,N_5504,N_5000);
nor U6886 (N_6886,N_5354,N_5734);
and U6887 (N_6887,N_4541,N_5138);
xor U6888 (N_6888,N_4747,N_4592);
or U6889 (N_6889,N_4862,N_5941);
nand U6890 (N_6890,N_5586,N_5057);
xor U6891 (N_6891,N_5881,N_5114);
nand U6892 (N_6892,N_5597,N_4843);
or U6893 (N_6893,N_4511,N_5900);
nand U6894 (N_6894,N_4861,N_4914);
and U6895 (N_6895,N_5293,N_5656);
nand U6896 (N_6896,N_5108,N_5322);
nand U6897 (N_6897,N_5461,N_5483);
xnor U6898 (N_6898,N_4833,N_5623);
or U6899 (N_6899,N_4962,N_5064);
or U6900 (N_6900,N_4605,N_5581);
nand U6901 (N_6901,N_5972,N_5083);
nand U6902 (N_6902,N_4577,N_4823);
nand U6903 (N_6903,N_5967,N_4703);
nor U6904 (N_6904,N_5814,N_5301);
nor U6905 (N_6905,N_5288,N_4862);
nand U6906 (N_6906,N_5289,N_5457);
nor U6907 (N_6907,N_5068,N_4930);
nor U6908 (N_6908,N_5528,N_5793);
and U6909 (N_6909,N_4892,N_5773);
nand U6910 (N_6910,N_5082,N_4957);
nand U6911 (N_6911,N_4743,N_5764);
or U6912 (N_6912,N_5726,N_5558);
and U6913 (N_6913,N_4721,N_4850);
nor U6914 (N_6914,N_5716,N_4719);
and U6915 (N_6915,N_4645,N_5992);
or U6916 (N_6916,N_5511,N_5987);
and U6917 (N_6917,N_5097,N_4707);
nand U6918 (N_6918,N_5405,N_5803);
nand U6919 (N_6919,N_5684,N_5937);
or U6920 (N_6920,N_4717,N_5134);
nand U6921 (N_6921,N_5140,N_5953);
or U6922 (N_6922,N_5319,N_5604);
nor U6923 (N_6923,N_5296,N_5558);
and U6924 (N_6924,N_5842,N_5211);
nor U6925 (N_6925,N_5714,N_4737);
nand U6926 (N_6926,N_5493,N_5219);
nor U6927 (N_6927,N_4902,N_4655);
nand U6928 (N_6928,N_5577,N_5077);
nand U6929 (N_6929,N_5094,N_5868);
nand U6930 (N_6930,N_5616,N_4804);
nand U6931 (N_6931,N_5817,N_5646);
and U6932 (N_6932,N_5876,N_5873);
or U6933 (N_6933,N_5267,N_5520);
xor U6934 (N_6934,N_4535,N_5936);
nor U6935 (N_6935,N_5913,N_5281);
nand U6936 (N_6936,N_4949,N_4983);
nor U6937 (N_6937,N_5535,N_5287);
or U6938 (N_6938,N_5036,N_4924);
and U6939 (N_6939,N_5819,N_4947);
or U6940 (N_6940,N_4868,N_5678);
and U6941 (N_6941,N_5446,N_4976);
or U6942 (N_6942,N_5543,N_5781);
nand U6943 (N_6943,N_5312,N_5725);
nand U6944 (N_6944,N_5158,N_4563);
and U6945 (N_6945,N_5942,N_5795);
or U6946 (N_6946,N_5396,N_5185);
and U6947 (N_6947,N_5758,N_4543);
or U6948 (N_6948,N_5135,N_4952);
nand U6949 (N_6949,N_4815,N_4641);
nor U6950 (N_6950,N_5318,N_5778);
nand U6951 (N_6951,N_5173,N_5299);
and U6952 (N_6952,N_5252,N_5745);
and U6953 (N_6953,N_5971,N_4524);
or U6954 (N_6954,N_5211,N_4847);
and U6955 (N_6955,N_5790,N_5041);
and U6956 (N_6956,N_5210,N_5775);
or U6957 (N_6957,N_5878,N_4508);
or U6958 (N_6958,N_5882,N_4670);
nand U6959 (N_6959,N_5948,N_5306);
nand U6960 (N_6960,N_5400,N_5128);
nand U6961 (N_6961,N_4699,N_4503);
nor U6962 (N_6962,N_5055,N_5375);
or U6963 (N_6963,N_5889,N_4845);
nand U6964 (N_6964,N_5448,N_4619);
or U6965 (N_6965,N_4672,N_5280);
nand U6966 (N_6966,N_5888,N_4850);
and U6967 (N_6967,N_5305,N_4945);
and U6968 (N_6968,N_5405,N_5847);
nor U6969 (N_6969,N_4622,N_5711);
nand U6970 (N_6970,N_4698,N_4930);
nor U6971 (N_6971,N_4595,N_4626);
or U6972 (N_6972,N_4662,N_4601);
or U6973 (N_6973,N_5502,N_4660);
and U6974 (N_6974,N_5073,N_5145);
nor U6975 (N_6975,N_5837,N_4978);
xnor U6976 (N_6976,N_5323,N_5847);
and U6977 (N_6977,N_5046,N_5689);
or U6978 (N_6978,N_5518,N_4650);
nor U6979 (N_6979,N_4538,N_5802);
or U6980 (N_6980,N_4582,N_5370);
or U6981 (N_6981,N_4918,N_5559);
nand U6982 (N_6982,N_5519,N_5540);
nand U6983 (N_6983,N_4693,N_5158);
or U6984 (N_6984,N_5345,N_5106);
or U6985 (N_6985,N_5345,N_4713);
or U6986 (N_6986,N_4513,N_4579);
and U6987 (N_6987,N_5831,N_4824);
nand U6988 (N_6988,N_4710,N_5551);
nand U6989 (N_6989,N_5718,N_5970);
nand U6990 (N_6990,N_5233,N_5316);
nand U6991 (N_6991,N_5846,N_4895);
nor U6992 (N_6992,N_5323,N_5023);
nand U6993 (N_6993,N_4932,N_5156);
nor U6994 (N_6994,N_4853,N_4767);
and U6995 (N_6995,N_5148,N_5161);
or U6996 (N_6996,N_4580,N_4696);
nor U6997 (N_6997,N_5706,N_4714);
nor U6998 (N_6998,N_5950,N_5697);
and U6999 (N_6999,N_5990,N_4850);
and U7000 (N_7000,N_5320,N_5257);
nor U7001 (N_7001,N_5795,N_4783);
nand U7002 (N_7002,N_5349,N_4798);
xnor U7003 (N_7003,N_5219,N_4728);
nand U7004 (N_7004,N_4508,N_4705);
or U7005 (N_7005,N_5864,N_4997);
or U7006 (N_7006,N_5815,N_5788);
nor U7007 (N_7007,N_4571,N_5642);
and U7008 (N_7008,N_5850,N_5483);
nor U7009 (N_7009,N_5563,N_5207);
nor U7010 (N_7010,N_4577,N_5249);
and U7011 (N_7011,N_5141,N_5917);
and U7012 (N_7012,N_4648,N_4713);
nor U7013 (N_7013,N_5714,N_5631);
nand U7014 (N_7014,N_4917,N_5794);
nor U7015 (N_7015,N_4611,N_4827);
or U7016 (N_7016,N_5574,N_5029);
and U7017 (N_7017,N_5154,N_5492);
and U7018 (N_7018,N_5717,N_5974);
nor U7019 (N_7019,N_4925,N_5861);
nor U7020 (N_7020,N_5020,N_5450);
nor U7021 (N_7021,N_5727,N_5949);
or U7022 (N_7022,N_5104,N_5754);
or U7023 (N_7023,N_5543,N_4639);
nor U7024 (N_7024,N_5120,N_4927);
and U7025 (N_7025,N_5079,N_4737);
or U7026 (N_7026,N_4925,N_5566);
nand U7027 (N_7027,N_4759,N_4684);
nand U7028 (N_7028,N_4940,N_5015);
nor U7029 (N_7029,N_4989,N_5832);
nand U7030 (N_7030,N_5084,N_5390);
nor U7031 (N_7031,N_5978,N_5606);
nor U7032 (N_7032,N_4651,N_4764);
and U7033 (N_7033,N_5142,N_5434);
and U7034 (N_7034,N_5576,N_5159);
and U7035 (N_7035,N_5254,N_5553);
nor U7036 (N_7036,N_5778,N_5806);
and U7037 (N_7037,N_5886,N_5385);
xnor U7038 (N_7038,N_4604,N_5430);
nand U7039 (N_7039,N_5592,N_5118);
nor U7040 (N_7040,N_4952,N_5609);
and U7041 (N_7041,N_4820,N_5542);
nand U7042 (N_7042,N_5936,N_5603);
or U7043 (N_7043,N_5979,N_4549);
and U7044 (N_7044,N_4543,N_5473);
nor U7045 (N_7045,N_5929,N_5072);
and U7046 (N_7046,N_5000,N_5614);
or U7047 (N_7047,N_4813,N_5422);
or U7048 (N_7048,N_5883,N_5544);
and U7049 (N_7049,N_5703,N_5882);
and U7050 (N_7050,N_5858,N_5800);
or U7051 (N_7051,N_5980,N_5837);
or U7052 (N_7052,N_5950,N_4902);
nand U7053 (N_7053,N_5080,N_4546);
nor U7054 (N_7054,N_5255,N_4935);
and U7055 (N_7055,N_5497,N_5072);
nand U7056 (N_7056,N_5607,N_5459);
nand U7057 (N_7057,N_5785,N_5349);
nand U7058 (N_7058,N_5477,N_5390);
and U7059 (N_7059,N_4665,N_5221);
nor U7060 (N_7060,N_5072,N_4683);
and U7061 (N_7061,N_5860,N_4711);
and U7062 (N_7062,N_5262,N_5328);
or U7063 (N_7063,N_5136,N_5347);
and U7064 (N_7064,N_4928,N_5583);
and U7065 (N_7065,N_4620,N_5420);
or U7066 (N_7066,N_4734,N_4657);
nand U7067 (N_7067,N_5352,N_4662);
and U7068 (N_7068,N_5049,N_4577);
or U7069 (N_7069,N_5230,N_5459);
nor U7070 (N_7070,N_5865,N_5006);
or U7071 (N_7071,N_5869,N_5383);
and U7072 (N_7072,N_5082,N_4984);
nor U7073 (N_7073,N_5126,N_4819);
or U7074 (N_7074,N_4972,N_5098);
nand U7075 (N_7075,N_5182,N_4700);
and U7076 (N_7076,N_4776,N_5569);
nor U7077 (N_7077,N_5947,N_5475);
nand U7078 (N_7078,N_5659,N_5571);
and U7079 (N_7079,N_5339,N_5804);
and U7080 (N_7080,N_5709,N_4997);
xor U7081 (N_7081,N_5085,N_5352);
xor U7082 (N_7082,N_4817,N_4607);
or U7083 (N_7083,N_5323,N_5771);
or U7084 (N_7084,N_5075,N_4559);
nand U7085 (N_7085,N_5477,N_5916);
nand U7086 (N_7086,N_4934,N_5609);
and U7087 (N_7087,N_5855,N_4955);
nand U7088 (N_7088,N_4805,N_5318);
nand U7089 (N_7089,N_5956,N_4753);
nor U7090 (N_7090,N_5911,N_4572);
and U7091 (N_7091,N_5972,N_5107);
and U7092 (N_7092,N_4655,N_5205);
nor U7093 (N_7093,N_4644,N_4897);
nor U7094 (N_7094,N_5510,N_5933);
nand U7095 (N_7095,N_5329,N_5227);
and U7096 (N_7096,N_4677,N_4687);
and U7097 (N_7097,N_5276,N_5479);
nor U7098 (N_7098,N_4737,N_5514);
and U7099 (N_7099,N_5656,N_4863);
nand U7100 (N_7100,N_5534,N_5082);
nor U7101 (N_7101,N_5659,N_5292);
nor U7102 (N_7102,N_5321,N_5933);
and U7103 (N_7103,N_5328,N_4703);
and U7104 (N_7104,N_5889,N_4757);
and U7105 (N_7105,N_4636,N_5856);
nor U7106 (N_7106,N_5660,N_5476);
nor U7107 (N_7107,N_5522,N_4986);
or U7108 (N_7108,N_4509,N_5803);
nor U7109 (N_7109,N_5281,N_4658);
or U7110 (N_7110,N_5791,N_5638);
nor U7111 (N_7111,N_5168,N_5725);
or U7112 (N_7112,N_5813,N_5608);
nor U7113 (N_7113,N_4852,N_5953);
nor U7114 (N_7114,N_5012,N_5753);
or U7115 (N_7115,N_5197,N_5199);
nor U7116 (N_7116,N_5429,N_5338);
or U7117 (N_7117,N_4601,N_5542);
nand U7118 (N_7118,N_4680,N_4912);
nand U7119 (N_7119,N_4527,N_4898);
and U7120 (N_7120,N_5187,N_4574);
or U7121 (N_7121,N_5939,N_5875);
or U7122 (N_7122,N_5785,N_4919);
nor U7123 (N_7123,N_5697,N_4604);
or U7124 (N_7124,N_5609,N_4691);
and U7125 (N_7125,N_5939,N_5317);
nand U7126 (N_7126,N_5255,N_4712);
and U7127 (N_7127,N_5959,N_5706);
and U7128 (N_7128,N_5827,N_4941);
and U7129 (N_7129,N_5436,N_4889);
and U7130 (N_7130,N_4629,N_4707);
nand U7131 (N_7131,N_4636,N_4811);
and U7132 (N_7132,N_4691,N_5011);
or U7133 (N_7133,N_5844,N_4778);
or U7134 (N_7134,N_5419,N_4897);
and U7135 (N_7135,N_4753,N_4706);
nor U7136 (N_7136,N_5758,N_5498);
nor U7137 (N_7137,N_5783,N_4743);
and U7138 (N_7138,N_5078,N_5009);
and U7139 (N_7139,N_5997,N_5156);
nand U7140 (N_7140,N_4714,N_5371);
nand U7141 (N_7141,N_5809,N_5421);
and U7142 (N_7142,N_4799,N_5076);
and U7143 (N_7143,N_4681,N_5336);
nor U7144 (N_7144,N_4540,N_5106);
or U7145 (N_7145,N_5986,N_5485);
and U7146 (N_7146,N_5489,N_5680);
nor U7147 (N_7147,N_4953,N_5994);
or U7148 (N_7148,N_4576,N_5696);
or U7149 (N_7149,N_4571,N_4916);
and U7150 (N_7150,N_5888,N_4733);
nand U7151 (N_7151,N_5107,N_5394);
and U7152 (N_7152,N_5287,N_4891);
and U7153 (N_7153,N_4764,N_4557);
nand U7154 (N_7154,N_5779,N_4610);
or U7155 (N_7155,N_5433,N_5483);
nor U7156 (N_7156,N_4901,N_5928);
nor U7157 (N_7157,N_5675,N_5262);
or U7158 (N_7158,N_5121,N_4578);
nor U7159 (N_7159,N_4775,N_4753);
or U7160 (N_7160,N_5408,N_5687);
or U7161 (N_7161,N_4537,N_5374);
nand U7162 (N_7162,N_5211,N_5414);
or U7163 (N_7163,N_5312,N_4748);
or U7164 (N_7164,N_5495,N_5427);
or U7165 (N_7165,N_4981,N_5061);
nand U7166 (N_7166,N_5125,N_5526);
or U7167 (N_7167,N_4627,N_5001);
nand U7168 (N_7168,N_5420,N_5358);
nor U7169 (N_7169,N_4946,N_5997);
nor U7170 (N_7170,N_5105,N_5119);
nand U7171 (N_7171,N_5495,N_5432);
and U7172 (N_7172,N_5077,N_5732);
nand U7173 (N_7173,N_5359,N_5423);
and U7174 (N_7174,N_5247,N_5847);
or U7175 (N_7175,N_4896,N_5066);
and U7176 (N_7176,N_5840,N_5965);
or U7177 (N_7177,N_5122,N_5518);
or U7178 (N_7178,N_5082,N_4836);
nand U7179 (N_7179,N_5448,N_4897);
nor U7180 (N_7180,N_5651,N_5564);
and U7181 (N_7181,N_5094,N_5613);
and U7182 (N_7182,N_4552,N_4540);
and U7183 (N_7183,N_5548,N_4634);
and U7184 (N_7184,N_5731,N_4527);
and U7185 (N_7185,N_4733,N_4925);
and U7186 (N_7186,N_4624,N_4682);
nand U7187 (N_7187,N_5717,N_4519);
and U7188 (N_7188,N_5481,N_5054);
and U7189 (N_7189,N_5951,N_5773);
and U7190 (N_7190,N_4503,N_5810);
and U7191 (N_7191,N_4863,N_5685);
and U7192 (N_7192,N_4776,N_5272);
and U7193 (N_7193,N_5186,N_5791);
nand U7194 (N_7194,N_5186,N_4738);
and U7195 (N_7195,N_5145,N_5467);
or U7196 (N_7196,N_5858,N_5482);
or U7197 (N_7197,N_4599,N_5199);
and U7198 (N_7198,N_5587,N_5504);
nand U7199 (N_7199,N_5482,N_5254);
or U7200 (N_7200,N_5441,N_4582);
nor U7201 (N_7201,N_4700,N_5922);
nor U7202 (N_7202,N_5634,N_4721);
nand U7203 (N_7203,N_4789,N_4787);
nand U7204 (N_7204,N_5249,N_5010);
nand U7205 (N_7205,N_5846,N_5400);
and U7206 (N_7206,N_5203,N_4506);
and U7207 (N_7207,N_4530,N_4935);
and U7208 (N_7208,N_5385,N_5916);
nand U7209 (N_7209,N_5997,N_4822);
nand U7210 (N_7210,N_5092,N_5173);
and U7211 (N_7211,N_5446,N_4554);
or U7212 (N_7212,N_4879,N_4861);
or U7213 (N_7213,N_5788,N_4955);
or U7214 (N_7214,N_5960,N_4797);
nand U7215 (N_7215,N_5405,N_5428);
and U7216 (N_7216,N_5662,N_5188);
and U7217 (N_7217,N_4601,N_5872);
or U7218 (N_7218,N_4999,N_5844);
nor U7219 (N_7219,N_5446,N_4986);
and U7220 (N_7220,N_5082,N_4864);
nor U7221 (N_7221,N_4916,N_5579);
nand U7222 (N_7222,N_5630,N_5025);
nor U7223 (N_7223,N_5940,N_5650);
nand U7224 (N_7224,N_5952,N_5989);
or U7225 (N_7225,N_4700,N_4506);
and U7226 (N_7226,N_4521,N_5502);
or U7227 (N_7227,N_5534,N_4956);
nand U7228 (N_7228,N_4718,N_5955);
nand U7229 (N_7229,N_5582,N_5328);
nor U7230 (N_7230,N_5382,N_5189);
or U7231 (N_7231,N_5234,N_5691);
nand U7232 (N_7232,N_5064,N_5434);
nor U7233 (N_7233,N_5155,N_5750);
nor U7234 (N_7234,N_5566,N_5111);
nor U7235 (N_7235,N_4511,N_5860);
nor U7236 (N_7236,N_5078,N_4861);
xor U7237 (N_7237,N_4972,N_4997);
nand U7238 (N_7238,N_5274,N_5320);
nor U7239 (N_7239,N_5946,N_4950);
and U7240 (N_7240,N_5137,N_5890);
nor U7241 (N_7241,N_5735,N_5898);
and U7242 (N_7242,N_5379,N_5649);
nor U7243 (N_7243,N_4601,N_4933);
nor U7244 (N_7244,N_5416,N_5747);
nand U7245 (N_7245,N_5505,N_4621);
nand U7246 (N_7246,N_4574,N_5643);
and U7247 (N_7247,N_5772,N_4764);
or U7248 (N_7248,N_5528,N_5324);
nand U7249 (N_7249,N_5987,N_4710);
xor U7250 (N_7250,N_5813,N_5740);
and U7251 (N_7251,N_5330,N_4853);
nor U7252 (N_7252,N_4966,N_4644);
or U7253 (N_7253,N_5841,N_5025);
nand U7254 (N_7254,N_5095,N_4740);
nand U7255 (N_7255,N_5039,N_4623);
nor U7256 (N_7256,N_5643,N_4569);
or U7257 (N_7257,N_5906,N_5944);
nand U7258 (N_7258,N_5510,N_5020);
nor U7259 (N_7259,N_5467,N_5889);
nor U7260 (N_7260,N_5970,N_5978);
nor U7261 (N_7261,N_5405,N_4769);
nor U7262 (N_7262,N_4914,N_4910);
and U7263 (N_7263,N_5776,N_4735);
nor U7264 (N_7264,N_4937,N_5913);
nor U7265 (N_7265,N_5074,N_4836);
and U7266 (N_7266,N_5941,N_4779);
xor U7267 (N_7267,N_5657,N_5575);
xnor U7268 (N_7268,N_5183,N_4810);
nor U7269 (N_7269,N_5839,N_5887);
nor U7270 (N_7270,N_4591,N_5295);
or U7271 (N_7271,N_5556,N_5087);
or U7272 (N_7272,N_5794,N_4704);
and U7273 (N_7273,N_5699,N_4681);
or U7274 (N_7274,N_5684,N_5871);
and U7275 (N_7275,N_5150,N_4552);
and U7276 (N_7276,N_4630,N_5437);
nor U7277 (N_7277,N_4615,N_4670);
and U7278 (N_7278,N_5966,N_4731);
nor U7279 (N_7279,N_4940,N_5723);
or U7280 (N_7280,N_5185,N_5983);
nor U7281 (N_7281,N_4688,N_5713);
nand U7282 (N_7282,N_5845,N_5367);
nand U7283 (N_7283,N_4684,N_5969);
nand U7284 (N_7284,N_5414,N_4739);
and U7285 (N_7285,N_5025,N_4704);
and U7286 (N_7286,N_4942,N_4959);
or U7287 (N_7287,N_5928,N_5643);
nand U7288 (N_7288,N_5853,N_4751);
xnor U7289 (N_7289,N_4883,N_5246);
and U7290 (N_7290,N_5770,N_5439);
nand U7291 (N_7291,N_5524,N_5449);
or U7292 (N_7292,N_4579,N_5680);
nand U7293 (N_7293,N_5111,N_4558);
or U7294 (N_7294,N_4687,N_5652);
or U7295 (N_7295,N_5854,N_5413);
nand U7296 (N_7296,N_4619,N_4648);
or U7297 (N_7297,N_4513,N_4673);
or U7298 (N_7298,N_5273,N_4802);
and U7299 (N_7299,N_5689,N_4823);
nand U7300 (N_7300,N_4528,N_4502);
or U7301 (N_7301,N_4999,N_4848);
or U7302 (N_7302,N_5135,N_5506);
nor U7303 (N_7303,N_5610,N_4870);
or U7304 (N_7304,N_5482,N_5624);
nor U7305 (N_7305,N_5619,N_4684);
or U7306 (N_7306,N_5542,N_5551);
nand U7307 (N_7307,N_4570,N_5528);
nand U7308 (N_7308,N_5249,N_4589);
or U7309 (N_7309,N_5892,N_5533);
nor U7310 (N_7310,N_5918,N_5707);
or U7311 (N_7311,N_5021,N_5145);
nor U7312 (N_7312,N_5573,N_5654);
nand U7313 (N_7313,N_5809,N_4591);
or U7314 (N_7314,N_4583,N_5186);
or U7315 (N_7315,N_5069,N_5034);
nor U7316 (N_7316,N_5182,N_4910);
nand U7317 (N_7317,N_4515,N_4957);
xnor U7318 (N_7318,N_5770,N_5028);
nand U7319 (N_7319,N_5054,N_5766);
or U7320 (N_7320,N_4893,N_4568);
or U7321 (N_7321,N_5182,N_4591);
and U7322 (N_7322,N_5364,N_5070);
nor U7323 (N_7323,N_5640,N_5012);
or U7324 (N_7324,N_5065,N_5611);
nor U7325 (N_7325,N_5113,N_5702);
and U7326 (N_7326,N_5119,N_5133);
nand U7327 (N_7327,N_5724,N_4671);
and U7328 (N_7328,N_4715,N_5877);
nand U7329 (N_7329,N_5373,N_4515);
or U7330 (N_7330,N_5688,N_5392);
or U7331 (N_7331,N_5085,N_5507);
xor U7332 (N_7332,N_5719,N_5160);
nand U7333 (N_7333,N_4660,N_5644);
nor U7334 (N_7334,N_5545,N_5445);
or U7335 (N_7335,N_5335,N_5787);
xnor U7336 (N_7336,N_5415,N_4501);
nor U7337 (N_7337,N_5260,N_4674);
and U7338 (N_7338,N_5343,N_5900);
or U7339 (N_7339,N_4807,N_4957);
or U7340 (N_7340,N_4883,N_5921);
or U7341 (N_7341,N_4893,N_4528);
and U7342 (N_7342,N_5689,N_5891);
xnor U7343 (N_7343,N_5980,N_5561);
and U7344 (N_7344,N_5846,N_5066);
or U7345 (N_7345,N_5877,N_4765);
and U7346 (N_7346,N_5892,N_4746);
and U7347 (N_7347,N_5060,N_4732);
and U7348 (N_7348,N_4555,N_5071);
nand U7349 (N_7349,N_5763,N_4510);
and U7350 (N_7350,N_5737,N_4662);
nand U7351 (N_7351,N_5661,N_5340);
nor U7352 (N_7352,N_5077,N_4523);
nor U7353 (N_7353,N_5921,N_5889);
nand U7354 (N_7354,N_4921,N_4552);
xnor U7355 (N_7355,N_5881,N_4795);
or U7356 (N_7356,N_5699,N_5119);
or U7357 (N_7357,N_5981,N_4752);
nor U7358 (N_7358,N_4690,N_4612);
and U7359 (N_7359,N_4870,N_4980);
nor U7360 (N_7360,N_5930,N_4593);
nor U7361 (N_7361,N_5144,N_5939);
nand U7362 (N_7362,N_5088,N_5737);
and U7363 (N_7363,N_5857,N_5416);
nand U7364 (N_7364,N_4929,N_5387);
nand U7365 (N_7365,N_4912,N_4549);
and U7366 (N_7366,N_5417,N_5330);
and U7367 (N_7367,N_4662,N_4988);
nand U7368 (N_7368,N_4684,N_5507);
or U7369 (N_7369,N_5118,N_5189);
nand U7370 (N_7370,N_4822,N_5596);
nand U7371 (N_7371,N_5050,N_4581);
nor U7372 (N_7372,N_5425,N_5658);
or U7373 (N_7373,N_5660,N_4861);
nor U7374 (N_7374,N_5701,N_4951);
nor U7375 (N_7375,N_5318,N_5820);
nand U7376 (N_7376,N_4564,N_5576);
or U7377 (N_7377,N_5226,N_5029);
and U7378 (N_7378,N_4911,N_5098);
or U7379 (N_7379,N_4546,N_5297);
and U7380 (N_7380,N_5808,N_4742);
nor U7381 (N_7381,N_5123,N_5099);
nor U7382 (N_7382,N_5514,N_5702);
and U7383 (N_7383,N_5468,N_4629);
nand U7384 (N_7384,N_5041,N_4885);
or U7385 (N_7385,N_5396,N_4954);
or U7386 (N_7386,N_4998,N_5013);
and U7387 (N_7387,N_5244,N_5232);
or U7388 (N_7388,N_5714,N_4861);
nand U7389 (N_7389,N_5529,N_4851);
nand U7390 (N_7390,N_4794,N_5557);
and U7391 (N_7391,N_5931,N_5210);
nor U7392 (N_7392,N_5583,N_5278);
and U7393 (N_7393,N_4820,N_5190);
nand U7394 (N_7394,N_5925,N_4536);
and U7395 (N_7395,N_4677,N_5468);
xnor U7396 (N_7396,N_4608,N_5680);
and U7397 (N_7397,N_5080,N_5395);
and U7398 (N_7398,N_4738,N_5784);
nand U7399 (N_7399,N_5004,N_4523);
nor U7400 (N_7400,N_5004,N_5895);
and U7401 (N_7401,N_5246,N_4979);
or U7402 (N_7402,N_5809,N_4781);
and U7403 (N_7403,N_4984,N_4852);
nor U7404 (N_7404,N_5681,N_5314);
and U7405 (N_7405,N_5774,N_5299);
nor U7406 (N_7406,N_4532,N_4701);
or U7407 (N_7407,N_4587,N_4556);
nand U7408 (N_7408,N_5469,N_5546);
or U7409 (N_7409,N_5607,N_4928);
nor U7410 (N_7410,N_5436,N_5838);
nor U7411 (N_7411,N_4781,N_4573);
and U7412 (N_7412,N_4793,N_5534);
nor U7413 (N_7413,N_5809,N_5903);
and U7414 (N_7414,N_4941,N_4765);
nand U7415 (N_7415,N_5589,N_5531);
or U7416 (N_7416,N_5841,N_4625);
nand U7417 (N_7417,N_5213,N_5620);
or U7418 (N_7418,N_4676,N_4949);
and U7419 (N_7419,N_5501,N_5328);
nor U7420 (N_7420,N_4704,N_5646);
and U7421 (N_7421,N_5962,N_5854);
xor U7422 (N_7422,N_5391,N_4541);
nand U7423 (N_7423,N_4786,N_4972);
nand U7424 (N_7424,N_4983,N_5824);
nand U7425 (N_7425,N_4903,N_4790);
nand U7426 (N_7426,N_5609,N_4676);
or U7427 (N_7427,N_4828,N_4872);
and U7428 (N_7428,N_5339,N_5851);
or U7429 (N_7429,N_5393,N_5281);
or U7430 (N_7430,N_5814,N_5679);
nand U7431 (N_7431,N_5637,N_5682);
or U7432 (N_7432,N_4898,N_5386);
and U7433 (N_7433,N_5136,N_4904);
nor U7434 (N_7434,N_5103,N_5491);
nor U7435 (N_7435,N_5344,N_5644);
or U7436 (N_7436,N_4751,N_5838);
or U7437 (N_7437,N_4569,N_5347);
or U7438 (N_7438,N_5501,N_5453);
and U7439 (N_7439,N_5635,N_4964);
nor U7440 (N_7440,N_5590,N_5283);
nand U7441 (N_7441,N_4966,N_4905);
nor U7442 (N_7442,N_5123,N_4926);
nand U7443 (N_7443,N_4567,N_5308);
and U7444 (N_7444,N_5161,N_5500);
nand U7445 (N_7445,N_5832,N_4578);
and U7446 (N_7446,N_5160,N_5531);
nand U7447 (N_7447,N_5381,N_5328);
nand U7448 (N_7448,N_5658,N_4780);
nand U7449 (N_7449,N_4753,N_5111);
or U7450 (N_7450,N_5122,N_5676);
and U7451 (N_7451,N_4784,N_4569);
or U7452 (N_7452,N_4976,N_5132);
nor U7453 (N_7453,N_5965,N_5768);
nand U7454 (N_7454,N_5142,N_4625);
nor U7455 (N_7455,N_5834,N_5547);
and U7456 (N_7456,N_5061,N_5168);
and U7457 (N_7457,N_5948,N_5838);
or U7458 (N_7458,N_5087,N_4621);
nor U7459 (N_7459,N_4759,N_4673);
or U7460 (N_7460,N_4996,N_4542);
and U7461 (N_7461,N_4658,N_5655);
nand U7462 (N_7462,N_5718,N_5782);
nor U7463 (N_7463,N_5805,N_5548);
nor U7464 (N_7464,N_5152,N_4578);
nand U7465 (N_7465,N_5606,N_4683);
or U7466 (N_7466,N_4550,N_4600);
or U7467 (N_7467,N_5213,N_5494);
nand U7468 (N_7468,N_4595,N_5638);
or U7469 (N_7469,N_5121,N_4680);
nand U7470 (N_7470,N_4520,N_5514);
nand U7471 (N_7471,N_5446,N_5284);
nand U7472 (N_7472,N_4878,N_4850);
and U7473 (N_7473,N_5250,N_5936);
and U7474 (N_7474,N_4519,N_4648);
nor U7475 (N_7475,N_5500,N_5751);
or U7476 (N_7476,N_5104,N_4862);
nand U7477 (N_7477,N_5974,N_4734);
or U7478 (N_7478,N_4720,N_5467);
and U7479 (N_7479,N_5695,N_5104);
or U7480 (N_7480,N_4638,N_5626);
and U7481 (N_7481,N_5670,N_5323);
or U7482 (N_7482,N_5589,N_5937);
and U7483 (N_7483,N_5153,N_5374);
or U7484 (N_7484,N_5615,N_4846);
nor U7485 (N_7485,N_4620,N_4574);
or U7486 (N_7486,N_5693,N_4708);
or U7487 (N_7487,N_5128,N_5639);
xor U7488 (N_7488,N_5631,N_4673);
and U7489 (N_7489,N_5559,N_5454);
and U7490 (N_7490,N_4812,N_5459);
nand U7491 (N_7491,N_5281,N_5239);
and U7492 (N_7492,N_5048,N_5187);
nand U7493 (N_7493,N_5725,N_4588);
and U7494 (N_7494,N_4537,N_4890);
nor U7495 (N_7495,N_5708,N_5034);
nand U7496 (N_7496,N_5670,N_5731);
nand U7497 (N_7497,N_4767,N_5841);
nand U7498 (N_7498,N_5621,N_5858);
or U7499 (N_7499,N_5049,N_5730);
or U7500 (N_7500,N_6204,N_6960);
or U7501 (N_7501,N_6834,N_7267);
nor U7502 (N_7502,N_6701,N_6451);
or U7503 (N_7503,N_6624,N_6211);
or U7504 (N_7504,N_6547,N_7279);
and U7505 (N_7505,N_7300,N_6179);
and U7506 (N_7506,N_6231,N_6038);
or U7507 (N_7507,N_7348,N_6140);
or U7508 (N_7508,N_7098,N_7456);
nand U7509 (N_7509,N_6257,N_7159);
and U7510 (N_7510,N_6468,N_6275);
nor U7511 (N_7511,N_7027,N_6082);
nor U7512 (N_7512,N_6386,N_7012);
nor U7513 (N_7513,N_6956,N_7221);
and U7514 (N_7514,N_6183,N_6627);
or U7515 (N_7515,N_7170,N_6587);
nand U7516 (N_7516,N_7096,N_6943);
and U7517 (N_7517,N_7337,N_6288);
nor U7518 (N_7518,N_6004,N_6416);
nand U7519 (N_7519,N_7014,N_7296);
and U7520 (N_7520,N_7498,N_7403);
or U7521 (N_7521,N_7242,N_6518);
nor U7522 (N_7522,N_6088,N_6483);
and U7523 (N_7523,N_6768,N_6585);
nor U7524 (N_7524,N_7350,N_6448);
or U7525 (N_7525,N_6572,N_6605);
and U7526 (N_7526,N_6591,N_6337);
nand U7527 (N_7527,N_6678,N_6658);
nand U7528 (N_7528,N_6042,N_6548);
and U7529 (N_7529,N_7390,N_7317);
nand U7530 (N_7530,N_6796,N_6091);
and U7531 (N_7531,N_6311,N_6266);
xnor U7532 (N_7532,N_6393,N_6463);
and U7533 (N_7533,N_7460,N_6002);
nor U7534 (N_7534,N_7053,N_6623);
and U7535 (N_7535,N_6663,N_7410);
nor U7536 (N_7536,N_7357,N_6369);
nand U7537 (N_7537,N_7040,N_6356);
nand U7538 (N_7538,N_6064,N_7274);
and U7539 (N_7539,N_6688,N_6824);
nand U7540 (N_7540,N_6090,N_6374);
and U7541 (N_7541,N_7062,N_6783);
and U7542 (N_7542,N_6507,N_7203);
nand U7543 (N_7543,N_6175,N_7426);
and U7544 (N_7544,N_6509,N_6519);
or U7545 (N_7545,N_6757,N_6776);
xor U7546 (N_7546,N_6437,N_6270);
and U7547 (N_7547,N_7257,N_7404);
nor U7548 (N_7548,N_6214,N_7320);
and U7549 (N_7549,N_6735,N_7204);
nor U7550 (N_7550,N_6366,N_7429);
and U7551 (N_7551,N_6722,N_6282);
and U7552 (N_7552,N_7104,N_6223);
or U7553 (N_7553,N_6084,N_6992);
nor U7554 (N_7554,N_6839,N_6945);
or U7555 (N_7555,N_7189,N_6545);
and U7556 (N_7556,N_6309,N_6018);
or U7557 (N_7557,N_7111,N_6077);
nor U7558 (N_7558,N_6474,N_7361);
and U7559 (N_7559,N_7423,N_6492);
and U7560 (N_7560,N_6958,N_6613);
nand U7561 (N_7561,N_7022,N_7194);
and U7562 (N_7562,N_6449,N_7230);
nand U7563 (N_7563,N_7331,N_6712);
nor U7564 (N_7564,N_7121,N_6932);
nor U7565 (N_7565,N_7285,N_6316);
or U7566 (N_7566,N_6893,N_7029);
or U7567 (N_7567,N_7148,N_6740);
or U7568 (N_7568,N_6693,N_7123);
nand U7569 (N_7569,N_7491,N_7328);
nor U7570 (N_7570,N_6075,N_6680);
nand U7571 (N_7571,N_6329,N_6138);
or U7572 (N_7572,N_6597,N_7037);
nand U7573 (N_7573,N_7118,N_6926);
and U7574 (N_7574,N_7011,N_6767);
nand U7575 (N_7575,N_7050,N_7485);
nor U7576 (N_7576,N_6130,N_6836);
nor U7577 (N_7577,N_6953,N_6383);
nand U7578 (N_7578,N_6788,N_6814);
nor U7579 (N_7579,N_6041,N_6418);
nor U7580 (N_7580,N_7464,N_7499);
or U7581 (N_7581,N_7487,N_7327);
nor U7582 (N_7582,N_6330,N_7420);
or U7583 (N_7583,N_6901,N_6208);
or U7584 (N_7584,N_7442,N_6424);
nor U7585 (N_7585,N_7183,N_6685);
nor U7586 (N_7586,N_7018,N_6125);
nand U7587 (N_7587,N_6371,N_6124);
nor U7588 (N_7588,N_7085,N_6970);
nand U7589 (N_7589,N_6738,N_6924);
and U7590 (N_7590,N_6414,N_6011);
nor U7591 (N_7591,N_6941,N_6340);
and U7592 (N_7592,N_6060,N_6532);
nand U7593 (N_7593,N_6874,N_6840);
and U7594 (N_7594,N_6989,N_6898);
or U7595 (N_7595,N_7351,N_6095);
nor U7596 (N_7596,N_7115,N_7192);
xor U7597 (N_7597,N_7056,N_6017);
nor U7598 (N_7598,N_6906,N_7241);
or U7599 (N_7599,N_6595,N_6219);
nor U7600 (N_7600,N_7432,N_7474);
and U7601 (N_7601,N_7117,N_6710);
or U7602 (N_7602,N_6815,N_7278);
and U7603 (N_7603,N_6037,N_6111);
nor U7604 (N_7604,N_6935,N_6035);
and U7605 (N_7605,N_6149,N_7217);
or U7606 (N_7606,N_6599,N_6045);
and U7607 (N_7607,N_6640,N_6147);
and U7608 (N_7608,N_6671,N_7273);
or U7609 (N_7609,N_6016,N_7075);
nor U7610 (N_7610,N_7486,N_6559);
and U7611 (N_7611,N_6533,N_6864);
nand U7612 (N_7612,N_7389,N_6165);
nor U7613 (N_7613,N_6803,N_6733);
or U7614 (N_7614,N_6642,N_6446);
nor U7615 (N_7615,N_7400,N_6635);
or U7616 (N_7616,N_7301,N_6283);
nand U7617 (N_7617,N_6452,N_6494);
and U7618 (N_7618,N_6552,N_7231);
or U7619 (N_7619,N_6965,N_7476);
or U7620 (N_7620,N_6290,N_7377);
nor U7621 (N_7621,N_7174,N_7421);
or U7622 (N_7622,N_7019,N_7459);
nand U7623 (N_7623,N_6305,N_7413);
nor U7624 (N_7624,N_7411,N_6825);
nor U7625 (N_7625,N_7463,N_6749);
and U7626 (N_7626,N_6530,N_6539);
nor U7627 (N_7627,N_6698,N_7313);
or U7628 (N_7628,N_6476,N_7276);
nor U7629 (N_7629,N_6308,N_7190);
nand U7630 (N_7630,N_7065,N_6745);
and U7631 (N_7631,N_6729,N_7295);
and U7632 (N_7632,N_6441,N_6537);
nand U7633 (N_7633,N_6774,N_6368);
or U7634 (N_7634,N_6040,N_6873);
nand U7635 (N_7635,N_6114,N_6780);
nand U7636 (N_7636,N_7240,N_6860);
nand U7637 (N_7637,N_6569,N_6711);
nand U7638 (N_7638,N_7478,N_6234);
and U7639 (N_7639,N_7051,N_6215);
or U7640 (N_7640,N_6927,N_6382);
and U7641 (N_7641,N_6500,N_7154);
nor U7642 (N_7642,N_6076,N_6473);
nor U7643 (N_7643,N_6736,N_6080);
nor U7644 (N_7644,N_7344,N_7430);
nor U7645 (N_7645,N_6412,N_6348);
nand U7646 (N_7646,N_7316,N_7208);
nor U7647 (N_7647,N_7439,N_7108);
and U7648 (N_7648,N_6431,N_6364);
and U7649 (N_7649,N_7393,N_6489);
or U7650 (N_7650,N_6122,N_7319);
or U7651 (N_7651,N_7131,N_6352);
or U7652 (N_7652,N_7071,N_6370);
nand U7653 (N_7653,N_7153,N_6996);
or U7654 (N_7654,N_7307,N_6297);
nand U7655 (N_7655,N_7150,N_6723);
nor U7656 (N_7656,N_6194,N_6377);
xor U7657 (N_7657,N_6339,N_7223);
nand U7658 (N_7658,N_6438,N_7347);
and U7659 (N_7659,N_6510,N_6014);
or U7660 (N_7660,N_6968,N_6844);
nor U7661 (N_7661,N_7321,N_7110);
nand U7662 (N_7662,N_7196,N_6287);
nor U7663 (N_7663,N_6879,N_6020);
nand U7664 (N_7664,N_6246,N_6975);
nor U7665 (N_7665,N_6294,N_7286);
or U7666 (N_7666,N_6912,N_6575);
or U7667 (N_7667,N_6400,N_7372);
and U7668 (N_7668,N_6614,N_6944);
and U7669 (N_7669,N_7078,N_6074);
nor U7670 (N_7670,N_6931,N_6302);
nand U7671 (N_7671,N_6265,N_7314);
and U7672 (N_7672,N_6062,N_7323);
and U7673 (N_7673,N_7382,N_7338);
xnor U7674 (N_7674,N_7120,N_7472);
and U7675 (N_7675,N_6579,N_6612);
nand U7676 (N_7676,N_6966,N_7101);
or U7677 (N_7677,N_6065,N_6460);
nor U7678 (N_7678,N_6816,N_6871);
and U7679 (N_7679,N_6779,N_7132);
or U7680 (N_7680,N_6154,N_6319);
and U7681 (N_7681,N_6362,N_6972);
nand U7682 (N_7682,N_6029,N_7137);
nor U7683 (N_7683,N_6298,N_7253);
nor U7684 (N_7684,N_6505,N_6962);
and U7685 (N_7685,N_6028,N_7356);
nand U7686 (N_7686,N_6728,N_6771);
or U7687 (N_7687,N_6413,N_6067);
and U7688 (N_7688,N_6556,N_7205);
xnor U7689 (N_7689,N_6869,N_7090);
or U7690 (N_7690,N_6128,N_6508);
and U7691 (N_7691,N_7184,N_6358);
nor U7692 (N_7692,N_7122,N_6964);
nand U7693 (N_7693,N_6727,N_6333);
nor U7694 (N_7694,N_7368,N_6529);
and U7695 (N_7695,N_7144,N_7129);
nor U7696 (N_7696,N_7312,N_6315);
or U7697 (N_7697,N_6566,N_7471);
nand U7698 (N_7698,N_6230,N_6027);
or U7699 (N_7699,N_7450,N_7431);
nand U7700 (N_7700,N_6984,N_6379);
nor U7701 (N_7701,N_6127,N_6544);
and U7702 (N_7702,N_6625,N_6969);
and U7703 (N_7703,N_6520,N_6359);
or U7704 (N_7704,N_6044,N_6367);
nand U7705 (N_7705,N_6577,N_6744);
nand U7706 (N_7706,N_6439,N_6596);
and U7707 (N_7707,N_6527,N_6714);
or U7708 (N_7708,N_6630,N_7467);
nand U7709 (N_7709,N_7335,N_6583);
or U7710 (N_7710,N_6853,N_7399);
nand U7711 (N_7711,N_6903,N_7023);
and U7712 (N_7712,N_6240,N_6787);
and U7713 (N_7713,N_6645,N_6277);
nand U7714 (N_7714,N_7156,N_6541);
and U7715 (N_7715,N_7255,N_6391);
or U7716 (N_7716,N_7169,N_6096);
and U7717 (N_7717,N_6797,N_6528);
nand U7718 (N_7718,N_6925,N_7172);
or U7719 (N_7719,N_6899,N_7398);
and U7720 (N_7720,N_6250,N_6313);
nand U7721 (N_7721,N_6506,N_6481);
or U7722 (N_7722,N_6497,N_6905);
nor U7723 (N_7723,N_6677,N_6328);
or U7724 (N_7724,N_6480,N_7305);
nor U7725 (N_7725,N_6521,N_7161);
or U7726 (N_7726,N_6963,N_6974);
nand U7727 (N_7727,N_7353,N_7375);
or U7728 (N_7728,N_6785,N_6856);
nor U7729 (N_7729,N_7376,N_6551);
or U7730 (N_7730,N_6058,N_7256);
nand U7731 (N_7731,N_6929,N_7374);
or U7732 (N_7732,N_6571,N_6775);
or U7733 (N_7733,N_6024,N_7386);
nor U7734 (N_7734,N_6384,N_6542);
nand U7735 (N_7735,N_6877,N_6454);
and U7736 (N_7736,N_6408,N_7373);
nand U7737 (N_7737,N_6007,N_6565);
and U7738 (N_7738,N_6069,N_6900);
and U7739 (N_7739,N_7366,N_6472);
and U7740 (N_7740,N_7187,N_6440);
or U7741 (N_7741,N_6576,N_6743);
nand U7742 (N_7742,N_6828,N_6887);
nor U7743 (N_7743,N_6716,N_6152);
and U7744 (N_7744,N_6255,N_7220);
nor U7745 (N_7745,N_7381,N_6057);
and U7746 (N_7746,N_6657,N_7440);
nor U7747 (N_7747,N_7039,N_7292);
nand U7748 (N_7748,N_6610,N_7270);
nor U7749 (N_7749,N_6669,N_6350);
nor U7750 (N_7750,N_6885,N_7482);
nor U7751 (N_7751,N_7036,N_6636);
and U7752 (N_7752,N_6469,N_6433);
nor U7753 (N_7753,N_7497,N_6137);
or U7754 (N_7754,N_6694,N_7182);
and U7755 (N_7755,N_6267,N_6558);
or U7756 (N_7756,N_6055,N_6388);
nor U7757 (N_7757,N_7162,N_6664);
and U7758 (N_7758,N_7380,N_6692);
and U7759 (N_7759,N_6911,N_6849);
nor U7760 (N_7760,N_6616,N_6325);
and U7761 (N_7761,N_6253,N_6564);
or U7762 (N_7762,N_6638,N_7128);
or U7763 (N_7763,N_7343,N_6052);
and U7764 (N_7764,N_7433,N_7007);
nand U7765 (N_7765,N_6777,N_6380);
and U7766 (N_7766,N_6923,N_6419);
nor U7767 (N_7767,N_6063,N_6157);
and U7768 (N_7768,N_6602,N_7177);
nor U7769 (N_7769,N_7477,N_6649);
or U7770 (N_7770,N_6643,N_6731);
nor U7771 (N_7771,N_6718,N_6878);
and U7772 (N_7772,N_6346,N_7297);
and U7773 (N_7773,N_6994,N_6141);
xor U7774 (N_7774,N_6155,N_6462);
nor U7775 (N_7775,N_7151,N_6392);
and U7776 (N_7776,N_6502,N_6739);
nor U7777 (N_7777,N_6724,N_7070);
nor U7778 (N_7778,N_7202,N_6407);
or U7779 (N_7779,N_7239,N_6991);
or U7780 (N_7780,N_7214,N_6237);
or U7781 (N_7781,N_6707,N_6485);
or U7782 (N_7782,N_7416,N_6523);
nand U7783 (N_7783,N_6951,N_6162);
and U7784 (N_7784,N_7138,N_6593);
nor U7785 (N_7785,N_6800,N_7142);
or U7786 (N_7786,N_6784,N_6660);
nand U7787 (N_7787,N_6586,N_7406);
or U7788 (N_7788,N_7346,N_7139);
or U7789 (N_7789,N_6928,N_7315);
and U7790 (N_7790,N_6273,N_7063);
and U7791 (N_7791,N_7141,N_7355);
nor U7792 (N_7792,N_6952,N_7397);
or U7793 (N_7793,N_6910,N_7052);
or U7794 (N_7794,N_6227,N_6228);
nand U7795 (N_7795,N_6977,N_7146);
or U7796 (N_7796,N_7035,N_6031);
or U7797 (N_7797,N_6673,N_7290);
or U7798 (N_7798,N_6381,N_6160);
nor U7799 (N_7799,N_6226,N_6332);
xnor U7800 (N_7800,N_7311,N_7195);
nor U7801 (N_7801,N_6517,N_6801);
and U7802 (N_7802,N_7457,N_7147);
and U7803 (N_7803,N_6713,N_7445);
and U7804 (N_7804,N_6734,N_7193);
nand U7805 (N_7805,N_7059,N_6761);
or U7806 (N_7806,N_6837,N_6904);
and U7807 (N_7807,N_7309,N_7465);
and U7808 (N_7808,N_6135,N_6661);
or U7809 (N_7809,N_7082,N_6026);
nand U7810 (N_7810,N_6192,N_6631);
or U7811 (N_7811,N_6396,N_6628);
or U7812 (N_7812,N_7124,N_6998);
and U7813 (N_7813,N_6808,N_6335);
and U7814 (N_7814,N_6511,N_6758);
nand U7815 (N_7815,N_6292,N_7001);
and U7816 (N_7816,N_6608,N_7268);
or U7817 (N_7817,N_6865,N_6197);
and U7818 (N_7818,N_6009,N_7009);
nand U7819 (N_7819,N_6762,N_6487);
nor U7820 (N_7820,N_7114,N_6322);
nor U7821 (N_7821,N_6882,N_6184);
and U7822 (N_7822,N_7178,N_6493);
and U7823 (N_7823,N_6909,N_6676);
and U7824 (N_7824,N_6567,N_7074);
nand U7825 (N_7825,N_6299,N_6401);
or U7826 (N_7826,N_6034,N_7045);
and U7827 (N_7827,N_6447,N_6629);
nand U7828 (N_7828,N_7013,N_6913);
nand U7829 (N_7829,N_6444,N_6997);
nor U7830 (N_7830,N_6557,N_7244);
nand U7831 (N_7831,N_7469,N_7281);
or U7832 (N_7832,N_7054,N_6217);
and U7833 (N_7833,N_7383,N_7125);
nand U7834 (N_7834,N_6831,N_6251);
nand U7835 (N_7835,N_6751,N_7091);
nand U7836 (N_7836,N_6106,N_6225);
nor U7837 (N_7837,N_6023,N_7489);
nor U7838 (N_7838,N_7370,N_6888);
xor U7839 (N_7839,N_6786,N_7167);
nand U7840 (N_7840,N_6512,N_6540);
or U7841 (N_7841,N_7107,N_6046);
nand U7842 (N_7842,N_7447,N_6684);
and U7843 (N_7843,N_7483,N_6142);
or U7844 (N_7844,N_6870,N_6987);
nand U7845 (N_7845,N_6458,N_6405);
nand U7846 (N_7846,N_7248,N_6104);
or U7847 (N_7847,N_6915,N_7302);
nor U7848 (N_7848,N_6752,N_6363);
and U7849 (N_7849,N_7448,N_7032);
or U7850 (N_7850,N_7043,N_7378);
or U7851 (N_7851,N_7462,N_7152);
nor U7852 (N_7852,N_7210,N_7102);
nand U7853 (N_7853,N_7234,N_6134);
or U7854 (N_7854,N_6536,N_6372);
and U7855 (N_7855,N_6349,N_6159);
and U7856 (N_7856,N_6341,N_6897);
and U7857 (N_7857,N_7233,N_6107);
nor U7858 (N_7858,N_7158,N_6939);
and U7859 (N_7859,N_7160,N_6504);
nand U7860 (N_7860,N_6272,N_6798);
and U7861 (N_7861,N_7261,N_6222);
nor U7862 (N_7862,N_6973,N_6553);
nand U7863 (N_7863,N_6429,N_7046);
nand U7864 (N_7864,N_6056,N_6889);
and U7865 (N_7865,N_6570,N_6967);
nand U7866 (N_7866,N_6995,N_6830);
and U7867 (N_7867,N_6102,N_6666);
nand U7868 (N_7868,N_7330,N_7222);
or U7869 (N_7869,N_7112,N_6687);
nand U7870 (N_7870,N_6858,N_6872);
and U7871 (N_7871,N_7092,N_7095);
nor U7872 (N_7872,N_6902,N_7494);
and U7873 (N_7873,N_7003,N_7488);
nand U7874 (N_7874,N_6121,N_6005);
nor U7875 (N_7875,N_7047,N_6703);
nand U7876 (N_7876,N_6286,N_6232);
or U7877 (N_7877,N_6705,N_6804);
nor U7878 (N_7878,N_7069,N_6262);
nor U7879 (N_7879,N_6229,N_6813);
and U7880 (N_7880,N_6248,N_6061);
or U7881 (N_7881,N_6478,N_7435);
or U7882 (N_7882,N_6675,N_6496);
nor U7883 (N_7883,N_7226,N_7392);
or U7884 (N_7884,N_6531,N_6886);
nand U7885 (N_7885,N_7310,N_6269);
or U7886 (N_7886,N_7164,N_6948);
and U7887 (N_7887,N_6659,N_6933);
or U7888 (N_7888,N_7388,N_7219);
and U7889 (N_7889,N_6279,N_6730);
and U7890 (N_7890,N_7237,N_7004);
nor U7891 (N_7891,N_6765,N_6003);
or U7892 (N_7892,N_7033,N_7318);
and U7893 (N_7893,N_7289,N_6781);
nor U7894 (N_7894,N_7198,N_7466);
nor U7895 (N_7895,N_6950,N_6621);
nor U7896 (N_7896,N_6841,N_6647);
or U7897 (N_7897,N_7280,N_6216);
nand U7898 (N_7898,N_6148,N_6515);
and U7899 (N_7899,N_6054,N_6750);
or U7900 (N_7900,N_6012,N_7298);
and U7901 (N_7901,N_6182,N_6385);
or U7902 (N_7902,N_6049,N_7266);
nand U7903 (N_7903,N_7171,N_7496);
and U7904 (N_7904,N_7087,N_6456);
nand U7905 (N_7905,N_6829,N_6174);
nand U7906 (N_7906,N_6000,N_6030);
nor U7907 (N_7907,N_6741,N_6826);
nor U7908 (N_7908,N_6940,N_6862);
nor U7909 (N_7909,N_7209,N_6854);
nand U7910 (N_7910,N_6013,N_6985);
and U7911 (N_7911,N_6696,N_7490);
nand U7912 (N_7912,N_6524,N_7395);
nor U7913 (N_7913,N_6453,N_6598);
and U7914 (N_7914,N_6938,N_7017);
nand U7915 (N_7915,N_6086,N_6592);
nor U7916 (N_7916,N_6426,N_7049);
nor U7917 (N_7917,N_7345,N_6981);
nand U7918 (N_7918,N_6395,N_6151);
and U7919 (N_7919,N_6285,N_6499);
and U7920 (N_7920,N_6327,N_6525);
nand U7921 (N_7921,N_6241,N_6810);
nor U7922 (N_7922,N_6113,N_6619);
nand U7923 (N_7923,N_7354,N_7021);
or U7924 (N_7924,N_6561,N_6318);
and U7925 (N_7925,N_6347,N_6185);
nor U7926 (N_7926,N_6891,N_6947);
nor U7927 (N_7927,N_7271,N_6930);
or U7928 (N_7928,N_6978,N_6725);
nand U7929 (N_7929,N_6772,N_6001);
or U7930 (N_7930,N_6846,N_6450);
or U7931 (N_7931,N_6143,N_6207);
or U7932 (N_7932,N_6809,N_6880);
nor U7933 (N_7933,N_6156,N_6291);
nor U7934 (N_7934,N_7088,N_7264);
nor U7935 (N_7935,N_6171,N_6949);
or U7936 (N_7936,N_6161,N_6847);
nor U7937 (N_7937,N_6656,N_7133);
nand U7938 (N_7938,N_6890,N_6976);
or U7939 (N_7939,N_6868,N_7005);
and U7940 (N_7940,N_6916,N_7369);
nand U7941 (N_7941,N_6081,N_6129);
or U7942 (N_7942,N_6176,N_6832);
or U7943 (N_7943,N_6420,N_6373);
nand U7944 (N_7944,N_7106,N_7409);
or U7945 (N_7945,N_6793,N_7275);
or U7946 (N_7946,N_7006,N_7042);
and U7947 (N_7947,N_6236,N_6015);
nor U7948 (N_7948,N_6402,N_7365);
nand U7949 (N_7949,N_7250,N_6306);
or U7950 (N_7950,N_6312,N_6674);
nand U7951 (N_7951,N_6079,N_7304);
and U7952 (N_7952,N_7197,N_6549);
and U7953 (N_7953,N_6099,N_7484);
nor U7954 (N_7954,N_6189,N_7434);
and U7955 (N_7955,N_7444,N_7436);
nand U7956 (N_7956,N_6908,N_7402);
nor U7957 (N_7957,N_6097,N_7061);
and U7958 (N_7958,N_7455,N_6195);
nand U7959 (N_7959,N_7135,N_7099);
nor U7960 (N_7960,N_7084,N_6427);
and U7961 (N_7961,N_7140,N_6261);
and U7962 (N_7962,N_7385,N_6150);
and U7963 (N_7963,N_6178,N_6957);
nor U7964 (N_7964,N_6699,N_7339);
and U7965 (N_7965,N_6823,N_6344);
and U7966 (N_7966,N_6522,N_6875);
nand U7967 (N_7967,N_7028,N_6503);
nor U7968 (N_7968,N_6415,N_6430);
nand U7969 (N_7969,N_6833,N_7294);
nand U7970 (N_7970,N_7438,N_6295);
or U7971 (N_7971,N_7468,N_7324);
nor U7972 (N_7972,N_6859,N_6259);
nand U7973 (N_7973,N_7058,N_6618);
nor U7974 (N_7974,N_6158,N_6554);
and U7975 (N_7975,N_6353,N_6720);
nor U7976 (N_7976,N_7419,N_7360);
and U7977 (N_7977,N_6988,N_6342);
and U7978 (N_7978,N_6651,N_6633);
nor U7979 (N_7979,N_6971,N_6284);
nor U7980 (N_7980,N_7422,N_6445);
or U7981 (N_7981,N_6146,N_6555);
xnor U7982 (N_7982,N_7081,N_6220);
or U7983 (N_7983,N_6094,N_7470);
or U7984 (N_7984,N_6498,N_6357);
or U7985 (N_7985,N_6177,N_7026);
nand U7986 (N_7986,N_6389,N_6486);
and U7987 (N_7987,N_7149,N_6457);
nand U7988 (N_7988,N_6378,N_7245);
or U7989 (N_7989,N_6406,N_7079);
nor U7990 (N_7990,N_7265,N_7227);
or U7991 (N_7991,N_6442,N_6239);
nor U7992 (N_7992,N_7405,N_6668);
and U7993 (N_7993,N_7113,N_6690);
nor U7994 (N_7994,N_7341,N_6033);
or U7995 (N_7995,N_6048,N_7322);
nand U7996 (N_7996,N_6857,N_6737);
nor U7997 (N_7997,N_6748,N_6314);
nor U7998 (N_7998,N_6403,N_6594);
nor U7999 (N_7999,N_6764,N_6578);
nor U8000 (N_8000,N_7401,N_6213);
nor U8001 (N_8001,N_7407,N_7340);
or U8002 (N_8002,N_6863,N_6773);
nand U8003 (N_8003,N_7452,N_6186);
and U8004 (N_8004,N_6068,N_7349);
and U8005 (N_8005,N_6098,N_7030);
and U8006 (N_8006,N_7086,N_7415);
and U8007 (N_8007,N_7130,N_6986);
nand U8008 (N_8008,N_6802,N_7126);
and U8009 (N_8009,N_6746,N_6936);
nor U8010 (N_8010,N_6163,N_6360);
or U8011 (N_8011,N_6488,N_6200);
nor U8012 (N_8012,N_6717,N_7427);
and U8013 (N_8013,N_6345,N_7020);
nand U8014 (N_8014,N_6101,N_6550);
nand U8015 (N_8015,N_6534,N_7200);
nand U8016 (N_8016,N_7394,N_7229);
nand U8017 (N_8017,N_6820,N_6025);
nor U8018 (N_8018,N_6654,N_7287);
nand U8019 (N_8019,N_7443,N_7097);
nor U8020 (N_8020,N_7364,N_7105);
nand U8021 (N_8021,N_6907,N_7277);
nand U8022 (N_8022,N_7191,N_6050);
and U8023 (N_8023,N_6807,N_7119);
and U8024 (N_8024,N_6324,N_7263);
nand U8025 (N_8025,N_7048,N_6100);
or U8026 (N_8026,N_7473,N_6085);
and U8027 (N_8027,N_6274,N_6181);
and U8028 (N_8028,N_7024,N_6980);
nand U8029 (N_8029,N_6336,N_6895);
nor U8030 (N_8030,N_6838,N_6700);
nor U8031 (N_8031,N_6421,N_6709);
or U8032 (N_8032,N_7475,N_6256);
nand U8033 (N_8033,N_6848,N_7358);
xnor U8034 (N_8034,N_6387,N_6747);
or U8035 (N_8035,N_7283,N_6193);
and U8036 (N_8036,N_6109,N_6582);
or U8037 (N_8037,N_6238,N_6047);
nand U8038 (N_8038,N_6589,N_7165);
or U8039 (N_8039,N_6855,N_6632);
and U8040 (N_8040,N_6679,N_6805);
nor U8041 (N_8041,N_6573,N_6852);
nor U8042 (N_8042,N_7299,N_6683);
nand U8043 (N_8043,N_6410,N_6172);
or U8044 (N_8044,N_7408,N_6959);
nor U8045 (N_8045,N_7016,N_7038);
and U8046 (N_8046,N_7057,N_6702);
nor U8047 (N_8047,N_6376,N_6249);
nor U8048 (N_8048,N_7002,N_7067);
or U8049 (N_8049,N_6112,N_7175);
nor U8050 (N_8050,N_6770,N_6320);
and U8051 (N_8051,N_6766,N_7143);
nand U8052 (N_8052,N_7068,N_6580);
nor U8053 (N_8053,N_6708,N_6326);
or U8054 (N_8054,N_6252,N_6490);
and U8055 (N_8055,N_6119,N_6317);
and U8056 (N_8056,N_7044,N_7163);
and U8057 (N_8057,N_6817,N_6861);
nor U8058 (N_8058,N_6351,N_6188);
or U8059 (N_8059,N_6423,N_6914);
and U8060 (N_8060,N_6338,N_7185);
nand U8061 (N_8061,N_6268,N_6584);
and U8062 (N_8062,N_6411,N_6681);
and U8063 (N_8063,N_7181,N_6168);
nand U8064 (N_8064,N_6417,N_6942);
nor U8065 (N_8065,N_7212,N_6422);
nand U8066 (N_8066,N_6600,N_6235);
or U8067 (N_8067,N_6842,N_6546);
nor U8068 (N_8068,N_6982,N_6394);
and U8069 (N_8069,N_6021,N_7293);
or U8070 (N_8070,N_7232,N_7428);
and U8071 (N_8071,N_7333,N_6078);
and U8072 (N_8072,N_6110,N_6670);
or U8073 (N_8073,N_6535,N_7359);
nor U8074 (N_8074,N_7254,N_7417);
or U8075 (N_8075,N_6581,N_7103);
or U8076 (N_8076,N_6242,N_6721);
nand U8077 (N_8077,N_6131,N_7288);
and U8078 (N_8078,N_7247,N_7213);
nand U8079 (N_8079,N_6954,N_7493);
or U8080 (N_8080,N_6513,N_6611);
and U8081 (N_8081,N_6881,N_6894);
nor U8082 (N_8082,N_7235,N_6843);
and U8083 (N_8083,N_6477,N_6759);
and U8084 (N_8084,N_6922,N_6271);
nor U8085 (N_8085,N_7173,N_6514);
nor U8086 (N_8086,N_6008,N_6845);
and U8087 (N_8087,N_6867,N_6233);
nand U8088 (N_8088,N_7396,N_6646);
nor U8089 (N_8089,N_6365,N_6672);
or U8090 (N_8090,N_6092,N_7243);
or U8091 (N_8091,N_7201,N_7387);
nor U8092 (N_8092,N_6662,N_6300);
and U8093 (N_8093,N_6032,N_6301);
or U8094 (N_8094,N_6918,N_7093);
nor U8095 (N_8095,N_6484,N_6244);
nor U8096 (N_8096,N_6153,N_7480);
nand U8097 (N_8097,N_6247,N_6467);
nor U8098 (N_8098,N_7246,N_6704);
nand U8099 (N_8099,N_6568,N_6999);
or U8100 (N_8100,N_6115,N_7176);
and U8101 (N_8101,N_6756,N_6221);
nand U8102 (N_8102,N_6053,N_6655);
nor U8103 (N_8103,N_7199,N_6432);
nor U8104 (N_8104,N_6398,N_6397);
nor U8105 (N_8105,N_7034,N_7325);
and U8106 (N_8106,N_6258,N_7166);
and U8107 (N_8107,N_6203,N_6732);
nor U8108 (N_8108,N_6126,N_6117);
nor U8109 (N_8109,N_7258,N_6822);
nor U8110 (N_8110,N_6205,N_7449);
nand U8111 (N_8111,N_7269,N_6218);
nor U8112 (N_8112,N_6039,N_7262);
or U8113 (N_8113,N_6920,N_7060);
and U8114 (N_8114,N_6209,N_6850);
xnor U8115 (N_8115,N_6281,N_7329);
nor U8116 (N_8116,N_7157,N_7249);
nand U8117 (N_8117,N_6116,N_6799);
or U8118 (N_8118,N_6491,N_6620);
nor U8119 (N_8119,N_6173,N_7481);
or U8120 (N_8120,N_7225,N_6790);
nand U8121 (N_8121,N_7260,N_7259);
or U8122 (N_8122,N_6639,N_6212);
nor U8123 (N_8123,N_6726,N_7492);
and U8124 (N_8124,N_6390,N_6083);
or U8125 (N_8125,N_6070,N_6145);
nand U8126 (N_8126,N_6763,N_6202);
nor U8127 (N_8127,N_6409,N_6166);
nor U8128 (N_8128,N_7424,N_7215);
nand U8129 (N_8129,N_6425,N_6190);
nand U8130 (N_8130,N_6955,N_6404);
and U8131 (N_8131,N_6892,N_6466);
nand U8132 (N_8132,N_6601,N_6778);
or U8133 (N_8133,N_6634,N_6224);
nor U8134 (N_8134,N_6051,N_6667);
nor U8135 (N_8135,N_6876,N_6697);
xnor U8136 (N_8136,N_7282,N_7224);
or U8137 (N_8137,N_7100,N_7116);
or U8138 (N_8138,N_7216,N_6133);
and U8139 (N_8139,N_7384,N_7008);
or U8140 (N_8140,N_7458,N_6435);
and U8141 (N_8141,N_6648,N_7109);
nand U8142 (N_8142,N_6132,N_6071);
or U8143 (N_8143,N_6590,N_6755);
and U8144 (N_8144,N_6979,N_7211);
nand U8145 (N_8145,N_6198,N_6543);
and U8146 (N_8146,N_7418,N_6334);
and U8147 (N_8147,N_7425,N_7168);
nand U8148 (N_8148,N_6361,N_6470);
nand U8149 (N_8149,N_6459,N_6818);
or U8150 (N_8150,N_7251,N_6812);
or U8151 (N_8151,N_6622,N_6883);
nand U8152 (N_8152,N_7180,N_6921);
nand U8153 (N_8153,N_6089,N_7454);
nand U8154 (N_8154,N_6303,N_7238);
nand U8155 (N_8155,N_7072,N_7077);
or U8156 (N_8156,N_6754,N_6574);
or U8157 (N_8157,N_7363,N_6010);
or U8158 (N_8158,N_6293,N_7080);
or U8159 (N_8159,N_6169,N_7303);
or U8160 (N_8160,N_7308,N_7186);
nor U8161 (N_8161,N_6495,N_6310);
and U8162 (N_8162,N_6103,N_6461);
nand U8163 (N_8163,N_6073,N_6245);
nand U8164 (N_8164,N_7145,N_6123);
and U8165 (N_8165,N_7437,N_6652);
and U8166 (N_8166,N_6795,N_6760);
nand U8167 (N_8167,N_6615,N_6604);
nor U8168 (N_8168,N_6607,N_6170);
or U8169 (N_8169,N_6896,N_6617);
nand U8170 (N_8170,N_6917,N_7218);
nand U8171 (N_8171,N_6637,N_6689);
nand U8172 (N_8172,N_6375,N_6254);
or U8173 (N_8173,N_7155,N_6206);
xnor U8174 (N_8174,N_6276,N_6479);
nand U8175 (N_8175,N_7055,N_6851);
nand U8176 (N_8176,N_7412,N_6465);
nand U8177 (N_8177,N_6821,N_7252);
or U8178 (N_8178,N_6196,N_7451);
or U8179 (N_8179,N_6343,N_6835);
nand U8180 (N_8180,N_7188,N_6782);
nand U8181 (N_8181,N_6562,N_6354);
or U8182 (N_8182,N_7025,N_6501);
nand U8183 (N_8183,N_6043,N_7228);
nand U8184 (N_8184,N_7306,N_7272);
nor U8185 (N_8185,N_6139,N_7066);
and U8186 (N_8186,N_6072,N_6471);
nor U8187 (N_8187,N_6264,N_6792);
or U8188 (N_8188,N_6641,N_7207);
or U8189 (N_8189,N_7332,N_6191);
or U8190 (N_8190,N_6482,N_6682);
and U8191 (N_8191,N_6819,N_6443);
nor U8192 (N_8192,N_6120,N_6475);
nand U8193 (N_8193,N_6019,N_6789);
and U8194 (N_8194,N_6983,N_6428);
nor U8195 (N_8195,N_6199,N_6136);
nand U8196 (N_8196,N_6210,N_6323);
or U8197 (N_8197,N_6087,N_6105);
nand U8198 (N_8198,N_6606,N_6108);
nor U8199 (N_8199,N_6937,N_7089);
and U8200 (N_8200,N_7371,N_7414);
nor U8201 (N_8201,N_7031,N_6464);
nor U8202 (N_8202,N_6455,N_6243);
nor U8203 (N_8203,N_6434,N_6827);
or U8204 (N_8204,N_6516,N_7367);
or U8205 (N_8205,N_6066,N_7094);
nor U8206 (N_8206,N_7015,N_6866);
and U8207 (N_8207,N_7336,N_6990);
and U8208 (N_8208,N_6180,N_7134);
nand U8209 (N_8209,N_7379,N_6644);
or U8210 (N_8210,N_6144,N_6695);
or U8211 (N_8211,N_7041,N_7352);
nand U8212 (N_8212,N_6560,N_6946);
and U8213 (N_8213,N_6653,N_6588);
nor U8214 (N_8214,N_6769,N_6289);
nand U8215 (N_8215,N_7326,N_7495);
and U8216 (N_8216,N_7453,N_6603);
and U8217 (N_8217,N_6650,N_6260);
and U8218 (N_8218,N_6563,N_6626);
and U8219 (N_8219,N_6742,N_7064);
and U8220 (N_8220,N_7010,N_7000);
nor U8221 (N_8221,N_6753,N_6201);
nor U8222 (N_8222,N_7136,N_7479);
nor U8223 (N_8223,N_6934,N_6059);
or U8224 (N_8224,N_7206,N_6436);
nor U8225 (N_8225,N_7127,N_7076);
nand U8226 (N_8226,N_6280,N_6691);
nor U8227 (N_8227,N_7284,N_6296);
nand U8228 (N_8228,N_6036,N_6919);
or U8229 (N_8229,N_6006,N_6355);
nor U8230 (N_8230,N_6167,N_6706);
and U8231 (N_8231,N_7236,N_7073);
nor U8232 (N_8232,N_7461,N_6715);
nand U8233 (N_8233,N_6609,N_6263);
or U8234 (N_8234,N_7342,N_6719);
or U8235 (N_8235,N_7291,N_6794);
nand U8236 (N_8236,N_7362,N_6884);
nor U8237 (N_8237,N_6993,N_6187);
nor U8238 (N_8238,N_7441,N_6526);
or U8239 (N_8239,N_7083,N_6278);
nor U8240 (N_8240,N_6811,N_6399);
nand U8241 (N_8241,N_7334,N_7179);
or U8242 (N_8242,N_6304,N_7446);
or U8243 (N_8243,N_6961,N_6806);
or U8244 (N_8244,N_6307,N_6791);
and U8245 (N_8245,N_6665,N_6538);
or U8246 (N_8246,N_6093,N_6164);
nor U8247 (N_8247,N_6118,N_6686);
nand U8248 (N_8248,N_6331,N_7391);
nor U8249 (N_8249,N_6321,N_6022);
nor U8250 (N_8250,N_6591,N_6941);
or U8251 (N_8251,N_6508,N_6365);
nor U8252 (N_8252,N_6026,N_7262);
nor U8253 (N_8253,N_6574,N_6198);
nand U8254 (N_8254,N_6928,N_7020);
and U8255 (N_8255,N_7022,N_7448);
nand U8256 (N_8256,N_6958,N_7363);
or U8257 (N_8257,N_7214,N_7114);
nand U8258 (N_8258,N_7061,N_6382);
and U8259 (N_8259,N_6769,N_6918);
and U8260 (N_8260,N_6930,N_7083);
or U8261 (N_8261,N_7082,N_6876);
nor U8262 (N_8262,N_6695,N_6762);
or U8263 (N_8263,N_6514,N_6301);
and U8264 (N_8264,N_6217,N_6239);
or U8265 (N_8265,N_6065,N_6549);
nand U8266 (N_8266,N_6597,N_6231);
nor U8267 (N_8267,N_6644,N_6166);
or U8268 (N_8268,N_6033,N_6047);
nand U8269 (N_8269,N_6459,N_7034);
nor U8270 (N_8270,N_6210,N_7214);
nor U8271 (N_8271,N_6308,N_7482);
or U8272 (N_8272,N_6217,N_7235);
or U8273 (N_8273,N_6278,N_6195);
and U8274 (N_8274,N_6643,N_6492);
or U8275 (N_8275,N_6627,N_6530);
nor U8276 (N_8276,N_6690,N_6234);
or U8277 (N_8277,N_6306,N_6756);
or U8278 (N_8278,N_6283,N_6726);
and U8279 (N_8279,N_6527,N_6346);
nand U8280 (N_8280,N_6445,N_6183);
and U8281 (N_8281,N_6972,N_6912);
or U8282 (N_8282,N_6858,N_7380);
nand U8283 (N_8283,N_6791,N_6880);
nor U8284 (N_8284,N_7333,N_6272);
nor U8285 (N_8285,N_7113,N_6610);
nor U8286 (N_8286,N_6597,N_6446);
and U8287 (N_8287,N_6662,N_6427);
or U8288 (N_8288,N_6765,N_7019);
nor U8289 (N_8289,N_7413,N_7467);
nor U8290 (N_8290,N_6027,N_6406);
xor U8291 (N_8291,N_6506,N_7445);
nor U8292 (N_8292,N_6761,N_6404);
or U8293 (N_8293,N_6714,N_6372);
xor U8294 (N_8294,N_7078,N_7334);
nor U8295 (N_8295,N_6206,N_7040);
nand U8296 (N_8296,N_6301,N_6543);
or U8297 (N_8297,N_6338,N_6531);
or U8298 (N_8298,N_7221,N_6685);
or U8299 (N_8299,N_7093,N_7204);
and U8300 (N_8300,N_6232,N_6590);
and U8301 (N_8301,N_7067,N_6800);
xnor U8302 (N_8302,N_6024,N_7380);
nor U8303 (N_8303,N_7211,N_6977);
xnor U8304 (N_8304,N_6860,N_7040);
nor U8305 (N_8305,N_6125,N_6771);
and U8306 (N_8306,N_6094,N_7432);
and U8307 (N_8307,N_6079,N_6346);
nor U8308 (N_8308,N_6284,N_7489);
nor U8309 (N_8309,N_6112,N_6368);
and U8310 (N_8310,N_6782,N_7476);
nand U8311 (N_8311,N_7001,N_7428);
and U8312 (N_8312,N_6836,N_6116);
or U8313 (N_8313,N_6952,N_6245);
or U8314 (N_8314,N_6511,N_6359);
or U8315 (N_8315,N_7163,N_6015);
and U8316 (N_8316,N_6955,N_6194);
nor U8317 (N_8317,N_6019,N_6908);
nor U8318 (N_8318,N_7292,N_6170);
nand U8319 (N_8319,N_6227,N_6765);
nor U8320 (N_8320,N_7421,N_6342);
or U8321 (N_8321,N_7326,N_6151);
or U8322 (N_8322,N_6031,N_6916);
nor U8323 (N_8323,N_7308,N_6121);
or U8324 (N_8324,N_6728,N_6734);
nor U8325 (N_8325,N_6457,N_7416);
and U8326 (N_8326,N_6941,N_6199);
nor U8327 (N_8327,N_6587,N_7008);
nor U8328 (N_8328,N_7132,N_6543);
or U8329 (N_8329,N_7422,N_6430);
or U8330 (N_8330,N_7490,N_6318);
nor U8331 (N_8331,N_6572,N_6833);
and U8332 (N_8332,N_6480,N_6948);
nand U8333 (N_8333,N_6756,N_6166);
nor U8334 (N_8334,N_7332,N_7385);
nor U8335 (N_8335,N_6948,N_6596);
nor U8336 (N_8336,N_6084,N_6248);
nand U8337 (N_8337,N_6701,N_7424);
nor U8338 (N_8338,N_6709,N_7109);
nor U8339 (N_8339,N_6523,N_6899);
nor U8340 (N_8340,N_6901,N_6872);
nand U8341 (N_8341,N_6545,N_7285);
and U8342 (N_8342,N_6186,N_6131);
nand U8343 (N_8343,N_7018,N_7139);
and U8344 (N_8344,N_6718,N_6694);
nor U8345 (N_8345,N_6356,N_7068);
nand U8346 (N_8346,N_6943,N_6895);
nor U8347 (N_8347,N_6647,N_6580);
nor U8348 (N_8348,N_7130,N_7299);
nor U8349 (N_8349,N_7366,N_6210);
nand U8350 (N_8350,N_6128,N_6264);
or U8351 (N_8351,N_6524,N_7477);
and U8352 (N_8352,N_6648,N_6219);
nor U8353 (N_8353,N_6466,N_6941);
nor U8354 (N_8354,N_7076,N_6093);
nand U8355 (N_8355,N_6468,N_7157);
and U8356 (N_8356,N_6183,N_6630);
or U8357 (N_8357,N_6056,N_6426);
or U8358 (N_8358,N_7127,N_6486);
nor U8359 (N_8359,N_7452,N_6964);
nor U8360 (N_8360,N_7059,N_6872);
and U8361 (N_8361,N_7341,N_7031);
nand U8362 (N_8362,N_6312,N_6875);
nor U8363 (N_8363,N_6428,N_6714);
or U8364 (N_8364,N_6154,N_7371);
nand U8365 (N_8365,N_6879,N_7164);
and U8366 (N_8366,N_7024,N_7489);
nand U8367 (N_8367,N_6368,N_6786);
nand U8368 (N_8368,N_7210,N_6938);
nor U8369 (N_8369,N_6760,N_7238);
nand U8370 (N_8370,N_6252,N_7257);
nand U8371 (N_8371,N_6669,N_6153);
nor U8372 (N_8372,N_6025,N_6764);
or U8373 (N_8373,N_7122,N_7084);
or U8374 (N_8374,N_7147,N_6359);
nand U8375 (N_8375,N_6802,N_6091);
nor U8376 (N_8376,N_6165,N_6930);
nor U8377 (N_8377,N_6533,N_6148);
or U8378 (N_8378,N_6949,N_7315);
nand U8379 (N_8379,N_6341,N_7083);
nor U8380 (N_8380,N_7142,N_7360);
xor U8381 (N_8381,N_7179,N_6671);
nand U8382 (N_8382,N_6410,N_6974);
and U8383 (N_8383,N_6468,N_6523);
and U8384 (N_8384,N_7473,N_6105);
nand U8385 (N_8385,N_6491,N_7012);
nand U8386 (N_8386,N_6991,N_6861);
or U8387 (N_8387,N_6621,N_7096);
and U8388 (N_8388,N_6414,N_7361);
nand U8389 (N_8389,N_6530,N_6262);
or U8390 (N_8390,N_7046,N_6887);
nand U8391 (N_8391,N_6241,N_6857);
or U8392 (N_8392,N_6039,N_6612);
and U8393 (N_8393,N_6468,N_6093);
and U8394 (N_8394,N_6765,N_7454);
or U8395 (N_8395,N_6596,N_6974);
xnor U8396 (N_8396,N_6969,N_6837);
or U8397 (N_8397,N_7044,N_7190);
nor U8398 (N_8398,N_6799,N_7138);
nor U8399 (N_8399,N_7037,N_6902);
nor U8400 (N_8400,N_6855,N_7341);
nor U8401 (N_8401,N_6331,N_7483);
nor U8402 (N_8402,N_6526,N_6229);
nand U8403 (N_8403,N_6211,N_6145);
and U8404 (N_8404,N_6068,N_6970);
nor U8405 (N_8405,N_6830,N_6210);
nor U8406 (N_8406,N_7345,N_6950);
or U8407 (N_8407,N_7313,N_6970);
and U8408 (N_8408,N_7446,N_6201);
nor U8409 (N_8409,N_6041,N_6899);
nor U8410 (N_8410,N_7167,N_6271);
and U8411 (N_8411,N_6113,N_6108);
xnor U8412 (N_8412,N_6815,N_6866);
or U8413 (N_8413,N_6403,N_6132);
nor U8414 (N_8414,N_6084,N_6841);
or U8415 (N_8415,N_6811,N_7478);
and U8416 (N_8416,N_7186,N_7364);
nor U8417 (N_8417,N_6441,N_7172);
or U8418 (N_8418,N_6803,N_7269);
or U8419 (N_8419,N_6458,N_6144);
nor U8420 (N_8420,N_7204,N_7144);
or U8421 (N_8421,N_7498,N_6155);
or U8422 (N_8422,N_7088,N_7166);
or U8423 (N_8423,N_7160,N_7230);
nand U8424 (N_8424,N_6817,N_7484);
nand U8425 (N_8425,N_6226,N_6074);
nand U8426 (N_8426,N_7218,N_6574);
nor U8427 (N_8427,N_7376,N_6107);
nand U8428 (N_8428,N_6420,N_6390);
or U8429 (N_8429,N_6364,N_6128);
nand U8430 (N_8430,N_7243,N_6097);
and U8431 (N_8431,N_6491,N_6935);
and U8432 (N_8432,N_6772,N_6445);
and U8433 (N_8433,N_7312,N_6841);
nor U8434 (N_8434,N_6420,N_6871);
nor U8435 (N_8435,N_6167,N_6110);
and U8436 (N_8436,N_6359,N_6759);
or U8437 (N_8437,N_7190,N_7104);
nand U8438 (N_8438,N_6260,N_7309);
or U8439 (N_8439,N_6981,N_6948);
nand U8440 (N_8440,N_7413,N_7258);
nand U8441 (N_8441,N_6581,N_7208);
and U8442 (N_8442,N_6285,N_7380);
or U8443 (N_8443,N_7214,N_6373);
or U8444 (N_8444,N_6741,N_6889);
or U8445 (N_8445,N_7481,N_7107);
nor U8446 (N_8446,N_7210,N_6797);
nand U8447 (N_8447,N_7479,N_7471);
nor U8448 (N_8448,N_6359,N_6718);
or U8449 (N_8449,N_6039,N_7268);
nand U8450 (N_8450,N_6090,N_6078);
nor U8451 (N_8451,N_6206,N_6231);
or U8452 (N_8452,N_6811,N_7055);
and U8453 (N_8453,N_7452,N_7176);
and U8454 (N_8454,N_7285,N_6681);
and U8455 (N_8455,N_6771,N_6763);
and U8456 (N_8456,N_7323,N_7499);
nand U8457 (N_8457,N_6323,N_6806);
and U8458 (N_8458,N_6361,N_6106);
or U8459 (N_8459,N_7132,N_6523);
or U8460 (N_8460,N_6109,N_6123);
nor U8461 (N_8461,N_6263,N_6403);
or U8462 (N_8462,N_7249,N_7242);
nor U8463 (N_8463,N_7186,N_6300);
and U8464 (N_8464,N_7463,N_6043);
nand U8465 (N_8465,N_6725,N_7350);
or U8466 (N_8466,N_6356,N_7377);
or U8467 (N_8467,N_6092,N_7035);
and U8468 (N_8468,N_6755,N_6406);
or U8469 (N_8469,N_6432,N_6180);
or U8470 (N_8470,N_6963,N_6891);
or U8471 (N_8471,N_7044,N_6554);
and U8472 (N_8472,N_6885,N_6718);
nand U8473 (N_8473,N_6462,N_7151);
nor U8474 (N_8474,N_6353,N_6778);
nor U8475 (N_8475,N_6331,N_7489);
nand U8476 (N_8476,N_6467,N_6747);
and U8477 (N_8477,N_6583,N_6471);
nor U8478 (N_8478,N_6926,N_7377);
and U8479 (N_8479,N_6006,N_6282);
nand U8480 (N_8480,N_6352,N_6643);
or U8481 (N_8481,N_6422,N_7083);
nand U8482 (N_8482,N_6944,N_6963);
nor U8483 (N_8483,N_7432,N_6351);
nor U8484 (N_8484,N_6182,N_7238);
nand U8485 (N_8485,N_7328,N_7481);
nand U8486 (N_8486,N_6874,N_7230);
nand U8487 (N_8487,N_7036,N_6815);
and U8488 (N_8488,N_6328,N_7270);
and U8489 (N_8489,N_7354,N_6861);
and U8490 (N_8490,N_6178,N_7147);
and U8491 (N_8491,N_6997,N_6293);
nor U8492 (N_8492,N_6777,N_6227);
nor U8493 (N_8493,N_7024,N_6180);
nor U8494 (N_8494,N_7192,N_7342);
nor U8495 (N_8495,N_6089,N_6304);
nand U8496 (N_8496,N_6138,N_7437);
nor U8497 (N_8497,N_6192,N_6364);
nor U8498 (N_8498,N_6948,N_7229);
or U8499 (N_8499,N_6652,N_7493);
nand U8500 (N_8500,N_6222,N_6084);
nand U8501 (N_8501,N_7411,N_7060);
nor U8502 (N_8502,N_7322,N_7349);
and U8503 (N_8503,N_6972,N_7421);
nor U8504 (N_8504,N_6229,N_6891);
or U8505 (N_8505,N_6747,N_7282);
or U8506 (N_8506,N_6814,N_7381);
or U8507 (N_8507,N_6898,N_7184);
nand U8508 (N_8508,N_6639,N_7073);
or U8509 (N_8509,N_7014,N_7137);
or U8510 (N_8510,N_6723,N_6803);
and U8511 (N_8511,N_6876,N_7063);
or U8512 (N_8512,N_7291,N_6592);
nor U8513 (N_8513,N_7188,N_7331);
and U8514 (N_8514,N_6007,N_6774);
and U8515 (N_8515,N_7432,N_6539);
nand U8516 (N_8516,N_6561,N_6295);
nor U8517 (N_8517,N_6658,N_6145);
nand U8518 (N_8518,N_7279,N_7147);
nor U8519 (N_8519,N_6210,N_6458);
and U8520 (N_8520,N_7048,N_6860);
nor U8521 (N_8521,N_7164,N_6863);
or U8522 (N_8522,N_7168,N_7188);
and U8523 (N_8523,N_6079,N_6446);
and U8524 (N_8524,N_6237,N_7014);
nand U8525 (N_8525,N_7360,N_6046);
or U8526 (N_8526,N_7248,N_7032);
or U8527 (N_8527,N_6492,N_6353);
and U8528 (N_8528,N_6317,N_7329);
nand U8529 (N_8529,N_6677,N_6737);
nor U8530 (N_8530,N_6487,N_6436);
or U8531 (N_8531,N_6859,N_7179);
or U8532 (N_8532,N_7362,N_6768);
nor U8533 (N_8533,N_6882,N_7455);
nor U8534 (N_8534,N_6443,N_6289);
and U8535 (N_8535,N_7111,N_6193);
and U8536 (N_8536,N_6501,N_6619);
or U8537 (N_8537,N_6123,N_6506);
and U8538 (N_8538,N_7398,N_7081);
and U8539 (N_8539,N_7384,N_7113);
or U8540 (N_8540,N_6641,N_6584);
nand U8541 (N_8541,N_6241,N_6218);
nand U8542 (N_8542,N_6339,N_6617);
and U8543 (N_8543,N_7045,N_6012);
nor U8544 (N_8544,N_6281,N_6088);
nand U8545 (N_8545,N_7038,N_6432);
nand U8546 (N_8546,N_6217,N_6094);
nor U8547 (N_8547,N_6810,N_6722);
or U8548 (N_8548,N_6911,N_6693);
xnor U8549 (N_8549,N_6851,N_6602);
and U8550 (N_8550,N_6758,N_7139);
nand U8551 (N_8551,N_7190,N_6368);
or U8552 (N_8552,N_6881,N_6433);
nor U8553 (N_8553,N_6275,N_6743);
and U8554 (N_8554,N_7159,N_6210);
and U8555 (N_8555,N_6504,N_6630);
and U8556 (N_8556,N_6299,N_6834);
nand U8557 (N_8557,N_7497,N_6605);
and U8558 (N_8558,N_6276,N_6843);
and U8559 (N_8559,N_7152,N_6611);
nand U8560 (N_8560,N_6537,N_6174);
xnor U8561 (N_8561,N_6373,N_7127);
and U8562 (N_8562,N_6192,N_6567);
or U8563 (N_8563,N_6968,N_6351);
nand U8564 (N_8564,N_6892,N_7350);
nand U8565 (N_8565,N_6637,N_6427);
and U8566 (N_8566,N_6561,N_6011);
or U8567 (N_8567,N_6020,N_7493);
and U8568 (N_8568,N_6846,N_6912);
or U8569 (N_8569,N_6325,N_6254);
nand U8570 (N_8570,N_6802,N_6631);
and U8571 (N_8571,N_6206,N_6592);
and U8572 (N_8572,N_6241,N_6631);
nand U8573 (N_8573,N_7435,N_6380);
nand U8574 (N_8574,N_6442,N_6405);
nor U8575 (N_8575,N_6654,N_6309);
nor U8576 (N_8576,N_6600,N_6014);
nand U8577 (N_8577,N_7110,N_6518);
or U8578 (N_8578,N_6977,N_7373);
nor U8579 (N_8579,N_7422,N_6527);
or U8580 (N_8580,N_6540,N_6995);
nand U8581 (N_8581,N_6360,N_6330);
and U8582 (N_8582,N_6362,N_6823);
nand U8583 (N_8583,N_6270,N_6414);
and U8584 (N_8584,N_6657,N_7123);
and U8585 (N_8585,N_6797,N_6620);
nor U8586 (N_8586,N_7250,N_6277);
nand U8587 (N_8587,N_6903,N_6095);
and U8588 (N_8588,N_6646,N_6193);
nor U8589 (N_8589,N_7402,N_6023);
or U8590 (N_8590,N_7328,N_6761);
or U8591 (N_8591,N_7070,N_6396);
and U8592 (N_8592,N_6471,N_6480);
or U8593 (N_8593,N_6177,N_7234);
nor U8594 (N_8594,N_6330,N_6078);
xnor U8595 (N_8595,N_7241,N_6793);
nor U8596 (N_8596,N_7279,N_6004);
or U8597 (N_8597,N_6285,N_6482);
nand U8598 (N_8598,N_7180,N_7120);
nor U8599 (N_8599,N_6634,N_6219);
nand U8600 (N_8600,N_6659,N_6660);
nand U8601 (N_8601,N_6127,N_6939);
nand U8602 (N_8602,N_7138,N_6730);
nor U8603 (N_8603,N_6502,N_6938);
or U8604 (N_8604,N_6794,N_7411);
nand U8605 (N_8605,N_6611,N_6017);
nor U8606 (N_8606,N_6122,N_6601);
nor U8607 (N_8607,N_7175,N_6391);
nor U8608 (N_8608,N_7418,N_6182);
or U8609 (N_8609,N_7278,N_6667);
or U8610 (N_8610,N_6256,N_6915);
nand U8611 (N_8611,N_6671,N_6217);
or U8612 (N_8612,N_6146,N_6297);
nand U8613 (N_8613,N_6089,N_7175);
and U8614 (N_8614,N_7392,N_6329);
nand U8615 (N_8615,N_6979,N_6341);
nor U8616 (N_8616,N_7098,N_6720);
or U8617 (N_8617,N_7422,N_7414);
nor U8618 (N_8618,N_7195,N_6472);
xor U8619 (N_8619,N_6891,N_6923);
and U8620 (N_8620,N_6295,N_6934);
nor U8621 (N_8621,N_6305,N_6831);
and U8622 (N_8622,N_7394,N_6794);
or U8623 (N_8623,N_6035,N_7044);
and U8624 (N_8624,N_7087,N_6208);
and U8625 (N_8625,N_6499,N_6811);
nor U8626 (N_8626,N_6224,N_6741);
nor U8627 (N_8627,N_6067,N_7341);
nand U8628 (N_8628,N_7020,N_6972);
nand U8629 (N_8629,N_6987,N_6125);
xor U8630 (N_8630,N_6499,N_6971);
and U8631 (N_8631,N_6622,N_6012);
and U8632 (N_8632,N_6462,N_6271);
nand U8633 (N_8633,N_7196,N_6110);
nand U8634 (N_8634,N_7079,N_6787);
and U8635 (N_8635,N_6686,N_7258);
nor U8636 (N_8636,N_6611,N_6782);
nor U8637 (N_8637,N_7377,N_7073);
nor U8638 (N_8638,N_7436,N_6454);
or U8639 (N_8639,N_7107,N_6650);
and U8640 (N_8640,N_7090,N_6930);
nand U8641 (N_8641,N_7348,N_6874);
and U8642 (N_8642,N_6932,N_7288);
nand U8643 (N_8643,N_7080,N_6923);
nor U8644 (N_8644,N_7134,N_6785);
nor U8645 (N_8645,N_7451,N_7302);
nand U8646 (N_8646,N_7217,N_6182);
nand U8647 (N_8647,N_6425,N_7096);
nand U8648 (N_8648,N_7258,N_6273);
nand U8649 (N_8649,N_7149,N_6317);
nand U8650 (N_8650,N_6327,N_6242);
or U8651 (N_8651,N_7201,N_7345);
nor U8652 (N_8652,N_7237,N_6533);
nand U8653 (N_8653,N_7102,N_6347);
nand U8654 (N_8654,N_7135,N_6545);
or U8655 (N_8655,N_7278,N_6573);
or U8656 (N_8656,N_6264,N_7040);
nand U8657 (N_8657,N_6995,N_7359);
nand U8658 (N_8658,N_6238,N_6403);
nand U8659 (N_8659,N_6897,N_7044);
and U8660 (N_8660,N_6125,N_7034);
and U8661 (N_8661,N_6507,N_6485);
nor U8662 (N_8662,N_7459,N_6027);
nand U8663 (N_8663,N_7019,N_6369);
or U8664 (N_8664,N_6763,N_7229);
nand U8665 (N_8665,N_7069,N_6961);
nand U8666 (N_8666,N_7258,N_6487);
nand U8667 (N_8667,N_7036,N_7172);
or U8668 (N_8668,N_7291,N_6750);
and U8669 (N_8669,N_6209,N_7088);
nor U8670 (N_8670,N_7150,N_6565);
nand U8671 (N_8671,N_7409,N_6721);
nor U8672 (N_8672,N_6446,N_6045);
nor U8673 (N_8673,N_6201,N_7336);
nor U8674 (N_8674,N_7032,N_6831);
or U8675 (N_8675,N_6893,N_7023);
nor U8676 (N_8676,N_7068,N_6079);
nor U8677 (N_8677,N_6221,N_7157);
nand U8678 (N_8678,N_6593,N_6674);
nand U8679 (N_8679,N_6566,N_6459);
nand U8680 (N_8680,N_7344,N_6941);
nor U8681 (N_8681,N_6346,N_6206);
or U8682 (N_8682,N_7178,N_6157);
nand U8683 (N_8683,N_6065,N_6199);
xor U8684 (N_8684,N_7330,N_6098);
nand U8685 (N_8685,N_7277,N_6392);
and U8686 (N_8686,N_6266,N_6098);
and U8687 (N_8687,N_6782,N_6271);
nand U8688 (N_8688,N_7431,N_7282);
or U8689 (N_8689,N_6698,N_6651);
nand U8690 (N_8690,N_6195,N_6718);
nor U8691 (N_8691,N_6871,N_7261);
and U8692 (N_8692,N_7161,N_7084);
nor U8693 (N_8693,N_6182,N_6084);
and U8694 (N_8694,N_6389,N_6717);
nor U8695 (N_8695,N_6820,N_7189);
and U8696 (N_8696,N_6618,N_7381);
nor U8697 (N_8697,N_6209,N_6371);
and U8698 (N_8698,N_6681,N_6870);
nand U8699 (N_8699,N_6440,N_7266);
or U8700 (N_8700,N_6590,N_6414);
nand U8701 (N_8701,N_6918,N_7106);
xor U8702 (N_8702,N_6955,N_7200);
or U8703 (N_8703,N_6007,N_6557);
nand U8704 (N_8704,N_7329,N_7016);
nor U8705 (N_8705,N_6511,N_6065);
or U8706 (N_8706,N_6080,N_6396);
or U8707 (N_8707,N_6273,N_7425);
or U8708 (N_8708,N_6052,N_7173);
or U8709 (N_8709,N_7297,N_6748);
nor U8710 (N_8710,N_6221,N_6398);
or U8711 (N_8711,N_6255,N_7321);
xor U8712 (N_8712,N_6333,N_7287);
or U8713 (N_8713,N_7450,N_7250);
nand U8714 (N_8714,N_6890,N_6645);
and U8715 (N_8715,N_7295,N_6096);
nor U8716 (N_8716,N_6709,N_6150);
nor U8717 (N_8717,N_7008,N_6013);
and U8718 (N_8718,N_6193,N_6190);
nand U8719 (N_8719,N_7090,N_7264);
nand U8720 (N_8720,N_6860,N_7257);
nor U8721 (N_8721,N_6111,N_6945);
nor U8722 (N_8722,N_6386,N_6968);
or U8723 (N_8723,N_6954,N_6184);
nand U8724 (N_8724,N_6274,N_6085);
and U8725 (N_8725,N_6789,N_6621);
and U8726 (N_8726,N_6007,N_6863);
or U8727 (N_8727,N_6437,N_6340);
and U8728 (N_8728,N_7409,N_6174);
and U8729 (N_8729,N_6345,N_6009);
nand U8730 (N_8730,N_6412,N_6815);
or U8731 (N_8731,N_6781,N_6244);
and U8732 (N_8732,N_6934,N_6262);
and U8733 (N_8733,N_6644,N_7272);
nor U8734 (N_8734,N_6437,N_6469);
nor U8735 (N_8735,N_6286,N_7489);
nor U8736 (N_8736,N_6025,N_6955);
nor U8737 (N_8737,N_6622,N_6938);
nand U8738 (N_8738,N_7013,N_6460);
nor U8739 (N_8739,N_7435,N_6251);
or U8740 (N_8740,N_6555,N_6678);
nor U8741 (N_8741,N_7433,N_7300);
or U8742 (N_8742,N_6291,N_6339);
or U8743 (N_8743,N_6742,N_7370);
nor U8744 (N_8744,N_6839,N_6087);
and U8745 (N_8745,N_6279,N_6485);
and U8746 (N_8746,N_6110,N_6096);
nand U8747 (N_8747,N_7428,N_6211);
nor U8748 (N_8748,N_7177,N_6091);
or U8749 (N_8749,N_6306,N_7168);
and U8750 (N_8750,N_6115,N_6675);
and U8751 (N_8751,N_6618,N_6815);
nor U8752 (N_8752,N_6421,N_7382);
nor U8753 (N_8753,N_7184,N_6928);
or U8754 (N_8754,N_6374,N_7499);
and U8755 (N_8755,N_6099,N_6264);
nand U8756 (N_8756,N_6448,N_7431);
or U8757 (N_8757,N_7045,N_6614);
or U8758 (N_8758,N_7279,N_7486);
nand U8759 (N_8759,N_6321,N_6357);
nor U8760 (N_8760,N_6061,N_7157);
nor U8761 (N_8761,N_6969,N_6304);
or U8762 (N_8762,N_6572,N_7246);
and U8763 (N_8763,N_6782,N_6190);
or U8764 (N_8764,N_6552,N_7002);
or U8765 (N_8765,N_6074,N_6048);
nand U8766 (N_8766,N_6310,N_6866);
and U8767 (N_8767,N_6815,N_6424);
nand U8768 (N_8768,N_6283,N_7403);
nand U8769 (N_8769,N_7335,N_6111);
nor U8770 (N_8770,N_6065,N_6340);
or U8771 (N_8771,N_6169,N_6139);
or U8772 (N_8772,N_6491,N_6275);
or U8773 (N_8773,N_7318,N_6261);
and U8774 (N_8774,N_7286,N_6730);
and U8775 (N_8775,N_6599,N_6777);
or U8776 (N_8776,N_7041,N_7204);
nand U8777 (N_8777,N_6609,N_6407);
or U8778 (N_8778,N_7084,N_6995);
nor U8779 (N_8779,N_6395,N_6315);
and U8780 (N_8780,N_6676,N_6403);
and U8781 (N_8781,N_6763,N_6219);
or U8782 (N_8782,N_6039,N_6416);
nand U8783 (N_8783,N_6395,N_6816);
nand U8784 (N_8784,N_6859,N_6396);
or U8785 (N_8785,N_6225,N_6280);
or U8786 (N_8786,N_7010,N_6428);
nand U8787 (N_8787,N_7450,N_6491);
nand U8788 (N_8788,N_6775,N_7444);
or U8789 (N_8789,N_7410,N_7216);
nand U8790 (N_8790,N_6709,N_6073);
and U8791 (N_8791,N_6849,N_6034);
nor U8792 (N_8792,N_6123,N_6865);
nand U8793 (N_8793,N_7073,N_6174);
nand U8794 (N_8794,N_6032,N_7315);
or U8795 (N_8795,N_6205,N_7250);
and U8796 (N_8796,N_6209,N_6144);
or U8797 (N_8797,N_6723,N_6638);
or U8798 (N_8798,N_6316,N_7370);
or U8799 (N_8799,N_6709,N_7325);
nand U8800 (N_8800,N_6529,N_6517);
and U8801 (N_8801,N_6061,N_6991);
and U8802 (N_8802,N_6869,N_6933);
or U8803 (N_8803,N_6698,N_6296);
nand U8804 (N_8804,N_6554,N_6972);
or U8805 (N_8805,N_6505,N_6532);
nand U8806 (N_8806,N_6326,N_7033);
nor U8807 (N_8807,N_6780,N_6225);
or U8808 (N_8808,N_6572,N_6174);
and U8809 (N_8809,N_6269,N_6106);
xnor U8810 (N_8810,N_6191,N_6117);
and U8811 (N_8811,N_7123,N_6332);
nor U8812 (N_8812,N_7494,N_6859);
or U8813 (N_8813,N_6179,N_6823);
nand U8814 (N_8814,N_6674,N_6427);
nor U8815 (N_8815,N_6952,N_7325);
and U8816 (N_8816,N_6450,N_7148);
and U8817 (N_8817,N_6989,N_7354);
nor U8818 (N_8818,N_7068,N_7404);
or U8819 (N_8819,N_6358,N_6782);
or U8820 (N_8820,N_6164,N_6042);
and U8821 (N_8821,N_7303,N_7485);
or U8822 (N_8822,N_6123,N_6755);
or U8823 (N_8823,N_6767,N_6421);
nor U8824 (N_8824,N_6914,N_6881);
and U8825 (N_8825,N_6262,N_6481);
or U8826 (N_8826,N_6973,N_7286);
or U8827 (N_8827,N_7152,N_6929);
or U8828 (N_8828,N_6368,N_7459);
nor U8829 (N_8829,N_7269,N_7235);
or U8830 (N_8830,N_6849,N_6332);
nand U8831 (N_8831,N_7383,N_7151);
nand U8832 (N_8832,N_6638,N_6207);
or U8833 (N_8833,N_6865,N_6420);
or U8834 (N_8834,N_6541,N_6007);
or U8835 (N_8835,N_7207,N_6401);
and U8836 (N_8836,N_6097,N_6526);
and U8837 (N_8837,N_6516,N_6013);
or U8838 (N_8838,N_7448,N_6316);
xor U8839 (N_8839,N_7252,N_6372);
nand U8840 (N_8840,N_6442,N_6928);
xor U8841 (N_8841,N_7018,N_6572);
nand U8842 (N_8842,N_6760,N_6437);
nor U8843 (N_8843,N_7457,N_6707);
and U8844 (N_8844,N_7491,N_7253);
nand U8845 (N_8845,N_6074,N_6966);
or U8846 (N_8846,N_6826,N_6895);
and U8847 (N_8847,N_6198,N_7483);
and U8848 (N_8848,N_6252,N_6620);
nor U8849 (N_8849,N_6084,N_6643);
nor U8850 (N_8850,N_6377,N_6228);
nand U8851 (N_8851,N_6248,N_6201);
nand U8852 (N_8852,N_7284,N_6235);
nand U8853 (N_8853,N_6543,N_7307);
or U8854 (N_8854,N_6991,N_6437);
nand U8855 (N_8855,N_7270,N_7101);
and U8856 (N_8856,N_7207,N_7048);
nor U8857 (N_8857,N_6076,N_6608);
and U8858 (N_8858,N_6676,N_6439);
xnor U8859 (N_8859,N_6587,N_6347);
nand U8860 (N_8860,N_6794,N_6597);
nor U8861 (N_8861,N_6341,N_6262);
nand U8862 (N_8862,N_6250,N_6043);
nor U8863 (N_8863,N_6561,N_7101);
or U8864 (N_8864,N_6789,N_6354);
or U8865 (N_8865,N_6812,N_6279);
nor U8866 (N_8866,N_6096,N_6076);
nand U8867 (N_8867,N_7193,N_6014);
nand U8868 (N_8868,N_7354,N_7403);
and U8869 (N_8869,N_6953,N_6854);
nor U8870 (N_8870,N_6436,N_6227);
nor U8871 (N_8871,N_7166,N_6603);
nor U8872 (N_8872,N_6102,N_6598);
and U8873 (N_8873,N_6026,N_6564);
and U8874 (N_8874,N_6064,N_6222);
nor U8875 (N_8875,N_6378,N_6345);
nand U8876 (N_8876,N_7387,N_6906);
or U8877 (N_8877,N_6517,N_6659);
and U8878 (N_8878,N_7047,N_7141);
or U8879 (N_8879,N_7496,N_7224);
and U8880 (N_8880,N_6917,N_7410);
or U8881 (N_8881,N_6933,N_7149);
nor U8882 (N_8882,N_6226,N_7465);
nand U8883 (N_8883,N_6779,N_6709);
nor U8884 (N_8884,N_6467,N_7049);
and U8885 (N_8885,N_6944,N_6449);
nand U8886 (N_8886,N_6181,N_7233);
nor U8887 (N_8887,N_6311,N_7077);
or U8888 (N_8888,N_6953,N_6105);
and U8889 (N_8889,N_7315,N_7058);
nor U8890 (N_8890,N_6801,N_6420);
and U8891 (N_8891,N_6019,N_6073);
or U8892 (N_8892,N_7401,N_7407);
nand U8893 (N_8893,N_7033,N_6021);
or U8894 (N_8894,N_7100,N_6895);
and U8895 (N_8895,N_6231,N_6165);
nor U8896 (N_8896,N_6260,N_6278);
or U8897 (N_8897,N_7216,N_6981);
and U8898 (N_8898,N_6380,N_6765);
nand U8899 (N_8899,N_6341,N_6472);
nand U8900 (N_8900,N_7417,N_7246);
and U8901 (N_8901,N_6422,N_7420);
or U8902 (N_8902,N_6963,N_6985);
nor U8903 (N_8903,N_6904,N_6232);
and U8904 (N_8904,N_6428,N_7455);
or U8905 (N_8905,N_6763,N_6660);
or U8906 (N_8906,N_6109,N_6679);
nand U8907 (N_8907,N_6187,N_6926);
and U8908 (N_8908,N_7333,N_6951);
or U8909 (N_8909,N_6370,N_6216);
nand U8910 (N_8910,N_7005,N_6576);
nand U8911 (N_8911,N_6326,N_7129);
and U8912 (N_8912,N_6619,N_6544);
nor U8913 (N_8913,N_6812,N_7409);
or U8914 (N_8914,N_6985,N_7152);
and U8915 (N_8915,N_6112,N_7150);
and U8916 (N_8916,N_6008,N_6616);
or U8917 (N_8917,N_6548,N_6619);
nor U8918 (N_8918,N_6284,N_6153);
or U8919 (N_8919,N_6325,N_6132);
nand U8920 (N_8920,N_6621,N_6350);
nand U8921 (N_8921,N_6034,N_7193);
nor U8922 (N_8922,N_6874,N_6820);
and U8923 (N_8923,N_6558,N_6415);
or U8924 (N_8924,N_6523,N_6457);
and U8925 (N_8925,N_7420,N_6340);
nand U8926 (N_8926,N_6415,N_6629);
or U8927 (N_8927,N_6888,N_6213);
and U8928 (N_8928,N_7451,N_6973);
nor U8929 (N_8929,N_6711,N_6424);
nor U8930 (N_8930,N_7075,N_6233);
or U8931 (N_8931,N_7382,N_6641);
nand U8932 (N_8932,N_6540,N_6350);
nor U8933 (N_8933,N_6898,N_6860);
and U8934 (N_8934,N_6894,N_6656);
and U8935 (N_8935,N_6150,N_7389);
or U8936 (N_8936,N_6962,N_7322);
and U8937 (N_8937,N_7309,N_6133);
and U8938 (N_8938,N_7055,N_7416);
or U8939 (N_8939,N_6236,N_6201);
xnor U8940 (N_8940,N_7100,N_6184);
and U8941 (N_8941,N_6607,N_6831);
or U8942 (N_8942,N_6733,N_6110);
nand U8943 (N_8943,N_6641,N_7082);
and U8944 (N_8944,N_6543,N_6694);
nand U8945 (N_8945,N_7104,N_6699);
nand U8946 (N_8946,N_6842,N_7292);
and U8947 (N_8947,N_7109,N_6003);
nand U8948 (N_8948,N_6149,N_6633);
and U8949 (N_8949,N_7182,N_7492);
or U8950 (N_8950,N_6698,N_6726);
or U8951 (N_8951,N_6414,N_7042);
or U8952 (N_8952,N_6258,N_6841);
or U8953 (N_8953,N_6046,N_7052);
nor U8954 (N_8954,N_7090,N_6692);
and U8955 (N_8955,N_7050,N_6214);
nand U8956 (N_8956,N_7086,N_7326);
nand U8957 (N_8957,N_6776,N_6349);
or U8958 (N_8958,N_7018,N_6061);
nor U8959 (N_8959,N_6614,N_7151);
nand U8960 (N_8960,N_7125,N_6656);
xnor U8961 (N_8961,N_7014,N_6272);
nand U8962 (N_8962,N_6561,N_6892);
or U8963 (N_8963,N_6710,N_7433);
nor U8964 (N_8964,N_7221,N_6429);
or U8965 (N_8965,N_6065,N_6667);
xnor U8966 (N_8966,N_6366,N_6570);
or U8967 (N_8967,N_7361,N_6587);
nand U8968 (N_8968,N_7271,N_7195);
nand U8969 (N_8969,N_7221,N_6918);
and U8970 (N_8970,N_7155,N_7389);
and U8971 (N_8971,N_7389,N_6044);
nand U8972 (N_8972,N_6075,N_6723);
or U8973 (N_8973,N_6269,N_6210);
nand U8974 (N_8974,N_6680,N_6484);
or U8975 (N_8975,N_7439,N_7279);
nor U8976 (N_8976,N_6449,N_6041);
nor U8977 (N_8977,N_6280,N_6527);
or U8978 (N_8978,N_6589,N_6560);
nor U8979 (N_8979,N_6391,N_6794);
nor U8980 (N_8980,N_7315,N_7248);
nand U8981 (N_8981,N_7055,N_7155);
and U8982 (N_8982,N_6314,N_7317);
and U8983 (N_8983,N_7003,N_6436);
nor U8984 (N_8984,N_7137,N_6293);
nand U8985 (N_8985,N_7352,N_7435);
or U8986 (N_8986,N_6923,N_7444);
and U8987 (N_8987,N_6034,N_6215);
nand U8988 (N_8988,N_7031,N_6156);
nand U8989 (N_8989,N_6672,N_7284);
and U8990 (N_8990,N_6435,N_6239);
nand U8991 (N_8991,N_6127,N_6327);
nor U8992 (N_8992,N_6352,N_6488);
or U8993 (N_8993,N_6712,N_6170);
and U8994 (N_8994,N_7213,N_6145);
nand U8995 (N_8995,N_6311,N_7049);
and U8996 (N_8996,N_6500,N_6102);
or U8997 (N_8997,N_6651,N_6815);
nand U8998 (N_8998,N_6680,N_6215);
and U8999 (N_8999,N_6651,N_6099);
and U9000 (N_9000,N_8919,N_7902);
and U9001 (N_9001,N_8081,N_8292);
or U9002 (N_9002,N_8949,N_8504);
nor U9003 (N_9003,N_8363,N_8410);
or U9004 (N_9004,N_8475,N_8820);
or U9005 (N_9005,N_7757,N_7506);
nand U9006 (N_9006,N_7652,N_8026);
and U9007 (N_9007,N_8498,N_8585);
and U9008 (N_9008,N_7713,N_8831);
or U9009 (N_9009,N_8177,N_8441);
and U9010 (N_9010,N_8672,N_8552);
nand U9011 (N_9011,N_7643,N_7969);
and U9012 (N_9012,N_8968,N_8809);
or U9013 (N_9013,N_8909,N_8027);
nor U9014 (N_9014,N_7801,N_7951);
or U9015 (N_9015,N_8036,N_8301);
and U9016 (N_9016,N_8602,N_8342);
or U9017 (N_9017,N_7870,N_8562);
and U9018 (N_9018,N_7532,N_7554);
or U9019 (N_9019,N_8325,N_8954);
and U9020 (N_9020,N_7621,N_7936);
nor U9021 (N_9021,N_8059,N_7933);
or U9022 (N_9022,N_8680,N_8063);
or U9023 (N_9023,N_7804,N_7930);
or U9024 (N_9024,N_8135,N_7913);
and U9025 (N_9025,N_8308,N_7600);
nand U9026 (N_9026,N_8957,N_8638);
nand U9027 (N_9027,N_8367,N_7788);
and U9028 (N_9028,N_8061,N_7709);
nand U9029 (N_9029,N_8448,N_8594);
nor U9030 (N_9030,N_7723,N_7727);
nor U9031 (N_9031,N_8629,N_8024);
nand U9032 (N_9032,N_8510,N_7985);
nand U9033 (N_9033,N_8781,N_7567);
and U9034 (N_9034,N_8920,N_7648);
nor U9035 (N_9035,N_7928,N_8001);
and U9036 (N_9036,N_8845,N_8269);
nor U9037 (N_9037,N_8144,N_8256);
nor U9038 (N_9038,N_8775,N_8616);
or U9039 (N_9039,N_7903,N_8897);
and U9040 (N_9040,N_8155,N_7961);
nor U9041 (N_9041,N_8537,N_8017);
or U9042 (N_9042,N_8999,N_8422);
nor U9043 (N_9043,N_8089,N_8451);
nor U9044 (N_9044,N_8543,N_8095);
nand U9045 (N_9045,N_8685,N_8418);
and U9046 (N_9046,N_8521,N_7883);
nor U9047 (N_9047,N_8804,N_8335);
or U9048 (N_9048,N_7500,N_8033);
or U9049 (N_9049,N_8208,N_8090);
or U9050 (N_9050,N_8706,N_8791);
or U9051 (N_9051,N_7995,N_8720);
or U9052 (N_9052,N_7521,N_8705);
nand U9053 (N_9053,N_7968,N_8823);
or U9054 (N_9054,N_7908,N_8558);
and U9055 (N_9055,N_8861,N_8306);
and U9056 (N_9056,N_7917,N_8664);
and U9057 (N_9057,N_8221,N_7948);
nor U9058 (N_9058,N_8064,N_8575);
and U9059 (N_9059,N_8379,N_7695);
nor U9060 (N_9060,N_8153,N_8931);
nand U9061 (N_9061,N_7862,N_7983);
nor U9062 (N_9062,N_7871,N_7994);
or U9063 (N_9063,N_7920,N_7632);
or U9064 (N_9064,N_8803,N_8567);
and U9065 (N_9065,N_7647,N_8644);
nand U9066 (N_9066,N_8245,N_8557);
or U9067 (N_9067,N_7697,N_7748);
or U9068 (N_9068,N_8646,N_7982);
nand U9069 (N_9069,N_8146,N_7775);
and U9070 (N_9070,N_8390,N_8354);
and U9071 (N_9071,N_8692,N_7832);
nor U9072 (N_9072,N_7977,N_7842);
or U9073 (N_9073,N_7747,N_8573);
nor U9074 (N_9074,N_7984,N_7691);
nand U9075 (N_9075,N_8223,N_8197);
nand U9076 (N_9076,N_8226,N_8873);
nand U9077 (N_9077,N_7759,N_8201);
or U9078 (N_9078,N_7593,N_8322);
nor U9079 (N_9079,N_8773,N_8730);
and U9080 (N_9080,N_8601,N_8523);
and U9081 (N_9081,N_8946,N_7702);
or U9082 (N_9082,N_8419,N_7729);
nand U9083 (N_9083,N_8735,N_8625);
nor U9084 (N_9084,N_8468,N_8477);
or U9085 (N_9085,N_7992,N_8595);
and U9086 (N_9086,N_8598,N_7745);
nand U9087 (N_9087,N_8959,N_7724);
and U9088 (N_9088,N_8290,N_7909);
nand U9089 (N_9089,N_8799,N_8670);
nand U9090 (N_9090,N_7603,N_7504);
nor U9091 (N_9091,N_8219,N_8532);
nor U9092 (N_9092,N_7566,N_7740);
or U9093 (N_9093,N_7588,N_7805);
nor U9094 (N_9094,N_8753,N_7750);
nor U9095 (N_9095,N_8125,N_8711);
nand U9096 (N_9096,N_7831,N_7587);
and U9097 (N_9097,N_8472,N_8016);
nor U9098 (N_9098,N_8827,N_8164);
nand U9099 (N_9099,N_7770,N_8715);
nor U9100 (N_9100,N_8307,N_8784);
and U9101 (N_9101,N_8224,N_8912);
or U9102 (N_9102,N_7630,N_7837);
and U9103 (N_9103,N_8856,N_7570);
and U9104 (N_9104,N_8875,N_7548);
or U9105 (N_9105,N_8811,N_7639);
or U9106 (N_9106,N_7999,N_8466);
nor U9107 (N_9107,N_7591,N_8790);
nor U9108 (N_9108,N_8172,N_7514);
and U9109 (N_9109,N_7797,N_7853);
nor U9110 (N_9110,N_7998,N_7865);
xor U9111 (N_9111,N_8134,N_7658);
nor U9112 (N_9112,N_8070,N_7615);
and U9113 (N_9113,N_7791,N_8123);
and U9114 (N_9114,N_7949,N_8106);
nand U9115 (N_9115,N_7519,N_8194);
or U9116 (N_9116,N_7612,N_7843);
nand U9117 (N_9117,N_7828,N_8128);
or U9118 (N_9118,N_8599,N_8238);
and U9119 (N_9119,N_8490,N_8348);
or U9120 (N_9120,N_8055,N_8826);
and U9121 (N_9121,N_8566,N_7705);
and U9122 (N_9122,N_8005,N_8182);
and U9123 (N_9123,N_8788,N_8321);
and U9124 (N_9124,N_7778,N_8295);
and U9125 (N_9125,N_8420,N_8358);
xor U9126 (N_9126,N_7619,N_8141);
nor U9127 (N_9127,N_7662,N_7905);
nand U9128 (N_9128,N_8161,N_7677);
or U9129 (N_9129,N_8339,N_8406);
and U9130 (N_9130,N_7594,N_7597);
or U9131 (N_9131,N_8641,N_8188);
or U9132 (N_9132,N_8841,N_8700);
or U9133 (N_9133,N_8288,N_7776);
nand U9134 (N_9134,N_8760,N_8916);
nand U9135 (N_9135,N_8396,N_7611);
or U9136 (N_9136,N_8818,N_7613);
or U9137 (N_9137,N_8789,N_7501);
or U9138 (N_9138,N_8000,N_7675);
or U9139 (N_9139,N_8277,N_7889);
or U9140 (N_9140,N_8872,N_8242);
nor U9141 (N_9141,N_7937,N_8654);
and U9142 (N_9142,N_7857,N_7838);
nor U9143 (N_9143,N_8832,N_8010);
nor U9144 (N_9144,N_8344,N_8671);
and U9145 (N_9145,N_7980,N_8075);
nor U9146 (N_9146,N_8854,N_7940);
xnor U9147 (N_9147,N_8052,N_7833);
nor U9148 (N_9148,N_8004,N_8699);
nor U9149 (N_9149,N_8237,N_8278);
or U9150 (N_9150,N_8539,N_8205);
nor U9151 (N_9151,N_7608,N_8855);
nor U9152 (N_9152,N_8553,N_8503);
and U9153 (N_9153,N_8446,N_8732);
nor U9154 (N_9154,N_8836,N_7565);
nor U9155 (N_9155,N_8716,N_8285);
nor U9156 (N_9156,N_8935,N_7574);
or U9157 (N_9157,N_7581,N_8035);
xor U9158 (N_9158,N_8282,N_8323);
or U9159 (N_9159,N_8907,N_8497);
or U9160 (N_9160,N_7773,N_8513);
nand U9161 (N_9161,N_8564,N_8812);
and U9162 (N_9162,N_8158,N_7605);
nand U9163 (N_9163,N_8686,N_7672);
nand U9164 (N_9164,N_8351,N_8357);
nand U9165 (N_9165,N_7529,N_7784);
nand U9166 (N_9166,N_7645,N_7845);
nand U9167 (N_9167,N_8244,N_8857);
and U9168 (N_9168,N_8372,N_8434);
or U9169 (N_9169,N_7888,N_8012);
nor U9170 (N_9170,N_8359,N_8154);
and U9171 (N_9171,N_8586,N_8159);
and U9172 (N_9172,N_8560,N_8987);
nand U9173 (N_9173,N_7993,N_8657);
nand U9174 (N_9174,N_8369,N_8364);
nor U9175 (N_9175,N_7796,N_8973);
or U9176 (N_9176,N_8209,N_8460);
and U9177 (N_9177,N_7543,N_8427);
and U9178 (N_9178,N_7683,N_7991);
nand U9179 (N_9179,N_8948,N_8750);
nand U9180 (N_9180,N_8019,N_8776);
nand U9181 (N_9181,N_8243,N_8408);
nor U9182 (N_9182,N_8737,N_7953);
nand U9183 (N_9183,N_8709,N_7684);
nand U9184 (N_9184,N_8330,N_8633);
nor U9185 (N_9185,N_7935,N_8584);
nor U9186 (N_9186,N_8681,N_8688);
nor U9187 (N_9187,N_7946,N_7622);
xnor U9188 (N_9188,N_8313,N_8212);
nor U9189 (N_9189,N_8530,N_7822);
and U9190 (N_9190,N_8527,N_8926);
and U9191 (N_9191,N_8696,N_7872);
and U9192 (N_9192,N_8758,N_8337);
nor U9193 (N_9193,N_7690,N_8470);
nor U9194 (N_9194,N_8943,N_8506);
nor U9195 (N_9195,N_8956,N_8051);
or U9196 (N_9196,N_7899,N_7829);
nand U9197 (N_9197,N_8701,N_8763);
nand U9198 (N_9198,N_7896,N_8590);
nand U9199 (N_9199,N_8800,N_8077);
or U9200 (N_9200,N_7628,N_7559);
nand U9201 (N_9201,N_8392,N_8755);
and U9202 (N_9202,N_8119,N_8381);
nand U9203 (N_9203,N_8045,N_8921);
or U9204 (N_9204,N_7868,N_7636);
or U9205 (N_9205,N_8041,N_8667);
nor U9206 (N_9206,N_8507,N_8961);
nand U9207 (N_9207,N_7809,N_8281);
or U9208 (N_9208,N_8828,N_7879);
and U9209 (N_9209,N_8574,N_8984);
nand U9210 (N_9210,N_8072,N_8170);
nand U9211 (N_9211,N_8496,N_8195);
nand U9212 (N_9212,N_7542,N_8186);
and U9213 (N_9213,N_8710,N_7954);
nand U9214 (N_9214,N_8632,N_8879);
and U9215 (N_9215,N_7975,N_8576);
nand U9216 (N_9216,N_7586,N_8794);
nand U9217 (N_9217,N_8399,N_8104);
nand U9218 (N_9218,N_8196,N_8871);
nor U9219 (N_9219,N_8156,N_8908);
or U9220 (N_9220,N_7766,N_8938);
and U9221 (N_9221,N_8866,N_8998);
xor U9222 (N_9222,N_7765,N_8502);
nand U9223 (N_9223,N_8349,N_7959);
nor U9224 (N_9224,N_8044,N_8228);
or U9225 (N_9225,N_8362,N_7812);
and U9226 (N_9226,N_8734,N_8631);
nor U9227 (N_9227,N_7701,N_7517);
nand U9228 (N_9228,N_8884,N_7717);
and U9229 (N_9229,N_8165,N_8694);
or U9230 (N_9230,N_7692,N_7551);
and U9231 (N_9231,N_8937,N_8137);
nor U9232 (N_9232,N_7798,N_7512);
nor U9233 (N_9233,N_8407,N_8189);
xnor U9234 (N_9234,N_7877,N_7525);
nand U9235 (N_9235,N_8317,N_7582);
or U9236 (N_9236,N_8492,N_8605);
and U9237 (N_9237,N_7781,N_8600);
or U9238 (N_9238,N_8930,N_7725);
and U9239 (N_9239,N_8541,N_8554);
or U9240 (N_9240,N_8689,N_8102);
nor U9241 (N_9241,N_7965,N_8176);
nor U9242 (N_9242,N_8084,N_8565);
nor U9243 (N_9243,N_8439,N_8080);
nand U9244 (N_9244,N_8082,N_8747);
or U9245 (N_9245,N_8993,N_8428);
nor U9246 (N_9246,N_8785,N_8368);
nand U9247 (N_9247,N_8536,N_7824);
nand U9248 (N_9248,N_8405,N_8953);
nor U9249 (N_9249,N_7650,N_8087);
and U9250 (N_9250,N_8848,N_8393);
or U9251 (N_9251,N_8813,N_8996);
nand U9252 (N_9252,N_8893,N_7642);
and U9253 (N_9253,N_8662,N_8661);
nor U9254 (N_9254,N_8780,N_8914);
and U9255 (N_9255,N_7919,N_8199);
nor U9256 (N_9256,N_7669,N_8065);
or U9257 (N_9257,N_8302,N_7817);
or U9258 (N_9258,N_8656,N_8712);
and U9259 (N_9259,N_8340,N_8976);
or U9260 (N_9260,N_8904,N_8822);
nor U9261 (N_9261,N_8819,N_8969);
and U9262 (N_9262,N_8821,N_8870);
nor U9263 (N_9263,N_8883,N_7922);
nor U9264 (N_9264,N_7846,N_7694);
and U9265 (N_9265,N_8037,N_7735);
or U9266 (N_9266,N_8910,N_8459);
nor U9267 (N_9267,N_8495,N_8548);
and U9268 (N_9268,N_7810,N_8022);
and U9269 (N_9269,N_8771,N_8531);
nand U9270 (N_9270,N_8814,N_8890);
or U9271 (N_9271,N_8842,N_8116);
or U9272 (N_9272,N_7947,N_8708);
or U9273 (N_9273,N_8388,N_7979);
nand U9274 (N_9274,N_8118,N_7821);
nor U9275 (N_9275,N_8555,N_8733);
and U9276 (N_9276,N_8371,N_8450);
and U9277 (N_9277,N_8778,N_8626);
nand U9278 (N_9278,N_8549,N_8556);
nor U9279 (N_9279,N_8484,N_7743);
nor U9280 (N_9280,N_8929,N_7808);
and U9281 (N_9281,N_8642,N_8550);
nand U9282 (N_9282,N_7732,N_8499);
nor U9283 (N_9283,N_8387,N_8328);
or U9284 (N_9284,N_7840,N_8166);
nand U9285 (N_9285,N_7646,N_8596);
or U9286 (N_9286,N_8860,N_8918);
and U9287 (N_9287,N_8142,N_8140);
or U9288 (N_9288,N_8666,N_7714);
or U9289 (N_9289,N_8143,N_8751);
nand U9290 (N_9290,N_8713,N_8018);
nor U9291 (N_9291,N_8382,N_8587);
nor U9292 (N_9292,N_8426,N_8375);
nand U9293 (N_9293,N_8997,N_7874);
nor U9294 (N_9294,N_8906,N_8787);
nor U9295 (N_9295,N_8376,N_8270);
or U9296 (N_9296,N_8391,N_7912);
or U9297 (N_9297,N_8683,N_8417);
and U9298 (N_9298,N_8132,N_8263);
xor U9299 (N_9299,N_8425,N_8105);
nand U9300 (N_9300,N_7848,N_8336);
nor U9301 (N_9301,N_8147,N_8621);
or U9302 (N_9302,N_7689,N_8698);
nor U9303 (N_9303,N_8529,N_8480);
nand U9304 (N_9304,N_8259,N_8752);
nor U9305 (N_9305,N_8677,N_8623);
nor U9306 (N_9306,N_7737,N_8056);
or U9307 (N_9307,N_7927,N_8284);
and U9308 (N_9308,N_8046,N_7986);
nand U9309 (N_9309,N_8464,N_8829);
and U9310 (N_9310,N_8062,N_8442);
or U9311 (N_9311,N_8885,N_8346);
or U9312 (N_9312,N_8639,N_8649);
or U9313 (N_9313,N_8637,N_7536);
nand U9314 (N_9314,N_8054,N_8014);
or U9315 (N_9315,N_8453,N_8286);
and U9316 (N_9316,N_8404,N_8798);
nand U9317 (N_9317,N_8665,N_8673);
nand U9318 (N_9318,N_7719,N_8786);
and U9319 (N_9319,N_8617,N_8707);
or U9320 (N_9320,N_8192,N_7564);
or U9321 (N_9321,N_8247,N_8184);
nor U9322 (N_9322,N_7556,N_8612);
nand U9323 (N_9323,N_7507,N_7753);
and U9324 (N_9324,N_8965,N_8169);
and U9325 (N_9325,N_8519,N_7782);
or U9326 (N_9326,N_8635,N_8876);
or U9327 (N_9327,N_7878,N_7509);
nor U9328 (N_9328,N_8473,N_7544);
or U9329 (N_9329,N_8374,N_8079);
nor U9330 (N_9330,N_7641,N_7774);
or U9331 (N_9331,N_8311,N_8461);
nand U9332 (N_9332,N_8679,N_8850);
or U9333 (N_9333,N_7561,N_7609);
and U9334 (N_9334,N_7718,N_8078);
and U9335 (N_9335,N_7602,N_7898);
and U9336 (N_9336,N_8456,N_7901);
nand U9337 (N_9337,N_8721,N_7962);
and U9338 (N_9338,N_8091,N_8613);
or U9339 (N_9339,N_8913,N_8267);
nand U9340 (N_9340,N_8048,N_8465);
or U9341 (N_9341,N_8108,N_8312);
and U9342 (N_9342,N_7681,N_8589);
nand U9343 (N_9343,N_8611,N_7785);
nor U9344 (N_9344,N_8924,N_7635);
nor U9345 (N_9345,N_7686,N_8726);
nor U9346 (N_9346,N_8252,N_8928);
or U9347 (N_9347,N_8991,N_8167);
nand U9348 (N_9348,N_7967,N_7864);
nor U9349 (N_9349,N_7955,N_8347);
and U9350 (N_9350,N_8314,N_8260);
or U9351 (N_9351,N_7764,N_8103);
nand U9352 (N_9352,N_8958,N_8859);
nand U9353 (N_9353,N_8604,N_8867);
or U9354 (N_9354,N_7925,N_8887);
nand U9355 (N_9355,N_8049,N_7726);
or U9356 (N_9356,N_8863,N_8443);
or U9357 (N_9357,N_7661,N_7720);
nor U9358 (N_9358,N_7617,N_7550);
nand U9359 (N_9359,N_7712,N_8849);
or U9360 (N_9360,N_8772,N_8741);
or U9361 (N_9361,N_8902,N_8462);
or U9362 (N_9362,N_8889,N_8236);
or U9363 (N_9363,N_8522,N_7976);
nor U9364 (N_9364,N_7891,N_7513);
nor U9365 (N_9365,N_8331,N_7510);
or U9366 (N_9366,N_8500,N_7873);
nand U9367 (N_9367,N_7783,N_8258);
nand U9368 (N_9368,N_8482,N_8289);
nand U9369 (N_9369,N_7671,N_8253);
xnor U9370 (N_9370,N_8006,N_7706);
nand U9371 (N_9371,N_8757,N_8501);
and U9372 (N_9372,N_8148,N_8467);
or U9373 (N_9373,N_7769,N_7606);
nor U9374 (N_9374,N_8927,N_7807);
nand U9375 (N_9375,N_8400,N_8768);
nor U9376 (N_9376,N_8844,N_8168);
or U9377 (N_9377,N_8742,N_7533);
nor U9378 (N_9378,N_8945,N_7547);
and U9379 (N_9379,N_7942,N_8511);
and U9380 (N_9380,N_8233,N_8719);
nor U9381 (N_9381,N_8676,N_8865);
nand U9382 (N_9382,N_7523,N_8942);
or U9383 (N_9383,N_8008,N_7861);
nor U9384 (N_9384,N_8653,N_8774);
nand U9385 (N_9385,N_8098,N_7827);
and U9386 (N_9386,N_7580,N_8248);
nand U9387 (N_9387,N_8932,N_8559);
nor U9388 (N_9388,N_8583,N_8761);
nor U9389 (N_9389,N_7858,N_8606);
nor U9390 (N_9390,N_8964,N_8038);
or U9391 (N_9391,N_8432,N_8533);
or U9392 (N_9392,N_7815,N_8833);
nand U9393 (N_9393,N_7813,N_8995);
and U9394 (N_9394,N_7849,N_8933);
and U9395 (N_9395,N_7644,N_8545);
and U9396 (N_9396,N_8512,N_8538);
or U9397 (N_9397,N_7830,N_7987);
nor U9398 (N_9398,N_7590,N_7884);
xnor U9399 (N_9399,N_8293,N_7502);
or U9400 (N_9400,N_8092,N_8915);
nor U9401 (N_9401,N_8327,N_8149);
nand U9402 (N_9402,N_8609,N_8454);
nand U9403 (N_9403,N_8725,N_8319);
and U9404 (N_9404,N_8028,N_8463);
and U9405 (N_9405,N_8231,N_8178);
nor U9406 (N_9406,N_8415,N_8950);
and U9407 (N_9407,N_8250,N_8268);
or U9408 (N_9408,N_7583,N_8972);
nor U9409 (N_9409,N_7989,N_8329);
nand U9410 (N_9410,N_8767,N_7880);
nor U9411 (N_9411,N_8514,N_8660);
and U9412 (N_9412,N_8074,N_8951);
or U9413 (N_9413,N_7971,N_7618);
and U9414 (N_9414,N_8191,N_7850);
nor U9415 (N_9415,N_8645,N_7741);
xnor U9416 (N_9416,N_8569,N_7614);
nand U9417 (N_9417,N_8175,N_7730);
and U9418 (N_9418,N_7860,N_8630);
and U9419 (N_9419,N_8690,N_8544);
and U9420 (N_9420,N_8944,N_7631);
nor U9421 (N_9421,N_7746,N_7904);
nand U9422 (N_9422,N_7792,N_8094);
and U9423 (N_9423,N_8678,N_7956);
nor U9424 (N_9424,N_8494,N_8207);
and U9425 (N_9425,N_8764,N_7793);
nor U9426 (N_9426,N_7634,N_8251);
nand U9427 (N_9427,N_8684,N_8988);
nor U9428 (N_9428,N_7761,N_8249);
and U9429 (N_9429,N_8911,N_8232);
and U9430 (N_9430,N_8736,N_8160);
nand U9431 (N_9431,N_8262,N_7907);
nor U9432 (N_9432,N_7760,N_8067);
nor U9433 (N_9433,N_8941,N_8838);
or U9434 (N_9434,N_8843,N_7515);
nor U9435 (N_9435,N_7772,N_8650);
nand U9436 (N_9436,N_8580,N_8840);
nor U9437 (N_9437,N_8085,N_7640);
nand U9438 (N_9438,N_7762,N_7978);
nor U9439 (N_9439,N_8607,N_8122);
nor U9440 (N_9440,N_8326,N_7893);
nor U9441 (N_9441,N_7676,N_8517);
or U9442 (N_9442,N_7520,N_7545);
nor U9443 (N_9443,N_7572,N_8411);
xnor U9444 (N_9444,N_8881,N_7596);
nor U9445 (N_9445,N_8577,N_8994);
and U9446 (N_9446,N_8754,N_7699);
nand U9447 (N_9447,N_8117,N_8015);
and U9448 (N_9448,N_7707,N_7887);
nor U9449 (N_9449,N_8275,N_8975);
or U9450 (N_9450,N_7876,N_7767);
and U9451 (N_9451,N_8271,N_7819);
nand U9452 (N_9452,N_8806,N_7667);
nor U9453 (N_9453,N_8303,N_8296);
and U9454 (N_9454,N_7897,N_7654);
or U9455 (N_9455,N_8985,N_8796);
xnor U9456 (N_9456,N_7685,N_8624);
and U9457 (N_9457,N_8888,N_8588);
nor U9458 (N_9458,N_7972,N_7633);
nor U9459 (N_9459,N_8515,N_8663);
nor U9460 (N_9460,N_7670,N_8341);
nor U9461 (N_9461,N_8316,N_8412);
and U9462 (N_9462,N_7926,N_7522);
xnor U9463 (N_9463,N_7818,N_8745);
or U9464 (N_9464,N_8489,N_7546);
nor U9465 (N_9465,N_8974,N_7918);
or U9466 (N_9466,N_8546,N_8220);
or U9467 (N_9467,N_8193,N_8516);
nor U9468 (N_9468,N_7906,N_8213);
and U9469 (N_9469,N_7673,N_8272);
nor U9470 (N_9470,N_8797,N_8053);
and U9471 (N_9471,N_8343,N_8651);
nor U9472 (N_9472,N_8210,N_7779);
and U9473 (N_9473,N_7915,N_8218);
or U9474 (N_9474,N_8839,N_8234);
nand U9475 (N_9475,N_7931,N_8488);
and U9476 (N_9476,N_7733,N_8825);
or U9477 (N_9477,N_8636,N_8471);
or U9478 (N_9478,N_8648,N_7771);
nor U9479 (N_9479,N_8628,N_8978);
nand U9480 (N_9480,N_7924,N_8977);
and U9481 (N_9481,N_7704,N_8421);
and U9482 (N_9482,N_7716,N_7851);
nand U9483 (N_9483,N_8486,N_7708);
or U9484 (N_9484,N_7952,N_8695);
nor U9485 (N_9485,N_8744,N_8955);
or U9486 (N_9486,N_8332,N_8276);
nand U9487 (N_9487,N_8687,N_7911);
and U9488 (N_9488,N_7749,N_8380);
nand U9489 (N_9489,N_7811,N_8891);
nand U9490 (N_9490,N_8824,N_7964);
nor U9491 (N_9491,N_7763,N_8206);
nor U9492 (N_9492,N_8099,N_8150);
nand U9493 (N_9493,N_8762,N_8060);
nor U9494 (N_9494,N_7816,N_8174);
nand U9495 (N_9495,N_7526,N_8805);
or U9496 (N_9496,N_8291,N_8877);
and U9497 (N_9497,N_8801,N_7659);
nand U9498 (N_9498,N_8703,N_7799);
nor U9499 (N_9499,N_8042,N_8578);
nor U9500 (N_9500,N_8614,N_8299);
nor U9501 (N_9501,N_7541,N_8403);
nor U9502 (N_9502,N_8173,N_7698);
or U9503 (N_9503,N_8592,N_8971);
or U9504 (N_9504,N_7534,N_8452);
and U9505 (N_9505,N_8409,N_7703);
nor U9506 (N_9506,N_7835,N_7620);
or U9507 (N_9507,N_8043,N_7950);
and U9508 (N_9508,N_8963,N_8066);
and U9509 (N_9509,N_7668,N_8402);
nor U9510 (N_9510,N_8743,N_7910);
nor U9511 (N_9511,N_8862,N_8273);
nor U9512 (N_9512,N_8069,N_7595);
and U9513 (N_9513,N_8793,N_8257);
and U9514 (N_9514,N_7895,N_7900);
nand U9515 (N_9515,N_8023,N_8179);
nor U9516 (N_9516,N_7834,N_8593);
nor U9517 (N_9517,N_7859,N_7592);
nor U9518 (N_9518,N_7638,N_8350);
and U9519 (N_9519,N_7794,N_7656);
or U9520 (N_9520,N_8917,N_7516);
nand U9521 (N_9521,N_7790,N_7738);
nor U9522 (N_9522,N_8746,N_8294);
or U9523 (N_9523,N_8163,N_7627);
nand U9524 (N_9524,N_8225,N_8280);
nand U9525 (N_9525,N_8647,N_8430);
and U9526 (N_9526,N_8183,N_8040);
nand U9527 (N_9527,N_8385,N_7552);
and U9528 (N_9528,N_7786,N_8520);
nand U9529 (N_9529,N_8187,N_8769);
nand U9530 (N_9530,N_8966,N_8373);
and U9531 (N_9531,N_8315,N_8892);
nor U9532 (N_9532,N_8096,N_7731);
nand U9533 (N_9533,N_8485,N_8962);
or U9534 (N_9534,N_8795,N_8655);
or U9535 (N_9535,N_8384,N_8619);
or U9536 (N_9536,N_8551,N_7966);
and U9537 (N_9537,N_8967,N_8455);
nand U9538 (N_9538,N_8127,N_7752);
nor U9539 (N_9539,N_8133,N_7736);
and U9540 (N_9540,N_8071,N_8704);
or U9541 (N_9541,N_8652,N_8643);
or U9542 (N_9542,N_8923,N_7939);
nand U9543 (N_9543,N_8216,N_8992);
or U9544 (N_9544,N_7693,N_8847);
nor U9545 (N_9545,N_8230,N_8185);
nor U9546 (N_9546,N_8834,N_7990);
nor U9547 (N_9547,N_8353,N_8723);
nor U9548 (N_9548,N_8124,N_7687);
nor U9549 (N_9549,N_7528,N_7663);
and U9550 (N_9550,N_8525,N_8429);
nor U9551 (N_9551,N_8886,N_7844);
nor U9552 (N_9552,N_7974,N_7610);
or U9553 (N_9553,N_7624,N_8007);
or U9554 (N_9554,N_8318,N_8121);
and U9555 (N_9555,N_7530,N_8765);
and U9556 (N_9556,N_8002,N_7996);
and U9557 (N_9557,N_8131,N_8030);
nor U9558 (N_9558,N_8365,N_7531);
nand U9559 (N_9559,N_8748,N_7885);
nor U9560 (N_9560,N_8395,N_8782);
or U9561 (N_9561,N_7538,N_8939);
nor U9562 (N_9562,N_8438,N_8481);
nor U9563 (N_9563,N_7875,N_8579);
nor U9564 (N_9564,N_7963,N_7734);
and U9565 (N_9565,N_8640,N_8940);
xor U9566 (N_9566,N_8980,N_7696);
nand U9567 (N_9567,N_8922,N_8487);
nor U9568 (N_9568,N_8298,N_8246);
or U9569 (N_9569,N_8868,N_7820);
nand U9570 (N_9570,N_8815,N_7728);
nor U9571 (N_9571,N_8440,N_7585);
or U9572 (N_9572,N_8279,N_8334);
and U9573 (N_9573,N_8130,N_8093);
nand U9574 (N_9574,N_7678,N_7576);
nor U9575 (N_9575,N_8970,N_8202);
nand U9576 (N_9576,N_7960,N_7881);
nor U9577 (N_9577,N_8524,N_8668);
nand U9578 (N_9578,N_8618,N_7768);
nand U9579 (N_9579,N_8397,N_8853);
nor U9580 (N_9580,N_8240,N_8627);
or U9581 (N_9581,N_8200,N_7589);
nand U9582 (N_9582,N_8483,N_8100);
and U9583 (N_9583,N_8802,N_7802);
nor U9584 (N_9584,N_7780,N_8416);
nor U9585 (N_9585,N_7680,N_7916);
nand U9586 (N_9586,N_8215,N_7777);
or U9587 (N_9587,N_7869,N_7505);
and U9588 (N_9588,N_7679,N_7890);
and U9589 (N_9589,N_8034,N_8882);
and U9590 (N_9590,N_8983,N_7944);
nand U9591 (N_9591,N_7665,N_8895);
or U9592 (N_9592,N_8718,N_8903);
or U9593 (N_9593,N_8032,N_7660);
and U9594 (N_9594,N_8851,N_8505);
and U9595 (N_9595,N_7649,N_7806);
or U9596 (N_9596,N_8355,N_8021);
nand U9597 (N_9597,N_8029,N_7508);
nor U9598 (N_9598,N_7839,N_7674);
nor U9599 (N_9599,N_8101,N_8157);
and U9600 (N_9600,N_7756,N_7549);
nand U9601 (N_9601,N_7932,N_7655);
or U9602 (N_9602,N_8360,N_7863);
or U9603 (N_9603,N_7558,N_8180);
nor U9604 (N_9604,N_8352,N_8571);
nor U9605 (N_9605,N_8729,N_8749);
and U9606 (N_9606,N_8020,N_8361);
nand U9607 (N_9607,N_7710,N_8568);
nor U9608 (N_9608,N_7599,N_7943);
nand U9609 (N_9609,N_8310,N_7664);
or U9610 (N_9610,N_7742,N_7892);
or U9611 (N_9611,N_7721,N_8986);
or U9612 (N_9612,N_8437,N_8126);
or U9613 (N_9613,N_8287,N_8846);
or U9614 (N_9614,N_8047,N_8107);
nor U9615 (N_9615,N_8255,N_8582);
or U9616 (N_9616,N_7836,N_8345);
and U9617 (N_9617,N_7823,N_8110);
and U9618 (N_9618,N_7569,N_7518);
or U9619 (N_9619,N_7934,N_7929);
or U9620 (N_9620,N_7527,N_7789);
and U9621 (N_9621,N_8982,N_7571);
nor U9622 (N_9622,N_8659,N_8979);
or U9623 (N_9623,N_7787,N_8386);
or U9624 (N_9624,N_8563,N_8476);
and U9625 (N_9625,N_7629,N_8254);
or U9626 (N_9626,N_8581,N_8398);
nor U9627 (N_9627,N_7795,N_8899);
and U9628 (N_9628,N_7938,N_7607);
nor U9629 (N_9629,N_8900,N_8003);
nor U9630 (N_9630,N_7945,N_8370);
nor U9631 (N_9631,N_8171,N_8111);
or U9632 (N_9632,N_7553,N_7653);
nand U9633 (N_9633,N_7511,N_7997);
and U9634 (N_9634,N_7882,N_7625);
and U9635 (N_9635,N_8073,N_8058);
nor U9636 (N_9636,N_7657,N_8697);
nand U9637 (N_9637,N_8324,N_8265);
and U9638 (N_9638,N_8431,N_8894);
and U9639 (N_9639,N_7970,N_7856);
nor U9640 (N_9640,N_8011,N_8777);
or U9641 (N_9641,N_8309,N_8542);
nand U9642 (N_9642,N_8724,N_8508);
or U9643 (N_9643,N_7847,N_7623);
or U9644 (N_9644,N_8086,N_8057);
and U9645 (N_9645,N_8305,N_8905);
and U9646 (N_9646,N_8989,N_8925);
and U9647 (N_9647,N_8414,N_8603);
nand U9648 (N_9648,N_8413,N_8835);
nand U9649 (N_9649,N_8615,N_7537);
nor U9650 (N_9650,N_7535,N_8947);
or U9651 (N_9651,N_8837,N_8674);
and U9652 (N_9652,N_7688,N_8478);
nand U9653 (N_9653,N_8852,N_8394);
or U9654 (N_9654,N_8151,N_8990);
nor U9655 (N_9655,N_7981,N_8658);
or U9656 (N_9656,N_8901,N_7560);
and U9657 (N_9657,N_7800,N_8702);
or U9658 (N_9658,N_8766,N_7957);
and U9659 (N_9659,N_8457,N_8112);
nor U9660 (N_9660,N_8547,N_8088);
nor U9661 (N_9661,N_7826,N_8675);
or U9662 (N_9662,N_8114,N_7867);
or U9663 (N_9663,N_8528,N_8669);
nand U9664 (N_9664,N_8436,N_8136);
nor U9665 (N_9665,N_8435,N_7744);
and U9666 (N_9666,N_8145,N_8981);
nand U9667 (N_9667,N_8540,N_7575);
and U9668 (N_9668,N_8138,N_8229);
and U9669 (N_9669,N_8241,N_7557);
and U9670 (N_9670,N_7988,N_8050);
or U9671 (N_9671,N_7715,N_8682);
and U9672 (N_9672,N_8068,N_7524);
and U9673 (N_9673,N_8792,N_8759);
or U9674 (N_9674,N_8740,N_8731);
nand U9675 (N_9675,N_8783,N_7852);
and U9676 (N_9676,N_8491,N_7637);
nor U9677 (N_9677,N_8526,N_8083);
or U9678 (N_9678,N_8591,N_8934);
or U9679 (N_9679,N_7722,N_8190);
nor U9680 (N_9680,N_8227,N_8808);
nand U9681 (N_9681,N_8266,N_8333);
or U9682 (N_9682,N_8445,N_7555);
nand U9683 (N_9683,N_8109,N_8816);
nor U9684 (N_9684,N_8261,N_8297);
or U9685 (N_9685,N_8817,N_8444);
and U9686 (N_9686,N_8493,N_7973);
nand U9687 (N_9687,N_8874,N_8727);
nor U9688 (N_9688,N_7814,N_7579);
or U9689 (N_9689,N_7626,N_7562);
nor U9690 (N_9690,N_7854,N_8561);
or U9691 (N_9691,N_8152,N_7651);
nand U9692 (N_9692,N_8756,N_8389);
and U9693 (N_9693,N_7584,N_8960);
and U9694 (N_9694,N_8509,N_8217);
nor U9695 (N_9695,N_8458,N_8535);
nand U9696 (N_9696,N_8728,N_8356);
nor U9697 (N_9697,N_8097,N_7803);
or U9698 (N_9698,N_8810,N_8869);
and U9699 (N_9699,N_8770,N_8572);
and U9700 (N_9700,N_8211,N_8479);
or U9701 (N_9701,N_7941,N_7503);
nor U9702 (N_9702,N_7923,N_8691);
nor U9703 (N_9703,N_8377,N_8722);
or U9704 (N_9704,N_7539,N_8693);
xnor U9705 (N_9705,N_8214,N_8235);
nand U9706 (N_9706,N_7886,N_8013);
nor U9707 (N_9707,N_7758,N_8113);
nor U9708 (N_9708,N_8779,N_7739);
nor U9709 (N_9709,N_7894,N_8858);
or U9710 (N_9710,N_8378,N_8283);
nor U9711 (N_9711,N_7568,N_8120);
nor U9712 (N_9712,N_8115,N_7573);
nand U9713 (N_9713,N_8383,N_8264);
or U9714 (N_9714,N_8896,N_8039);
nor U9715 (N_9715,N_8222,N_8423);
nand U9716 (N_9716,N_8518,N_7700);
nand U9717 (N_9717,N_8807,N_8129);
xor U9718 (N_9718,N_8424,N_8622);
or U9719 (N_9719,N_8300,N_7866);
and U9720 (N_9720,N_8717,N_8447);
or U9721 (N_9721,N_8366,N_8864);
or U9722 (N_9722,N_7666,N_8620);
or U9723 (N_9723,N_7754,N_8449);
and U9724 (N_9724,N_8534,N_8597);
nand U9725 (N_9725,N_8570,N_7577);
nand U9726 (N_9726,N_8181,N_7921);
or U9727 (N_9727,N_7958,N_7604);
nand U9728 (N_9728,N_8076,N_8880);
and U9729 (N_9729,N_7616,N_8936);
nor U9730 (N_9730,N_7751,N_8203);
and U9731 (N_9731,N_8009,N_7578);
and U9732 (N_9732,N_8198,N_8610);
or U9733 (N_9733,N_8469,N_7914);
nand U9734 (N_9734,N_8304,N_7598);
nand U9735 (N_9735,N_8162,N_8474);
nor U9736 (N_9736,N_7855,N_8320);
nor U9737 (N_9737,N_8204,N_8274);
or U9738 (N_9738,N_8031,N_7711);
nand U9739 (N_9739,N_8830,N_8433);
nand U9740 (N_9740,N_8739,N_7563);
nor U9741 (N_9741,N_8139,N_8634);
nor U9742 (N_9742,N_7825,N_7682);
and U9743 (N_9743,N_8714,N_8608);
and U9744 (N_9744,N_8401,N_7601);
xnor U9745 (N_9745,N_8239,N_8338);
or U9746 (N_9746,N_8738,N_8898);
and U9747 (N_9747,N_7540,N_7755);
or U9748 (N_9748,N_8952,N_7841);
or U9749 (N_9749,N_8878,N_8025);
or U9750 (N_9750,N_8473,N_8013);
or U9751 (N_9751,N_8462,N_8547);
nand U9752 (N_9752,N_7946,N_8964);
or U9753 (N_9753,N_8382,N_8114);
nand U9754 (N_9754,N_8964,N_8744);
and U9755 (N_9755,N_8036,N_8756);
and U9756 (N_9756,N_8059,N_7868);
nor U9757 (N_9757,N_8238,N_8911);
nor U9758 (N_9758,N_7908,N_8466);
nand U9759 (N_9759,N_8142,N_8949);
or U9760 (N_9760,N_7804,N_8366);
nor U9761 (N_9761,N_8537,N_8413);
nand U9762 (N_9762,N_8268,N_8683);
nor U9763 (N_9763,N_8222,N_8010);
nand U9764 (N_9764,N_8434,N_8489);
and U9765 (N_9765,N_8238,N_7720);
and U9766 (N_9766,N_8667,N_8304);
and U9767 (N_9767,N_7817,N_8738);
nand U9768 (N_9768,N_7569,N_8304);
and U9769 (N_9769,N_7532,N_7701);
xnor U9770 (N_9770,N_8277,N_7763);
or U9771 (N_9771,N_8551,N_8179);
nand U9772 (N_9772,N_8351,N_7922);
or U9773 (N_9773,N_8317,N_8676);
and U9774 (N_9774,N_8509,N_8992);
nand U9775 (N_9775,N_7674,N_8652);
nand U9776 (N_9776,N_8790,N_8384);
and U9777 (N_9777,N_8289,N_7932);
and U9778 (N_9778,N_7618,N_8654);
or U9779 (N_9779,N_8981,N_7756);
nor U9780 (N_9780,N_7693,N_7630);
or U9781 (N_9781,N_8376,N_8899);
and U9782 (N_9782,N_7993,N_8075);
and U9783 (N_9783,N_8203,N_8362);
nor U9784 (N_9784,N_8592,N_7992);
nor U9785 (N_9785,N_8630,N_8112);
nor U9786 (N_9786,N_8893,N_8415);
nand U9787 (N_9787,N_8500,N_8114);
or U9788 (N_9788,N_7738,N_8946);
nor U9789 (N_9789,N_8681,N_8504);
and U9790 (N_9790,N_8226,N_8616);
and U9791 (N_9791,N_7612,N_8766);
nor U9792 (N_9792,N_7951,N_7937);
and U9793 (N_9793,N_8234,N_7651);
and U9794 (N_9794,N_7818,N_7527);
or U9795 (N_9795,N_7774,N_8045);
nand U9796 (N_9796,N_7944,N_8750);
nor U9797 (N_9797,N_7806,N_8006);
nand U9798 (N_9798,N_7775,N_8562);
nor U9799 (N_9799,N_8869,N_8466);
nor U9800 (N_9800,N_8852,N_8091);
nor U9801 (N_9801,N_7757,N_8285);
nand U9802 (N_9802,N_8116,N_8950);
nand U9803 (N_9803,N_7771,N_8533);
nor U9804 (N_9804,N_8021,N_7725);
nand U9805 (N_9805,N_8507,N_8004);
nor U9806 (N_9806,N_8150,N_8808);
nand U9807 (N_9807,N_8051,N_7655);
nor U9808 (N_9808,N_8484,N_8080);
nand U9809 (N_9809,N_7852,N_7534);
or U9810 (N_9810,N_8705,N_8318);
nand U9811 (N_9811,N_8632,N_8147);
and U9812 (N_9812,N_7725,N_7936);
or U9813 (N_9813,N_7537,N_7970);
nand U9814 (N_9814,N_8427,N_8990);
and U9815 (N_9815,N_7903,N_8226);
or U9816 (N_9816,N_7792,N_8208);
or U9817 (N_9817,N_8702,N_8546);
nand U9818 (N_9818,N_7547,N_8170);
or U9819 (N_9819,N_8159,N_8542);
or U9820 (N_9820,N_8416,N_8214);
nor U9821 (N_9821,N_8462,N_8082);
and U9822 (N_9822,N_7899,N_7610);
nor U9823 (N_9823,N_8598,N_8223);
nor U9824 (N_9824,N_7570,N_8556);
or U9825 (N_9825,N_8097,N_7644);
or U9826 (N_9826,N_7598,N_8772);
nor U9827 (N_9827,N_8946,N_8452);
nor U9828 (N_9828,N_8702,N_8291);
nand U9829 (N_9829,N_8115,N_8754);
or U9830 (N_9830,N_8754,N_8475);
nor U9831 (N_9831,N_8909,N_8902);
nand U9832 (N_9832,N_8628,N_8879);
or U9833 (N_9833,N_8492,N_7973);
nor U9834 (N_9834,N_8210,N_8123);
or U9835 (N_9835,N_8157,N_7793);
and U9836 (N_9836,N_7810,N_8545);
nor U9837 (N_9837,N_7693,N_8256);
nor U9838 (N_9838,N_8504,N_8415);
nor U9839 (N_9839,N_7937,N_8153);
nor U9840 (N_9840,N_8064,N_7782);
nand U9841 (N_9841,N_8475,N_8068);
and U9842 (N_9842,N_8185,N_8511);
nand U9843 (N_9843,N_7884,N_8350);
and U9844 (N_9844,N_8455,N_8911);
or U9845 (N_9845,N_8355,N_8034);
nand U9846 (N_9846,N_7888,N_8497);
nor U9847 (N_9847,N_8355,N_8884);
nand U9848 (N_9848,N_8921,N_7864);
or U9849 (N_9849,N_7667,N_8988);
nor U9850 (N_9850,N_7641,N_7513);
or U9851 (N_9851,N_8544,N_7990);
nor U9852 (N_9852,N_7685,N_7740);
or U9853 (N_9853,N_8833,N_8665);
and U9854 (N_9854,N_8421,N_7942);
nand U9855 (N_9855,N_8149,N_7988);
nor U9856 (N_9856,N_7923,N_7924);
nand U9857 (N_9857,N_7554,N_7918);
nand U9858 (N_9858,N_8001,N_8708);
or U9859 (N_9859,N_8227,N_8219);
or U9860 (N_9860,N_8920,N_8818);
nor U9861 (N_9861,N_7620,N_8319);
or U9862 (N_9862,N_8243,N_8785);
and U9863 (N_9863,N_8997,N_8158);
and U9864 (N_9864,N_8062,N_8300);
nor U9865 (N_9865,N_8852,N_7937);
nor U9866 (N_9866,N_8575,N_7503);
nand U9867 (N_9867,N_8357,N_7910);
nand U9868 (N_9868,N_8213,N_7597);
or U9869 (N_9869,N_7510,N_8938);
and U9870 (N_9870,N_8166,N_7673);
and U9871 (N_9871,N_8471,N_8931);
or U9872 (N_9872,N_8975,N_8448);
and U9873 (N_9873,N_8425,N_8921);
or U9874 (N_9874,N_7758,N_8315);
nor U9875 (N_9875,N_7843,N_8468);
or U9876 (N_9876,N_8788,N_8936);
nand U9877 (N_9877,N_8382,N_8223);
and U9878 (N_9878,N_8387,N_7795);
or U9879 (N_9879,N_8665,N_8661);
nand U9880 (N_9880,N_8228,N_8081);
nor U9881 (N_9881,N_8305,N_7965);
nor U9882 (N_9882,N_7785,N_8880);
and U9883 (N_9883,N_8737,N_8766);
or U9884 (N_9884,N_7912,N_7536);
nand U9885 (N_9885,N_8924,N_7749);
and U9886 (N_9886,N_7549,N_8503);
or U9887 (N_9887,N_8187,N_7609);
nor U9888 (N_9888,N_7749,N_8487);
and U9889 (N_9889,N_8760,N_8704);
nand U9890 (N_9890,N_7542,N_8647);
nand U9891 (N_9891,N_8573,N_7974);
nor U9892 (N_9892,N_7894,N_7853);
or U9893 (N_9893,N_8149,N_7880);
nor U9894 (N_9894,N_8489,N_7654);
nor U9895 (N_9895,N_8935,N_8596);
or U9896 (N_9896,N_8913,N_7719);
nand U9897 (N_9897,N_8097,N_8294);
and U9898 (N_9898,N_8448,N_8636);
and U9899 (N_9899,N_8117,N_8048);
nand U9900 (N_9900,N_7965,N_8026);
nand U9901 (N_9901,N_8354,N_8630);
and U9902 (N_9902,N_8549,N_8928);
and U9903 (N_9903,N_7713,N_8148);
or U9904 (N_9904,N_8826,N_8524);
or U9905 (N_9905,N_8268,N_7866);
nand U9906 (N_9906,N_7671,N_7680);
nand U9907 (N_9907,N_8021,N_8702);
or U9908 (N_9908,N_7669,N_8335);
or U9909 (N_9909,N_8573,N_7532);
and U9910 (N_9910,N_8852,N_7884);
or U9911 (N_9911,N_8104,N_8885);
nor U9912 (N_9912,N_8279,N_7553);
nand U9913 (N_9913,N_8525,N_7965);
nor U9914 (N_9914,N_7901,N_8922);
and U9915 (N_9915,N_8061,N_8558);
and U9916 (N_9916,N_8697,N_8300);
and U9917 (N_9917,N_7789,N_8248);
and U9918 (N_9918,N_8256,N_7825);
and U9919 (N_9919,N_7837,N_7523);
nand U9920 (N_9920,N_7677,N_7594);
nand U9921 (N_9921,N_8954,N_8245);
nor U9922 (N_9922,N_7592,N_7656);
and U9923 (N_9923,N_7556,N_7736);
nor U9924 (N_9924,N_8995,N_8248);
nor U9925 (N_9925,N_8339,N_7855);
or U9926 (N_9926,N_8320,N_7864);
or U9927 (N_9927,N_8354,N_8431);
or U9928 (N_9928,N_8685,N_8594);
or U9929 (N_9929,N_8264,N_8698);
nand U9930 (N_9930,N_8497,N_8480);
or U9931 (N_9931,N_7595,N_8781);
or U9932 (N_9932,N_8815,N_7719);
and U9933 (N_9933,N_8532,N_7948);
nand U9934 (N_9934,N_8490,N_8272);
xnor U9935 (N_9935,N_7986,N_8306);
and U9936 (N_9936,N_8811,N_7974);
nor U9937 (N_9937,N_8054,N_8333);
nand U9938 (N_9938,N_8297,N_8636);
and U9939 (N_9939,N_8140,N_7755);
or U9940 (N_9940,N_7986,N_8859);
nor U9941 (N_9941,N_8320,N_8881);
and U9942 (N_9942,N_8256,N_7818);
nor U9943 (N_9943,N_8484,N_8118);
or U9944 (N_9944,N_7882,N_8413);
or U9945 (N_9945,N_8944,N_7532);
or U9946 (N_9946,N_8668,N_8394);
and U9947 (N_9947,N_8359,N_8186);
nor U9948 (N_9948,N_8187,N_8097);
or U9949 (N_9949,N_7735,N_8702);
or U9950 (N_9950,N_8047,N_8327);
nor U9951 (N_9951,N_8290,N_7781);
or U9952 (N_9952,N_8773,N_8868);
nor U9953 (N_9953,N_7881,N_8663);
nor U9954 (N_9954,N_8829,N_7547);
nor U9955 (N_9955,N_7724,N_8017);
nand U9956 (N_9956,N_8255,N_7760);
and U9957 (N_9957,N_8209,N_8466);
nor U9958 (N_9958,N_8105,N_7828);
nand U9959 (N_9959,N_7624,N_8765);
or U9960 (N_9960,N_8560,N_7550);
and U9961 (N_9961,N_8404,N_8051);
nor U9962 (N_9962,N_8302,N_7578);
and U9963 (N_9963,N_8215,N_8915);
and U9964 (N_9964,N_7545,N_7848);
nand U9965 (N_9965,N_8266,N_8405);
and U9966 (N_9966,N_8360,N_8838);
nand U9967 (N_9967,N_8596,N_7940);
or U9968 (N_9968,N_7796,N_7567);
or U9969 (N_9969,N_8179,N_8623);
nand U9970 (N_9970,N_8472,N_7797);
or U9971 (N_9971,N_8395,N_8528);
or U9972 (N_9972,N_8715,N_8562);
or U9973 (N_9973,N_8508,N_8439);
nand U9974 (N_9974,N_8021,N_7971);
nand U9975 (N_9975,N_8690,N_7803);
and U9976 (N_9976,N_7970,N_7883);
and U9977 (N_9977,N_7958,N_7959);
and U9978 (N_9978,N_8611,N_8724);
or U9979 (N_9979,N_8245,N_8713);
and U9980 (N_9980,N_8964,N_8383);
and U9981 (N_9981,N_7956,N_8424);
or U9982 (N_9982,N_8582,N_8711);
and U9983 (N_9983,N_7958,N_8174);
or U9984 (N_9984,N_8520,N_8328);
nand U9985 (N_9985,N_8660,N_8080);
and U9986 (N_9986,N_7660,N_8631);
or U9987 (N_9987,N_8062,N_7865);
and U9988 (N_9988,N_7541,N_7876);
xnor U9989 (N_9989,N_7529,N_7606);
nor U9990 (N_9990,N_7722,N_8062);
nor U9991 (N_9991,N_8231,N_7753);
and U9992 (N_9992,N_7608,N_8859);
nand U9993 (N_9993,N_7688,N_7847);
or U9994 (N_9994,N_8678,N_8397);
nand U9995 (N_9995,N_8263,N_8691);
or U9996 (N_9996,N_8854,N_8058);
or U9997 (N_9997,N_8866,N_8072);
or U9998 (N_9998,N_8799,N_8222);
nand U9999 (N_9999,N_8035,N_8418);
nor U10000 (N_10000,N_7961,N_7872);
or U10001 (N_10001,N_7802,N_8114);
nor U10002 (N_10002,N_8858,N_8679);
and U10003 (N_10003,N_7816,N_7595);
or U10004 (N_10004,N_8834,N_8805);
nand U10005 (N_10005,N_8297,N_8196);
nor U10006 (N_10006,N_8341,N_8083);
nand U10007 (N_10007,N_8591,N_8709);
nor U10008 (N_10008,N_7951,N_7586);
nor U10009 (N_10009,N_8883,N_8166);
nor U10010 (N_10010,N_7949,N_7780);
xor U10011 (N_10011,N_8811,N_8404);
or U10012 (N_10012,N_7786,N_7836);
nor U10013 (N_10013,N_8528,N_8363);
and U10014 (N_10014,N_7733,N_7624);
nand U10015 (N_10015,N_8974,N_8421);
nand U10016 (N_10016,N_8731,N_7609);
nor U10017 (N_10017,N_7519,N_8768);
or U10018 (N_10018,N_8668,N_8428);
or U10019 (N_10019,N_8711,N_8733);
or U10020 (N_10020,N_7603,N_8197);
or U10021 (N_10021,N_8180,N_8531);
or U10022 (N_10022,N_8992,N_8243);
and U10023 (N_10023,N_7629,N_8119);
nor U10024 (N_10024,N_8937,N_7899);
nand U10025 (N_10025,N_7643,N_8204);
nand U10026 (N_10026,N_7768,N_7513);
and U10027 (N_10027,N_7883,N_8062);
nor U10028 (N_10028,N_7777,N_8924);
or U10029 (N_10029,N_8804,N_7862);
and U10030 (N_10030,N_8673,N_8321);
or U10031 (N_10031,N_8688,N_8352);
nand U10032 (N_10032,N_8974,N_7879);
or U10033 (N_10033,N_8952,N_7554);
nand U10034 (N_10034,N_7619,N_8610);
nor U10035 (N_10035,N_8275,N_8187);
and U10036 (N_10036,N_7615,N_8608);
or U10037 (N_10037,N_7855,N_8677);
nand U10038 (N_10038,N_8129,N_8875);
and U10039 (N_10039,N_8832,N_8505);
and U10040 (N_10040,N_8872,N_7757);
and U10041 (N_10041,N_8442,N_8597);
nor U10042 (N_10042,N_8864,N_8442);
nor U10043 (N_10043,N_7571,N_8562);
nor U10044 (N_10044,N_8363,N_7677);
and U10045 (N_10045,N_7742,N_8363);
nor U10046 (N_10046,N_8556,N_8099);
nor U10047 (N_10047,N_8822,N_7788);
nand U10048 (N_10048,N_8385,N_7924);
nor U10049 (N_10049,N_8211,N_7948);
nand U10050 (N_10050,N_8178,N_8416);
nand U10051 (N_10051,N_8120,N_8038);
nand U10052 (N_10052,N_7849,N_7699);
nor U10053 (N_10053,N_8418,N_8911);
nand U10054 (N_10054,N_8088,N_7584);
and U10055 (N_10055,N_8329,N_8753);
nor U10056 (N_10056,N_7546,N_8486);
and U10057 (N_10057,N_8117,N_8812);
or U10058 (N_10058,N_8957,N_7501);
nor U10059 (N_10059,N_8210,N_8961);
nand U10060 (N_10060,N_8384,N_8189);
or U10061 (N_10061,N_8218,N_8756);
and U10062 (N_10062,N_8938,N_8057);
nand U10063 (N_10063,N_7995,N_8566);
or U10064 (N_10064,N_8911,N_8902);
or U10065 (N_10065,N_8452,N_8650);
and U10066 (N_10066,N_8807,N_8075);
nor U10067 (N_10067,N_7539,N_8027);
and U10068 (N_10068,N_7861,N_7774);
nor U10069 (N_10069,N_7780,N_8855);
nor U10070 (N_10070,N_7776,N_8799);
and U10071 (N_10071,N_8511,N_8490);
or U10072 (N_10072,N_8399,N_7559);
or U10073 (N_10073,N_7542,N_8883);
and U10074 (N_10074,N_7699,N_7909);
or U10075 (N_10075,N_7925,N_8191);
or U10076 (N_10076,N_8872,N_8906);
nor U10077 (N_10077,N_8159,N_8592);
nor U10078 (N_10078,N_8013,N_7678);
nand U10079 (N_10079,N_8963,N_8359);
nor U10080 (N_10080,N_7895,N_8118);
nand U10081 (N_10081,N_8459,N_8645);
or U10082 (N_10082,N_8305,N_8076);
nand U10083 (N_10083,N_8023,N_8184);
nor U10084 (N_10084,N_7945,N_7593);
and U10085 (N_10085,N_8232,N_8560);
nand U10086 (N_10086,N_8311,N_8459);
nand U10087 (N_10087,N_7774,N_8964);
and U10088 (N_10088,N_8132,N_8585);
or U10089 (N_10089,N_7794,N_8973);
and U10090 (N_10090,N_7752,N_8655);
and U10091 (N_10091,N_7640,N_8555);
nor U10092 (N_10092,N_8824,N_8410);
nor U10093 (N_10093,N_7737,N_8762);
nand U10094 (N_10094,N_8078,N_8298);
and U10095 (N_10095,N_8340,N_7791);
and U10096 (N_10096,N_8424,N_8714);
and U10097 (N_10097,N_8916,N_8334);
nor U10098 (N_10098,N_7541,N_8440);
and U10099 (N_10099,N_8947,N_8659);
or U10100 (N_10100,N_7665,N_8836);
or U10101 (N_10101,N_8643,N_8850);
and U10102 (N_10102,N_8381,N_8474);
and U10103 (N_10103,N_8116,N_8135);
nand U10104 (N_10104,N_8665,N_8797);
nor U10105 (N_10105,N_8160,N_7703);
and U10106 (N_10106,N_7594,N_8545);
nor U10107 (N_10107,N_8797,N_8088);
xor U10108 (N_10108,N_8731,N_8049);
nor U10109 (N_10109,N_7606,N_7781);
nor U10110 (N_10110,N_8110,N_7709);
and U10111 (N_10111,N_8618,N_8770);
or U10112 (N_10112,N_7954,N_8999);
or U10113 (N_10113,N_8658,N_7760);
and U10114 (N_10114,N_8894,N_8577);
nor U10115 (N_10115,N_8865,N_8819);
nand U10116 (N_10116,N_7515,N_7994);
nand U10117 (N_10117,N_8911,N_8876);
nand U10118 (N_10118,N_8519,N_8746);
and U10119 (N_10119,N_8035,N_8037);
nand U10120 (N_10120,N_7556,N_8712);
nand U10121 (N_10121,N_8776,N_8413);
nand U10122 (N_10122,N_7993,N_8170);
or U10123 (N_10123,N_7619,N_8948);
nor U10124 (N_10124,N_8128,N_8915);
or U10125 (N_10125,N_8223,N_8222);
or U10126 (N_10126,N_8324,N_8009);
nand U10127 (N_10127,N_8450,N_7739);
nor U10128 (N_10128,N_7855,N_8939);
or U10129 (N_10129,N_8592,N_8440);
and U10130 (N_10130,N_8246,N_7849);
and U10131 (N_10131,N_8496,N_8346);
nor U10132 (N_10132,N_8717,N_8909);
nand U10133 (N_10133,N_7685,N_7691);
nor U10134 (N_10134,N_8344,N_7636);
or U10135 (N_10135,N_8565,N_8818);
and U10136 (N_10136,N_8312,N_7652);
nor U10137 (N_10137,N_7768,N_8373);
nand U10138 (N_10138,N_8952,N_7732);
or U10139 (N_10139,N_8570,N_8836);
nor U10140 (N_10140,N_8935,N_8303);
nor U10141 (N_10141,N_8230,N_8721);
or U10142 (N_10142,N_7618,N_8316);
and U10143 (N_10143,N_8288,N_8010);
nor U10144 (N_10144,N_7616,N_8188);
or U10145 (N_10145,N_8424,N_8475);
nor U10146 (N_10146,N_7884,N_8543);
nor U10147 (N_10147,N_8693,N_8714);
or U10148 (N_10148,N_8684,N_7513);
nor U10149 (N_10149,N_8188,N_8950);
or U10150 (N_10150,N_8841,N_8024);
nor U10151 (N_10151,N_7690,N_7908);
nand U10152 (N_10152,N_8262,N_7825);
and U10153 (N_10153,N_7974,N_7810);
nand U10154 (N_10154,N_8284,N_7793);
nor U10155 (N_10155,N_8208,N_8248);
and U10156 (N_10156,N_8412,N_8977);
or U10157 (N_10157,N_8745,N_8847);
or U10158 (N_10158,N_8687,N_8988);
or U10159 (N_10159,N_8666,N_8785);
nand U10160 (N_10160,N_8822,N_8213);
or U10161 (N_10161,N_8063,N_8603);
and U10162 (N_10162,N_8017,N_7888);
and U10163 (N_10163,N_7514,N_8123);
or U10164 (N_10164,N_8354,N_8622);
nand U10165 (N_10165,N_7694,N_8914);
and U10166 (N_10166,N_7779,N_8006);
nand U10167 (N_10167,N_7729,N_8873);
and U10168 (N_10168,N_8099,N_8574);
nor U10169 (N_10169,N_8406,N_7707);
and U10170 (N_10170,N_7696,N_7770);
nor U10171 (N_10171,N_7827,N_8352);
nand U10172 (N_10172,N_8079,N_7541);
nor U10173 (N_10173,N_8734,N_8132);
nor U10174 (N_10174,N_8909,N_8045);
and U10175 (N_10175,N_8007,N_8798);
nand U10176 (N_10176,N_7720,N_7501);
or U10177 (N_10177,N_7728,N_8224);
and U10178 (N_10178,N_8641,N_7548);
xnor U10179 (N_10179,N_8415,N_7579);
nand U10180 (N_10180,N_8170,N_7580);
and U10181 (N_10181,N_8118,N_7966);
nor U10182 (N_10182,N_7951,N_7572);
nor U10183 (N_10183,N_8002,N_8148);
nand U10184 (N_10184,N_8880,N_7653);
nor U10185 (N_10185,N_7547,N_8950);
nand U10186 (N_10186,N_8734,N_7731);
or U10187 (N_10187,N_7693,N_7884);
nor U10188 (N_10188,N_8251,N_7887);
nand U10189 (N_10189,N_8697,N_8931);
and U10190 (N_10190,N_8919,N_7979);
or U10191 (N_10191,N_8844,N_8303);
nor U10192 (N_10192,N_8346,N_8744);
nand U10193 (N_10193,N_8329,N_8768);
nor U10194 (N_10194,N_8250,N_7746);
nor U10195 (N_10195,N_8318,N_8165);
and U10196 (N_10196,N_8922,N_8244);
or U10197 (N_10197,N_8309,N_7906);
nand U10198 (N_10198,N_7947,N_7826);
nand U10199 (N_10199,N_8089,N_8685);
nor U10200 (N_10200,N_7873,N_8739);
nor U10201 (N_10201,N_8100,N_8250);
nand U10202 (N_10202,N_8157,N_7853);
nor U10203 (N_10203,N_8759,N_8563);
or U10204 (N_10204,N_8912,N_7503);
nand U10205 (N_10205,N_8462,N_8904);
nand U10206 (N_10206,N_7908,N_8978);
or U10207 (N_10207,N_8214,N_8754);
and U10208 (N_10208,N_7985,N_8391);
nor U10209 (N_10209,N_8211,N_8337);
nand U10210 (N_10210,N_8887,N_7582);
nor U10211 (N_10211,N_8678,N_8783);
and U10212 (N_10212,N_8036,N_8850);
and U10213 (N_10213,N_8220,N_7608);
nor U10214 (N_10214,N_8115,N_8206);
xnor U10215 (N_10215,N_7841,N_8575);
or U10216 (N_10216,N_7753,N_8471);
or U10217 (N_10217,N_8714,N_8445);
nand U10218 (N_10218,N_8664,N_8040);
nand U10219 (N_10219,N_8374,N_7990);
nor U10220 (N_10220,N_8528,N_8368);
or U10221 (N_10221,N_7521,N_8249);
nand U10222 (N_10222,N_8596,N_8978);
or U10223 (N_10223,N_8276,N_8226);
and U10224 (N_10224,N_7860,N_8505);
and U10225 (N_10225,N_8519,N_8982);
and U10226 (N_10226,N_8005,N_7973);
or U10227 (N_10227,N_8609,N_7899);
and U10228 (N_10228,N_7910,N_8361);
nor U10229 (N_10229,N_7635,N_8345);
or U10230 (N_10230,N_8366,N_7968);
nand U10231 (N_10231,N_8072,N_8028);
or U10232 (N_10232,N_7723,N_8314);
and U10233 (N_10233,N_8381,N_8760);
nor U10234 (N_10234,N_7701,N_8279);
and U10235 (N_10235,N_7518,N_8072);
nor U10236 (N_10236,N_8958,N_8202);
or U10237 (N_10237,N_7945,N_8221);
nor U10238 (N_10238,N_7506,N_8872);
nor U10239 (N_10239,N_8172,N_8041);
nor U10240 (N_10240,N_8309,N_8943);
or U10241 (N_10241,N_7502,N_7920);
and U10242 (N_10242,N_8121,N_8918);
nor U10243 (N_10243,N_7975,N_8377);
nor U10244 (N_10244,N_8298,N_7955);
and U10245 (N_10245,N_8741,N_8252);
nand U10246 (N_10246,N_8503,N_7586);
nor U10247 (N_10247,N_7594,N_7566);
and U10248 (N_10248,N_8797,N_8695);
and U10249 (N_10249,N_8090,N_8109);
and U10250 (N_10250,N_8174,N_8990);
or U10251 (N_10251,N_7943,N_7759);
nor U10252 (N_10252,N_8508,N_8455);
nor U10253 (N_10253,N_8808,N_8856);
and U10254 (N_10254,N_8981,N_7861);
nor U10255 (N_10255,N_8824,N_7638);
and U10256 (N_10256,N_8803,N_8532);
nand U10257 (N_10257,N_8552,N_8604);
and U10258 (N_10258,N_7924,N_7846);
xnor U10259 (N_10259,N_7992,N_8723);
and U10260 (N_10260,N_7779,N_7796);
nor U10261 (N_10261,N_7519,N_7961);
and U10262 (N_10262,N_8959,N_7689);
nor U10263 (N_10263,N_8418,N_8945);
and U10264 (N_10264,N_7832,N_8273);
and U10265 (N_10265,N_8538,N_8844);
nor U10266 (N_10266,N_8995,N_8491);
and U10267 (N_10267,N_8527,N_8275);
nor U10268 (N_10268,N_7752,N_7689);
or U10269 (N_10269,N_7856,N_8929);
nand U10270 (N_10270,N_8146,N_8484);
or U10271 (N_10271,N_8476,N_8956);
nand U10272 (N_10272,N_8541,N_8848);
or U10273 (N_10273,N_8465,N_8996);
nand U10274 (N_10274,N_8592,N_7913);
and U10275 (N_10275,N_8568,N_8434);
nand U10276 (N_10276,N_8970,N_7923);
nor U10277 (N_10277,N_8267,N_8299);
and U10278 (N_10278,N_8566,N_7597);
and U10279 (N_10279,N_8567,N_8635);
nand U10280 (N_10280,N_8435,N_7807);
nand U10281 (N_10281,N_8999,N_8110);
or U10282 (N_10282,N_8621,N_8078);
or U10283 (N_10283,N_8557,N_7622);
nand U10284 (N_10284,N_7676,N_7956);
and U10285 (N_10285,N_8193,N_7619);
or U10286 (N_10286,N_8087,N_7924);
or U10287 (N_10287,N_7820,N_7595);
or U10288 (N_10288,N_8264,N_8527);
or U10289 (N_10289,N_7890,N_8036);
or U10290 (N_10290,N_8599,N_8442);
or U10291 (N_10291,N_8880,N_8999);
nand U10292 (N_10292,N_8767,N_7751);
or U10293 (N_10293,N_8332,N_8483);
nor U10294 (N_10294,N_8668,N_8600);
nor U10295 (N_10295,N_8001,N_8103);
or U10296 (N_10296,N_8581,N_7600);
or U10297 (N_10297,N_8981,N_8205);
or U10298 (N_10298,N_7995,N_8244);
or U10299 (N_10299,N_8056,N_8414);
or U10300 (N_10300,N_8289,N_8320);
or U10301 (N_10301,N_7791,N_8223);
and U10302 (N_10302,N_8244,N_7815);
and U10303 (N_10303,N_7624,N_8949);
and U10304 (N_10304,N_7875,N_8146);
and U10305 (N_10305,N_7920,N_8687);
nand U10306 (N_10306,N_7817,N_7700);
nor U10307 (N_10307,N_8740,N_7867);
nand U10308 (N_10308,N_7767,N_7859);
and U10309 (N_10309,N_7832,N_7706);
or U10310 (N_10310,N_8167,N_8475);
and U10311 (N_10311,N_8519,N_7639);
nand U10312 (N_10312,N_7778,N_8359);
nand U10313 (N_10313,N_8620,N_8437);
or U10314 (N_10314,N_8158,N_8605);
or U10315 (N_10315,N_8249,N_7652);
nor U10316 (N_10316,N_8158,N_8121);
and U10317 (N_10317,N_8607,N_8061);
nor U10318 (N_10318,N_8452,N_8227);
and U10319 (N_10319,N_8636,N_8660);
nand U10320 (N_10320,N_8202,N_7619);
and U10321 (N_10321,N_8440,N_8728);
or U10322 (N_10322,N_7833,N_8582);
and U10323 (N_10323,N_7964,N_8298);
and U10324 (N_10324,N_8889,N_8754);
nand U10325 (N_10325,N_8391,N_8213);
and U10326 (N_10326,N_8512,N_7845);
and U10327 (N_10327,N_7792,N_8446);
xnor U10328 (N_10328,N_7923,N_7793);
nor U10329 (N_10329,N_8848,N_7862);
or U10330 (N_10330,N_8511,N_8975);
nand U10331 (N_10331,N_8440,N_8908);
nand U10332 (N_10332,N_8156,N_8466);
or U10333 (N_10333,N_8595,N_8129);
or U10334 (N_10334,N_8066,N_8537);
nand U10335 (N_10335,N_8267,N_8564);
or U10336 (N_10336,N_8717,N_7760);
nand U10337 (N_10337,N_8004,N_8266);
and U10338 (N_10338,N_7665,N_8721);
nand U10339 (N_10339,N_8596,N_8765);
and U10340 (N_10340,N_8694,N_7753);
or U10341 (N_10341,N_8709,N_7678);
nand U10342 (N_10342,N_7509,N_8224);
and U10343 (N_10343,N_8703,N_8216);
nand U10344 (N_10344,N_7727,N_8346);
nor U10345 (N_10345,N_7820,N_7766);
nand U10346 (N_10346,N_8491,N_8060);
nand U10347 (N_10347,N_7770,N_8544);
nor U10348 (N_10348,N_7978,N_8405);
and U10349 (N_10349,N_8967,N_7537);
and U10350 (N_10350,N_8415,N_7581);
and U10351 (N_10351,N_8886,N_8600);
nor U10352 (N_10352,N_8205,N_8900);
nand U10353 (N_10353,N_7694,N_7848);
nor U10354 (N_10354,N_7890,N_7704);
or U10355 (N_10355,N_7618,N_8432);
nand U10356 (N_10356,N_7883,N_7623);
nor U10357 (N_10357,N_8583,N_7785);
or U10358 (N_10358,N_7779,N_7780);
and U10359 (N_10359,N_8498,N_8707);
or U10360 (N_10360,N_8252,N_8743);
or U10361 (N_10361,N_7958,N_8442);
and U10362 (N_10362,N_8919,N_7862);
or U10363 (N_10363,N_8622,N_7658);
and U10364 (N_10364,N_7903,N_7593);
nor U10365 (N_10365,N_8887,N_8348);
and U10366 (N_10366,N_8600,N_8906);
nor U10367 (N_10367,N_8825,N_7961);
xor U10368 (N_10368,N_8491,N_8949);
and U10369 (N_10369,N_8147,N_7856);
nor U10370 (N_10370,N_8393,N_8597);
and U10371 (N_10371,N_8670,N_8146);
nand U10372 (N_10372,N_8098,N_8699);
and U10373 (N_10373,N_7696,N_7992);
or U10374 (N_10374,N_8982,N_7669);
nor U10375 (N_10375,N_8897,N_8821);
nand U10376 (N_10376,N_8177,N_7949);
and U10377 (N_10377,N_8394,N_8216);
and U10378 (N_10378,N_8425,N_7646);
nor U10379 (N_10379,N_7594,N_8957);
and U10380 (N_10380,N_8669,N_7927);
and U10381 (N_10381,N_8468,N_7509);
and U10382 (N_10382,N_8750,N_7938);
nand U10383 (N_10383,N_7914,N_7804);
nor U10384 (N_10384,N_8507,N_8895);
and U10385 (N_10385,N_8709,N_8566);
or U10386 (N_10386,N_7910,N_7575);
or U10387 (N_10387,N_7514,N_8441);
or U10388 (N_10388,N_7551,N_8696);
nor U10389 (N_10389,N_8322,N_8848);
and U10390 (N_10390,N_8127,N_8233);
or U10391 (N_10391,N_7680,N_8773);
nor U10392 (N_10392,N_7561,N_8428);
or U10393 (N_10393,N_7965,N_7966);
nor U10394 (N_10394,N_7919,N_8888);
and U10395 (N_10395,N_8953,N_7779);
nor U10396 (N_10396,N_8894,N_8186);
or U10397 (N_10397,N_8595,N_8929);
or U10398 (N_10398,N_8339,N_7642);
and U10399 (N_10399,N_8953,N_8005);
nor U10400 (N_10400,N_8447,N_8595);
and U10401 (N_10401,N_8080,N_8363);
or U10402 (N_10402,N_7609,N_7548);
or U10403 (N_10403,N_7676,N_8853);
nand U10404 (N_10404,N_8920,N_8919);
and U10405 (N_10405,N_7793,N_7748);
and U10406 (N_10406,N_8354,N_8204);
and U10407 (N_10407,N_7848,N_8381);
or U10408 (N_10408,N_7742,N_8627);
and U10409 (N_10409,N_8173,N_7883);
nand U10410 (N_10410,N_8956,N_8035);
and U10411 (N_10411,N_8986,N_8893);
or U10412 (N_10412,N_8357,N_8689);
nand U10413 (N_10413,N_8497,N_7825);
and U10414 (N_10414,N_8020,N_7763);
nor U10415 (N_10415,N_8280,N_8409);
and U10416 (N_10416,N_8491,N_8902);
and U10417 (N_10417,N_7898,N_8330);
or U10418 (N_10418,N_8174,N_8456);
nor U10419 (N_10419,N_7650,N_8837);
nand U10420 (N_10420,N_8608,N_8973);
nand U10421 (N_10421,N_8345,N_7963);
nand U10422 (N_10422,N_8166,N_8709);
nor U10423 (N_10423,N_7550,N_8156);
and U10424 (N_10424,N_8519,N_8816);
nand U10425 (N_10425,N_7688,N_8054);
or U10426 (N_10426,N_7880,N_8565);
nor U10427 (N_10427,N_8488,N_8028);
nand U10428 (N_10428,N_8066,N_8223);
nor U10429 (N_10429,N_8682,N_8018);
and U10430 (N_10430,N_7609,N_8464);
nor U10431 (N_10431,N_8030,N_8620);
nor U10432 (N_10432,N_7760,N_7690);
nor U10433 (N_10433,N_8356,N_7868);
nor U10434 (N_10434,N_8604,N_7706);
and U10435 (N_10435,N_8999,N_8569);
or U10436 (N_10436,N_7668,N_7709);
nand U10437 (N_10437,N_8948,N_8962);
nor U10438 (N_10438,N_8221,N_8615);
nand U10439 (N_10439,N_7634,N_8685);
or U10440 (N_10440,N_8765,N_8088);
nor U10441 (N_10441,N_7535,N_8478);
nor U10442 (N_10442,N_8493,N_7541);
xor U10443 (N_10443,N_8495,N_8133);
nor U10444 (N_10444,N_8279,N_8893);
or U10445 (N_10445,N_8564,N_7551);
nand U10446 (N_10446,N_7559,N_7914);
nor U10447 (N_10447,N_8327,N_7646);
or U10448 (N_10448,N_8900,N_8671);
and U10449 (N_10449,N_7575,N_8178);
nand U10450 (N_10450,N_8154,N_8116);
and U10451 (N_10451,N_7950,N_7862);
nor U10452 (N_10452,N_8236,N_8871);
or U10453 (N_10453,N_7507,N_8834);
nand U10454 (N_10454,N_8761,N_8479);
nor U10455 (N_10455,N_8493,N_8262);
nor U10456 (N_10456,N_8975,N_7532);
nor U10457 (N_10457,N_7705,N_8216);
nor U10458 (N_10458,N_7595,N_7763);
nand U10459 (N_10459,N_7920,N_8400);
nand U10460 (N_10460,N_7763,N_7760);
or U10461 (N_10461,N_7913,N_7531);
nor U10462 (N_10462,N_8136,N_8724);
nor U10463 (N_10463,N_7696,N_8594);
and U10464 (N_10464,N_7582,N_7716);
and U10465 (N_10465,N_8526,N_7647);
or U10466 (N_10466,N_8404,N_8859);
nand U10467 (N_10467,N_8841,N_7989);
nand U10468 (N_10468,N_8460,N_8289);
nor U10469 (N_10469,N_8161,N_7563);
or U10470 (N_10470,N_8120,N_7581);
nor U10471 (N_10471,N_7996,N_8425);
nand U10472 (N_10472,N_8731,N_8631);
and U10473 (N_10473,N_8569,N_7540);
or U10474 (N_10474,N_8017,N_7639);
or U10475 (N_10475,N_7659,N_8445);
nor U10476 (N_10476,N_8092,N_7787);
nand U10477 (N_10477,N_7750,N_8532);
or U10478 (N_10478,N_8988,N_8427);
and U10479 (N_10479,N_8222,N_7742);
and U10480 (N_10480,N_8407,N_8474);
nand U10481 (N_10481,N_7601,N_7890);
or U10482 (N_10482,N_7926,N_7833);
or U10483 (N_10483,N_8123,N_7671);
nor U10484 (N_10484,N_7851,N_7586);
nand U10485 (N_10485,N_8853,N_8846);
nor U10486 (N_10486,N_8796,N_7597);
or U10487 (N_10487,N_8791,N_8999);
nand U10488 (N_10488,N_7693,N_7783);
or U10489 (N_10489,N_8656,N_8743);
or U10490 (N_10490,N_8299,N_8608);
and U10491 (N_10491,N_7616,N_8314);
and U10492 (N_10492,N_8387,N_8613);
or U10493 (N_10493,N_8368,N_7528);
nor U10494 (N_10494,N_7899,N_8689);
or U10495 (N_10495,N_7762,N_8605);
and U10496 (N_10496,N_7605,N_7852);
and U10497 (N_10497,N_8039,N_7901);
or U10498 (N_10498,N_8537,N_7759);
nand U10499 (N_10499,N_7621,N_8894);
nor U10500 (N_10500,N_10225,N_9871);
or U10501 (N_10501,N_10039,N_9117);
nor U10502 (N_10502,N_9238,N_9365);
nand U10503 (N_10503,N_9360,N_9408);
or U10504 (N_10504,N_9152,N_9173);
and U10505 (N_10505,N_9830,N_10353);
or U10506 (N_10506,N_9386,N_9693);
or U10507 (N_10507,N_9392,N_10394);
nor U10508 (N_10508,N_10105,N_10324);
nand U10509 (N_10509,N_9624,N_9636);
and U10510 (N_10510,N_9083,N_9865);
nor U10511 (N_10511,N_10262,N_9981);
nand U10512 (N_10512,N_9121,N_10348);
nand U10513 (N_10513,N_10271,N_10159);
nand U10514 (N_10514,N_9047,N_10310);
nand U10515 (N_10515,N_10061,N_9382);
nor U10516 (N_10516,N_10493,N_9081);
nand U10517 (N_10517,N_9148,N_10465);
and U10518 (N_10518,N_9899,N_9416);
or U10519 (N_10519,N_9685,N_9485);
nand U10520 (N_10520,N_9023,N_10045);
and U10521 (N_10521,N_10043,N_9112);
or U10522 (N_10522,N_9293,N_10067);
nor U10523 (N_10523,N_10021,N_10094);
nor U10524 (N_10524,N_9477,N_9602);
nor U10525 (N_10525,N_10453,N_9944);
or U10526 (N_10526,N_9491,N_9253);
and U10527 (N_10527,N_9827,N_9336);
and U10528 (N_10528,N_10468,N_9858);
or U10529 (N_10529,N_9545,N_10035);
nand U10530 (N_10530,N_9998,N_9806);
nand U10531 (N_10531,N_9974,N_9953);
nand U10532 (N_10532,N_9913,N_9243);
xnor U10533 (N_10533,N_10008,N_9887);
nand U10534 (N_10534,N_9123,N_9478);
nor U10535 (N_10535,N_10054,N_9839);
or U10536 (N_10536,N_10098,N_9412);
and U10537 (N_10537,N_9332,N_10230);
nor U10538 (N_10538,N_9694,N_9218);
and U10539 (N_10539,N_9810,N_9769);
nor U10540 (N_10540,N_10025,N_10487);
or U10541 (N_10541,N_9284,N_9828);
nand U10542 (N_10542,N_10483,N_10250);
nand U10543 (N_10543,N_9215,N_9251);
or U10544 (N_10544,N_10325,N_10417);
and U10545 (N_10545,N_9580,N_10029);
nor U10546 (N_10546,N_9384,N_9246);
and U10547 (N_10547,N_9846,N_10090);
and U10548 (N_10548,N_10333,N_10226);
and U10549 (N_10549,N_10293,N_9468);
nor U10550 (N_10550,N_10488,N_9889);
and U10551 (N_10551,N_10278,N_9156);
nand U10552 (N_10552,N_10221,N_9305);
nand U10553 (N_10553,N_9473,N_9038);
nand U10554 (N_10554,N_9767,N_9629);
nand U10555 (N_10555,N_9594,N_9460);
nand U10556 (N_10556,N_9711,N_10119);
and U10557 (N_10557,N_9667,N_9946);
xor U10558 (N_10558,N_9054,N_9572);
or U10559 (N_10559,N_10466,N_9560);
and U10560 (N_10560,N_9228,N_9638);
nand U10561 (N_10561,N_9760,N_9955);
nand U10562 (N_10562,N_9322,N_9640);
and U10563 (N_10563,N_9024,N_9978);
nand U10564 (N_10564,N_9684,N_10138);
nand U10565 (N_10565,N_10038,N_10260);
or U10566 (N_10566,N_9682,N_9958);
and U10567 (N_10567,N_9564,N_9690);
or U10568 (N_10568,N_10192,N_9613);
or U10569 (N_10569,N_10133,N_9809);
nand U10570 (N_10570,N_9351,N_9844);
nor U10571 (N_10571,N_9942,N_9194);
or U10572 (N_10572,N_9724,N_10136);
nand U10573 (N_10573,N_10314,N_9597);
nand U10574 (N_10574,N_9713,N_9573);
and U10575 (N_10575,N_9774,N_9619);
nand U10576 (N_10576,N_9838,N_9183);
nor U10577 (N_10577,N_9303,N_9877);
nand U10578 (N_10578,N_9364,N_9330);
and U10579 (N_10579,N_9237,N_9453);
nor U10580 (N_10580,N_9455,N_10007);
and U10581 (N_10581,N_9298,N_10342);
nand U10582 (N_10582,N_10413,N_10396);
nor U10583 (N_10583,N_9107,N_10459);
or U10584 (N_10584,N_9299,N_9199);
and U10585 (N_10585,N_9239,N_9113);
or U10586 (N_10586,N_9527,N_10254);
nand U10587 (N_10587,N_9281,N_9983);
or U10588 (N_10588,N_9815,N_9072);
or U10589 (N_10589,N_9352,N_10452);
and U10590 (N_10590,N_10251,N_10264);
or U10591 (N_10591,N_9610,N_9224);
or U10592 (N_10592,N_9357,N_9862);
and U10593 (N_10593,N_10202,N_9503);
and U10594 (N_10594,N_9935,N_9302);
and U10595 (N_10595,N_10256,N_10084);
or U10596 (N_10596,N_10229,N_10241);
and U10597 (N_10597,N_9812,N_9067);
nand U10598 (N_10598,N_9504,N_9703);
nor U10599 (N_10599,N_9297,N_9556);
or U10600 (N_10600,N_9964,N_9449);
nor U10601 (N_10601,N_9311,N_9791);
and U10602 (N_10602,N_10438,N_9006);
and U10603 (N_10603,N_10183,N_9221);
nor U10604 (N_10604,N_9292,N_9617);
and U10605 (N_10605,N_9499,N_9139);
and U10606 (N_10606,N_9973,N_10266);
and U10607 (N_10607,N_9529,N_10199);
nor U10608 (N_10608,N_9487,N_9980);
nand U10609 (N_10609,N_9244,N_9456);
or U10610 (N_10610,N_9538,N_9732);
nand U10611 (N_10611,N_9296,N_9103);
nor U10612 (N_10612,N_10104,N_10498);
nand U10613 (N_10613,N_9821,N_9544);
nand U10614 (N_10614,N_9263,N_9999);
or U10615 (N_10615,N_9376,N_9648);
nor U10616 (N_10616,N_10321,N_9639);
nand U10617 (N_10617,N_10153,N_10197);
nor U10618 (N_10618,N_10435,N_10194);
and U10619 (N_10619,N_10462,N_9531);
nor U10620 (N_10620,N_9326,N_9581);
nor U10621 (N_10621,N_9756,N_9407);
nor U10622 (N_10622,N_9035,N_9454);
nand U10623 (N_10623,N_10288,N_10042);
nand U10624 (N_10624,N_10106,N_9133);
or U10625 (N_10625,N_9993,N_9982);
nor U10626 (N_10626,N_9151,N_10268);
nand U10627 (N_10627,N_9334,N_9200);
nor U10628 (N_10628,N_9055,N_9323);
nand U10629 (N_10629,N_9960,N_9938);
or U10630 (N_10630,N_9320,N_9385);
and U10631 (N_10631,N_9891,N_9344);
or U10632 (N_10632,N_9698,N_9071);
or U10633 (N_10633,N_9957,N_9161);
or U10634 (N_10634,N_9276,N_9442);
or U10635 (N_10635,N_10450,N_10274);
nor U10636 (N_10636,N_9971,N_9525);
nand U10637 (N_10637,N_9337,N_10422);
nor U10638 (N_10638,N_10441,N_9631);
or U10639 (N_10639,N_9737,N_9632);
nor U10640 (N_10640,N_9131,N_9608);
xnor U10641 (N_10641,N_9095,N_9533);
or U10642 (N_10642,N_10469,N_9190);
nand U10643 (N_10643,N_9446,N_9420);
or U10644 (N_10644,N_9819,N_9659);
or U10645 (N_10645,N_10014,N_9645);
or U10646 (N_10646,N_9945,N_10280);
nor U10647 (N_10647,N_10012,N_9683);
and U10648 (N_10648,N_9319,N_10201);
nand U10649 (N_10649,N_10088,N_9108);
nor U10650 (N_10650,N_9225,N_9751);
and U10651 (N_10651,N_9833,N_9291);
nand U10652 (N_10652,N_9169,N_10227);
nor U10653 (N_10653,N_9702,N_9059);
and U10654 (N_10654,N_9132,N_9542);
or U10655 (N_10655,N_9289,N_9753);
or U10656 (N_10656,N_9170,N_9716);
or U10657 (N_10657,N_10100,N_10215);
nor U10658 (N_10658,N_10033,N_9843);
nor U10659 (N_10659,N_9462,N_9733);
nor U10660 (N_10660,N_9579,N_10247);
nand U10661 (N_10661,N_10036,N_9179);
or U10662 (N_10662,N_10113,N_10055);
nand U10663 (N_10663,N_9187,N_9193);
nor U10664 (N_10664,N_9158,N_9532);
or U10665 (N_10665,N_10429,N_9817);
nand U10666 (N_10666,N_9075,N_9849);
and U10667 (N_10667,N_10270,N_9260);
and U10668 (N_10668,N_9497,N_9762);
and U10669 (N_10669,N_9977,N_10491);
and U10670 (N_10670,N_9787,N_9128);
nand U10671 (N_10671,N_10212,N_9441);
nor U10672 (N_10672,N_10190,N_10019);
nand U10673 (N_10673,N_10312,N_9486);
nand U10674 (N_10674,N_10299,N_10392);
or U10675 (N_10675,N_9353,N_10272);
nor U10676 (N_10676,N_10248,N_10114);
or U10677 (N_10677,N_10016,N_9424);
and U10678 (N_10678,N_9135,N_9451);
xnor U10679 (N_10679,N_10072,N_9707);
nand U10680 (N_10680,N_9100,N_9991);
or U10681 (N_10681,N_10307,N_10406);
and U10682 (N_10682,N_10470,N_9350);
and U10683 (N_10683,N_10283,N_9091);
or U10684 (N_10684,N_10123,N_9509);
nand U10685 (N_10685,N_10085,N_10147);
or U10686 (N_10686,N_10380,N_9926);
or U10687 (N_10687,N_9752,N_10034);
nor U10688 (N_10688,N_10287,N_9582);
nand U10689 (N_10689,N_9310,N_10244);
xor U10690 (N_10690,N_10242,N_9906);
or U10691 (N_10691,N_9073,N_10075);
xnor U10692 (N_10692,N_10330,N_10347);
or U10693 (N_10693,N_10243,N_9650);
or U10694 (N_10694,N_9885,N_10379);
or U10695 (N_10695,N_9379,N_10475);
nor U10696 (N_10696,N_9188,N_10276);
and U10697 (N_10697,N_10471,N_9140);
or U10698 (N_10698,N_10297,N_10208);
or U10699 (N_10699,N_10162,N_9842);
or U10700 (N_10700,N_9901,N_10040);
nor U10701 (N_10701,N_10472,N_10158);
or U10702 (N_10702,N_9457,N_9514);
nand U10703 (N_10703,N_10128,N_10200);
nor U10704 (N_10704,N_9498,N_10286);
and U10705 (N_10705,N_9670,N_9633);
or U10706 (N_10706,N_10204,N_9155);
or U10707 (N_10707,N_9781,N_9057);
and U10708 (N_10708,N_10175,N_9275);
or U10709 (N_10709,N_9832,N_10397);
or U10710 (N_10710,N_9658,N_9403);
and U10711 (N_10711,N_10388,N_9782);
nand U10712 (N_10712,N_10446,N_9105);
nor U10713 (N_10713,N_9834,N_9101);
and U10714 (N_10714,N_9411,N_9929);
nor U10715 (N_10715,N_10077,N_10418);
or U10716 (N_10716,N_10117,N_9773);
or U10717 (N_10717,N_9226,N_9149);
and U10718 (N_10718,N_10161,N_9984);
or U10719 (N_10719,N_9110,N_9150);
nand U10720 (N_10720,N_9211,N_9589);
or U10721 (N_10721,N_9668,N_9082);
nand U10722 (N_10722,N_10426,N_9470);
nand U10723 (N_10723,N_9587,N_9327);
nand U10724 (N_10724,N_9779,N_9956);
nand U10725 (N_10725,N_9571,N_9546);
nand U10726 (N_10726,N_9409,N_9458);
nand U10727 (N_10727,N_10156,N_9518);
and U10728 (N_10728,N_10044,N_10357);
or U10729 (N_10729,N_10344,N_9765);
or U10730 (N_10730,N_10024,N_9472);
nor U10731 (N_10731,N_10411,N_10425);
nor U10732 (N_10732,N_10401,N_9666);
or U10733 (N_10733,N_10002,N_10367);
and U10734 (N_10734,N_10432,N_10037);
nor U10735 (N_10735,N_9595,N_9143);
and U10736 (N_10736,N_9195,N_9181);
and U10737 (N_10737,N_9242,N_9616);
or U10738 (N_10738,N_10494,N_10474);
or U10739 (N_10739,N_9268,N_9679);
nand U10740 (N_10740,N_9034,N_9259);
or U10741 (N_10741,N_10387,N_10328);
nand U10742 (N_10742,N_10004,N_9256);
nor U10743 (N_10743,N_9878,N_10070);
nand U10744 (N_10744,N_10294,N_9895);
nor U10745 (N_10745,N_9723,N_9970);
or U10746 (N_10746,N_10051,N_9176);
or U10747 (N_10747,N_10370,N_9697);
nand U10748 (N_10748,N_10107,N_9427);
nand U10749 (N_10749,N_9689,N_9966);
nand U10750 (N_10750,N_10371,N_9406);
and U10751 (N_10751,N_9641,N_9736);
and U10752 (N_10752,N_10116,N_10188);
nor U10753 (N_10753,N_10144,N_9814);
or U10754 (N_10754,N_9943,N_9593);
nand U10755 (N_10755,N_9085,N_10336);
xor U10756 (N_10756,N_9717,N_9206);
xnor U10757 (N_10757,N_9250,N_9037);
nand U10758 (N_10758,N_10449,N_9807);
nand U10759 (N_10759,N_10073,N_9696);
and U10760 (N_10760,N_10434,N_10031);
or U10761 (N_10761,N_9300,N_9254);
nand U10762 (N_10762,N_9309,N_9512);
nor U10763 (N_10763,N_9157,N_9663);
and U10764 (N_10764,N_10281,N_10329);
and U10765 (N_10765,N_10155,N_9996);
or U10766 (N_10766,N_9489,N_10277);
and U10767 (N_10767,N_10216,N_9362);
and U10768 (N_10768,N_10020,N_10490);
nor U10769 (N_10769,N_10124,N_9163);
or U10770 (N_10770,N_9315,N_9046);
nor U10771 (N_10771,N_10393,N_10298);
nor U10772 (N_10772,N_9086,N_9501);
and U10773 (N_10773,N_9010,N_9431);
nand U10774 (N_10774,N_9502,N_9635);
nand U10775 (N_10775,N_10065,N_9063);
nand U10776 (N_10776,N_9672,N_10146);
and U10777 (N_10777,N_10390,N_9719);
and U10778 (N_10778,N_10028,N_9359);
or U10779 (N_10779,N_9099,N_10381);
nor U10780 (N_10780,N_10210,N_9644);
and U10781 (N_10781,N_10068,N_9989);
or U10782 (N_10782,N_9708,N_9675);
and U10783 (N_10783,N_9372,N_10206);
or U10784 (N_10784,N_10140,N_9264);
and U10785 (N_10785,N_9596,N_10332);
and U10786 (N_10786,N_9339,N_10364);
and U10787 (N_10787,N_10340,N_10050);
or U10788 (N_10788,N_9285,N_10318);
nor U10789 (N_10789,N_10081,N_9664);
nor U10790 (N_10790,N_9876,N_9045);
and U10791 (N_10791,N_10480,N_9488);
nor U10792 (N_10792,N_10399,N_9102);
or U10793 (N_10793,N_9443,N_9918);
and U10794 (N_10794,N_9134,N_9177);
nor U10795 (N_10795,N_9077,N_9153);
nand U10796 (N_10796,N_10032,N_9872);
and U10797 (N_10797,N_9585,N_9080);
and U10798 (N_10798,N_9393,N_9890);
or U10799 (N_10799,N_9069,N_10093);
nor U10800 (N_10800,N_9591,N_9550);
or U10801 (N_10801,N_10126,N_9643);
nor U10802 (N_10802,N_9611,N_9534);
or U10803 (N_10803,N_9031,N_9825);
or U10804 (N_10804,N_9463,N_10327);
nor U10805 (N_10805,N_9798,N_9931);
nand U10806 (N_10806,N_10245,N_9620);
nand U10807 (N_10807,N_10120,N_10207);
nand U10808 (N_10808,N_10409,N_10414);
and U10809 (N_10809,N_10198,N_10178);
nor U10810 (N_10810,N_9419,N_9348);
nor U10811 (N_10811,N_9119,N_9937);
nor U10812 (N_10812,N_9954,N_9005);
nand U10813 (N_10813,N_9043,N_10455);
nand U10814 (N_10814,N_9325,N_9007);
nor U10815 (N_10815,N_9160,N_9936);
and U10816 (N_10816,N_10150,N_9576);
or U10817 (N_10817,N_10302,N_9106);
nand U10818 (N_10818,N_10377,N_9854);
or U10819 (N_10819,N_10022,N_9425);
nand U10820 (N_10820,N_9882,N_9855);
and U10821 (N_10821,N_9262,N_10315);
and U10822 (N_10822,N_10009,N_9673);
and U10823 (N_10823,N_9328,N_9317);
nand U10824 (N_10824,N_10129,N_9900);
nor U10825 (N_10825,N_10087,N_9400);
or U10826 (N_10826,N_9897,N_10499);
and U10827 (N_10827,N_9543,N_9241);
nor U10828 (N_10828,N_10171,N_9232);
nand U10829 (N_10829,N_9469,N_9851);
and U10830 (N_10830,N_9346,N_9797);
and U10831 (N_10831,N_9418,N_9087);
nor U10832 (N_10832,N_9680,N_9314);
nand U10833 (N_10833,N_9415,N_9599);
and U10834 (N_10834,N_9840,N_9884);
and U10835 (N_10835,N_9536,N_9764);
nand U10836 (N_10836,N_10376,N_9642);
nand U10837 (N_10837,N_9939,N_10440);
nand U10838 (N_10838,N_10013,N_9092);
nor U10839 (N_10839,N_9661,N_9614);
nand U10840 (N_10840,N_10282,N_9304);
nor U10841 (N_10841,N_9528,N_9896);
or U10842 (N_10842,N_10448,N_9569);
nor U10843 (N_10843,N_9748,N_9600);
nor U10844 (N_10844,N_10052,N_10006);
and U10845 (N_10845,N_9266,N_9568);
and U10846 (N_10846,N_10258,N_9714);
nor U10847 (N_10847,N_9623,N_9508);
or U10848 (N_10848,N_9381,N_9358);
and U10849 (N_10849,N_9866,N_9231);
nor U10850 (N_10850,N_9162,N_9584);
nand U10851 (N_10851,N_9207,N_9892);
nand U10852 (N_10852,N_9349,N_9009);
or U10853 (N_10853,N_10373,N_9577);
nor U10854 (N_10854,N_9335,N_10337);
nor U10855 (N_10855,N_10056,N_9802);
and U10856 (N_10856,N_9338,N_9772);
or U10857 (N_10857,N_9391,N_9167);
and U10858 (N_10858,N_9720,N_9811);
nor U10859 (N_10859,N_10363,N_9480);
nand U10860 (N_10860,N_9141,N_10358);
nand U10861 (N_10861,N_9992,N_9565);
nand U10862 (N_10862,N_9868,N_10424);
nand U10863 (N_10863,N_10064,N_9089);
or U10864 (N_10864,N_9535,N_10041);
nand U10865 (N_10865,N_10407,N_9541);
nor U10866 (N_10866,N_10122,N_9345);
nor U10867 (N_10867,N_9212,N_9027);
or U10868 (N_10868,N_9387,N_9261);
and U10869 (N_10869,N_9930,N_10182);
or U10870 (N_10870,N_9459,N_9062);
and U10871 (N_10871,N_9744,N_9789);
nand U10872 (N_10872,N_9097,N_9513);
nand U10873 (N_10873,N_10412,N_10359);
and U10874 (N_10874,N_9307,N_9726);
nand U10875 (N_10875,N_10301,N_10195);
or U10876 (N_10876,N_10209,N_9793);
and U10877 (N_10877,N_9985,N_9410);
nor U10878 (N_10878,N_10430,N_9873);
or U10879 (N_10879,N_9656,N_9380);
nor U10880 (N_10880,N_9125,N_9066);
nor U10881 (N_10881,N_9405,N_10305);
nand U10882 (N_10882,N_9537,N_9084);
nor U10883 (N_10883,N_9677,N_9144);
and U10884 (N_10884,N_9312,N_9607);
or U10885 (N_10885,N_9399,N_10423);
and U10886 (N_10886,N_9742,N_9847);
nor U10887 (N_10887,N_9621,N_9574);
and U10888 (N_10888,N_9860,N_9279);
and U10889 (N_10889,N_9695,N_9864);
and U10890 (N_10890,N_9709,N_9692);
and U10891 (N_10891,N_10167,N_9539);
and U10892 (N_10892,N_9522,N_10484);
and U10893 (N_10893,N_9822,N_10354);
and U10894 (N_10894,N_9178,N_10460);
and U10895 (N_10895,N_9495,N_9021);
nor U10896 (N_10896,N_9561,N_9433);
and U10897 (N_10897,N_10110,N_10132);
nand U10898 (N_10898,N_10289,N_9191);
nand U10899 (N_10899,N_9961,N_9551);
nor U10900 (N_10900,N_9549,N_9356);
and U10901 (N_10901,N_10464,N_10157);
and U10902 (N_10902,N_9728,N_9968);
nor U10903 (N_10903,N_9761,N_9039);
or U10904 (N_10904,N_9388,N_9988);
and U10905 (N_10905,N_10378,N_10476);
or U10906 (N_10906,N_10095,N_10053);
or U10907 (N_10907,N_9559,N_9725);
nand U10908 (N_10908,N_9374,N_10148);
and U10909 (N_10909,N_9870,N_9915);
nor U10910 (N_10910,N_9547,N_9222);
nor U10911 (N_10911,N_10352,N_9515);
and U10912 (N_10912,N_9919,N_9363);
nand U10913 (N_10913,N_10317,N_9898);
nand U10914 (N_10914,N_10458,N_10109);
nand U10915 (N_10915,N_10486,N_10145);
nand U10916 (N_10916,N_9464,N_10279);
or U10917 (N_10917,N_9783,N_10439);
and U10918 (N_10918,N_9567,N_10421);
nor U10919 (N_10919,N_9686,N_9647);
and U10920 (N_10920,N_10232,N_10005);
or U10921 (N_10921,N_9479,N_9562);
nor U10922 (N_10922,N_9867,N_10482);
nand U10923 (N_10923,N_9688,N_9601);
and U10924 (N_10924,N_10125,N_9739);
nor U10925 (N_10925,N_9004,N_9492);
nor U10926 (N_10926,N_10436,N_9016);
nor U10927 (N_10927,N_9258,N_10320);
and U10928 (N_10928,N_9025,N_10026);
or U10929 (N_10929,N_9794,N_9578);
nor U10930 (N_10930,N_10442,N_9118);
nor U10931 (N_10931,N_9355,N_9058);
nor U10932 (N_10932,N_10071,N_9625);
nand U10933 (N_10933,N_10366,N_9452);
or U10934 (N_10934,N_9096,N_9159);
nor U10935 (N_10935,N_10092,N_10431);
nand U10936 (N_10936,N_9282,N_10463);
nor U10937 (N_10937,N_9450,N_9033);
nand U10938 (N_10938,N_10181,N_9776);
nor U10939 (N_10939,N_10027,N_9757);
nand U10940 (N_10940,N_9145,N_9439);
nor U10941 (N_10941,N_9088,N_9920);
or U10942 (N_10942,N_9775,N_10419);
and U10943 (N_10943,N_9653,N_10224);
nand U10944 (N_10944,N_10383,N_9941);
and U10945 (N_10945,N_9367,N_9831);
nand U10946 (N_10946,N_9997,N_10049);
nand U10947 (N_10947,N_9361,N_9301);
nor U10948 (N_10948,N_9051,N_9969);
or U10949 (N_10949,N_10141,N_10010);
nor U10950 (N_10950,N_9521,N_9235);
or U10951 (N_10951,N_10495,N_9654);
or U10952 (N_10952,N_9705,N_9008);
or U10953 (N_10953,N_9507,N_10391);
and U10954 (N_10954,N_10172,N_9566);
or U10955 (N_10955,N_9612,N_10351);
and U10956 (N_10956,N_9875,N_9510);
nand U10957 (N_10957,N_9448,N_9049);
nor U10958 (N_10958,N_9219,N_10000);
or U10959 (N_10959,N_9011,N_9548);
or U10960 (N_10960,N_9164,N_9044);
or U10961 (N_10961,N_9820,N_10334);
nor U10962 (N_10962,N_10236,N_9061);
or U10963 (N_10963,N_10295,N_10205);
and U10964 (N_10964,N_9848,N_9715);
nand U10965 (N_10965,N_9951,N_9921);
nand U10966 (N_10966,N_10345,N_9657);
nor U10967 (N_10967,N_10233,N_10222);
and U10968 (N_10968,N_9652,N_9604);
and U10969 (N_10969,N_9116,N_10285);
or U10970 (N_10970,N_9029,N_9669);
nor U10971 (N_10971,N_9272,N_10478);
or U10972 (N_10972,N_9563,N_9947);
nor U10973 (N_10973,N_9001,N_9979);
and U10974 (N_10974,N_9270,N_10214);
nand U10975 (N_10975,N_9681,N_9098);
nor U10976 (N_10976,N_9208,N_9429);
and U10977 (N_10977,N_10184,N_9000);
or U10978 (N_10978,N_10382,N_9127);
nor U10979 (N_10979,N_9466,N_9922);
and U10980 (N_10980,N_9972,N_9013);
nand U10981 (N_10981,N_9465,N_10457);
nand U10982 (N_10982,N_9710,N_9586);
nor U10983 (N_10983,N_9395,N_9925);
nand U10984 (N_10984,N_9210,N_9180);
and U10985 (N_10985,N_10433,N_9785);
nand U10986 (N_10986,N_9014,N_10203);
nand U10987 (N_10987,N_10121,N_10074);
nor U10988 (N_10988,N_10234,N_9287);
nand U10989 (N_10989,N_9800,N_9354);
or U10990 (N_10990,N_9438,N_10118);
nand U10991 (N_10991,N_10444,N_9402);
or U10992 (N_10992,N_9295,N_10135);
nor U10993 (N_10993,N_9198,N_10384);
or U10994 (N_10994,N_9036,N_9759);
nand U10995 (N_10995,N_10089,N_9240);
nor U10996 (N_10996,N_9904,N_9530);
or U10997 (N_10997,N_9394,N_9401);
or U10998 (N_10998,N_10160,N_9962);
nand U10999 (N_10999,N_10265,N_9126);
nand U11000 (N_11000,N_9417,N_9740);
nand U11001 (N_11001,N_10017,N_9908);
xor U11002 (N_11002,N_9124,N_9343);
and U11003 (N_11003,N_9881,N_9074);
nand U11004 (N_11004,N_9928,N_9022);
nand U11005 (N_11005,N_9383,N_10180);
nand U11006 (N_11006,N_9888,N_9869);
nor U11007 (N_11007,N_10079,N_10322);
xnor U11008 (N_11008,N_9630,N_9893);
or U11009 (N_11009,N_9369,N_9646);
nor U11010 (N_11010,N_9165,N_9853);
nand U11011 (N_11011,N_9204,N_10372);
nand U11012 (N_11012,N_10228,N_10001);
xor U11013 (N_11013,N_10130,N_10408);
or U11014 (N_11014,N_10261,N_9366);
or U11015 (N_11015,N_10416,N_10253);
and U11016 (N_11016,N_10300,N_9627);
nor U11017 (N_11017,N_10349,N_9552);
nand U11018 (N_11018,N_10030,N_9712);
and U11019 (N_11019,N_9104,N_9475);
nor U11020 (N_11020,N_9248,N_9189);
xnor U11021 (N_11021,N_10246,N_10403);
and U11022 (N_11022,N_10223,N_9662);
nand U11023 (N_11023,N_9687,N_9070);
and U11024 (N_11024,N_10196,N_9422);
nand U11025 (N_11025,N_9932,N_9371);
nor U11026 (N_11026,N_9306,N_9770);
nand U11027 (N_11027,N_9805,N_9605);
nand U11028 (N_11028,N_9727,N_10492);
nor U11029 (N_11029,N_9265,N_10023);
or U11030 (N_11030,N_9389,N_9755);
nand U11031 (N_11031,N_9856,N_10477);
xor U11032 (N_11032,N_9483,N_9390);
and U11033 (N_11033,N_10395,N_10356);
and U11034 (N_11034,N_9963,N_9437);
nor U11035 (N_11035,N_10179,N_10291);
nor U11036 (N_11036,N_9018,N_9699);
nor U11037 (N_11037,N_9671,N_10083);
and U11038 (N_11038,N_9283,N_9575);
or U11039 (N_11039,N_10443,N_10211);
and U11040 (N_11040,N_10360,N_9230);
and U11041 (N_11041,N_9691,N_9115);
nand U11042 (N_11042,N_10143,N_10060);
or U11043 (N_11043,N_10316,N_9166);
nand U11044 (N_11044,N_10082,N_10341);
nand U11045 (N_11045,N_9286,N_9130);
nor U11046 (N_11046,N_9064,N_9467);
and U11047 (N_11047,N_9818,N_9940);
nor U11048 (N_11048,N_9933,N_10185);
or U11049 (N_11049,N_10428,N_10165);
or U11050 (N_11050,N_9990,N_9269);
or U11051 (N_11051,N_9701,N_10176);
or U11052 (N_11052,N_9333,N_10168);
and U11053 (N_11053,N_9729,N_9368);
and U11054 (N_11054,N_9280,N_10217);
nor U11055 (N_11055,N_10374,N_9859);
and U11056 (N_11056,N_10189,N_9373);
and U11057 (N_11057,N_10096,N_9175);
or U11058 (N_11058,N_9094,N_9592);
and U11059 (N_11059,N_9674,N_10127);
nand U11060 (N_11060,N_10059,N_10108);
nor U11061 (N_11061,N_10149,N_9078);
or U11062 (N_11062,N_10375,N_9090);
or U11063 (N_11063,N_10398,N_9015);
or U11064 (N_11064,N_9003,N_10103);
and U11065 (N_11065,N_10218,N_9040);
and U11066 (N_11066,N_10309,N_10134);
and U11067 (N_11067,N_10187,N_9223);
nand U11068 (N_11068,N_10292,N_10306);
or U11069 (N_11069,N_9731,N_9902);
nor U11070 (N_11070,N_10240,N_9801);
or U11071 (N_11071,N_9766,N_9655);
or U11072 (N_11072,N_9590,N_9277);
and U11073 (N_11073,N_9795,N_9622);
or U11074 (N_11074,N_10368,N_9857);
and U11075 (N_11075,N_9288,N_9205);
or U11076 (N_11076,N_9432,N_9136);
or U11077 (N_11077,N_9803,N_9026);
nand U11078 (N_11078,N_10112,N_9257);
and U11079 (N_11079,N_10220,N_9267);
nand U11080 (N_11080,N_9850,N_10018);
nor U11081 (N_11081,N_9331,N_9845);
nor U11082 (N_11082,N_10011,N_10238);
nor U11083 (N_11083,N_10400,N_9706);
nand U11084 (N_11084,N_9196,N_9768);
nor U11085 (N_11085,N_9628,N_9516);
nor U11086 (N_11086,N_9184,N_10164);
nor U11087 (N_11087,N_10235,N_9447);
or U11088 (N_11088,N_9234,N_10296);
and U11089 (N_11089,N_9493,N_10447);
and U11090 (N_11090,N_10219,N_10099);
or U11091 (N_11091,N_10338,N_10257);
or U11092 (N_11092,N_9829,N_10497);
and U11093 (N_11093,N_9987,N_9020);
and U11094 (N_11094,N_9217,N_10361);
or U11095 (N_11095,N_9002,N_10275);
or U11096 (N_11096,N_9378,N_10076);
or U11097 (N_11097,N_9271,N_9986);
nor U11098 (N_11098,N_10323,N_9142);
nor U11099 (N_11099,N_10063,N_10249);
nand U11100 (N_11100,N_9273,N_9375);
nor U11101 (N_11101,N_10259,N_9780);
nand U11102 (N_11102,N_9721,N_9274);
nand U11103 (N_11103,N_9750,N_9749);
or U11104 (N_11104,N_9500,N_9434);
nor U11105 (N_11105,N_9056,N_9730);
nor U11106 (N_11106,N_9959,N_9397);
nor U11107 (N_11107,N_9626,N_10091);
nand U11108 (N_11108,N_9786,N_9496);
nand U11109 (N_11109,N_9213,N_9743);
nor U11110 (N_11110,N_9916,N_10461);
or U11111 (N_11111,N_9934,N_9093);
or U11112 (N_11112,N_9482,N_9517);
and U11113 (N_11113,N_9948,N_9676);
nand U11114 (N_11114,N_9168,N_10069);
nor U11115 (N_11115,N_9771,N_10313);
and U11116 (N_11116,N_9554,N_9197);
and U11117 (N_11117,N_9174,N_10365);
nand U11118 (N_11118,N_9700,N_10191);
and U11119 (N_11119,N_9428,N_9852);
nor U11120 (N_11120,N_10003,N_9894);
nand U11121 (N_11121,N_10269,N_9079);
nand U11122 (N_11122,N_9111,N_9606);
and U11123 (N_11123,N_9255,N_9880);
nor U11124 (N_11124,N_9245,N_10131);
and U11125 (N_11125,N_10451,N_9841);
nor U11126 (N_11126,N_9746,N_10078);
or U11127 (N_11127,N_10355,N_9120);
xnor U11128 (N_11128,N_9050,N_9490);
nand U11129 (N_11129,N_9995,N_9792);
or U11130 (N_11130,N_10402,N_9065);
nand U11131 (N_11131,N_10267,N_9813);
or U11132 (N_11132,N_9558,N_10405);
or U11133 (N_11133,N_9796,N_10467);
or U11134 (N_11134,N_9994,N_9484);
nand U11135 (N_11135,N_9436,N_9526);
and U11136 (N_11136,N_9520,N_9147);
and U11137 (N_11137,N_10369,N_10137);
nor U11138 (N_11138,N_9863,N_9347);
nand U11139 (N_11139,N_9874,N_9032);
and U11140 (N_11140,N_9660,N_9171);
and U11141 (N_11141,N_9398,N_10496);
and U11142 (N_11142,N_10166,N_9523);
nand U11143 (N_11143,N_9028,N_9540);
nand U11144 (N_11144,N_9214,N_9837);
and U11145 (N_11145,N_9861,N_9423);
or U11146 (N_11146,N_10335,N_9911);
and U11147 (N_11147,N_9053,N_10057);
and U11148 (N_11148,N_9377,N_9421);
nor U11149 (N_11149,N_9665,N_10152);
nand U11150 (N_11150,N_9233,N_9278);
and U11151 (N_11151,N_10177,N_10362);
or U11152 (N_11152,N_9370,N_10481);
nor U11153 (N_11153,N_10346,N_9216);
nor U11154 (N_11154,N_9758,N_9952);
nor U11155 (N_11155,N_10319,N_9912);
xnor U11156 (N_11156,N_9060,N_10102);
nor U11157 (N_11157,N_9076,N_10303);
or U11158 (N_11158,N_9471,N_9886);
nor U11159 (N_11159,N_10111,N_10326);
and U11160 (N_11160,N_9430,N_9907);
nand U11161 (N_11161,N_9445,N_9048);
nand U11162 (N_11162,N_9603,N_9340);
or U11163 (N_11163,N_9201,N_10193);
or U11164 (N_11164,N_9735,N_9553);
nor U11165 (N_11165,N_9976,N_9444);
nand U11166 (N_11166,N_10163,N_10213);
nor U11167 (N_11167,N_9012,N_10308);
nand U11168 (N_11168,N_10445,N_10410);
nor U11169 (N_11169,N_10046,N_10485);
nand U11170 (N_11170,N_9588,N_9290);
nand U11171 (N_11171,N_10255,N_10252);
nand U11172 (N_11172,N_9324,N_10142);
or U11173 (N_11173,N_9318,N_9505);
xor U11174 (N_11174,N_9678,N_10066);
xnor U11175 (N_11175,N_9435,N_9042);
or U11176 (N_11176,N_9790,N_9185);
nand U11177 (N_11177,N_9316,N_9718);
nor U11178 (N_11178,N_9909,N_9778);
or U11179 (N_11179,N_9236,N_9308);
or U11180 (N_11180,N_9052,N_9519);
and U11181 (N_11181,N_9570,N_9555);
nand U11182 (N_11182,N_10290,N_9763);
or U11183 (N_11183,N_9914,N_10139);
nor U11184 (N_11184,N_9905,N_10154);
nor U11185 (N_11185,N_9313,N_9738);
nor U11186 (N_11186,N_10489,N_9414);
and U11187 (N_11187,N_9799,N_9341);
nor U11188 (N_11188,N_9461,N_9440);
and U11189 (N_11189,N_9154,N_9754);
nand U11190 (N_11190,N_9114,N_10174);
or U11191 (N_11191,N_9109,N_9924);
or U11192 (N_11192,N_10273,N_10151);
and U11193 (N_11193,N_9804,N_9192);
or U11194 (N_11194,N_9474,N_10284);
and U11195 (N_11195,N_9637,N_9784);
and U11196 (N_11196,N_9618,N_9329);
nand U11197 (N_11197,N_9129,N_10415);
or U11198 (N_11198,N_9704,N_9017);
nand U11199 (N_11199,N_10331,N_9511);
nand U11200 (N_11200,N_9722,N_9321);
nand U11201 (N_11201,N_10173,N_9122);
nand U11202 (N_11202,N_10169,N_9583);
or U11203 (N_11203,N_9203,N_9835);
nand U11204 (N_11204,N_10339,N_10404);
nand U11205 (N_11205,N_9404,N_10115);
nor U11206 (N_11206,N_9609,N_9615);
xor U11207 (N_11207,N_10350,N_10456);
nor U11208 (N_11208,N_9879,N_9950);
nand U11209 (N_11209,N_9734,N_9209);
and U11210 (N_11210,N_9826,N_10048);
and U11211 (N_11211,N_10427,N_10385);
nand U11212 (N_11212,N_9651,N_10454);
nor U11213 (N_11213,N_9824,N_10097);
and U11214 (N_11214,N_9138,N_10231);
or U11215 (N_11215,N_9836,N_9788);
and U11216 (N_11216,N_9186,N_10343);
or U11217 (N_11217,N_9649,N_9247);
or U11218 (N_11218,N_9249,N_10237);
and U11219 (N_11219,N_9949,N_10437);
nand U11220 (N_11220,N_9476,N_9227);
and U11221 (N_11221,N_10170,N_9137);
nand U11222 (N_11222,N_9777,N_9903);
nand U11223 (N_11223,N_9927,N_9741);
nor U11224 (N_11224,N_10062,N_9634);
nand U11225 (N_11225,N_9068,N_10304);
and U11226 (N_11226,N_10058,N_9524);
or U11227 (N_11227,N_10311,N_10386);
nand U11228 (N_11228,N_9967,N_9146);
or U11229 (N_11229,N_10015,N_10080);
and U11230 (N_11230,N_9910,N_9202);
and U11231 (N_11231,N_10186,N_9923);
nor U11232 (N_11232,N_10263,N_10047);
or U11233 (N_11233,N_9481,N_10473);
or U11234 (N_11234,N_9019,N_9426);
or U11235 (N_11235,N_10101,N_9413);
nor U11236 (N_11236,N_9823,N_9506);
xor U11237 (N_11237,N_9965,N_9229);
or U11238 (N_11238,N_9975,N_9396);
or U11239 (N_11239,N_9252,N_9182);
nand U11240 (N_11240,N_9745,N_9883);
and U11241 (N_11241,N_9598,N_9494);
or U11242 (N_11242,N_9747,N_9342);
and U11243 (N_11243,N_10420,N_9808);
or U11244 (N_11244,N_10239,N_9917);
and U11245 (N_11245,N_10086,N_9557);
or U11246 (N_11246,N_9294,N_9172);
or U11247 (N_11247,N_9816,N_10479);
nor U11248 (N_11248,N_10389,N_9030);
nand U11249 (N_11249,N_9041,N_9220);
and U11250 (N_11250,N_9659,N_9317);
or U11251 (N_11251,N_9491,N_10336);
nor U11252 (N_11252,N_9562,N_9773);
nand U11253 (N_11253,N_9749,N_10236);
or U11254 (N_11254,N_10052,N_9345);
or U11255 (N_11255,N_10224,N_10048);
nor U11256 (N_11256,N_9060,N_9579);
nor U11257 (N_11257,N_10026,N_9002);
nand U11258 (N_11258,N_10308,N_9569);
nor U11259 (N_11259,N_10359,N_9993);
and U11260 (N_11260,N_9202,N_10037);
and U11261 (N_11261,N_10393,N_9941);
and U11262 (N_11262,N_9868,N_10177);
nand U11263 (N_11263,N_9198,N_9528);
or U11264 (N_11264,N_9072,N_9833);
xor U11265 (N_11265,N_9719,N_9237);
nand U11266 (N_11266,N_9705,N_10188);
nor U11267 (N_11267,N_9765,N_9095);
or U11268 (N_11268,N_9123,N_9498);
or U11269 (N_11269,N_10217,N_10012);
nor U11270 (N_11270,N_9261,N_9775);
or U11271 (N_11271,N_9885,N_10271);
nor U11272 (N_11272,N_10330,N_9401);
and U11273 (N_11273,N_9528,N_9639);
and U11274 (N_11274,N_9418,N_9148);
or U11275 (N_11275,N_9468,N_10249);
nor U11276 (N_11276,N_9669,N_9526);
nand U11277 (N_11277,N_9018,N_9767);
nor U11278 (N_11278,N_10119,N_9353);
or U11279 (N_11279,N_10474,N_10265);
or U11280 (N_11280,N_9310,N_9329);
and U11281 (N_11281,N_9612,N_9282);
or U11282 (N_11282,N_10368,N_9184);
nand U11283 (N_11283,N_9613,N_9873);
nor U11284 (N_11284,N_10306,N_9070);
or U11285 (N_11285,N_9564,N_9789);
nand U11286 (N_11286,N_9098,N_9192);
and U11287 (N_11287,N_9504,N_9962);
or U11288 (N_11288,N_9089,N_9502);
or U11289 (N_11289,N_10488,N_10176);
nand U11290 (N_11290,N_10213,N_9352);
xnor U11291 (N_11291,N_9598,N_9017);
or U11292 (N_11292,N_9988,N_10297);
and U11293 (N_11293,N_9598,N_9094);
and U11294 (N_11294,N_10403,N_10173);
nor U11295 (N_11295,N_9463,N_9755);
or U11296 (N_11296,N_10488,N_10319);
and U11297 (N_11297,N_9252,N_9351);
or U11298 (N_11298,N_9323,N_9184);
or U11299 (N_11299,N_10447,N_9874);
and U11300 (N_11300,N_9617,N_9670);
or U11301 (N_11301,N_9896,N_10384);
nand U11302 (N_11302,N_9418,N_9600);
nand U11303 (N_11303,N_10064,N_10193);
or U11304 (N_11304,N_9805,N_9682);
xnor U11305 (N_11305,N_9806,N_9443);
and U11306 (N_11306,N_10024,N_10118);
xnor U11307 (N_11307,N_9712,N_9009);
nand U11308 (N_11308,N_9544,N_9535);
nor U11309 (N_11309,N_9043,N_10088);
nor U11310 (N_11310,N_9656,N_9322);
and U11311 (N_11311,N_10351,N_9918);
nand U11312 (N_11312,N_9029,N_9131);
nor U11313 (N_11313,N_10001,N_10215);
nor U11314 (N_11314,N_10436,N_9450);
nor U11315 (N_11315,N_10263,N_9425);
and U11316 (N_11316,N_9070,N_10326);
or U11317 (N_11317,N_9315,N_9001);
nor U11318 (N_11318,N_9857,N_10163);
or U11319 (N_11319,N_10313,N_10429);
nand U11320 (N_11320,N_9149,N_9050);
and U11321 (N_11321,N_9308,N_9462);
or U11322 (N_11322,N_9359,N_10042);
and U11323 (N_11323,N_10064,N_9816);
nand U11324 (N_11324,N_9687,N_10140);
nor U11325 (N_11325,N_9336,N_9303);
nor U11326 (N_11326,N_9438,N_10310);
nand U11327 (N_11327,N_9397,N_9968);
or U11328 (N_11328,N_10371,N_9535);
nand U11329 (N_11329,N_9614,N_9714);
nor U11330 (N_11330,N_9325,N_9953);
and U11331 (N_11331,N_9509,N_9694);
and U11332 (N_11332,N_9456,N_9132);
nand U11333 (N_11333,N_9073,N_10216);
and U11334 (N_11334,N_10443,N_9967);
nor U11335 (N_11335,N_9259,N_9035);
or U11336 (N_11336,N_9552,N_10212);
nor U11337 (N_11337,N_9462,N_9761);
nor U11338 (N_11338,N_9092,N_9181);
or U11339 (N_11339,N_10325,N_10212);
nor U11340 (N_11340,N_10364,N_9602);
or U11341 (N_11341,N_9609,N_9367);
and U11342 (N_11342,N_10289,N_10296);
and U11343 (N_11343,N_9849,N_9431);
or U11344 (N_11344,N_9284,N_10373);
or U11345 (N_11345,N_9322,N_10186);
and U11346 (N_11346,N_9015,N_10293);
nor U11347 (N_11347,N_10198,N_9691);
and U11348 (N_11348,N_9688,N_10292);
nor U11349 (N_11349,N_9730,N_10488);
nor U11350 (N_11350,N_9565,N_10150);
xnor U11351 (N_11351,N_10332,N_9586);
nand U11352 (N_11352,N_10054,N_9378);
nand U11353 (N_11353,N_9351,N_9954);
and U11354 (N_11354,N_9008,N_9707);
and U11355 (N_11355,N_9413,N_9547);
nand U11356 (N_11356,N_9273,N_9463);
and U11357 (N_11357,N_9560,N_9609);
xnor U11358 (N_11358,N_9366,N_9893);
nor U11359 (N_11359,N_10304,N_9534);
nand U11360 (N_11360,N_9286,N_9832);
or U11361 (N_11361,N_9565,N_9896);
nand U11362 (N_11362,N_9004,N_9129);
nor U11363 (N_11363,N_9188,N_9348);
nor U11364 (N_11364,N_9326,N_9373);
or U11365 (N_11365,N_9752,N_9281);
nand U11366 (N_11366,N_9122,N_9448);
and U11367 (N_11367,N_9997,N_10355);
nor U11368 (N_11368,N_9717,N_9964);
nand U11369 (N_11369,N_9618,N_9475);
nand U11370 (N_11370,N_9788,N_9605);
nor U11371 (N_11371,N_9214,N_10079);
nand U11372 (N_11372,N_9463,N_10444);
xnor U11373 (N_11373,N_9005,N_10319);
nand U11374 (N_11374,N_9445,N_9437);
nand U11375 (N_11375,N_10432,N_9660);
nor U11376 (N_11376,N_9924,N_10234);
or U11377 (N_11377,N_9934,N_9054);
nand U11378 (N_11378,N_9518,N_9574);
nand U11379 (N_11379,N_9247,N_9137);
and U11380 (N_11380,N_10243,N_9012);
nor U11381 (N_11381,N_9052,N_9198);
and U11382 (N_11382,N_9582,N_9649);
and U11383 (N_11383,N_9894,N_9314);
nor U11384 (N_11384,N_9294,N_10123);
nand U11385 (N_11385,N_10441,N_9705);
nor U11386 (N_11386,N_10226,N_10406);
nor U11387 (N_11387,N_9019,N_9201);
or U11388 (N_11388,N_9099,N_9233);
and U11389 (N_11389,N_9348,N_10294);
nor U11390 (N_11390,N_9749,N_9479);
and U11391 (N_11391,N_9663,N_10341);
and U11392 (N_11392,N_9371,N_10166);
nand U11393 (N_11393,N_10247,N_10266);
or U11394 (N_11394,N_10287,N_9492);
nor U11395 (N_11395,N_10075,N_9181);
and U11396 (N_11396,N_9191,N_9920);
and U11397 (N_11397,N_10154,N_9775);
nor U11398 (N_11398,N_10413,N_9166);
nand U11399 (N_11399,N_9580,N_9544);
and U11400 (N_11400,N_9889,N_9148);
nand U11401 (N_11401,N_9662,N_9725);
and U11402 (N_11402,N_10000,N_9125);
nand U11403 (N_11403,N_9087,N_9816);
or U11404 (N_11404,N_9301,N_10001);
nand U11405 (N_11405,N_9635,N_10461);
nand U11406 (N_11406,N_9961,N_9504);
nand U11407 (N_11407,N_9588,N_9903);
nand U11408 (N_11408,N_10270,N_9525);
nand U11409 (N_11409,N_9509,N_9150);
nor U11410 (N_11410,N_9426,N_10147);
or U11411 (N_11411,N_9293,N_9056);
nand U11412 (N_11412,N_9905,N_9999);
nand U11413 (N_11413,N_9220,N_10394);
and U11414 (N_11414,N_9506,N_10283);
and U11415 (N_11415,N_10052,N_10313);
nor U11416 (N_11416,N_9647,N_9654);
nor U11417 (N_11417,N_9448,N_9076);
and U11418 (N_11418,N_10285,N_10179);
nor U11419 (N_11419,N_9725,N_10170);
xor U11420 (N_11420,N_9842,N_9648);
and U11421 (N_11421,N_9455,N_9483);
or U11422 (N_11422,N_9933,N_9182);
or U11423 (N_11423,N_10141,N_9440);
or U11424 (N_11424,N_9217,N_9980);
nand U11425 (N_11425,N_9383,N_9048);
nand U11426 (N_11426,N_9484,N_9046);
nand U11427 (N_11427,N_9023,N_9179);
nor U11428 (N_11428,N_9225,N_9038);
or U11429 (N_11429,N_9588,N_9106);
nand U11430 (N_11430,N_10340,N_10293);
nor U11431 (N_11431,N_9169,N_10150);
nor U11432 (N_11432,N_9101,N_9822);
xor U11433 (N_11433,N_9767,N_10099);
nor U11434 (N_11434,N_9512,N_9667);
and U11435 (N_11435,N_10123,N_9170);
and U11436 (N_11436,N_9352,N_9330);
or U11437 (N_11437,N_10454,N_9370);
nand U11438 (N_11438,N_9424,N_9498);
nand U11439 (N_11439,N_9635,N_9019);
and U11440 (N_11440,N_10203,N_10310);
nor U11441 (N_11441,N_9186,N_10193);
and U11442 (N_11442,N_10417,N_9015);
nor U11443 (N_11443,N_9937,N_9712);
or U11444 (N_11444,N_9081,N_9910);
nand U11445 (N_11445,N_10446,N_9611);
and U11446 (N_11446,N_10109,N_10214);
nand U11447 (N_11447,N_10231,N_9492);
or U11448 (N_11448,N_9812,N_9322);
or U11449 (N_11449,N_10441,N_9476);
and U11450 (N_11450,N_9274,N_9799);
nand U11451 (N_11451,N_10176,N_9020);
or U11452 (N_11452,N_9402,N_9665);
or U11453 (N_11453,N_10080,N_9790);
nor U11454 (N_11454,N_10233,N_9466);
and U11455 (N_11455,N_9637,N_10142);
nor U11456 (N_11456,N_9081,N_10042);
and U11457 (N_11457,N_9508,N_9177);
nor U11458 (N_11458,N_9471,N_9871);
nor U11459 (N_11459,N_9963,N_9407);
nand U11460 (N_11460,N_10461,N_9315);
or U11461 (N_11461,N_10484,N_9217);
or U11462 (N_11462,N_10416,N_10231);
nor U11463 (N_11463,N_9966,N_9265);
nand U11464 (N_11464,N_9001,N_10234);
nand U11465 (N_11465,N_10000,N_10258);
nand U11466 (N_11466,N_9647,N_9814);
nor U11467 (N_11467,N_10343,N_9357);
nand U11468 (N_11468,N_9960,N_9187);
or U11469 (N_11469,N_9482,N_9366);
nand U11470 (N_11470,N_9255,N_10446);
nor U11471 (N_11471,N_10485,N_9750);
or U11472 (N_11472,N_9208,N_9057);
or U11473 (N_11473,N_9041,N_9259);
nor U11474 (N_11474,N_9107,N_9746);
nor U11475 (N_11475,N_9014,N_10460);
or U11476 (N_11476,N_9602,N_10069);
or U11477 (N_11477,N_9049,N_10216);
nor U11478 (N_11478,N_10253,N_10204);
nand U11479 (N_11479,N_9501,N_10158);
or U11480 (N_11480,N_10014,N_9328);
nor U11481 (N_11481,N_10116,N_10186);
or U11482 (N_11482,N_9717,N_10278);
nor U11483 (N_11483,N_9505,N_9799);
and U11484 (N_11484,N_10330,N_9140);
nand U11485 (N_11485,N_9978,N_9207);
nor U11486 (N_11486,N_10357,N_10438);
and U11487 (N_11487,N_9635,N_9067);
and U11488 (N_11488,N_9364,N_10330);
and U11489 (N_11489,N_9587,N_9507);
and U11490 (N_11490,N_10053,N_9062);
or U11491 (N_11491,N_9707,N_9375);
nor U11492 (N_11492,N_9598,N_9608);
nor U11493 (N_11493,N_9781,N_9873);
or U11494 (N_11494,N_10038,N_9525);
and U11495 (N_11495,N_9122,N_10147);
or U11496 (N_11496,N_10470,N_9773);
and U11497 (N_11497,N_9051,N_10464);
or U11498 (N_11498,N_9604,N_10449);
nor U11499 (N_11499,N_10371,N_9140);
or U11500 (N_11500,N_9781,N_10314);
or U11501 (N_11501,N_9339,N_9824);
or U11502 (N_11502,N_9013,N_10011);
nor U11503 (N_11503,N_9929,N_9887);
or U11504 (N_11504,N_10251,N_9133);
nand U11505 (N_11505,N_9830,N_9749);
or U11506 (N_11506,N_9760,N_9977);
nand U11507 (N_11507,N_10237,N_10115);
nand U11508 (N_11508,N_10189,N_10225);
nor U11509 (N_11509,N_9533,N_9425);
nor U11510 (N_11510,N_9747,N_10357);
or U11511 (N_11511,N_9328,N_9305);
nor U11512 (N_11512,N_10005,N_9060);
nor U11513 (N_11513,N_10186,N_9379);
or U11514 (N_11514,N_10133,N_9726);
nor U11515 (N_11515,N_9798,N_9032);
nor U11516 (N_11516,N_10031,N_10499);
nor U11517 (N_11517,N_9804,N_10172);
nand U11518 (N_11518,N_10147,N_9903);
and U11519 (N_11519,N_10153,N_9916);
nor U11520 (N_11520,N_9334,N_9659);
nand U11521 (N_11521,N_10099,N_9065);
nor U11522 (N_11522,N_10258,N_10246);
and U11523 (N_11523,N_9830,N_9589);
nor U11524 (N_11524,N_10430,N_9449);
or U11525 (N_11525,N_10153,N_9548);
nor U11526 (N_11526,N_10023,N_10039);
nor U11527 (N_11527,N_9695,N_9138);
and U11528 (N_11528,N_9426,N_10146);
nor U11529 (N_11529,N_10445,N_9403);
nand U11530 (N_11530,N_9092,N_10218);
nor U11531 (N_11531,N_10440,N_10406);
and U11532 (N_11532,N_9944,N_9831);
nand U11533 (N_11533,N_9342,N_9391);
and U11534 (N_11534,N_10105,N_9520);
nand U11535 (N_11535,N_10242,N_9962);
and U11536 (N_11536,N_9827,N_9824);
or U11537 (N_11537,N_10108,N_9057);
and U11538 (N_11538,N_9535,N_10000);
nor U11539 (N_11539,N_9785,N_9112);
or U11540 (N_11540,N_10439,N_9428);
and U11541 (N_11541,N_9256,N_9279);
nand U11542 (N_11542,N_10364,N_10252);
and U11543 (N_11543,N_10436,N_10246);
nor U11544 (N_11544,N_10017,N_9879);
nor U11545 (N_11545,N_10446,N_9340);
nor U11546 (N_11546,N_10027,N_10360);
nand U11547 (N_11547,N_10002,N_9083);
or U11548 (N_11548,N_9195,N_10192);
or U11549 (N_11549,N_9327,N_9357);
and U11550 (N_11550,N_9279,N_9028);
and U11551 (N_11551,N_10258,N_9121);
nor U11552 (N_11552,N_9441,N_9646);
nor U11553 (N_11553,N_9716,N_9551);
nand U11554 (N_11554,N_10416,N_10032);
nor U11555 (N_11555,N_10223,N_9770);
nor U11556 (N_11556,N_10352,N_9144);
or U11557 (N_11557,N_9436,N_9262);
or U11558 (N_11558,N_9419,N_9755);
or U11559 (N_11559,N_9546,N_9357);
nand U11560 (N_11560,N_10278,N_9326);
and U11561 (N_11561,N_10015,N_9666);
or U11562 (N_11562,N_9854,N_9592);
or U11563 (N_11563,N_10369,N_10053);
and U11564 (N_11564,N_10323,N_9563);
nand U11565 (N_11565,N_9288,N_9456);
and U11566 (N_11566,N_9842,N_10219);
nand U11567 (N_11567,N_9050,N_9211);
nand U11568 (N_11568,N_9832,N_9011);
nor U11569 (N_11569,N_10322,N_10404);
nor U11570 (N_11570,N_9920,N_9337);
and U11571 (N_11571,N_10235,N_10088);
nand U11572 (N_11572,N_9970,N_9069);
and U11573 (N_11573,N_9348,N_9624);
and U11574 (N_11574,N_9416,N_10009);
or U11575 (N_11575,N_9471,N_10233);
and U11576 (N_11576,N_9638,N_10341);
or U11577 (N_11577,N_9395,N_9086);
nor U11578 (N_11578,N_10079,N_9927);
and U11579 (N_11579,N_9832,N_10243);
or U11580 (N_11580,N_9077,N_9291);
nand U11581 (N_11581,N_9115,N_9802);
and U11582 (N_11582,N_9553,N_9524);
nand U11583 (N_11583,N_9961,N_9484);
or U11584 (N_11584,N_9689,N_9142);
or U11585 (N_11585,N_9050,N_10165);
nor U11586 (N_11586,N_9688,N_10031);
nand U11587 (N_11587,N_10263,N_9674);
nor U11588 (N_11588,N_9100,N_10209);
or U11589 (N_11589,N_10084,N_9488);
or U11590 (N_11590,N_9434,N_9082);
or U11591 (N_11591,N_10018,N_10104);
nand U11592 (N_11592,N_9228,N_9277);
nand U11593 (N_11593,N_9086,N_9242);
nor U11594 (N_11594,N_9324,N_10486);
or U11595 (N_11595,N_10369,N_10478);
or U11596 (N_11596,N_9006,N_10283);
nand U11597 (N_11597,N_9825,N_9634);
nor U11598 (N_11598,N_10002,N_9877);
nand U11599 (N_11599,N_10195,N_10108);
or U11600 (N_11600,N_9822,N_9390);
or U11601 (N_11601,N_9858,N_9273);
nor U11602 (N_11602,N_10394,N_9440);
nor U11603 (N_11603,N_10117,N_10212);
nand U11604 (N_11604,N_9554,N_9285);
or U11605 (N_11605,N_9366,N_9081);
or U11606 (N_11606,N_9401,N_9443);
or U11607 (N_11607,N_9521,N_9574);
and U11608 (N_11608,N_9436,N_9671);
nand U11609 (N_11609,N_9223,N_9883);
and U11610 (N_11610,N_9879,N_10327);
nand U11611 (N_11611,N_10346,N_9676);
and U11612 (N_11612,N_9514,N_9565);
and U11613 (N_11613,N_9480,N_10010);
and U11614 (N_11614,N_10376,N_9456);
nor U11615 (N_11615,N_9117,N_9374);
and U11616 (N_11616,N_10213,N_9156);
and U11617 (N_11617,N_9456,N_10229);
and U11618 (N_11618,N_9433,N_9195);
and U11619 (N_11619,N_9336,N_9664);
and U11620 (N_11620,N_10278,N_9237);
and U11621 (N_11621,N_9785,N_9252);
or U11622 (N_11622,N_9438,N_9165);
or U11623 (N_11623,N_10313,N_9030);
and U11624 (N_11624,N_9610,N_9981);
or U11625 (N_11625,N_10228,N_10112);
nand U11626 (N_11626,N_9351,N_10426);
and U11627 (N_11627,N_9575,N_9766);
or U11628 (N_11628,N_10109,N_9468);
nand U11629 (N_11629,N_9768,N_10103);
nand U11630 (N_11630,N_9691,N_10399);
nand U11631 (N_11631,N_10131,N_9469);
or U11632 (N_11632,N_9688,N_10300);
nor U11633 (N_11633,N_9331,N_9473);
nand U11634 (N_11634,N_9653,N_9060);
nand U11635 (N_11635,N_9118,N_10085);
and U11636 (N_11636,N_10038,N_10443);
and U11637 (N_11637,N_9734,N_9642);
nand U11638 (N_11638,N_9518,N_9720);
nor U11639 (N_11639,N_9601,N_9768);
nor U11640 (N_11640,N_10292,N_9247);
or U11641 (N_11641,N_9859,N_9658);
nor U11642 (N_11642,N_9106,N_9340);
nor U11643 (N_11643,N_10320,N_9810);
and U11644 (N_11644,N_9034,N_10447);
or U11645 (N_11645,N_10089,N_9252);
nand U11646 (N_11646,N_9265,N_10273);
or U11647 (N_11647,N_9119,N_9564);
and U11648 (N_11648,N_10315,N_9737);
nand U11649 (N_11649,N_10209,N_9864);
nand U11650 (N_11650,N_9986,N_10067);
nand U11651 (N_11651,N_9787,N_9755);
nor U11652 (N_11652,N_9935,N_9961);
and U11653 (N_11653,N_10250,N_9969);
nor U11654 (N_11654,N_9959,N_9489);
and U11655 (N_11655,N_9550,N_10257);
or U11656 (N_11656,N_9276,N_10375);
nor U11657 (N_11657,N_10063,N_9456);
nand U11658 (N_11658,N_9998,N_9930);
nor U11659 (N_11659,N_9939,N_10389);
or U11660 (N_11660,N_9138,N_9913);
nor U11661 (N_11661,N_10399,N_9628);
or U11662 (N_11662,N_10122,N_9678);
xor U11663 (N_11663,N_9221,N_9283);
nor U11664 (N_11664,N_10493,N_9398);
nor U11665 (N_11665,N_9731,N_9618);
and U11666 (N_11666,N_9729,N_10374);
or U11667 (N_11667,N_9906,N_9008);
nor U11668 (N_11668,N_9410,N_9574);
or U11669 (N_11669,N_9139,N_9401);
or U11670 (N_11670,N_10132,N_10409);
and U11671 (N_11671,N_9128,N_9000);
nor U11672 (N_11672,N_9846,N_10412);
or U11673 (N_11673,N_10441,N_9710);
nor U11674 (N_11674,N_10298,N_9195);
nand U11675 (N_11675,N_9579,N_10291);
or U11676 (N_11676,N_10205,N_9939);
and U11677 (N_11677,N_9184,N_9336);
or U11678 (N_11678,N_10051,N_10456);
and U11679 (N_11679,N_9855,N_9511);
nand U11680 (N_11680,N_9650,N_9147);
or U11681 (N_11681,N_9764,N_9835);
and U11682 (N_11682,N_9891,N_9937);
nand U11683 (N_11683,N_9003,N_9103);
and U11684 (N_11684,N_10152,N_9800);
and U11685 (N_11685,N_9006,N_9286);
nor U11686 (N_11686,N_9839,N_9756);
nand U11687 (N_11687,N_9315,N_9890);
and U11688 (N_11688,N_9460,N_9135);
nor U11689 (N_11689,N_9244,N_10268);
nand U11690 (N_11690,N_9858,N_9904);
nor U11691 (N_11691,N_9900,N_9909);
and U11692 (N_11692,N_10117,N_10196);
and U11693 (N_11693,N_9308,N_10426);
nand U11694 (N_11694,N_9645,N_9711);
nand U11695 (N_11695,N_9880,N_9688);
and U11696 (N_11696,N_9904,N_9094);
or U11697 (N_11697,N_10024,N_9616);
and U11698 (N_11698,N_9978,N_9666);
or U11699 (N_11699,N_9149,N_9172);
nand U11700 (N_11700,N_9857,N_9562);
nor U11701 (N_11701,N_9824,N_9008);
and U11702 (N_11702,N_10036,N_9335);
or U11703 (N_11703,N_10296,N_9155);
or U11704 (N_11704,N_9202,N_9884);
or U11705 (N_11705,N_9098,N_10485);
and U11706 (N_11706,N_9742,N_9760);
nand U11707 (N_11707,N_9973,N_9541);
and U11708 (N_11708,N_9339,N_10192);
nor U11709 (N_11709,N_10411,N_10094);
or U11710 (N_11710,N_9272,N_9960);
and U11711 (N_11711,N_10344,N_9430);
nor U11712 (N_11712,N_10407,N_9928);
or U11713 (N_11713,N_9001,N_9521);
and U11714 (N_11714,N_9001,N_9493);
and U11715 (N_11715,N_9260,N_10261);
or U11716 (N_11716,N_9171,N_10153);
and U11717 (N_11717,N_10165,N_9246);
or U11718 (N_11718,N_10012,N_10473);
or U11719 (N_11719,N_9334,N_10314);
nor U11720 (N_11720,N_9795,N_10177);
nor U11721 (N_11721,N_10045,N_9552);
and U11722 (N_11722,N_9021,N_9117);
and U11723 (N_11723,N_9018,N_10453);
nand U11724 (N_11724,N_10345,N_9689);
and U11725 (N_11725,N_9658,N_10058);
nand U11726 (N_11726,N_10431,N_9836);
or U11727 (N_11727,N_9151,N_9301);
nand U11728 (N_11728,N_9300,N_10167);
or U11729 (N_11729,N_10284,N_10137);
and U11730 (N_11730,N_9276,N_10201);
or U11731 (N_11731,N_9807,N_9951);
nand U11732 (N_11732,N_9141,N_10487);
nor U11733 (N_11733,N_9447,N_9026);
or U11734 (N_11734,N_10220,N_9763);
and U11735 (N_11735,N_9871,N_10039);
nand U11736 (N_11736,N_9929,N_10344);
or U11737 (N_11737,N_10044,N_9621);
nand U11738 (N_11738,N_9430,N_9759);
nor U11739 (N_11739,N_9041,N_9437);
nor U11740 (N_11740,N_10300,N_9305);
nand U11741 (N_11741,N_9184,N_9519);
and U11742 (N_11742,N_9140,N_10357);
nand U11743 (N_11743,N_10051,N_9819);
and U11744 (N_11744,N_9243,N_9490);
and U11745 (N_11745,N_9466,N_9105);
nor U11746 (N_11746,N_9111,N_10337);
nor U11747 (N_11747,N_9279,N_9224);
or U11748 (N_11748,N_9065,N_9926);
nor U11749 (N_11749,N_9768,N_9992);
nor U11750 (N_11750,N_10098,N_9191);
nand U11751 (N_11751,N_9321,N_10170);
nor U11752 (N_11752,N_9790,N_9206);
nor U11753 (N_11753,N_9272,N_9055);
nor U11754 (N_11754,N_10412,N_9128);
and U11755 (N_11755,N_10453,N_9721);
nor U11756 (N_11756,N_9886,N_10323);
or U11757 (N_11757,N_9122,N_9747);
nand U11758 (N_11758,N_10054,N_9653);
nand U11759 (N_11759,N_9244,N_9938);
nand U11760 (N_11760,N_10299,N_9415);
nand U11761 (N_11761,N_10010,N_9356);
or U11762 (N_11762,N_9115,N_10377);
and U11763 (N_11763,N_10422,N_9027);
or U11764 (N_11764,N_9405,N_9092);
nand U11765 (N_11765,N_9941,N_9367);
nand U11766 (N_11766,N_9319,N_9713);
nand U11767 (N_11767,N_9388,N_9044);
and U11768 (N_11768,N_10293,N_9176);
nand U11769 (N_11769,N_10045,N_9744);
or U11770 (N_11770,N_10346,N_10143);
or U11771 (N_11771,N_10413,N_10239);
or U11772 (N_11772,N_10251,N_10246);
nand U11773 (N_11773,N_10348,N_10447);
nor U11774 (N_11774,N_10149,N_9524);
and U11775 (N_11775,N_9353,N_10184);
nand U11776 (N_11776,N_9116,N_9217);
and U11777 (N_11777,N_9149,N_9115);
or U11778 (N_11778,N_10236,N_10493);
or U11779 (N_11779,N_9741,N_10075);
or U11780 (N_11780,N_10487,N_9796);
nand U11781 (N_11781,N_9007,N_9046);
or U11782 (N_11782,N_9138,N_9893);
or U11783 (N_11783,N_9169,N_9748);
nand U11784 (N_11784,N_9547,N_9296);
and U11785 (N_11785,N_10382,N_9966);
or U11786 (N_11786,N_9834,N_9018);
or U11787 (N_11787,N_9975,N_10427);
nand U11788 (N_11788,N_9695,N_9957);
nand U11789 (N_11789,N_9177,N_9543);
and U11790 (N_11790,N_10261,N_9699);
nor U11791 (N_11791,N_9163,N_9024);
nor U11792 (N_11792,N_9179,N_9562);
or U11793 (N_11793,N_10287,N_9462);
and U11794 (N_11794,N_10221,N_9697);
or U11795 (N_11795,N_9767,N_9874);
or U11796 (N_11796,N_10479,N_9248);
and U11797 (N_11797,N_10198,N_10003);
and U11798 (N_11798,N_9317,N_9012);
or U11799 (N_11799,N_9597,N_10268);
or U11800 (N_11800,N_10178,N_9049);
or U11801 (N_11801,N_9932,N_9019);
or U11802 (N_11802,N_9039,N_10326);
or U11803 (N_11803,N_10095,N_9851);
or U11804 (N_11804,N_10437,N_9113);
or U11805 (N_11805,N_9287,N_9444);
nand U11806 (N_11806,N_9315,N_9945);
and U11807 (N_11807,N_10321,N_10148);
and U11808 (N_11808,N_9439,N_9656);
nand U11809 (N_11809,N_9393,N_9542);
nand U11810 (N_11810,N_9090,N_10439);
and U11811 (N_11811,N_9267,N_9378);
nand U11812 (N_11812,N_9530,N_10237);
or U11813 (N_11813,N_10431,N_10161);
nand U11814 (N_11814,N_10325,N_9639);
nor U11815 (N_11815,N_9668,N_9144);
and U11816 (N_11816,N_9643,N_9756);
and U11817 (N_11817,N_9675,N_10360);
and U11818 (N_11818,N_10347,N_9532);
nor U11819 (N_11819,N_9391,N_9299);
nand U11820 (N_11820,N_10258,N_10005);
and U11821 (N_11821,N_9776,N_9021);
nor U11822 (N_11822,N_10467,N_9505);
nand U11823 (N_11823,N_10107,N_9356);
or U11824 (N_11824,N_9355,N_9521);
and U11825 (N_11825,N_9192,N_10108);
or U11826 (N_11826,N_9378,N_9563);
and U11827 (N_11827,N_9715,N_9567);
and U11828 (N_11828,N_10150,N_9766);
and U11829 (N_11829,N_9410,N_10328);
nor U11830 (N_11830,N_9618,N_10105);
nand U11831 (N_11831,N_9472,N_9339);
nand U11832 (N_11832,N_10264,N_10335);
nor U11833 (N_11833,N_10398,N_10402);
nor U11834 (N_11834,N_9007,N_9898);
and U11835 (N_11835,N_9422,N_10100);
nor U11836 (N_11836,N_9890,N_10134);
nand U11837 (N_11837,N_9790,N_9661);
nand U11838 (N_11838,N_9079,N_9424);
nor U11839 (N_11839,N_9228,N_10280);
nand U11840 (N_11840,N_9037,N_10056);
nor U11841 (N_11841,N_9577,N_9131);
nand U11842 (N_11842,N_9322,N_9105);
nand U11843 (N_11843,N_10144,N_10124);
nor U11844 (N_11844,N_9449,N_9509);
or U11845 (N_11845,N_10282,N_9554);
nand U11846 (N_11846,N_9334,N_10156);
or U11847 (N_11847,N_9595,N_10166);
or U11848 (N_11848,N_9888,N_9601);
nor U11849 (N_11849,N_10475,N_10446);
and U11850 (N_11850,N_9094,N_9613);
or U11851 (N_11851,N_9379,N_9058);
nand U11852 (N_11852,N_9997,N_9668);
nor U11853 (N_11853,N_10178,N_9682);
xnor U11854 (N_11854,N_10442,N_10041);
or U11855 (N_11855,N_9407,N_9105);
or U11856 (N_11856,N_9583,N_9511);
and U11857 (N_11857,N_9328,N_10475);
and U11858 (N_11858,N_9597,N_10024);
nand U11859 (N_11859,N_10308,N_9169);
and U11860 (N_11860,N_10122,N_9343);
and U11861 (N_11861,N_9618,N_9483);
nor U11862 (N_11862,N_9043,N_9509);
or U11863 (N_11863,N_10198,N_9164);
nand U11864 (N_11864,N_9472,N_9002);
and U11865 (N_11865,N_9899,N_9731);
nand U11866 (N_11866,N_10420,N_9868);
or U11867 (N_11867,N_10285,N_9243);
and U11868 (N_11868,N_10193,N_10309);
and U11869 (N_11869,N_9479,N_10008);
nor U11870 (N_11870,N_10262,N_10304);
or U11871 (N_11871,N_9226,N_9465);
nor U11872 (N_11872,N_9588,N_10241);
nand U11873 (N_11873,N_9290,N_9925);
nand U11874 (N_11874,N_9286,N_10128);
and U11875 (N_11875,N_10307,N_10402);
or U11876 (N_11876,N_9228,N_10007);
and U11877 (N_11877,N_9582,N_9014);
nand U11878 (N_11878,N_9860,N_10114);
nand U11879 (N_11879,N_9493,N_9543);
nand U11880 (N_11880,N_9324,N_9865);
nor U11881 (N_11881,N_9775,N_9615);
nand U11882 (N_11882,N_9897,N_9757);
or U11883 (N_11883,N_9131,N_10049);
nor U11884 (N_11884,N_9032,N_9348);
or U11885 (N_11885,N_9834,N_10336);
nand U11886 (N_11886,N_9999,N_9071);
or U11887 (N_11887,N_9442,N_10164);
or U11888 (N_11888,N_9715,N_10492);
and U11889 (N_11889,N_9464,N_10346);
nor U11890 (N_11890,N_9814,N_10391);
nand U11891 (N_11891,N_9616,N_9111);
nor U11892 (N_11892,N_9438,N_10305);
and U11893 (N_11893,N_9200,N_9551);
nand U11894 (N_11894,N_10221,N_10319);
or U11895 (N_11895,N_9892,N_9759);
or U11896 (N_11896,N_10333,N_10350);
nand U11897 (N_11897,N_9584,N_10385);
or U11898 (N_11898,N_10161,N_9104);
and U11899 (N_11899,N_9335,N_9772);
nand U11900 (N_11900,N_9663,N_9371);
or U11901 (N_11901,N_9738,N_9677);
nor U11902 (N_11902,N_9934,N_10055);
nand U11903 (N_11903,N_9888,N_9822);
nand U11904 (N_11904,N_9231,N_9870);
nor U11905 (N_11905,N_9352,N_9659);
nand U11906 (N_11906,N_9677,N_9057);
or U11907 (N_11907,N_10045,N_10291);
or U11908 (N_11908,N_9220,N_9087);
nor U11909 (N_11909,N_9185,N_9359);
or U11910 (N_11910,N_9512,N_9229);
nand U11911 (N_11911,N_9860,N_10066);
xor U11912 (N_11912,N_9361,N_9155);
and U11913 (N_11913,N_10205,N_10449);
and U11914 (N_11914,N_9224,N_9090);
nand U11915 (N_11915,N_9400,N_10352);
nand U11916 (N_11916,N_9346,N_9468);
nor U11917 (N_11917,N_9992,N_9085);
or U11918 (N_11918,N_9539,N_9229);
nand U11919 (N_11919,N_9866,N_10006);
or U11920 (N_11920,N_10307,N_9201);
nor U11921 (N_11921,N_10186,N_9126);
nor U11922 (N_11922,N_9714,N_9574);
nor U11923 (N_11923,N_9622,N_9379);
nand U11924 (N_11924,N_9744,N_10248);
nor U11925 (N_11925,N_9197,N_9756);
nand U11926 (N_11926,N_10233,N_10274);
and U11927 (N_11927,N_9762,N_9912);
nand U11928 (N_11928,N_9215,N_10119);
nor U11929 (N_11929,N_10052,N_9940);
nand U11930 (N_11930,N_10016,N_10271);
or U11931 (N_11931,N_9832,N_9855);
nand U11932 (N_11932,N_10106,N_9479);
nor U11933 (N_11933,N_9992,N_9594);
nand U11934 (N_11934,N_9766,N_9318);
nand U11935 (N_11935,N_9836,N_9218);
nand U11936 (N_11936,N_9676,N_9257);
nor U11937 (N_11937,N_9428,N_10033);
nor U11938 (N_11938,N_9150,N_9593);
nand U11939 (N_11939,N_9868,N_9576);
or U11940 (N_11940,N_9313,N_9407);
nor U11941 (N_11941,N_9024,N_10041);
and U11942 (N_11942,N_9056,N_9350);
nor U11943 (N_11943,N_9814,N_9898);
nand U11944 (N_11944,N_9336,N_9978);
or U11945 (N_11945,N_9181,N_10422);
and U11946 (N_11946,N_10225,N_10391);
nand U11947 (N_11947,N_10407,N_9370);
or U11948 (N_11948,N_9877,N_9495);
nor U11949 (N_11949,N_9686,N_10103);
nor U11950 (N_11950,N_9188,N_9248);
and U11951 (N_11951,N_9627,N_9204);
nor U11952 (N_11952,N_9388,N_9137);
nand U11953 (N_11953,N_10189,N_10306);
and U11954 (N_11954,N_9881,N_10345);
and U11955 (N_11955,N_10227,N_9640);
and U11956 (N_11956,N_9396,N_10269);
nor U11957 (N_11957,N_9838,N_9285);
and U11958 (N_11958,N_10072,N_9082);
or U11959 (N_11959,N_10376,N_10443);
nand U11960 (N_11960,N_9069,N_9097);
and U11961 (N_11961,N_9142,N_10404);
and U11962 (N_11962,N_10211,N_9978);
nor U11963 (N_11963,N_9561,N_9169);
or U11964 (N_11964,N_10027,N_10277);
or U11965 (N_11965,N_9337,N_9496);
and U11966 (N_11966,N_9180,N_10292);
and U11967 (N_11967,N_10259,N_10458);
or U11968 (N_11968,N_10413,N_9766);
and U11969 (N_11969,N_10003,N_9123);
and U11970 (N_11970,N_9666,N_9458);
or U11971 (N_11971,N_10144,N_9507);
and U11972 (N_11972,N_9803,N_9902);
and U11973 (N_11973,N_9500,N_10433);
or U11974 (N_11974,N_9978,N_9744);
and U11975 (N_11975,N_9896,N_9772);
and U11976 (N_11976,N_10376,N_9054);
nor U11977 (N_11977,N_9015,N_9341);
nor U11978 (N_11978,N_9072,N_10171);
nor U11979 (N_11979,N_9971,N_9552);
or U11980 (N_11980,N_9997,N_10447);
nand U11981 (N_11981,N_10343,N_9836);
nand U11982 (N_11982,N_10328,N_9438);
nand U11983 (N_11983,N_9307,N_9800);
nand U11984 (N_11984,N_9135,N_9417);
nand U11985 (N_11985,N_10338,N_9261);
and U11986 (N_11986,N_10149,N_9566);
nand U11987 (N_11987,N_9015,N_9960);
nand U11988 (N_11988,N_9100,N_10226);
or U11989 (N_11989,N_9020,N_10348);
nor U11990 (N_11990,N_9410,N_9464);
nor U11991 (N_11991,N_9356,N_9789);
and U11992 (N_11992,N_9058,N_9352);
nand U11993 (N_11993,N_9464,N_9971);
nor U11994 (N_11994,N_9742,N_10217);
or U11995 (N_11995,N_10409,N_9863);
nand U11996 (N_11996,N_10054,N_9792);
nand U11997 (N_11997,N_9395,N_9186);
xor U11998 (N_11998,N_10074,N_9571);
and U11999 (N_11999,N_10226,N_10385);
or U12000 (N_12000,N_11747,N_10932);
and U12001 (N_12001,N_10632,N_10969);
or U12002 (N_12002,N_11920,N_10901);
and U12003 (N_12003,N_10896,N_10703);
nor U12004 (N_12004,N_10535,N_11054);
or U12005 (N_12005,N_11847,N_11102);
or U12006 (N_12006,N_11228,N_10908);
xor U12007 (N_12007,N_11925,N_11866);
or U12008 (N_12008,N_11771,N_11446);
nand U12009 (N_12009,N_11786,N_11049);
and U12010 (N_12010,N_10858,N_11700);
or U12011 (N_12011,N_11275,N_10973);
nor U12012 (N_12012,N_11519,N_10546);
nand U12013 (N_12013,N_10501,N_10603);
or U12014 (N_12014,N_10729,N_11950);
nor U12015 (N_12015,N_11809,N_11114);
nor U12016 (N_12016,N_11587,N_11900);
nor U12017 (N_12017,N_11047,N_11190);
or U12018 (N_12018,N_10686,N_11041);
nor U12019 (N_12019,N_10984,N_10558);
nand U12020 (N_12020,N_11953,N_10889);
nor U12021 (N_12021,N_10562,N_11735);
nor U12022 (N_12022,N_11766,N_11635);
and U12023 (N_12023,N_11973,N_11144);
xor U12024 (N_12024,N_11202,N_11949);
and U12025 (N_12025,N_11590,N_11894);
or U12026 (N_12026,N_10977,N_10534);
nand U12027 (N_12027,N_10665,N_11475);
nand U12028 (N_12028,N_10699,N_10823);
nand U12029 (N_12029,N_11038,N_10745);
or U12030 (N_12030,N_11146,N_10503);
nor U12031 (N_12031,N_11929,N_11922);
nor U12032 (N_12032,N_11581,N_11983);
and U12033 (N_12033,N_10882,N_10862);
and U12034 (N_12034,N_10829,N_10884);
nand U12035 (N_12035,N_11611,N_11760);
nand U12036 (N_12036,N_10514,N_10926);
nor U12037 (N_12037,N_11783,N_10551);
nand U12038 (N_12038,N_10717,N_11250);
or U12039 (N_12039,N_11103,N_10772);
and U12040 (N_12040,N_11307,N_11153);
nor U12041 (N_12041,N_10892,N_11396);
and U12042 (N_12042,N_11895,N_11659);
or U12043 (N_12043,N_11946,N_11821);
or U12044 (N_12044,N_11754,N_11424);
nor U12045 (N_12045,N_11174,N_11425);
nor U12046 (N_12046,N_11876,N_11763);
nand U12047 (N_12047,N_11348,N_11397);
or U12048 (N_12048,N_11568,N_11770);
and U12049 (N_12049,N_11533,N_11552);
nand U12050 (N_12050,N_10521,N_10851);
or U12051 (N_12051,N_10671,N_11569);
and U12052 (N_12052,N_10592,N_11789);
nand U12053 (N_12053,N_11717,N_11991);
and U12054 (N_12054,N_11057,N_11784);
and U12055 (N_12055,N_11395,N_11506);
and U12056 (N_12056,N_10584,N_11402);
nand U12057 (N_12057,N_11488,N_11999);
and U12058 (N_12058,N_11882,N_11594);
nand U12059 (N_12059,N_11933,N_11811);
nor U12060 (N_12060,N_10854,N_11565);
nand U12061 (N_12061,N_11357,N_11914);
or U12062 (N_12062,N_11903,N_11217);
nor U12063 (N_12063,N_10769,N_10867);
nand U12064 (N_12064,N_11223,N_10903);
nand U12065 (N_12065,N_10661,N_11797);
nor U12066 (N_12066,N_11740,N_11582);
and U12067 (N_12067,N_11767,N_11042);
nand U12068 (N_12068,N_10972,N_10777);
nor U12069 (N_12069,N_10989,N_11753);
nor U12070 (N_12070,N_11640,N_11387);
nand U12071 (N_12071,N_11342,N_10611);
nand U12072 (N_12072,N_11714,N_10790);
or U12073 (N_12073,N_11065,N_11277);
nor U12074 (N_12074,N_11340,N_11936);
and U12075 (N_12075,N_11529,N_11432);
and U12076 (N_12076,N_10741,N_11222);
and U12077 (N_12077,N_11654,N_10815);
nor U12078 (N_12078,N_10707,N_10948);
nor U12079 (N_12079,N_11386,N_10561);
nor U12080 (N_12080,N_11334,N_11015);
nand U12081 (N_12081,N_11410,N_11155);
nand U12082 (N_12082,N_11713,N_10904);
and U12083 (N_12083,N_10833,N_11596);
nand U12084 (N_12084,N_11429,N_10590);
nand U12085 (N_12085,N_11186,N_11508);
nand U12086 (N_12086,N_11361,N_11076);
or U12087 (N_12087,N_11695,N_11551);
and U12088 (N_12088,N_11863,N_11382);
nor U12089 (N_12089,N_11848,N_11672);
and U12090 (N_12090,N_10791,N_10993);
nand U12091 (N_12091,N_11218,N_11235);
or U12092 (N_12092,N_11852,N_10610);
nand U12093 (N_12093,N_11563,N_11215);
nor U12094 (N_12094,N_10831,N_10813);
nand U12095 (N_12095,N_11749,N_11591);
nand U12096 (N_12096,N_10623,N_11282);
and U12097 (N_12097,N_11294,N_10869);
nand U12098 (N_12098,N_11002,N_11776);
and U12099 (N_12099,N_11743,N_11299);
nor U12100 (N_12100,N_11748,N_11927);
nand U12101 (N_12101,N_11124,N_11972);
nand U12102 (N_12102,N_10957,N_10995);
or U12103 (N_12103,N_11035,N_11706);
nor U12104 (N_12104,N_10848,N_11270);
or U12105 (N_12105,N_11795,N_10510);
and U12106 (N_12106,N_11355,N_11471);
nand U12107 (N_12107,N_11916,N_11673);
or U12108 (N_12108,N_11941,N_11616);
and U12109 (N_12109,N_10511,N_11491);
nand U12110 (N_12110,N_10976,N_11535);
nor U12111 (N_12111,N_10881,N_11824);
and U12112 (N_12112,N_10887,N_11530);
or U12113 (N_12113,N_11136,N_11774);
and U12114 (N_12114,N_11457,N_10682);
nand U12115 (N_12115,N_11430,N_10742);
or U12116 (N_12116,N_11990,N_10974);
nand U12117 (N_12117,N_11944,N_11333);
and U12118 (N_12118,N_10515,N_10537);
or U12119 (N_12119,N_11943,N_11321);
nor U12120 (N_12120,N_11390,N_11130);
nand U12121 (N_12121,N_11481,N_11969);
nand U12122 (N_12122,N_11661,N_11435);
xnor U12123 (N_12123,N_11165,N_10599);
nand U12124 (N_12124,N_11668,N_11674);
xor U12125 (N_12125,N_11658,N_11806);
or U12126 (N_12126,N_11602,N_11249);
xor U12127 (N_12127,N_11070,N_11585);
nor U12128 (N_12128,N_11653,N_10504);
nor U12129 (N_12129,N_11856,N_11992);
nand U12130 (N_12130,N_11884,N_11233);
or U12131 (N_12131,N_11704,N_11945);
nand U12132 (N_12132,N_11595,N_11669);
xor U12133 (N_12133,N_11864,N_11243);
and U12134 (N_12134,N_10847,N_10606);
or U12135 (N_12135,N_10685,N_10695);
nand U12136 (N_12136,N_10556,N_11648);
or U12137 (N_12137,N_10630,N_10753);
or U12138 (N_12138,N_11158,N_11421);
nand U12139 (N_12139,N_11139,N_11870);
nand U12140 (N_12140,N_11531,N_11675);
nor U12141 (N_12141,N_10966,N_11617);
nor U12142 (N_12142,N_11409,N_10722);
or U12143 (N_12143,N_10803,N_11378);
or U12144 (N_12144,N_11636,N_10960);
and U12145 (N_12145,N_11147,N_11314);
nor U12146 (N_12146,N_10523,N_10597);
and U12147 (N_12147,N_11162,N_10783);
and U12148 (N_12148,N_11733,N_11248);
and U12149 (N_12149,N_11460,N_11203);
and U12150 (N_12150,N_11752,N_10965);
nand U12151 (N_12151,N_11919,N_11601);
nand U12152 (N_12152,N_11731,N_10639);
or U12153 (N_12153,N_11997,N_11645);
and U12154 (N_12154,N_11651,N_11344);
nor U12155 (N_12155,N_11014,N_10645);
nand U12156 (N_12156,N_11678,N_11417);
nor U12157 (N_12157,N_11796,N_11204);
or U12158 (N_12158,N_11613,N_10620);
nand U12159 (N_12159,N_11461,N_10721);
nand U12160 (N_12160,N_11512,N_10517);
or U12161 (N_12161,N_11930,N_10560);
or U12162 (N_12162,N_11129,N_11918);
nor U12163 (N_12163,N_11172,N_11521);
nand U12164 (N_12164,N_11152,N_10657);
xor U12165 (N_12165,N_10547,N_11718);
or U12166 (N_12166,N_11027,N_10849);
nor U12167 (N_12167,N_11817,N_11295);
nor U12168 (N_12168,N_10894,N_11479);
nor U12169 (N_12169,N_10680,N_11939);
nand U12170 (N_12170,N_10767,N_10757);
and U12171 (N_12171,N_10575,N_10841);
nor U12172 (N_12172,N_11650,N_10796);
and U12173 (N_12173,N_10865,N_10668);
or U12174 (N_12174,N_11951,N_10990);
and U12175 (N_12175,N_11093,N_10746);
nor U12176 (N_12176,N_11280,N_11293);
or U12177 (N_12177,N_11180,N_10626);
nor U12178 (N_12178,N_10795,N_11309);
nor U12179 (N_12179,N_10621,N_11703);
or U12180 (N_12180,N_10735,N_11317);
nor U12181 (N_12181,N_11934,N_11720);
nor U12182 (N_12182,N_11626,N_10935);
nor U12183 (N_12183,N_11988,N_10733);
nor U12184 (N_12184,N_11211,N_11744);
and U12185 (N_12185,N_11554,N_11170);
nand U12186 (N_12186,N_11656,N_11520);
or U12187 (N_12187,N_11493,N_10988);
and U12188 (N_12188,N_11572,N_11257);
nand U12189 (N_12189,N_11405,N_11341);
and U12190 (N_12190,N_11517,N_11021);
and U12191 (N_12191,N_11845,N_11039);
nand U12192 (N_12192,N_11686,N_10542);
nor U12193 (N_12193,N_10540,N_11287);
or U12194 (N_12194,N_11095,N_11161);
and U12195 (N_12195,N_10507,N_11584);
and U12196 (N_12196,N_11547,N_10702);
xnor U12197 (N_12197,N_11935,N_11087);
nand U12198 (N_12198,N_11874,N_10637);
nor U12199 (N_12199,N_11148,N_10789);
nand U12200 (N_12200,N_10782,N_11841);
nor U12201 (N_12201,N_11464,N_11986);
and U12202 (N_12202,N_10730,N_11666);
nor U12203 (N_12203,N_11163,N_11906);
or U12204 (N_12204,N_10660,N_10825);
nor U12205 (N_12205,N_11016,N_10885);
or U12206 (N_12206,N_10585,N_10765);
nand U12207 (N_12207,N_11509,N_10697);
nor U12208 (N_12208,N_10544,N_11639);
nand U12209 (N_12209,N_11854,N_11351);
nor U12210 (N_12210,N_11522,N_11001);
and U12211 (N_12211,N_11226,N_10526);
and U12212 (N_12212,N_10962,N_11982);
nand U12213 (N_12213,N_10747,N_11259);
nor U12214 (N_12214,N_11137,N_11398);
and U12215 (N_12215,N_11790,N_11019);
and U12216 (N_12216,N_10898,N_11234);
and U12217 (N_12217,N_11971,N_10594);
nand U12218 (N_12218,N_11262,N_10710);
or U12219 (N_12219,N_10915,N_10955);
and U12220 (N_12220,N_10936,N_10567);
nor U12221 (N_12221,N_11091,N_11184);
or U12222 (N_12222,N_11444,N_11476);
and U12223 (N_12223,N_10835,N_11484);
and U12224 (N_12224,N_10586,N_10604);
or U12225 (N_12225,N_11928,N_10548);
or U12226 (N_12226,N_11423,N_11955);
or U12227 (N_12227,N_10737,N_11513);
nor U12228 (N_12228,N_11434,N_11059);
nor U12229 (N_12229,N_11289,N_11210);
nor U12230 (N_12230,N_10756,N_10947);
and U12231 (N_12231,N_11502,N_11119);
or U12232 (N_12232,N_10525,N_11561);
or U12233 (N_12233,N_11045,N_10840);
nor U12234 (N_12234,N_11465,N_11123);
or U12235 (N_12235,N_10805,N_10899);
and U12236 (N_12236,N_11367,N_11698);
nand U12237 (N_12237,N_10927,N_11082);
and U12238 (N_12238,N_11993,N_10814);
and U12239 (N_12239,N_11677,N_10797);
nand U12240 (N_12240,N_11800,N_10824);
nor U12241 (N_12241,N_11276,N_11187);
nor U12242 (N_12242,N_10607,N_11623);
nor U12243 (N_12243,N_10930,N_11791);
and U12244 (N_12244,N_10696,N_10786);
nor U12245 (N_12245,N_10612,N_11643);
nor U12246 (N_12246,N_10982,N_11680);
or U12247 (N_12247,N_10888,N_11505);
nand U12248 (N_12248,N_11849,N_11185);
nand U12249 (N_12249,N_10587,N_10555);
nor U12250 (N_12250,N_11160,N_10807);
nand U12251 (N_12251,N_11480,N_11813);
nand U12252 (N_12252,N_11330,N_11958);
and U12253 (N_12253,N_10543,N_11173);
and U12254 (N_12254,N_11579,N_10509);
and U12255 (N_12255,N_11808,N_11501);
or U12256 (N_12256,N_11498,N_11556);
or U12257 (N_12257,N_10785,N_10574);
and U12258 (N_12258,N_11838,N_11339);
nand U12259 (N_12259,N_11762,N_11459);
nand U12260 (N_12260,N_10978,N_11143);
and U12261 (N_12261,N_10979,N_11024);
and U12262 (N_12262,N_11792,N_11078);
or U12263 (N_12263,N_10700,N_11712);
or U12264 (N_12264,N_11592,N_11212);
or U12265 (N_12265,N_11956,N_10781);
nand U12266 (N_12266,N_11614,N_10940);
nand U12267 (N_12267,N_11157,N_11332);
nor U12268 (N_12268,N_11527,N_10941);
or U12269 (N_12269,N_11769,N_11877);
or U12270 (N_12270,N_11660,N_10655);
nand U12271 (N_12271,N_11105,N_11033);
and U12272 (N_12272,N_10541,N_11567);
and U12273 (N_12273,N_10763,N_10600);
and U12274 (N_12274,N_10837,N_11998);
nand U12275 (N_12275,N_11060,N_11192);
nor U12276 (N_12276,N_10975,N_11979);
nand U12277 (N_12277,N_10649,N_11092);
or U12278 (N_12278,N_10705,N_11963);
and U12279 (N_12279,N_11449,N_11369);
xnor U12280 (N_12280,N_10793,N_11657);
and U12281 (N_12281,N_10608,N_11883);
and U12282 (N_12282,N_11872,N_10669);
nand U12283 (N_12283,N_11633,N_11727);
nand U12284 (N_12284,N_11478,N_11085);
nor U12285 (N_12285,N_10718,N_11413);
or U12286 (N_12286,N_11031,N_11886);
and U12287 (N_12287,N_11837,N_11365);
xor U12288 (N_12288,N_11954,N_11236);
nor U12289 (N_12289,N_10748,N_10943);
nor U12290 (N_12290,N_11537,N_11490);
xor U12291 (N_12291,N_11468,N_11499);
nor U12292 (N_12292,N_11921,N_11026);
nor U12293 (N_12293,N_11067,N_10713);
and U12294 (N_12294,N_11115,N_10624);
or U12295 (N_12295,N_11063,N_11071);
or U12296 (N_12296,N_10647,N_10934);
nor U12297 (N_12297,N_11641,N_10684);
or U12298 (N_12298,N_10998,N_11156);
nor U12299 (N_12299,N_11634,N_11380);
nor U12300 (N_12300,N_11676,N_11777);
or U12301 (N_12301,N_10583,N_10743);
and U12302 (N_12302,N_10997,N_10714);
nand U12303 (N_12303,N_11216,N_11904);
and U12304 (N_12304,N_11406,N_11965);
nor U12305 (N_12305,N_11597,N_10569);
nor U12306 (N_12306,N_10709,N_11696);
and U12307 (N_12307,N_11815,N_10613);
or U12308 (N_12308,N_11758,N_10780);
or U12309 (N_12309,N_11495,N_10893);
nor U12310 (N_12310,N_10822,N_11588);
nor U12311 (N_12311,N_11354,N_11832);
nand U12312 (N_12312,N_10963,N_11685);
or U12313 (N_12313,N_11532,N_11924);
nor U12314 (N_12314,N_11843,N_11012);
xor U12315 (N_12315,N_10897,N_11559);
nand U12316 (N_12316,N_10983,N_11005);
nand U12317 (N_12317,N_10576,N_11878);
and U12318 (N_12318,N_11716,N_11463);
or U12319 (N_12319,N_11857,N_11542);
and U12320 (N_12320,N_11662,N_11942);
and U12321 (N_12321,N_11399,N_11141);
or U12322 (N_12322,N_11337,N_10673);
nand U12323 (N_12323,N_11319,N_11100);
and U12324 (N_12324,N_11244,N_11737);
nor U12325 (N_12325,N_11166,N_10866);
nand U12326 (N_12326,N_11548,N_11000);
or U12327 (N_12327,N_11072,N_11006);
nand U12328 (N_12328,N_10890,N_11169);
nand U12329 (N_12329,N_10616,N_11489);
nand U12330 (N_12330,N_11785,N_11349);
or U12331 (N_12331,N_11245,N_11231);
or U12332 (N_12332,N_10635,N_10528);
or U12333 (N_12333,N_11379,N_11073);
or U12334 (N_12334,N_11976,N_11593);
nand U12335 (N_12335,N_11994,N_11007);
and U12336 (N_12336,N_10716,N_10950);
and U12337 (N_12337,N_11394,N_11431);
nand U12338 (N_12338,N_11196,N_10817);
nand U12339 (N_12339,N_11497,N_11371);
nand U12340 (N_12340,N_10951,N_11177);
or U12341 (N_12341,N_10656,N_10931);
and U12342 (N_12342,N_10529,N_10986);
nor U12343 (N_12343,N_11194,N_11738);
nand U12344 (N_12344,N_11504,N_10627);
nand U12345 (N_12345,N_11765,N_11691);
or U12346 (N_12346,N_11948,N_10659);
or U12347 (N_12347,N_11286,N_10895);
and U12348 (N_12348,N_11603,N_11422);
nand U12349 (N_12349,N_10605,N_11631);
nor U12350 (N_12350,N_11437,N_11881);
nor U12351 (N_12351,N_10758,N_11492);
nor U12352 (N_12352,N_11909,N_11393);
or U12353 (N_12353,N_11198,N_11981);
and U12354 (N_12354,N_11246,N_11232);
or U12355 (N_12355,N_11885,N_10839);
or U12356 (N_12356,N_11473,N_11515);
and U12357 (N_12357,N_11775,N_11850);
nand U12358 (N_12358,N_11096,N_10954);
nor U12359 (N_12359,N_10877,N_11324);
nor U12360 (N_12360,N_10875,N_11412);
nor U12361 (N_12361,N_10956,N_11283);
or U12362 (N_12362,N_11618,N_11729);
or U12363 (N_12363,N_11830,N_10619);
and U12364 (N_12364,N_11020,N_10539);
and U12365 (N_12365,N_10643,N_11404);
or U12366 (N_12366,N_10910,N_10860);
nand U12367 (N_12367,N_10816,N_11284);
nor U12368 (N_12368,N_11191,N_11350);
nand U12369 (N_12369,N_11199,N_11400);
and U12370 (N_12370,N_10856,N_10698);
or U12371 (N_12371,N_10964,N_10683);
nor U12372 (N_12372,N_10646,N_10838);
nor U12373 (N_12373,N_10572,N_11606);
or U12374 (N_12374,N_11574,N_11609);
or U12375 (N_12375,N_11426,N_11443);
and U12376 (N_12376,N_10900,N_11964);
nand U12377 (N_12377,N_10644,N_11710);
or U12378 (N_12378,N_11570,N_10545);
nor U12379 (N_12379,N_11290,N_11195);
nor U12380 (N_12380,N_11818,N_11755);
nor U12381 (N_12381,N_11408,N_11528);
or U12382 (N_12382,N_11225,N_11514);
and U12383 (N_12383,N_11858,N_11401);
or U12384 (N_12384,N_10563,N_11987);
or U12385 (N_12385,N_11362,N_10651);
and U12386 (N_12386,N_11154,N_11627);
nand U12387 (N_12387,N_10640,N_11008);
nand U12388 (N_12388,N_10994,N_11684);
or U12389 (N_12389,N_10692,N_10826);
nand U12390 (N_12390,N_11168,N_11253);
nor U12391 (N_12391,N_10519,N_10842);
nor U12392 (N_12392,N_10844,N_11189);
nand U12393 (N_12393,N_10532,N_11466);
and U12394 (N_12394,N_11030,N_11229);
nor U12395 (N_12395,N_11995,N_11138);
nand U12396 (N_12396,N_11966,N_11441);
nor U12397 (N_12397,N_11834,N_10663);
and U12398 (N_12398,N_10734,N_11764);
and U12399 (N_12399,N_11266,N_11227);
or U12400 (N_12400,N_11923,N_11892);
nor U12401 (N_12401,N_10751,N_11725);
and U12402 (N_12402,N_11037,N_10725);
or U12403 (N_12403,N_10727,N_11470);
nand U12404 (N_12404,N_11311,N_10513);
nand U12405 (N_12405,N_10766,N_11086);
nor U12406 (N_12406,N_10773,N_11176);
and U12407 (N_12407,N_11018,N_11108);
nor U12408 (N_12408,N_11782,N_11325);
nor U12409 (N_12409,N_11912,N_10808);
and U12410 (N_12410,N_10634,N_10596);
nand U12411 (N_12411,N_11017,N_10723);
nor U12412 (N_12412,N_11428,N_11681);
nor U12413 (N_12413,N_11264,N_10670);
nor U12414 (N_12414,N_11305,N_10538);
and U12415 (N_12415,N_11442,N_11113);
or U12416 (N_12416,N_11241,N_10878);
and U12417 (N_12417,N_11080,N_10809);
or U12418 (N_12418,N_11901,N_11252);
nor U12419 (N_12419,N_10872,N_10873);
nor U12420 (N_12420,N_11118,N_10968);
and U12421 (N_12421,N_10715,N_11183);
nand U12422 (N_12422,N_10602,N_10739);
or U12423 (N_12423,N_11134,N_11828);
nand U12424 (N_12424,N_11860,N_11109);
and U12425 (N_12425,N_11302,N_11384);
and U12426 (N_12426,N_10502,N_10689);
nand U12427 (N_12427,N_11967,N_11296);
and U12428 (N_12428,N_11975,N_11077);
nand U12429 (N_12429,N_10724,N_10629);
nand U12430 (N_12430,N_11214,N_10706);
and U12431 (N_12431,N_11540,N_10638);
and U12432 (N_12432,N_10880,N_11873);
nand U12433 (N_12433,N_11897,N_11208);
or U12434 (N_12434,N_11193,N_11663);
nor U12435 (N_12435,N_10571,N_11539);
nand U12436 (N_12436,N_11411,N_11051);
nor U12437 (N_12437,N_11306,N_11074);
nor U12438 (N_12438,N_11871,N_10861);
or U12439 (N_12439,N_11826,N_11642);
and U12440 (N_12440,N_11458,N_10531);
and U12441 (N_12441,N_10759,N_10768);
nand U12442 (N_12442,N_11794,N_11612);
or U12443 (N_12443,N_10731,N_11316);
or U12444 (N_12444,N_10749,N_11022);
nor U12445 (N_12445,N_10701,N_10999);
and U12446 (N_12446,N_11932,N_10593);
and U12447 (N_12447,N_11523,N_10863);
or U12448 (N_12448,N_11805,N_11525);
xor U12449 (N_12449,N_11261,N_11343);
or U12450 (N_12450,N_11482,N_11439);
nand U12451 (N_12451,N_11297,N_11238);
nand U12452 (N_12452,N_11624,N_11391);
nand U12453 (N_12453,N_11798,N_10553);
nand U12454 (N_12454,N_10530,N_11915);
nor U12455 (N_12455,N_10879,N_10764);
and U12456 (N_12456,N_11197,N_11793);
and U12457 (N_12457,N_10949,N_10917);
nand U12458 (N_12458,N_11880,N_11996);
and U12459 (N_12459,N_11959,N_11589);
nor U12460 (N_12460,N_11200,N_10928);
nand U12461 (N_12461,N_11736,N_11911);
nor U12462 (N_12462,N_11075,N_11558);
or U12463 (N_12463,N_10843,N_10981);
or U12464 (N_12464,N_11630,N_11107);
nor U12465 (N_12465,N_11910,N_11511);
nor U12466 (N_12466,N_10810,N_10580);
nor U12467 (N_12467,N_11167,N_10588);
and U12468 (N_12468,N_10920,N_10991);
or U12469 (N_12469,N_11814,N_11761);
or U12470 (N_12470,N_11013,N_11907);
or U12471 (N_12471,N_11106,N_10775);
nand U12472 (N_12472,N_11003,N_11048);
or U12473 (N_12473,N_11781,N_11719);
and U12474 (N_12474,N_11750,N_11009);
nand U12475 (N_12475,N_10818,N_11285);
nand U12476 (N_12476,N_11110,N_11621);
or U12477 (N_12477,N_11455,N_10970);
nor U12478 (N_12478,N_11483,N_11576);
nand U12479 (N_12479,N_10578,N_10598);
xor U12480 (N_12480,N_11968,N_10985);
nand U12481 (N_12481,N_11632,N_11879);
nand U12482 (N_12482,N_10711,N_11940);
nor U12483 (N_12483,N_11836,N_10836);
and U12484 (N_12484,N_10883,N_10508);
nand U12485 (N_12485,N_11052,N_11112);
or U12486 (N_12486,N_11890,N_10771);
nand U12487 (N_12487,N_11345,N_11328);
and U12488 (N_12488,N_10520,N_11757);
nor U12489 (N_12489,N_11580,N_10688);
or U12490 (N_12490,N_11827,N_10601);
nor U12491 (N_12491,N_10615,N_10577);
nor U12492 (N_12492,N_11810,N_11705);
nand U12493 (N_12493,N_11577,N_10944);
nor U12494 (N_12494,N_11825,N_10568);
nand U12495 (N_12495,N_10552,N_11802);
or U12496 (N_12496,N_11573,N_11178);
and U12497 (N_12497,N_10516,N_11977);
and U12498 (N_12498,N_11534,N_10664);
or U12499 (N_12499,N_11619,N_10874);
and U12500 (N_12500,N_10812,N_11853);
nor U12501 (N_12501,N_11416,N_11844);
nor U12502 (N_12502,N_10828,N_10961);
nand U12503 (N_12503,N_11260,N_11089);
and U12504 (N_12504,N_10726,N_11628);
nor U12505 (N_12505,N_11242,N_10570);
nand U12506 (N_12506,N_11715,N_11181);
nand U12507 (N_12507,N_10762,N_10609);
or U12508 (N_12508,N_11902,N_10591);
nand U12509 (N_12509,N_10937,N_11472);
and U12510 (N_12510,N_10738,N_10752);
and U12511 (N_12511,N_11831,N_11058);
and U12512 (N_12512,N_10693,N_11304);
nand U12513 (N_12513,N_10933,N_11851);
nor U12514 (N_12514,N_11622,N_11575);
and U12515 (N_12515,N_11164,N_11046);
and U12516 (N_12516,N_10675,N_11440);
or U12517 (N_12517,N_11315,N_11679);
and U12518 (N_12518,N_10559,N_11247);
and U12519 (N_12519,N_10720,N_10736);
nand U12520 (N_12520,N_10918,N_11445);
nor U12521 (N_12521,N_11646,N_11420);
or U12522 (N_12522,N_11739,N_11553);
nor U12523 (N_12523,N_11607,N_11418);
nand U12524 (N_12524,N_10652,N_10614);
nand U12525 (N_12525,N_11835,N_11044);
or U12526 (N_12526,N_11145,N_11751);
nand U12527 (N_12527,N_10914,N_11980);
or U12528 (N_12528,N_11313,N_11926);
nor U12529 (N_12529,N_10784,N_11376);
and U12530 (N_12530,N_11462,N_11694);
or U12531 (N_12531,N_10681,N_11846);
and U12532 (N_12532,N_11823,N_10549);
and U12533 (N_12533,N_11723,N_11331);
nor U12534 (N_12534,N_11029,N_10524);
or U12535 (N_12535,N_10846,N_11543);
or U12536 (N_12536,N_11487,N_11448);
and U12537 (N_12537,N_11649,N_10924);
and U12538 (N_12538,N_10674,N_10617);
or U12539 (N_12539,N_10891,N_11084);
nor U12540 (N_12540,N_11383,N_11724);
nand U12541 (N_12541,N_11224,N_10633);
nor U12542 (N_12542,N_10834,N_11583);
nand U12543 (N_12543,N_11812,N_11010);
and U12544 (N_12544,N_11670,N_11056);
nand U12545 (N_12545,N_11905,N_10876);
and U12546 (N_12546,N_11358,N_11374);
nand U12547 (N_12547,N_10518,N_11230);
nand U12548 (N_12548,N_11557,N_11629);
nand U12549 (N_12549,N_11258,N_11855);
and U12550 (N_12550,N_11083,N_11300);
nand U12551 (N_12551,N_11875,N_11549);
nor U12552 (N_12552,N_11206,N_11507);
nor U12553 (N_12553,N_11151,N_11373);
or U12554 (N_12554,N_10536,N_11599);
nor U12555 (N_12555,N_11667,N_11278);
and U12556 (N_12556,N_11689,N_11291);
and U12557 (N_12557,N_10800,N_11709);
nor U12558 (N_12558,N_10958,N_10907);
nand U12559 (N_12559,N_10618,N_10820);
nand U12560 (N_12560,N_11773,N_11268);
nand U12561 (N_12561,N_11256,N_11213);
and U12562 (N_12562,N_10821,N_10802);
nor U12563 (N_12563,N_11370,N_11069);
nor U12564 (N_12564,N_11079,N_11862);
or U12565 (N_12565,N_11989,N_10589);
and U12566 (N_12566,N_11220,N_11887);
and U12567 (N_12567,N_11081,N_11389);
nand U12568 (N_12568,N_11687,N_10760);
and U12569 (N_12569,N_11707,N_10666);
nor U12570 (N_12570,N_10658,N_11545);
and U12571 (N_12571,N_11407,N_11359);
and U12572 (N_12572,N_11962,N_11388);
xnor U12573 (N_12573,N_11500,N_11840);
nand U12574 (N_12574,N_11598,N_10929);
nor U12575 (N_12575,N_11171,N_10533);
nand U12576 (N_12576,N_11899,N_10650);
nand U12577 (N_12577,N_11415,N_11833);
nand U12578 (N_12578,N_11518,N_11829);
nor U12579 (N_12579,N_11615,N_11127);
nor U12580 (N_12580,N_10565,N_11759);
nor U12581 (N_12581,N_10811,N_11023);
or U12582 (N_12582,N_10761,N_11061);
or U12583 (N_12583,N_10776,N_10704);
nand U12584 (N_12584,N_11188,N_11279);
and U12585 (N_12585,N_11891,N_11353);
nor U12586 (N_12586,N_10952,N_11111);
nor U12587 (N_12587,N_11839,N_11702);
and U12588 (N_12588,N_10636,N_10845);
and U12589 (N_12589,N_11043,N_11125);
nand U12590 (N_12590,N_10996,N_10916);
nor U12591 (N_12591,N_11372,N_11272);
nor U12592 (N_12592,N_11467,N_10708);
and U12593 (N_12593,N_11638,N_11697);
nand U12594 (N_12594,N_11427,N_11436);
or U12595 (N_12595,N_10566,N_11801);
nand U12596 (N_12596,N_11240,N_11064);
or U12597 (N_12597,N_10679,N_11721);
nand U12598 (N_12598,N_11456,N_10654);
nand U12599 (N_12599,N_11032,N_11780);
nor U12600 (N_12600,N_11620,N_11931);
nor U12601 (N_12601,N_11947,N_11356);
nand U12602 (N_12602,N_11360,N_11768);
nand U12603 (N_12603,N_11779,N_11366);
nand U12604 (N_12604,N_11693,N_11126);
or U12605 (N_12605,N_10971,N_11338);
or U12606 (N_12606,N_10864,N_11133);
or U12607 (N_12607,N_10579,N_11322);
or U12608 (N_12608,N_11474,N_11438);
nor U12609 (N_12609,N_11560,N_11269);
or U12610 (N_12610,N_10923,N_11098);
nor U12611 (N_12611,N_11336,N_10853);
and U12612 (N_12612,N_11335,N_11536);
or U12613 (N_12613,N_10987,N_11961);
or U12614 (N_12614,N_10755,N_11756);
nor U12615 (N_12615,N_11034,N_11869);
nand U12616 (N_12616,N_11665,N_10806);
nor U12617 (N_12617,N_10625,N_11055);
or U12618 (N_12618,N_11952,N_10938);
or U12619 (N_12619,N_11375,N_11053);
or U12620 (N_12620,N_10687,N_10564);
and U12621 (N_12621,N_11451,N_10527);
nor U12622 (N_12622,N_10788,N_11730);
and U12623 (N_12623,N_11889,N_11816);
and U12624 (N_12624,N_11453,N_10804);
and U12625 (N_12625,N_10909,N_10728);
nand U12626 (N_12626,N_11159,N_11555);
nor U12627 (N_12627,N_10919,N_11040);
nor U12628 (N_12628,N_11526,N_11728);
xor U12629 (N_12629,N_10770,N_10801);
xnor U12630 (N_12630,N_11004,N_11861);
nor U12631 (N_12631,N_10942,N_11647);
nand U12632 (N_12632,N_11312,N_11265);
nor U12633 (N_12633,N_11893,N_11711);
nand U12634 (N_12634,N_10628,N_11608);
and U12635 (N_12635,N_11699,N_10631);
nor U12636 (N_12636,N_10905,N_10672);
nor U12637 (N_12637,N_10522,N_11320);
or U12638 (N_12638,N_11985,N_10921);
nand U12639 (N_12639,N_11804,N_10792);
or U12640 (N_12640,N_11510,N_10855);
and U12641 (N_12641,N_11454,N_11363);
and U12642 (N_12642,N_10959,N_11352);
nor U12643 (N_12643,N_11516,N_10754);
nand U12644 (N_12644,N_11538,N_11447);
and U12645 (N_12645,N_11150,N_10678);
or U12646 (N_12646,N_10925,N_11094);
nand U12647 (N_12647,N_11419,N_10913);
nor U12648 (N_12648,N_10799,N_11726);
or U12649 (N_12649,N_11741,N_11062);
or U12650 (N_12650,N_11550,N_11414);
nand U12651 (N_12651,N_11722,N_11381);
or U12652 (N_12652,N_10505,N_10830);
nand U12653 (N_12653,N_11149,N_10744);
or U12654 (N_12654,N_11140,N_10550);
nor U12655 (N_12655,N_11571,N_11822);
nor U12656 (N_12656,N_11271,N_11025);
and U12657 (N_12657,N_11960,N_10676);
and U12658 (N_12658,N_11274,N_11368);
and U12659 (N_12659,N_11868,N_11564);
nor U12660 (N_12660,N_11820,N_11066);
and U12661 (N_12661,N_11131,N_11255);
nor U12662 (N_12662,N_10992,N_11655);
nand U12663 (N_12663,N_11068,N_11347);
nand U12664 (N_12664,N_11205,N_11310);
or U12665 (N_12665,N_11541,N_11524);
nor U12666 (N_12666,N_10557,N_10622);
and U12667 (N_12667,N_10740,N_11819);
and U12668 (N_12668,N_10852,N_11600);
nand U12669 (N_12669,N_11970,N_11267);
nand U12670 (N_12670,N_10857,N_11896);
nor U12671 (N_12671,N_10500,N_11403);
or U12672 (N_12672,N_11732,N_11690);
nand U12673 (N_12673,N_11683,N_11219);
nor U12674 (N_12674,N_11128,N_11708);
nand U12675 (N_12675,N_11308,N_10667);
nor U12676 (N_12676,N_10859,N_10581);
or U12677 (N_12677,N_10691,N_11135);
nor U12678 (N_12678,N_11298,N_11254);
and U12679 (N_12679,N_11544,N_11239);
nor U12680 (N_12680,N_11898,N_10886);
nand U12681 (N_12681,N_10642,N_10850);
or U12682 (N_12682,N_11605,N_11122);
or U12683 (N_12683,N_11503,N_10794);
nor U12684 (N_12684,N_11908,N_11664);
and U12685 (N_12685,N_10662,N_11859);
and U12686 (N_12686,N_10573,N_11701);
nor U12687 (N_12687,N_11938,N_10774);
nor U12688 (N_12688,N_10945,N_11099);
or U12689 (N_12689,N_10712,N_11807);
nor U12690 (N_12690,N_11392,N_11385);
nor U12691 (N_12691,N_11090,N_10798);
xnor U12692 (N_12692,N_11097,N_11292);
nand U12693 (N_12693,N_11496,N_11799);
or U12694 (N_12694,N_11546,N_10554);
nand U12695 (N_12695,N_11477,N_11562);
nor U12696 (N_12696,N_11209,N_10912);
or U12697 (N_12697,N_10911,N_11984);
nand U12698 (N_12698,N_10506,N_11772);
nor U12699 (N_12699,N_11842,N_11327);
and U12700 (N_12700,N_10870,N_11364);
nor U12701 (N_12701,N_11088,N_10980);
nand U12702 (N_12702,N_11652,N_11303);
or U12703 (N_12703,N_11301,N_11117);
xor U12704 (N_12704,N_11175,N_11787);
nor U12705 (N_12705,N_11865,N_11104);
or U12706 (N_12706,N_10819,N_10778);
nor U12707 (N_12707,N_11323,N_11028);
nor U12708 (N_12708,N_11888,N_10732);
nor U12709 (N_12709,N_10582,N_11251);
nor U12710 (N_12710,N_11671,N_11221);
nor U12711 (N_12711,N_11637,N_10871);
nand U12712 (N_12712,N_10750,N_11610);
or U12713 (N_12713,N_11746,N_11329);
or U12714 (N_12714,N_11318,N_11486);
or U12715 (N_12715,N_11377,N_10719);
or U12716 (N_12716,N_11625,N_11742);
and U12717 (N_12717,N_10779,N_10953);
nand U12718 (N_12718,N_11682,N_11011);
nand U12719 (N_12719,N_11263,N_11803);
and U12720 (N_12720,N_10868,N_11433);
nand U12721 (N_12721,N_10906,N_10939);
and U12722 (N_12722,N_11957,N_10827);
or U12723 (N_12723,N_11586,N_11237);
and U12724 (N_12724,N_10641,N_10648);
nor U12725 (N_12725,N_11452,N_11913);
or U12726 (N_12726,N_10677,N_10694);
or U12727 (N_12727,N_10946,N_11692);
or U12728 (N_12728,N_11566,N_11450);
and U12729 (N_12729,N_10653,N_11281);
or U12730 (N_12730,N_11132,N_11745);
nand U12731 (N_12731,N_11974,N_10690);
nor U12732 (N_12732,N_11346,N_11788);
or U12733 (N_12733,N_11494,N_11978);
and U12734 (N_12734,N_11101,N_11207);
nor U12735 (N_12735,N_11036,N_11469);
nand U12736 (N_12736,N_11578,N_11688);
or U12737 (N_12737,N_11116,N_11485);
or U12738 (N_12738,N_11050,N_11734);
or U12739 (N_12739,N_10787,N_10902);
or U12740 (N_12740,N_11120,N_11182);
nand U12741 (N_12741,N_11604,N_11778);
nor U12742 (N_12742,N_11179,N_10967);
xor U12743 (N_12743,N_11917,N_10832);
xor U12744 (N_12744,N_11121,N_11288);
nand U12745 (N_12745,N_11273,N_11867);
nand U12746 (N_12746,N_11201,N_11142);
or U12747 (N_12747,N_10595,N_11326);
nor U12748 (N_12748,N_11644,N_11937);
xor U12749 (N_12749,N_10512,N_10922);
nor U12750 (N_12750,N_10803,N_10893);
nor U12751 (N_12751,N_11734,N_11461);
and U12752 (N_12752,N_11545,N_11492);
or U12753 (N_12753,N_11522,N_11246);
nand U12754 (N_12754,N_11451,N_11962);
or U12755 (N_12755,N_11080,N_10889);
or U12756 (N_12756,N_10944,N_11642);
nor U12757 (N_12757,N_10903,N_10820);
nor U12758 (N_12758,N_10690,N_11252);
and U12759 (N_12759,N_11545,N_10533);
or U12760 (N_12760,N_11356,N_11515);
and U12761 (N_12761,N_11077,N_11497);
nand U12762 (N_12762,N_11499,N_11882);
and U12763 (N_12763,N_10506,N_11837);
and U12764 (N_12764,N_11915,N_10815);
nand U12765 (N_12765,N_10838,N_11028);
or U12766 (N_12766,N_11091,N_11217);
nand U12767 (N_12767,N_11795,N_11160);
and U12768 (N_12768,N_10814,N_10777);
nand U12769 (N_12769,N_11714,N_11828);
nor U12770 (N_12770,N_11297,N_10753);
or U12771 (N_12771,N_10798,N_11831);
and U12772 (N_12772,N_11887,N_11764);
or U12773 (N_12773,N_10801,N_10852);
nand U12774 (N_12774,N_10510,N_11888);
nand U12775 (N_12775,N_10855,N_11436);
or U12776 (N_12776,N_11344,N_11842);
and U12777 (N_12777,N_11262,N_11835);
nand U12778 (N_12778,N_10794,N_11929);
nand U12779 (N_12779,N_10671,N_11953);
or U12780 (N_12780,N_11471,N_11058);
nor U12781 (N_12781,N_10806,N_11387);
and U12782 (N_12782,N_11792,N_11749);
or U12783 (N_12783,N_11515,N_11377);
nand U12784 (N_12784,N_11064,N_11159);
nor U12785 (N_12785,N_11668,N_11445);
nand U12786 (N_12786,N_10783,N_11309);
and U12787 (N_12787,N_11233,N_11800);
or U12788 (N_12788,N_11166,N_11683);
nand U12789 (N_12789,N_11401,N_11938);
and U12790 (N_12790,N_11237,N_11888);
or U12791 (N_12791,N_10893,N_11688);
and U12792 (N_12792,N_11259,N_11773);
nor U12793 (N_12793,N_11887,N_10815);
nor U12794 (N_12794,N_11163,N_11490);
nor U12795 (N_12795,N_10706,N_11617);
nand U12796 (N_12796,N_11239,N_10887);
and U12797 (N_12797,N_11516,N_11367);
nand U12798 (N_12798,N_11717,N_10770);
nand U12799 (N_12799,N_11827,N_11676);
and U12800 (N_12800,N_11916,N_10692);
or U12801 (N_12801,N_10791,N_11797);
nor U12802 (N_12802,N_11837,N_10721);
or U12803 (N_12803,N_11639,N_11190);
or U12804 (N_12804,N_10614,N_11394);
or U12805 (N_12805,N_11273,N_11649);
or U12806 (N_12806,N_10557,N_11532);
and U12807 (N_12807,N_10821,N_11611);
nand U12808 (N_12808,N_10999,N_11656);
or U12809 (N_12809,N_11622,N_11479);
nand U12810 (N_12810,N_10948,N_11316);
nor U12811 (N_12811,N_11002,N_10830);
and U12812 (N_12812,N_11731,N_11053);
nand U12813 (N_12813,N_11201,N_11310);
or U12814 (N_12814,N_11571,N_10509);
or U12815 (N_12815,N_11602,N_11225);
or U12816 (N_12816,N_11321,N_11596);
or U12817 (N_12817,N_11023,N_11865);
nand U12818 (N_12818,N_10539,N_10737);
nor U12819 (N_12819,N_11223,N_11292);
nand U12820 (N_12820,N_10569,N_11429);
and U12821 (N_12821,N_10682,N_11963);
nor U12822 (N_12822,N_10558,N_10572);
and U12823 (N_12823,N_11753,N_11348);
nand U12824 (N_12824,N_10785,N_11343);
xnor U12825 (N_12825,N_10924,N_10932);
or U12826 (N_12826,N_11475,N_10846);
nand U12827 (N_12827,N_10916,N_11085);
nand U12828 (N_12828,N_11157,N_11447);
nor U12829 (N_12829,N_10738,N_11037);
and U12830 (N_12830,N_10985,N_11839);
nand U12831 (N_12831,N_11321,N_11855);
and U12832 (N_12832,N_10735,N_10803);
or U12833 (N_12833,N_11327,N_10837);
nand U12834 (N_12834,N_10941,N_10673);
or U12835 (N_12835,N_11769,N_10802);
nor U12836 (N_12836,N_10793,N_11724);
nand U12837 (N_12837,N_11353,N_10614);
and U12838 (N_12838,N_11094,N_10830);
and U12839 (N_12839,N_11677,N_10776);
nand U12840 (N_12840,N_10640,N_11432);
nand U12841 (N_12841,N_11084,N_10623);
and U12842 (N_12842,N_11046,N_10836);
or U12843 (N_12843,N_11482,N_11603);
and U12844 (N_12844,N_11249,N_11876);
nand U12845 (N_12845,N_11607,N_11464);
nand U12846 (N_12846,N_10675,N_10574);
or U12847 (N_12847,N_10599,N_11809);
nand U12848 (N_12848,N_10984,N_11587);
or U12849 (N_12849,N_10870,N_10842);
nand U12850 (N_12850,N_11758,N_10821);
nand U12851 (N_12851,N_10521,N_11075);
or U12852 (N_12852,N_11791,N_11316);
nor U12853 (N_12853,N_10898,N_10625);
nand U12854 (N_12854,N_11933,N_11148);
nand U12855 (N_12855,N_11268,N_11782);
nand U12856 (N_12856,N_11029,N_10818);
nor U12857 (N_12857,N_11654,N_11738);
and U12858 (N_12858,N_11856,N_11022);
and U12859 (N_12859,N_11535,N_11026);
or U12860 (N_12860,N_11480,N_11299);
or U12861 (N_12861,N_11135,N_11385);
and U12862 (N_12862,N_11558,N_11616);
nand U12863 (N_12863,N_11601,N_11178);
nor U12864 (N_12864,N_10914,N_11719);
and U12865 (N_12865,N_10760,N_10663);
nor U12866 (N_12866,N_10529,N_10947);
or U12867 (N_12867,N_10795,N_10605);
or U12868 (N_12868,N_11498,N_10768);
nor U12869 (N_12869,N_11450,N_11884);
and U12870 (N_12870,N_10584,N_11064);
nor U12871 (N_12871,N_11200,N_11306);
or U12872 (N_12872,N_10860,N_11155);
and U12873 (N_12873,N_11036,N_11657);
nor U12874 (N_12874,N_11592,N_10871);
and U12875 (N_12875,N_10616,N_10512);
nor U12876 (N_12876,N_11361,N_11659);
nor U12877 (N_12877,N_11390,N_11740);
and U12878 (N_12878,N_11190,N_10929);
and U12879 (N_12879,N_11598,N_10990);
nor U12880 (N_12880,N_11230,N_11772);
or U12881 (N_12881,N_11577,N_11306);
nand U12882 (N_12882,N_11205,N_11290);
nor U12883 (N_12883,N_11261,N_11488);
and U12884 (N_12884,N_10900,N_10998);
and U12885 (N_12885,N_11469,N_10959);
nand U12886 (N_12886,N_11902,N_11743);
nand U12887 (N_12887,N_11568,N_11075);
or U12888 (N_12888,N_11488,N_11303);
or U12889 (N_12889,N_11510,N_11310);
and U12890 (N_12890,N_10834,N_11062);
nor U12891 (N_12891,N_11235,N_11207);
nor U12892 (N_12892,N_10700,N_11049);
and U12893 (N_12893,N_10656,N_11395);
or U12894 (N_12894,N_11172,N_11130);
nand U12895 (N_12895,N_11560,N_10931);
nand U12896 (N_12896,N_11603,N_10612);
nand U12897 (N_12897,N_10876,N_11209);
or U12898 (N_12898,N_10879,N_11884);
nand U12899 (N_12899,N_11877,N_11109);
nor U12900 (N_12900,N_11412,N_11174);
or U12901 (N_12901,N_10790,N_10514);
nor U12902 (N_12902,N_11360,N_11060);
nor U12903 (N_12903,N_11634,N_11189);
or U12904 (N_12904,N_10537,N_10521);
nor U12905 (N_12905,N_11898,N_11954);
and U12906 (N_12906,N_11373,N_11939);
or U12907 (N_12907,N_10797,N_11976);
and U12908 (N_12908,N_11648,N_10729);
nand U12909 (N_12909,N_11700,N_11447);
nand U12910 (N_12910,N_11705,N_11341);
and U12911 (N_12911,N_11323,N_11935);
nor U12912 (N_12912,N_11040,N_11335);
or U12913 (N_12913,N_11660,N_11684);
and U12914 (N_12914,N_11614,N_10817);
and U12915 (N_12915,N_11377,N_10535);
nor U12916 (N_12916,N_10934,N_11319);
and U12917 (N_12917,N_10846,N_11848);
nand U12918 (N_12918,N_11242,N_10723);
nor U12919 (N_12919,N_11378,N_11229);
nor U12920 (N_12920,N_11369,N_10792);
and U12921 (N_12921,N_11656,N_10684);
and U12922 (N_12922,N_11509,N_11103);
or U12923 (N_12923,N_11999,N_11474);
nor U12924 (N_12924,N_11461,N_11476);
and U12925 (N_12925,N_10774,N_11846);
or U12926 (N_12926,N_11660,N_10825);
or U12927 (N_12927,N_11189,N_10885);
nand U12928 (N_12928,N_11848,N_11633);
and U12929 (N_12929,N_11852,N_10891);
or U12930 (N_12930,N_11120,N_11653);
or U12931 (N_12931,N_10855,N_11113);
nand U12932 (N_12932,N_10993,N_10947);
nor U12933 (N_12933,N_11468,N_11181);
or U12934 (N_12934,N_10605,N_11710);
nand U12935 (N_12935,N_11760,N_11027);
nand U12936 (N_12936,N_11299,N_10689);
nor U12937 (N_12937,N_11223,N_11304);
and U12938 (N_12938,N_11052,N_10693);
or U12939 (N_12939,N_11837,N_11594);
nor U12940 (N_12940,N_10638,N_10724);
nand U12941 (N_12941,N_11904,N_10532);
nor U12942 (N_12942,N_10663,N_10995);
or U12943 (N_12943,N_11370,N_10785);
and U12944 (N_12944,N_11539,N_10547);
nor U12945 (N_12945,N_11076,N_11750);
and U12946 (N_12946,N_10941,N_11965);
or U12947 (N_12947,N_10603,N_10637);
xor U12948 (N_12948,N_11145,N_11459);
nor U12949 (N_12949,N_11521,N_11786);
and U12950 (N_12950,N_10700,N_11296);
nor U12951 (N_12951,N_11686,N_11131);
xnor U12952 (N_12952,N_11994,N_11389);
and U12953 (N_12953,N_11071,N_11599);
nor U12954 (N_12954,N_11782,N_10950);
nand U12955 (N_12955,N_11914,N_10915);
and U12956 (N_12956,N_11607,N_10793);
nand U12957 (N_12957,N_10996,N_11416);
nor U12958 (N_12958,N_11278,N_11383);
and U12959 (N_12959,N_11844,N_11476);
and U12960 (N_12960,N_11230,N_10848);
or U12961 (N_12961,N_10971,N_10965);
or U12962 (N_12962,N_10956,N_11871);
and U12963 (N_12963,N_10694,N_11254);
or U12964 (N_12964,N_10878,N_11714);
nor U12965 (N_12965,N_10559,N_10754);
nand U12966 (N_12966,N_10598,N_11606);
or U12967 (N_12967,N_10646,N_10630);
and U12968 (N_12968,N_10508,N_11781);
and U12969 (N_12969,N_10611,N_10877);
nand U12970 (N_12970,N_10810,N_11403);
and U12971 (N_12971,N_10715,N_11071);
nand U12972 (N_12972,N_11467,N_11723);
and U12973 (N_12973,N_11506,N_11567);
nor U12974 (N_12974,N_11570,N_10853);
nor U12975 (N_12975,N_10777,N_11485);
or U12976 (N_12976,N_11059,N_10941);
nor U12977 (N_12977,N_10992,N_10750);
nor U12978 (N_12978,N_11541,N_11774);
and U12979 (N_12979,N_11714,N_10928);
nor U12980 (N_12980,N_11911,N_11778);
nand U12981 (N_12981,N_11893,N_11413);
nor U12982 (N_12982,N_11264,N_11560);
nand U12983 (N_12983,N_11418,N_11911);
and U12984 (N_12984,N_11268,N_11346);
or U12985 (N_12985,N_11145,N_11207);
and U12986 (N_12986,N_10679,N_10942);
nand U12987 (N_12987,N_11213,N_11536);
or U12988 (N_12988,N_11163,N_10574);
or U12989 (N_12989,N_11409,N_10505);
nor U12990 (N_12990,N_11301,N_11351);
and U12991 (N_12991,N_11056,N_11681);
nand U12992 (N_12992,N_11515,N_11438);
and U12993 (N_12993,N_10611,N_10614);
and U12994 (N_12994,N_11802,N_10554);
and U12995 (N_12995,N_11893,N_11642);
nand U12996 (N_12996,N_11363,N_11356);
or U12997 (N_12997,N_11048,N_10946);
nor U12998 (N_12998,N_11188,N_11863);
nor U12999 (N_12999,N_10819,N_11015);
and U13000 (N_13000,N_11822,N_10560);
nor U13001 (N_13001,N_11437,N_11053);
nor U13002 (N_13002,N_11855,N_11836);
nor U13003 (N_13003,N_11051,N_11029);
nand U13004 (N_13004,N_11377,N_11699);
and U13005 (N_13005,N_11179,N_11351);
nand U13006 (N_13006,N_11299,N_11442);
and U13007 (N_13007,N_10921,N_11886);
and U13008 (N_13008,N_10743,N_11838);
nor U13009 (N_13009,N_10897,N_11018);
or U13010 (N_13010,N_11124,N_10516);
nor U13011 (N_13011,N_11173,N_11137);
and U13012 (N_13012,N_11411,N_10661);
and U13013 (N_13013,N_11448,N_10573);
nand U13014 (N_13014,N_10649,N_11398);
nand U13015 (N_13015,N_11149,N_10559);
and U13016 (N_13016,N_10653,N_11838);
and U13017 (N_13017,N_11936,N_11623);
nor U13018 (N_13018,N_10652,N_11755);
and U13019 (N_13019,N_11805,N_10840);
nand U13020 (N_13020,N_11123,N_11397);
and U13021 (N_13021,N_11180,N_11076);
xor U13022 (N_13022,N_11236,N_11296);
nor U13023 (N_13023,N_10512,N_10514);
nor U13024 (N_13024,N_11290,N_11188);
or U13025 (N_13025,N_10673,N_11073);
and U13026 (N_13026,N_10984,N_11810);
or U13027 (N_13027,N_10647,N_10530);
or U13028 (N_13028,N_10843,N_11679);
or U13029 (N_13029,N_11725,N_11763);
nor U13030 (N_13030,N_11508,N_11401);
nor U13031 (N_13031,N_11499,N_11464);
or U13032 (N_13032,N_11488,N_11930);
and U13033 (N_13033,N_11822,N_11734);
nand U13034 (N_13034,N_10768,N_10772);
or U13035 (N_13035,N_11155,N_10919);
xnor U13036 (N_13036,N_10820,N_11452);
nor U13037 (N_13037,N_11665,N_11732);
or U13038 (N_13038,N_10801,N_11838);
or U13039 (N_13039,N_11875,N_11453);
or U13040 (N_13040,N_10601,N_11389);
and U13041 (N_13041,N_11057,N_11455);
or U13042 (N_13042,N_10655,N_11860);
and U13043 (N_13043,N_10885,N_11295);
and U13044 (N_13044,N_11765,N_11757);
or U13045 (N_13045,N_10692,N_10966);
or U13046 (N_13046,N_11323,N_11942);
nor U13047 (N_13047,N_11824,N_11794);
nand U13048 (N_13048,N_11963,N_11053);
or U13049 (N_13049,N_10527,N_11668);
nand U13050 (N_13050,N_10671,N_11104);
or U13051 (N_13051,N_11681,N_11143);
and U13052 (N_13052,N_10987,N_11112);
or U13053 (N_13053,N_10975,N_11198);
or U13054 (N_13054,N_11353,N_11253);
nor U13055 (N_13055,N_11041,N_11779);
or U13056 (N_13056,N_11194,N_11825);
nor U13057 (N_13057,N_10858,N_11192);
nand U13058 (N_13058,N_11755,N_11711);
nor U13059 (N_13059,N_11429,N_11469);
nor U13060 (N_13060,N_11868,N_11566);
and U13061 (N_13061,N_11688,N_11961);
and U13062 (N_13062,N_11860,N_10898);
and U13063 (N_13063,N_11263,N_11902);
or U13064 (N_13064,N_11025,N_11674);
nor U13065 (N_13065,N_10807,N_10604);
or U13066 (N_13066,N_11012,N_11089);
or U13067 (N_13067,N_11540,N_10942);
nand U13068 (N_13068,N_10853,N_10711);
nand U13069 (N_13069,N_10973,N_11477);
nand U13070 (N_13070,N_11173,N_11915);
nor U13071 (N_13071,N_11012,N_11412);
or U13072 (N_13072,N_11459,N_10825);
or U13073 (N_13073,N_10994,N_10568);
nand U13074 (N_13074,N_11304,N_11629);
nand U13075 (N_13075,N_10507,N_10713);
nor U13076 (N_13076,N_11870,N_10784);
nor U13077 (N_13077,N_11614,N_11169);
nor U13078 (N_13078,N_10758,N_11382);
and U13079 (N_13079,N_11066,N_10939);
or U13080 (N_13080,N_10947,N_10671);
or U13081 (N_13081,N_11876,N_10628);
or U13082 (N_13082,N_11337,N_11809);
or U13083 (N_13083,N_10806,N_10772);
or U13084 (N_13084,N_11285,N_10687);
and U13085 (N_13085,N_11468,N_11903);
nand U13086 (N_13086,N_11742,N_10556);
nor U13087 (N_13087,N_11094,N_10636);
nor U13088 (N_13088,N_11743,N_10598);
nand U13089 (N_13089,N_11555,N_11514);
nand U13090 (N_13090,N_11627,N_11234);
or U13091 (N_13091,N_11157,N_11635);
nor U13092 (N_13092,N_10530,N_11045);
or U13093 (N_13093,N_10685,N_11327);
nor U13094 (N_13094,N_10631,N_11184);
or U13095 (N_13095,N_11907,N_11699);
and U13096 (N_13096,N_11927,N_11373);
nor U13097 (N_13097,N_11749,N_10698);
and U13098 (N_13098,N_11292,N_10671);
or U13099 (N_13099,N_11020,N_11318);
nor U13100 (N_13100,N_11625,N_11941);
nor U13101 (N_13101,N_11054,N_10729);
nor U13102 (N_13102,N_10604,N_11406);
and U13103 (N_13103,N_11822,N_11588);
nand U13104 (N_13104,N_11866,N_11513);
nor U13105 (N_13105,N_11790,N_11400);
or U13106 (N_13106,N_10971,N_10979);
nand U13107 (N_13107,N_11245,N_10782);
nand U13108 (N_13108,N_10909,N_10852);
nand U13109 (N_13109,N_11616,N_11396);
or U13110 (N_13110,N_10828,N_11993);
nand U13111 (N_13111,N_11075,N_10735);
and U13112 (N_13112,N_11633,N_11182);
and U13113 (N_13113,N_10720,N_11326);
and U13114 (N_13114,N_10732,N_10799);
and U13115 (N_13115,N_10692,N_11907);
or U13116 (N_13116,N_11238,N_10679);
nor U13117 (N_13117,N_11202,N_10966);
or U13118 (N_13118,N_11850,N_10635);
nor U13119 (N_13119,N_11029,N_10859);
nand U13120 (N_13120,N_11650,N_10992);
nor U13121 (N_13121,N_11938,N_11906);
and U13122 (N_13122,N_10779,N_10679);
or U13123 (N_13123,N_11800,N_10871);
or U13124 (N_13124,N_11800,N_11943);
and U13125 (N_13125,N_10723,N_11563);
and U13126 (N_13126,N_11825,N_11331);
nand U13127 (N_13127,N_11025,N_11798);
or U13128 (N_13128,N_10898,N_11066);
nor U13129 (N_13129,N_10764,N_10724);
nor U13130 (N_13130,N_11739,N_10910);
and U13131 (N_13131,N_11409,N_11944);
nor U13132 (N_13132,N_11665,N_11492);
or U13133 (N_13133,N_11191,N_10711);
nand U13134 (N_13134,N_10925,N_10740);
nor U13135 (N_13135,N_10754,N_11438);
nand U13136 (N_13136,N_10977,N_10606);
nor U13137 (N_13137,N_11516,N_11970);
or U13138 (N_13138,N_11920,N_11900);
and U13139 (N_13139,N_11212,N_11083);
nor U13140 (N_13140,N_10753,N_11208);
nand U13141 (N_13141,N_11936,N_11396);
nor U13142 (N_13142,N_11079,N_11721);
or U13143 (N_13143,N_11888,N_11043);
nand U13144 (N_13144,N_11428,N_10925);
xor U13145 (N_13145,N_11594,N_11660);
nand U13146 (N_13146,N_10693,N_10539);
nor U13147 (N_13147,N_10597,N_11782);
and U13148 (N_13148,N_10717,N_11726);
nand U13149 (N_13149,N_10701,N_11490);
xnor U13150 (N_13150,N_10916,N_11276);
nor U13151 (N_13151,N_11673,N_11599);
nor U13152 (N_13152,N_11825,N_10855);
nor U13153 (N_13153,N_10505,N_10974);
and U13154 (N_13154,N_10622,N_11379);
nor U13155 (N_13155,N_11013,N_11748);
nor U13156 (N_13156,N_11241,N_10654);
nor U13157 (N_13157,N_11730,N_11314);
nor U13158 (N_13158,N_11795,N_11905);
and U13159 (N_13159,N_11748,N_11993);
and U13160 (N_13160,N_11741,N_11033);
or U13161 (N_13161,N_10907,N_10960);
nand U13162 (N_13162,N_11061,N_11017);
or U13163 (N_13163,N_11379,N_11620);
and U13164 (N_13164,N_11205,N_10594);
nand U13165 (N_13165,N_11517,N_11689);
nor U13166 (N_13166,N_10510,N_11214);
and U13167 (N_13167,N_11447,N_11858);
and U13168 (N_13168,N_10714,N_11651);
or U13169 (N_13169,N_11416,N_11187);
nor U13170 (N_13170,N_10940,N_10723);
nand U13171 (N_13171,N_10584,N_11676);
or U13172 (N_13172,N_11345,N_11447);
and U13173 (N_13173,N_10590,N_11217);
and U13174 (N_13174,N_11026,N_11968);
nor U13175 (N_13175,N_11655,N_11644);
nor U13176 (N_13176,N_11088,N_10743);
or U13177 (N_13177,N_11089,N_11346);
nand U13178 (N_13178,N_11150,N_10771);
nor U13179 (N_13179,N_11719,N_10997);
or U13180 (N_13180,N_11598,N_11121);
or U13181 (N_13181,N_10572,N_11640);
or U13182 (N_13182,N_11627,N_10709);
nor U13183 (N_13183,N_10640,N_11514);
nor U13184 (N_13184,N_11581,N_11795);
nand U13185 (N_13185,N_11789,N_11525);
nand U13186 (N_13186,N_11496,N_11696);
and U13187 (N_13187,N_11160,N_11999);
xnor U13188 (N_13188,N_11479,N_11421);
or U13189 (N_13189,N_10760,N_10928);
or U13190 (N_13190,N_10622,N_10660);
or U13191 (N_13191,N_11577,N_10661);
nand U13192 (N_13192,N_11363,N_11838);
or U13193 (N_13193,N_10626,N_11223);
nand U13194 (N_13194,N_11703,N_10762);
nor U13195 (N_13195,N_11437,N_11448);
and U13196 (N_13196,N_11226,N_11842);
nand U13197 (N_13197,N_11475,N_11678);
nand U13198 (N_13198,N_10660,N_10818);
or U13199 (N_13199,N_11112,N_11660);
and U13200 (N_13200,N_11960,N_11204);
or U13201 (N_13201,N_11233,N_11155);
or U13202 (N_13202,N_10786,N_11616);
nor U13203 (N_13203,N_11621,N_11434);
or U13204 (N_13204,N_11324,N_11903);
and U13205 (N_13205,N_11423,N_11068);
and U13206 (N_13206,N_10972,N_11372);
nand U13207 (N_13207,N_11673,N_10579);
nor U13208 (N_13208,N_11993,N_11323);
and U13209 (N_13209,N_11503,N_11683);
nor U13210 (N_13210,N_11410,N_10809);
or U13211 (N_13211,N_11816,N_11583);
or U13212 (N_13212,N_10887,N_10532);
and U13213 (N_13213,N_11497,N_10819);
nor U13214 (N_13214,N_10958,N_11863);
and U13215 (N_13215,N_11563,N_10535);
nor U13216 (N_13216,N_11075,N_11726);
nand U13217 (N_13217,N_11266,N_10924);
and U13218 (N_13218,N_10995,N_10865);
nand U13219 (N_13219,N_11397,N_11161);
or U13220 (N_13220,N_11150,N_11055);
nor U13221 (N_13221,N_10912,N_10852);
nor U13222 (N_13222,N_10555,N_11431);
and U13223 (N_13223,N_11185,N_10980);
and U13224 (N_13224,N_11074,N_11136);
and U13225 (N_13225,N_10691,N_11516);
nand U13226 (N_13226,N_10892,N_10857);
or U13227 (N_13227,N_10506,N_11369);
or U13228 (N_13228,N_11887,N_10938);
nand U13229 (N_13229,N_11781,N_11316);
nor U13230 (N_13230,N_11030,N_11881);
and U13231 (N_13231,N_11579,N_11985);
and U13232 (N_13232,N_10756,N_11457);
or U13233 (N_13233,N_11994,N_11889);
or U13234 (N_13234,N_11377,N_11470);
nor U13235 (N_13235,N_11872,N_11438);
nand U13236 (N_13236,N_11488,N_10632);
nor U13237 (N_13237,N_10906,N_11284);
and U13238 (N_13238,N_11472,N_11851);
and U13239 (N_13239,N_11804,N_11350);
or U13240 (N_13240,N_10761,N_11289);
nor U13241 (N_13241,N_11179,N_11001);
nor U13242 (N_13242,N_11661,N_11461);
nor U13243 (N_13243,N_10740,N_11695);
nand U13244 (N_13244,N_10983,N_10731);
and U13245 (N_13245,N_11092,N_11660);
nand U13246 (N_13246,N_10628,N_11359);
or U13247 (N_13247,N_10682,N_11063);
or U13248 (N_13248,N_11272,N_11564);
nand U13249 (N_13249,N_10540,N_11610);
xnor U13250 (N_13250,N_11144,N_11040);
nand U13251 (N_13251,N_11372,N_11173);
and U13252 (N_13252,N_10935,N_10555);
nor U13253 (N_13253,N_11934,N_10979);
and U13254 (N_13254,N_11793,N_11027);
nand U13255 (N_13255,N_11061,N_11863);
nor U13256 (N_13256,N_11660,N_11995);
nand U13257 (N_13257,N_11626,N_11614);
nor U13258 (N_13258,N_10660,N_10885);
nand U13259 (N_13259,N_11992,N_10686);
nor U13260 (N_13260,N_11807,N_10563);
nand U13261 (N_13261,N_11863,N_11081);
and U13262 (N_13262,N_11798,N_11689);
and U13263 (N_13263,N_10503,N_10661);
nor U13264 (N_13264,N_11954,N_11071);
nor U13265 (N_13265,N_11106,N_11864);
nand U13266 (N_13266,N_10785,N_11337);
nor U13267 (N_13267,N_10614,N_10769);
or U13268 (N_13268,N_11690,N_11346);
and U13269 (N_13269,N_11396,N_11280);
and U13270 (N_13270,N_10762,N_10791);
nand U13271 (N_13271,N_11837,N_11003);
or U13272 (N_13272,N_10864,N_11765);
nand U13273 (N_13273,N_11346,N_11768);
nor U13274 (N_13274,N_10811,N_11692);
and U13275 (N_13275,N_11062,N_10836);
or U13276 (N_13276,N_11901,N_10948);
nand U13277 (N_13277,N_10852,N_11491);
nor U13278 (N_13278,N_11100,N_11028);
nand U13279 (N_13279,N_11722,N_10886);
and U13280 (N_13280,N_11446,N_11972);
or U13281 (N_13281,N_11791,N_11366);
and U13282 (N_13282,N_11038,N_11172);
and U13283 (N_13283,N_11336,N_11996);
nand U13284 (N_13284,N_10954,N_11214);
nand U13285 (N_13285,N_11368,N_10923);
and U13286 (N_13286,N_11236,N_10663);
or U13287 (N_13287,N_11541,N_10897);
and U13288 (N_13288,N_11110,N_11497);
nand U13289 (N_13289,N_11668,N_10939);
or U13290 (N_13290,N_10866,N_10824);
and U13291 (N_13291,N_10733,N_11543);
and U13292 (N_13292,N_11200,N_11000);
nand U13293 (N_13293,N_10937,N_11520);
and U13294 (N_13294,N_11340,N_11365);
nor U13295 (N_13295,N_11007,N_11416);
and U13296 (N_13296,N_11283,N_11876);
and U13297 (N_13297,N_11838,N_11077);
nand U13298 (N_13298,N_10895,N_10745);
nand U13299 (N_13299,N_10889,N_11242);
or U13300 (N_13300,N_11344,N_11193);
or U13301 (N_13301,N_11429,N_10571);
nor U13302 (N_13302,N_11948,N_11977);
nand U13303 (N_13303,N_11088,N_11583);
and U13304 (N_13304,N_11093,N_11383);
nor U13305 (N_13305,N_11058,N_10911);
nor U13306 (N_13306,N_11796,N_10792);
nand U13307 (N_13307,N_10516,N_11042);
nand U13308 (N_13308,N_10826,N_10977);
or U13309 (N_13309,N_11963,N_10761);
or U13310 (N_13310,N_11933,N_10941);
nor U13311 (N_13311,N_11652,N_11761);
nor U13312 (N_13312,N_10863,N_11486);
or U13313 (N_13313,N_10574,N_10898);
and U13314 (N_13314,N_11747,N_11157);
or U13315 (N_13315,N_11546,N_10743);
nand U13316 (N_13316,N_11265,N_11900);
and U13317 (N_13317,N_11210,N_11168);
and U13318 (N_13318,N_11337,N_11161);
nor U13319 (N_13319,N_11468,N_11754);
nand U13320 (N_13320,N_10646,N_11310);
and U13321 (N_13321,N_10979,N_10903);
or U13322 (N_13322,N_10599,N_10857);
or U13323 (N_13323,N_10822,N_11856);
or U13324 (N_13324,N_10851,N_11151);
nand U13325 (N_13325,N_11345,N_11744);
and U13326 (N_13326,N_10978,N_11999);
and U13327 (N_13327,N_11789,N_11538);
or U13328 (N_13328,N_10993,N_11197);
nand U13329 (N_13329,N_11101,N_11851);
and U13330 (N_13330,N_10636,N_10664);
nor U13331 (N_13331,N_11607,N_11821);
and U13332 (N_13332,N_11797,N_11612);
nand U13333 (N_13333,N_10622,N_11806);
nor U13334 (N_13334,N_10599,N_11894);
or U13335 (N_13335,N_11538,N_11191);
nand U13336 (N_13336,N_11733,N_11664);
or U13337 (N_13337,N_10648,N_11078);
or U13338 (N_13338,N_10922,N_11669);
xor U13339 (N_13339,N_11069,N_10725);
nor U13340 (N_13340,N_10726,N_11060);
or U13341 (N_13341,N_10868,N_11880);
and U13342 (N_13342,N_11854,N_10780);
or U13343 (N_13343,N_11574,N_11706);
and U13344 (N_13344,N_11773,N_11231);
or U13345 (N_13345,N_11867,N_11745);
or U13346 (N_13346,N_11612,N_11819);
nor U13347 (N_13347,N_11325,N_11343);
or U13348 (N_13348,N_10714,N_10556);
nand U13349 (N_13349,N_11437,N_10744);
or U13350 (N_13350,N_10930,N_11530);
nor U13351 (N_13351,N_10534,N_11125);
nand U13352 (N_13352,N_10903,N_11351);
and U13353 (N_13353,N_11561,N_11762);
or U13354 (N_13354,N_11029,N_11054);
nor U13355 (N_13355,N_11825,N_10967);
nand U13356 (N_13356,N_11157,N_11449);
or U13357 (N_13357,N_11087,N_11401);
nand U13358 (N_13358,N_11947,N_11970);
and U13359 (N_13359,N_11110,N_10954);
nor U13360 (N_13360,N_11636,N_11270);
and U13361 (N_13361,N_10897,N_11247);
or U13362 (N_13362,N_10953,N_11358);
nand U13363 (N_13363,N_10929,N_11117);
and U13364 (N_13364,N_10570,N_10538);
and U13365 (N_13365,N_11253,N_10755);
nand U13366 (N_13366,N_11566,N_11310);
nor U13367 (N_13367,N_11876,N_11183);
nand U13368 (N_13368,N_11183,N_11920);
and U13369 (N_13369,N_10853,N_11180);
nor U13370 (N_13370,N_10688,N_11856);
nor U13371 (N_13371,N_11994,N_11960);
nor U13372 (N_13372,N_10839,N_11361);
and U13373 (N_13373,N_11883,N_11185);
and U13374 (N_13374,N_10879,N_11844);
or U13375 (N_13375,N_11179,N_10949);
nand U13376 (N_13376,N_11837,N_10742);
and U13377 (N_13377,N_10556,N_11695);
or U13378 (N_13378,N_10841,N_10668);
nor U13379 (N_13379,N_11195,N_11786);
nand U13380 (N_13380,N_11453,N_11671);
or U13381 (N_13381,N_11364,N_11420);
or U13382 (N_13382,N_11739,N_11110);
and U13383 (N_13383,N_10921,N_10989);
or U13384 (N_13384,N_11476,N_11998);
nor U13385 (N_13385,N_11472,N_11215);
or U13386 (N_13386,N_11380,N_11930);
nor U13387 (N_13387,N_10787,N_10863);
or U13388 (N_13388,N_11980,N_11973);
nand U13389 (N_13389,N_10850,N_11091);
nor U13390 (N_13390,N_10709,N_11535);
and U13391 (N_13391,N_10877,N_11138);
nor U13392 (N_13392,N_11792,N_11905);
or U13393 (N_13393,N_11104,N_11150);
nor U13394 (N_13394,N_11990,N_11270);
nand U13395 (N_13395,N_11840,N_11231);
nand U13396 (N_13396,N_11179,N_11497);
nand U13397 (N_13397,N_10666,N_11723);
and U13398 (N_13398,N_11787,N_11202);
and U13399 (N_13399,N_10696,N_11354);
and U13400 (N_13400,N_11591,N_11945);
nor U13401 (N_13401,N_11913,N_11677);
nor U13402 (N_13402,N_11106,N_11288);
xnor U13403 (N_13403,N_10500,N_10855);
nor U13404 (N_13404,N_11291,N_11660);
or U13405 (N_13405,N_11141,N_11532);
and U13406 (N_13406,N_11067,N_10827);
nand U13407 (N_13407,N_10783,N_11558);
or U13408 (N_13408,N_11848,N_11341);
nand U13409 (N_13409,N_11893,N_11079);
nor U13410 (N_13410,N_10542,N_11886);
nand U13411 (N_13411,N_10739,N_11360);
or U13412 (N_13412,N_10759,N_11316);
and U13413 (N_13413,N_10514,N_10670);
and U13414 (N_13414,N_11605,N_10852);
nor U13415 (N_13415,N_11077,N_11904);
nor U13416 (N_13416,N_10735,N_10602);
and U13417 (N_13417,N_10819,N_11391);
nor U13418 (N_13418,N_10706,N_11273);
or U13419 (N_13419,N_11163,N_11386);
and U13420 (N_13420,N_10553,N_11090);
nor U13421 (N_13421,N_11699,N_10797);
nor U13422 (N_13422,N_11399,N_11468);
nor U13423 (N_13423,N_11240,N_11591);
and U13424 (N_13424,N_11672,N_11682);
nand U13425 (N_13425,N_10762,N_11610);
nor U13426 (N_13426,N_10829,N_11903);
and U13427 (N_13427,N_11086,N_10692);
nand U13428 (N_13428,N_10810,N_10926);
xnor U13429 (N_13429,N_11489,N_11279);
and U13430 (N_13430,N_10563,N_11932);
and U13431 (N_13431,N_11027,N_11619);
xnor U13432 (N_13432,N_11574,N_10907);
nand U13433 (N_13433,N_10678,N_11207);
nor U13434 (N_13434,N_11793,N_11006);
or U13435 (N_13435,N_10908,N_11186);
nand U13436 (N_13436,N_11914,N_10822);
nor U13437 (N_13437,N_10739,N_11740);
and U13438 (N_13438,N_11447,N_11026);
or U13439 (N_13439,N_10837,N_11937);
nand U13440 (N_13440,N_10542,N_10872);
nand U13441 (N_13441,N_10803,N_11240);
or U13442 (N_13442,N_11116,N_11342);
nand U13443 (N_13443,N_11784,N_10532);
nor U13444 (N_13444,N_11069,N_11375);
nor U13445 (N_13445,N_11633,N_11236);
nor U13446 (N_13446,N_10982,N_10966);
nor U13447 (N_13447,N_10572,N_11826);
nand U13448 (N_13448,N_10918,N_11508);
nand U13449 (N_13449,N_10603,N_11844);
nor U13450 (N_13450,N_11729,N_11858);
nor U13451 (N_13451,N_11522,N_10734);
or U13452 (N_13452,N_11931,N_11213);
nor U13453 (N_13453,N_11838,N_10798);
or U13454 (N_13454,N_11254,N_11969);
and U13455 (N_13455,N_11888,N_10659);
nor U13456 (N_13456,N_11264,N_11646);
nor U13457 (N_13457,N_10879,N_10963);
nor U13458 (N_13458,N_10982,N_11735);
nor U13459 (N_13459,N_11324,N_11442);
nand U13460 (N_13460,N_11359,N_11783);
nand U13461 (N_13461,N_10945,N_11904);
or U13462 (N_13462,N_11813,N_10625);
and U13463 (N_13463,N_11426,N_11608);
or U13464 (N_13464,N_11290,N_10840);
nand U13465 (N_13465,N_10771,N_11645);
and U13466 (N_13466,N_11566,N_11528);
nand U13467 (N_13467,N_10890,N_11373);
nor U13468 (N_13468,N_10826,N_11191);
nand U13469 (N_13469,N_10759,N_11921);
and U13470 (N_13470,N_11159,N_11682);
nor U13471 (N_13471,N_10932,N_10939);
nor U13472 (N_13472,N_11307,N_10537);
and U13473 (N_13473,N_11067,N_10544);
nand U13474 (N_13474,N_10799,N_11152);
nor U13475 (N_13475,N_11813,N_10960);
or U13476 (N_13476,N_11607,N_10592);
and U13477 (N_13477,N_11457,N_10829);
nor U13478 (N_13478,N_11056,N_10583);
and U13479 (N_13479,N_11194,N_11604);
and U13480 (N_13480,N_11504,N_11496);
and U13481 (N_13481,N_11720,N_11741);
nor U13482 (N_13482,N_10536,N_11570);
xnor U13483 (N_13483,N_11539,N_10684);
and U13484 (N_13484,N_11498,N_10645);
or U13485 (N_13485,N_11510,N_11901);
nand U13486 (N_13486,N_11779,N_11907);
or U13487 (N_13487,N_10511,N_11364);
and U13488 (N_13488,N_11879,N_11882);
nor U13489 (N_13489,N_11116,N_11268);
nand U13490 (N_13490,N_11367,N_10946);
nor U13491 (N_13491,N_11059,N_11495);
nand U13492 (N_13492,N_10663,N_11676);
or U13493 (N_13493,N_10692,N_11817);
nand U13494 (N_13494,N_11121,N_10883);
and U13495 (N_13495,N_11579,N_11912);
and U13496 (N_13496,N_11051,N_11750);
and U13497 (N_13497,N_11294,N_11395);
nor U13498 (N_13498,N_10578,N_11940);
nand U13499 (N_13499,N_11052,N_11144);
nor U13500 (N_13500,N_12787,N_13178);
and U13501 (N_13501,N_12033,N_13195);
and U13502 (N_13502,N_12455,N_12139);
or U13503 (N_13503,N_12107,N_12793);
or U13504 (N_13504,N_13437,N_13462);
or U13505 (N_13505,N_12443,N_12045);
nor U13506 (N_13506,N_12598,N_12270);
and U13507 (N_13507,N_12495,N_13340);
or U13508 (N_13508,N_12095,N_12730);
and U13509 (N_13509,N_13423,N_12281);
nor U13510 (N_13510,N_13339,N_12723);
nor U13511 (N_13511,N_13306,N_13447);
nand U13512 (N_13512,N_13264,N_13409);
xor U13513 (N_13513,N_12459,N_12397);
and U13514 (N_13514,N_13427,N_12812);
and U13515 (N_13515,N_13267,N_12437);
and U13516 (N_13516,N_12530,N_13002);
nand U13517 (N_13517,N_12317,N_13023);
or U13518 (N_13518,N_12616,N_12451);
and U13519 (N_13519,N_12359,N_13068);
and U13520 (N_13520,N_13345,N_12135);
and U13521 (N_13521,N_12828,N_12626);
or U13522 (N_13522,N_12020,N_12168);
nor U13523 (N_13523,N_12146,N_12234);
or U13524 (N_13524,N_13280,N_12917);
nand U13525 (N_13525,N_13472,N_12386);
nor U13526 (N_13526,N_13136,N_12357);
or U13527 (N_13527,N_12923,N_12804);
or U13528 (N_13528,N_13322,N_12946);
and U13529 (N_13529,N_12779,N_12861);
or U13530 (N_13530,N_13343,N_13457);
or U13531 (N_13531,N_12452,N_13065);
and U13532 (N_13532,N_12218,N_13269);
or U13533 (N_13533,N_12873,N_13405);
and U13534 (N_13534,N_12585,N_13109);
or U13535 (N_13535,N_12278,N_13238);
nand U13536 (N_13536,N_12065,N_12192);
nand U13537 (N_13537,N_12915,N_12128);
nor U13538 (N_13538,N_12658,N_13055);
nor U13539 (N_13539,N_12739,N_13126);
and U13540 (N_13540,N_13358,N_12433);
nor U13541 (N_13541,N_12737,N_13144);
and U13542 (N_13542,N_12389,N_12345);
nand U13543 (N_13543,N_12222,N_12843);
or U13544 (N_13544,N_12354,N_13402);
and U13545 (N_13545,N_12963,N_12333);
or U13546 (N_13546,N_12235,N_12629);
and U13547 (N_13547,N_12034,N_12327);
and U13548 (N_13548,N_12975,N_12987);
nand U13549 (N_13549,N_12978,N_12889);
nand U13550 (N_13550,N_12456,N_12693);
nand U13551 (N_13551,N_13478,N_12162);
or U13552 (N_13552,N_12047,N_12927);
and U13553 (N_13553,N_12605,N_13040);
nor U13554 (N_13554,N_13170,N_12838);
and U13555 (N_13555,N_13367,N_12201);
nand U13556 (N_13556,N_12157,N_12290);
and U13557 (N_13557,N_13203,N_13008);
nor U13558 (N_13558,N_12934,N_12972);
xnor U13559 (N_13559,N_12367,N_12332);
nand U13560 (N_13560,N_12628,N_13207);
nand U13561 (N_13561,N_12876,N_12574);
nor U13562 (N_13562,N_13298,N_13141);
or U13563 (N_13563,N_12249,N_12104);
nor U13564 (N_13564,N_12092,N_12618);
nand U13565 (N_13565,N_13095,N_13487);
nand U13566 (N_13566,N_13096,N_12719);
or U13567 (N_13567,N_12085,N_12758);
nand U13568 (N_13568,N_13027,N_13153);
or U13569 (N_13569,N_12712,N_13110);
nor U13570 (N_13570,N_12622,N_12973);
nor U13571 (N_13571,N_12394,N_12700);
nor U13572 (N_13572,N_13154,N_13300);
and U13573 (N_13573,N_13104,N_12111);
nand U13574 (N_13574,N_12297,N_12038);
and U13575 (N_13575,N_12884,N_12143);
nor U13576 (N_13576,N_12043,N_12477);
and U13577 (N_13577,N_12924,N_13060);
or U13578 (N_13578,N_12362,N_13081);
or U13579 (N_13579,N_12767,N_13274);
or U13580 (N_13580,N_12421,N_12959);
nand U13581 (N_13581,N_13440,N_13128);
and U13582 (N_13582,N_12687,N_12048);
nor U13583 (N_13583,N_12307,N_13341);
and U13584 (N_13584,N_12424,N_12287);
or U13585 (N_13585,N_12770,N_13059);
and U13586 (N_13586,N_13281,N_12053);
nand U13587 (N_13587,N_12331,N_13385);
or U13588 (N_13588,N_12961,N_12590);
nand U13589 (N_13589,N_13448,N_12244);
or U13590 (N_13590,N_12405,N_13377);
nand U13591 (N_13591,N_12060,N_12503);
and U13592 (N_13592,N_13276,N_12832);
nor U13593 (N_13593,N_12600,N_12059);
and U13594 (N_13594,N_12565,N_12588);
or U13595 (N_13595,N_13185,N_13466);
or U13596 (N_13596,N_12229,N_13268);
nand U13597 (N_13597,N_12520,N_13296);
or U13598 (N_13598,N_12369,N_12734);
nand U13599 (N_13599,N_12123,N_12254);
and U13600 (N_13600,N_13356,N_12831);
nand U13601 (N_13601,N_13025,N_12497);
nand U13602 (N_13602,N_12606,N_13217);
and U13603 (N_13603,N_13482,N_13188);
nor U13604 (N_13604,N_12458,N_12300);
nand U13605 (N_13605,N_12089,N_13214);
nor U13606 (N_13606,N_12350,N_13278);
and U13607 (N_13607,N_12099,N_12240);
nor U13608 (N_13608,N_13132,N_13253);
or U13609 (N_13609,N_13432,N_12990);
nor U13610 (N_13610,N_12132,N_12093);
and U13611 (N_13611,N_12129,N_12356);
nor U13612 (N_13612,N_12119,N_13176);
nand U13613 (N_13613,N_12877,N_13140);
nand U13614 (N_13614,N_13378,N_12248);
nor U13615 (N_13615,N_13460,N_12875);
and U13616 (N_13616,N_13493,N_12371);
and U13617 (N_13617,N_12390,N_13229);
or U13618 (N_13618,N_12088,N_12196);
nand U13619 (N_13619,N_13164,N_13393);
nand U13620 (N_13620,N_12262,N_12989);
and U13621 (N_13621,N_12220,N_12153);
nor U13622 (N_13622,N_12524,N_13082);
nand U13623 (N_13623,N_13221,N_13445);
nor U13624 (N_13624,N_13388,N_12611);
nand U13625 (N_13625,N_12860,N_13312);
nor U13626 (N_13626,N_13106,N_12736);
xnor U13627 (N_13627,N_13004,N_13183);
and U13628 (N_13628,N_12098,N_12136);
and U13629 (N_13629,N_13206,N_12049);
and U13630 (N_13630,N_12462,N_12137);
or U13631 (N_13631,N_12032,N_12316);
nand U13632 (N_13632,N_12880,N_12149);
nand U13633 (N_13633,N_12003,N_12492);
nor U13634 (N_13634,N_12985,N_12695);
nand U13635 (N_13635,N_13254,N_13215);
xor U13636 (N_13636,N_12822,N_12453);
or U13637 (N_13637,N_12133,N_13193);
and U13638 (N_13638,N_13028,N_13381);
nand U13639 (N_13639,N_12579,N_12246);
and U13640 (N_13640,N_12182,N_12580);
and U13641 (N_13641,N_12778,N_12226);
and U13642 (N_13642,N_13467,N_12722);
nor U13643 (N_13643,N_12050,N_12555);
nor U13644 (N_13644,N_12352,N_13320);
and U13645 (N_13645,N_12475,N_13047);
nand U13646 (N_13646,N_12856,N_13205);
or U13647 (N_13647,N_12745,N_13013);
or U13648 (N_13648,N_12465,N_12378);
or U13649 (N_13649,N_12466,N_12215);
or U13650 (N_13650,N_13498,N_12183);
nor U13651 (N_13651,N_12620,N_12148);
nor U13652 (N_13652,N_12957,N_12850);
nand U13653 (N_13653,N_13048,N_12061);
nor U13654 (N_13654,N_12663,N_12268);
or U13655 (N_13655,N_12733,N_13014);
nand U13656 (N_13656,N_13124,N_12273);
nor U13657 (N_13657,N_12691,N_12072);
nor U13658 (N_13658,N_12340,N_12926);
or U13659 (N_13659,N_13228,N_12920);
nand U13660 (N_13660,N_13160,N_12334);
and U13661 (N_13661,N_12062,N_12160);
nor U13662 (N_13662,N_12170,N_13067);
and U13663 (N_13663,N_12147,N_12392);
nor U13664 (N_13664,N_12493,N_13441);
or U13665 (N_13665,N_13012,N_13087);
nand U13666 (N_13666,N_12057,N_13252);
and U13667 (N_13667,N_12950,N_13000);
and U13668 (N_13668,N_12193,N_13194);
nand U13669 (N_13669,N_12208,N_13456);
or U13670 (N_13670,N_13469,N_13330);
or U13671 (N_13671,N_12223,N_13387);
and U13672 (N_13672,N_12991,N_12699);
nor U13673 (N_13673,N_12621,N_12266);
nand U13674 (N_13674,N_12964,N_12771);
nor U13675 (N_13675,N_12158,N_12083);
and U13676 (N_13676,N_12250,N_13054);
and U13677 (N_13677,N_12772,N_12374);
xor U13678 (N_13678,N_12603,N_12538);
and U13679 (N_13679,N_13138,N_12021);
and U13680 (N_13680,N_12644,N_12916);
nand U13681 (N_13681,N_12097,N_12776);
and U13682 (N_13682,N_12472,N_13116);
nand U13683 (N_13683,N_12159,N_13332);
or U13684 (N_13684,N_12597,N_13061);
and U13685 (N_13685,N_12432,N_12754);
nand U13686 (N_13686,N_12905,N_12656);
nand U13687 (N_13687,N_13291,N_12680);
nand U13688 (N_13688,N_12797,N_12411);
or U13689 (N_13689,N_12649,N_12842);
nand U13690 (N_13690,N_12635,N_12706);
nor U13691 (N_13691,N_12030,N_13303);
or U13692 (N_13692,N_12785,N_12702);
and U13693 (N_13693,N_13352,N_12756);
nand U13694 (N_13694,N_12602,N_12631);
xnor U13695 (N_13695,N_12904,N_13213);
nand U13696 (N_13696,N_12557,N_12848);
and U13697 (N_13697,N_12811,N_13090);
and U13698 (N_13698,N_12398,N_12716);
or U13699 (N_13699,N_13108,N_12871);
nand U13700 (N_13700,N_12217,N_12903);
nor U13701 (N_13701,N_12750,N_12866);
or U13702 (N_13702,N_13244,N_12552);
nor U13703 (N_13703,N_12295,N_12006);
and U13704 (N_13704,N_12988,N_12084);
nor U13705 (N_13705,N_13143,N_12541);
nor U13706 (N_13706,N_12931,N_13318);
or U13707 (N_13707,N_12485,N_12079);
nand U13708 (N_13708,N_12642,N_12741);
nand U13709 (N_13709,N_13382,N_13145);
nand U13710 (N_13710,N_13302,N_12806);
or U13711 (N_13711,N_12522,N_12315);
nor U13712 (N_13712,N_12526,N_12319);
or U13713 (N_13713,N_12001,N_12766);
nor U13714 (N_13714,N_13473,N_12419);
or U13715 (N_13715,N_12849,N_12696);
or U13716 (N_13716,N_12803,N_13257);
nand U13717 (N_13717,N_12948,N_12156);
or U13718 (N_13718,N_12109,N_12259);
and U13719 (N_13719,N_12569,N_12054);
or U13720 (N_13720,N_12939,N_13459);
nor U13721 (N_13721,N_12929,N_12018);
and U13722 (N_13722,N_12535,N_12800);
nand U13723 (N_13723,N_12118,N_12910);
nor U13724 (N_13724,N_13271,N_12301);
and U13725 (N_13725,N_12376,N_12527);
nor U13726 (N_13726,N_12174,N_12824);
or U13727 (N_13727,N_12799,N_12761);
and U13728 (N_13728,N_12531,N_12066);
or U13729 (N_13729,N_13050,N_13497);
or U13730 (N_13730,N_13197,N_12124);
nand U13731 (N_13731,N_13184,N_12480);
nor U13732 (N_13732,N_13121,N_12979);
nand U13733 (N_13733,N_12499,N_12036);
and U13734 (N_13734,N_12473,N_13314);
nand U13735 (N_13735,N_13286,N_12593);
nor U13736 (N_13736,N_13255,N_13098);
nand U13737 (N_13737,N_12496,N_12909);
or U13738 (N_13738,N_13173,N_12388);
nand U13739 (N_13739,N_13245,N_12257);
or U13740 (N_13740,N_13035,N_12847);
nand U13741 (N_13741,N_13389,N_12130);
and U13742 (N_13742,N_13074,N_12063);
and U13743 (N_13743,N_12589,N_13349);
or U13744 (N_13744,N_12373,N_13461);
or U13745 (N_13745,N_12969,N_12511);
and U13746 (N_13746,N_12363,N_13401);
or U13747 (N_13747,N_12074,N_12450);
nor U13748 (N_13748,N_12955,N_13411);
or U13749 (N_13749,N_12228,N_13250);
or U13750 (N_13750,N_12841,N_12942);
or U13751 (N_13751,N_12339,N_12467);
and U13752 (N_13752,N_13416,N_13248);
nand U13753 (N_13753,N_13293,N_12186);
and U13754 (N_13754,N_12711,N_12925);
nand U13755 (N_13755,N_12851,N_12484);
or U13756 (N_13756,N_13155,N_13275);
nand U13757 (N_13757,N_12474,N_13292);
and U13758 (N_13758,N_12227,N_13235);
and U13759 (N_13759,N_12654,N_13446);
or U13760 (N_13760,N_13438,N_12643);
and U13761 (N_13761,N_13357,N_12471);
nand U13762 (N_13762,N_13191,N_12670);
and U13763 (N_13763,N_12069,N_12191);
and U13764 (N_13764,N_12478,N_12500);
or U13765 (N_13765,N_12154,N_13233);
and U13766 (N_13766,N_12769,N_13125);
or U13767 (N_13767,N_12966,N_12679);
nand U13768 (N_13768,N_12864,N_12205);
and U13769 (N_13769,N_12404,N_12648);
or U13770 (N_13770,N_12528,N_13425);
nand U13771 (N_13771,N_13383,N_12343);
nor U13772 (N_13772,N_12686,N_12862);
nand U13773 (N_13773,N_12998,N_12314);
or U13774 (N_13774,N_13396,N_12540);
or U13775 (N_13775,N_12284,N_12891);
and U13776 (N_13776,N_13216,N_13371);
nand U13777 (N_13777,N_13260,N_13336);
nor U13778 (N_13778,N_12713,N_12516);
nand U13779 (N_13779,N_12140,N_12303);
nor U13780 (N_13780,N_12814,N_12683);
nand U13781 (N_13781,N_12023,N_13152);
and U13782 (N_13782,N_12650,N_13372);
nor U13783 (N_13783,N_12042,N_13316);
or U13784 (N_13784,N_12134,N_12344);
or U13785 (N_13785,N_13078,N_13403);
nor U13786 (N_13786,N_12651,N_13102);
xor U13787 (N_13787,N_12839,N_12276);
and U13788 (N_13788,N_12116,N_12409);
and U13789 (N_13789,N_12892,N_12566);
and U13790 (N_13790,N_12563,N_12090);
nand U13791 (N_13791,N_13202,N_12940);
and U13792 (N_13792,N_12040,N_13421);
nor U13793 (N_13793,N_12836,N_13100);
or U13794 (N_13794,N_12992,N_13288);
nor U13795 (N_13795,N_12641,N_13429);
nor U13796 (N_13796,N_12415,N_12429);
or U13797 (N_13797,N_13265,N_13398);
nor U13798 (N_13798,N_12922,N_12073);
nand U13799 (N_13799,N_12056,N_12935);
nor U13800 (N_13800,N_12245,N_13305);
or U13801 (N_13801,N_13272,N_13323);
nor U13802 (N_13802,N_13072,N_13365);
nor U13803 (N_13803,N_13499,N_12029);
nand U13804 (N_13804,N_12529,N_13210);
or U13805 (N_13805,N_13005,N_12692);
and U13806 (N_13806,N_13394,N_12630);
and U13807 (N_13807,N_12490,N_13212);
nand U13808 (N_13808,N_12735,N_12619);
or U13809 (N_13809,N_12640,N_12044);
or U13810 (N_13810,N_12578,N_12385);
and U13811 (N_13811,N_12690,N_12977);
nand U13812 (N_13812,N_12592,N_12852);
or U13813 (N_13813,N_12292,N_12788);
xor U13814 (N_13814,N_13444,N_12813);
and U13815 (N_13815,N_12584,N_13076);
nand U13816 (N_13816,N_13051,N_13057);
nand U13817 (N_13817,N_13430,N_12582);
nor U13818 (N_13818,N_12994,N_13259);
nand U13819 (N_13819,N_13375,N_12665);
nor U13820 (N_13820,N_12688,N_12587);
and U13821 (N_13821,N_13251,N_12945);
nor U13822 (N_13822,N_12607,N_13391);
and U13823 (N_13823,N_13166,N_13239);
or U13824 (N_13824,N_13015,N_13242);
nand U13825 (N_13825,N_12594,N_12610);
nor U13826 (N_13826,N_12308,N_13315);
and U13827 (N_13827,N_12460,N_12161);
or U13828 (N_13828,N_13410,N_12697);
and U13829 (N_13829,N_13159,N_13018);
and U13830 (N_13830,N_12285,N_12412);
or U13831 (N_13831,N_13325,N_13169);
nor U13832 (N_13832,N_12035,N_13370);
nand U13833 (N_13833,N_12764,N_13118);
or U13834 (N_13834,N_13384,N_13080);
and U13835 (N_13835,N_12731,N_13485);
nor U13836 (N_13836,N_12231,N_12199);
nor U13837 (N_13837,N_13158,N_13156);
and U13838 (N_13838,N_12324,N_12845);
nand U13839 (N_13839,N_12637,N_12322);
or U13840 (N_13840,N_12962,N_13354);
nor U13841 (N_13841,N_12982,N_13464);
nand U13842 (N_13842,N_13418,N_12907);
nor U13843 (N_13843,N_12835,N_12489);
nand U13844 (N_13844,N_13366,N_12064);
nand U13845 (N_13845,N_13465,N_12403);
nand U13846 (N_13846,N_12105,N_12560);
nand U13847 (N_13847,N_12729,N_13187);
or U13848 (N_13848,N_13168,N_12506);
nand U13849 (N_13849,N_12781,N_13246);
and U13850 (N_13850,N_12138,N_12025);
nand U13851 (N_13851,N_12189,N_13415);
and U13852 (N_13852,N_12486,N_13227);
and U13853 (N_13853,N_12202,N_13039);
or U13854 (N_13854,N_12476,N_13199);
or U13855 (N_13855,N_12689,N_13263);
nor U13856 (N_13856,N_12243,N_13105);
nand U13857 (N_13857,N_12536,N_12853);
nor U13858 (N_13858,N_12338,N_12173);
nand U13859 (N_13859,N_12625,N_12740);
and U13860 (N_13860,N_13192,N_12360);
nor U13861 (N_13861,N_12256,N_12823);
and U13862 (N_13862,N_12242,N_12913);
nand U13863 (N_13863,N_13196,N_12971);
and U13864 (N_13864,N_12177,N_12518);
nand U13865 (N_13865,N_12275,N_12328);
and U13866 (N_13866,N_13439,N_12615);
nor U13867 (N_13867,N_12559,N_12510);
or U13868 (N_13868,N_13020,N_13162);
nand U13869 (N_13869,N_13480,N_13443);
or U13870 (N_13870,N_13026,N_12011);
and U13871 (N_13871,N_12100,N_13313);
or U13872 (N_13872,N_12967,N_12523);
and U13873 (N_13873,N_12595,N_12534);
and U13874 (N_13874,N_12944,N_12009);
and U13875 (N_13875,N_12968,N_13258);
and U13876 (N_13876,N_12930,N_12941);
nor U13877 (N_13877,N_13127,N_12817);
nand U13878 (N_13878,N_13111,N_12525);
or U13879 (N_13879,N_13309,N_13030);
nand U13880 (N_13880,N_12678,N_12166);
nor U13881 (N_13881,N_12727,N_12184);
or U13882 (N_13882,N_12746,N_12422);
nand U13883 (N_13883,N_12883,N_13165);
nand U13884 (N_13884,N_12279,N_12329);
and U13885 (N_13885,N_12645,N_13119);
nor U13886 (N_13886,N_12291,N_13380);
and U13887 (N_13887,N_13204,N_13019);
or U13888 (N_13888,N_12311,N_12763);
nand U13889 (N_13889,N_12387,N_12827);
and U13890 (N_13890,N_12790,N_12002);
nor U13891 (N_13891,N_12260,N_12313);
nand U13892 (N_13892,N_13256,N_13333);
xor U13893 (N_13893,N_12881,N_12375);
or U13894 (N_13894,N_12568,N_13094);
nor U13895 (N_13895,N_12532,N_12431);
or U13896 (N_13896,N_12368,N_12464);
and U13897 (N_13897,N_13120,N_13007);
and U13898 (N_13898,N_12572,N_12694);
nand U13899 (N_13899,N_12704,N_13231);
nor U13900 (N_13900,N_12743,N_13043);
nand U13901 (N_13901,N_12914,N_12310);
or U13902 (N_13902,N_13492,N_13428);
or U13903 (N_13903,N_12608,N_12951);
nand U13904 (N_13904,N_13317,N_12238);
nor U13905 (N_13905,N_12206,N_12976);
nand U13906 (N_13906,N_13071,N_12361);
nor U13907 (N_13907,N_13045,N_13112);
or U13908 (N_13908,N_12498,N_12251);
or U13909 (N_13909,N_12720,N_13359);
nand U13910 (N_13910,N_12401,N_12647);
nor U13911 (N_13911,N_13022,N_12780);
nand U13912 (N_13912,N_13084,N_12636);
xor U13913 (N_13913,N_12479,N_13468);
nor U13914 (N_13914,N_12633,N_12171);
nand U13915 (N_13915,N_12890,N_12627);
nand U13916 (N_13916,N_12786,N_12701);
and U13917 (N_13917,N_13079,N_13001);
or U13918 (N_13918,N_13435,N_12067);
nor U13919 (N_13919,N_12094,N_13321);
and U13920 (N_13920,N_13009,N_12013);
nor U13921 (N_13921,N_12491,N_12197);
nor U13922 (N_13922,N_12445,N_12236);
and U13923 (N_13923,N_12172,N_13338);
nor U13924 (N_13924,N_12481,N_12899);
nor U13925 (N_13925,N_12673,N_13364);
nand U13926 (N_13926,N_12718,N_12221);
nor U13927 (N_13927,N_12068,N_12708);
nand U13928 (N_13928,N_13240,N_12789);
or U13929 (N_13929,N_12113,N_12482);
or U13930 (N_13930,N_12423,N_13122);
nand U13931 (N_13931,N_12886,N_12624);
nor U13932 (N_13932,N_12117,N_12102);
nor U13933 (N_13933,N_13284,N_13142);
or U13934 (N_13934,N_12399,N_12908);
and U13935 (N_13935,N_12661,N_13412);
nor U13936 (N_13936,N_12457,N_12768);
nand U13937 (N_13937,N_12122,N_12077);
nor U13938 (N_13938,N_12165,N_13088);
and U13939 (N_13939,N_12819,N_13208);
nand U13940 (N_13940,N_12652,N_13335);
nor U13941 (N_13941,N_12114,N_12685);
nor U13942 (N_13942,N_12115,N_12380);
nor U13943 (N_13943,N_13362,N_12426);
or U13944 (N_13944,N_12142,N_13167);
nand U13945 (N_13945,N_13133,N_12384);
nand U13946 (N_13946,N_12655,N_12349);
or U13947 (N_13947,N_12952,N_12372);
or U13948 (N_13948,N_12936,N_13406);
nor U13949 (N_13949,N_12112,N_12086);
or U13950 (N_13950,N_13182,N_12164);
nand U13951 (N_13951,N_12573,N_13413);
nand U13952 (N_13952,N_13097,N_13331);
or U13953 (N_13953,N_12406,N_13075);
or U13954 (N_13954,N_12576,N_13151);
nor U13955 (N_13955,N_12494,N_12765);
or U13956 (N_13956,N_12668,N_12550);
nand U13957 (N_13957,N_13350,N_12468);
nand U13958 (N_13958,N_13011,N_13147);
nor U13959 (N_13959,N_12277,N_12264);
and U13960 (N_13960,N_12760,N_12857);
or U13961 (N_13961,N_13400,N_12239);
nand U13962 (N_13962,N_13032,N_13036);
and U13963 (N_13963,N_13101,N_13351);
xnor U13964 (N_13964,N_12017,N_12681);
or U13965 (N_13965,N_12407,N_12078);
or U13966 (N_13966,N_13360,N_12747);
nand U13967 (N_13967,N_12859,N_13277);
nand U13968 (N_13968,N_12055,N_12570);
or U13969 (N_13969,N_12698,N_13016);
or U13970 (N_13970,N_12505,N_13234);
nand U13971 (N_13971,N_12519,N_12725);
nand U13972 (N_13972,N_12178,N_13450);
and U13973 (N_13973,N_12774,N_13107);
nor U13974 (N_13974,N_13150,N_12051);
nor U13975 (N_13975,N_12646,N_12402);
or U13976 (N_13976,N_13049,N_13407);
and U13977 (N_13977,N_12381,N_12997);
or U13978 (N_13978,N_12783,N_13474);
nor U13979 (N_13979,N_13186,N_13038);
or U13980 (N_13980,N_12271,N_13181);
and U13981 (N_13981,N_13033,N_13010);
nand U13982 (N_13982,N_13175,N_12798);
nor U13983 (N_13983,N_12441,N_12393);
nor U13984 (N_13984,N_13017,N_12609);
or U13985 (N_13985,N_12757,N_12304);
nor U13986 (N_13986,N_13149,N_13374);
nor U13987 (N_13987,N_12840,N_13052);
and U13988 (N_13988,N_13174,N_12351);
or U13989 (N_13989,N_13363,N_13021);
and U13990 (N_13990,N_13424,N_12010);
nand U13991 (N_13991,N_12703,N_12395);
nand U13992 (N_13992,N_12863,N_13342);
or U13993 (N_13993,N_13337,N_13433);
nand U13994 (N_13994,N_12918,N_12306);
or U13995 (N_13995,N_12542,N_12037);
or U13996 (N_13996,N_12553,N_12413);
and U13997 (N_13997,N_12601,N_12547);
and U13998 (N_13998,N_12818,N_12854);
nor U13999 (N_13999,N_13361,N_12470);
or U14000 (N_14000,N_12288,N_13129);
or U14001 (N_14001,N_13077,N_12224);
nor U14002 (N_14002,N_12007,N_12732);
nor U14003 (N_14003,N_12348,N_13376);
and U14004 (N_14004,N_13198,N_12653);
nor U14005 (N_14005,N_12543,N_12921);
nand U14006 (N_14006,N_13290,N_13180);
nor U14007 (N_14007,N_12999,N_12483);
nand U14008 (N_14008,N_13266,N_12179);
or U14009 (N_14009,N_13434,N_12539);
or U14010 (N_14010,N_13092,N_12659);
or U14011 (N_14011,N_12318,N_13179);
nand U14012 (N_14012,N_13373,N_12996);
nor U14013 (N_14013,N_13327,N_12617);
and U14014 (N_14014,N_12662,N_13093);
nor U14015 (N_14015,N_12956,N_12502);
and U14016 (N_14016,N_12082,N_12436);
nor U14017 (N_14017,N_12749,N_12282);
and U14018 (N_14018,N_12004,N_12382);
or U14019 (N_14019,N_12544,N_12855);
and U14020 (N_14020,N_12571,N_12188);
nand U14021 (N_14021,N_12705,N_12258);
nand U14022 (N_14022,N_13355,N_13044);
nand U14023 (N_14023,N_12879,N_12439);
and U14024 (N_14024,N_12517,N_13283);
and U14025 (N_14025,N_12549,N_12995);
nand U14026 (N_14026,N_12808,N_13114);
nand U14027 (N_14027,N_12501,N_13003);
or U14028 (N_14028,N_12355,N_12575);
and U14029 (N_14029,N_13064,N_13146);
nand U14030 (N_14030,N_12742,N_13417);
or U14031 (N_14031,N_13476,N_12567);
nand U14032 (N_14032,N_13042,N_12634);
or U14033 (N_14033,N_12717,N_13369);
nand U14034 (N_14034,N_12448,N_12366);
or U14035 (N_14035,N_12509,N_12212);
or U14036 (N_14036,N_12983,N_12709);
nand U14037 (N_14037,N_12041,N_13496);
and U14038 (N_14038,N_13294,N_13491);
nor U14039 (N_14039,N_12726,N_12198);
nor U14040 (N_14040,N_13301,N_13053);
nor U14041 (N_14041,N_13297,N_12302);
or U14042 (N_14042,N_12087,N_13470);
or U14043 (N_14043,N_12901,N_12396);
or U14044 (N_14044,N_12417,N_12155);
and U14045 (N_14045,N_13397,N_12280);
nand U14046 (N_14046,N_13353,N_12027);
or U14047 (N_14047,N_12885,N_13171);
nor U14048 (N_14048,N_12241,N_12181);
nor U14049 (N_14049,N_12435,N_12335);
and U14050 (N_14050,N_12993,N_12682);
or U14051 (N_14051,N_12632,N_13226);
and U14052 (N_14052,N_12261,N_12427);
nand U14053 (N_14053,N_13477,N_12346);
nand U14054 (N_14054,N_12127,N_12613);
nor U14055 (N_14055,N_12533,N_12965);
or U14056 (N_14056,N_12219,N_12336);
nand U14057 (N_14057,N_12752,N_13137);
and U14058 (N_14058,N_12816,N_12974);
or U14059 (N_14059,N_12954,N_12434);
and U14060 (N_14060,N_13344,N_13308);
nand U14061 (N_14061,N_13189,N_13241);
or U14062 (N_14062,N_13243,N_13172);
nor U14063 (N_14063,N_13310,N_12024);
nor U14064 (N_14064,N_13117,N_12897);
or U14065 (N_14065,N_12755,N_13436);
or U14066 (N_14066,N_12126,N_12383);
and U14067 (N_14067,N_13029,N_12773);
nor U14068 (N_14068,N_13452,N_13386);
nor U14069 (N_14069,N_13285,N_13494);
nor U14070 (N_14070,N_13046,N_12377);
and U14071 (N_14071,N_13115,N_12943);
and U14072 (N_14072,N_12305,N_13037);
xnor U14073 (N_14073,N_13218,N_12537);
nor U14074 (N_14074,N_13139,N_12830);
nor U14075 (N_14075,N_12211,N_12209);
nand U14076 (N_14076,N_13130,N_13449);
nand U14077 (N_14077,N_12337,N_13161);
nor U14078 (N_14078,N_12513,N_13201);
nand U14079 (N_14079,N_13034,N_12896);
and U14080 (N_14080,N_12504,N_13451);
or U14081 (N_14081,N_12309,N_13190);
nand U14082 (N_14082,N_12933,N_13249);
nand U14083 (N_14083,N_13103,N_13495);
and U14084 (N_14084,N_12145,N_13455);
nand U14085 (N_14085,N_12391,N_12190);
nor U14086 (N_14086,N_12639,N_12096);
nand U14087 (N_14087,N_12805,N_12986);
and U14088 (N_14088,N_12442,N_12012);
and U14089 (N_14089,N_13488,N_12194);
nand U14090 (N_14090,N_12753,N_13348);
and U14091 (N_14091,N_12325,N_12400);
nor U14092 (N_14092,N_12091,N_12269);
and U14093 (N_14093,N_12488,N_12657);
nand U14094 (N_14094,N_12596,N_13289);
nand U14095 (N_14095,N_13458,N_13490);
or U14096 (N_14096,N_12947,N_12449);
and U14097 (N_14097,N_13058,N_12900);
xnor U14098 (N_14098,N_12289,N_12809);
and U14099 (N_14099,N_12714,N_13083);
and U14100 (N_14100,N_12326,N_13085);
nor U14101 (N_14101,N_12826,N_12577);
nand U14102 (N_14102,N_12512,N_13326);
nor U14103 (N_14103,N_12420,N_12283);
nand U14104 (N_14104,N_12028,N_12751);
or U14105 (N_14105,N_12833,N_13273);
and U14106 (N_14106,N_12846,N_12815);
nor U14107 (N_14107,N_13287,N_12213);
nand U14108 (N_14108,N_13390,N_13113);
or U14109 (N_14109,N_12103,N_12237);
nand U14110 (N_14110,N_12919,N_12370);
and U14111 (N_14111,N_12425,N_12810);
or U14112 (N_14112,N_12844,N_12440);
and U14113 (N_14113,N_13148,N_12016);
nor U14114 (N_14114,N_13307,N_12101);
nand U14115 (N_14115,N_12347,N_12152);
nand U14116 (N_14116,N_13484,N_12120);
xnor U14117 (N_14117,N_13279,N_12710);
nor U14118 (N_14118,N_12167,N_12233);
and U14119 (N_14119,N_13219,N_12834);
or U14120 (N_14120,N_13070,N_13069);
or U14121 (N_14121,N_12430,N_12545);
or U14122 (N_14122,N_12561,N_12014);
or U14123 (N_14123,N_12562,N_12379);
and U14124 (N_14124,N_13073,N_13282);
and U14125 (N_14125,N_12782,N_12131);
nor U14126 (N_14126,N_13123,N_13420);
nand U14127 (N_14127,N_12121,N_12341);
nand U14128 (N_14128,N_12265,N_12599);
and U14129 (N_14129,N_12583,N_13091);
and U14130 (N_14130,N_12775,N_12724);
nor U14131 (N_14131,N_13270,N_13024);
and U14132 (N_14132,N_12556,N_12671);
nand U14133 (N_14133,N_12794,N_13157);
nor U14134 (N_14134,N_12195,N_12604);
nand U14135 (N_14135,N_12895,N_12638);
nor U14136 (N_14136,N_12902,N_13220);
nor U14137 (N_14137,N_13463,N_13483);
and U14138 (N_14138,N_12558,N_12293);
or U14139 (N_14139,N_12554,N_12795);
nor U14140 (N_14140,N_12323,N_12108);
and U14141 (N_14141,N_12911,N_12748);
or U14142 (N_14142,N_12081,N_12169);
nand U14143 (N_14143,N_12408,N_12807);
or U14144 (N_14144,N_12872,N_12252);
nor U14145 (N_14145,N_12715,N_13489);
nor U14146 (N_14146,N_12802,N_12507);
nor U14147 (N_14147,N_13395,N_12286);
xor U14148 (N_14148,N_12255,N_12882);
nand U14149 (N_14149,N_12187,N_12667);
nand U14150 (N_14150,N_13346,N_12141);
or U14151 (N_14151,N_12365,N_12203);
nor U14152 (N_14152,N_12820,N_12612);
or U14153 (N_14153,N_12207,N_12669);
and U14154 (N_14154,N_13399,N_12046);
and U14155 (N_14155,N_13062,N_12867);
or U14156 (N_14156,N_12586,N_12912);
and U14157 (N_14157,N_13368,N_13419);
and U14158 (N_14158,N_12672,N_12125);
and U14159 (N_14159,N_12777,N_12937);
nor U14160 (N_14160,N_13442,N_12960);
or U14161 (N_14161,N_12296,N_12591);
nand U14162 (N_14162,N_12676,N_12564);
or U14163 (N_14163,N_12151,N_12981);
nand U14164 (N_14164,N_13324,N_12052);
nand U14165 (N_14165,N_13328,N_12870);
and U14166 (N_14166,N_13056,N_13230);
or U14167 (N_14167,N_12321,N_12878);
and U14168 (N_14168,N_13063,N_12008);
or U14169 (N_14169,N_12185,N_12022);
nand U14170 (N_14170,N_13261,N_12949);
and U14171 (N_14171,N_12728,N_13408);
or U14172 (N_14172,N_12548,N_12469);
nor U14173 (N_14173,N_12175,N_13177);
nor U14174 (N_14174,N_12791,N_13225);
or U14175 (N_14175,N_12837,N_12438);
nor U14176 (N_14176,N_12080,N_13414);
nor U14177 (N_14177,N_12225,N_12546);
and U14178 (N_14178,N_13319,N_12163);
and U14179 (N_14179,N_12888,N_12330);
or U14180 (N_14180,N_13262,N_12869);
and U14181 (N_14181,N_12026,N_12000);
and U14182 (N_14182,N_12019,N_12358);
or U14183 (N_14183,N_12515,N_13475);
and U14184 (N_14184,N_12664,N_12454);
nand U14185 (N_14185,N_12759,N_12015);
nand U14186 (N_14186,N_12551,N_12660);
nor U14187 (N_14187,N_12176,N_13089);
nor U14188 (N_14188,N_12298,N_13031);
and U14189 (N_14189,N_13453,N_12521);
and U14190 (N_14190,N_12796,N_12932);
or U14191 (N_14191,N_12508,N_13232);
nor U14192 (N_14192,N_12180,N_13209);
and U14193 (N_14193,N_13131,N_12893);
xor U14194 (N_14194,N_12210,N_12514);
and U14195 (N_14195,N_12076,N_13426);
nor U14196 (N_14196,N_12829,N_13347);
and U14197 (N_14197,N_13041,N_12581);
nand U14198 (N_14198,N_12267,N_12970);
nor U14199 (N_14199,N_12216,N_12444);
nor U14200 (N_14200,N_12858,N_13422);
or U14201 (N_14201,N_12364,N_12938);
or U14202 (N_14202,N_12263,N_12232);
and U14203 (N_14203,N_13200,N_12410);
or U14204 (N_14204,N_12874,N_12274);
and U14205 (N_14205,N_13404,N_12894);
or U14206 (N_14206,N_13311,N_12666);
or U14207 (N_14207,N_12058,N_12784);
or U14208 (N_14208,N_12272,N_12247);
and U14209 (N_14209,N_13247,N_12684);
nand U14210 (N_14210,N_12825,N_12744);
and U14211 (N_14211,N_12868,N_13304);
or U14212 (N_14212,N_12312,N_12071);
and U14213 (N_14213,N_13481,N_12031);
nor U14214 (N_14214,N_13479,N_13329);
nand U14215 (N_14215,N_12428,N_13295);
nand U14216 (N_14216,N_12353,N_12677);
or U14217 (N_14217,N_12070,N_12200);
and U14218 (N_14218,N_13486,N_12342);
and U14219 (N_14219,N_12953,N_13299);
or U14220 (N_14220,N_12898,N_12463);
and U14221 (N_14221,N_12204,N_12106);
nand U14222 (N_14222,N_13163,N_13086);
xnor U14223 (N_14223,N_12614,N_12674);
and U14224 (N_14224,N_12294,N_12416);
or U14225 (N_14225,N_12928,N_13431);
and U14226 (N_14226,N_12110,N_12792);
nand U14227 (N_14227,N_12414,N_13134);
and U14228 (N_14228,N_13236,N_13135);
nand U14229 (N_14229,N_12299,N_12980);
or U14230 (N_14230,N_13454,N_12958);
nand U14231 (N_14231,N_12801,N_13471);
xor U14232 (N_14232,N_12418,N_13099);
nand U14233 (N_14233,N_12253,N_12144);
nand U14234 (N_14234,N_12230,N_13066);
or U14235 (N_14235,N_13237,N_12623);
and U14236 (N_14236,N_12762,N_12675);
nand U14237 (N_14237,N_12984,N_12446);
and U14238 (N_14238,N_13222,N_12005);
or U14239 (N_14239,N_13006,N_12487);
or U14240 (N_14240,N_13211,N_12738);
nor U14241 (N_14241,N_13334,N_12887);
nor U14242 (N_14242,N_12707,N_12821);
or U14243 (N_14243,N_12906,N_13392);
nor U14244 (N_14244,N_13223,N_12039);
nor U14245 (N_14245,N_12447,N_12075);
nand U14246 (N_14246,N_12721,N_13224);
or U14247 (N_14247,N_12214,N_12150);
or U14248 (N_14248,N_13379,N_12865);
and U14249 (N_14249,N_12461,N_12320);
nand U14250 (N_14250,N_12031,N_12556);
nand U14251 (N_14251,N_13088,N_13107);
or U14252 (N_14252,N_13344,N_12242);
or U14253 (N_14253,N_12212,N_13389);
or U14254 (N_14254,N_12216,N_12162);
or U14255 (N_14255,N_13451,N_13489);
nor U14256 (N_14256,N_12668,N_12103);
and U14257 (N_14257,N_12725,N_12445);
nand U14258 (N_14258,N_12435,N_12935);
and U14259 (N_14259,N_13064,N_12641);
and U14260 (N_14260,N_12041,N_12436);
or U14261 (N_14261,N_12432,N_13314);
nor U14262 (N_14262,N_12513,N_12096);
nor U14263 (N_14263,N_12370,N_13267);
nor U14264 (N_14264,N_12495,N_13449);
or U14265 (N_14265,N_12860,N_13333);
or U14266 (N_14266,N_12447,N_12688);
and U14267 (N_14267,N_12654,N_12882);
nor U14268 (N_14268,N_12535,N_12589);
nor U14269 (N_14269,N_13306,N_12786);
nand U14270 (N_14270,N_12128,N_12492);
and U14271 (N_14271,N_12836,N_12699);
nor U14272 (N_14272,N_12712,N_12105);
nor U14273 (N_14273,N_13020,N_12592);
and U14274 (N_14274,N_13022,N_13329);
and U14275 (N_14275,N_12772,N_13258);
nor U14276 (N_14276,N_13102,N_12130);
or U14277 (N_14277,N_12830,N_12268);
or U14278 (N_14278,N_13311,N_12906);
nand U14279 (N_14279,N_13314,N_12016);
nor U14280 (N_14280,N_13327,N_12896);
nor U14281 (N_14281,N_12927,N_12826);
nor U14282 (N_14282,N_12310,N_12147);
or U14283 (N_14283,N_12347,N_13056);
xnor U14284 (N_14284,N_12363,N_13453);
and U14285 (N_14285,N_12478,N_12985);
or U14286 (N_14286,N_12917,N_12363);
nand U14287 (N_14287,N_12990,N_12624);
or U14288 (N_14288,N_13298,N_12168);
and U14289 (N_14289,N_13443,N_13321);
and U14290 (N_14290,N_12816,N_12751);
and U14291 (N_14291,N_12785,N_13443);
or U14292 (N_14292,N_12800,N_12192);
and U14293 (N_14293,N_13409,N_12362);
or U14294 (N_14294,N_13156,N_12571);
and U14295 (N_14295,N_12852,N_12010);
or U14296 (N_14296,N_13091,N_13458);
and U14297 (N_14297,N_13276,N_12687);
and U14298 (N_14298,N_13411,N_12783);
nor U14299 (N_14299,N_12725,N_12110);
or U14300 (N_14300,N_13280,N_12919);
nand U14301 (N_14301,N_13127,N_13467);
and U14302 (N_14302,N_13266,N_12446);
or U14303 (N_14303,N_13040,N_12940);
and U14304 (N_14304,N_12542,N_12927);
nand U14305 (N_14305,N_12767,N_12744);
and U14306 (N_14306,N_12842,N_13250);
and U14307 (N_14307,N_12024,N_12177);
or U14308 (N_14308,N_12954,N_13158);
and U14309 (N_14309,N_13251,N_12236);
nor U14310 (N_14310,N_13402,N_12959);
nor U14311 (N_14311,N_13296,N_13270);
nor U14312 (N_14312,N_13078,N_13138);
or U14313 (N_14313,N_12277,N_12275);
and U14314 (N_14314,N_13279,N_12916);
nor U14315 (N_14315,N_12148,N_13315);
and U14316 (N_14316,N_13498,N_12130);
nand U14317 (N_14317,N_12189,N_13271);
nor U14318 (N_14318,N_12945,N_13469);
and U14319 (N_14319,N_12570,N_12691);
nand U14320 (N_14320,N_12790,N_12692);
nor U14321 (N_14321,N_13310,N_13159);
nand U14322 (N_14322,N_13493,N_12330);
nor U14323 (N_14323,N_13168,N_13050);
or U14324 (N_14324,N_12434,N_13108);
and U14325 (N_14325,N_13037,N_12600);
nor U14326 (N_14326,N_12769,N_12105);
xnor U14327 (N_14327,N_12701,N_13064);
nor U14328 (N_14328,N_13118,N_12744);
nor U14329 (N_14329,N_12814,N_12064);
nor U14330 (N_14330,N_13091,N_12949);
and U14331 (N_14331,N_13382,N_13127);
and U14332 (N_14332,N_13358,N_12855);
or U14333 (N_14333,N_12996,N_13021);
and U14334 (N_14334,N_12693,N_12837);
nor U14335 (N_14335,N_12229,N_13030);
nand U14336 (N_14336,N_12276,N_12971);
xnor U14337 (N_14337,N_13091,N_13169);
nand U14338 (N_14338,N_13410,N_13367);
nor U14339 (N_14339,N_13227,N_13372);
nor U14340 (N_14340,N_12114,N_13300);
and U14341 (N_14341,N_12043,N_12335);
or U14342 (N_14342,N_12603,N_12133);
nand U14343 (N_14343,N_12641,N_12857);
and U14344 (N_14344,N_12130,N_12787);
and U14345 (N_14345,N_13122,N_12726);
nor U14346 (N_14346,N_12308,N_13121);
nand U14347 (N_14347,N_12619,N_12912);
nand U14348 (N_14348,N_13075,N_12186);
or U14349 (N_14349,N_12008,N_12553);
or U14350 (N_14350,N_12380,N_12313);
nand U14351 (N_14351,N_12541,N_13088);
nand U14352 (N_14352,N_12064,N_12904);
nand U14353 (N_14353,N_12524,N_12243);
nand U14354 (N_14354,N_12323,N_13454);
nand U14355 (N_14355,N_12656,N_12699);
nor U14356 (N_14356,N_13248,N_12115);
nor U14357 (N_14357,N_13408,N_12396);
or U14358 (N_14358,N_12134,N_12642);
nand U14359 (N_14359,N_12559,N_12980);
and U14360 (N_14360,N_12606,N_12663);
nor U14361 (N_14361,N_12571,N_12947);
or U14362 (N_14362,N_13147,N_13488);
and U14363 (N_14363,N_13298,N_13314);
or U14364 (N_14364,N_12972,N_12901);
or U14365 (N_14365,N_12761,N_12396);
or U14366 (N_14366,N_13286,N_12920);
and U14367 (N_14367,N_12447,N_12295);
xor U14368 (N_14368,N_12455,N_13492);
and U14369 (N_14369,N_12469,N_12881);
or U14370 (N_14370,N_12006,N_12928);
or U14371 (N_14371,N_12375,N_13423);
nand U14372 (N_14372,N_12840,N_12713);
nand U14373 (N_14373,N_12810,N_13288);
nor U14374 (N_14374,N_12451,N_12604);
and U14375 (N_14375,N_12388,N_12948);
and U14376 (N_14376,N_12454,N_13100);
nor U14377 (N_14377,N_12392,N_12882);
nor U14378 (N_14378,N_12453,N_12103);
nor U14379 (N_14379,N_12179,N_12779);
nand U14380 (N_14380,N_12320,N_12403);
nor U14381 (N_14381,N_12578,N_13355);
or U14382 (N_14382,N_12962,N_12902);
and U14383 (N_14383,N_12543,N_12028);
and U14384 (N_14384,N_13349,N_13246);
nand U14385 (N_14385,N_12738,N_13490);
nand U14386 (N_14386,N_12372,N_12660);
nand U14387 (N_14387,N_12229,N_13346);
and U14388 (N_14388,N_12233,N_12929);
and U14389 (N_14389,N_13475,N_12458);
or U14390 (N_14390,N_12099,N_13198);
nor U14391 (N_14391,N_13345,N_13342);
xnor U14392 (N_14392,N_12879,N_13493);
nand U14393 (N_14393,N_13459,N_13135);
xor U14394 (N_14394,N_12185,N_12743);
or U14395 (N_14395,N_13005,N_13485);
and U14396 (N_14396,N_12503,N_13041);
nor U14397 (N_14397,N_12585,N_12713);
and U14398 (N_14398,N_12223,N_12293);
nand U14399 (N_14399,N_12551,N_12640);
or U14400 (N_14400,N_12460,N_12816);
xor U14401 (N_14401,N_12654,N_12279);
nor U14402 (N_14402,N_13412,N_12766);
and U14403 (N_14403,N_12490,N_12454);
or U14404 (N_14404,N_13092,N_12668);
and U14405 (N_14405,N_12470,N_13189);
nor U14406 (N_14406,N_13202,N_13010);
or U14407 (N_14407,N_12436,N_12348);
and U14408 (N_14408,N_13412,N_13187);
and U14409 (N_14409,N_12633,N_12504);
nor U14410 (N_14410,N_12533,N_12191);
or U14411 (N_14411,N_12852,N_12974);
and U14412 (N_14412,N_12588,N_12509);
nand U14413 (N_14413,N_13279,N_12782);
or U14414 (N_14414,N_13497,N_12120);
nor U14415 (N_14415,N_13061,N_13134);
nor U14416 (N_14416,N_12963,N_12235);
and U14417 (N_14417,N_12786,N_12942);
or U14418 (N_14418,N_13078,N_12440);
and U14419 (N_14419,N_13443,N_12458);
nand U14420 (N_14420,N_12578,N_12556);
and U14421 (N_14421,N_12869,N_13195);
nor U14422 (N_14422,N_13415,N_12421);
nand U14423 (N_14423,N_13390,N_13470);
nor U14424 (N_14424,N_12436,N_13453);
and U14425 (N_14425,N_12778,N_12497);
nand U14426 (N_14426,N_12250,N_13315);
and U14427 (N_14427,N_12982,N_12258);
and U14428 (N_14428,N_12607,N_13448);
or U14429 (N_14429,N_12083,N_13495);
nand U14430 (N_14430,N_12254,N_12819);
nor U14431 (N_14431,N_12773,N_12310);
or U14432 (N_14432,N_13442,N_12874);
and U14433 (N_14433,N_13196,N_12576);
or U14434 (N_14434,N_12031,N_12345);
nand U14435 (N_14435,N_12055,N_13490);
nand U14436 (N_14436,N_12357,N_12119);
nand U14437 (N_14437,N_12059,N_13107);
and U14438 (N_14438,N_13097,N_12125);
or U14439 (N_14439,N_13123,N_12141);
and U14440 (N_14440,N_13464,N_12776);
nand U14441 (N_14441,N_12526,N_12238);
or U14442 (N_14442,N_13264,N_12488);
and U14443 (N_14443,N_12353,N_12523);
nand U14444 (N_14444,N_12606,N_12241);
nor U14445 (N_14445,N_13031,N_12823);
or U14446 (N_14446,N_12616,N_12346);
nand U14447 (N_14447,N_13282,N_13155);
or U14448 (N_14448,N_12589,N_13036);
and U14449 (N_14449,N_12312,N_12027);
nand U14450 (N_14450,N_12811,N_12949);
nand U14451 (N_14451,N_13248,N_13471);
nand U14452 (N_14452,N_13090,N_12178);
nor U14453 (N_14453,N_12987,N_12696);
nor U14454 (N_14454,N_12685,N_12057);
nand U14455 (N_14455,N_12600,N_12854);
or U14456 (N_14456,N_13338,N_12711);
and U14457 (N_14457,N_12288,N_12228);
nand U14458 (N_14458,N_13081,N_13114);
or U14459 (N_14459,N_12588,N_12691);
nor U14460 (N_14460,N_13489,N_12209);
nor U14461 (N_14461,N_12579,N_12140);
nor U14462 (N_14462,N_12981,N_12759);
nor U14463 (N_14463,N_12166,N_12709);
or U14464 (N_14464,N_12537,N_13302);
or U14465 (N_14465,N_12585,N_12115);
and U14466 (N_14466,N_12065,N_12167);
nor U14467 (N_14467,N_12406,N_13093);
or U14468 (N_14468,N_12240,N_13265);
and U14469 (N_14469,N_12289,N_13076);
or U14470 (N_14470,N_13157,N_13454);
or U14471 (N_14471,N_12024,N_13332);
and U14472 (N_14472,N_12125,N_12230);
and U14473 (N_14473,N_12758,N_12113);
and U14474 (N_14474,N_12834,N_12609);
nand U14475 (N_14475,N_12044,N_12355);
nand U14476 (N_14476,N_12883,N_12438);
nor U14477 (N_14477,N_12569,N_12824);
nand U14478 (N_14478,N_13294,N_13474);
or U14479 (N_14479,N_12236,N_12347);
nand U14480 (N_14480,N_12805,N_12958);
or U14481 (N_14481,N_13394,N_13163);
or U14482 (N_14482,N_13025,N_12089);
xnor U14483 (N_14483,N_12000,N_12187);
nand U14484 (N_14484,N_13321,N_12017);
or U14485 (N_14485,N_12719,N_12955);
nor U14486 (N_14486,N_13260,N_12584);
or U14487 (N_14487,N_13493,N_13159);
or U14488 (N_14488,N_12990,N_12307);
and U14489 (N_14489,N_12620,N_12836);
and U14490 (N_14490,N_12317,N_12277);
or U14491 (N_14491,N_12423,N_13006);
and U14492 (N_14492,N_12707,N_13348);
nand U14493 (N_14493,N_12915,N_13374);
and U14494 (N_14494,N_12996,N_12511);
nand U14495 (N_14495,N_13267,N_12337);
or U14496 (N_14496,N_13346,N_12129);
nand U14497 (N_14497,N_13355,N_13396);
and U14498 (N_14498,N_12998,N_12781);
nor U14499 (N_14499,N_12727,N_13332);
nor U14500 (N_14500,N_13449,N_12878);
nor U14501 (N_14501,N_12387,N_13355);
nor U14502 (N_14502,N_12707,N_12803);
nand U14503 (N_14503,N_12561,N_12007);
and U14504 (N_14504,N_13319,N_13335);
and U14505 (N_14505,N_13272,N_13298);
or U14506 (N_14506,N_12462,N_12743);
and U14507 (N_14507,N_13103,N_13354);
nor U14508 (N_14508,N_12654,N_12641);
nand U14509 (N_14509,N_12487,N_12389);
nor U14510 (N_14510,N_13186,N_12086);
nand U14511 (N_14511,N_13142,N_12013);
or U14512 (N_14512,N_12045,N_13197);
or U14513 (N_14513,N_13201,N_12025);
nand U14514 (N_14514,N_12385,N_13374);
or U14515 (N_14515,N_12396,N_12943);
and U14516 (N_14516,N_12210,N_13153);
and U14517 (N_14517,N_12955,N_13420);
and U14518 (N_14518,N_13195,N_13496);
nand U14519 (N_14519,N_13075,N_12911);
nand U14520 (N_14520,N_13359,N_12070);
or U14521 (N_14521,N_12081,N_12899);
nor U14522 (N_14522,N_12747,N_12783);
and U14523 (N_14523,N_13015,N_12795);
nor U14524 (N_14524,N_12211,N_13488);
and U14525 (N_14525,N_12864,N_12181);
and U14526 (N_14526,N_12885,N_12886);
nor U14527 (N_14527,N_12127,N_12679);
nand U14528 (N_14528,N_12878,N_13418);
and U14529 (N_14529,N_13107,N_12303);
and U14530 (N_14530,N_12330,N_12045);
or U14531 (N_14531,N_12935,N_13198);
or U14532 (N_14532,N_13071,N_12555);
and U14533 (N_14533,N_13269,N_13497);
or U14534 (N_14534,N_13120,N_12223);
and U14535 (N_14535,N_13074,N_12917);
nor U14536 (N_14536,N_13032,N_12443);
nand U14537 (N_14537,N_12404,N_12426);
or U14538 (N_14538,N_13328,N_12084);
nor U14539 (N_14539,N_13093,N_12270);
or U14540 (N_14540,N_13253,N_12548);
nand U14541 (N_14541,N_12733,N_12875);
and U14542 (N_14542,N_12209,N_13243);
or U14543 (N_14543,N_12786,N_12249);
nor U14544 (N_14544,N_12510,N_13487);
nand U14545 (N_14545,N_13165,N_13185);
or U14546 (N_14546,N_12973,N_12182);
nand U14547 (N_14547,N_12362,N_12925);
nand U14548 (N_14548,N_12281,N_13422);
nand U14549 (N_14549,N_12228,N_13070);
nand U14550 (N_14550,N_12886,N_12857);
nor U14551 (N_14551,N_12652,N_12144);
nor U14552 (N_14552,N_13403,N_13368);
nand U14553 (N_14553,N_12366,N_12605);
or U14554 (N_14554,N_12161,N_13061);
nor U14555 (N_14555,N_12724,N_13306);
nor U14556 (N_14556,N_12204,N_13477);
nand U14557 (N_14557,N_12066,N_13470);
nand U14558 (N_14558,N_12856,N_12369);
or U14559 (N_14559,N_12142,N_12122);
nor U14560 (N_14560,N_12343,N_12808);
and U14561 (N_14561,N_13160,N_12303);
nor U14562 (N_14562,N_13371,N_12414);
nand U14563 (N_14563,N_12071,N_12852);
nor U14564 (N_14564,N_12180,N_12857);
nand U14565 (N_14565,N_12356,N_13003);
nor U14566 (N_14566,N_13451,N_13386);
or U14567 (N_14567,N_12723,N_13383);
nand U14568 (N_14568,N_12429,N_12331);
and U14569 (N_14569,N_12821,N_12001);
nor U14570 (N_14570,N_12822,N_13143);
and U14571 (N_14571,N_12080,N_12150);
nor U14572 (N_14572,N_12640,N_12801);
nand U14573 (N_14573,N_12583,N_12845);
and U14574 (N_14574,N_12136,N_12368);
and U14575 (N_14575,N_12966,N_13148);
or U14576 (N_14576,N_12934,N_12093);
nand U14577 (N_14577,N_12885,N_12929);
nand U14578 (N_14578,N_13305,N_13015);
and U14579 (N_14579,N_13436,N_12864);
and U14580 (N_14580,N_13159,N_12626);
xor U14581 (N_14581,N_13053,N_12532);
or U14582 (N_14582,N_12860,N_12490);
or U14583 (N_14583,N_12612,N_13026);
and U14584 (N_14584,N_12691,N_12354);
and U14585 (N_14585,N_12088,N_12108);
and U14586 (N_14586,N_12129,N_12171);
or U14587 (N_14587,N_12400,N_12602);
nand U14588 (N_14588,N_12268,N_13424);
and U14589 (N_14589,N_12176,N_12046);
or U14590 (N_14590,N_12995,N_12567);
and U14591 (N_14591,N_12977,N_12066);
nand U14592 (N_14592,N_12814,N_12860);
or U14593 (N_14593,N_12746,N_12661);
or U14594 (N_14594,N_12324,N_12168);
or U14595 (N_14595,N_12331,N_12785);
and U14596 (N_14596,N_12979,N_12403);
and U14597 (N_14597,N_12213,N_13314);
or U14598 (N_14598,N_12321,N_12405);
and U14599 (N_14599,N_13167,N_13260);
or U14600 (N_14600,N_12363,N_12743);
nor U14601 (N_14601,N_12217,N_12037);
and U14602 (N_14602,N_12170,N_12466);
nand U14603 (N_14603,N_12265,N_13020);
nand U14604 (N_14604,N_12684,N_13051);
and U14605 (N_14605,N_13337,N_12398);
nand U14606 (N_14606,N_12351,N_12147);
nand U14607 (N_14607,N_12642,N_12704);
nor U14608 (N_14608,N_13063,N_12642);
nand U14609 (N_14609,N_12194,N_12432);
nand U14610 (N_14610,N_12694,N_12321);
or U14611 (N_14611,N_13463,N_12584);
nand U14612 (N_14612,N_13205,N_13207);
xor U14613 (N_14613,N_13280,N_12908);
or U14614 (N_14614,N_12304,N_12959);
and U14615 (N_14615,N_12019,N_13465);
and U14616 (N_14616,N_12224,N_12757);
and U14617 (N_14617,N_12802,N_13369);
nand U14618 (N_14618,N_13457,N_12261);
and U14619 (N_14619,N_12258,N_12666);
nor U14620 (N_14620,N_12256,N_12156);
and U14621 (N_14621,N_12068,N_12649);
nand U14622 (N_14622,N_12543,N_12173);
nand U14623 (N_14623,N_12041,N_12035);
nand U14624 (N_14624,N_12502,N_13079);
nor U14625 (N_14625,N_12537,N_13135);
or U14626 (N_14626,N_12064,N_12416);
nor U14627 (N_14627,N_12401,N_12038);
or U14628 (N_14628,N_13480,N_12913);
nor U14629 (N_14629,N_13252,N_12105);
and U14630 (N_14630,N_12623,N_12161);
and U14631 (N_14631,N_12697,N_13298);
and U14632 (N_14632,N_13458,N_13497);
nor U14633 (N_14633,N_13259,N_13471);
and U14634 (N_14634,N_12008,N_13398);
and U14635 (N_14635,N_13400,N_13280);
or U14636 (N_14636,N_12289,N_12803);
or U14637 (N_14637,N_12798,N_12593);
or U14638 (N_14638,N_12403,N_12748);
and U14639 (N_14639,N_13131,N_12822);
nor U14640 (N_14640,N_12313,N_12710);
or U14641 (N_14641,N_12418,N_12324);
and U14642 (N_14642,N_12411,N_12603);
and U14643 (N_14643,N_13495,N_12154);
nor U14644 (N_14644,N_12947,N_13421);
nand U14645 (N_14645,N_13415,N_12536);
or U14646 (N_14646,N_12092,N_12324);
and U14647 (N_14647,N_12107,N_12361);
nand U14648 (N_14648,N_12960,N_13228);
nor U14649 (N_14649,N_12165,N_12135);
and U14650 (N_14650,N_12267,N_12898);
nand U14651 (N_14651,N_12202,N_13020);
nand U14652 (N_14652,N_12098,N_13377);
nor U14653 (N_14653,N_12750,N_12618);
or U14654 (N_14654,N_12080,N_12325);
nand U14655 (N_14655,N_12523,N_12358);
nor U14656 (N_14656,N_12792,N_13471);
or U14657 (N_14657,N_13138,N_13334);
and U14658 (N_14658,N_12958,N_12322);
nor U14659 (N_14659,N_13394,N_12215);
and U14660 (N_14660,N_12923,N_12521);
or U14661 (N_14661,N_12515,N_13059);
nand U14662 (N_14662,N_13103,N_12672);
and U14663 (N_14663,N_12931,N_13491);
nor U14664 (N_14664,N_13424,N_12331);
or U14665 (N_14665,N_13284,N_12038);
nand U14666 (N_14666,N_12016,N_12962);
nand U14667 (N_14667,N_13033,N_12416);
nor U14668 (N_14668,N_12156,N_12000);
or U14669 (N_14669,N_12099,N_13129);
or U14670 (N_14670,N_13024,N_13042);
nor U14671 (N_14671,N_12223,N_12089);
or U14672 (N_14672,N_12916,N_12786);
or U14673 (N_14673,N_12608,N_12212);
nand U14674 (N_14674,N_13271,N_12260);
or U14675 (N_14675,N_12021,N_12058);
nor U14676 (N_14676,N_12847,N_12184);
and U14677 (N_14677,N_12197,N_13134);
nor U14678 (N_14678,N_12911,N_12478);
or U14679 (N_14679,N_12115,N_12467);
and U14680 (N_14680,N_13411,N_13126);
or U14681 (N_14681,N_13336,N_13174);
nand U14682 (N_14682,N_12375,N_13357);
nor U14683 (N_14683,N_12544,N_12634);
nor U14684 (N_14684,N_13280,N_12577);
xnor U14685 (N_14685,N_13314,N_12450);
nor U14686 (N_14686,N_12888,N_12638);
nand U14687 (N_14687,N_13323,N_12469);
nor U14688 (N_14688,N_12313,N_12376);
or U14689 (N_14689,N_13073,N_12572);
nand U14690 (N_14690,N_12264,N_12897);
nand U14691 (N_14691,N_12710,N_12650);
or U14692 (N_14692,N_12152,N_12885);
or U14693 (N_14693,N_13079,N_13035);
or U14694 (N_14694,N_12362,N_12461);
and U14695 (N_14695,N_13075,N_12463);
nor U14696 (N_14696,N_12987,N_12649);
nor U14697 (N_14697,N_12685,N_13256);
nor U14698 (N_14698,N_13303,N_12386);
and U14699 (N_14699,N_12091,N_12641);
or U14700 (N_14700,N_12727,N_12283);
or U14701 (N_14701,N_12183,N_12919);
nand U14702 (N_14702,N_12986,N_12860);
or U14703 (N_14703,N_13144,N_13457);
nand U14704 (N_14704,N_12125,N_13306);
and U14705 (N_14705,N_12668,N_12950);
nand U14706 (N_14706,N_12315,N_12463);
nor U14707 (N_14707,N_13313,N_12970);
and U14708 (N_14708,N_12861,N_12379);
and U14709 (N_14709,N_13391,N_13254);
and U14710 (N_14710,N_12927,N_12131);
nand U14711 (N_14711,N_13262,N_12675);
or U14712 (N_14712,N_12527,N_13039);
nand U14713 (N_14713,N_12931,N_12486);
nor U14714 (N_14714,N_12425,N_12907);
or U14715 (N_14715,N_13221,N_12570);
and U14716 (N_14716,N_12225,N_13185);
or U14717 (N_14717,N_13044,N_13009);
and U14718 (N_14718,N_13098,N_12835);
or U14719 (N_14719,N_12984,N_12149);
nand U14720 (N_14720,N_12303,N_13272);
nand U14721 (N_14721,N_12999,N_13372);
nand U14722 (N_14722,N_13140,N_13424);
or U14723 (N_14723,N_12571,N_12522);
nor U14724 (N_14724,N_12497,N_12122);
nor U14725 (N_14725,N_13095,N_13349);
nor U14726 (N_14726,N_13330,N_13210);
nand U14727 (N_14727,N_12484,N_12092);
or U14728 (N_14728,N_13435,N_12357);
nor U14729 (N_14729,N_12659,N_12098);
nor U14730 (N_14730,N_13018,N_12533);
nand U14731 (N_14731,N_12502,N_12175);
and U14732 (N_14732,N_12313,N_12255);
nor U14733 (N_14733,N_13302,N_13432);
nand U14734 (N_14734,N_12259,N_12607);
or U14735 (N_14735,N_13159,N_12251);
and U14736 (N_14736,N_12531,N_12658);
nor U14737 (N_14737,N_12945,N_12663);
nand U14738 (N_14738,N_12062,N_12272);
or U14739 (N_14739,N_12029,N_12486);
nand U14740 (N_14740,N_12265,N_13332);
or U14741 (N_14741,N_12122,N_13271);
and U14742 (N_14742,N_12902,N_13149);
and U14743 (N_14743,N_12498,N_13197);
or U14744 (N_14744,N_13154,N_13112);
nor U14745 (N_14745,N_13070,N_13257);
nand U14746 (N_14746,N_12433,N_12158);
nand U14747 (N_14747,N_12698,N_12365);
or U14748 (N_14748,N_12302,N_13038);
or U14749 (N_14749,N_12191,N_12287);
nor U14750 (N_14750,N_12329,N_12889);
nor U14751 (N_14751,N_13249,N_12105);
nor U14752 (N_14752,N_13327,N_13420);
nand U14753 (N_14753,N_12811,N_12612);
nor U14754 (N_14754,N_12324,N_13497);
nand U14755 (N_14755,N_12525,N_13156);
or U14756 (N_14756,N_12321,N_12729);
xor U14757 (N_14757,N_12439,N_12932);
nand U14758 (N_14758,N_12167,N_13204);
nand U14759 (N_14759,N_13155,N_12093);
or U14760 (N_14760,N_12861,N_12001);
nor U14761 (N_14761,N_13249,N_12095);
or U14762 (N_14762,N_13124,N_13147);
nor U14763 (N_14763,N_12247,N_12273);
and U14764 (N_14764,N_12840,N_13343);
nand U14765 (N_14765,N_13129,N_13418);
nor U14766 (N_14766,N_12725,N_12728);
nand U14767 (N_14767,N_12978,N_13128);
and U14768 (N_14768,N_13086,N_13252);
or U14769 (N_14769,N_12008,N_13378);
nand U14770 (N_14770,N_12835,N_12272);
nand U14771 (N_14771,N_12776,N_12642);
or U14772 (N_14772,N_12067,N_12306);
and U14773 (N_14773,N_12614,N_12434);
and U14774 (N_14774,N_12152,N_13246);
nand U14775 (N_14775,N_12557,N_12563);
or U14776 (N_14776,N_12160,N_13102);
or U14777 (N_14777,N_12795,N_13122);
or U14778 (N_14778,N_13144,N_12110);
and U14779 (N_14779,N_13408,N_12620);
nand U14780 (N_14780,N_12578,N_12276);
and U14781 (N_14781,N_13014,N_13099);
and U14782 (N_14782,N_12954,N_12886);
nand U14783 (N_14783,N_12833,N_13191);
nor U14784 (N_14784,N_13235,N_12019);
or U14785 (N_14785,N_12393,N_12517);
nor U14786 (N_14786,N_12810,N_13029);
xor U14787 (N_14787,N_12775,N_13028);
nor U14788 (N_14788,N_13428,N_12101);
nor U14789 (N_14789,N_12213,N_12378);
or U14790 (N_14790,N_12556,N_12867);
or U14791 (N_14791,N_13210,N_12770);
nand U14792 (N_14792,N_12393,N_13395);
nor U14793 (N_14793,N_12028,N_13293);
nand U14794 (N_14794,N_13025,N_13436);
or U14795 (N_14795,N_12854,N_12306);
or U14796 (N_14796,N_13384,N_12735);
nand U14797 (N_14797,N_12193,N_12955);
and U14798 (N_14798,N_12502,N_12537);
or U14799 (N_14799,N_12871,N_12393);
and U14800 (N_14800,N_12768,N_12903);
or U14801 (N_14801,N_12716,N_12121);
or U14802 (N_14802,N_13248,N_12249);
nand U14803 (N_14803,N_12565,N_12337);
or U14804 (N_14804,N_12246,N_12030);
and U14805 (N_14805,N_12299,N_12891);
or U14806 (N_14806,N_12493,N_13081);
nor U14807 (N_14807,N_13380,N_12437);
xnor U14808 (N_14808,N_12223,N_12657);
nor U14809 (N_14809,N_13431,N_13338);
and U14810 (N_14810,N_12665,N_12127);
or U14811 (N_14811,N_13093,N_12046);
nor U14812 (N_14812,N_13408,N_12928);
or U14813 (N_14813,N_12170,N_13384);
or U14814 (N_14814,N_13082,N_13144);
and U14815 (N_14815,N_12470,N_12320);
nor U14816 (N_14816,N_13458,N_13334);
nor U14817 (N_14817,N_12389,N_13464);
nand U14818 (N_14818,N_12427,N_13237);
nor U14819 (N_14819,N_12565,N_12680);
nand U14820 (N_14820,N_12554,N_12378);
nand U14821 (N_14821,N_13487,N_12668);
nand U14822 (N_14822,N_12366,N_13326);
nor U14823 (N_14823,N_13306,N_13103);
or U14824 (N_14824,N_12702,N_12391);
or U14825 (N_14825,N_12221,N_12700);
and U14826 (N_14826,N_12484,N_12675);
nor U14827 (N_14827,N_12572,N_12852);
and U14828 (N_14828,N_12846,N_12574);
nand U14829 (N_14829,N_13384,N_12556);
nor U14830 (N_14830,N_13478,N_12672);
and U14831 (N_14831,N_12378,N_12529);
nand U14832 (N_14832,N_13231,N_12931);
and U14833 (N_14833,N_12773,N_13191);
and U14834 (N_14834,N_12180,N_13321);
or U14835 (N_14835,N_13112,N_12128);
nand U14836 (N_14836,N_13058,N_12058);
and U14837 (N_14837,N_12414,N_12210);
and U14838 (N_14838,N_13008,N_13230);
and U14839 (N_14839,N_12575,N_12271);
or U14840 (N_14840,N_12527,N_13239);
or U14841 (N_14841,N_12552,N_12363);
nor U14842 (N_14842,N_12659,N_12432);
and U14843 (N_14843,N_12671,N_13136);
and U14844 (N_14844,N_12058,N_12478);
or U14845 (N_14845,N_12126,N_13130);
nand U14846 (N_14846,N_12515,N_12594);
and U14847 (N_14847,N_12661,N_12198);
nand U14848 (N_14848,N_12439,N_13056);
xor U14849 (N_14849,N_12493,N_12282);
and U14850 (N_14850,N_13393,N_12224);
nand U14851 (N_14851,N_12154,N_13039);
or U14852 (N_14852,N_12646,N_12624);
and U14853 (N_14853,N_13059,N_12753);
and U14854 (N_14854,N_13439,N_13011);
and U14855 (N_14855,N_12262,N_13364);
nor U14856 (N_14856,N_13088,N_12852);
or U14857 (N_14857,N_12286,N_12746);
nand U14858 (N_14858,N_13098,N_12582);
xor U14859 (N_14859,N_12908,N_12193);
and U14860 (N_14860,N_13196,N_13018);
nor U14861 (N_14861,N_12397,N_12812);
xor U14862 (N_14862,N_13376,N_12217);
nor U14863 (N_14863,N_12789,N_12425);
nor U14864 (N_14864,N_12421,N_12511);
and U14865 (N_14865,N_12543,N_12958);
nand U14866 (N_14866,N_12461,N_13365);
or U14867 (N_14867,N_12418,N_12261);
and U14868 (N_14868,N_12273,N_12744);
nor U14869 (N_14869,N_13374,N_13010);
nand U14870 (N_14870,N_13289,N_12306);
nand U14871 (N_14871,N_12962,N_13471);
or U14872 (N_14872,N_13370,N_12757);
nor U14873 (N_14873,N_13186,N_12243);
and U14874 (N_14874,N_12949,N_12465);
and U14875 (N_14875,N_13417,N_12435);
and U14876 (N_14876,N_12409,N_12820);
nor U14877 (N_14877,N_12088,N_12326);
or U14878 (N_14878,N_12373,N_12308);
or U14879 (N_14879,N_12758,N_13300);
and U14880 (N_14880,N_12310,N_12576);
or U14881 (N_14881,N_12995,N_13083);
xnor U14882 (N_14882,N_12310,N_13062);
nor U14883 (N_14883,N_12798,N_12694);
and U14884 (N_14884,N_12831,N_13442);
nor U14885 (N_14885,N_12521,N_12055);
and U14886 (N_14886,N_12367,N_13268);
nor U14887 (N_14887,N_12339,N_12501);
nor U14888 (N_14888,N_12866,N_12544);
nor U14889 (N_14889,N_13039,N_12622);
or U14890 (N_14890,N_13275,N_13206);
nand U14891 (N_14891,N_13261,N_13180);
or U14892 (N_14892,N_12679,N_13467);
nor U14893 (N_14893,N_12859,N_12431);
and U14894 (N_14894,N_12153,N_12322);
and U14895 (N_14895,N_13182,N_12082);
or U14896 (N_14896,N_12934,N_13427);
or U14897 (N_14897,N_13100,N_13241);
and U14898 (N_14898,N_12126,N_12876);
nand U14899 (N_14899,N_13387,N_12805);
xnor U14900 (N_14900,N_12728,N_12521);
or U14901 (N_14901,N_12787,N_13174);
or U14902 (N_14902,N_13289,N_12426);
nand U14903 (N_14903,N_12045,N_12434);
nand U14904 (N_14904,N_12259,N_13089);
nand U14905 (N_14905,N_12819,N_12151);
or U14906 (N_14906,N_12478,N_12342);
nor U14907 (N_14907,N_12146,N_13189);
nand U14908 (N_14908,N_13167,N_12811);
nand U14909 (N_14909,N_13265,N_12293);
nor U14910 (N_14910,N_12943,N_12578);
xnor U14911 (N_14911,N_13027,N_13046);
or U14912 (N_14912,N_13068,N_12730);
nor U14913 (N_14913,N_13279,N_13286);
and U14914 (N_14914,N_13308,N_12269);
and U14915 (N_14915,N_12380,N_13320);
nor U14916 (N_14916,N_12098,N_12663);
nand U14917 (N_14917,N_13175,N_13293);
and U14918 (N_14918,N_12506,N_12556);
or U14919 (N_14919,N_12682,N_12229);
nor U14920 (N_14920,N_13005,N_13311);
nand U14921 (N_14921,N_12769,N_12034);
or U14922 (N_14922,N_12379,N_12203);
or U14923 (N_14923,N_12573,N_12670);
nor U14924 (N_14924,N_12061,N_13126);
and U14925 (N_14925,N_13367,N_12990);
nor U14926 (N_14926,N_12552,N_13091);
and U14927 (N_14927,N_13317,N_12404);
nor U14928 (N_14928,N_12620,N_12178);
and U14929 (N_14929,N_13398,N_12087);
or U14930 (N_14930,N_12620,N_12266);
nor U14931 (N_14931,N_13398,N_12731);
nor U14932 (N_14932,N_12584,N_12646);
xor U14933 (N_14933,N_12819,N_12668);
or U14934 (N_14934,N_12813,N_12142);
and U14935 (N_14935,N_12603,N_12358);
nor U14936 (N_14936,N_12676,N_12273);
nand U14937 (N_14937,N_13152,N_13020);
or U14938 (N_14938,N_13335,N_13210);
or U14939 (N_14939,N_12167,N_12099);
or U14940 (N_14940,N_13139,N_12289);
and U14941 (N_14941,N_12082,N_12194);
or U14942 (N_14942,N_13484,N_12933);
nor U14943 (N_14943,N_13259,N_12342);
or U14944 (N_14944,N_12270,N_12533);
or U14945 (N_14945,N_12752,N_12110);
nand U14946 (N_14946,N_13354,N_12690);
and U14947 (N_14947,N_12934,N_12584);
nand U14948 (N_14948,N_13272,N_12349);
or U14949 (N_14949,N_13222,N_12560);
nor U14950 (N_14950,N_12080,N_13091);
or U14951 (N_14951,N_12300,N_12692);
and U14952 (N_14952,N_12541,N_12720);
nor U14953 (N_14953,N_13216,N_13183);
and U14954 (N_14954,N_12815,N_13308);
and U14955 (N_14955,N_12842,N_13124);
or U14956 (N_14956,N_12152,N_13021);
and U14957 (N_14957,N_12927,N_13307);
or U14958 (N_14958,N_12385,N_12454);
or U14959 (N_14959,N_12270,N_13392);
or U14960 (N_14960,N_13310,N_12423);
nand U14961 (N_14961,N_12676,N_12649);
or U14962 (N_14962,N_12685,N_12363);
nand U14963 (N_14963,N_12053,N_12370);
nor U14964 (N_14964,N_12475,N_12777);
nand U14965 (N_14965,N_12333,N_13057);
nand U14966 (N_14966,N_12346,N_12711);
nor U14967 (N_14967,N_12135,N_13499);
nand U14968 (N_14968,N_12766,N_13464);
or U14969 (N_14969,N_12628,N_12256);
or U14970 (N_14970,N_13175,N_13278);
and U14971 (N_14971,N_12899,N_12297);
nor U14972 (N_14972,N_12003,N_12740);
nor U14973 (N_14973,N_12305,N_12223);
nand U14974 (N_14974,N_12598,N_12104);
nand U14975 (N_14975,N_12476,N_12587);
nand U14976 (N_14976,N_13091,N_12687);
nor U14977 (N_14977,N_13330,N_13345);
nand U14978 (N_14978,N_12286,N_12930);
nor U14979 (N_14979,N_12273,N_12049);
nor U14980 (N_14980,N_13010,N_12213);
or U14981 (N_14981,N_13428,N_12405);
or U14982 (N_14982,N_12329,N_13245);
nand U14983 (N_14983,N_13479,N_13105);
nand U14984 (N_14984,N_12290,N_12318);
nor U14985 (N_14985,N_12745,N_13037);
or U14986 (N_14986,N_12228,N_13430);
and U14987 (N_14987,N_13414,N_12068);
nand U14988 (N_14988,N_13022,N_12798);
nor U14989 (N_14989,N_12903,N_12961);
nor U14990 (N_14990,N_13178,N_12565);
nor U14991 (N_14991,N_12369,N_13050);
or U14992 (N_14992,N_12315,N_12000);
nand U14993 (N_14993,N_13075,N_13269);
nor U14994 (N_14994,N_12562,N_13228);
nor U14995 (N_14995,N_12930,N_13126);
and U14996 (N_14996,N_12558,N_12198);
nand U14997 (N_14997,N_12107,N_12074);
nor U14998 (N_14998,N_13264,N_12555);
or U14999 (N_14999,N_12938,N_12831);
nand UO_0 (O_0,N_13712,N_14742);
or UO_1 (O_1,N_14077,N_13881);
nor UO_2 (O_2,N_14531,N_13619);
nand UO_3 (O_3,N_14306,N_14540);
or UO_4 (O_4,N_14922,N_14165);
or UO_5 (O_5,N_13863,N_14498);
or UO_6 (O_6,N_14716,N_13890);
nand UO_7 (O_7,N_14856,N_14002);
and UO_8 (O_8,N_13629,N_13570);
or UO_9 (O_9,N_14224,N_13649);
and UO_10 (O_10,N_13675,N_14510);
nand UO_11 (O_11,N_14397,N_14894);
nand UO_12 (O_12,N_14217,N_13578);
or UO_13 (O_13,N_14288,N_14519);
nor UO_14 (O_14,N_14882,N_14652);
nand UO_15 (O_15,N_13746,N_14668);
nand UO_16 (O_16,N_14578,N_13818);
nor UO_17 (O_17,N_13513,N_14827);
or UO_18 (O_18,N_14683,N_13831);
nand UO_19 (O_19,N_14547,N_14718);
nand UO_20 (O_20,N_14130,N_14211);
or UO_21 (O_21,N_14817,N_14191);
and UO_22 (O_22,N_14596,N_13856);
xnor UO_23 (O_23,N_13534,N_14579);
or UO_24 (O_24,N_14842,N_14630);
nor UO_25 (O_25,N_14560,N_13916);
or UO_26 (O_26,N_14699,N_14163);
nor UO_27 (O_27,N_13545,N_14441);
nor UO_28 (O_28,N_14851,N_14651);
nand UO_29 (O_29,N_14686,N_14290);
nor UO_30 (O_30,N_14528,N_14685);
or UO_31 (O_31,N_14183,N_13820);
and UO_32 (O_32,N_13880,N_14773);
nand UO_33 (O_33,N_14634,N_13735);
nor UO_34 (O_34,N_13584,N_14705);
and UO_35 (O_35,N_13964,N_14226);
or UO_36 (O_36,N_14524,N_13718);
nor UO_37 (O_37,N_14957,N_14810);
or UO_38 (O_38,N_14327,N_14446);
and UO_39 (O_39,N_13620,N_13812);
nand UO_40 (O_40,N_14932,N_14990);
and UO_41 (O_41,N_14607,N_14299);
nand UO_42 (O_42,N_13983,N_14914);
nand UO_43 (O_43,N_14302,N_14335);
nor UO_44 (O_44,N_14366,N_14019);
nand UO_45 (O_45,N_13661,N_14247);
nand UO_46 (O_46,N_14762,N_14253);
nor UO_47 (O_47,N_14935,N_14076);
nor UO_48 (O_48,N_13908,N_14889);
nand UO_49 (O_49,N_14746,N_14362);
nand UO_50 (O_50,N_13806,N_13763);
nor UO_51 (O_51,N_13854,N_14166);
xor UO_52 (O_52,N_14044,N_14964);
nor UO_53 (O_53,N_14045,N_13689);
nor UO_54 (O_54,N_13679,N_14633);
and UO_55 (O_55,N_14172,N_14029);
or UO_56 (O_56,N_14244,N_14337);
nand UO_57 (O_57,N_13824,N_14920);
nor UO_58 (O_58,N_14317,N_13753);
and UO_59 (O_59,N_13760,N_13727);
or UO_60 (O_60,N_14860,N_14496);
or UO_61 (O_61,N_14318,N_13791);
or UO_62 (O_62,N_14050,N_14240);
or UO_63 (O_63,N_14774,N_14022);
or UO_64 (O_64,N_14344,N_13607);
and UO_65 (O_65,N_13776,N_14939);
nor UO_66 (O_66,N_14322,N_13569);
or UO_67 (O_67,N_14963,N_14636);
or UO_68 (O_68,N_13531,N_14180);
and UO_69 (O_69,N_14236,N_14698);
or UO_70 (O_70,N_14602,N_14262);
and UO_71 (O_71,N_13774,N_14612);
and UO_72 (O_72,N_14261,N_13590);
or UO_73 (O_73,N_13556,N_13621);
and UO_74 (O_74,N_14576,N_14499);
and UO_75 (O_75,N_14380,N_13747);
nor UO_76 (O_76,N_14311,N_13628);
nor UO_77 (O_77,N_14201,N_14987);
nand UO_78 (O_78,N_14071,N_14902);
nor UO_79 (O_79,N_14893,N_13794);
and UO_80 (O_80,N_13775,N_14493);
nand UO_81 (O_81,N_14783,N_13589);
nor UO_82 (O_82,N_13785,N_13742);
or UO_83 (O_83,N_13795,N_14800);
and UO_84 (O_84,N_14017,N_14459);
or UO_85 (O_85,N_14820,N_14843);
nand UO_86 (O_86,N_13648,N_13973);
and UO_87 (O_87,N_14557,N_14754);
or UO_88 (O_88,N_14532,N_14556);
or UO_89 (O_89,N_13547,N_13840);
nor UO_90 (O_90,N_14456,N_13886);
or UO_91 (O_91,N_14753,N_13662);
and UO_92 (O_92,N_14118,N_14844);
nand UO_93 (O_93,N_14927,N_14109);
nor UO_94 (O_94,N_14482,N_14156);
and UO_95 (O_95,N_13919,N_14066);
and UO_96 (O_96,N_14133,N_14890);
nor UO_97 (O_97,N_14016,N_14548);
and UO_98 (O_98,N_14874,N_14233);
nand UO_99 (O_99,N_13520,N_13700);
or UO_100 (O_100,N_14931,N_13814);
or UO_101 (O_101,N_13627,N_14792);
nand UO_102 (O_102,N_14878,N_14877);
nor UO_103 (O_103,N_14825,N_13713);
nor UO_104 (O_104,N_14582,N_13924);
nand UO_105 (O_105,N_13858,N_14151);
or UO_106 (O_106,N_14487,N_14449);
nor UO_107 (O_107,N_14372,N_13568);
nor UO_108 (O_108,N_13960,N_14907);
xnor UO_109 (O_109,N_14714,N_14631);
and UO_110 (O_110,N_14128,N_14309);
nand UO_111 (O_111,N_14134,N_13722);
and UO_112 (O_112,N_13910,N_13710);
or UO_113 (O_113,N_13626,N_14241);
nand UO_114 (O_114,N_13514,N_13725);
nand UO_115 (O_115,N_14808,N_14291);
nand UO_116 (O_116,N_13643,N_13929);
nor UO_117 (O_117,N_14996,N_13579);
and UO_118 (O_118,N_14178,N_14048);
nand UO_119 (O_119,N_13652,N_14719);
nor UO_120 (O_120,N_14912,N_14876);
xor UO_121 (O_121,N_14030,N_14841);
and UO_122 (O_122,N_14323,N_14120);
or UO_123 (O_123,N_14938,N_13839);
or UO_124 (O_124,N_13728,N_13934);
or UO_125 (O_125,N_13985,N_14517);
and UO_126 (O_126,N_14569,N_13507);
or UO_127 (O_127,N_13804,N_14729);
or UO_128 (O_128,N_14425,N_14770);
and UO_129 (O_129,N_14102,N_14896);
nand UO_130 (O_130,N_14084,N_14884);
and UO_131 (O_131,N_13731,N_14021);
or UO_132 (O_132,N_14757,N_13826);
nor UO_133 (O_133,N_14167,N_14953);
and UO_134 (O_134,N_13943,N_14189);
and UO_135 (O_135,N_13587,N_14554);
and UO_136 (O_136,N_14069,N_14514);
nand UO_137 (O_137,N_14563,N_14671);
and UO_138 (O_138,N_14260,N_13810);
and UO_139 (O_139,N_13878,N_14955);
nor UO_140 (O_140,N_14307,N_14732);
nand UO_141 (O_141,N_13936,N_14779);
or UO_142 (O_142,N_14092,N_14586);
nand UO_143 (O_143,N_14834,N_14750);
and UO_144 (O_144,N_14188,N_14003);
nand UO_145 (O_145,N_14011,N_13622);
nand UO_146 (O_146,N_13846,N_14570);
nor UO_147 (O_147,N_14433,N_14155);
and UO_148 (O_148,N_14251,N_14766);
nor UO_149 (O_149,N_14505,N_14369);
and UO_150 (O_150,N_14845,N_14515);
and UO_151 (O_151,N_13549,N_14013);
and UO_152 (O_152,N_14930,N_13623);
or UO_153 (O_153,N_14246,N_14041);
or UO_154 (O_154,N_14836,N_14315);
and UO_155 (O_155,N_14078,N_14124);
nor UO_156 (O_156,N_14606,N_14678);
or UO_157 (O_157,N_14897,N_14175);
nor UO_158 (O_158,N_14662,N_14007);
nand UO_159 (O_159,N_14743,N_13615);
nor UO_160 (O_160,N_14345,N_13743);
and UO_161 (O_161,N_14734,N_14488);
nand UO_162 (O_162,N_14553,N_14873);
nor UO_163 (O_163,N_13571,N_14802);
nand UO_164 (O_164,N_14292,N_14936);
nand UO_165 (O_165,N_14919,N_13935);
nor UO_166 (O_166,N_14974,N_14584);
nand UO_167 (O_167,N_13738,N_13502);
nand UO_168 (O_168,N_14075,N_13769);
nand UO_169 (O_169,N_14072,N_14129);
or UO_170 (O_170,N_14485,N_13918);
or UO_171 (O_171,N_14853,N_14564);
nand UO_172 (O_172,N_14502,N_13773);
or UO_173 (O_173,N_14014,N_14739);
and UO_174 (O_174,N_13896,N_14414);
nor UO_175 (O_175,N_13690,N_14983);
nor UO_176 (O_176,N_14395,N_13759);
and UO_177 (O_177,N_14872,N_14168);
nand UO_178 (O_178,N_14985,N_14095);
nor UO_179 (O_179,N_13975,N_14803);
nand UO_180 (O_180,N_14279,N_13640);
nor UO_181 (O_181,N_14006,N_13741);
nor UO_182 (O_182,N_13749,N_14467);
or UO_183 (O_183,N_14921,N_14535);
or UO_184 (O_184,N_14127,N_14212);
nand UO_185 (O_185,N_14759,N_13971);
and UO_186 (O_186,N_14815,N_14207);
or UO_187 (O_187,N_14094,N_14160);
nor UO_188 (O_188,N_13530,N_14284);
and UO_189 (O_189,N_13697,N_13696);
nor UO_190 (O_190,N_13512,N_14255);
nor UO_191 (O_191,N_13517,N_13724);
nand UO_192 (O_192,N_14360,N_14644);
nand UO_193 (O_193,N_14899,N_13860);
and UO_194 (O_194,N_14658,N_13865);
nor UO_195 (O_195,N_13944,N_14703);
nand UO_196 (O_196,N_13974,N_14767);
nand UO_197 (O_197,N_14138,N_14994);
nand UO_198 (O_198,N_13827,N_14649);
nor UO_199 (O_199,N_13551,N_14629);
or UO_200 (O_200,N_14616,N_13913);
nand UO_201 (O_201,N_14351,N_14988);
nor UO_202 (O_202,N_14501,N_14057);
nand UO_203 (O_203,N_14096,N_13683);
or UO_204 (O_204,N_13548,N_13630);
and UO_205 (O_205,N_14799,N_14545);
and UO_206 (O_206,N_14484,N_14239);
or UO_207 (O_207,N_13909,N_14981);
nand UO_208 (O_208,N_14313,N_14677);
and UO_209 (O_209,N_13976,N_13601);
or UO_210 (O_210,N_13602,N_14653);
and UO_211 (O_211,N_14438,N_14023);
or UO_212 (O_212,N_13966,N_13585);
and UO_213 (O_213,N_14132,N_14628);
or UO_214 (O_214,N_13819,N_14647);
nor UO_215 (O_215,N_13647,N_14620);
or UO_216 (O_216,N_14837,N_14061);
nor UO_217 (O_217,N_13981,N_14525);
or UO_218 (O_218,N_14506,N_14551);
nand UO_219 (O_219,N_14982,N_13844);
nand UO_220 (O_220,N_14150,N_14424);
nor UO_221 (O_221,N_14355,N_14674);
and UO_222 (O_222,N_14812,N_14354);
nor UO_223 (O_223,N_13750,N_13947);
or UO_224 (O_224,N_14926,N_14418);
nand UO_225 (O_225,N_14148,N_14198);
or UO_226 (O_226,N_13594,N_13667);
and UO_227 (O_227,N_14934,N_14585);
and UO_228 (O_228,N_14141,N_14403);
and UO_229 (O_229,N_13616,N_14377);
or UO_230 (O_230,N_13891,N_14363);
nor UO_231 (O_231,N_14452,N_14552);
and UO_232 (O_232,N_14135,N_13907);
and UO_233 (O_233,N_14225,N_13631);
nand UO_234 (O_234,N_14826,N_14243);
nand UO_235 (O_235,N_14608,N_14451);
nor UO_236 (O_236,N_13893,N_14149);
or UO_237 (O_237,N_14474,N_13565);
nor UO_238 (O_238,N_13635,N_13861);
nand UO_239 (O_239,N_14303,N_13838);
and UO_240 (O_240,N_13555,N_14070);
and UO_241 (O_241,N_14090,N_13633);
nor UO_242 (O_242,N_13949,N_14371);
and UO_243 (O_243,N_14818,N_13799);
nor UO_244 (O_244,N_13748,N_14656);
nor UO_245 (O_245,N_14806,N_14059);
nor UO_246 (O_246,N_14654,N_13639);
nand UO_247 (O_247,N_14062,N_14642);
nor UO_248 (O_248,N_13836,N_14571);
nand UO_249 (O_249,N_13539,N_14724);
or UO_250 (O_250,N_13942,N_14434);
and UO_251 (O_251,N_14618,N_13613);
nand UO_252 (O_252,N_14237,N_13522);
nand UO_253 (O_253,N_14301,N_14319);
and UO_254 (O_254,N_14170,N_13906);
and UO_255 (O_255,N_13752,N_14330);
nor UO_256 (O_256,N_13686,N_13707);
nor UO_257 (O_257,N_13636,N_13811);
nand UO_258 (O_258,N_14108,N_13925);
or UO_259 (O_259,N_13702,N_14305);
nor UO_260 (O_260,N_13659,N_14063);
or UO_261 (O_261,N_14232,N_14966);
or UO_262 (O_262,N_14694,N_14264);
or UO_263 (O_263,N_14392,N_14892);
nor UO_264 (O_264,N_14436,N_13876);
and UO_265 (O_265,N_14031,N_13766);
or UO_266 (O_266,N_13699,N_14886);
nor UO_267 (O_267,N_14000,N_14598);
nand UO_268 (O_268,N_14967,N_14831);
nand UO_269 (O_269,N_14619,N_14866);
nor UO_270 (O_270,N_14638,N_14708);
nor UO_271 (O_271,N_14087,N_14727);
and UO_272 (O_272,N_13991,N_13848);
or UO_273 (O_273,N_14416,N_14854);
or UO_274 (O_274,N_14187,N_14913);
or UO_275 (O_275,N_14869,N_14676);
or UO_276 (O_276,N_14033,N_14943);
nand UO_277 (O_277,N_14895,N_13542);
and UO_278 (O_278,N_14641,N_13870);
or UO_279 (O_279,N_14942,N_13573);
or UO_280 (O_280,N_14526,N_14669);
nand UO_281 (O_281,N_13701,N_14503);
and UO_282 (O_282,N_14796,N_14153);
or UO_283 (O_283,N_14911,N_14946);
and UO_284 (O_284,N_14468,N_14435);
or UO_285 (O_285,N_14546,N_13955);
or UO_286 (O_286,N_14483,N_14404);
nor UO_287 (O_287,N_14600,N_14804);
and UO_288 (O_288,N_14389,N_14736);
and UO_289 (O_289,N_13789,N_14763);
nand UO_290 (O_290,N_14223,N_13708);
and UO_291 (O_291,N_14326,N_14680);
or UO_292 (O_292,N_14152,N_14756);
or UO_293 (O_293,N_14206,N_14965);
or UO_294 (O_294,N_14793,N_14572);
or UO_295 (O_295,N_13611,N_13845);
and UO_296 (O_296,N_14807,N_14537);
nand UO_297 (O_297,N_14621,N_14368);
nand UO_298 (O_298,N_14916,N_14480);
xnor UO_299 (O_299,N_13898,N_14209);
or UO_300 (O_300,N_14738,N_13581);
nor UO_301 (O_301,N_14373,N_14347);
nand UO_302 (O_302,N_13656,N_14511);
nand UO_303 (O_303,N_14972,N_14702);
and UO_304 (O_304,N_14681,N_13676);
nor UO_305 (O_305,N_14005,N_14272);
nor UO_306 (O_306,N_14390,N_14463);
and UO_307 (O_307,N_14382,N_13998);
or UO_308 (O_308,N_14768,N_14879);
and UO_309 (O_309,N_14682,N_13755);
nor UO_310 (O_310,N_14394,N_14276);
and UO_311 (O_311,N_13957,N_14508);
nand UO_312 (O_312,N_13723,N_14971);
and UO_313 (O_313,N_13688,N_13600);
nand UO_314 (O_314,N_14056,N_14234);
and UO_315 (O_315,N_14402,N_14868);
or UO_316 (O_316,N_14847,N_14772);
nor UO_317 (O_317,N_14701,N_13516);
and UO_318 (O_318,N_13550,N_14666);
and UO_319 (O_319,N_14464,N_14962);
or UO_320 (O_320,N_14864,N_14871);
nor UO_321 (O_321,N_14374,N_14364);
nand UO_322 (O_322,N_13698,N_14115);
and UO_323 (O_323,N_13945,N_14399);
and UO_324 (O_324,N_14018,N_13681);
and UO_325 (O_325,N_13829,N_14901);
or UO_326 (O_326,N_13851,N_14158);
nand UO_327 (O_327,N_13855,N_13801);
nor UO_328 (O_328,N_14639,N_14422);
or UO_329 (O_329,N_14959,N_13521);
nand UO_330 (O_330,N_14604,N_13901);
and UO_331 (O_331,N_13754,N_13808);
and UO_332 (O_332,N_14945,N_13946);
and UO_333 (O_333,N_13536,N_14393);
and UO_334 (O_334,N_13927,N_14590);
nor UO_335 (O_335,N_13694,N_14089);
nor UO_336 (O_336,N_14909,N_14358);
and UO_337 (O_337,N_14980,N_13950);
nor UO_338 (O_338,N_14448,N_14038);
and UO_339 (O_339,N_14164,N_14405);
nor UO_340 (O_340,N_14867,N_13761);
nand UO_341 (O_341,N_14862,N_13889);
or UO_342 (O_342,N_13882,N_14093);
nor UO_343 (O_343,N_14849,N_14162);
nand UO_344 (O_344,N_14082,N_13937);
nand UO_345 (O_345,N_14771,N_14123);
nor UO_346 (O_346,N_14192,N_14915);
and UO_347 (O_347,N_14067,N_14737);
nor UO_348 (O_348,N_13872,N_14733);
or UO_349 (O_349,N_13798,N_13897);
or UO_350 (O_350,N_13711,N_13892);
nor UO_351 (O_351,N_13511,N_14544);
nand UO_352 (O_352,N_14139,N_13693);
or UO_353 (O_353,N_13519,N_14906);
and UO_354 (O_354,N_14352,N_13610);
or UO_355 (O_355,N_14489,N_14083);
and UO_356 (O_356,N_13745,N_13980);
nand UO_357 (O_357,N_13771,N_13797);
nand UO_358 (O_358,N_14214,N_14320);
or UO_359 (O_359,N_14529,N_13654);
or UO_360 (O_360,N_14850,N_13560);
or UO_361 (O_361,N_14052,N_14780);
nand UO_362 (O_362,N_13952,N_14523);
nand UO_363 (O_363,N_14785,N_14710);
nor UO_364 (O_364,N_14367,N_14898);
or UO_365 (O_365,N_14199,N_14880);
or UO_366 (O_366,N_14462,N_14855);
nor UO_367 (O_367,N_14784,N_14891);
or UO_368 (O_368,N_14024,N_13715);
nor UO_369 (O_369,N_14473,N_14396);
nand UO_370 (O_370,N_13997,N_14058);
nand UO_371 (O_371,N_13767,N_14200);
nor UO_372 (O_372,N_14614,N_14781);
or UO_373 (O_373,N_13650,N_14098);
and UO_374 (O_374,N_14176,N_13895);
or UO_375 (O_375,N_14970,N_14695);
nor UO_376 (O_376,N_14238,N_13503);
or UO_377 (O_377,N_14297,N_14581);
nand UO_378 (O_378,N_14221,N_14624);
nor UO_379 (O_379,N_14749,N_14865);
or UO_380 (O_380,N_14637,N_14944);
nor UO_381 (O_381,N_14903,N_14775);
and UO_382 (O_382,N_14491,N_13540);
nand UO_383 (O_383,N_14177,N_14043);
or UO_384 (O_384,N_14110,N_13692);
nor UO_385 (O_385,N_13672,N_14020);
or UO_386 (O_386,N_13885,N_14379);
and UO_387 (O_387,N_14137,N_13515);
nand UO_388 (O_388,N_14388,N_14925);
or UO_389 (O_389,N_14472,N_14242);
nor UO_390 (O_390,N_14998,N_14343);
nand UO_391 (O_391,N_13657,N_14755);
and UO_392 (O_392,N_14740,N_14648);
and UO_393 (O_393,N_14193,N_14386);
and UO_394 (O_394,N_13821,N_14341);
nand UO_395 (O_395,N_13967,N_14444);
or UO_396 (O_396,N_13670,N_13866);
nor UO_397 (O_397,N_14977,N_13655);
and UO_398 (O_398,N_13716,N_13671);
or UO_399 (O_399,N_14885,N_14053);
or UO_400 (O_400,N_14601,N_13730);
and UO_401 (O_401,N_13911,N_14310);
nor UO_402 (O_402,N_14426,N_13900);
nand UO_403 (O_403,N_14409,N_13920);
nand UO_404 (O_404,N_13951,N_13765);
nand UO_405 (O_405,N_14136,N_14412);
nor UO_406 (O_406,N_14179,N_14659);
nor UO_407 (O_407,N_14114,N_14333);
or UO_408 (O_408,N_14227,N_13786);
and UO_409 (O_409,N_14574,N_14252);
and UO_410 (O_410,N_14248,N_14125);
nand UO_411 (O_411,N_14027,N_14764);
and UO_412 (O_412,N_13884,N_14777);
or UO_413 (O_413,N_14445,N_13958);
nor UO_414 (O_414,N_13835,N_13720);
nor UO_415 (O_415,N_14004,N_13687);
nor UO_416 (O_416,N_14720,N_13574);
nor UO_417 (O_417,N_13717,N_13782);
nor UO_418 (O_418,N_14431,N_13930);
nor UO_419 (O_419,N_14408,N_13703);
nor UO_420 (O_420,N_14010,N_14336);
and UO_421 (O_421,N_14481,N_14265);
nand UO_422 (O_422,N_14460,N_14492);
nor UO_423 (O_423,N_13779,N_14204);
and UO_424 (O_424,N_14324,N_14900);
and UO_425 (O_425,N_14692,N_14555);
or UO_426 (O_426,N_14410,N_13847);
nor UO_427 (O_427,N_13928,N_14427);
nor UO_428 (O_428,N_14859,N_14747);
or UO_429 (O_429,N_14790,N_13658);
or UO_430 (O_430,N_14278,N_14542);
or UO_431 (O_431,N_14910,N_13537);
and UO_432 (O_432,N_13841,N_13803);
and UO_433 (O_433,N_14101,N_14250);
nor UO_434 (O_434,N_14144,N_14952);
nor UO_435 (O_435,N_13558,N_14593);
or UO_436 (O_436,N_14042,N_13962);
nand UO_437 (O_437,N_14507,N_13500);
or UO_438 (O_438,N_14028,N_13714);
and UO_439 (O_439,N_13988,N_14561);
nand UO_440 (O_440,N_14951,N_14329);
nand UO_441 (O_441,N_14116,N_14331);
or UO_442 (O_442,N_14186,N_13862);
or UO_443 (O_443,N_13805,N_14384);
nor UO_444 (O_444,N_13857,N_13526);
nor UO_445 (O_445,N_13993,N_13682);
nor UO_446 (O_446,N_14839,N_13781);
or UO_447 (O_447,N_14821,N_13546);
nor UO_448 (O_448,N_14989,N_14049);
nand UO_449 (O_449,N_14956,N_14157);
or UO_450 (O_450,N_13783,N_14249);
and UO_451 (O_451,N_14627,N_14625);
nor UO_452 (O_452,N_14254,N_13843);
or UO_453 (O_453,N_13637,N_13674);
nor UO_454 (O_454,N_14263,N_14174);
nand UO_455 (O_455,N_14673,N_13625);
nor UO_456 (O_456,N_14091,N_13948);
and UO_457 (O_457,N_14591,N_14937);
nand UO_458 (O_458,N_14992,N_14142);
or UO_459 (O_459,N_14428,N_14566);
nor UO_460 (O_460,N_13653,N_13523);
nor UO_461 (O_461,N_14287,N_14086);
and UO_462 (O_462,N_14470,N_13923);
or UO_463 (O_463,N_14640,N_14184);
nand UO_464 (O_464,N_13850,N_13543);
nand UO_465 (O_465,N_14840,N_13984);
nor UO_466 (O_466,N_13926,N_13931);
nor UO_467 (O_467,N_14979,N_14940);
and UO_468 (O_468,N_13796,N_13953);
nand UO_469 (O_469,N_14280,N_14823);
nor UO_470 (O_470,N_14423,N_14266);
or UO_471 (O_471,N_14154,N_14104);
or UO_472 (O_472,N_13664,N_13562);
or UO_473 (O_473,N_14245,N_13978);
nor UO_474 (O_474,N_14672,N_14968);
or UO_475 (O_475,N_13849,N_13505);
or UO_476 (O_476,N_13504,N_14328);
nand UO_477 (O_477,N_14978,N_13852);
and UO_478 (O_478,N_14219,N_13595);
nand UO_479 (O_479,N_14210,N_14228);
nand UO_480 (O_480,N_14852,N_14617);
and UO_481 (O_481,N_14999,N_14034);
and UO_482 (O_482,N_14811,N_13915);
nor UO_483 (O_483,N_13894,N_14690);
xnor UO_484 (O_484,N_13875,N_13591);
nor UO_485 (O_485,N_14081,N_13588);
or UO_486 (O_486,N_14285,N_13739);
or UO_487 (O_487,N_13566,N_14991);
and UO_488 (O_488,N_14858,N_14294);
and UO_489 (O_489,N_14450,N_14819);
nand UO_490 (O_490,N_14465,N_14430);
nand UO_491 (O_491,N_13559,N_14447);
or UO_492 (O_492,N_13992,N_14295);
and UO_493 (O_493,N_13904,N_13704);
and UO_494 (O_494,N_14097,N_14721);
nand UO_495 (O_495,N_13995,N_13859);
or UO_496 (O_496,N_13762,N_14594);
and UO_497 (O_497,N_13583,N_14696);
or UO_498 (O_498,N_13941,N_13816);
and UO_499 (O_499,N_13614,N_14469);
nand UO_500 (O_500,N_14829,N_13986);
nand UO_501 (O_501,N_14623,N_14832);
nor UO_502 (O_502,N_14235,N_13641);
and UO_503 (O_503,N_14530,N_14222);
nor UO_504 (O_504,N_14281,N_13645);
nor UO_505 (O_505,N_14486,N_14975);
or UO_506 (O_506,N_14300,N_14776);
and UO_507 (O_507,N_14597,N_14039);
and UO_508 (O_508,N_14615,N_13634);
nand UO_509 (O_509,N_14745,N_14413);
and UO_510 (O_510,N_14924,N_14997);
nand UO_511 (O_511,N_14587,N_14271);
nand UO_512 (O_512,N_14202,N_14929);
and UO_513 (O_513,N_14259,N_14182);
and UO_514 (O_514,N_14933,N_14411);
or UO_515 (O_515,N_13832,N_13580);
nor UO_516 (O_516,N_14230,N_14918);
nor UO_517 (O_517,N_13970,N_14522);
nor UO_518 (O_518,N_14205,N_13586);
or UO_519 (O_519,N_14798,N_14442);
nor UO_520 (O_520,N_14609,N_14687);
nor UO_521 (O_521,N_14559,N_14870);
or UO_522 (O_522,N_13666,N_14376);
nor UO_523 (O_523,N_14008,N_13939);
and UO_524 (O_524,N_14385,N_14477);
and UO_525 (O_525,N_14035,N_14357);
or UO_526 (O_526,N_14976,N_13669);
nor UO_527 (O_527,N_13758,N_14904);
and UO_528 (O_528,N_14375,N_14282);
nand UO_529 (O_529,N_14941,N_14119);
nand UO_530 (O_530,N_14700,N_13564);
nor UO_531 (O_531,N_13987,N_14969);
nand UO_532 (O_532,N_14947,N_14613);
or UO_533 (O_533,N_13940,N_13969);
or UO_534 (O_534,N_14605,N_14478);
and UO_535 (O_535,N_14171,N_13533);
nor UO_536 (O_536,N_13576,N_14443);
or UO_537 (O_537,N_14679,N_14797);
nand UO_538 (O_538,N_14466,N_14117);
or UO_539 (O_539,N_14905,N_13879);
nand UO_540 (O_540,N_14316,N_13706);
nor UO_541 (O_541,N_13557,N_13778);
or UO_542 (O_542,N_14356,N_14269);
nand UO_543 (O_543,N_13651,N_14986);
nand UO_544 (O_544,N_13777,N_13695);
nor UO_545 (O_545,N_13632,N_13554);
and UO_546 (O_546,N_14813,N_14711);
and UO_547 (O_547,N_14312,N_13788);
nor UO_548 (O_548,N_14643,N_13938);
nand UO_549 (O_549,N_14054,N_14103);
and UO_550 (O_550,N_14748,N_14541);
nand UO_551 (O_551,N_13599,N_14208);
nand UO_552 (O_552,N_14401,N_14213);
nand UO_553 (O_553,N_13665,N_14398);
or UO_554 (O_554,N_13990,N_14814);
nor UO_555 (O_555,N_14454,N_14744);
nand UO_556 (O_556,N_14495,N_14025);
or UO_557 (O_557,N_14500,N_14830);
nor UO_558 (O_558,N_14599,N_14824);
nand UO_559 (O_559,N_14074,N_14381);
nor UO_560 (O_560,N_14107,N_14848);
or UO_561 (O_561,N_14846,N_14461);
nor UO_562 (O_562,N_13660,N_13740);
nand UO_563 (O_563,N_14215,N_14661);
or UO_564 (O_564,N_14112,N_14549);
nor UO_565 (O_565,N_14610,N_14195);
nand UO_566 (O_566,N_14715,N_14314);
nand UO_567 (O_567,N_14709,N_13751);
nor UO_568 (O_568,N_13677,N_14805);
nor UO_569 (O_569,N_14726,N_14664);
or UO_570 (O_570,N_14816,N_14741);
nor UO_571 (O_571,N_13606,N_14274);
nor UO_572 (O_572,N_14420,N_14595);
nand UO_573 (O_573,N_14592,N_14961);
xnor UO_574 (O_574,N_13853,N_14194);
nor UO_575 (O_575,N_14065,N_14875);
and UO_576 (O_576,N_13994,N_14917);
nor UO_577 (O_577,N_13837,N_14688);
nand UO_578 (O_578,N_13552,N_13528);
and UO_579 (O_579,N_14220,N_14973);
or UO_580 (O_580,N_14432,N_14655);
nand UO_581 (O_581,N_14203,N_13609);
and UO_582 (O_582,N_13617,N_14346);
nor UO_583 (O_583,N_13646,N_14835);
or UO_584 (O_584,N_14100,N_14348);
nand UO_585 (O_585,N_14415,N_14181);
or UO_586 (O_586,N_14378,N_14752);
nor UO_587 (O_587,N_14550,N_13541);
or UO_588 (O_588,N_13644,N_14713);
and UO_589 (O_589,N_13527,N_14521);
or UO_590 (O_590,N_14960,N_13871);
xnor UO_591 (O_591,N_14778,N_13705);
or UO_592 (O_592,N_14185,N_14760);
nor UO_593 (O_593,N_14801,N_14289);
nor UO_594 (O_594,N_14349,N_14993);
nor UO_595 (O_595,N_13917,N_13977);
nand UO_596 (O_596,N_14332,N_13518);
or UO_597 (O_597,N_14321,N_14995);
nor UO_598 (O_598,N_14122,N_13638);
nand UO_599 (O_599,N_14789,N_13834);
and UO_600 (O_600,N_14504,N_14196);
and UO_601 (O_601,N_14888,N_14458);
and UO_602 (O_602,N_14632,N_14169);
nand UO_603 (O_603,N_14573,N_14575);
nand UO_604 (O_604,N_14457,N_13510);
or UO_605 (O_605,N_14286,N_14717);
and UO_606 (O_606,N_13800,N_14334);
nor UO_607 (O_607,N_13965,N_14417);
nor UO_608 (O_608,N_14562,N_13532);
nand UO_609 (O_609,N_14693,N_14543);
and UO_610 (O_610,N_14769,N_14490);
nand UO_611 (O_611,N_13887,N_14455);
nor UO_612 (O_612,N_14140,N_14794);
and UO_613 (O_613,N_14229,N_14113);
xnor UO_614 (O_614,N_14660,N_13729);
and UO_615 (O_615,N_14051,N_13603);
nand UO_616 (O_616,N_14722,N_13921);
nand UO_617 (O_617,N_14383,N_13642);
nand UO_618 (O_618,N_14626,N_14475);
and UO_619 (O_619,N_14231,N_14786);
nor UO_620 (O_620,N_13793,N_13868);
nand UO_621 (O_621,N_14040,N_13737);
nor UO_622 (O_622,N_14338,N_14948);
or UO_623 (O_623,N_14161,N_14047);
nand UO_624 (O_624,N_14015,N_14131);
nand UO_625 (O_625,N_14603,N_14536);
or UO_626 (O_626,N_14984,N_14787);
and UO_627 (O_627,N_13721,N_13501);
nand UO_628 (O_628,N_14589,N_13593);
nand UO_629 (O_629,N_14611,N_14512);
and UO_630 (O_630,N_13932,N_14293);
nand UO_631 (O_631,N_14106,N_13605);
nor UO_632 (O_632,N_13678,N_13506);
nor UO_633 (O_633,N_13525,N_13572);
nand UO_634 (O_634,N_14111,N_14928);
or UO_635 (O_635,N_13509,N_13903);
nand UO_636 (O_636,N_13809,N_14667);
and UO_637 (O_637,N_13912,N_14419);
or UO_638 (O_638,N_14268,N_13813);
or UO_639 (O_639,N_13673,N_13979);
nand UO_640 (O_640,N_14731,N_14675);
nor UO_641 (O_641,N_14080,N_13732);
nor UO_642 (O_642,N_14725,N_14064);
and UO_643 (O_643,N_14126,N_14365);
or UO_644 (O_644,N_14147,N_14538);
nand UO_645 (O_645,N_14577,N_13922);
or UO_646 (O_646,N_14340,N_13902);
or UO_647 (O_647,N_14256,N_14159);
or UO_648 (O_648,N_13538,N_14706);
nand UO_649 (O_649,N_13764,N_14908);
nand UO_650 (O_650,N_14751,N_14439);
nand UO_651 (O_651,N_14697,N_14001);
nand UO_652 (O_652,N_13817,N_14958);
nor UO_653 (O_653,N_13582,N_13597);
and UO_654 (O_654,N_14646,N_14509);
and UO_655 (O_655,N_13888,N_13663);
nor UO_656 (O_656,N_13757,N_13982);
or UO_657 (O_657,N_13596,N_13604);
nand UO_658 (O_658,N_14520,N_13823);
or UO_659 (O_659,N_13864,N_14949);
and UO_660 (O_660,N_14622,N_14650);
or UO_661 (O_661,N_14881,N_13685);
and UO_662 (O_662,N_14568,N_13736);
nor UO_663 (O_663,N_14684,N_14361);
xnor UO_664 (O_664,N_14273,N_13989);
or UO_665 (O_665,N_14534,N_13999);
nand UO_666 (O_666,N_14437,N_14099);
nand UO_667 (O_667,N_14421,N_13784);
and UO_668 (O_668,N_14822,N_13833);
nor UO_669 (O_669,N_14350,N_13575);
nand UO_670 (O_670,N_13956,N_14406);
or UO_671 (O_671,N_14765,N_14954);
nand UO_672 (O_672,N_14707,N_14105);
or UO_673 (O_673,N_14275,N_13544);
and UO_674 (O_674,N_13933,N_13961);
and UO_675 (O_675,N_14216,N_13772);
and UO_676 (O_676,N_13592,N_13873);
nand UO_677 (O_677,N_14788,N_14723);
nor UO_678 (O_678,N_14863,N_14277);
nor UO_679 (O_679,N_13802,N_13842);
or UO_680 (O_680,N_13815,N_13529);
or UO_681 (O_681,N_14296,N_14085);
and UO_682 (O_682,N_13954,N_14453);
or UO_683 (O_683,N_13905,N_13959);
or UO_684 (O_684,N_14791,N_14258);
and UO_685 (O_685,N_14645,N_14391);
or UO_686 (O_686,N_14190,N_14146);
and UO_687 (O_687,N_14479,N_14012);
nand UO_688 (O_688,N_13770,N_13691);
or UO_689 (O_689,N_14055,N_14588);
or UO_690 (O_690,N_14670,N_13792);
or UO_691 (O_691,N_14663,N_14689);
or UO_692 (O_692,N_14838,N_13553);
and UO_693 (O_693,N_13822,N_13624);
nor UO_694 (O_694,N_14565,N_14009);
or UO_695 (O_695,N_14567,N_14121);
and UO_696 (O_696,N_13963,N_13867);
or UO_697 (O_697,N_14518,N_14060);
and UO_698 (O_698,N_14068,N_14143);
or UO_699 (O_699,N_14429,N_13869);
nor UO_700 (O_700,N_13996,N_14036);
or UO_701 (O_701,N_13830,N_14861);
nand UO_702 (O_702,N_14197,N_14325);
and UO_703 (O_703,N_13719,N_14883);
and UO_704 (O_704,N_13787,N_14298);
nand UO_705 (O_705,N_13877,N_14353);
nand UO_706 (O_706,N_14032,N_13524);
xor UO_707 (O_707,N_14387,N_14712);
nor UO_708 (O_708,N_13567,N_14471);
or UO_709 (O_709,N_14073,N_13598);
xor UO_710 (O_710,N_14476,N_14359);
and UO_711 (O_711,N_13608,N_13828);
nand UO_712 (O_712,N_14950,N_14407);
and UO_713 (O_713,N_13734,N_14539);
nor UO_714 (O_714,N_14857,N_13968);
nand UO_715 (O_715,N_13508,N_13874);
nor UO_716 (O_716,N_14761,N_13744);
nor UO_717 (O_717,N_14267,N_14923);
nand UO_718 (O_718,N_13618,N_14339);
and UO_719 (O_719,N_14580,N_13563);
nand UO_720 (O_720,N_14735,N_13825);
and UO_721 (O_721,N_14728,N_13684);
and UO_722 (O_722,N_14513,N_14527);
nor UO_723 (O_723,N_14887,N_14173);
or UO_724 (O_724,N_13577,N_14145);
or UO_725 (O_725,N_14782,N_13726);
xor UO_726 (O_726,N_13709,N_14046);
nor UO_727 (O_727,N_13680,N_13790);
nand UO_728 (O_728,N_14704,N_14758);
or UO_729 (O_729,N_14691,N_13668);
nor UO_730 (O_730,N_13561,N_14440);
and UO_731 (O_731,N_13914,N_13733);
and UO_732 (O_732,N_14270,N_13535);
or UO_733 (O_733,N_13756,N_14283);
and UO_734 (O_734,N_14304,N_14400);
or UO_735 (O_735,N_14809,N_13899);
nor UO_736 (O_736,N_14342,N_14583);
or UO_737 (O_737,N_14730,N_14665);
nor UO_738 (O_738,N_14558,N_14657);
nor UO_739 (O_739,N_14026,N_13807);
nor UO_740 (O_740,N_14533,N_13883);
or UO_741 (O_741,N_13780,N_14516);
xnor UO_742 (O_742,N_14079,N_13612);
nor UO_743 (O_743,N_14088,N_14497);
nand UO_744 (O_744,N_14257,N_13972);
and UO_745 (O_745,N_14308,N_14218);
nor UO_746 (O_746,N_14828,N_13768);
nand UO_747 (O_747,N_14037,N_14370);
nand UO_748 (O_748,N_14833,N_14795);
nand UO_749 (O_749,N_14494,N_14635);
nand UO_750 (O_750,N_13714,N_14169);
or UO_751 (O_751,N_14580,N_13843);
and UO_752 (O_752,N_14133,N_14997);
nor UO_753 (O_753,N_13675,N_13684);
nor UO_754 (O_754,N_13595,N_13625);
nor UO_755 (O_755,N_14587,N_13734);
and UO_756 (O_756,N_14695,N_13529);
or UO_757 (O_757,N_13998,N_13993);
nand UO_758 (O_758,N_14446,N_14586);
nand UO_759 (O_759,N_14959,N_14436);
and UO_760 (O_760,N_14575,N_13777);
nor UO_761 (O_761,N_13892,N_13960);
nand UO_762 (O_762,N_13574,N_14543);
xnor UO_763 (O_763,N_14403,N_14036);
nand UO_764 (O_764,N_14962,N_13862);
nand UO_765 (O_765,N_14411,N_13677);
and UO_766 (O_766,N_14845,N_14092);
nand UO_767 (O_767,N_14977,N_14791);
nor UO_768 (O_768,N_14441,N_14453);
nand UO_769 (O_769,N_14188,N_13846);
nand UO_770 (O_770,N_14949,N_14599);
nor UO_771 (O_771,N_14754,N_13803);
nand UO_772 (O_772,N_13789,N_14858);
and UO_773 (O_773,N_14191,N_13623);
nor UO_774 (O_774,N_14295,N_14456);
or UO_775 (O_775,N_14375,N_13807);
and UO_776 (O_776,N_14897,N_14503);
nand UO_777 (O_777,N_14966,N_14017);
and UO_778 (O_778,N_14209,N_13585);
or UO_779 (O_779,N_14517,N_14798);
and UO_780 (O_780,N_13615,N_14118);
nand UO_781 (O_781,N_14756,N_14690);
xor UO_782 (O_782,N_13981,N_13697);
nor UO_783 (O_783,N_14289,N_14884);
nor UO_784 (O_784,N_14792,N_13532);
nor UO_785 (O_785,N_14105,N_14291);
and UO_786 (O_786,N_13740,N_14901);
nor UO_787 (O_787,N_14262,N_14403);
nor UO_788 (O_788,N_14053,N_14530);
nand UO_789 (O_789,N_14722,N_14339);
and UO_790 (O_790,N_13839,N_13778);
nor UO_791 (O_791,N_13516,N_14200);
xnor UO_792 (O_792,N_14608,N_14812);
nor UO_793 (O_793,N_14948,N_14127);
or UO_794 (O_794,N_13631,N_14171);
nor UO_795 (O_795,N_14684,N_13687);
nor UO_796 (O_796,N_14356,N_14313);
xor UO_797 (O_797,N_14789,N_13531);
nor UO_798 (O_798,N_14821,N_14481);
and UO_799 (O_799,N_14246,N_14413);
nor UO_800 (O_800,N_14691,N_13897);
and UO_801 (O_801,N_14130,N_14026);
and UO_802 (O_802,N_14683,N_13988);
nand UO_803 (O_803,N_14127,N_14010);
and UO_804 (O_804,N_13659,N_14394);
and UO_805 (O_805,N_14323,N_14012);
and UO_806 (O_806,N_14896,N_14441);
or UO_807 (O_807,N_14252,N_14422);
or UO_808 (O_808,N_13800,N_14028);
and UO_809 (O_809,N_14110,N_14296);
or UO_810 (O_810,N_14771,N_13965);
or UO_811 (O_811,N_13954,N_14055);
or UO_812 (O_812,N_13846,N_13988);
and UO_813 (O_813,N_13861,N_13946);
and UO_814 (O_814,N_14479,N_14787);
and UO_815 (O_815,N_13594,N_13852);
nor UO_816 (O_816,N_14914,N_13986);
nand UO_817 (O_817,N_14224,N_14390);
or UO_818 (O_818,N_14307,N_14347);
nor UO_819 (O_819,N_13962,N_14430);
or UO_820 (O_820,N_14047,N_13657);
nor UO_821 (O_821,N_13793,N_14674);
nand UO_822 (O_822,N_14936,N_13772);
nand UO_823 (O_823,N_14429,N_14741);
nor UO_824 (O_824,N_13746,N_13807);
and UO_825 (O_825,N_14700,N_14825);
nand UO_826 (O_826,N_14837,N_14389);
xor UO_827 (O_827,N_13779,N_14128);
or UO_828 (O_828,N_14231,N_13684);
or UO_829 (O_829,N_13883,N_14706);
or UO_830 (O_830,N_14840,N_14054);
nand UO_831 (O_831,N_14021,N_14312);
and UO_832 (O_832,N_14644,N_13522);
and UO_833 (O_833,N_14664,N_13744);
nand UO_834 (O_834,N_14565,N_13759);
and UO_835 (O_835,N_14772,N_13862);
and UO_836 (O_836,N_14952,N_13979);
or UO_837 (O_837,N_14704,N_13936);
nand UO_838 (O_838,N_13553,N_14111);
or UO_839 (O_839,N_14503,N_14479);
or UO_840 (O_840,N_13809,N_14271);
or UO_841 (O_841,N_14783,N_14709);
or UO_842 (O_842,N_13811,N_14494);
or UO_843 (O_843,N_14528,N_14906);
nand UO_844 (O_844,N_13673,N_14218);
nor UO_845 (O_845,N_13603,N_13722);
nor UO_846 (O_846,N_13988,N_13886);
or UO_847 (O_847,N_13937,N_13984);
and UO_848 (O_848,N_13784,N_14465);
or UO_849 (O_849,N_14318,N_13763);
nand UO_850 (O_850,N_13579,N_13932);
or UO_851 (O_851,N_14533,N_14013);
nand UO_852 (O_852,N_13856,N_14961);
or UO_853 (O_853,N_13589,N_14482);
nor UO_854 (O_854,N_14305,N_14501);
nand UO_855 (O_855,N_13812,N_14501);
nand UO_856 (O_856,N_14124,N_14452);
nor UO_857 (O_857,N_13724,N_14339);
or UO_858 (O_858,N_14171,N_14442);
and UO_859 (O_859,N_14746,N_14982);
nand UO_860 (O_860,N_14236,N_14585);
nand UO_861 (O_861,N_14286,N_13901);
nor UO_862 (O_862,N_14299,N_14172);
and UO_863 (O_863,N_14230,N_14225);
nor UO_864 (O_864,N_14699,N_13638);
xor UO_865 (O_865,N_14054,N_13672);
xnor UO_866 (O_866,N_13905,N_13714);
nor UO_867 (O_867,N_14031,N_14055);
and UO_868 (O_868,N_14264,N_14895);
nand UO_869 (O_869,N_14392,N_14053);
or UO_870 (O_870,N_14929,N_14385);
or UO_871 (O_871,N_14598,N_14329);
nor UO_872 (O_872,N_14118,N_13504);
or UO_873 (O_873,N_13996,N_14804);
nor UO_874 (O_874,N_13691,N_13509);
and UO_875 (O_875,N_13760,N_13519);
nor UO_876 (O_876,N_14845,N_14417);
nor UO_877 (O_877,N_14892,N_13573);
nor UO_878 (O_878,N_14373,N_13624);
nand UO_879 (O_879,N_14896,N_14897);
or UO_880 (O_880,N_14534,N_14702);
or UO_881 (O_881,N_14922,N_13532);
and UO_882 (O_882,N_14723,N_14717);
nand UO_883 (O_883,N_14184,N_13965);
nor UO_884 (O_884,N_13567,N_13551);
nor UO_885 (O_885,N_14516,N_14687);
nor UO_886 (O_886,N_13904,N_13537);
or UO_887 (O_887,N_14973,N_13745);
or UO_888 (O_888,N_13679,N_13633);
and UO_889 (O_889,N_13772,N_14663);
nand UO_890 (O_890,N_14021,N_14119);
and UO_891 (O_891,N_14749,N_14472);
and UO_892 (O_892,N_13619,N_14491);
nor UO_893 (O_893,N_14648,N_14606);
and UO_894 (O_894,N_13810,N_13724);
or UO_895 (O_895,N_13547,N_14565);
or UO_896 (O_896,N_14855,N_13608);
or UO_897 (O_897,N_14011,N_14865);
and UO_898 (O_898,N_13812,N_14171);
nor UO_899 (O_899,N_14251,N_13932);
nor UO_900 (O_900,N_14546,N_14633);
and UO_901 (O_901,N_14851,N_14336);
nor UO_902 (O_902,N_14803,N_13783);
and UO_903 (O_903,N_14639,N_14971);
and UO_904 (O_904,N_13925,N_13837);
or UO_905 (O_905,N_14262,N_14081);
nor UO_906 (O_906,N_14570,N_14315);
or UO_907 (O_907,N_14488,N_14206);
or UO_908 (O_908,N_14274,N_13852);
nand UO_909 (O_909,N_13527,N_14824);
and UO_910 (O_910,N_13665,N_14538);
and UO_911 (O_911,N_14629,N_13725);
nand UO_912 (O_912,N_13919,N_14242);
nor UO_913 (O_913,N_13793,N_14394);
nand UO_914 (O_914,N_13694,N_14379);
nor UO_915 (O_915,N_13560,N_13970);
nand UO_916 (O_916,N_14609,N_14717);
and UO_917 (O_917,N_14080,N_14655);
and UO_918 (O_918,N_14846,N_13903);
or UO_919 (O_919,N_14658,N_14874);
nand UO_920 (O_920,N_14863,N_14056);
nand UO_921 (O_921,N_14488,N_14236);
nor UO_922 (O_922,N_14813,N_13661);
nor UO_923 (O_923,N_14869,N_13555);
nor UO_924 (O_924,N_14924,N_14785);
nor UO_925 (O_925,N_14730,N_14469);
or UO_926 (O_926,N_13640,N_13736);
nor UO_927 (O_927,N_14413,N_13861);
nor UO_928 (O_928,N_14190,N_13617);
or UO_929 (O_929,N_14402,N_13886);
nand UO_930 (O_930,N_14939,N_13940);
and UO_931 (O_931,N_14777,N_14750);
and UO_932 (O_932,N_14142,N_14212);
nand UO_933 (O_933,N_14352,N_14519);
or UO_934 (O_934,N_14995,N_13700);
nand UO_935 (O_935,N_14062,N_13889);
nand UO_936 (O_936,N_14154,N_14832);
nor UO_937 (O_937,N_14122,N_14872);
and UO_938 (O_938,N_14862,N_13665);
nand UO_939 (O_939,N_14477,N_13683);
or UO_940 (O_940,N_13798,N_14094);
or UO_941 (O_941,N_14527,N_13580);
and UO_942 (O_942,N_14810,N_14950);
nor UO_943 (O_943,N_14524,N_14260);
nor UO_944 (O_944,N_14235,N_14550);
or UO_945 (O_945,N_14439,N_13659);
nand UO_946 (O_946,N_13850,N_14248);
and UO_947 (O_947,N_14374,N_14939);
or UO_948 (O_948,N_14694,N_13544);
and UO_949 (O_949,N_14012,N_14875);
nor UO_950 (O_950,N_14242,N_13899);
nand UO_951 (O_951,N_13699,N_13538);
or UO_952 (O_952,N_13743,N_14190);
or UO_953 (O_953,N_14064,N_14731);
nand UO_954 (O_954,N_14272,N_13507);
nand UO_955 (O_955,N_13894,N_14374);
nand UO_956 (O_956,N_14787,N_13557);
xnor UO_957 (O_957,N_14014,N_13868);
nor UO_958 (O_958,N_13829,N_14767);
nand UO_959 (O_959,N_14455,N_13684);
nand UO_960 (O_960,N_14208,N_13611);
and UO_961 (O_961,N_14965,N_14565);
xnor UO_962 (O_962,N_13560,N_14821);
and UO_963 (O_963,N_14734,N_13956);
nand UO_964 (O_964,N_14704,N_14485);
nand UO_965 (O_965,N_13864,N_14459);
nand UO_966 (O_966,N_14903,N_14300);
or UO_967 (O_967,N_14289,N_14446);
nand UO_968 (O_968,N_14242,N_14104);
nand UO_969 (O_969,N_14032,N_14941);
nor UO_970 (O_970,N_14189,N_14563);
nor UO_971 (O_971,N_13573,N_14788);
and UO_972 (O_972,N_13957,N_14095);
nor UO_973 (O_973,N_14349,N_14991);
nand UO_974 (O_974,N_14065,N_13798);
and UO_975 (O_975,N_14877,N_13985);
nor UO_976 (O_976,N_13647,N_14604);
nor UO_977 (O_977,N_14654,N_14820);
nand UO_978 (O_978,N_13691,N_13546);
nor UO_979 (O_979,N_14388,N_13694);
or UO_980 (O_980,N_14936,N_13602);
and UO_981 (O_981,N_14483,N_14886);
and UO_982 (O_982,N_14220,N_14440);
or UO_983 (O_983,N_13855,N_14826);
nand UO_984 (O_984,N_14461,N_14628);
nor UO_985 (O_985,N_14998,N_14496);
or UO_986 (O_986,N_13910,N_14127);
and UO_987 (O_987,N_14646,N_14970);
nand UO_988 (O_988,N_14176,N_14122);
or UO_989 (O_989,N_14606,N_14017);
nand UO_990 (O_990,N_14794,N_14691);
and UO_991 (O_991,N_14880,N_14758);
and UO_992 (O_992,N_13502,N_13935);
and UO_993 (O_993,N_14733,N_14471);
and UO_994 (O_994,N_13685,N_13849);
nand UO_995 (O_995,N_14765,N_13808);
and UO_996 (O_996,N_14028,N_14865);
or UO_997 (O_997,N_14468,N_14568);
or UO_998 (O_998,N_14620,N_14277);
or UO_999 (O_999,N_13995,N_14759);
or UO_1000 (O_1000,N_14655,N_14141);
nor UO_1001 (O_1001,N_14762,N_14916);
nand UO_1002 (O_1002,N_13618,N_14310);
or UO_1003 (O_1003,N_14836,N_14541);
or UO_1004 (O_1004,N_14174,N_14864);
nand UO_1005 (O_1005,N_13832,N_13751);
nand UO_1006 (O_1006,N_14732,N_14626);
and UO_1007 (O_1007,N_13901,N_13537);
nand UO_1008 (O_1008,N_13847,N_13820);
and UO_1009 (O_1009,N_14363,N_14262);
or UO_1010 (O_1010,N_14235,N_13731);
and UO_1011 (O_1011,N_14185,N_14558);
or UO_1012 (O_1012,N_13842,N_14409);
and UO_1013 (O_1013,N_14367,N_13607);
nor UO_1014 (O_1014,N_14933,N_14406);
and UO_1015 (O_1015,N_14508,N_14946);
nor UO_1016 (O_1016,N_14691,N_14115);
or UO_1017 (O_1017,N_13537,N_14353);
nor UO_1018 (O_1018,N_14995,N_14942);
and UO_1019 (O_1019,N_13785,N_14707);
nor UO_1020 (O_1020,N_14670,N_14645);
nand UO_1021 (O_1021,N_14260,N_14791);
or UO_1022 (O_1022,N_14992,N_14565);
nor UO_1023 (O_1023,N_14580,N_14096);
and UO_1024 (O_1024,N_13569,N_14296);
and UO_1025 (O_1025,N_14352,N_14912);
nand UO_1026 (O_1026,N_14766,N_14764);
nor UO_1027 (O_1027,N_14838,N_14962);
nor UO_1028 (O_1028,N_14809,N_14205);
or UO_1029 (O_1029,N_14360,N_14137);
and UO_1030 (O_1030,N_14591,N_14335);
nor UO_1031 (O_1031,N_14413,N_13503);
and UO_1032 (O_1032,N_13734,N_14072);
and UO_1033 (O_1033,N_14916,N_14834);
or UO_1034 (O_1034,N_13968,N_14778);
or UO_1035 (O_1035,N_13527,N_14799);
nand UO_1036 (O_1036,N_13744,N_14010);
or UO_1037 (O_1037,N_14149,N_14174);
nand UO_1038 (O_1038,N_14002,N_14083);
nor UO_1039 (O_1039,N_14871,N_14420);
nor UO_1040 (O_1040,N_13911,N_14412);
nand UO_1041 (O_1041,N_14403,N_14234);
nor UO_1042 (O_1042,N_14043,N_14594);
nand UO_1043 (O_1043,N_13607,N_14307);
or UO_1044 (O_1044,N_13677,N_14708);
and UO_1045 (O_1045,N_14917,N_14720);
or UO_1046 (O_1046,N_14940,N_13606);
or UO_1047 (O_1047,N_13690,N_14142);
and UO_1048 (O_1048,N_14615,N_13999);
nor UO_1049 (O_1049,N_13673,N_14431);
and UO_1050 (O_1050,N_13525,N_14514);
and UO_1051 (O_1051,N_14624,N_14173);
or UO_1052 (O_1052,N_13592,N_14380);
nand UO_1053 (O_1053,N_14646,N_14797);
and UO_1054 (O_1054,N_14729,N_14294);
nand UO_1055 (O_1055,N_14968,N_13641);
nand UO_1056 (O_1056,N_14796,N_13947);
and UO_1057 (O_1057,N_14559,N_14258);
nand UO_1058 (O_1058,N_13663,N_14807);
nand UO_1059 (O_1059,N_14593,N_13762);
nor UO_1060 (O_1060,N_14792,N_14554);
nor UO_1061 (O_1061,N_14092,N_14598);
or UO_1062 (O_1062,N_14614,N_14995);
nor UO_1063 (O_1063,N_13847,N_14777);
or UO_1064 (O_1064,N_13543,N_14248);
nand UO_1065 (O_1065,N_13552,N_14306);
nor UO_1066 (O_1066,N_14457,N_14594);
and UO_1067 (O_1067,N_13597,N_14088);
or UO_1068 (O_1068,N_14385,N_13651);
nand UO_1069 (O_1069,N_14856,N_14478);
or UO_1070 (O_1070,N_13712,N_14062);
or UO_1071 (O_1071,N_14098,N_13516);
nand UO_1072 (O_1072,N_14882,N_14691);
and UO_1073 (O_1073,N_13516,N_14147);
or UO_1074 (O_1074,N_13712,N_14384);
or UO_1075 (O_1075,N_14107,N_13618);
nor UO_1076 (O_1076,N_14895,N_13918);
or UO_1077 (O_1077,N_14465,N_14514);
nor UO_1078 (O_1078,N_14973,N_14051);
nand UO_1079 (O_1079,N_14878,N_14959);
or UO_1080 (O_1080,N_14646,N_14717);
and UO_1081 (O_1081,N_14623,N_14030);
nor UO_1082 (O_1082,N_13992,N_14545);
xor UO_1083 (O_1083,N_14483,N_14367);
nor UO_1084 (O_1084,N_14924,N_13814);
xor UO_1085 (O_1085,N_13732,N_13518);
or UO_1086 (O_1086,N_14991,N_14942);
nor UO_1087 (O_1087,N_14840,N_14150);
or UO_1088 (O_1088,N_14459,N_13571);
and UO_1089 (O_1089,N_14171,N_14072);
or UO_1090 (O_1090,N_14203,N_14721);
nand UO_1091 (O_1091,N_14555,N_13671);
nand UO_1092 (O_1092,N_14328,N_14967);
or UO_1093 (O_1093,N_13792,N_13682);
and UO_1094 (O_1094,N_13700,N_14905);
or UO_1095 (O_1095,N_13833,N_13872);
and UO_1096 (O_1096,N_14729,N_13811);
nor UO_1097 (O_1097,N_14149,N_14307);
nor UO_1098 (O_1098,N_14018,N_14779);
nand UO_1099 (O_1099,N_14495,N_14157);
and UO_1100 (O_1100,N_14923,N_14721);
nor UO_1101 (O_1101,N_14461,N_14855);
nor UO_1102 (O_1102,N_14475,N_14259);
nor UO_1103 (O_1103,N_14876,N_14466);
and UO_1104 (O_1104,N_13896,N_14473);
or UO_1105 (O_1105,N_14406,N_13528);
and UO_1106 (O_1106,N_14986,N_14407);
nor UO_1107 (O_1107,N_14066,N_14388);
nor UO_1108 (O_1108,N_13748,N_14355);
nand UO_1109 (O_1109,N_14480,N_14505);
and UO_1110 (O_1110,N_13869,N_14220);
nand UO_1111 (O_1111,N_13552,N_14796);
or UO_1112 (O_1112,N_14985,N_14294);
nor UO_1113 (O_1113,N_14796,N_14832);
and UO_1114 (O_1114,N_14254,N_13619);
nor UO_1115 (O_1115,N_14157,N_13869);
nand UO_1116 (O_1116,N_14824,N_13687);
and UO_1117 (O_1117,N_13914,N_14624);
or UO_1118 (O_1118,N_14072,N_14032);
and UO_1119 (O_1119,N_14185,N_14046);
or UO_1120 (O_1120,N_14898,N_13572);
nor UO_1121 (O_1121,N_13782,N_14696);
and UO_1122 (O_1122,N_14167,N_14686);
xnor UO_1123 (O_1123,N_13674,N_14053);
nor UO_1124 (O_1124,N_14580,N_13567);
or UO_1125 (O_1125,N_13676,N_14195);
nand UO_1126 (O_1126,N_14959,N_14317);
or UO_1127 (O_1127,N_14857,N_14443);
nor UO_1128 (O_1128,N_14399,N_14115);
or UO_1129 (O_1129,N_14788,N_14329);
or UO_1130 (O_1130,N_14389,N_14109);
nand UO_1131 (O_1131,N_14675,N_14209);
or UO_1132 (O_1132,N_14277,N_13801);
and UO_1133 (O_1133,N_13549,N_14444);
nor UO_1134 (O_1134,N_13706,N_14560);
nor UO_1135 (O_1135,N_14984,N_14012);
nand UO_1136 (O_1136,N_14719,N_13641);
or UO_1137 (O_1137,N_14645,N_14250);
or UO_1138 (O_1138,N_13989,N_14679);
nor UO_1139 (O_1139,N_14284,N_14909);
nor UO_1140 (O_1140,N_14591,N_14269);
and UO_1141 (O_1141,N_14659,N_14136);
or UO_1142 (O_1142,N_14351,N_14000);
nor UO_1143 (O_1143,N_14424,N_14800);
and UO_1144 (O_1144,N_14959,N_14782);
or UO_1145 (O_1145,N_13512,N_14371);
and UO_1146 (O_1146,N_13625,N_14380);
nand UO_1147 (O_1147,N_14061,N_14468);
nor UO_1148 (O_1148,N_14473,N_14423);
nand UO_1149 (O_1149,N_14591,N_14433);
nand UO_1150 (O_1150,N_14514,N_14366);
nand UO_1151 (O_1151,N_14896,N_14707);
and UO_1152 (O_1152,N_14079,N_14837);
nand UO_1153 (O_1153,N_14795,N_14445);
nand UO_1154 (O_1154,N_14166,N_14763);
or UO_1155 (O_1155,N_14224,N_14758);
nand UO_1156 (O_1156,N_13580,N_14795);
nand UO_1157 (O_1157,N_14527,N_14156);
nand UO_1158 (O_1158,N_13739,N_14990);
or UO_1159 (O_1159,N_14635,N_14531);
nor UO_1160 (O_1160,N_13999,N_14329);
and UO_1161 (O_1161,N_14442,N_13882);
nand UO_1162 (O_1162,N_14615,N_14200);
or UO_1163 (O_1163,N_14871,N_14244);
or UO_1164 (O_1164,N_13611,N_14297);
nand UO_1165 (O_1165,N_13919,N_14015);
nor UO_1166 (O_1166,N_13736,N_14240);
nand UO_1167 (O_1167,N_14677,N_14925);
and UO_1168 (O_1168,N_14260,N_13643);
nand UO_1169 (O_1169,N_14879,N_14956);
and UO_1170 (O_1170,N_13683,N_13990);
or UO_1171 (O_1171,N_14339,N_14488);
or UO_1172 (O_1172,N_13905,N_13831);
or UO_1173 (O_1173,N_14166,N_14159);
nand UO_1174 (O_1174,N_14892,N_14198);
or UO_1175 (O_1175,N_14758,N_14975);
xor UO_1176 (O_1176,N_13503,N_13533);
nor UO_1177 (O_1177,N_14564,N_14332);
or UO_1178 (O_1178,N_14920,N_13512);
or UO_1179 (O_1179,N_13875,N_13982);
nand UO_1180 (O_1180,N_13939,N_14333);
nand UO_1181 (O_1181,N_14480,N_13526);
or UO_1182 (O_1182,N_14614,N_14906);
or UO_1183 (O_1183,N_13974,N_14540);
or UO_1184 (O_1184,N_14459,N_14438);
nor UO_1185 (O_1185,N_13930,N_14810);
nor UO_1186 (O_1186,N_14336,N_14051);
and UO_1187 (O_1187,N_14421,N_13985);
nor UO_1188 (O_1188,N_14538,N_14817);
or UO_1189 (O_1189,N_14375,N_14219);
nand UO_1190 (O_1190,N_13645,N_14208);
and UO_1191 (O_1191,N_14849,N_14952);
and UO_1192 (O_1192,N_13768,N_13525);
and UO_1193 (O_1193,N_14775,N_14526);
or UO_1194 (O_1194,N_14177,N_13987);
nor UO_1195 (O_1195,N_14620,N_14204);
nand UO_1196 (O_1196,N_14468,N_14770);
nand UO_1197 (O_1197,N_14948,N_13716);
and UO_1198 (O_1198,N_14384,N_14333);
or UO_1199 (O_1199,N_14575,N_13797);
nand UO_1200 (O_1200,N_14566,N_14473);
nor UO_1201 (O_1201,N_14189,N_14271);
and UO_1202 (O_1202,N_14893,N_13953);
or UO_1203 (O_1203,N_13751,N_14547);
or UO_1204 (O_1204,N_14615,N_14367);
or UO_1205 (O_1205,N_14682,N_14955);
or UO_1206 (O_1206,N_14074,N_13935);
nand UO_1207 (O_1207,N_14924,N_14609);
or UO_1208 (O_1208,N_13536,N_14582);
or UO_1209 (O_1209,N_13879,N_14179);
nor UO_1210 (O_1210,N_14916,N_14751);
and UO_1211 (O_1211,N_13645,N_14080);
nor UO_1212 (O_1212,N_13860,N_14878);
and UO_1213 (O_1213,N_13584,N_14957);
or UO_1214 (O_1214,N_14505,N_13763);
or UO_1215 (O_1215,N_14211,N_13850);
or UO_1216 (O_1216,N_14663,N_13561);
or UO_1217 (O_1217,N_14029,N_13605);
nor UO_1218 (O_1218,N_13964,N_14217);
and UO_1219 (O_1219,N_14951,N_13587);
nor UO_1220 (O_1220,N_14117,N_14169);
or UO_1221 (O_1221,N_14387,N_14265);
and UO_1222 (O_1222,N_14485,N_14707);
nand UO_1223 (O_1223,N_14365,N_14132);
nor UO_1224 (O_1224,N_13748,N_14523);
nor UO_1225 (O_1225,N_14319,N_13878);
nor UO_1226 (O_1226,N_13511,N_13554);
nor UO_1227 (O_1227,N_14050,N_14937);
and UO_1228 (O_1228,N_14431,N_14085);
and UO_1229 (O_1229,N_13726,N_14299);
and UO_1230 (O_1230,N_14036,N_13693);
or UO_1231 (O_1231,N_14720,N_14566);
and UO_1232 (O_1232,N_14837,N_13680);
or UO_1233 (O_1233,N_13593,N_14076);
nor UO_1234 (O_1234,N_14693,N_14915);
nor UO_1235 (O_1235,N_14114,N_13774);
and UO_1236 (O_1236,N_14315,N_13853);
nor UO_1237 (O_1237,N_14636,N_13967);
nor UO_1238 (O_1238,N_14041,N_14331);
nor UO_1239 (O_1239,N_13960,N_14888);
or UO_1240 (O_1240,N_14683,N_14135);
nand UO_1241 (O_1241,N_13846,N_14291);
nor UO_1242 (O_1242,N_14149,N_14081);
nand UO_1243 (O_1243,N_13732,N_14803);
nor UO_1244 (O_1244,N_14954,N_13706);
or UO_1245 (O_1245,N_14148,N_13562);
nand UO_1246 (O_1246,N_14403,N_13757);
nor UO_1247 (O_1247,N_14941,N_13597);
or UO_1248 (O_1248,N_14715,N_13885);
and UO_1249 (O_1249,N_13960,N_14537);
or UO_1250 (O_1250,N_13838,N_14929);
and UO_1251 (O_1251,N_14464,N_13741);
nor UO_1252 (O_1252,N_13770,N_14438);
nand UO_1253 (O_1253,N_14661,N_14426);
or UO_1254 (O_1254,N_14900,N_14241);
and UO_1255 (O_1255,N_14780,N_13923);
or UO_1256 (O_1256,N_13668,N_14378);
and UO_1257 (O_1257,N_14391,N_14069);
nand UO_1258 (O_1258,N_13935,N_14457);
nor UO_1259 (O_1259,N_14971,N_14939);
nor UO_1260 (O_1260,N_13776,N_14123);
and UO_1261 (O_1261,N_14203,N_14042);
and UO_1262 (O_1262,N_14738,N_14039);
and UO_1263 (O_1263,N_14237,N_14866);
or UO_1264 (O_1264,N_13822,N_13571);
or UO_1265 (O_1265,N_13648,N_13726);
or UO_1266 (O_1266,N_13800,N_14481);
nor UO_1267 (O_1267,N_13780,N_14997);
and UO_1268 (O_1268,N_13903,N_14631);
nor UO_1269 (O_1269,N_14153,N_14346);
or UO_1270 (O_1270,N_13809,N_14491);
or UO_1271 (O_1271,N_14326,N_14996);
nor UO_1272 (O_1272,N_13603,N_13817);
nor UO_1273 (O_1273,N_14806,N_14065);
or UO_1274 (O_1274,N_14397,N_14318);
and UO_1275 (O_1275,N_14438,N_14497);
nor UO_1276 (O_1276,N_14080,N_14257);
and UO_1277 (O_1277,N_14710,N_13644);
nand UO_1278 (O_1278,N_14352,N_14586);
and UO_1279 (O_1279,N_13836,N_14464);
and UO_1280 (O_1280,N_14157,N_14208);
and UO_1281 (O_1281,N_14431,N_14888);
nor UO_1282 (O_1282,N_14485,N_14962);
xnor UO_1283 (O_1283,N_13924,N_13657);
nand UO_1284 (O_1284,N_13726,N_14753);
or UO_1285 (O_1285,N_13825,N_14461);
xnor UO_1286 (O_1286,N_14092,N_13837);
nor UO_1287 (O_1287,N_14573,N_13776);
nand UO_1288 (O_1288,N_14026,N_14286);
and UO_1289 (O_1289,N_13690,N_14775);
nand UO_1290 (O_1290,N_14336,N_13804);
nor UO_1291 (O_1291,N_14610,N_14570);
or UO_1292 (O_1292,N_14677,N_14720);
nand UO_1293 (O_1293,N_14173,N_14761);
nand UO_1294 (O_1294,N_13872,N_13781);
nand UO_1295 (O_1295,N_14191,N_14350);
nand UO_1296 (O_1296,N_14093,N_14294);
nor UO_1297 (O_1297,N_14729,N_14651);
and UO_1298 (O_1298,N_14933,N_14663);
and UO_1299 (O_1299,N_13673,N_14243);
and UO_1300 (O_1300,N_14686,N_14429);
nor UO_1301 (O_1301,N_14492,N_13568);
or UO_1302 (O_1302,N_14021,N_14009);
nor UO_1303 (O_1303,N_14539,N_13766);
nand UO_1304 (O_1304,N_14989,N_13824);
nor UO_1305 (O_1305,N_13764,N_13762);
nor UO_1306 (O_1306,N_13961,N_14803);
nor UO_1307 (O_1307,N_14500,N_13567);
or UO_1308 (O_1308,N_13650,N_14689);
nand UO_1309 (O_1309,N_14685,N_14715);
or UO_1310 (O_1310,N_13658,N_14915);
and UO_1311 (O_1311,N_13643,N_14065);
nor UO_1312 (O_1312,N_14447,N_14874);
nor UO_1313 (O_1313,N_13802,N_13940);
nor UO_1314 (O_1314,N_14737,N_13986);
nand UO_1315 (O_1315,N_14110,N_13794);
nand UO_1316 (O_1316,N_14285,N_14932);
nor UO_1317 (O_1317,N_13875,N_14314);
and UO_1318 (O_1318,N_14966,N_14168);
or UO_1319 (O_1319,N_13501,N_14365);
nor UO_1320 (O_1320,N_13526,N_13792);
nor UO_1321 (O_1321,N_13800,N_13813);
or UO_1322 (O_1322,N_14150,N_14990);
nor UO_1323 (O_1323,N_13734,N_14185);
and UO_1324 (O_1324,N_14422,N_14631);
nor UO_1325 (O_1325,N_14966,N_14452);
or UO_1326 (O_1326,N_13509,N_14853);
nor UO_1327 (O_1327,N_14392,N_14951);
nand UO_1328 (O_1328,N_13741,N_14458);
or UO_1329 (O_1329,N_14064,N_13871);
and UO_1330 (O_1330,N_14208,N_14065);
and UO_1331 (O_1331,N_14780,N_14335);
or UO_1332 (O_1332,N_14083,N_14075);
nor UO_1333 (O_1333,N_13620,N_13524);
and UO_1334 (O_1334,N_14598,N_14424);
or UO_1335 (O_1335,N_14036,N_14307);
and UO_1336 (O_1336,N_14290,N_14164);
nor UO_1337 (O_1337,N_14551,N_14973);
and UO_1338 (O_1338,N_14738,N_14424);
and UO_1339 (O_1339,N_13925,N_13620);
nand UO_1340 (O_1340,N_14158,N_14223);
and UO_1341 (O_1341,N_14047,N_13568);
nor UO_1342 (O_1342,N_14674,N_14059);
nand UO_1343 (O_1343,N_13625,N_14585);
nand UO_1344 (O_1344,N_13993,N_14495);
nor UO_1345 (O_1345,N_14035,N_14291);
nand UO_1346 (O_1346,N_14354,N_14832);
nor UO_1347 (O_1347,N_14398,N_14773);
nand UO_1348 (O_1348,N_14680,N_14378);
or UO_1349 (O_1349,N_13551,N_14579);
and UO_1350 (O_1350,N_13668,N_14010);
or UO_1351 (O_1351,N_14363,N_14091);
nor UO_1352 (O_1352,N_14626,N_14020);
nand UO_1353 (O_1353,N_14770,N_13537);
or UO_1354 (O_1354,N_13969,N_13727);
nand UO_1355 (O_1355,N_14691,N_14006);
or UO_1356 (O_1356,N_14757,N_14858);
xor UO_1357 (O_1357,N_14420,N_14425);
or UO_1358 (O_1358,N_14848,N_14845);
and UO_1359 (O_1359,N_14336,N_14210);
or UO_1360 (O_1360,N_13773,N_14118);
and UO_1361 (O_1361,N_13653,N_13521);
and UO_1362 (O_1362,N_14730,N_14677);
or UO_1363 (O_1363,N_14320,N_13923);
or UO_1364 (O_1364,N_14416,N_13827);
or UO_1365 (O_1365,N_13619,N_13845);
nand UO_1366 (O_1366,N_14263,N_13728);
or UO_1367 (O_1367,N_14283,N_14147);
nor UO_1368 (O_1368,N_14457,N_14649);
nor UO_1369 (O_1369,N_14268,N_14549);
and UO_1370 (O_1370,N_14211,N_14423);
or UO_1371 (O_1371,N_14372,N_14132);
nor UO_1372 (O_1372,N_14941,N_13978);
and UO_1373 (O_1373,N_14579,N_14057);
nand UO_1374 (O_1374,N_14781,N_13813);
or UO_1375 (O_1375,N_14325,N_14695);
or UO_1376 (O_1376,N_13748,N_13796);
nor UO_1377 (O_1377,N_14950,N_13873);
and UO_1378 (O_1378,N_13828,N_14768);
or UO_1379 (O_1379,N_13822,N_14677);
nand UO_1380 (O_1380,N_14241,N_13547);
or UO_1381 (O_1381,N_13915,N_14384);
nor UO_1382 (O_1382,N_13552,N_13916);
and UO_1383 (O_1383,N_14938,N_14130);
and UO_1384 (O_1384,N_14183,N_13831);
or UO_1385 (O_1385,N_14670,N_14301);
and UO_1386 (O_1386,N_14836,N_13551);
nand UO_1387 (O_1387,N_13551,N_14733);
and UO_1388 (O_1388,N_14365,N_14210);
or UO_1389 (O_1389,N_13532,N_13822);
xor UO_1390 (O_1390,N_14950,N_13933);
nand UO_1391 (O_1391,N_14312,N_14782);
nor UO_1392 (O_1392,N_13973,N_13721);
nor UO_1393 (O_1393,N_13581,N_14205);
and UO_1394 (O_1394,N_14203,N_14509);
nand UO_1395 (O_1395,N_14389,N_14593);
or UO_1396 (O_1396,N_13528,N_14031);
nor UO_1397 (O_1397,N_13500,N_13771);
nand UO_1398 (O_1398,N_14087,N_14565);
or UO_1399 (O_1399,N_14838,N_14945);
or UO_1400 (O_1400,N_14212,N_14954);
or UO_1401 (O_1401,N_13923,N_14515);
nand UO_1402 (O_1402,N_14350,N_14290);
and UO_1403 (O_1403,N_14379,N_14478);
nand UO_1404 (O_1404,N_14608,N_14500);
nand UO_1405 (O_1405,N_14779,N_13974);
xor UO_1406 (O_1406,N_14577,N_14698);
nor UO_1407 (O_1407,N_14015,N_14506);
and UO_1408 (O_1408,N_14609,N_14182);
or UO_1409 (O_1409,N_14374,N_14195);
and UO_1410 (O_1410,N_14538,N_14924);
or UO_1411 (O_1411,N_14843,N_13859);
nor UO_1412 (O_1412,N_14129,N_14748);
or UO_1413 (O_1413,N_14087,N_13949);
or UO_1414 (O_1414,N_14646,N_14467);
or UO_1415 (O_1415,N_13784,N_14230);
nor UO_1416 (O_1416,N_14939,N_13602);
nor UO_1417 (O_1417,N_14848,N_13970);
and UO_1418 (O_1418,N_13722,N_14291);
or UO_1419 (O_1419,N_13937,N_13545);
or UO_1420 (O_1420,N_14168,N_14738);
and UO_1421 (O_1421,N_14167,N_13531);
or UO_1422 (O_1422,N_14089,N_14030);
or UO_1423 (O_1423,N_14892,N_14243);
and UO_1424 (O_1424,N_14871,N_14251);
and UO_1425 (O_1425,N_14593,N_13931);
or UO_1426 (O_1426,N_14696,N_14486);
nor UO_1427 (O_1427,N_14599,N_13857);
nor UO_1428 (O_1428,N_14745,N_13702);
nor UO_1429 (O_1429,N_13806,N_14817);
nand UO_1430 (O_1430,N_14526,N_14787);
nand UO_1431 (O_1431,N_13925,N_14059);
nor UO_1432 (O_1432,N_14295,N_13569);
nor UO_1433 (O_1433,N_14173,N_14112);
and UO_1434 (O_1434,N_13964,N_13962);
and UO_1435 (O_1435,N_14532,N_14977);
nand UO_1436 (O_1436,N_14083,N_14832);
or UO_1437 (O_1437,N_14768,N_14387);
nand UO_1438 (O_1438,N_14650,N_14654);
nand UO_1439 (O_1439,N_14488,N_14327);
and UO_1440 (O_1440,N_13809,N_14140);
or UO_1441 (O_1441,N_14728,N_14441);
nand UO_1442 (O_1442,N_14820,N_14011);
and UO_1443 (O_1443,N_14147,N_13682);
or UO_1444 (O_1444,N_13653,N_14726);
nor UO_1445 (O_1445,N_14015,N_13846);
nor UO_1446 (O_1446,N_13652,N_14080);
nor UO_1447 (O_1447,N_13692,N_14570);
and UO_1448 (O_1448,N_14927,N_13766);
nand UO_1449 (O_1449,N_14050,N_14462);
nor UO_1450 (O_1450,N_13717,N_13849);
or UO_1451 (O_1451,N_14826,N_14743);
nor UO_1452 (O_1452,N_14120,N_13927);
nor UO_1453 (O_1453,N_14918,N_13586);
nor UO_1454 (O_1454,N_14168,N_13625);
nor UO_1455 (O_1455,N_14497,N_14956);
and UO_1456 (O_1456,N_13911,N_14594);
nor UO_1457 (O_1457,N_13603,N_14077);
nor UO_1458 (O_1458,N_13938,N_14235);
and UO_1459 (O_1459,N_14532,N_14720);
and UO_1460 (O_1460,N_14967,N_14537);
or UO_1461 (O_1461,N_13611,N_14748);
or UO_1462 (O_1462,N_14189,N_14500);
or UO_1463 (O_1463,N_14885,N_14319);
or UO_1464 (O_1464,N_14868,N_14285);
and UO_1465 (O_1465,N_13635,N_14201);
or UO_1466 (O_1466,N_14684,N_14447);
nor UO_1467 (O_1467,N_13949,N_14297);
nand UO_1468 (O_1468,N_13962,N_13882);
nand UO_1469 (O_1469,N_13955,N_13502);
or UO_1470 (O_1470,N_13923,N_14452);
and UO_1471 (O_1471,N_14522,N_14640);
nand UO_1472 (O_1472,N_14660,N_14220);
nor UO_1473 (O_1473,N_14723,N_14209);
or UO_1474 (O_1474,N_14737,N_14920);
nor UO_1475 (O_1475,N_14663,N_14089);
or UO_1476 (O_1476,N_14143,N_14191);
or UO_1477 (O_1477,N_14241,N_14573);
and UO_1478 (O_1478,N_14697,N_14778);
nand UO_1479 (O_1479,N_14944,N_14035);
nand UO_1480 (O_1480,N_13726,N_14766);
nand UO_1481 (O_1481,N_13659,N_14449);
xor UO_1482 (O_1482,N_14116,N_14213);
and UO_1483 (O_1483,N_14158,N_13805);
nand UO_1484 (O_1484,N_14947,N_14338);
nand UO_1485 (O_1485,N_14275,N_13784);
nand UO_1486 (O_1486,N_13913,N_13783);
or UO_1487 (O_1487,N_14739,N_14550);
nand UO_1488 (O_1488,N_13625,N_14586);
or UO_1489 (O_1489,N_13505,N_13691);
and UO_1490 (O_1490,N_14969,N_14598);
nor UO_1491 (O_1491,N_14443,N_14248);
nor UO_1492 (O_1492,N_14126,N_14667);
and UO_1493 (O_1493,N_13940,N_14245);
nor UO_1494 (O_1494,N_14264,N_13997);
and UO_1495 (O_1495,N_14908,N_14103);
or UO_1496 (O_1496,N_13711,N_13945);
and UO_1497 (O_1497,N_14025,N_14900);
nor UO_1498 (O_1498,N_13861,N_14438);
nand UO_1499 (O_1499,N_13653,N_13784);
nor UO_1500 (O_1500,N_14652,N_14958);
or UO_1501 (O_1501,N_14085,N_14729);
and UO_1502 (O_1502,N_14892,N_14927);
and UO_1503 (O_1503,N_14453,N_14164);
and UO_1504 (O_1504,N_14282,N_14843);
nor UO_1505 (O_1505,N_13575,N_14490);
nand UO_1506 (O_1506,N_14729,N_13550);
nor UO_1507 (O_1507,N_14101,N_14715);
and UO_1508 (O_1508,N_14388,N_13671);
nor UO_1509 (O_1509,N_14046,N_13683);
nor UO_1510 (O_1510,N_13620,N_14403);
and UO_1511 (O_1511,N_13646,N_14518);
nor UO_1512 (O_1512,N_13754,N_14315);
nand UO_1513 (O_1513,N_13772,N_14211);
nand UO_1514 (O_1514,N_14281,N_14970);
and UO_1515 (O_1515,N_14770,N_14061);
or UO_1516 (O_1516,N_14529,N_13834);
and UO_1517 (O_1517,N_14468,N_14520);
nand UO_1518 (O_1518,N_13769,N_13717);
nand UO_1519 (O_1519,N_13844,N_13546);
nor UO_1520 (O_1520,N_14290,N_13865);
or UO_1521 (O_1521,N_14461,N_14486);
or UO_1522 (O_1522,N_13614,N_14930);
nand UO_1523 (O_1523,N_13633,N_14878);
nor UO_1524 (O_1524,N_14571,N_13643);
nor UO_1525 (O_1525,N_14287,N_13956);
nor UO_1526 (O_1526,N_14216,N_13787);
or UO_1527 (O_1527,N_13813,N_14620);
nor UO_1528 (O_1528,N_13824,N_14429);
and UO_1529 (O_1529,N_14541,N_14881);
or UO_1530 (O_1530,N_13869,N_14473);
or UO_1531 (O_1531,N_13635,N_13932);
or UO_1532 (O_1532,N_14785,N_13760);
nor UO_1533 (O_1533,N_14554,N_13781);
nand UO_1534 (O_1534,N_13961,N_14989);
nand UO_1535 (O_1535,N_14769,N_13867);
and UO_1536 (O_1536,N_14454,N_13930);
and UO_1537 (O_1537,N_14262,N_14167);
nand UO_1538 (O_1538,N_13794,N_13837);
and UO_1539 (O_1539,N_14585,N_14391);
or UO_1540 (O_1540,N_13748,N_14435);
and UO_1541 (O_1541,N_14108,N_14622);
nor UO_1542 (O_1542,N_14725,N_13642);
nand UO_1543 (O_1543,N_14189,N_13825);
nand UO_1544 (O_1544,N_14942,N_13651);
and UO_1545 (O_1545,N_13959,N_14892);
or UO_1546 (O_1546,N_14397,N_14968);
nand UO_1547 (O_1547,N_14933,N_13500);
or UO_1548 (O_1548,N_14099,N_14498);
and UO_1549 (O_1549,N_14777,N_13659);
or UO_1550 (O_1550,N_14917,N_13851);
nor UO_1551 (O_1551,N_13644,N_14339);
and UO_1552 (O_1552,N_13784,N_14821);
or UO_1553 (O_1553,N_14612,N_14138);
and UO_1554 (O_1554,N_14858,N_14828);
and UO_1555 (O_1555,N_13639,N_13790);
nand UO_1556 (O_1556,N_14243,N_14089);
nor UO_1557 (O_1557,N_14667,N_14393);
nor UO_1558 (O_1558,N_14167,N_13978);
nand UO_1559 (O_1559,N_14161,N_14302);
nor UO_1560 (O_1560,N_13576,N_14554);
nor UO_1561 (O_1561,N_14300,N_14771);
nor UO_1562 (O_1562,N_14748,N_14345);
nand UO_1563 (O_1563,N_13989,N_14522);
or UO_1564 (O_1564,N_13905,N_14225);
or UO_1565 (O_1565,N_13505,N_13608);
or UO_1566 (O_1566,N_13637,N_14930);
or UO_1567 (O_1567,N_13824,N_14723);
and UO_1568 (O_1568,N_14129,N_14408);
and UO_1569 (O_1569,N_14092,N_14109);
nand UO_1570 (O_1570,N_14396,N_14912);
xor UO_1571 (O_1571,N_14767,N_14034);
nand UO_1572 (O_1572,N_13706,N_13991);
and UO_1573 (O_1573,N_13869,N_13953);
nand UO_1574 (O_1574,N_13817,N_14259);
nor UO_1575 (O_1575,N_14483,N_14620);
or UO_1576 (O_1576,N_14143,N_14178);
nor UO_1577 (O_1577,N_14718,N_13856);
nor UO_1578 (O_1578,N_13946,N_13995);
and UO_1579 (O_1579,N_13758,N_14302);
and UO_1580 (O_1580,N_13821,N_14458);
nand UO_1581 (O_1581,N_13826,N_13916);
and UO_1582 (O_1582,N_14492,N_14858);
nand UO_1583 (O_1583,N_14086,N_14962);
nor UO_1584 (O_1584,N_13959,N_14889);
and UO_1585 (O_1585,N_13599,N_14956);
nor UO_1586 (O_1586,N_14812,N_14351);
or UO_1587 (O_1587,N_13530,N_14759);
or UO_1588 (O_1588,N_14372,N_14048);
nand UO_1589 (O_1589,N_13956,N_14456);
and UO_1590 (O_1590,N_14726,N_13552);
and UO_1591 (O_1591,N_13563,N_13533);
nand UO_1592 (O_1592,N_14898,N_14049);
or UO_1593 (O_1593,N_14181,N_14724);
or UO_1594 (O_1594,N_13581,N_13750);
and UO_1595 (O_1595,N_13870,N_14093);
nor UO_1596 (O_1596,N_14767,N_14755);
and UO_1597 (O_1597,N_13843,N_14354);
nor UO_1598 (O_1598,N_14307,N_14245);
nor UO_1599 (O_1599,N_14029,N_14415);
or UO_1600 (O_1600,N_14226,N_14223);
nor UO_1601 (O_1601,N_13600,N_14786);
and UO_1602 (O_1602,N_14745,N_14649);
or UO_1603 (O_1603,N_14639,N_14544);
and UO_1604 (O_1604,N_14188,N_13908);
or UO_1605 (O_1605,N_14353,N_14633);
and UO_1606 (O_1606,N_14879,N_13649);
nor UO_1607 (O_1607,N_14114,N_14749);
nor UO_1608 (O_1608,N_13546,N_14114);
nand UO_1609 (O_1609,N_13881,N_13686);
nor UO_1610 (O_1610,N_13742,N_13530);
xor UO_1611 (O_1611,N_13603,N_13652);
nor UO_1612 (O_1612,N_13546,N_14555);
nor UO_1613 (O_1613,N_13962,N_14402);
and UO_1614 (O_1614,N_14806,N_13543);
and UO_1615 (O_1615,N_13883,N_14148);
nand UO_1616 (O_1616,N_14141,N_14913);
or UO_1617 (O_1617,N_14302,N_14591);
nor UO_1618 (O_1618,N_13807,N_14481);
or UO_1619 (O_1619,N_13785,N_14452);
nor UO_1620 (O_1620,N_14827,N_13623);
and UO_1621 (O_1621,N_14153,N_14471);
or UO_1622 (O_1622,N_13669,N_13775);
and UO_1623 (O_1623,N_14588,N_13726);
nand UO_1624 (O_1624,N_13761,N_14506);
or UO_1625 (O_1625,N_14051,N_14633);
nor UO_1626 (O_1626,N_14184,N_14863);
and UO_1627 (O_1627,N_14167,N_14231);
nor UO_1628 (O_1628,N_14021,N_14861);
and UO_1629 (O_1629,N_13931,N_14329);
or UO_1630 (O_1630,N_14416,N_14038);
nor UO_1631 (O_1631,N_14154,N_14682);
or UO_1632 (O_1632,N_14927,N_14962);
nand UO_1633 (O_1633,N_13521,N_14029);
nand UO_1634 (O_1634,N_14280,N_14066);
nor UO_1635 (O_1635,N_14797,N_14040);
or UO_1636 (O_1636,N_14291,N_13502);
nor UO_1637 (O_1637,N_14204,N_14232);
nand UO_1638 (O_1638,N_14685,N_14309);
xnor UO_1639 (O_1639,N_14811,N_14114);
nor UO_1640 (O_1640,N_13831,N_14946);
and UO_1641 (O_1641,N_14506,N_14556);
and UO_1642 (O_1642,N_13948,N_13662);
or UO_1643 (O_1643,N_14805,N_13990);
nand UO_1644 (O_1644,N_14397,N_14062);
nand UO_1645 (O_1645,N_13703,N_13521);
and UO_1646 (O_1646,N_13574,N_14672);
nand UO_1647 (O_1647,N_14532,N_13794);
nand UO_1648 (O_1648,N_14190,N_14720);
nand UO_1649 (O_1649,N_13951,N_13880);
nor UO_1650 (O_1650,N_14617,N_14867);
and UO_1651 (O_1651,N_14847,N_14739);
and UO_1652 (O_1652,N_14012,N_14946);
nor UO_1653 (O_1653,N_14488,N_14104);
or UO_1654 (O_1654,N_14047,N_14394);
or UO_1655 (O_1655,N_14243,N_13917);
and UO_1656 (O_1656,N_14703,N_14864);
nand UO_1657 (O_1657,N_14700,N_13706);
nand UO_1658 (O_1658,N_14829,N_13720);
nand UO_1659 (O_1659,N_14218,N_14910);
or UO_1660 (O_1660,N_14226,N_14575);
nor UO_1661 (O_1661,N_14700,N_14290);
nor UO_1662 (O_1662,N_13591,N_13554);
or UO_1663 (O_1663,N_14990,N_14919);
and UO_1664 (O_1664,N_14112,N_14426);
nand UO_1665 (O_1665,N_14160,N_14487);
nor UO_1666 (O_1666,N_13709,N_14854);
xnor UO_1667 (O_1667,N_14760,N_14482);
and UO_1668 (O_1668,N_13625,N_13523);
or UO_1669 (O_1669,N_14191,N_13919);
and UO_1670 (O_1670,N_14252,N_13776);
and UO_1671 (O_1671,N_14756,N_14210);
nand UO_1672 (O_1672,N_14688,N_14182);
nand UO_1673 (O_1673,N_14359,N_14677);
nor UO_1674 (O_1674,N_14005,N_14689);
nor UO_1675 (O_1675,N_13824,N_13964);
and UO_1676 (O_1676,N_14267,N_13530);
nand UO_1677 (O_1677,N_14992,N_13935);
and UO_1678 (O_1678,N_14731,N_13976);
nor UO_1679 (O_1679,N_13979,N_14679);
nor UO_1680 (O_1680,N_14506,N_13723);
nor UO_1681 (O_1681,N_14203,N_13754);
nand UO_1682 (O_1682,N_14138,N_13863);
and UO_1683 (O_1683,N_14590,N_13632);
or UO_1684 (O_1684,N_14644,N_13839);
or UO_1685 (O_1685,N_14041,N_14239);
or UO_1686 (O_1686,N_14932,N_14219);
and UO_1687 (O_1687,N_13664,N_13804);
and UO_1688 (O_1688,N_14351,N_14779);
nand UO_1689 (O_1689,N_14148,N_13602);
and UO_1690 (O_1690,N_13735,N_14592);
or UO_1691 (O_1691,N_13819,N_13797);
nor UO_1692 (O_1692,N_14117,N_14825);
or UO_1693 (O_1693,N_13963,N_14536);
nor UO_1694 (O_1694,N_14209,N_14394);
nand UO_1695 (O_1695,N_14570,N_14519);
or UO_1696 (O_1696,N_14583,N_14781);
and UO_1697 (O_1697,N_14223,N_14098);
and UO_1698 (O_1698,N_14375,N_13913);
nor UO_1699 (O_1699,N_13857,N_13893);
or UO_1700 (O_1700,N_14077,N_14397);
and UO_1701 (O_1701,N_14563,N_14528);
nor UO_1702 (O_1702,N_14297,N_14266);
and UO_1703 (O_1703,N_13884,N_13526);
or UO_1704 (O_1704,N_14621,N_13684);
or UO_1705 (O_1705,N_14529,N_13569);
and UO_1706 (O_1706,N_13947,N_14755);
xnor UO_1707 (O_1707,N_14607,N_14170);
or UO_1708 (O_1708,N_14756,N_14944);
or UO_1709 (O_1709,N_14481,N_14022);
nand UO_1710 (O_1710,N_14932,N_13782);
or UO_1711 (O_1711,N_14051,N_14580);
nand UO_1712 (O_1712,N_14401,N_13868);
nand UO_1713 (O_1713,N_14532,N_14019);
nor UO_1714 (O_1714,N_13890,N_13569);
or UO_1715 (O_1715,N_13519,N_13622);
nand UO_1716 (O_1716,N_14291,N_14420);
nor UO_1717 (O_1717,N_13585,N_13736);
or UO_1718 (O_1718,N_14896,N_13650);
and UO_1719 (O_1719,N_14908,N_14217);
xnor UO_1720 (O_1720,N_13872,N_13622);
or UO_1721 (O_1721,N_14560,N_13947);
nor UO_1722 (O_1722,N_13969,N_14289);
or UO_1723 (O_1723,N_14428,N_14008);
or UO_1724 (O_1724,N_14493,N_13800);
nand UO_1725 (O_1725,N_14195,N_14231);
or UO_1726 (O_1726,N_14941,N_13840);
and UO_1727 (O_1727,N_13827,N_14303);
nor UO_1728 (O_1728,N_14982,N_14749);
nand UO_1729 (O_1729,N_14513,N_14657);
nand UO_1730 (O_1730,N_14805,N_13577);
or UO_1731 (O_1731,N_14174,N_14680);
or UO_1732 (O_1732,N_14837,N_14230);
nand UO_1733 (O_1733,N_14117,N_14903);
nor UO_1734 (O_1734,N_14308,N_14883);
or UO_1735 (O_1735,N_14759,N_14293);
nor UO_1736 (O_1736,N_14840,N_14190);
and UO_1737 (O_1737,N_14142,N_14506);
nand UO_1738 (O_1738,N_14777,N_14136);
nand UO_1739 (O_1739,N_14437,N_13999);
nor UO_1740 (O_1740,N_14986,N_13550);
nor UO_1741 (O_1741,N_14789,N_14313);
nand UO_1742 (O_1742,N_14157,N_13967);
and UO_1743 (O_1743,N_14897,N_14446);
and UO_1744 (O_1744,N_14057,N_14925);
or UO_1745 (O_1745,N_13775,N_14373);
and UO_1746 (O_1746,N_14651,N_14237);
and UO_1747 (O_1747,N_13910,N_13760);
and UO_1748 (O_1748,N_13762,N_13927);
and UO_1749 (O_1749,N_13673,N_13956);
and UO_1750 (O_1750,N_14065,N_14941);
nand UO_1751 (O_1751,N_14112,N_13978);
nor UO_1752 (O_1752,N_14178,N_14476);
or UO_1753 (O_1753,N_14470,N_13563);
and UO_1754 (O_1754,N_14708,N_13789);
and UO_1755 (O_1755,N_14723,N_14294);
nand UO_1756 (O_1756,N_14662,N_14638);
nor UO_1757 (O_1757,N_14350,N_14378);
nand UO_1758 (O_1758,N_14982,N_14430);
nor UO_1759 (O_1759,N_14108,N_14058);
or UO_1760 (O_1760,N_13799,N_13614);
and UO_1761 (O_1761,N_14871,N_13533);
or UO_1762 (O_1762,N_14653,N_14290);
nand UO_1763 (O_1763,N_13835,N_14296);
xnor UO_1764 (O_1764,N_14575,N_14419);
or UO_1765 (O_1765,N_13573,N_14284);
nand UO_1766 (O_1766,N_14527,N_14646);
nand UO_1767 (O_1767,N_13994,N_13503);
and UO_1768 (O_1768,N_14580,N_14892);
or UO_1769 (O_1769,N_13508,N_14373);
nor UO_1770 (O_1770,N_13633,N_14833);
nand UO_1771 (O_1771,N_13614,N_13845);
or UO_1772 (O_1772,N_14066,N_14114);
or UO_1773 (O_1773,N_14663,N_14194);
nand UO_1774 (O_1774,N_14842,N_13672);
and UO_1775 (O_1775,N_14910,N_13984);
nand UO_1776 (O_1776,N_14501,N_14174);
and UO_1777 (O_1777,N_14830,N_13636);
or UO_1778 (O_1778,N_14127,N_13564);
nor UO_1779 (O_1779,N_14752,N_13623);
nor UO_1780 (O_1780,N_14563,N_14409);
nand UO_1781 (O_1781,N_14956,N_14968);
nand UO_1782 (O_1782,N_14184,N_14214);
nand UO_1783 (O_1783,N_14407,N_13504);
or UO_1784 (O_1784,N_14392,N_14531);
and UO_1785 (O_1785,N_14651,N_14974);
and UO_1786 (O_1786,N_14744,N_14741);
nor UO_1787 (O_1787,N_14584,N_14486);
and UO_1788 (O_1788,N_14382,N_13932);
nand UO_1789 (O_1789,N_14004,N_14835);
nand UO_1790 (O_1790,N_14947,N_14098);
nand UO_1791 (O_1791,N_13897,N_13520);
and UO_1792 (O_1792,N_13860,N_13913);
nand UO_1793 (O_1793,N_13619,N_13535);
or UO_1794 (O_1794,N_13752,N_13821);
and UO_1795 (O_1795,N_14687,N_14442);
and UO_1796 (O_1796,N_13608,N_14951);
nor UO_1797 (O_1797,N_14382,N_14290);
and UO_1798 (O_1798,N_14669,N_13813);
and UO_1799 (O_1799,N_14856,N_14235);
and UO_1800 (O_1800,N_13662,N_13588);
and UO_1801 (O_1801,N_14611,N_14708);
nor UO_1802 (O_1802,N_14915,N_13843);
nor UO_1803 (O_1803,N_13779,N_14752);
nand UO_1804 (O_1804,N_14618,N_14841);
or UO_1805 (O_1805,N_13991,N_14272);
and UO_1806 (O_1806,N_13656,N_13511);
nand UO_1807 (O_1807,N_14086,N_13507);
nor UO_1808 (O_1808,N_14942,N_14687);
nand UO_1809 (O_1809,N_13931,N_13821);
nor UO_1810 (O_1810,N_13765,N_14125);
and UO_1811 (O_1811,N_14494,N_14966);
nor UO_1812 (O_1812,N_14016,N_13746);
nand UO_1813 (O_1813,N_13856,N_14301);
and UO_1814 (O_1814,N_14078,N_14709);
nor UO_1815 (O_1815,N_14161,N_14889);
nor UO_1816 (O_1816,N_14433,N_13751);
or UO_1817 (O_1817,N_14856,N_14630);
nor UO_1818 (O_1818,N_14108,N_14358);
or UO_1819 (O_1819,N_14183,N_13741);
nor UO_1820 (O_1820,N_14859,N_14521);
nor UO_1821 (O_1821,N_14395,N_14415);
nor UO_1822 (O_1822,N_13952,N_13745);
or UO_1823 (O_1823,N_14411,N_13899);
or UO_1824 (O_1824,N_14641,N_14130);
nor UO_1825 (O_1825,N_14133,N_14209);
or UO_1826 (O_1826,N_13883,N_14367);
nor UO_1827 (O_1827,N_14885,N_14127);
nand UO_1828 (O_1828,N_13644,N_14654);
nand UO_1829 (O_1829,N_13973,N_13843);
and UO_1830 (O_1830,N_13662,N_14746);
and UO_1831 (O_1831,N_14953,N_14705);
and UO_1832 (O_1832,N_14983,N_14220);
nor UO_1833 (O_1833,N_14090,N_14456);
or UO_1834 (O_1834,N_14338,N_14084);
nor UO_1835 (O_1835,N_14795,N_13541);
and UO_1836 (O_1836,N_14581,N_14649);
nor UO_1837 (O_1837,N_13651,N_14377);
nor UO_1838 (O_1838,N_14413,N_14443);
and UO_1839 (O_1839,N_13555,N_14049);
nand UO_1840 (O_1840,N_14144,N_14956);
or UO_1841 (O_1841,N_14282,N_13763);
or UO_1842 (O_1842,N_13715,N_13834);
or UO_1843 (O_1843,N_14238,N_14784);
and UO_1844 (O_1844,N_14620,N_14043);
nand UO_1845 (O_1845,N_14108,N_14005);
and UO_1846 (O_1846,N_13815,N_13708);
and UO_1847 (O_1847,N_14827,N_14384);
nand UO_1848 (O_1848,N_14737,N_14488);
or UO_1849 (O_1849,N_14869,N_13679);
or UO_1850 (O_1850,N_14109,N_13790);
nor UO_1851 (O_1851,N_13830,N_13781);
and UO_1852 (O_1852,N_14204,N_14366);
or UO_1853 (O_1853,N_13854,N_13820);
and UO_1854 (O_1854,N_13697,N_13508);
and UO_1855 (O_1855,N_14339,N_13764);
and UO_1856 (O_1856,N_13551,N_13763);
or UO_1857 (O_1857,N_14407,N_13938);
or UO_1858 (O_1858,N_14553,N_13637);
nor UO_1859 (O_1859,N_13686,N_14577);
nor UO_1860 (O_1860,N_14052,N_13539);
nand UO_1861 (O_1861,N_13833,N_14639);
nor UO_1862 (O_1862,N_13721,N_14748);
and UO_1863 (O_1863,N_14084,N_13794);
nor UO_1864 (O_1864,N_14857,N_14820);
nor UO_1865 (O_1865,N_13955,N_13908);
nand UO_1866 (O_1866,N_14707,N_13511);
or UO_1867 (O_1867,N_13806,N_14174);
and UO_1868 (O_1868,N_14960,N_13638);
and UO_1869 (O_1869,N_14357,N_14552);
nand UO_1870 (O_1870,N_14116,N_14473);
nand UO_1871 (O_1871,N_13881,N_14304);
nand UO_1872 (O_1872,N_14021,N_13833);
and UO_1873 (O_1873,N_14943,N_14372);
nor UO_1874 (O_1874,N_13547,N_14929);
nand UO_1875 (O_1875,N_13991,N_14376);
or UO_1876 (O_1876,N_14783,N_14857);
and UO_1877 (O_1877,N_14014,N_14240);
nand UO_1878 (O_1878,N_14644,N_14328);
nand UO_1879 (O_1879,N_13745,N_14952);
and UO_1880 (O_1880,N_13656,N_14907);
nand UO_1881 (O_1881,N_13892,N_14111);
nand UO_1882 (O_1882,N_14204,N_14465);
and UO_1883 (O_1883,N_14113,N_14864);
nor UO_1884 (O_1884,N_14982,N_13604);
nor UO_1885 (O_1885,N_14616,N_13529);
nor UO_1886 (O_1886,N_13522,N_14573);
or UO_1887 (O_1887,N_14423,N_13623);
nand UO_1888 (O_1888,N_14533,N_14304);
and UO_1889 (O_1889,N_14662,N_14935);
and UO_1890 (O_1890,N_14984,N_14668);
nor UO_1891 (O_1891,N_14056,N_14054);
or UO_1892 (O_1892,N_14712,N_14448);
nor UO_1893 (O_1893,N_13726,N_13868);
nand UO_1894 (O_1894,N_13805,N_13694);
nor UO_1895 (O_1895,N_13925,N_14616);
and UO_1896 (O_1896,N_13555,N_14721);
or UO_1897 (O_1897,N_14944,N_13692);
nor UO_1898 (O_1898,N_13669,N_14052);
or UO_1899 (O_1899,N_14289,N_13550);
and UO_1900 (O_1900,N_14471,N_14023);
or UO_1901 (O_1901,N_13933,N_14156);
nor UO_1902 (O_1902,N_13823,N_14116);
nand UO_1903 (O_1903,N_13863,N_13663);
or UO_1904 (O_1904,N_14508,N_13970);
nor UO_1905 (O_1905,N_14109,N_13581);
or UO_1906 (O_1906,N_14590,N_13934);
nor UO_1907 (O_1907,N_14054,N_14580);
and UO_1908 (O_1908,N_14314,N_14013);
or UO_1909 (O_1909,N_14738,N_14277);
nand UO_1910 (O_1910,N_13517,N_14411);
nor UO_1911 (O_1911,N_14475,N_14907);
nand UO_1912 (O_1912,N_13564,N_13863);
nand UO_1913 (O_1913,N_13530,N_14337);
or UO_1914 (O_1914,N_14907,N_14893);
nor UO_1915 (O_1915,N_13707,N_14527);
nand UO_1916 (O_1916,N_14054,N_14215);
and UO_1917 (O_1917,N_13635,N_14368);
nor UO_1918 (O_1918,N_14406,N_13849);
or UO_1919 (O_1919,N_13551,N_14622);
and UO_1920 (O_1920,N_14291,N_14040);
or UO_1921 (O_1921,N_14830,N_13608);
nor UO_1922 (O_1922,N_14864,N_14674);
and UO_1923 (O_1923,N_14008,N_13567);
and UO_1924 (O_1924,N_13576,N_14385);
or UO_1925 (O_1925,N_14773,N_13730);
nor UO_1926 (O_1926,N_14891,N_13749);
and UO_1927 (O_1927,N_14761,N_14820);
nor UO_1928 (O_1928,N_13811,N_14136);
nand UO_1929 (O_1929,N_14332,N_14980);
or UO_1930 (O_1930,N_14040,N_14118);
xnor UO_1931 (O_1931,N_13928,N_13876);
nand UO_1932 (O_1932,N_14956,N_13932);
and UO_1933 (O_1933,N_13559,N_14910);
or UO_1934 (O_1934,N_13889,N_13595);
or UO_1935 (O_1935,N_13950,N_14071);
nand UO_1936 (O_1936,N_14187,N_14616);
nand UO_1937 (O_1937,N_13905,N_14527);
or UO_1938 (O_1938,N_14651,N_14191);
xnor UO_1939 (O_1939,N_14076,N_13852);
and UO_1940 (O_1940,N_14173,N_14837);
and UO_1941 (O_1941,N_13504,N_14971);
and UO_1942 (O_1942,N_13984,N_14422);
or UO_1943 (O_1943,N_14065,N_14954);
and UO_1944 (O_1944,N_14171,N_14169);
nand UO_1945 (O_1945,N_13747,N_14293);
or UO_1946 (O_1946,N_14045,N_13646);
nand UO_1947 (O_1947,N_14339,N_13804);
nand UO_1948 (O_1948,N_14721,N_14068);
and UO_1949 (O_1949,N_14782,N_14857);
nor UO_1950 (O_1950,N_14997,N_14239);
and UO_1951 (O_1951,N_14730,N_14110);
and UO_1952 (O_1952,N_14117,N_14271);
xnor UO_1953 (O_1953,N_13512,N_14909);
and UO_1954 (O_1954,N_14774,N_14746);
nand UO_1955 (O_1955,N_14580,N_14120);
or UO_1956 (O_1956,N_14543,N_14848);
nand UO_1957 (O_1957,N_14700,N_14721);
nand UO_1958 (O_1958,N_14989,N_13700);
nand UO_1959 (O_1959,N_14463,N_14057);
nand UO_1960 (O_1960,N_14902,N_14585);
and UO_1961 (O_1961,N_14716,N_14569);
or UO_1962 (O_1962,N_14253,N_14811);
nand UO_1963 (O_1963,N_14418,N_13713);
or UO_1964 (O_1964,N_13888,N_14062);
xor UO_1965 (O_1965,N_14673,N_14286);
nand UO_1966 (O_1966,N_14909,N_13586);
nand UO_1967 (O_1967,N_14788,N_13982);
nand UO_1968 (O_1968,N_13903,N_14182);
nor UO_1969 (O_1969,N_13749,N_13562);
or UO_1970 (O_1970,N_14402,N_13910);
nor UO_1971 (O_1971,N_14743,N_14389);
nand UO_1972 (O_1972,N_14789,N_13946);
and UO_1973 (O_1973,N_13846,N_14936);
nor UO_1974 (O_1974,N_13538,N_14842);
or UO_1975 (O_1975,N_14455,N_14961);
nor UO_1976 (O_1976,N_14400,N_14049);
nor UO_1977 (O_1977,N_14324,N_14767);
and UO_1978 (O_1978,N_14186,N_14809);
nand UO_1979 (O_1979,N_13613,N_13709);
nand UO_1980 (O_1980,N_14104,N_14609);
nor UO_1981 (O_1981,N_14294,N_14913);
or UO_1982 (O_1982,N_14436,N_14624);
or UO_1983 (O_1983,N_14738,N_13779);
and UO_1984 (O_1984,N_14231,N_14642);
and UO_1985 (O_1985,N_14274,N_13661);
or UO_1986 (O_1986,N_14741,N_14123);
or UO_1987 (O_1987,N_13798,N_14223);
nand UO_1988 (O_1988,N_13856,N_14650);
nor UO_1989 (O_1989,N_14669,N_14784);
and UO_1990 (O_1990,N_14259,N_14094);
and UO_1991 (O_1991,N_13549,N_14496);
nand UO_1992 (O_1992,N_14281,N_13699);
nand UO_1993 (O_1993,N_14436,N_14487);
and UO_1994 (O_1994,N_14460,N_13970);
nor UO_1995 (O_1995,N_13872,N_13955);
or UO_1996 (O_1996,N_13621,N_14460);
nand UO_1997 (O_1997,N_14834,N_13965);
nand UO_1998 (O_1998,N_13864,N_14544);
or UO_1999 (O_1999,N_13876,N_13622);
endmodule