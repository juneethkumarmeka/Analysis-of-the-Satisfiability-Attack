module basic_750_5000_1000_25_levels_2xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
nand U0 (N_0,In_128,In_687);
or U1 (N_1,In_417,In_173);
nor U2 (N_2,In_555,In_0);
and U3 (N_3,In_342,In_537);
nor U4 (N_4,In_209,In_386);
or U5 (N_5,In_730,In_235);
nor U6 (N_6,In_266,In_189);
or U7 (N_7,In_253,In_36);
nand U8 (N_8,In_264,In_135);
and U9 (N_9,In_679,In_638);
nor U10 (N_10,In_736,In_32);
and U11 (N_11,In_713,In_343);
nor U12 (N_12,In_81,In_338);
or U13 (N_13,In_605,In_484);
nand U14 (N_14,In_291,In_402);
nand U15 (N_15,In_457,In_734);
or U16 (N_16,In_357,In_503);
nor U17 (N_17,In_702,In_241);
nor U18 (N_18,In_579,In_504);
nor U19 (N_19,In_126,In_482);
or U20 (N_20,In_118,In_589);
nand U21 (N_21,In_155,In_377);
nor U22 (N_22,In_448,In_424);
and U23 (N_23,In_90,In_304);
or U24 (N_24,In_184,In_525);
nand U25 (N_25,In_57,In_334);
or U26 (N_26,In_230,In_522);
nand U27 (N_27,In_204,In_636);
nand U28 (N_28,In_65,In_33);
and U29 (N_29,In_540,In_285);
xor U30 (N_30,In_728,In_551);
xnor U31 (N_31,In_621,In_177);
nand U32 (N_32,In_320,In_564);
nand U33 (N_33,In_236,In_528);
nor U34 (N_34,In_481,In_314);
nand U35 (N_35,In_444,In_646);
nor U36 (N_36,In_624,In_14);
nand U37 (N_37,In_244,In_558);
and U38 (N_38,In_627,In_170);
nand U39 (N_39,In_460,In_632);
or U40 (N_40,In_573,In_480);
nand U41 (N_41,In_127,In_399);
nand U42 (N_42,In_634,In_328);
nand U43 (N_43,In_310,In_592);
nand U44 (N_44,In_13,In_221);
and U45 (N_45,In_473,In_447);
or U46 (N_46,In_688,In_131);
nand U47 (N_47,In_628,In_231);
and U48 (N_48,In_239,In_167);
nor U49 (N_49,In_296,In_647);
and U50 (N_50,In_681,In_576);
nand U51 (N_51,In_607,In_745);
nor U52 (N_52,In_722,In_563);
and U53 (N_53,In_349,In_711);
nor U54 (N_54,In_600,In_159);
nand U55 (N_55,In_415,In_698);
or U56 (N_56,In_570,In_298);
or U57 (N_57,In_387,In_526);
and U58 (N_58,In_88,In_651);
or U59 (N_59,In_3,In_265);
nor U60 (N_60,In_141,In_657);
nand U61 (N_61,In_4,In_259);
and U62 (N_62,In_217,In_436);
nor U63 (N_63,In_86,In_39);
xnor U64 (N_64,In_613,In_534);
xor U65 (N_65,In_198,In_140);
xnor U66 (N_66,In_455,In_717);
and U67 (N_67,In_527,In_445);
nor U68 (N_68,In_375,In_658);
nor U69 (N_69,In_201,In_323);
or U70 (N_70,In_418,In_603);
nor U71 (N_71,In_523,In_749);
nand U72 (N_72,In_403,In_517);
nand U73 (N_73,In_674,In_79);
or U74 (N_74,In_676,In_544);
nand U75 (N_75,In_222,In_58);
nor U76 (N_76,In_468,In_142);
nand U77 (N_77,In_149,In_132);
and U78 (N_78,In_109,In_125);
nand U79 (N_79,In_391,In_166);
nor U80 (N_80,In_359,In_505);
nor U81 (N_81,In_590,In_367);
nor U82 (N_82,In_156,In_656);
nor U83 (N_83,In_542,In_407);
and U84 (N_84,In_55,In_92);
and U85 (N_85,In_178,In_566);
nor U86 (N_86,In_684,In_620);
nor U87 (N_87,In_242,In_732);
or U88 (N_88,In_179,In_479);
or U89 (N_89,In_188,In_735);
nand U90 (N_90,In_390,In_196);
nor U91 (N_91,In_116,In_669);
and U92 (N_92,In_597,In_238);
nor U93 (N_93,In_234,In_440);
and U94 (N_94,In_616,In_219);
nor U95 (N_95,In_335,In_267);
nor U96 (N_96,In_382,In_274);
nor U97 (N_97,In_599,In_532);
or U98 (N_98,In_397,In_28);
nand U99 (N_99,In_565,In_587);
or U100 (N_100,In_560,In_153);
nand U101 (N_101,In_195,In_213);
nor U102 (N_102,In_164,In_695);
nand U103 (N_103,In_136,In_427);
and U104 (N_104,In_20,In_748);
or U105 (N_105,In_240,In_429);
and U106 (N_106,In_268,In_718);
or U107 (N_107,In_495,In_146);
nor U108 (N_108,In_705,In_277);
or U109 (N_109,In_258,In_451);
or U110 (N_110,In_594,In_609);
or U111 (N_111,In_10,In_630);
or U112 (N_112,In_8,In_344);
and U113 (N_113,In_223,In_53);
or U114 (N_114,In_106,In_514);
or U115 (N_115,In_215,In_644);
or U116 (N_116,In_461,In_625);
and U117 (N_117,In_2,In_207);
or U118 (N_118,In_324,In_261);
and U119 (N_119,In_193,In_413);
or U120 (N_120,In_553,In_17);
or U121 (N_121,In_64,In_59);
or U122 (N_122,In_355,In_746);
nor U123 (N_123,In_80,In_100);
nand U124 (N_124,In_224,In_708);
nor U125 (N_125,In_337,In_331);
nor U126 (N_126,In_313,In_409);
or U127 (N_127,In_21,In_162);
or U128 (N_128,In_103,In_442);
nand U129 (N_129,In_353,In_247);
nor U130 (N_130,In_61,In_76);
nand U131 (N_131,In_346,In_69);
and U132 (N_132,In_692,In_400);
and U133 (N_133,In_562,In_330);
nor U134 (N_134,In_124,In_245);
nor U135 (N_135,In_639,In_216);
and U136 (N_136,In_364,In_568);
or U137 (N_137,In_250,In_388);
or U138 (N_138,In_332,In_273);
and U139 (N_139,In_694,In_358);
and U140 (N_140,In_99,In_411);
nor U141 (N_141,In_666,In_428);
and U142 (N_142,In_114,In_721);
nand U143 (N_143,In_663,In_82);
nand U144 (N_144,In_425,In_742);
and U145 (N_145,In_452,In_303);
nand U146 (N_146,In_25,In_70);
or U147 (N_147,In_71,In_716);
xor U148 (N_148,In_383,In_501);
nor U149 (N_149,In_408,In_535);
and U150 (N_150,In_185,In_622);
or U151 (N_151,In_567,In_459);
or U152 (N_152,In_430,In_392);
or U153 (N_153,In_301,In_673);
nand U154 (N_154,In_472,In_180);
nand U155 (N_155,In_700,In_182);
and U156 (N_156,In_653,In_37);
and U157 (N_157,In_212,In_228);
nand U158 (N_158,In_263,In_302);
nor U159 (N_159,In_642,In_211);
nor U160 (N_160,In_699,In_243);
nor U161 (N_161,In_252,In_287);
nand U162 (N_162,In_168,In_214);
and U163 (N_163,In_706,In_601);
nand U164 (N_164,In_665,In_208);
nand U165 (N_165,In_414,In_516);
nor U166 (N_166,In_366,In_691);
or U167 (N_167,In_200,In_731);
nand U168 (N_168,In_161,In_279);
nand U169 (N_169,In_311,In_50);
nand U170 (N_170,In_499,In_197);
nor U171 (N_171,In_278,In_376);
nor U172 (N_172,In_175,In_134);
nor U173 (N_173,In_333,In_450);
or U174 (N_174,In_42,In_640);
or U175 (N_175,In_119,In_370);
nor U176 (N_176,In_496,In_95);
or U177 (N_177,In_519,In_297);
nor U178 (N_178,In_325,In_191);
or U179 (N_179,In_405,In_582);
nand U180 (N_180,In_633,In_435);
nor U181 (N_181,In_690,In_584);
nand U182 (N_182,In_7,In_1);
nor U183 (N_183,In_105,In_449);
nor U184 (N_184,In_580,In_678);
nor U185 (N_185,In_115,In_44);
or U186 (N_186,In_77,In_586);
nor U187 (N_187,In_741,In_282);
nor U188 (N_188,In_352,In_150);
or U189 (N_189,In_533,In_737);
or U190 (N_190,In_596,In_571);
nor U191 (N_191,In_111,In_422);
nand U192 (N_192,In_139,In_143);
nand U193 (N_193,In_321,In_183);
nor U194 (N_194,In_374,In_423);
nor U195 (N_195,In_255,In_262);
nor U196 (N_196,In_538,In_471);
or U197 (N_197,In_74,In_662);
and U198 (N_198,In_612,In_675);
nor U199 (N_199,In_347,In_606);
nand U200 (N_200,N_170,N_5);
and U201 (N_201,In_561,In_45);
xor U202 (N_202,N_85,In_194);
or U203 (N_203,In_689,In_454);
nor U204 (N_204,In_341,In_290);
and U205 (N_205,In_610,N_80);
nor U206 (N_206,N_40,In_110);
and U207 (N_207,In_23,In_133);
nand U208 (N_208,In_203,In_385);
nor U209 (N_209,In_598,In_29);
nor U210 (N_210,In_548,In_165);
nor U211 (N_211,In_510,In_434);
and U212 (N_212,In_617,In_248);
and U213 (N_213,N_69,N_67);
nand U214 (N_214,N_151,N_175);
xor U215 (N_215,N_88,In_744);
nor U216 (N_216,In_350,N_86);
and U217 (N_217,In_130,In_56);
or U218 (N_218,N_190,In_35);
nor U219 (N_219,In_643,In_372);
nand U220 (N_220,In_486,In_648);
nor U221 (N_221,In_93,N_46);
nand U222 (N_222,In_112,In_477);
nand U223 (N_223,In_664,In_365);
and U224 (N_224,In_467,In_724);
nand U225 (N_225,In_719,In_148);
nand U226 (N_226,In_233,In_438);
and U227 (N_227,In_465,In_659);
and U228 (N_228,In_257,N_16);
nand U229 (N_229,N_78,N_118);
and U230 (N_230,In_122,N_149);
nor U231 (N_231,N_177,In_368);
or U232 (N_232,In_498,N_96);
nor U233 (N_233,In_300,In_379);
nand U234 (N_234,In_163,In_701);
or U235 (N_235,In_476,In_431);
nor U236 (N_236,In_18,N_173);
or U237 (N_237,In_635,N_34);
nor U238 (N_238,N_17,In_319);
and U239 (N_239,In_577,In_229);
nor U240 (N_240,N_114,N_104);
nand U241 (N_241,N_4,N_108);
nand U242 (N_242,In_545,In_186);
nor U243 (N_243,In_40,In_11);
nand U244 (N_244,N_30,N_139);
nor U245 (N_245,In_453,In_595);
or U246 (N_246,In_104,In_412);
nand U247 (N_247,In_326,In_671);
and U248 (N_248,In_145,In_710);
and U249 (N_249,In_672,N_100);
and U250 (N_250,In_715,In_67);
nand U251 (N_251,In_157,N_122);
nand U252 (N_252,In_547,In_720);
and U253 (N_253,N_130,In_470);
and U254 (N_254,N_196,In_176);
xnor U255 (N_255,In_645,In_406);
or U256 (N_256,N_8,In_22);
nand U257 (N_257,N_11,N_60);
and U258 (N_258,N_43,In_41);
or U259 (N_259,In_611,In_318);
and U260 (N_260,In_462,In_312);
xor U261 (N_261,In_464,In_463);
nor U262 (N_262,In_16,In_500);
nand U263 (N_263,N_193,In_491);
and U264 (N_264,In_512,In_351);
nand U265 (N_265,N_141,In_206);
or U266 (N_266,In_541,In_62);
or U267 (N_267,In_593,N_155);
or U268 (N_268,In_360,In_747);
nand U269 (N_269,N_159,In_117);
and U270 (N_270,In_373,In_329);
or U271 (N_271,N_6,N_39);
nand U272 (N_272,In_509,In_295);
and U273 (N_273,In_98,In_288);
xor U274 (N_274,In_668,In_696);
nand U275 (N_275,In_660,N_101);
nor U276 (N_276,N_72,N_162);
xor U277 (N_277,In_475,N_158);
or U278 (N_278,In_72,N_110);
and U279 (N_279,In_623,N_195);
nor U280 (N_280,In_441,In_322);
nand U281 (N_281,In_123,In_437);
nor U282 (N_282,In_19,N_160);
and U283 (N_283,In_270,In_152);
or U284 (N_284,In_738,N_64);
and U285 (N_285,N_111,In_536);
nor U286 (N_286,In_220,In_726);
nor U287 (N_287,In_588,N_153);
nor U288 (N_288,In_380,In_91);
nand U289 (N_289,In_641,In_327);
nand U290 (N_290,In_218,In_138);
and U291 (N_291,In_280,In_256);
nand U292 (N_292,N_24,In_78);
nand U293 (N_293,In_539,In_269);
and U294 (N_294,In_410,In_107);
nand U295 (N_295,In_308,N_25);
or U296 (N_296,In_73,N_164);
nor U297 (N_297,In_232,N_48);
nand U298 (N_298,N_35,In_733);
and U299 (N_299,In_543,In_246);
or U300 (N_300,N_47,N_156);
or U301 (N_301,N_150,N_112);
and U302 (N_302,N_188,In_316);
and U303 (N_303,In_384,N_90);
nor U304 (N_304,In_446,N_1);
and U305 (N_305,N_65,In_650);
xnor U306 (N_306,N_103,N_81);
nand U307 (N_307,N_152,N_185);
or U308 (N_308,N_77,In_511);
and U309 (N_309,N_95,In_556);
nor U310 (N_310,In_96,N_157);
nor U311 (N_311,In_443,In_637);
and U312 (N_312,In_94,N_174);
and U313 (N_313,In_31,In_549);
or U314 (N_314,In_293,In_614);
and U315 (N_315,In_661,N_113);
nor U316 (N_316,In_552,In_707);
nand U317 (N_317,In_395,In_181);
nand U318 (N_318,In_550,N_136);
nand U319 (N_319,In_608,In_557);
nand U320 (N_320,N_76,In_469);
and U321 (N_321,In_354,In_369);
and U322 (N_322,In_685,In_15);
and U323 (N_323,N_171,In_362);
and U324 (N_324,In_12,N_137);
nand U325 (N_325,N_50,In_281);
or U326 (N_326,N_140,In_75);
and U327 (N_327,N_125,In_85);
nand U328 (N_328,In_348,N_128);
xnor U329 (N_329,N_93,In_574);
and U330 (N_330,In_546,In_652);
nand U331 (N_331,N_26,In_381);
and U332 (N_332,In_210,In_284);
or U333 (N_333,N_166,In_283);
nand U334 (N_334,In_654,In_339);
nor U335 (N_335,In_294,In_158);
nand U336 (N_336,In_680,In_416);
and U337 (N_337,N_165,In_420);
or U338 (N_338,In_68,In_160);
or U339 (N_339,In_393,In_389);
or U340 (N_340,In_494,In_485);
nor U341 (N_341,N_194,In_490);
nand U342 (N_342,N_42,In_83);
nand U343 (N_343,N_124,In_682);
nand U344 (N_344,In_137,In_740);
or U345 (N_345,In_489,In_289);
nor U346 (N_346,N_168,In_426);
and U347 (N_347,N_163,In_559);
and U348 (N_348,In_38,N_172);
nor U349 (N_349,In_292,In_508);
nand U350 (N_350,N_37,In_629);
nor U351 (N_351,N_148,In_506);
or U352 (N_352,N_129,N_145);
nor U353 (N_353,In_488,N_121);
nand U354 (N_354,In_371,In_478);
nand U355 (N_355,N_120,N_109);
or U356 (N_356,N_138,In_174);
and U357 (N_357,N_61,In_52);
nor U358 (N_358,In_101,N_198);
nand U359 (N_359,N_186,N_178);
or U360 (N_360,In_47,In_725);
and U361 (N_361,N_29,In_520);
nor U362 (N_362,In_121,N_89);
nor U363 (N_363,In_89,In_306);
and U364 (N_364,N_71,In_345);
and U365 (N_365,In_419,In_585);
nand U366 (N_366,N_31,N_83);
or U367 (N_367,In_226,In_202);
or U368 (N_368,In_6,N_117);
and U369 (N_369,In_683,N_36);
or U370 (N_370,In_97,In_497);
nand U371 (N_371,N_189,N_147);
and U372 (N_372,In_286,In_439);
and U373 (N_373,N_197,N_53);
nand U374 (N_374,In_26,In_108);
nand U375 (N_375,In_171,In_515);
and U376 (N_376,In_66,In_272);
and U377 (N_377,In_396,N_91);
nor U378 (N_378,In_271,In_199);
nand U379 (N_379,In_456,In_686);
nand U380 (N_380,In_655,In_483);
or U381 (N_381,N_97,In_205);
or U382 (N_382,In_492,In_474);
nand U383 (N_383,In_237,In_521);
nand U384 (N_384,In_63,In_363);
nor U385 (N_385,N_59,N_123);
nand U386 (N_386,In_336,In_649);
nand U387 (N_387,N_62,N_12);
nor U388 (N_388,N_181,In_361);
and U389 (N_389,In_575,N_146);
or U390 (N_390,N_22,N_115);
and U391 (N_391,N_27,N_51);
or U392 (N_392,In_305,N_0);
nor U393 (N_393,In_714,N_132);
or U394 (N_394,In_487,In_187);
and U395 (N_395,In_315,N_92);
and U396 (N_396,In_260,In_531);
nor U397 (N_397,In_693,In_46);
nor U398 (N_398,N_73,In_583);
and U399 (N_399,N_10,N_75);
nand U400 (N_400,N_281,N_386);
nor U401 (N_401,In_618,N_299);
xor U402 (N_402,N_82,N_396);
or U403 (N_403,N_23,N_28);
nor U404 (N_404,N_254,In_677);
nor U405 (N_405,N_240,N_388);
or U406 (N_406,N_350,N_342);
nand U407 (N_407,N_106,N_220);
nor U408 (N_408,In_9,N_57);
or U409 (N_409,N_169,In_432);
and U410 (N_410,N_102,N_217);
and U411 (N_411,N_357,N_143);
nand U412 (N_412,N_325,N_366);
nand U413 (N_413,In_84,N_55);
or U414 (N_414,N_283,N_383);
and U415 (N_415,N_337,In_249);
nor U416 (N_416,In_192,N_329);
nand U417 (N_417,In_727,In_458);
nand U418 (N_418,N_205,N_302);
or U419 (N_419,In_275,N_127);
nor U420 (N_420,In_378,N_345);
and U421 (N_421,N_56,N_243);
nand U422 (N_422,N_183,N_87);
nor U423 (N_423,N_225,N_266);
and U424 (N_424,In_739,N_353);
nand U425 (N_425,In_172,N_297);
nand U426 (N_426,N_211,N_9);
or U427 (N_427,N_192,N_310);
nor U428 (N_428,N_135,N_282);
nor U429 (N_429,N_308,In_667);
nor U430 (N_430,N_379,In_697);
nor U431 (N_431,N_293,N_371);
and U432 (N_432,N_355,N_213);
or U433 (N_433,In_43,In_619);
or U434 (N_434,N_214,N_176);
and U435 (N_435,N_203,N_394);
nor U436 (N_436,N_280,N_259);
nand U437 (N_437,In_227,N_290);
nor U438 (N_438,N_311,N_269);
nor U439 (N_439,N_369,N_99);
or U440 (N_440,N_235,N_74);
nand U441 (N_441,In_225,In_144);
and U442 (N_442,N_326,N_304);
nor U443 (N_443,In_340,N_3);
nand U444 (N_444,In_276,N_319);
nand U445 (N_445,N_107,In_48);
or U446 (N_446,N_66,In_102);
or U447 (N_447,N_336,N_248);
or U448 (N_448,In_147,N_250);
or U449 (N_449,In_54,N_273);
nand U450 (N_450,In_113,In_615);
or U451 (N_451,N_21,N_309);
and U452 (N_452,In_356,In_317);
and U453 (N_453,N_258,N_378);
or U454 (N_454,N_54,In_631);
nand U455 (N_455,N_237,In_704);
or U456 (N_456,N_348,N_208);
nand U457 (N_457,N_44,N_224);
or U458 (N_458,N_391,In_34);
and U459 (N_459,N_340,N_13);
nand U460 (N_460,N_382,N_314);
nor U461 (N_461,In_729,N_318);
nand U462 (N_462,N_260,N_294);
nor U463 (N_463,In_712,N_352);
and U464 (N_464,N_301,N_305);
nand U465 (N_465,N_351,N_49);
nand U466 (N_466,N_328,N_94);
nor U467 (N_467,N_347,N_359);
nand U468 (N_468,N_229,In_401);
and U469 (N_469,N_268,In_518);
or U470 (N_470,In_24,N_200);
nand U471 (N_471,In_394,N_334);
or U472 (N_472,N_333,In_299);
xnor U473 (N_473,N_244,N_343);
nand U474 (N_474,N_84,In_529);
and U475 (N_475,In_602,N_33);
xor U476 (N_476,N_313,N_286);
nand U477 (N_477,N_234,N_218);
and U478 (N_478,N_320,In_49);
nor U479 (N_479,N_68,N_372);
or U480 (N_480,N_327,N_14);
and U481 (N_481,N_278,N_144);
nor U482 (N_482,N_276,N_38);
and U483 (N_483,N_230,N_226);
nor U484 (N_484,N_322,N_374);
and U485 (N_485,N_58,N_330);
and U486 (N_486,N_18,N_399);
nor U487 (N_487,N_354,In_743);
and U488 (N_488,N_331,N_385);
and U489 (N_489,N_232,N_377);
or U490 (N_490,N_338,N_364);
nor U491 (N_491,In_670,N_277);
nand U492 (N_492,N_257,N_332);
or U493 (N_493,N_381,N_380);
and U494 (N_494,N_270,In_120);
nor U495 (N_495,N_251,In_626);
xnor U496 (N_496,N_375,N_368);
nor U497 (N_497,N_393,N_209);
and U498 (N_498,N_238,N_228);
or U499 (N_499,N_264,N_344);
and U500 (N_500,N_362,In_502);
nor U501 (N_501,N_161,In_513);
and U502 (N_502,N_79,In_581);
xnor U503 (N_503,N_201,In_60);
nor U504 (N_504,N_133,N_323);
nand U505 (N_505,In_30,N_45);
or U506 (N_506,N_363,In_466);
or U507 (N_507,N_154,N_216);
nand U508 (N_508,In_493,N_184);
nand U509 (N_509,N_134,N_223);
nand U510 (N_510,In_569,In_530);
nand U511 (N_511,N_315,In_591);
nor U512 (N_512,N_346,N_300);
xnor U513 (N_513,In_709,N_131);
nand U514 (N_514,N_262,In_404);
or U515 (N_515,N_215,N_247);
and U516 (N_516,In_572,N_349);
or U517 (N_517,N_365,N_292);
nor U518 (N_518,N_275,N_389);
and U519 (N_519,N_390,N_370);
or U520 (N_520,N_252,N_265);
and U521 (N_521,N_236,N_63);
nor U522 (N_522,N_307,N_256);
and U523 (N_523,N_119,In_309);
or U524 (N_524,N_261,In_524);
and U525 (N_525,N_397,N_398);
nand U526 (N_526,N_255,N_241);
nand U527 (N_527,N_2,N_20);
and U528 (N_528,In_154,N_356);
and U529 (N_529,N_288,In_398);
and U530 (N_530,N_298,In_433);
or U531 (N_531,N_245,N_335);
nor U532 (N_532,In_129,In_254);
nand U533 (N_533,N_239,In_723);
or U534 (N_534,N_306,N_180);
or U535 (N_535,In_151,N_312);
nor U536 (N_536,N_295,N_222);
xor U537 (N_537,N_341,N_202);
and U538 (N_538,N_274,In_507);
nor U539 (N_539,N_339,N_142);
nand U540 (N_540,N_287,N_384);
or U541 (N_541,In_554,N_227);
and U542 (N_542,N_116,N_70);
nand U543 (N_543,N_296,N_32);
nor U544 (N_544,N_376,N_212);
nand U545 (N_545,N_367,N_231);
nand U546 (N_546,N_291,N_242);
and U547 (N_547,In_578,N_182);
nand U548 (N_548,N_41,N_15);
or U549 (N_549,N_373,N_204);
nand U550 (N_550,In_87,N_179);
nand U551 (N_551,In_703,N_52);
nand U552 (N_552,N_199,In_251);
nor U553 (N_553,N_360,N_324);
nand U554 (N_554,N_387,N_285);
and U555 (N_555,In_421,N_207);
nor U556 (N_556,N_233,N_167);
nand U557 (N_557,N_358,N_316);
nand U558 (N_558,N_267,N_272);
and U559 (N_559,N_191,N_289);
or U560 (N_560,N_303,N_219);
and U561 (N_561,N_284,N_321);
and U562 (N_562,N_253,In_169);
or U563 (N_563,In_604,N_98);
nor U564 (N_564,N_263,N_105);
and U565 (N_565,In_307,N_206);
nor U566 (N_566,N_126,N_19);
and U567 (N_567,N_7,In_5);
nor U568 (N_568,N_221,N_210);
or U569 (N_569,N_361,N_392);
and U570 (N_570,In_51,N_317);
nor U571 (N_571,N_395,In_27);
nand U572 (N_572,N_279,N_246);
or U573 (N_573,N_249,In_190);
nor U574 (N_574,N_187,N_271);
nor U575 (N_575,N_356,N_126);
nand U576 (N_576,N_58,N_390);
or U577 (N_577,In_172,N_387);
and U578 (N_578,In_172,N_323);
xnor U579 (N_579,In_49,N_199);
or U580 (N_580,N_358,In_309);
nand U581 (N_581,N_285,N_15);
nand U582 (N_582,N_293,N_232);
and U583 (N_583,N_260,N_272);
or U584 (N_584,N_255,In_378);
nor U585 (N_585,N_257,In_48);
nand U586 (N_586,In_493,In_102);
or U587 (N_587,N_224,In_401);
nor U588 (N_588,N_274,N_290);
xnor U589 (N_589,N_169,N_306);
and U590 (N_590,N_259,N_376);
xor U591 (N_591,N_200,N_368);
and U592 (N_592,N_226,N_242);
or U593 (N_593,N_398,In_154);
nand U594 (N_594,N_364,In_703);
and U595 (N_595,N_267,N_328);
nand U596 (N_596,N_215,N_299);
or U597 (N_597,N_380,N_257);
nand U598 (N_598,N_235,N_79);
or U599 (N_599,In_433,N_269);
nand U600 (N_600,N_456,N_433);
nand U601 (N_601,N_581,N_544);
nor U602 (N_602,N_539,N_506);
xor U603 (N_603,N_569,N_520);
and U604 (N_604,N_494,N_548);
or U605 (N_605,N_546,N_503);
nand U606 (N_606,N_526,N_573);
nand U607 (N_607,N_462,N_452);
nand U608 (N_608,N_448,N_413);
or U609 (N_609,N_465,N_488);
or U610 (N_610,N_458,N_449);
or U611 (N_611,N_455,N_407);
nand U612 (N_612,N_599,N_565);
nor U613 (N_613,N_467,N_580);
and U614 (N_614,N_487,N_571);
or U615 (N_615,N_424,N_527);
nand U616 (N_616,N_441,N_509);
or U617 (N_617,N_475,N_552);
or U618 (N_618,N_400,N_493);
nor U619 (N_619,N_550,N_478);
and U620 (N_620,N_499,N_575);
xor U621 (N_621,N_432,N_583);
nor U622 (N_622,N_572,N_560);
nor U623 (N_623,N_577,N_439);
or U624 (N_624,N_409,N_557);
nand U625 (N_625,N_477,N_419);
or U626 (N_626,N_496,N_464);
nor U627 (N_627,N_531,N_563);
nand U628 (N_628,N_574,N_521);
or U629 (N_629,N_590,N_474);
or U630 (N_630,N_576,N_584);
or U631 (N_631,N_404,N_481);
or U632 (N_632,N_547,N_512);
nand U633 (N_633,N_533,N_588);
and U634 (N_634,N_453,N_502);
xnor U635 (N_635,N_442,N_529);
and U636 (N_636,N_589,N_587);
nor U637 (N_637,N_492,N_535);
nor U638 (N_638,N_558,N_598);
or U639 (N_639,N_554,N_418);
nand U640 (N_640,N_483,N_408);
or U641 (N_641,N_594,N_579);
or U642 (N_642,N_450,N_405);
nor U643 (N_643,N_412,N_578);
nor U644 (N_644,N_513,N_505);
and U645 (N_645,N_507,N_417);
or U646 (N_646,N_402,N_470);
or U647 (N_647,N_485,N_463);
or U648 (N_648,N_431,N_454);
or U649 (N_649,N_518,N_426);
nand U650 (N_650,N_444,N_516);
and U651 (N_651,N_446,N_422);
nor U652 (N_652,N_498,N_472);
and U653 (N_653,N_482,N_504);
xnor U654 (N_654,N_425,N_415);
nor U655 (N_655,N_559,N_410);
nor U656 (N_656,N_500,N_476);
nand U657 (N_657,N_551,N_491);
nand U658 (N_658,N_420,N_484);
nand U659 (N_659,N_468,N_423);
nand U660 (N_660,N_510,N_495);
and U661 (N_661,N_416,N_515);
nand U662 (N_662,N_480,N_597);
and U663 (N_663,N_523,N_428);
and U664 (N_664,N_469,N_460);
nand U665 (N_665,N_591,N_501);
nand U666 (N_666,N_543,N_530);
and U667 (N_667,N_568,N_430);
or U668 (N_668,N_545,N_592);
nor U669 (N_669,N_522,N_435);
or U670 (N_670,N_451,N_508);
or U671 (N_671,N_489,N_461);
and U672 (N_672,N_403,N_427);
and U673 (N_673,N_541,N_564);
nand U674 (N_674,N_537,N_479);
nor U675 (N_675,N_406,N_471);
or U676 (N_676,N_528,N_536);
nand U677 (N_677,N_582,N_538);
nand U678 (N_678,N_561,N_562);
and U679 (N_679,N_553,N_445);
nor U680 (N_680,N_542,N_429);
nand U681 (N_681,N_438,N_497);
and U682 (N_682,N_486,N_401);
or U683 (N_683,N_532,N_593);
nor U684 (N_684,N_586,N_443);
nand U685 (N_685,N_436,N_473);
or U686 (N_686,N_525,N_490);
nand U687 (N_687,N_595,N_411);
nand U688 (N_688,N_556,N_447);
or U689 (N_689,N_517,N_421);
xnor U690 (N_690,N_459,N_524);
nor U691 (N_691,N_540,N_457);
and U692 (N_692,N_511,N_437);
nor U693 (N_693,N_534,N_440);
nand U694 (N_694,N_585,N_570);
or U695 (N_695,N_549,N_514);
nand U696 (N_696,N_519,N_414);
nor U697 (N_697,N_466,N_555);
nor U698 (N_698,N_596,N_567);
nand U699 (N_699,N_434,N_566);
and U700 (N_700,N_580,N_581);
and U701 (N_701,N_539,N_505);
nand U702 (N_702,N_401,N_461);
and U703 (N_703,N_473,N_540);
or U704 (N_704,N_584,N_571);
nor U705 (N_705,N_498,N_431);
or U706 (N_706,N_412,N_538);
or U707 (N_707,N_506,N_442);
and U708 (N_708,N_458,N_452);
and U709 (N_709,N_489,N_587);
and U710 (N_710,N_560,N_541);
and U711 (N_711,N_570,N_479);
nand U712 (N_712,N_540,N_449);
nand U713 (N_713,N_454,N_539);
nand U714 (N_714,N_561,N_482);
nor U715 (N_715,N_417,N_538);
and U716 (N_716,N_422,N_597);
nand U717 (N_717,N_587,N_420);
nor U718 (N_718,N_483,N_469);
nand U719 (N_719,N_587,N_462);
or U720 (N_720,N_584,N_596);
nor U721 (N_721,N_464,N_481);
nor U722 (N_722,N_402,N_531);
nand U723 (N_723,N_482,N_592);
nor U724 (N_724,N_480,N_550);
and U725 (N_725,N_515,N_422);
and U726 (N_726,N_562,N_587);
nor U727 (N_727,N_475,N_576);
or U728 (N_728,N_551,N_508);
and U729 (N_729,N_501,N_507);
nor U730 (N_730,N_505,N_439);
nand U731 (N_731,N_501,N_401);
and U732 (N_732,N_463,N_413);
and U733 (N_733,N_532,N_466);
or U734 (N_734,N_500,N_490);
nand U735 (N_735,N_492,N_551);
or U736 (N_736,N_414,N_422);
nor U737 (N_737,N_512,N_584);
and U738 (N_738,N_577,N_579);
or U739 (N_739,N_509,N_562);
nand U740 (N_740,N_484,N_580);
or U741 (N_741,N_553,N_536);
nand U742 (N_742,N_558,N_466);
or U743 (N_743,N_585,N_415);
nand U744 (N_744,N_566,N_463);
nor U745 (N_745,N_553,N_474);
or U746 (N_746,N_435,N_441);
and U747 (N_747,N_595,N_450);
or U748 (N_748,N_513,N_573);
or U749 (N_749,N_506,N_458);
and U750 (N_750,N_466,N_574);
or U751 (N_751,N_408,N_406);
nor U752 (N_752,N_404,N_565);
or U753 (N_753,N_599,N_559);
nor U754 (N_754,N_526,N_541);
and U755 (N_755,N_435,N_541);
and U756 (N_756,N_521,N_513);
xnor U757 (N_757,N_495,N_592);
nor U758 (N_758,N_400,N_549);
and U759 (N_759,N_454,N_568);
and U760 (N_760,N_552,N_418);
and U761 (N_761,N_479,N_514);
nand U762 (N_762,N_570,N_595);
nor U763 (N_763,N_466,N_510);
and U764 (N_764,N_539,N_465);
and U765 (N_765,N_448,N_434);
nand U766 (N_766,N_416,N_500);
nand U767 (N_767,N_425,N_466);
and U768 (N_768,N_533,N_467);
and U769 (N_769,N_413,N_477);
nor U770 (N_770,N_463,N_507);
nor U771 (N_771,N_424,N_539);
nor U772 (N_772,N_584,N_430);
xor U773 (N_773,N_443,N_459);
nand U774 (N_774,N_517,N_535);
nor U775 (N_775,N_491,N_438);
or U776 (N_776,N_457,N_546);
nor U777 (N_777,N_498,N_536);
and U778 (N_778,N_530,N_411);
and U779 (N_779,N_571,N_484);
and U780 (N_780,N_444,N_405);
nor U781 (N_781,N_492,N_494);
nand U782 (N_782,N_544,N_402);
xor U783 (N_783,N_524,N_427);
nand U784 (N_784,N_411,N_483);
nand U785 (N_785,N_437,N_452);
and U786 (N_786,N_443,N_425);
and U787 (N_787,N_590,N_493);
and U788 (N_788,N_477,N_423);
nand U789 (N_789,N_471,N_402);
nor U790 (N_790,N_456,N_598);
or U791 (N_791,N_496,N_412);
nor U792 (N_792,N_458,N_583);
nand U793 (N_793,N_535,N_579);
nand U794 (N_794,N_545,N_419);
nor U795 (N_795,N_514,N_463);
or U796 (N_796,N_421,N_580);
and U797 (N_797,N_428,N_542);
and U798 (N_798,N_406,N_436);
nand U799 (N_799,N_418,N_413);
or U800 (N_800,N_678,N_797);
or U801 (N_801,N_722,N_632);
or U802 (N_802,N_753,N_617);
nand U803 (N_803,N_609,N_696);
or U804 (N_804,N_630,N_629);
or U805 (N_805,N_718,N_721);
or U806 (N_806,N_776,N_655);
xnor U807 (N_807,N_711,N_787);
nand U808 (N_808,N_642,N_663);
and U809 (N_809,N_786,N_717);
or U810 (N_810,N_633,N_656);
nor U811 (N_811,N_731,N_756);
nand U812 (N_812,N_713,N_667);
and U813 (N_813,N_768,N_765);
or U814 (N_814,N_605,N_638);
or U815 (N_815,N_720,N_612);
nand U816 (N_816,N_671,N_739);
or U817 (N_817,N_631,N_697);
and U818 (N_818,N_646,N_686);
nand U819 (N_819,N_737,N_716);
xor U820 (N_820,N_723,N_749);
nand U821 (N_821,N_637,N_674);
nor U822 (N_822,N_691,N_659);
and U823 (N_823,N_645,N_715);
and U824 (N_824,N_784,N_788);
nand U825 (N_825,N_771,N_729);
or U826 (N_826,N_750,N_602);
nand U827 (N_827,N_708,N_685);
or U828 (N_828,N_651,N_608);
or U829 (N_829,N_618,N_647);
nor U830 (N_830,N_625,N_763);
or U831 (N_831,N_764,N_735);
nor U832 (N_832,N_798,N_707);
nand U833 (N_833,N_702,N_782);
nand U834 (N_834,N_773,N_772);
and U835 (N_835,N_619,N_622);
or U836 (N_836,N_610,N_687);
nor U837 (N_837,N_639,N_699);
nor U838 (N_838,N_653,N_675);
nand U839 (N_839,N_614,N_693);
and U840 (N_840,N_760,N_726);
and U841 (N_841,N_751,N_741);
and U842 (N_842,N_635,N_725);
and U843 (N_843,N_681,N_620);
nor U844 (N_844,N_689,N_601);
nand U845 (N_845,N_661,N_613);
or U846 (N_846,N_746,N_793);
nor U847 (N_847,N_742,N_775);
and U848 (N_848,N_727,N_740);
and U849 (N_849,N_759,N_606);
or U850 (N_850,N_748,N_701);
nand U851 (N_851,N_666,N_781);
or U852 (N_852,N_660,N_774);
nand U853 (N_853,N_744,N_680);
nor U854 (N_854,N_624,N_700);
nor U855 (N_855,N_709,N_785);
and U856 (N_856,N_615,N_662);
or U857 (N_857,N_692,N_728);
and U858 (N_858,N_743,N_752);
or U859 (N_859,N_669,N_683);
nor U860 (N_860,N_791,N_623);
and U861 (N_861,N_652,N_698);
nand U862 (N_862,N_626,N_736);
nand U863 (N_863,N_790,N_799);
or U864 (N_864,N_688,N_738);
nand U865 (N_865,N_673,N_650);
nand U866 (N_866,N_732,N_611);
nand U867 (N_867,N_757,N_754);
nand U868 (N_868,N_644,N_794);
nor U869 (N_869,N_677,N_648);
and U870 (N_870,N_694,N_734);
and U871 (N_871,N_766,N_628);
or U872 (N_872,N_657,N_770);
nor U873 (N_873,N_724,N_719);
nand U874 (N_874,N_780,N_733);
nand U875 (N_875,N_649,N_640);
and U876 (N_876,N_796,N_695);
nor U877 (N_877,N_705,N_676);
and U878 (N_878,N_747,N_710);
nand U879 (N_879,N_714,N_758);
and U880 (N_880,N_665,N_634);
nor U881 (N_881,N_603,N_712);
or U882 (N_882,N_636,N_703);
and U883 (N_883,N_641,N_745);
nand U884 (N_884,N_654,N_682);
xnor U885 (N_885,N_706,N_627);
or U886 (N_886,N_643,N_684);
or U887 (N_887,N_679,N_621);
and U888 (N_888,N_761,N_730);
nor U889 (N_889,N_769,N_600);
or U890 (N_890,N_704,N_783);
and U891 (N_891,N_779,N_658);
nor U892 (N_892,N_690,N_616);
nor U893 (N_893,N_795,N_670);
and U894 (N_894,N_668,N_777);
or U895 (N_895,N_672,N_607);
and U896 (N_896,N_778,N_604);
nor U897 (N_897,N_767,N_664);
and U898 (N_898,N_792,N_789);
xor U899 (N_899,N_762,N_755);
nor U900 (N_900,N_618,N_625);
nand U901 (N_901,N_775,N_656);
or U902 (N_902,N_758,N_734);
xnor U903 (N_903,N_611,N_663);
nand U904 (N_904,N_692,N_638);
nand U905 (N_905,N_697,N_641);
nand U906 (N_906,N_678,N_773);
or U907 (N_907,N_777,N_651);
nand U908 (N_908,N_778,N_723);
and U909 (N_909,N_653,N_657);
or U910 (N_910,N_684,N_795);
nor U911 (N_911,N_617,N_635);
nand U912 (N_912,N_677,N_798);
xor U913 (N_913,N_718,N_701);
or U914 (N_914,N_794,N_661);
nor U915 (N_915,N_725,N_784);
nand U916 (N_916,N_793,N_788);
or U917 (N_917,N_723,N_767);
or U918 (N_918,N_688,N_638);
and U919 (N_919,N_719,N_607);
or U920 (N_920,N_678,N_698);
or U921 (N_921,N_739,N_669);
or U922 (N_922,N_739,N_765);
or U923 (N_923,N_798,N_699);
or U924 (N_924,N_748,N_676);
nor U925 (N_925,N_687,N_760);
xor U926 (N_926,N_621,N_605);
nor U927 (N_927,N_648,N_622);
or U928 (N_928,N_630,N_699);
nor U929 (N_929,N_745,N_609);
nor U930 (N_930,N_793,N_649);
and U931 (N_931,N_736,N_661);
nand U932 (N_932,N_727,N_730);
nand U933 (N_933,N_674,N_741);
nor U934 (N_934,N_749,N_718);
and U935 (N_935,N_673,N_794);
nand U936 (N_936,N_601,N_733);
or U937 (N_937,N_762,N_682);
nand U938 (N_938,N_600,N_719);
or U939 (N_939,N_666,N_620);
or U940 (N_940,N_687,N_609);
nor U941 (N_941,N_735,N_753);
nor U942 (N_942,N_615,N_778);
nand U943 (N_943,N_655,N_628);
nand U944 (N_944,N_737,N_753);
nor U945 (N_945,N_601,N_766);
nor U946 (N_946,N_772,N_739);
nand U947 (N_947,N_624,N_699);
and U948 (N_948,N_727,N_724);
or U949 (N_949,N_665,N_620);
nor U950 (N_950,N_662,N_761);
nand U951 (N_951,N_742,N_675);
nand U952 (N_952,N_687,N_755);
or U953 (N_953,N_632,N_624);
and U954 (N_954,N_643,N_769);
nor U955 (N_955,N_685,N_701);
and U956 (N_956,N_630,N_695);
nand U957 (N_957,N_779,N_631);
or U958 (N_958,N_651,N_640);
and U959 (N_959,N_793,N_647);
nor U960 (N_960,N_754,N_632);
or U961 (N_961,N_673,N_674);
nand U962 (N_962,N_735,N_650);
and U963 (N_963,N_688,N_770);
nand U964 (N_964,N_796,N_789);
nand U965 (N_965,N_632,N_757);
or U966 (N_966,N_744,N_696);
nand U967 (N_967,N_609,N_771);
or U968 (N_968,N_747,N_644);
and U969 (N_969,N_613,N_736);
or U970 (N_970,N_732,N_682);
or U971 (N_971,N_778,N_666);
nor U972 (N_972,N_728,N_723);
and U973 (N_973,N_654,N_627);
nor U974 (N_974,N_645,N_785);
nand U975 (N_975,N_690,N_643);
nor U976 (N_976,N_699,N_663);
nand U977 (N_977,N_730,N_647);
or U978 (N_978,N_734,N_692);
nor U979 (N_979,N_723,N_739);
nand U980 (N_980,N_615,N_744);
nor U981 (N_981,N_670,N_740);
or U982 (N_982,N_646,N_654);
nor U983 (N_983,N_730,N_668);
nand U984 (N_984,N_625,N_646);
or U985 (N_985,N_683,N_641);
or U986 (N_986,N_692,N_748);
nand U987 (N_987,N_742,N_692);
xnor U988 (N_988,N_750,N_645);
nand U989 (N_989,N_733,N_796);
and U990 (N_990,N_641,N_739);
or U991 (N_991,N_633,N_610);
xor U992 (N_992,N_636,N_741);
or U993 (N_993,N_683,N_694);
nor U994 (N_994,N_642,N_752);
nand U995 (N_995,N_607,N_783);
nand U996 (N_996,N_696,N_672);
nand U997 (N_997,N_717,N_771);
or U998 (N_998,N_721,N_749);
or U999 (N_999,N_722,N_671);
nor U1000 (N_1000,N_918,N_989);
nand U1001 (N_1001,N_987,N_895);
and U1002 (N_1002,N_964,N_879);
nor U1003 (N_1003,N_859,N_944);
nand U1004 (N_1004,N_864,N_839);
nand U1005 (N_1005,N_829,N_940);
nand U1006 (N_1006,N_965,N_926);
or U1007 (N_1007,N_919,N_809);
nor U1008 (N_1008,N_922,N_976);
and U1009 (N_1009,N_907,N_913);
or U1010 (N_1010,N_961,N_805);
nand U1011 (N_1011,N_868,N_885);
nand U1012 (N_1012,N_953,N_818);
nor U1013 (N_1013,N_883,N_932);
nand U1014 (N_1014,N_956,N_977);
nand U1015 (N_1015,N_901,N_996);
and U1016 (N_1016,N_933,N_851);
nand U1017 (N_1017,N_929,N_857);
nand U1018 (N_1018,N_832,N_936);
nand U1019 (N_1019,N_867,N_894);
nand U1020 (N_1020,N_998,N_840);
or U1021 (N_1021,N_821,N_955);
and U1022 (N_1022,N_822,N_993);
nor U1023 (N_1023,N_988,N_862);
nor U1024 (N_1024,N_899,N_824);
or U1025 (N_1025,N_905,N_957);
and U1026 (N_1026,N_937,N_860);
nor U1027 (N_1027,N_872,N_952);
and U1028 (N_1028,N_896,N_854);
and U1029 (N_1029,N_935,N_808);
and U1030 (N_1030,N_915,N_865);
or U1031 (N_1031,N_878,N_975);
nor U1032 (N_1032,N_980,N_877);
and U1033 (N_1033,N_902,N_984);
nand U1034 (N_1034,N_870,N_900);
nand U1035 (N_1035,N_881,N_819);
nand U1036 (N_1036,N_991,N_814);
or U1037 (N_1037,N_921,N_817);
xnor U1038 (N_1038,N_835,N_999);
nor U1039 (N_1039,N_972,N_973);
nand U1040 (N_1040,N_982,N_880);
or U1041 (N_1041,N_853,N_960);
or U1042 (N_1042,N_904,N_979);
nand U1043 (N_1043,N_820,N_855);
nand U1044 (N_1044,N_992,N_962);
or U1045 (N_1045,N_866,N_924);
nor U1046 (N_1046,N_847,N_946);
nor U1047 (N_1047,N_945,N_848);
nand U1048 (N_1048,N_836,N_861);
or U1049 (N_1049,N_898,N_858);
nor U1050 (N_1050,N_920,N_897);
nor U1051 (N_1051,N_838,N_951);
or U1052 (N_1052,N_888,N_931);
nand U1053 (N_1053,N_806,N_971);
and U1054 (N_1054,N_974,N_815);
and U1055 (N_1055,N_846,N_909);
or U1056 (N_1056,N_802,N_947);
nand U1057 (N_1057,N_810,N_893);
nor U1058 (N_1058,N_834,N_903);
nor U1059 (N_1059,N_990,N_930);
nor U1060 (N_1060,N_911,N_830);
or U1061 (N_1061,N_890,N_925);
xnor U1062 (N_1062,N_912,N_831);
nand U1063 (N_1063,N_950,N_923);
or U1064 (N_1064,N_869,N_811);
nand U1065 (N_1065,N_871,N_967);
and U1066 (N_1066,N_826,N_997);
and U1067 (N_1067,N_886,N_934);
or U1068 (N_1068,N_954,N_966);
or U1069 (N_1069,N_943,N_889);
or U1070 (N_1070,N_842,N_876);
xnor U1071 (N_1071,N_882,N_985);
nand U1072 (N_1072,N_978,N_875);
nor U1073 (N_1073,N_927,N_849);
nand U1074 (N_1074,N_969,N_908);
or U1075 (N_1075,N_887,N_917);
or U1076 (N_1076,N_823,N_843);
xor U1077 (N_1077,N_884,N_828);
and U1078 (N_1078,N_833,N_910);
nand U1079 (N_1079,N_959,N_995);
nor U1080 (N_1080,N_941,N_916);
nand U1081 (N_1081,N_892,N_825);
and U1082 (N_1082,N_873,N_928);
and U1083 (N_1083,N_939,N_981);
nor U1084 (N_1084,N_942,N_845);
xor U1085 (N_1085,N_856,N_906);
or U1086 (N_1086,N_807,N_958);
and U1087 (N_1087,N_837,N_804);
or U1088 (N_1088,N_983,N_914);
nor U1089 (N_1089,N_852,N_949);
or U1090 (N_1090,N_863,N_968);
nor U1091 (N_1091,N_948,N_850);
and U1092 (N_1092,N_812,N_970);
nor U1093 (N_1093,N_986,N_827);
nand U1094 (N_1094,N_938,N_844);
nand U1095 (N_1095,N_801,N_891);
nand U1096 (N_1096,N_874,N_963);
or U1097 (N_1097,N_803,N_800);
and U1098 (N_1098,N_841,N_994);
nor U1099 (N_1099,N_813,N_816);
nand U1100 (N_1100,N_829,N_838);
nand U1101 (N_1101,N_876,N_883);
and U1102 (N_1102,N_822,N_838);
and U1103 (N_1103,N_873,N_812);
nand U1104 (N_1104,N_965,N_942);
or U1105 (N_1105,N_831,N_936);
nand U1106 (N_1106,N_976,N_989);
nand U1107 (N_1107,N_861,N_804);
nand U1108 (N_1108,N_852,N_918);
nand U1109 (N_1109,N_847,N_882);
and U1110 (N_1110,N_869,N_890);
nand U1111 (N_1111,N_868,N_942);
and U1112 (N_1112,N_868,N_923);
and U1113 (N_1113,N_863,N_886);
or U1114 (N_1114,N_836,N_985);
xor U1115 (N_1115,N_925,N_882);
nand U1116 (N_1116,N_990,N_835);
or U1117 (N_1117,N_895,N_806);
nor U1118 (N_1118,N_815,N_857);
nor U1119 (N_1119,N_842,N_848);
nor U1120 (N_1120,N_960,N_863);
nand U1121 (N_1121,N_914,N_937);
and U1122 (N_1122,N_980,N_922);
nor U1123 (N_1123,N_887,N_872);
or U1124 (N_1124,N_974,N_807);
and U1125 (N_1125,N_979,N_911);
nand U1126 (N_1126,N_882,N_801);
or U1127 (N_1127,N_895,N_804);
and U1128 (N_1128,N_903,N_910);
nor U1129 (N_1129,N_999,N_907);
and U1130 (N_1130,N_870,N_919);
nand U1131 (N_1131,N_945,N_896);
nor U1132 (N_1132,N_970,N_956);
and U1133 (N_1133,N_907,N_937);
or U1134 (N_1134,N_977,N_963);
and U1135 (N_1135,N_955,N_964);
and U1136 (N_1136,N_985,N_941);
nor U1137 (N_1137,N_818,N_939);
nand U1138 (N_1138,N_992,N_822);
or U1139 (N_1139,N_891,N_984);
nand U1140 (N_1140,N_804,N_834);
and U1141 (N_1141,N_881,N_843);
and U1142 (N_1142,N_868,N_859);
nor U1143 (N_1143,N_944,N_974);
or U1144 (N_1144,N_998,N_999);
nand U1145 (N_1145,N_903,N_918);
nand U1146 (N_1146,N_978,N_974);
or U1147 (N_1147,N_919,N_859);
nand U1148 (N_1148,N_904,N_876);
nand U1149 (N_1149,N_829,N_910);
nand U1150 (N_1150,N_948,N_933);
nor U1151 (N_1151,N_982,N_863);
or U1152 (N_1152,N_829,N_887);
and U1153 (N_1153,N_898,N_914);
or U1154 (N_1154,N_802,N_949);
and U1155 (N_1155,N_833,N_885);
and U1156 (N_1156,N_825,N_997);
nor U1157 (N_1157,N_975,N_853);
or U1158 (N_1158,N_917,N_975);
or U1159 (N_1159,N_919,N_824);
and U1160 (N_1160,N_872,N_846);
nand U1161 (N_1161,N_889,N_919);
nor U1162 (N_1162,N_895,N_924);
and U1163 (N_1163,N_966,N_894);
or U1164 (N_1164,N_878,N_800);
and U1165 (N_1165,N_835,N_930);
and U1166 (N_1166,N_831,N_844);
and U1167 (N_1167,N_857,N_908);
nand U1168 (N_1168,N_985,N_948);
or U1169 (N_1169,N_876,N_976);
nor U1170 (N_1170,N_907,N_860);
nand U1171 (N_1171,N_885,N_986);
nor U1172 (N_1172,N_892,N_908);
or U1173 (N_1173,N_938,N_880);
and U1174 (N_1174,N_980,N_921);
or U1175 (N_1175,N_929,N_996);
or U1176 (N_1176,N_942,N_822);
nand U1177 (N_1177,N_879,N_833);
nand U1178 (N_1178,N_867,N_921);
or U1179 (N_1179,N_911,N_804);
nor U1180 (N_1180,N_922,N_826);
and U1181 (N_1181,N_880,N_999);
or U1182 (N_1182,N_923,N_833);
or U1183 (N_1183,N_833,N_802);
nand U1184 (N_1184,N_964,N_807);
nand U1185 (N_1185,N_829,N_929);
and U1186 (N_1186,N_823,N_827);
and U1187 (N_1187,N_938,N_916);
xnor U1188 (N_1188,N_991,N_804);
nand U1189 (N_1189,N_839,N_994);
nor U1190 (N_1190,N_962,N_924);
and U1191 (N_1191,N_875,N_981);
or U1192 (N_1192,N_931,N_954);
nor U1193 (N_1193,N_827,N_819);
nand U1194 (N_1194,N_828,N_893);
and U1195 (N_1195,N_951,N_895);
nand U1196 (N_1196,N_901,N_841);
or U1197 (N_1197,N_845,N_804);
nor U1198 (N_1198,N_928,N_858);
nor U1199 (N_1199,N_930,N_848);
and U1200 (N_1200,N_1143,N_1100);
and U1201 (N_1201,N_1130,N_1071);
or U1202 (N_1202,N_1061,N_1060);
nand U1203 (N_1203,N_1015,N_1162);
or U1204 (N_1204,N_1000,N_1118);
nand U1205 (N_1205,N_1055,N_1051);
nand U1206 (N_1206,N_1020,N_1086);
or U1207 (N_1207,N_1067,N_1117);
nor U1208 (N_1208,N_1093,N_1003);
nor U1209 (N_1209,N_1062,N_1195);
nand U1210 (N_1210,N_1053,N_1039);
nor U1211 (N_1211,N_1121,N_1108);
nand U1212 (N_1212,N_1097,N_1024);
nand U1213 (N_1213,N_1157,N_1150);
or U1214 (N_1214,N_1198,N_1132);
and U1215 (N_1215,N_1068,N_1038);
nand U1216 (N_1216,N_1165,N_1006);
and U1217 (N_1217,N_1169,N_1016);
nor U1218 (N_1218,N_1023,N_1002);
nand U1219 (N_1219,N_1173,N_1104);
or U1220 (N_1220,N_1095,N_1014);
and U1221 (N_1221,N_1171,N_1145);
nor U1222 (N_1222,N_1153,N_1184);
nand U1223 (N_1223,N_1052,N_1054);
xor U1224 (N_1224,N_1126,N_1156);
or U1225 (N_1225,N_1098,N_1012);
and U1226 (N_1226,N_1158,N_1091);
nand U1227 (N_1227,N_1137,N_1042);
xor U1228 (N_1228,N_1070,N_1072);
nor U1229 (N_1229,N_1155,N_1044);
and U1230 (N_1230,N_1112,N_1160);
xnor U1231 (N_1231,N_1176,N_1084);
nor U1232 (N_1232,N_1167,N_1017);
nor U1233 (N_1233,N_1058,N_1078);
nand U1234 (N_1234,N_1115,N_1107);
or U1235 (N_1235,N_1131,N_1057);
nor U1236 (N_1236,N_1110,N_1151);
nand U1237 (N_1237,N_1037,N_1188);
or U1238 (N_1238,N_1141,N_1147);
nor U1239 (N_1239,N_1133,N_1127);
and U1240 (N_1240,N_1082,N_1076);
nand U1241 (N_1241,N_1085,N_1013);
and U1242 (N_1242,N_1026,N_1036);
and U1243 (N_1243,N_1181,N_1090);
nand U1244 (N_1244,N_1103,N_1134);
or U1245 (N_1245,N_1140,N_1018);
and U1246 (N_1246,N_1030,N_1029);
and U1247 (N_1247,N_1106,N_1022);
nor U1248 (N_1248,N_1081,N_1119);
nor U1249 (N_1249,N_1152,N_1066);
or U1250 (N_1250,N_1142,N_1019);
or U1251 (N_1251,N_1166,N_1148);
nor U1252 (N_1252,N_1089,N_1077);
nor U1253 (N_1253,N_1175,N_1164);
nand U1254 (N_1254,N_1114,N_1008);
or U1255 (N_1255,N_1028,N_1128);
nand U1256 (N_1256,N_1179,N_1087);
nand U1257 (N_1257,N_1180,N_1083);
nor U1258 (N_1258,N_1190,N_1174);
nand U1259 (N_1259,N_1170,N_1080);
nand U1260 (N_1260,N_1111,N_1079);
nor U1261 (N_1261,N_1031,N_1113);
nor U1262 (N_1262,N_1161,N_1043);
and U1263 (N_1263,N_1004,N_1194);
nand U1264 (N_1264,N_1009,N_1059);
and U1265 (N_1265,N_1183,N_1001);
xnor U1266 (N_1266,N_1191,N_1138);
or U1267 (N_1267,N_1032,N_1050);
and U1268 (N_1268,N_1049,N_1047);
nand U1269 (N_1269,N_1199,N_1189);
nor U1270 (N_1270,N_1005,N_1123);
nand U1271 (N_1271,N_1092,N_1192);
or U1272 (N_1272,N_1186,N_1048);
or U1273 (N_1273,N_1196,N_1064);
and U1274 (N_1274,N_1056,N_1159);
or U1275 (N_1275,N_1094,N_1125);
nor U1276 (N_1276,N_1177,N_1146);
and U1277 (N_1277,N_1025,N_1109);
nor U1278 (N_1278,N_1099,N_1011);
or U1279 (N_1279,N_1010,N_1124);
or U1280 (N_1280,N_1073,N_1007);
or U1281 (N_1281,N_1120,N_1033);
or U1282 (N_1282,N_1197,N_1172);
or U1283 (N_1283,N_1101,N_1045);
or U1284 (N_1284,N_1187,N_1041);
or U1285 (N_1285,N_1027,N_1096);
nand U1286 (N_1286,N_1065,N_1040);
or U1287 (N_1287,N_1129,N_1182);
or U1288 (N_1288,N_1122,N_1034);
or U1289 (N_1289,N_1144,N_1035);
xnor U1290 (N_1290,N_1088,N_1075);
nor U1291 (N_1291,N_1178,N_1074);
and U1292 (N_1292,N_1149,N_1069);
and U1293 (N_1293,N_1185,N_1021);
nand U1294 (N_1294,N_1046,N_1136);
or U1295 (N_1295,N_1168,N_1102);
and U1296 (N_1296,N_1105,N_1154);
xnor U1297 (N_1297,N_1135,N_1193);
or U1298 (N_1298,N_1139,N_1116);
nor U1299 (N_1299,N_1163,N_1063);
and U1300 (N_1300,N_1066,N_1093);
and U1301 (N_1301,N_1197,N_1052);
nor U1302 (N_1302,N_1063,N_1029);
nor U1303 (N_1303,N_1198,N_1157);
and U1304 (N_1304,N_1059,N_1037);
nand U1305 (N_1305,N_1124,N_1065);
nor U1306 (N_1306,N_1171,N_1079);
and U1307 (N_1307,N_1031,N_1197);
nand U1308 (N_1308,N_1037,N_1161);
or U1309 (N_1309,N_1094,N_1155);
nor U1310 (N_1310,N_1090,N_1150);
and U1311 (N_1311,N_1121,N_1055);
nor U1312 (N_1312,N_1074,N_1166);
nand U1313 (N_1313,N_1164,N_1071);
or U1314 (N_1314,N_1185,N_1018);
nor U1315 (N_1315,N_1169,N_1160);
and U1316 (N_1316,N_1117,N_1017);
or U1317 (N_1317,N_1165,N_1132);
nand U1318 (N_1318,N_1023,N_1158);
or U1319 (N_1319,N_1149,N_1139);
nand U1320 (N_1320,N_1191,N_1155);
nand U1321 (N_1321,N_1017,N_1052);
nor U1322 (N_1322,N_1024,N_1107);
nor U1323 (N_1323,N_1005,N_1109);
nand U1324 (N_1324,N_1019,N_1055);
and U1325 (N_1325,N_1199,N_1040);
nor U1326 (N_1326,N_1162,N_1005);
nand U1327 (N_1327,N_1182,N_1134);
nand U1328 (N_1328,N_1147,N_1018);
nand U1329 (N_1329,N_1094,N_1197);
nor U1330 (N_1330,N_1010,N_1123);
nand U1331 (N_1331,N_1100,N_1190);
nor U1332 (N_1332,N_1013,N_1041);
nor U1333 (N_1333,N_1156,N_1090);
and U1334 (N_1334,N_1091,N_1066);
nand U1335 (N_1335,N_1174,N_1107);
nor U1336 (N_1336,N_1063,N_1189);
nand U1337 (N_1337,N_1117,N_1131);
and U1338 (N_1338,N_1051,N_1147);
nand U1339 (N_1339,N_1153,N_1168);
nor U1340 (N_1340,N_1079,N_1067);
nand U1341 (N_1341,N_1032,N_1016);
or U1342 (N_1342,N_1040,N_1002);
xor U1343 (N_1343,N_1104,N_1017);
nand U1344 (N_1344,N_1159,N_1046);
and U1345 (N_1345,N_1178,N_1115);
or U1346 (N_1346,N_1013,N_1068);
nand U1347 (N_1347,N_1065,N_1021);
nand U1348 (N_1348,N_1116,N_1103);
nor U1349 (N_1349,N_1196,N_1093);
or U1350 (N_1350,N_1067,N_1179);
nand U1351 (N_1351,N_1156,N_1154);
nand U1352 (N_1352,N_1092,N_1137);
and U1353 (N_1353,N_1029,N_1177);
nor U1354 (N_1354,N_1189,N_1031);
nor U1355 (N_1355,N_1074,N_1194);
nor U1356 (N_1356,N_1078,N_1022);
or U1357 (N_1357,N_1065,N_1066);
nor U1358 (N_1358,N_1028,N_1156);
nor U1359 (N_1359,N_1012,N_1071);
and U1360 (N_1360,N_1115,N_1116);
nand U1361 (N_1361,N_1062,N_1199);
and U1362 (N_1362,N_1110,N_1033);
nand U1363 (N_1363,N_1036,N_1177);
nor U1364 (N_1364,N_1036,N_1160);
nor U1365 (N_1365,N_1030,N_1120);
or U1366 (N_1366,N_1198,N_1120);
nand U1367 (N_1367,N_1198,N_1129);
nor U1368 (N_1368,N_1149,N_1151);
nand U1369 (N_1369,N_1115,N_1058);
nand U1370 (N_1370,N_1195,N_1013);
nor U1371 (N_1371,N_1046,N_1158);
and U1372 (N_1372,N_1073,N_1076);
nand U1373 (N_1373,N_1161,N_1172);
xnor U1374 (N_1374,N_1095,N_1100);
nand U1375 (N_1375,N_1073,N_1154);
or U1376 (N_1376,N_1135,N_1101);
nor U1377 (N_1377,N_1058,N_1069);
and U1378 (N_1378,N_1101,N_1037);
and U1379 (N_1379,N_1196,N_1123);
nor U1380 (N_1380,N_1103,N_1188);
nor U1381 (N_1381,N_1065,N_1031);
or U1382 (N_1382,N_1105,N_1002);
or U1383 (N_1383,N_1017,N_1074);
and U1384 (N_1384,N_1111,N_1048);
nor U1385 (N_1385,N_1137,N_1023);
nand U1386 (N_1386,N_1023,N_1080);
nand U1387 (N_1387,N_1134,N_1163);
and U1388 (N_1388,N_1172,N_1066);
nand U1389 (N_1389,N_1036,N_1137);
nand U1390 (N_1390,N_1183,N_1120);
and U1391 (N_1391,N_1188,N_1157);
nor U1392 (N_1392,N_1006,N_1087);
nand U1393 (N_1393,N_1080,N_1101);
nand U1394 (N_1394,N_1102,N_1021);
nor U1395 (N_1395,N_1101,N_1082);
or U1396 (N_1396,N_1198,N_1000);
nor U1397 (N_1397,N_1107,N_1007);
nand U1398 (N_1398,N_1089,N_1090);
nand U1399 (N_1399,N_1040,N_1154);
and U1400 (N_1400,N_1309,N_1338);
or U1401 (N_1401,N_1241,N_1378);
or U1402 (N_1402,N_1208,N_1250);
and U1403 (N_1403,N_1304,N_1365);
or U1404 (N_1404,N_1222,N_1300);
and U1405 (N_1405,N_1218,N_1217);
nand U1406 (N_1406,N_1370,N_1322);
nand U1407 (N_1407,N_1392,N_1281);
and U1408 (N_1408,N_1349,N_1390);
or U1409 (N_1409,N_1221,N_1228);
and U1410 (N_1410,N_1227,N_1280);
nand U1411 (N_1411,N_1274,N_1331);
and U1412 (N_1412,N_1240,N_1375);
or U1413 (N_1413,N_1282,N_1332);
or U1414 (N_1414,N_1377,N_1284);
xnor U1415 (N_1415,N_1290,N_1333);
nand U1416 (N_1416,N_1383,N_1330);
xnor U1417 (N_1417,N_1379,N_1318);
and U1418 (N_1418,N_1277,N_1291);
xnor U1419 (N_1419,N_1200,N_1275);
and U1420 (N_1420,N_1233,N_1232);
or U1421 (N_1421,N_1235,N_1276);
and U1422 (N_1422,N_1323,N_1261);
nand U1423 (N_1423,N_1213,N_1388);
nand U1424 (N_1424,N_1285,N_1385);
nand U1425 (N_1425,N_1267,N_1381);
nor U1426 (N_1426,N_1348,N_1342);
or U1427 (N_1427,N_1212,N_1236);
or U1428 (N_1428,N_1289,N_1354);
nand U1429 (N_1429,N_1363,N_1269);
and U1430 (N_1430,N_1335,N_1319);
nor U1431 (N_1431,N_1268,N_1367);
or U1432 (N_1432,N_1242,N_1345);
nand U1433 (N_1433,N_1223,N_1373);
nor U1434 (N_1434,N_1328,N_1359);
and U1435 (N_1435,N_1211,N_1288);
and U1436 (N_1436,N_1397,N_1203);
or U1437 (N_1437,N_1204,N_1247);
nand U1438 (N_1438,N_1272,N_1329);
nor U1439 (N_1439,N_1244,N_1382);
nor U1440 (N_1440,N_1380,N_1337);
or U1441 (N_1441,N_1362,N_1327);
and U1442 (N_1442,N_1237,N_1395);
and U1443 (N_1443,N_1265,N_1339);
and U1444 (N_1444,N_1286,N_1202);
nand U1445 (N_1445,N_1372,N_1316);
nor U1446 (N_1446,N_1279,N_1324);
xor U1447 (N_1447,N_1243,N_1283);
nand U1448 (N_1448,N_1389,N_1302);
or U1449 (N_1449,N_1303,N_1201);
nand U1450 (N_1450,N_1371,N_1253);
or U1451 (N_1451,N_1234,N_1256);
or U1452 (N_1452,N_1229,N_1313);
nand U1453 (N_1453,N_1273,N_1312);
nor U1454 (N_1454,N_1317,N_1364);
and U1455 (N_1455,N_1393,N_1245);
or U1456 (N_1456,N_1311,N_1287);
nor U1457 (N_1457,N_1344,N_1366);
nand U1458 (N_1458,N_1216,N_1399);
nand U1459 (N_1459,N_1266,N_1356);
or U1460 (N_1460,N_1310,N_1258);
or U1461 (N_1461,N_1321,N_1326);
nand U1462 (N_1462,N_1263,N_1355);
nor U1463 (N_1463,N_1357,N_1398);
nor U1464 (N_1464,N_1320,N_1219);
and U1465 (N_1465,N_1301,N_1376);
and U1466 (N_1466,N_1278,N_1308);
or U1467 (N_1467,N_1350,N_1210);
nand U1468 (N_1468,N_1226,N_1297);
nor U1469 (N_1469,N_1358,N_1340);
nand U1470 (N_1470,N_1295,N_1346);
nor U1471 (N_1471,N_1343,N_1205);
nand U1472 (N_1472,N_1292,N_1239);
or U1473 (N_1473,N_1293,N_1207);
or U1474 (N_1474,N_1246,N_1214);
and U1475 (N_1475,N_1351,N_1353);
nor U1476 (N_1476,N_1225,N_1255);
nand U1477 (N_1477,N_1209,N_1386);
and U1478 (N_1478,N_1259,N_1252);
nor U1479 (N_1479,N_1260,N_1238);
and U1480 (N_1480,N_1249,N_1257);
nor U1481 (N_1481,N_1341,N_1206);
xor U1482 (N_1482,N_1306,N_1220);
nand U1483 (N_1483,N_1271,N_1325);
nor U1484 (N_1484,N_1387,N_1262);
or U1485 (N_1485,N_1299,N_1254);
xnor U1486 (N_1486,N_1314,N_1360);
and U1487 (N_1487,N_1315,N_1298);
nand U1488 (N_1488,N_1384,N_1215);
nor U1489 (N_1489,N_1361,N_1305);
nor U1490 (N_1490,N_1391,N_1264);
and U1491 (N_1491,N_1231,N_1369);
or U1492 (N_1492,N_1368,N_1374);
and U1493 (N_1493,N_1270,N_1294);
and U1494 (N_1494,N_1251,N_1296);
or U1495 (N_1495,N_1248,N_1336);
and U1496 (N_1496,N_1396,N_1224);
or U1497 (N_1497,N_1307,N_1334);
or U1498 (N_1498,N_1394,N_1230);
and U1499 (N_1499,N_1352,N_1347);
nor U1500 (N_1500,N_1212,N_1323);
nor U1501 (N_1501,N_1266,N_1241);
nand U1502 (N_1502,N_1344,N_1370);
nor U1503 (N_1503,N_1396,N_1288);
and U1504 (N_1504,N_1397,N_1297);
or U1505 (N_1505,N_1342,N_1393);
nand U1506 (N_1506,N_1252,N_1257);
nand U1507 (N_1507,N_1296,N_1311);
nor U1508 (N_1508,N_1370,N_1317);
and U1509 (N_1509,N_1284,N_1364);
nor U1510 (N_1510,N_1206,N_1233);
or U1511 (N_1511,N_1235,N_1200);
nor U1512 (N_1512,N_1225,N_1210);
or U1513 (N_1513,N_1369,N_1201);
nand U1514 (N_1514,N_1223,N_1287);
and U1515 (N_1515,N_1241,N_1392);
nor U1516 (N_1516,N_1216,N_1264);
and U1517 (N_1517,N_1378,N_1360);
nor U1518 (N_1518,N_1214,N_1283);
or U1519 (N_1519,N_1350,N_1285);
or U1520 (N_1520,N_1318,N_1225);
or U1521 (N_1521,N_1279,N_1229);
nand U1522 (N_1522,N_1233,N_1286);
nor U1523 (N_1523,N_1368,N_1355);
nor U1524 (N_1524,N_1309,N_1369);
nor U1525 (N_1525,N_1392,N_1375);
nor U1526 (N_1526,N_1389,N_1275);
and U1527 (N_1527,N_1331,N_1335);
nand U1528 (N_1528,N_1373,N_1204);
xor U1529 (N_1529,N_1382,N_1248);
xor U1530 (N_1530,N_1346,N_1238);
nand U1531 (N_1531,N_1380,N_1343);
or U1532 (N_1532,N_1211,N_1269);
or U1533 (N_1533,N_1396,N_1325);
or U1534 (N_1534,N_1217,N_1272);
or U1535 (N_1535,N_1388,N_1200);
or U1536 (N_1536,N_1396,N_1230);
or U1537 (N_1537,N_1226,N_1383);
nor U1538 (N_1538,N_1277,N_1311);
nand U1539 (N_1539,N_1292,N_1203);
nand U1540 (N_1540,N_1257,N_1338);
xor U1541 (N_1541,N_1266,N_1393);
nor U1542 (N_1542,N_1247,N_1242);
and U1543 (N_1543,N_1220,N_1349);
nor U1544 (N_1544,N_1236,N_1388);
nand U1545 (N_1545,N_1308,N_1276);
and U1546 (N_1546,N_1386,N_1304);
nand U1547 (N_1547,N_1370,N_1309);
or U1548 (N_1548,N_1269,N_1345);
nor U1549 (N_1549,N_1367,N_1273);
and U1550 (N_1550,N_1215,N_1322);
nor U1551 (N_1551,N_1220,N_1200);
nand U1552 (N_1552,N_1214,N_1362);
and U1553 (N_1553,N_1372,N_1291);
and U1554 (N_1554,N_1358,N_1357);
and U1555 (N_1555,N_1236,N_1399);
or U1556 (N_1556,N_1370,N_1278);
or U1557 (N_1557,N_1351,N_1343);
and U1558 (N_1558,N_1364,N_1209);
and U1559 (N_1559,N_1245,N_1369);
or U1560 (N_1560,N_1300,N_1360);
nor U1561 (N_1561,N_1206,N_1240);
nor U1562 (N_1562,N_1299,N_1260);
nor U1563 (N_1563,N_1300,N_1337);
and U1564 (N_1564,N_1373,N_1364);
and U1565 (N_1565,N_1257,N_1310);
nor U1566 (N_1566,N_1215,N_1219);
or U1567 (N_1567,N_1236,N_1224);
and U1568 (N_1568,N_1244,N_1387);
or U1569 (N_1569,N_1336,N_1275);
nand U1570 (N_1570,N_1212,N_1389);
or U1571 (N_1571,N_1276,N_1316);
nor U1572 (N_1572,N_1201,N_1258);
nand U1573 (N_1573,N_1318,N_1316);
or U1574 (N_1574,N_1364,N_1374);
or U1575 (N_1575,N_1375,N_1212);
and U1576 (N_1576,N_1222,N_1314);
nor U1577 (N_1577,N_1336,N_1226);
nand U1578 (N_1578,N_1313,N_1326);
and U1579 (N_1579,N_1275,N_1212);
nand U1580 (N_1580,N_1282,N_1292);
and U1581 (N_1581,N_1201,N_1357);
or U1582 (N_1582,N_1280,N_1237);
nand U1583 (N_1583,N_1266,N_1349);
or U1584 (N_1584,N_1355,N_1389);
nand U1585 (N_1585,N_1277,N_1274);
or U1586 (N_1586,N_1211,N_1324);
and U1587 (N_1587,N_1246,N_1231);
and U1588 (N_1588,N_1372,N_1207);
nand U1589 (N_1589,N_1233,N_1205);
nand U1590 (N_1590,N_1240,N_1337);
xor U1591 (N_1591,N_1380,N_1249);
nor U1592 (N_1592,N_1390,N_1201);
and U1593 (N_1593,N_1217,N_1278);
nand U1594 (N_1594,N_1203,N_1214);
and U1595 (N_1595,N_1242,N_1259);
nand U1596 (N_1596,N_1279,N_1395);
and U1597 (N_1597,N_1268,N_1371);
and U1598 (N_1598,N_1380,N_1211);
nand U1599 (N_1599,N_1253,N_1248);
nand U1600 (N_1600,N_1572,N_1441);
nand U1601 (N_1601,N_1417,N_1416);
nor U1602 (N_1602,N_1539,N_1565);
nand U1603 (N_1603,N_1511,N_1433);
nor U1604 (N_1604,N_1567,N_1466);
and U1605 (N_1605,N_1506,N_1402);
nand U1606 (N_1606,N_1525,N_1429);
nand U1607 (N_1607,N_1467,N_1522);
and U1608 (N_1608,N_1596,N_1528);
and U1609 (N_1609,N_1403,N_1412);
nand U1610 (N_1610,N_1468,N_1534);
or U1611 (N_1611,N_1457,N_1447);
or U1612 (N_1612,N_1418,N_1589);
nor U1613 (N_1613,N_1570,N_1432);
xor U1614 (N_1614,N_1547,N_1507);
nand U1615 (N_1615,N_1569,N_1576);
nor U1616 (N_1616,N_1553,N_1439);
or U1617 (N_1617,N_1427,N_1509);
and U1618 (N_1618,N_1410,N_1558);
or U1619 (N_1619,N_1471,N_1420);
or U1620 (N_1620,N_1422,N_1518);
and U1621 (N_1621,N_1544,N_1404);
nor U1622 (N_1622,N_1520,N_1446);
and U1623 (N_1623,N_1533,N_1411);
or U1624 (N_1624,N_1409,N_1462);
nor U1625 (N_1625,N_1542,N_1571);
and U1626 (N_1626,N_1414,N_1495);
nand U1627 (N_1627,N_1543,N_1426);
nand U1628 (N_1628,N_1578,N_1405);
nand U1629 (N_1629,N_1541,N_1434);
nor U1630 (N_1630,N_1524,N_1552);
nand U1631 (N_1631,N_1440,N_1537);
nor U1632 (N_1632,N_1475,N_1566);
or U1633 (N_1633,N_1563,N_1500);
or U1634 (N_1634,N_1555,N_1483);
and U1635 (N_1635,N_1595,N_1470);
or U1636 (N_1636,N_1477,N_1556);
and U1637 (N_1637,N_1549,N_1406);
nor U1638 (N_1638,N_1592,N_1591);
nand U1639 (N_1639,N_1562,N_1488);
nand U1640 (N_1640,N_1517,N_1529);
or U1641 (N_1641,N_1564,N_1586);
xor U1642 (N_1642,N_1512,N_1492);
nand U1643 (N_1643,N_1516,N_1487);
nor U1644 (N_1644,N_1455,N_1550);
or U1645 (N_1645,N_1400,N_1575);
or U1646 (N_1646,N_1526,N_1536);
or U1647 (N_1647,N_1430,N_1450);
or U1648 (N_1648,N_1415,N_1599);
nand U1649 (N_1649,N_1590,N_1453);
nand U1650 (N_1650,N_1535,N_1448);
nand U1651 (N_1651,N_1435,N_1421);
or U1652 (N_1652,N_1597,N_1478);
nand U1653 (N_1653,N_1489,N_1408);
and U1654 (N_1654,N_1557,N_1501);
nor U1655 (N_1655,N_1491,N_1463);
or U1656 (N_1656,N_1551,N_1548);
nor U1657 (N_1657,N_1493,N_1481);
nor U1658 (N_1658,N_1513,N_1454);
or U1659 (N_1659,N_1469,N_1532);
xor U1660 (N_1660,N_1464,N_1581);
and U1661 (N_1661,N_1425,N_1498);
nor U1662 (N_1662,N_1484,N_1444);
and U1663 (N_1663,N_1527,N_1401);
and U1664 (N_1664,N_1504,N_1583);
nand U1665 (N_1665,N_1458,N_1428);
or U1666 (N_1666,N_1456,N_1442);
or U1667 (N_1667,N_1445,N_1554);
and U1668 (N_1668,N_1560,N_1459);
nor U1669 (N_1669,N_1505,N_1582);
nand U1670 (N_1670,N_1476,N_1460);
and U1671 (N_1671,N_1587,N_1502);
and U1672 (N_1672,N_1574,N_1530);
and U1673 (N_1673,N_1490,N_1423);
or U1674 (N_1674,N_1531,N_1443);
and U1675 (N_1675,N_1474,N_1485);
nand U1676 (N_1676,N_1438,N_1479);
nor U1677 (N_1677,N_1514,N_1436);
nand U1678 (N_1678,N_1449,N_1573);
nand U1679 (N_1679,N_1584,N_1451);
and U1680 (N_1680,N_1546,N_1496);
or U1681 (N_1681,N_1521,N_1424);
or U1682 (N_1682,N_1568,N_1579);
nor U1683 (N_1683,N_1494,N_1497);
nand U1684 (N_1684,N_1515,N_1503);
or U1685 (N_1685,N_1419,N_1561);
nand U1686 (N_1686,N_1510,N_1545);
and U1687 (N_1687,N_1480,N_1598);
nor U1688 (N_1688,N_1486,N_1594);
nor U1689 (N_1689,N_1538,N_1585);
or U1690 (N_1690,N_1523,N_1472);
nand U1691 (N_1691,N_1580,N_1593);
and U1692 (N_1692,N_1588,N_1461);
or U1693 (N_1693,N_1540,N_1431);
or U1694 (N_1694,N_1577,N_1452);
xor U1695 (N_1695,N_1508,N_1559);
xor U1696 (N_1696,N_1482,N_1473);
nor U1697 (N_1697,N_1413,N_1437);
nor U1698 (N_1698,N_1499,N_1465);
xnor U1699 (N_1699,N_1407,N_1519);
and U1700 (N_1700,N_1564,N_1421);
and U1701 (N_1701,N_1500,N_1507);
and U1702 (N_1702,N_1568,N_1451);
and U1703 (N_1703,N_1457,N_1487);
nor U1704 (N_1704,N_1475,N_1452);
and U1705 (N_1705,N_1448,N_1558);
or U1706 (N_1706,N_1501,N_1461);
xnor U1707 (N_1707,N_1565,N_1531);
and U1708 (N_1708,N_1557,N_1430);
nor U1709 (N_1709,N_1573,N_1534);
and U1710 (N_1710,N_1451,N_1509);
nand U1711 (N_1711,N_1445,N_1407);
nor U1712 (N_1712,N_1512,N_1482);
and U1713 (N_1713,N_1418,N_1541);
or U1714 (N_1714,N_1497,N_1557);
and U1715 (N_1715,N_1545,N_1425);
or U1716 (N_1716,N_1403,N_1404);
nor U1717 (N_1717,N_1478,N_1554);
nand U1718 (N_1718,N_1492,N_1474);
xnor U1719 (N_1719,N_1409,N_1516);
xor U1720 (N_1720,N_1457,N_1406);
and U1721 (N_1721,N_1502,N_1544);
or U1722 (N_1722,N_1457,N_1503);
nor U1723 (N_1723,N_1506,N_1403);
nand U1724 (N_1724,N_1460,N_1543);
or U1725 (N_1725,N_1582,N_1428);
nor U1726 (N_1726,N_1476,N_1549);
nor U1727 (N_1727,N_1407,N_1593);
nand U1728 (N_1728,N_1502,N_1503);
nand U1729 (N_1729,N_1567,N_1599);
xnor U1730 (N_1730,N_1527,N_1480);
nand U1731 (N_1731,N_1559,N_1400);
nand U1732 (N_1732,N_1429,N_1508);
or U1733 (N_1733,N_1491,N_1420);
or U1734 (N_1734,N_1531,N_1490);
nand U1735 (N_1735,N_1451,N_1540);
nor U1736 (N_1736,N_1441,N_1536);
and U1737 (N_1737,N_1463,N_1485);
nand U1738 (N_1738,N_1468,N_1511);
nor U1739 (N_1739,N_1467,N_1551);
nor U1740 (N_1740,N_1406,N_1546);
xor U1741 (N_1741,N_1550,N_1515);
nand U1742 (N_1742,N_1411,N_1584);
and U1743 (N_1743,N_1505,N_1448);
or U1744 (N_1744,N_1444,N_1424);
and U1745 (N_1745,N_1463,N_1456);
and U1746 (N_1746,N_1531,N_1510);
nor U1747 (N_1747,N_1484,N_1579);
or U1748 (N_1748,N_1458,N_1567);
nand U1749 (N_1749,N_1584,N_1514);
or U1750 (N_1750,N_1565,N_1593);
nor U1751 (N_1751,N_1534,N_1574);
nand U1752 (N_1752,N_1582,N_1437);
nand U1753 (N_1753,N_1438,N_1451);
and U1754 (N_1754,N_1487,N_1545);
or U1755 (N_1755,N_1407,N_1500);
and U1756 (N_1756,N_1451,N_1548);
nand U1757 (N_1757,N_1513,N_1482);
or U1758 (N_1758,N_1400,N_1508);
nand U1759 (N_1759,N_1439,N_1552);
nand U1760 (N_1760,N_1481,N_1592);
and U1761 (N_1761,N_1598,N_1534);
nor U1762 (N_1762,N_1518,N_1568);
or U1763 (N_1763,N_1578,N_1556);
or U1764 (N_1764,N_1577,N_1426);
or U1765 (N_1765,N_1537,N_1471);
nor U1766 (N_1766,N_1513,N_1410);
nor U1767 (N_1767,N_1594,N_1473);
nand U1768 (N_1768,N_1550,N_1591);
or U1769 (N_1769,N_1463,N_1499);
nand U1770 (N_1770,N_1403,N_1400);
and U1771 (N_1771,N_1560,N_1558);
or U1772 (N_1772,N_1440,N_1480);
and U1773 (N_1773,N_1488,N_1586);
nor U1774 (N_1774,N_1453,N_1514);
or U1775 (N_1775,N_1452,N_1513);
and U1776 (N_1776,N_1555,N_1549);
nand U1777 (N_1777,N_1530,N_1498);
nand U1778 (N_1778,N_1457,N_1542);
nand U1779 (N_1779,N_1466,N_1533);
nor U1780 (N_1780,N_1540,N_1448);
nor U1781 (N_1781,N_1549,N_1467);
nor U1782 (N_1782,N_1579,N_1425);
nor U1783 (N_1783,N_1421,N_1598);
nand U1784 (N_1784,N_1443,N_1595);
or U1785 (N_1785,N_1470,N_1534);
nand U1786 (N_1786,N_1472,N_1539);
nor U1787 (N_1787,N_1484,N_1539);
and U1788 (N_1788,N_1565,N_1577);
and U1789 (N_1789,N_1449,N_1434);
and U1790 (N_1790,N_1451,N_1466);
and U1791 (N_1791,N_1598,N_1415);
or U1792 (N_1792,N_1535,N_1425);
and U1793 (N_1793,N_1520,N_1529);
or U1794 (N_1794,N_1574,N_1461);
or U1795 (N_1795,N_1562,N_1425);
nor U1796 (N_1796,N_1594,N_1495);
and U1797 (N_1797,N_1503,N_1415);
xnor U1798 (N_1798,N_1508,N_1560);
or U1799 (N_1799,N_1445,N_1491);
and U1800 (N_1800,N_1746,N_1733);
and U1801 (N_1801,N_1796,N_1783);
nand U1802 (N_1802,N_1643,N_1690);
nand U1803 (N_1803,N_1611,N_1658);
or U1804 (N_1804,N_1628,N_1730);
and U1805 (N_1805,N_1716,N_1788);
nand U1806 (N_1806,N_1747,N_1654);
nor U1807 (N_1807,N_1792,N_1770);
nor U1808 (N_1808,N_1629,N_1714);
and U1809 (N_1809,N_1739,N_1630);
nand U1810 (N_1810,N_1638,N_1648);
nor U1811 (N_1811,N_1639,N_1720);
xnor U1812 (N_1812,N_1793,N_1672);
and U1813 (N_1813,N_1734,N_1797);
nand U1814 (N_1814,N_1736,N_1708);
nand U1815 (N_1815,N_1606,N_1673);
xnor U1816 (N_1816,N_1735,N_1689);
or U1817 (N_1817,N_1795,N_1757);
nor U1818 (N_1818,N_1622,N_1728);
nand U1819 (N_1819,N_1702,N_1687);
or U1820 (N_1820,N_1646,N_1756);
or U1821 (N_1821,N_1692,N_1614);
and U1822 (N_1822,N_1670,N_1766);
or U1823 (N_1823,N_1647,N_1762);
xor U1824 (N_1824,N_1699,N_1613);
and U1825 (N_1825,N_1752,N_1683);
nand U1826 (N_1826,N_1680,N_1635);
nand U1827 (N_1827,N_1655,N_1659);
and U1828 (N_1828,N_1789,N_1765);
nor U1829 (N_1829,N_1755,N_1676);
nand U1830 (N_1830,N_1688,N_1607);
and U1831 (N_1831,N_1769,N_1706);
or U1832 (N_1832,N_1603,N_1604);
or U1833 (N_1833,N_1740,N_1693);
or U1834 (N_1834,N_1799,N_1612);
nand U1835 (N_1835,N_1753,N_1675);
or U1836 (N_1836,N_1704,N_1634);
nand U1837 (N_1837,N_1653,N_1618);
nor U1838 (N_1838,N_1656,N_1600);
nand U1839 (N_1839,N_1621,N_1785);
and U1840 (N_1840,N_1726,N_1652);
or U1841 (N_1841,N_1678,N_1758);
nor U1842 (N_1842,N_1731,N_1729);
nor U1843 (N_1843,N_1778,N_1760);
and U1844 (N_1844,N_1723,N_1691);
nand U1845 (N_1845,N_1751,N_1636);
and U1846 (N_1846,N_1772,N_1617);
or U1847 (N_1847,N_1657,N_1707);
and U1848 (N_1848,N_1696,N_1645);
or U1849 (N_1849,N_1697,N_1698);
and U1850 (N_1850,N_1665,N_1668);
xnor U1851 (N_1851,N_1743,N_1794);
nand U1852 (N_1852,N_1651,N_1623);
or U1853 (N_1853,N_1694,N_1798);
nand U1854 (N_1854,N_1786,N_1649);
nor U1855 (N_1855,N_1767,N_1724);
nor U1856 (N_1856,N_1650,N_1715);
or U1857 (N_1857,N_1749,N_1667);
xnor U1858 (N_1858,N_1709,N_1602);
and U1859 (N_1859,N_1664,N_1713);
nor U1860 (N_1860,N_1776,N_1608);
xnor U1861 (N_1861,N_1782,N_1609);
nand U1862 (N_1862,N_1632,N_1601);
xnor U1863 (N_1863,N_1679,N_1727);
or U1864 (N_1864,N_1779,N_1784);
or U1865 (N_1865,N_1711,N_1775);
nand U1866 (N_1866,N_1700,N_1761);
or U1867 (N_1867,N_1764,N_1748);
nor U1868 (N_1868,N_1620,N_1663);
nand U1869 (N_1869,N_1781,N_1666);
nor U1870 (N_1870,N_1717,N_1791);
or U1871 (N_1871,N_1644,N_1725);
and U1872 (N_1872,N_1624,N_1610);
nand U1873 (N_1873,N_1669,N_1732);
nor U1874 (N_1874,N_1615,N_1637);
or U1875 (N_1875,N_1774,N_1684);
nand U1876 (N_1876,N_1641,N_1737);
nor U1877 (N_1877,N_1619,N_1777);
nand U1878 (N_1878,N_1759,N_1744);
and U1879 (N_1879,N_1662,N_1640);
and U1880 (N_1880,N_1677,N_1627);
nor U1881 (N_1881,N_1721,N_1642);
nor U1882 (N_1882,N_1633,N_1754);
and U1883 (N_1883,N_1703,N_1685);
nor U1884 (N_1884,N_1741,N_1616);
and U1885 (N_1885,N_1719,N_1631);
nand U1886 (N_1886,N_1718,N_1661);
or U1887 (N_1887,N_1773,N_1674);
xnor U1888 (N_1888,N_1710,N_1722);
and U1889 (N_1889,N_1780,N_1742);
nor U1890 (N_1890,N_1625,N_1681);
and U1891 (N_1891,N_1745,N_1671);
or U1892 (N_1892,N_1605,N_1771);
nor U1893 (N_1893,N_1738,N_1695);
nor U1894 (N_1894,N_1682,N_1701);
nand U1895 (N_1895,N_1712,N_1790);
and U1896 (N_1896,N_1626,N_1763);
or U1897 (N_1897,N_1750,N_1787);
nor U1898 (N_1898,N_1686,N_1705);
nor U1899 (N_1899,N_1768,N_1660);
or U1900 (N_1900,N_1759,N_1721);
nand U1901 (N_1901,N_1667,N_1601);
nand U1902 (N_1902,N_1672,N_1754);
or U1903 (N_1903,N_1622,N_1684);
and U1904 (N_1904,N_1654,N_1755);
nor U1905 (N_1905,N_1679,N_1693);
or U1906 (N_1906,N_1770,N_1665);
nand U1907 (N_1907,N_1736,N_1758);
nor U1908 (N_1908,N_1768,N_1690);
nor U1909 (N_1909,N_1615,N_1661);
and U1910 (N_1910,N_1637,N_1642);
nand U1911 (N_1911,N_1729,N_1741);
nand U1912 (N_1912,N_1748,N_1727);
and U1913 (N_1913,N_1631,N_1729);
nor U1914 (N_1914,N_1757,N_1712);
nor U1915 (N_1915,N_1738,N_1656);
nor U1916 (N_1916,N_1773,N_1634);
nand U1917 (N_1917,N_1704,N_1600);
nor U1918 (N_1918,N_1632,N_1759);
nand U1919 (N_1919,N_1742,N_1743);
and U1920 (N_1920,N_1715,N_1756);
or U1921 (N_1921,N_1688,N_1730);
and U1922 (N_1922,N_1626,N_1682);
nand U1923 (N_1923,N_1698,N_1655);
nand U1924 (N_1924,N_1784,N_1689);
nand U1925 (N_1925,N_1785,N_1602);
or U1926 (N_1926,N_1691,N_1664);
and U1927 (N_1927,N_1696,N_1653);
or U1928 (N_1928,N_1726,N_1642);
nor U1929 (N_1929,N_1720,N_1657);
or U1930 (N_1930,N_1616,N_1717);
or U1931 (N_1931,N_1774,N_1636);
nand U1932 (N_1932,N_1771,N_1672);
and U1933 (N_1933,N_1752,N_1629);
nor U1934 (N_1934,N_1768,N_1711);
nor U1935 (N_1935,N_1694,N_1790);
nand U1936 (N_1936,N_1763,N_1724);
or U1937 (N_1937,N_1649,N_1617);
or U1938 (N_1938,N_1600,N_1601);
nor U1939 (N_1939,N_1700,N_1684);
nand U1940 (N_1940,N_1604,N_1624);
nor U1941 (N_1941,N_1606,N_1626);
and U1942 (N_1942,N_1731,N_1774);
and U1943 (N_1943,N_1698,N_1648);
and U1944 (N_1944,N_1694,N_1701);
and U1945 (N_1945,N_1739,N_1728);
or U1946 (N_1946,N_1707,N_1785);
or U1947 (N_1947,N_1772,N_1622);
nor U1948 (N_1948,N_1762,N_1767);
and U1949 (N_1949,N_1623,N_1758);
or U1950 (N_1950,N_1721,N_1640);
and U1951 (N_1951,N_1764,N_1738);
nor U1952 (N_1952,N_1737,N_1708);
and U1953 (N_1953,N_1699,N_1662);
nand U1954 (N_1954,N_1767,N_1634);
nand U1955 (N_1955,N_1606,N_1654);
nand U1956 (N_1956,N_1668,N_1659);
nor U1957 (N_1957,N_1681,N_1612);
nor U1958 (N_1958,N_1768,N_1703);
nor U1959 (N_1959,N_1658,N_1644);
or U1960 (N_1960,N_1749,N_1788);
nor U1961 (N_1961,N_1680,N_1762);
nand U1962 (N_1962,N_1769,N_1606);
nor U1963 (N_1963,N_1667,N_1615);
nor U1964 (N_1964,N_1693,N_1694);
and U1965 (N_1965,N_1665,N_1714);
nor U1966 (N_1966,N_1631,N_1716);
or U1967 (N_1967,N_1695,N_1663);
nand U1968 (N_1968,N_1775,N_1604);
nand U1969 (N_1969,N_1787,N_1772);
nor U1970 (N_1970,N_1791,N_1774);
xnor U1971 (N_1971,N_1700,N_1664);
or U1972 (N_1972,N_1785,N_1653);
or U1973 (N_1973,N_1617,N_1681);
and U1974 (N_1974,N_1670,N_1743);
or U1975 (N_1975,N_1606,N_1748);
or U1976 (N_1976,N_1716,N_1609);
nand U1977 (N_1977,N_1745,N_1740);
nand U1978 (N_1978,N_1630,N_1772);
nand U1979 (N_1979,N_1766,N_1651);
and U1980 (N_1980,N_1665,N_1721);
nor U1981 (N_1981,N_1738,N_1798);
nor U1982 (N_1982,N_1645,N_1734);
nor U1983 (N_1983,N_1738,N_1611);
and U1984 (N_1984,N_1717,N_1665);
nor U1985 (N_1985,N_1753,N_1654);
nor U1986 (N_1986,N_1753,N_1727);
nor U1987 (N_1987,N_1714,N_1619);
nor U1988 (N_1988,N_1796,N_1789);
and U1989 (N_1989,N_1699,N_1770);
nor U1990 (N_1990,N_1643,N_1677);
nor U1991 (N_1991,N_1687,N_1686);
xnor U1992 (N_1992,N_1761,N_1631);
and U1993 (N_1993,N_1726,N_1788);
and U1994 (N_1994,N_1684,N_1747);
nor U1995 (N_1995,N_1775,N_1653);
and U1996 (N_1996,N_1745,N_1607);
nand U1997 (N_1997,N_1609,N_1631);
nand U1998 (N_1998,N_1614,N_1777);
or U1999 (N_1999,N_1667,N_1727);
nand U2000 (N_2000,N_1844,N_1828);
nor U2001 (N_2001,N_1882,N_1863);
and U2002 (N_2002,N_1916,N_1905);
and U2003 (N_2003,N_1912,N_1881);
nand U2004 (N_2004,N_1996,N_1929);
nor U2005 (N_2005,N_1928,N_1953);
or U2006 (N_2006,N_1981,N_1920);
xor U2007 (N_2007,N_1966,N_1873);
or U2008 (N_2008,N_1838,N_1821);
or U2009 (N_2009,N_1994,N_1807);
nor U2010 (N_2010,N_1813,N_1880);
and U2011 (N_2011,N_1803,N_1919);
and U2012 (N_2012,N_1884,N_1924);
or U2013 (N_2013,N_1876,N_1904);
or U2014 (N_2014,N_1941,N_1978);
xnor U2015 (N_2015,N_1982,N_1959);
nor U2016 (N_2016,N_1865,N_1859);
nand U2017 (N_2017,N_1954,N_1870);
nor U2018 (N_2018,N_1974,N_1977);
and U2019 (N_2019,N_1906,N_1985);
nor U2020 (N_2020,N_1841,N_1915);
or U2021 (N_2021,N_1948,N_1900);
nand U2022 (N_2022,N_1864,N_1816);
nor U2023 (N_2023,N_1814,N_1903);
and U2024 (N_2024,N_1979,N_1855);
nand U2025 (N_2025,N_1914,N_1856);
and U2026 (N_2026,N_1877,N_1949);
or U2027 (N_2027,N_1832,N_1888);
or U2028 (N_2028,N_1874,N_1925);
or U2029 (N_2029,N_1893,N_1883);
or U2030 (N_2030,N_1896,N_1890);
nor U2031 (N_2031,N_1836,N_1886);
and U2032 (N_2032,N_1899,N_1895);
nand U2033 (N_2033,N_1802,N_1940);
or U2034 (N_2034,N_1871,N_1848);
and U2035 (N_2035,N_1989,N_1971);
or U2036 (N_2036,N_1812,N_1818);
xnor U2037 (N_2037,N_1851,N_1969);
and U2038 (N_2038,N_1967,N_1849);
and U2039 (N_2039,N_1897,N_1885);
nor U2040 (N_2040,N_1972,N_1853);
and U2041 (N_2041,N_1957,N_1991);
nand U2042 (N_2042,N_1943,N_1858);
nand U2043 (N_2043,N_1922,N_1847);
xor U2044 (N_2044,N_1857,N_1962);
or U2045 (N_2045,N_1990,N_1800);
nand U2046 (N_2046,N_1805,N_1843);
or U2047 (N_2047,N_1937,N_1921);
nor U2048 (N_2048,N_1997,N_1879);
nand U2049 (N_2049,N_1842,N_1926);
xor U2050 (N_2050,N_1917,N_1965);
or U2051 (N_2051,N_1998,N_1891);
nor U2052 (N_2052,N_1932,N_1930);
nor U2053 (N_2053,N_1983,N_1834);
and U2054 (N_2054,N_1939,N_1823);
nand U2055 (N_2055,N_1833,N_1898);
nand U2056 (N_2056,N_1936,N_1866);
or U2057 (N_2057,N_1801,N_1992);
nor U2058 (N_2058,N_1980,N_1935);
or U2059 (N_2059,N_1889,N_1942);
nand U2060 (N_2060,N_1923,N_1826);
nor U2061 (N_2061,N_1934,N_1809);
and U2062 (N_2062,N_1909,N_1976);
and U2063 (N_2063,N_1835,N_1867);
or U2064 (N_2064,N_1846,N_1845);
or U2065 (N_2065,N_1829,N_1840);
xnor U2066 (N_2066,N_1830,N_1810);
or U2067 (N_2067,N_1944,N_1975);
nor U2068 (N_2068,N_1875,N_1984);
nand U2069 (N_2069,N_1824,N_1894);
or U2070 (N_2070,N_1815,N_1952);
or U2071 (N_2071,N_1958,N_1987);
nand U2072 (N_2072,N_1804,N_1933);
nand U2073 (N_2073,N_1970,N_1938);
and U2074 (N_2074,N_1973,N_1999);
and U2075 (N_2075,N_1995,N_1839);
nand U2076 (N_2076,N_1817,N_1945);
and U2077 (N_2077,N_1901,N_1902);
nor U2078 (N_2078,N_1950,N_1887);
and U2079 (N_2079,N_1908,N_1872);
or U2080 (N_2080,N_1951,N_1811);
nor U2081 (N_2081,N_1852,N_1911);
or U2082 (N_2082,N_1993,N_1907);
and U2083 (N_2083,N_1956,N_1827);
or U2084 (N_2084,N_1955,N_1913);
nand U2085 (N_2085,N_1850,N_1862);
nand U2086 (N_2086,N_1819,N_1960);
nand U2087 (N_2087,N_1860,N_1837);
or U2088 (N_2088,N_1931,N_1927);
and U2089 (N_2089,N_1918,N_1964);
nand U2090 (N_2090,N_1825,N_1986);
nand U2091 (N_2091,N_1988,N_1946);
or U2092 (N_2092,N_1910,N_1868);
nor U2093 (N_2093,N_1854,N_1892);
nor U2094 (N_2094,N_1820,N_1861);
nand U2095 (N_2095,N_1961,N_1808);
xnor U2096 (N_2096,N_1968,N_1963);
and U2097 (N_2097,N_1869,N_1806);
or U2098 (N_2098,N_1822,N_1947);
nand U2099 (N_2099,N_1878,N_1831);
and U2100 (N_2100,N_1803,N_1954);
nand U2101 (N_2101,N_1998,N_1991);
nand U2102 (N_2102,N_1907,N_1806);
and U2103 (N_2103,N_1869,N_1997);
nor U2104 (N_2104,N_1867,N_1984);
or U2105 (N_2105,N_1829,N_1975);
nand U2106 (N_2106,N_1932,N_1964);
nor U2107 (N_2107,N_1812,N_1898);
nor U2108 (N_2108,N_1850,N_1889);
nand U2109 (N_2109,N_1917,N_1972);
and U2110 (N_2110,N_1981,N_1934);
or U2111 (N_2111,N_1805,N_1837);
and U2112 (N_2112,N_1830,N_1925);
and U2113 (N_2113,N_1800,N_1855);
nand U2114 (N_2114,N_1810,N_1893);
nor U2115 (N_2115,N_1907,N_1821);
and U2116 (N_2116,N_1979,N_1970);
and U2117 (N_2117,N_1980,N_1846);
or U2118 (N_2118,N_1866,N_1880);
nand U2119 (N_2119,N_1898,N_1991);
and U2120 (N_2120,N_1991,N_1848);
nand U2121 (N_2121,N_1873,N_1820);
nand U2122 (N_2122,N_1917,N_1884);
nor U2123 (N_2123,N_1855,N_1871);
and U2124 (N_2124,N_1996,N_1973);
nor U2125 (N_2125,N_1817,N_1814);
nand U2126 (N_2126,N_1840,N_1970);
and U2127 (N_2127,N_1922,N_1848);
xnor U2128 (N_2128,N_1839,N_1810);
or U2129 (N_2129,N_1871,N_1957);
or U2130 (N_2130,N_1973,N_1847);
nor U2131 (N_2131,N_1849,N_1836);
or U2132 (N_2132,N_1979,N_1934);
or U2133 (N_2133,N_1870,N_1841);
nor U2134 (N_2134,N_1830,N_1915);
nor U2135 (N_2135,N_1830,N_1860);
and U2136 (N_2136,N_1830,N_1919);
or U2137 (N_2137,N_1892,N_1988);
nor U2138 (N_2138,N_1856,N_1891);
or U2139 (N_2139,N_1906,N_1922);
and U2140 (N_2140,N_1898,N_1986);
and U2141 (N_2141,N_1854,N_1802);
and U2142 (N_2142,N_1942,N_1951);
and U2143 (N_2143,N_1853,N_1950);
or U2144 (N_2144,N_1981,N_1895);
nand U2145 (N_2145,N_1943,N_1865);
or U2146 (N_2146,N_1826,N_1835);
and U2147 (N_2147,N_1938,N_1901);
nor U2148 (N_2148,N_1896,N_1831);
nor U2149 (N_2149,N_1965,N_1964);
or U2150 (N_2150,N_1804,N_1843);
nor U2151 (N_2151,N_1856,N_1870);
or U2152 (N_2152,N_1850,N_1952);
or U2153 (N_2153,N_1808,N_1905);
nor U2154 (N_2154,N_1954,N_1942);
nand U2155 (N_2155,N_1858,N_1819);
and U2156 (N_2156,N_1818,N_1887);
and U2157 (N_2157,N_1855,N_1833);
nor U2158 (N_2158,N_1800,N_1995);
or U2159 (N_2159,N_1843,N_1970);
or U2160 (N_2160,N_1889,N_1824);
nor U2161 (N_2161,N_1977,N_1834);
and U2162 (N_2162,N_1992,N_1990);
xnor U2163 (N_2163,N_1902,N_1847);
and U2164 (N_2164,N_1829,N_1934);
and U2165 (N_2165,N_1849,N_1937);
and U2166 (N_2166,N_1821,N_1893);
or U2167 (N_2167,N_1993,N_1894);
and U2168 (N_2168,N_1854,N_1924);
or U2169 (N_2169,N_1918,N_1947);
or U2170 (N_2170,N_1820,N_1838);
or U2171 (N_2171,N_1897,N_1886);
nand U2172 (N_2172,N_1825,N_1908);
nand U2173 (N_2173,N_1903,N_1936);
or U2174 (N_2174,N_1929,N_1912);
and U2175 (N_2175,N_1802,N_1818);
and U2176 (N_2176,N_1925,N_1890);
and U2177 (N_2177,N_1978,N_1896);
nor U2178 (N_2178,N_1849,N_1958);
or U2179 (N_2179,N_1814,N_1897);
xnor U2180 (N_2180,N_1988,N_1821);
and U2181 (N_2181,N_1956,N_1945);
or U2182 (N_2182,N_1825,N_1922);
or U2183 (N_2183,N_1886,N_1955);
or U2184 (N_2184,N_1926,N_1965);
or U2185 (N_2185,N_1802,N_1859);
nand U2186 (N_2186,N_1985,N_1980);
nand U2187 (N_2187,N_1812,N_1979);
nand U2188 (N_2188,N_1940,N_1939);
or U2189 (N_2189,N_1995,N_1862);
and U2190 (N_2190,N_1865,N_1860);
nor U2191 (N_2191,N_1975,N_1858);
nor U2192 (N_2192,N_1983,N_1914);
nand U2193 (N_2193,N_1859,N_1873);
nand U2194 (N_2194,N_1828,N_1826);
and U2195 (N_2195,N_1818,N_1829);
nand U2196 (N_2196,N_1902,N_1835);
nor U2197 (N_2197,N_1993,N_1990);
or U2198 (N_2198,N_1845,N_1918);
nand U2199 (N_2199,N_1954,N_1923);
or U2200 (N_2200,N_2125,N_2089);
nand U2201 (N_2201,N_2149,N_2197);
nand U2202 (N_2202,N_2077,N_2059);
nand U2203 (N_2203,N_2045,N_2140);
and U2204 (N_2204,N_2072,N_2136);
nor U2205 (N_2205,N_2175,N_2027);
and U2206 (N_2206,N_2085,N_2053);
and U2207 (N_2207,N_2123,N_2129);
nand U2208 (N_2208,N_2086,N_2084);
nor U2209 (N_2209,N_2018,N_2071);
nand U2210 (N_2210,N_2099,N_2025);
and U2211 (N_2211,N_2049,N_2141);
nor U2212 (N_2212,N_2035,N_2154);
xor U2213 (N_2213,N_2050,N_2198);
nor U2214 (N_2214,N_2160,N_2060);
and U2215 (N_2215,N_2032,N_2096);
nand U2216 (N_2216,N_2065,N_2196);
or U2217 (N_2217,N_2002,N_2168);
nor U2218 (N_2218,N_2006,N_2155);
nand U2219 (N_2219,N_2159,N_2177);
nor U2220 (N_2220,N_2088,N_2098);
nor U2221 (N_2221,N_2067,N_2000);
nand U2222 (N_2222,N_2031,N_2130);
nor U2223 (N_2223,N_2188,N_2063);
or U2224 (N_2224,N_2144,N_2162);
nor U2225 (N_2225,N_2132,N_2070);
xnor U2226 (N_2226,N_2126,N_2112);
and U2227 (N_2227,N_2157,N_2034);
nor U2228 (N_2228,N_2116,N_2021);
or U2229 (N_2229,N_2104,N_2172);
and U2230 (N_2230,N_2047,N_2183);
nand U2231 (N_2231,N_2164,N_2022);
and U2232 (N_2232,N_2080,N_2124);
or U2233 (N_2233,N_2093,N_2026);
and U2234 (N_2234,N_2173,N_2010);
nand U2235 (N_2235,N_2083,N_2058);
nor U2236 (N_2236,N_2171,N_2165);
nor U2237 (N_2237,N_2119,N_2014);
xor U2238 (N_2238,N_2192,N_2023);
nor U2239 (N_2239,N_2107,N_2127);
and U2240 (N_2240,N_2131,N_2174);
nand U2241 (N_2241,N_2040,N_2161);
or U2242 (N_2242,N_2087,N_2147);
and U2243 (N_2243,N_2015,N_2038);
or U2244 (N_2244,N_2078,N_2179);
or U2245 (N_2245,N_2054,N_2181);
and U2246 (N_2246,N_2122,N_2004);
nand U2247 (N_2247,N_2020,N_2128);
or U2248 (N_2248,N_2097,N_2139);
and U2249 (N_2249,N_2094,N_2069);
nor U2250 (N_2250,N_2052,N_2199);
xor U2251 (N_2251,N_2191,N_2037);
and U2252 (N_2252,N_2117,N_2103);
nand U2253 (N_2253,N_2146,N_2153);
and U2254 (N_2254,N_2143,N_2007);
or U2255 (N_2255,N_2092,N_2075);
nand U2256 (N_2256,N_2073,N_2145);
nand U2257 (N_2257,N_2019,N_2148);
and U2258 (N_2258,N_2042,N_2113);
or U2259 (N_2259,N_2182,N_2151);
and U2260 (N_2260,N_2044,N_2091);
nor U2261 (N_2261,N_2184,N_2135);
nand U2262 (N_2262,N_2194,N_2079);
and U2263 (N_2263,N_2013,N_2185);
and U2264 (N_2264,N_2115,N_2195);
nand U2265 (N_2265,N_2120,N_2189);
nor U2266 (N_2266,N_2005,N_2158);
or U2267 (N_2267,N_2012,N_2193);
and U2268 (N_2268,N_2064,N_2137);
nand U2269 (N_2269,N_2169,N_2066);
and U2270 (N_2270,N_2156,N_2024);
or U2271 (N_2271,N_2105,N_2142);
and U2272 (N_2272,N_2001,N_2150);
nor U2273 (N_2273,N_2055,N_2163);
and U2274 (N_2274,N_2102,N_2048);
nor U2275 (N_2275,N_2152,N_2003);
nand U2276 (N_2276,N_2109,N_2166);
or U2277 (N_2277,N_2187,N_2180);
or U2278 (N_2278,N_2029,N_2090);
or U2279 (N_2279,N_2108,N_2134);
nor U2280 (N_2280,N_2076,N_2008);
nor U2281 (N_2281,N_2056,N_2017);
nand U2282 (N_2282,N_2082,N_2095);
or U2283 (N_2283,N_2167,N_2114);
and U2284 (N_2284,N_2074,N_2190);
and U2285 (N_2285,N_2051,N_2133);
nand U2286 (N_2286,N_2033,N_2170);
and U2287 (N_2287,N_2101,N_2046);
nor U2288 (N_2288,N_2039,N_2068);
nand U2289 (N_2289,N_2062,N_2028);
and U2290 (N_2290,N_2100,N_2030);
and U2291 (N_2291,N_2118,N_2186);
or U2292 (N_2292,N_2106,N_2043);
nand U2293 (N_2293,N_2011,N_2041);
or U2294 (N_2294,N_2121,N_2061);
or U2295 (N_2295,N_2138,N_2057);
nand U2296 (N_2296,N_2110,N_2176);
nor U2297 (N_2297,N_2178,N_2016);
and U2298 (N_2298,N_2009,N_2111);
and U2299 (N_2299,N_2036,N_2081);
nand U2300 (N_2300,N_2018,N_2051);
and U2301 (N_2301,N_2184,N_2058);
nor U2302 (N_2302,N_2103,N_2189);
nor U2303 (N_2303,N_2084,N_2011);
nand U2304 (N_2304,N_2099,N_2170);
nand U2305 (N_2305,N_2193,N_2054);
and U2306 (N_2306,N_2078,N_2034);
nand U2307 (N_2307,N_2056,N_2011);
nor U2308 (N_2308,N_2130,N_2046);
nor U2309 (N_2309,N_2001,N_2037);
or U2310 (N_2310,N_2142,N_2095);
or U2311 (N_2311,N_2115,N_2019);
nor U2312 (N_2312,N_2028,N_2040);
nor U2313 (N_2313,N_2019,N_2103);
or U2314 (N_2314,N_2066,N_2157);
nand U2315 (N_2315,N_2086,N_2114);
nand U2316 (N_2316,N_2147,N_2118);
nand U2317 (N_2317,N_2157,N_2009);
or U2318 (N_2318,N_2003,N_2162);
xor U2319 (N_2319,N_2155,N_2017);
or U2320 (N_2320,N_2183,N_2016);
and U2321 (N_2321,N_2076,N_2049);
xor U2322 (N_2322,N_2140,N_2030);
and U2323 (N_2323,N_2095,N_2034);
or U2324 (N_2324,N_2107,N_2077);
or U2325 (N_2325,N_2054,N_2043);
or U2326 (N_2326,N_2070,N_2042);
nor U2327 (N_2327,N_2022,N_2146);
nand U2328 (N_2328,N_2139,N_2126);
and U2329 (N_2329,N_2062,N_2070);
and U2330 (N_2330,N_2087,N_2021);
nand U2331 (N_2331,N_2065,N_2011);
nand U2332 (N_2332,N_2052,N_2054);
nor U2333 (N_2333,N_2050,N_2055);
nand U2334 (N_2334,N_2101,N_2186);
and U2335 (N_2335,N_2111,N_2167);
and U2336 (N_2336,N_2163,N_2075);
nand U2337 (N_2337,N_2019,N_2165);
nor U2338 (N_2338,N_2039,N_2139);
nor U2339 (N_2339,N_2137,N_2143);
nand U2340 (N_2340,N_2025,N_2163);
nor U2341 (N_2341,N_2139,N_2178);
and U2342 (N_2342,N_2115,N_2163);
nand U2343 (N_2343,N_2168,N_2085);
and U2344 (N_2344,N_2159,N_2008);
and U2345 (N_2345,N_2033,N_2057);
nand U2346 (N_2346,N_2096,N_2066);
and U2347 (N_2347,N_2123,N_2070);
or U2348 (N_2348,N_2009,N_2171);
nor U2349 (N_2349,N_2069,N_2051);
nand U2350 (N_2350,N_2191,N_2070);
nand U2351 (N_2351,N_2123,N_2188);
nand U2352 (N_2352,N_2020,N_2032);
or U2353 (N_2353,N_2020,N_2010);
or U2354 (N_2354,N_2041,N_2118);
nor U2355 (N_2355,N_2197,N_2041);
and U2356 (N_2356,N_2076,N_2016);
xnor U2357 (N_2357,N_2183,N_2156);
nor U2358 (N_2358,N_2105,N_2048);
or U2359 (N_2359,N_2010,N_2158);
nor U2360 (N_2360,N_2182,N_2022);
nor U2361 (N_2361,N_2027,N_2006);
nand U2362 (N_2362,N_2107,N_2051);
nand U2363 (N_2363,N_2093,N_2001);
nor U2364 (N_2364,N_2180,N_2008);
nor U2365 (N_2365,N_2062,N_2138);
nand U2366 (N_2366,N_2148,N_2141);
and U2367 (N_2367,N_2123,N_2141);
or U2368 (N_2368,N_2019,N_2126);
or U2369 (N_2369,N_2032,N_2140);
xnor U2370 (N_2370,N_2082,N_2191);
or U2371 (N_2371,N_2013,N_2196);
xor U2372 (N_2372,N_2148,N_2009);
and U2373 (N_2373,N_2116,N_2003);
nand U2374 (N_2374,N_2084,N_2021);
xnor U2375 (N_2375,N_2016,N_2002);
nand U2376 (N_2376,N_2001,N_2041);
xor U2377 (N_2377,N_2068,N_2161);
or U2378 (N_2378,N_2165,N_2018);
and U2379 (N_2379,N_2021,N_2111);
or U2380 (N_2380,N_2143,N_2159);
nor U2381 (N_2381,N_2142,N_2072);
nand U2382 (N_2382,N_2123,N_2025);
nor U2383 (N_2383,N_2132,N_2079);
nor U2384 (N_2384,N_2081,N_2045);
nand U2385 (N_2385,N_2110,N_2075);
or U2386 (N_2386,N_2140,N_2028);
nor U2387 (N_2387,N_2124,N_2086);
and U2388 (N_2388,N_2041,N_2117);
and U2389 (N_2389,N_2038,N_2157);
nand U2390 (N_2390,N_2172,N_2096);
xnor U2391 (N_2391,N_2178,N_2008);
nand U2392 (N_2392,N_2197,N_2030);
xor U2393 (N_2393,N_2182,N_2049);
nor U2394 (N_2394,N_2148,N_2139);
or U2395 (N_2395,N_2041,N_2081);
or U2396 (N_2396,N_2190,N_2061);
nand U2397 (N_2397,N_2036,N_2132);
nand U2398 (N_2398,N_2088,N_2134);
and U2399 (N_2399,N_2151,N_2074);
nand U2400 (N_2400,N_2224,N_2328);
nor U2401 (N_2401,N_2389,N_2292);
nor U2402 (N_2402,N_2387,N_2322);
nor U2403 (N_2403,N_2234,N_2313);
and U2404 (N_2404,N_2399,N_2232);
nor U2405 (N_2405,N_2372,N_2369);
nand U2406 (N_2406,N_2339,N_2351);
nor U2407 (N_2407,N_2265,N_2381);
or U2408 (N_2408,N_2255,N_2310);
or U2409 (N_2409,N_2337,N_2312);
nand U2410 (N_2410,N_2227,N_2386);
and U2411 (N_2411,N_2223,N_2233);
nor U2412 (N_2412,N_2258,N_2338);
nand U2413 (N_2413,N_2382,N_2349);
nand U2414 (N_2414,N_2286,N_2331);
xnor U2415 (N_2415,N_2362,N_2316);
nor U2416 (N_2416,N_2323,N_2391);
and U2417 (N_2417,N_2345,N_2268);
nor U2418 (N_2418,N_2273,N_2275);
and U2419 (N_2419,N_2370,N_2200);
or U2420 (N_2420,N_2251,N_2226);
nor U2421 (N_2421,N_2211,N_2367);
nand U2422 (N_2422,N_2340,N_2267);
nor U2423 (N_2423,N_2347,N_2308);
and U2424 (N_2424,N_2332,N_2278);
or U2425 (N_2425,N_2284,N_2207);
xnor U2426 (N_2426,N_2301,N_2379);
nor U2427 (N_2427,N_2385,N_2212);
and U2428 (N_2428,N_2383,N_2368);
or U2429 (N_2429,N_2342,N_2361);
or U2430 (N_2430,N_2243,N_2204);
and U2431 (N_2431,N_2398,N_2335);
or U2432 (N_2432,N_2250,N_2376);
or U2433 (N_2433,N_2326,N_2246);
nand U2434 (N_2434,N_2282,N_2293);
and U2435 (N_2435,N_2249,N_2299);
nor U2436 (N_2436,N_2309,N_2291);
nand U2437 (N_2437,N_2203,N_2215);
or U2438 (N_2438,N_2244,N_2231);
nand U2439 (N_2439,N_2289,N_2311);
and U2440 (N_2440,N_2348,N_2393);
nand U2441 (N_2441,N_2355,N_2346);
nor U2442 (N_2442,N_2336,N_2294);
nor U2443 (N_2443,N_2240,N_2350);
or U2444 (N_2444,N_2271,N_2247);
and U2445 (N_2445,N_2274,N_2295);
or U2446 (N_2446,N_2205,N_2390);
or U2447 (N_2447,N_2356,N_2279);
nand U2448 (N_2448,N_2300,N_2360);
nand U2449 (N_2449,N_2334,N_2364);
and U2450 (N_2450,N_2283,N_2214);
and U2451 (N_2451,N_2314,N_2307);
or U2452 (N_2452,N_2290,N_2395);
xor U2453 (N_2453,N_2357,N_2230);
nor U2454 (N_2454,N_2218,N_2374);
and U2455 (N_2455,N_2353,N_2280);
nand U2456 (N_2456,N_2239,N_2330);
nor U2457 (N_2457,N_2354,N_2261);
nand U2458 (N_2458,N_2343,N_2321);
or U2459 (N_2459,N_2325,N_2394);
nand U2460 (N_2460,N_2285,N_2371);
or U2461 (N_2461,N_2298,N_2296);
nor U2462 (N_2462,N_2363,N_2373);
nor U2463 (N_2463,N_2315,N_2235);
and U2464 (N_2464,N_2222,N_2229);
nand U2465 (N_2465,N_2236,N_2306);
and U2466 (N_2466,N_2358,N_2397);
nand U2467 (N_2467,N_2329,N_2388);
nand U2468 (N_2468,N_2201,N_2257);
and U2469 (N_2469,N_2375,N_2396);
or U2470 (N_2470,N_2366,N_2209);
nand U2471 (N_2471,N_2262,N_2272);
nor U2472 (N_2472,N_2318,N_2287);
or U2473 (N_2473,N_2206,N_2263);
or U2474 (N_2474,N_2324,N_2210);
and U2475 (N_2475,N_2319,N_2320);
or U2476 (N_2476,N_2253,N_2392);
or U2477 (N_2477,N_2256,N_2359);
nand U2478 (N_2478,N_2352,N_2252);
nand U2479 (N_2479,N_2213,N_2377);
and U2480 (N_2480,N_2365,N_2266);
nand U2481 (N_2481,N_2259,N_2202);
or U2482 (N_2482,N_2333,N_2254);
and U2483 (N_2483,N_2216,N_2219);
nand U2484 (N_2484,N_2270,N_2237);
nand U2485 (N_2485,N_2277,N_2221);
nor U2486 (N_2486,N_2303,N_2304);
or U2487 (N_2487,N_2341,N_2269);
or U2488 (N_2488,N_2248,N_2344);
nor U2489 (N_2489,N_2208,N_2297);
or U2490 (N_2490,N_2238,N_2305);
and U2491 (N_2491,N_2317,N_2220);
nand U2492 (N_2492,N_2260,N_2228);
xor U2493 (N_2493,N_2378,N_2245);
nor U2494 (N_2494,N_2302,N_2276);
or U2495 (N_2495,N_2217,N_2281);
nor U2496 (N_2496,N_2327,N_2380);
or U2497 (N_2497,N_2241,N_2384);
and U2498 (N_2498,N_2264,N_2288);
and U2499 (N_2499,N_2242,N_2225);
nand U2500 (N_2500,N_2271,N_2360);
and U2501 (N_2501,N_2397,N_2391);
and U2502 (N_2502,N_2258,N_2283);
nand U2503 (N_2503,N_2280,N_2222);
or U2504 (N_2504,N_2308,N_2216);
or U2505 (N_2505,N_2301,N_2224);
and U2506 (N_2506,N_2307,N_2322);
or U2507 (N_2507,N_2266,N_2353);
nand U2508 (N_2508,N_2296,N_2287);
nand U2509 (N_2509,N_2206,N_2306);
nand U2510 (N_2510,N_2220,N_2207);
or U2511 (N_2511,N_2282,N_2280);
and U2512 (N_2512,N_2243,N_2242);
and U2513 (N_2513,N_2264,N_2240);
and U2514 (N_2514,N_2329,N_2231);
nor U2515 (N_2515,N_2236,N_2320);
nand U2516 (N_2516,N_2309,N_2288);
nand U2517 (N_2517,N_2284,N_2235);
and U2518 (N_2518,N_2291,N_2302);
nand U2519 (N_2519,N_2302,N_2374);
nor U2520 (N_2520,N_2271,N_2209);
or U2521 (N_2521,N_2357,N_2280);
nand U2522 (N_2522,N_2389,N_2371);
xnor U2523 (N_2523,N_2202,N_2218);
and U2524 (N_2524,N_2211,N_2284);
or U2525 (N_2525,N_2392,N_2246);
xor U2526 (N_2526,N_2386,N_2394);
or U2527 (N_2527,N_2245,N_2323);
nor U2528 (N_2528,N_2326,N_2267);
and U2529 (N_2529,N_2335,N_2290);
or U2530 (N_2530,N_2283,N_2322);
nand U2531 (N_2531,N_2237,N_2243);
and U2532 (N_2532,N_2256,N_2395);
nand U2533 (N_2533,N_2217,N_2227);
or U2534 (N_2534,N_2365,N_2220);
nand U2535 (N_2535,N_2255,N_2365);
nand U2536 (N_2536,N_2340,N_2241);
xor U2537 (N_2537,N_2302,N_2301);
or U2538 (N_2538,N_2306,N_2203);
and U2539 (N_2539,N_2376,N_2221);
or U2540 (N_2540,N_2358,N_2243);
nand U2541 (N_2541,N_2376,N_2281);
and U2542 (N_2542,N_2290,N_2329);
nor U2543 (N_2543,N_2228,N_2208);
or U2544 (N_2544,N_2267,N_2216);
nor U2545 (N_2545,N_2359,N_2220);
nand U2546 (N_2546,N_2361,N_2359);
and U2547 (N_2547,N_2376,N_2211);
nor U2548 (N_2548,N_2398,N_2281);
or U2549 (N_2549,N_2395,N_2327);
xnor U2550 (N_2550,N_2335,N_2382);
nor U2551 (N_2551,N_2266,N_2206);
nor U2552 (N_2552,N_2390,N_2310);
nor U2553 (N_2553,N_2265,N_2391);
and U2554 (N_2554,N_2283,N_2274);
and U2555 (N_2555,N_2326,N_2211);
nand U2556 (N_2556,N_2347,N_2387);
and U2557 (N_2557,N_2371,N_2272);
nor U2558 (N_2558,N_2393,N_2351);
nor U2559 (N_2559,N_2348,N_2343);
or U2560 (N_2560,N_2230,N_2337);
or U2561 (N_2561,N_2204,N_2237);
and U2562 (N_2562,N_2245,N_2381);
and U2563 (N_2563,N_2345,N_2269);
nand U2564 (N_2564,N_2366,N_2397);
or U2565 (N_2565,N_2280,N_2399);
nand U2566 (N_2566,N_2296,N_2304);
or U2567 (N_2567,N_2283,N_2260);
and U2568 (N_2568,N_2384,N_2202);
and U2569 (N_2569,N_2249,N_2238);
nand U2570 (N_2570,N_2265,N_2356);
nand U2571 (N_2571,N_2378,N_2385);
and U2572 (N_2572,N_2346,N_2324);
and U2573 (N_2573,N_2349,N_2316);
and U2574 (N_2574,N_2283,N_2327);
nor U2575 (N_2575,N_2213,N_2356);
nor U2576 (N_2576,N_2391,N_2217);
and U2577 (N_2577,N_2338,N_2210);
and U2578 (N_2578,N_2211,N_2257);
and U2579 (N_2579,N_2284,N_2264);
nor U2580 (N_2580,N_2257,N_2336);
and U2581 (N_2581,N_2278,N_2232);
nor U2582 (N_2582,N_2208,N_2248);
xor U2583 (N_2583,N_2304,N_2305);
or U2584 (N_2584,N_2312,N_2245);
or U2585 (N_2585,N_2242,N_2384);
nand U2586 (N_2586,N_2244,N_2328);
or U2587 (N_2587,N_2333,N_2300);
nand U2588 (N_2588,N_2241,N_2378);
or U2589 (N_2589,N_2315,N_2277);
and U2590 (N_2590,N_2312,N_2267);
xor U2591 (N_2591,N_2215,N_2244);
and U2592 (N_2592,N_2325,N_2355);
or U2593 (N_2593,N_2291,N_2268);
nand U2594 (N_2594,N_2332,N_2379);
nor U2595 (N_2595,N_2376,N_2362);
and U2596 (N_2596,N_2379,N_2398);
or U2597 (N_2597,N_2391,N_2272);
nor U2598 (N_2598,N_2279,N_2257);
nand U2599 (N_2599,N_2368,N_2253);
or U2600 (N_2600,N_2573,N_2560);
nand U2601 (N_2601,N_2456,N_2414);
nand U2602 (N_2602,N_2546,N_2450);
nand U2603 (N_2603,N_2502,N_2498);
nand U2604 (N_2604,N_2478,N_2572);
nand U2605 (N_2605,N_2599,N_2420);
or U2606 (N_2606,N_2593,N_2537);
nand U2607 (N_2607,N_2596,N_2513);
or U2608 (N_2608,N_2407,N_2511);
and U2609 (N_2609,N_2459,N_2532);
and U2610 (N_2610,N_2578,N_2512);
and U2611 (N_2611,N_2460,N_2433);
nand U2612 (N_2612,N_2439,N_2554);
and U2613 (N_2613,N_2449,N_2455);
and U2614 (N_2614,N_2542,N_2481);
or U2615 (N_2615,N_2592,N_2557);
nand U2616 (N_2616,N_2567,N_2504);
nand U2617 (N_2617,N_2571,N_2538);
or U2618 (N_2618,N_2473,N_2522);
nand U2619 (N_2619,N_2539,N_2448);
nor U2620 (N_2620,N_2496,N_2415);
and U2621 (N_2621,N_2462,N_2527);
nand U2622 (N_2622,N_2404,N_2427);
or U2623 (N_2623,N_2566,N_2470);
or U2624 (N_2624,N_2432,N_2417);
and U2625 (N_2625,N_2469,N_2597);
or U2626 (N_2626,N_2438,N_2519);
or U2627 (N_2627,N_2403,N_2493);
or U2628 (N_2628,N_2520,N_2463);
or U2629 (N_2629,N_2525,N_2485);
nor U2630 (N_2630,N_2594,N_2589);
and U2631 (N_2631,N_2416,N_2418);
or U2632 (N_2632,N_2558,N_2491);
nor U2633 (N_2633,N_2484,N_2428);
nor U2634 (N_2634,N_2552,N_2430);
or U2635 (N_2635,N_2521,N_2591);
nand U2636 (N_2636,N_2503,N_2454);
nand U2637 (N_2637,N_2501,N_2435);
nor U2638 (N_2638,N_2531,N_2547);
nor U2639 (N_2639,N_2561,N_2526);
nand U2640 (N_2640,N_2423,N_2541);
xor U2641 (N_2641,N_2411,N_2523);
or U2642 (N_2642,N_2426,N_2429);
or U2643 (N_2643,N_2564,N_2528);
and U2644 (N_2644,N_2515,N_2408);
nand U2645 (N_2645,N_2476,N_2495);
nor U2646 (N_2646,N_2577,N_2500);
and U2647 (N_2647,N_2490,N_2482);
and U2648 (N_2648,N_2505,N_2529);
nand U2649 (N_2649,N_2464,N_2590);
or U2650 (N_2650,N_2444,N_2436);
nand U2651 (N_2651,N_2486,N_2575);
nor U2652 (N_2652,N_2524,N_2556);
nor U2653 (N_2653,N_2517,N_2437);
and U2654 (N_2654,N_2583,N_2580);
nand U2655 (N_2655,N_2425,N_2570);
nand U2656 (N_2656,N_2559,N_2550);
or U2657 (N_2657,N_2534,N_2494);
and U2658 (N_2658,N_2412,N_2492);
nand U2659 (N_2659,N_2509,N_2434);
or U2660 (N_2660,N_2544,N_2488);
and U2661 (N_2661,N_2442,N_2598);
nand U2662 (N_2662,N_2543,N_2533);
nand U2663 (N_2663,N_2402,N_2409);
or U2664 (N_2664,N_2585,N_2555);
nand U2665 (N_2665,N_2458,N_2562);
nand U2666 (N_2666,N_2480,N_2474);
nand U2667 (N_2667,N_2540,N_2466);
nand U2668 (N_2668,N_2453,N_2467);
and U2669 (N_2669,N_2483,N_2406);
or U2670 (N_2670,N_2447,N_2400);
nand U2671 (N_2671,N_2584,N_2569);
nand U2672 (N_2672,N_2465,N_2440);
or U2673 (N_2673,N_2421,N_2587);
nor U2674 (N_2674,N_2545,N_2499);
xnor U2675 (N_2675,N_2468,N_2431);
and U2676 (N_2676,N_2497,N_2588);
xnor U2677 (N_2677,N_2401,N_2475);
nand U2678 (N_2678,N_2530,N_2451);
and U2679 (N_2679,N_2506,N_2446);
nor U2680 (N_2680,N_2574,N_2568);
nor U2681 (N_2681,N_2548,N_2452);
or U2682 (N_2682,N_2479,N_2507);
nand U2683 (N_2683,N_2445,N_2461);
or U2684 (N_2684,N_2422,N_2516);
nand U2685 (N_2685,N_2443,N_2457);
and U2686 (N_2686,N_2441,N_2581);
nor U2687 (N_2687,N_2510,N_2565);
nand U2688 (N_2688,N_2424,N_2595);
nand U2689 (N_2689,N_2487,N_2405);
nor U2690 (N_2690,N_2582,N_2586);
xnor U2691 (N_2691,N_2576,N_2413);
nand U2692 (N_2692,N_2471,N_2477);
nand U2693 (N_2693,N_2518,N_2472);
and U2694 (N_2694,N_2579,N_2563);
and U2695 (N_2695,N_2489,N_2514);
nor U2696 (N_2696,N_2508,N_2551);
nand U2697 (N_2697,N_2419,N_2536);
nand U2698 (N_2698,N_2535,N_2549);
and U2699 (N_2699,N_2553,N_2410);
or U2700 (N_2700,N_2579,N_2469);
and U2701 (N_2701,N_2423,N_2519);
and U2702 (N_2702,N_2541,N_2503);
or U2703 (N_2703,N_2505,N_2494);
nand U2704 (N_2704,N_2594,N_2423);
nor U2705 (N_2705,N_2491,N_2494);
and U2706 (N_2706,N_2517,N_2571);
nor U2707 (N_2707,N_2517,N_2576);
nor U2708 (N_2708,N_2547,N_2514);
nor U2709 (N_2709,N_2461,N_2591);
or U2710 (N_2710,N_2409,N_2504);
and U2711 (N_2711,N_2483,N_2449);
or U2712 (N_2712,N_2513,N_2422);
and U2713 (N_2713,N_2457,N_2547);
or U2714 (N_2714,N_2561,N_2508);
or U2715 (N_2715,N_2530,N_2433);
nor U2716 (N_2716,N_2550,N_2551);
or U2717 (N_2717,N_2403,N_2533);
and U2718 (N_2718,N_2454,N_2470);
or U2719 (N_2719,N_2483,N_2434);
nand U2720 (N_2720,N_2497,N_2514);
and U2721 (N_2721,N_2430,N_2572);
nand U2722 (N_2722,N_2559,N_2407);
nand U2723 (N_2723,N_2512,N_2546);
nand U2724 (N_2724,N_2529,N_2539);
or U2725 (N_2725,N_2462,N_2415);
or U2726 (N_2726,N_2503,N_2556);
nor U2727 (N_2727,N_2554,N_2432);
nor U2728 (N_2728,N_2507,N_2427);
and U2729 (N_2729,N_2489,N_2499);
nand U2730 (N_2730,N_2573,N_2552);
nor U2731 (N_2731,N_2531,N_2489);
and U2732 (N_2732,N_2551,N_2552);
nand U2733 (N_2733,N_2544,N_2491);
nand U2734 (N_2734,N_2559,N_2487);
and U2735 (N_2735,N_2423,N_2502);
and U2736 (N_2736,N_2591,N_2438);
or U2737 (N_2737,N_2510,N_2526);
nand U2738 (N_2738,N_2409,N_2429);
and U2739 (N_2739,N_2450,N_2589);
nor U2740 (N_2740,N_2550,N_2594);
and U2741 (N_2741,N_2563,N_2523);
or U2742 (N_2742,N_2420,N_2445);
nand U2743 (N_2743,N_2568,N_2424);
nor U2744 (N_2744,N_2404,N_2589);
nor U2745 (N_2745,N_2477,N_2585);
nand U2746 (N_2746,N_2508,N_2465);
and U2747 (N_2747,N_2430,N_2579);
and U2748 (N_2748,N_2523,N_2467);
xor U2749 (N_2749,N_2530,N_2571);
nand U2750 (N_2750,N_2489,N_2512);
or U2751 (N_2751,N_2541,N_2537);
nand U2752 (N_2752,N_2415,N_2598);
or U2753 (N_2753,N_2436,N_2582);
or U2754 (N_2754,N_2527,N_2536);
nor U2755 (N_2755,N_2485,N_2404);
or U2756 (N_2756,N_2525,N_2555);
and U2757 (N_2757,N_2423,N_2434);
nor U2758 (N_2758,N_2495,N_2453);
and U2759 (N_2759,N_2477,N_2543);
and U2760 (N_2760,N_2464,N_2559);
nor U2761 (N_2761,N_2553,N_2599);
or U2762 (N_2762,N_2498,N_2454);
or U2763 (N_2763,N_2509,N_2591);
nand U2764 (N_2764,N_2491,N_2573);
nor U2765 (N_2765,N_2502,N_2580);
or U2766 (N_2766,N_2445,N_2528);
or U2767 (N_2767,N_2511,N_2515);
nor U2768 (N_2768,N_2406,N_2584);
and U2769 (N_2769,N_2486,N_2542);
nor U2770 (N_2770,N_2522,N_2504);
nor U2771 (N_2771,N_2432,N_2552);
or U2772 (N_2772,N_2444,N_2531);
or U2773 (N_2773,N_2596,N_2550);
and U2774 (N_2774,N_2407,N_2578);
and U2775 (N_2775,N_2448,N_2496);
or U2776 (N_2776,N_2504,N_2437);
or U2777 (N_2777,N_2470,N_2424);
or U2778 (N_2778,N_2528,N_2567);
and U2779 (N_2779,N_2503,N_2555);
nor U2780 (N_2780,N_2524,N_2422);
nand U2781 (N_2781,N_2415,N_2580);
or U2782 (N_2782,N_2590,N_2548);
xnor U2783 (N_2783,N_2499,N_2524);
nand U2784 (N_2784,N_2504,N_2439);
nor U2785 (N_2785,N_2430,N_2422);
nand U2786 (N_2786,N_2522,N_2589);
or U2787 (N_2787,N_2499,N_2540);
or U2788 (N_2788,N_2555,N_2504);
and U2789 (N_2789,N_2573,N_2577);
or U2790 (N_2790,N_2513,N_2516);
nor U2791 (N_2791,N_2563,N_2434);
or U2792 (N_2792,N_2401,N_2594);
xnor U2793 (N_2793,N_2594,N_2435);
and U2794 (N_2794,N_2537,N_2455);
nor U2795 (N_2795,N_2544,N_2495);
nand U2796 (N_2796,N_2467,N_2598);
nand U2797 (N_2797,N_2518,N_2441);
and U2798 (N_2798,N_2426,N_2558);
or U2799 (N_2799,N_2572,N_2584);
nor U2800 (N_2800,N_2765,N_2776);
xor U2801 (N_2801,N_2748,N_2724);
nand U2802 (N_2802,N_2601,N_2628);
nand U2803 (N_2803,N_2751,N_2605);
nand U2804 (N_2804,N_2727,N_2718);
nand U2805 (N_2805,N_2784,N_2614);
or U2806 (N_2806,N_2721,N_2680);
nand U2807 (N_2807,N_2760,N_2633);
or U2808 (N_2808,N_2719,N_2720);
nor U2809 (N_2809,N_2637,N_2791);
nand U2810 (N_2810,N_2741,N_2612);
nor U2811 (N_2811,N_2665,N_2667);
and U2812 (N_2812,N_2725,N_2624);
and U2813 (N_2813,N_2795,N_2689);
or U2814 (N_2814,N_2656,N_2668);
or U2815 (N_2815,N_2622,N_2794);
or U2816 (N_2816,N_2644,N_2691);
nand U2817 (N_2817,N_2669,N_2723);
nor U2818 (N_2818,N_2742,N_2722);
and U2819 (N_2819,N_2702,N_2648);
nand U2820 (N_2820,N_2636,N_2639);
nor U2821 (N_2821,N_2693,N_2683);
nor U2822 (N_2822,N_2659,N_2615);
nand U2823 (N_2823,N_2651,N_2733);
nor U2824 (N_2824,N_2726,N_2707);
or U2825 (N_2825,N_2678,N_2793);
and U2826 (N_2826,N_2682,N_2746);
nand U2827 (N_2827,N_2641,N_2664);
nand U2828 (N_2828,N_2740,N_2697);
or U2829 (N_2829,N_2767,N_2688);
nor U2830 (N_2830,N_2757,N_2634);
and U2831 (N_2831,N_2700,N_2621);
and U2832 (N_2832,N_2695,N_2755);
or U2833 (N_2833,N_2786,N_2731);
nand U2834 (N_2834,N_2657,N_2705);
nor U2835 (N_2835,N_2763,N_2645);
nand U2836 (N_2836,N_2674,N_2745);
or U2837 (N_2837,N_2773,N_2609);
nand U2838 (N_2838,N_2796,N_2711);
nand U2839 (N_2839,N_2646,N_2654);
or U2840 (N_2840,N_2606,N_2635);
xnor U2841 (N_2841,N_2736,N_2632);
nand U2842 (N_2842,N_2714,N_2782);
and U2843 (N_2843,N_2788,N_2777);
and U2844 (N_2844,N_2687,N_2739);
or U2845 (N_2845,N_2709,N_2708);
nor U2846 (N_2846,N_2710,N_2647);
and U2847 (N_2847,N_2608,N_2677);
nand U2848 (N_2848,N_2670,N_2660);
nand U2849 (N_2849,N_2713,N_2630);
and U2850 (N_2850,N_2747,N_2610);
and U2851 (N_2851,N_2618,N_2643);
or U2852 (N_2852,N_2696,N_2712);
or U2853 (N_2853,N_2769,N_2735);
or U2854 (N_2854,N_2704,N_2640);
nor U2855 (N_2855,N_2698,N_2729);
or U2856 (N_2856,N_2662,N_2778);
nand U2857 (N_2857,N_2616,N_2602);
xnor U2858 (N_2858,N_2672,N_2715);
nand U2859 (N_2859,N_2686,N_2768);
or U2860 (N_2860,N_2797,N_2758);
nand U2861 (N_2861,N_2770,N_2781);
or U2862 (N_2862,N_2625,N_2658);
nand U2863 (N_2863,N_2734,N_2732);
or U2864 (N_2864,N_2642,N_2623);
xor U2865 (N_2865,N_2706,N_2716);
nand U2866 (N_2866,N_2701,N_2620);
or U2867 (N_2867,N_2761,N_2611);
or U2868 (N_2868,N_2603,N_2737);
or U2869 (N_2869,N_2750,N_2613);
nand U2870 (N_2870,N_2792,N_2787);
nor U2871 (N_2871,N_2617,N_2604);
or U2872 (N_2872,N_2774,N_2790);
or U2873 (N_2873,N_2749,N_2779);
nor U2874 (N_2874,N_2783,N_2679);
nor U2875 (N_2875,N_2743,N_2775);
or U2876 (N_2876,N_2692,N_2789);
or U2877 (N_2877,N_2728,N_2607);
nor U2878 (N_2878,N_2762,N_2753);
nor U2879 (N_2879,N_2744,N_2600);
nor U2880 (N_2880,N_2650,N_2652);
and U2881 (N_2881,N_2699,N_2785);
and U2882 (N_2882,N_2694,N_2681);
nor U2883 (N_2883,N_2631,N_2626);
and U2884 (N_2884,N_2663,N_2655);
nand U2885 (N_2885,N_2780,N_2685);
nor U2886 (N_2886,N_2684,N_2619);
nor U2887 (N_2887,N_2754,N_2772);
or U2888 (N_2888,N_2676,N_2730);
nand U2889 (N_2889,N_2690,N_2756);
or U2890 (N_2890,N_2766,N_2738);
or U2891 (N_2891,N_2771,N_2798);
and U2892 (N_2892,N_2764,N_2666);
or U2893 (N_2893,N_2638,N_2629);
nor U2894 (N_2894,N_2675,N_2752);
nand U2895 (N_2895,N_2649,N_2717);
and U2896 (N_2896,N_2653,N_2799);
nor U2897 (N_2897,N_2759,N_2671);
nor U2898 (N_2898,N_2627,N_2673);
nand U2899 (N_2899,N_2661,N_2703);
and U2900 (N_2900,N_2677,N_2737);
or U2901 (N_2901,N_2668,N_2662);
and U2902 (N_2902,N_2764,N_2789);
nor U2903 (N_2903,N_2734,N_2652);
and U2904 (N_2904,N_2752,N_2645);
nor U2905 (N_2905,N_2742,N_2601);
nand U2906 (N_2906,N_2729,N_2716);
and U2907 (N_2907,N_2700,N_2799);
nand U2908 (N_2908,N_2674,N_2654);
nand U2909 (N_2909,N_2786,N_2754);
and U2910 (N_2910,N_2601,N_2703);
nor U2911 (N_2911,N_2641,N_2706);
or U2912 (N_2912,N_2669,N_2741);
and U2913 (N_2913,N_2664,N_2700);
or U2914 (N_2914,N_2703,N_2786);
or U2915 (N_2915,N_2765,N_2768);
and U2916 (N_2916,N_2731,N_2666);
or U2917 (N_2917,N_2605,N_2756);
nor U2918 (N_2918,N_2684,N_2767);
or U2919 (N_2919,N_2781,N_2600);
nor U2920 (N_2920,N_2601,N_2680);
nand U2921 (N_2921,N_2687,N_2663);
and U2922 (N_2922,N_2693,N_2747);
nor U2923 (N_2923,N_2752,N_2720);
and U2924 (N_2924,N_2750,N_2642);
nand U2925 (N_2925,N_2782,N_2601);
nor U2926 (N_2926,N_2658,N_2708);
nor U2927 (N_2927,N_2743,N_2608);
nor U2928 (N_2928,N_2702,N_2750);
or U2929 (N_2929,N_2695,N_2606);
nor U2930 (N_2930,N_2765,N_2798);
nand U2931 (N_2931,N_2767,N_2781);
and U2932 (N_2932,N_2787,N_2749);
or U2933 (N_2933,N_2757,N_2775);
or U2934 (N_2934,N_2620,N_2623);
nor U2935 (N_2935,N_2671,N_2650);
and U2936 (N_2936,N_2790,N_2691);
nor U2937 (N_2937,N_2691,N_2768);
or U2938 (N_2938,N_2774,N_2745);
xor U2939 (N_2939,N_2782,N_2791);
or U2940 (N_2940,N_2679,N_2792);
nand U2941 (N_2941,N_2738,N_2608);
or U2942 (N_2942,N_2759,N_2792);
or U2943 (N_2943,N_2692,N_2780);
and U2944 (N_2944,N_2698,N_2697);
nand U2945 (N_2945,N_2665,N_2669);
nor U2946 (N_2946,N_2697,N_2781);
and U2947 (N_2947,N_2667,N_2728);
nand U2948 (N_2948,N_2718,N_2781);
or U2949 (N_2949,N_2604,N_2752);
nand U2950 (N_2950,N_2723,N_2774);
or U2951 (N_2951,N_2620,N_2739);
nand U2952 (N_2952,N_2605,N_2735);
or U2953 (N_2953,N_2743,N_2605);
nand U2954 (N_2954,N_2624,N_2715);
xor U2955 (N_2955,N_2741,N_2799);
nor U2956 (N_2956,N_2718,N_2654);
nand U2957 (N_2957,N_2613,N_2645);
or U2958 (N_2958,N_2757,N_2764);
nand U2959 (N_2959,N_2753,N_2688);
nand U2960 (N_2960,N_2613,N_2684);
nand U2961 (N_2961,N_2742,N_2793);
nand U2962 (N_2962,N_2796,N_2700);
and U2963 (N_2963,N_2772,N_2782);
nor U2964 (N_2964,N_2682,N_2735);
nand U2965 (N_2965,N_2767,N_2625);
nand U2966 (N_2966,N_2788,N_2738);
or U2967 (N_2967,N_2648,N_2764);
and U2968 (N_2968,N_2667,N_2748);
and U2969 (N_2969,N_2717,N_2780);
and U2970 (N_2970,N_2684,N_2707);
and U2971 (N_2971,N_2661,N_2605);
and U2972 (N_2972,N_2796,N_2764);
xor U2973 (N_2973,N_2784,N_2799);
nand U2974 (N_2974,N_2629,N_2656);
nand U2975 (N_2975,N_2707,N_2613);
nand U2976 (N_2976,N_2618,N_2759);
nand U2977 (N_2977,N_2609,N_2656);
nor U2978 (N_2978,N_2705,N_2669);
nor U2979 (N_2979,N_2673,N_2721);
nand U2980 (N_2980,N_2631,N_2756);
nor U2981 (N_2981,N_2675,N_2685);
nand U2982 (N_2982,N_2791,N_2696);
or U2983 (N_2983,N_2603,N_2738);
nand U2984 (N_2984,N_2787,N_2679);
and U2985 (N_2985,N_2611,N_2681);
or U2986 (N_2986,N_2738,N_2697);
nor U2987 (N_2987,N_2673,N_2646);
nand U2988 (N_2988,N_2667,N_2740);
and U2989 (N_2989,N_2715,N_2664);
nand U2990 (N_2990,N_2652,N_2700);
or U2991 (N_2991,N_2649,N_2605);
nand U2992 (N_2992,N_2657,N_2658);
and U2993 (N_2993,N_2793,N_2757);
or U2994 (N_2994,N_2654,N_2762);
or U2995 (N_2995,N_2696,N_2755);
and U2996 (N_2996,N_2654,N_2781);
nor U2997 (N_2997,N_2638,N_2613);
xnor U2998 (N_2998,N_2751,N_2711);
nor U2999 (N_2999,N_2631,N_2682);
and U3000 (N_3000,N_2856,N_2874);
nand U3001 (N_3001,N_2859,N_2946);
or U3002 (N_3002,N_2961,N_2833);
nor U3003 (N_3003,N_2953,N_2929);
nand U3004 (N_3004,N_2814,N_2873);
nand U3005 (N_3005,N_2800,N_2891);
nor U3006 (N_3006,N_2981,N_2885);
or U3007 (N_3007,N_2869,N_2995);
or U3008 (N_3008,N_2998,N_2912);
nand U3009 (N_3009,N_2960,N_2922);
nor U3010 (N_3010,N_2824,N_2906);
and U3011 (N_3011,N_2997,N_2955);
nor U3012 (N_3012,N_2808,N_2902);
and U3013 (N_3013,N_2936,N_2820);
and U3014 (N_3014,N_2849,N_2894);
and U3015 (N_3015,N_2973,N_2903);
nor U3016 (N_3016,N_2887,N_2803);
nand U3017 (N_3017,N_2957,N_2971);
nand U3018 (N_3018,N_2816,N_2880);
or U3019 (N_3019,N_2951,N_2937);
or U3020 (N_3020,N_2990,N_2974);
nor U3021 (N_3021,N_2879,N_2886);
and U3022 (N_3022,N_2934,N_2994);
nand U3023 (N_3023,N_2949,N_2930);
nand U3024 (N_3024,N_2901,N_2966);
nand U3025 (N_3025,N_2989,N_2977);
nor U3026 (N_3026,N_2918,N_2809);
nand U3027 (N_3027,N_2825,N_2813);
and U3028 (N_3028,N_2913,N_2892);
nor U3029 (N_3029,N_2802,N_2923);
nand U3030 (N_3030,N_2840,N_2991);
or U3031 (N_3031,N_2841,N_2948);
nand U3032 (N_3032,N_2890,N_2927);
nand U3033 (N_3033,N_2863,N_2867);
nand U3034 (N_3034,N_2862,N_2958);
nor U3035 (N_3035,N_2865,N_2805);
or U3036 (N_3036,N_2920,N_2895);
nand U3037 (N_3037,N_2806,N_2963);
nor U3038 (N_3038,N_2975,N_2804);
nand U3039 (N_3039,N_2871,N_2943);
nor U3040 (N_3040,N_2819,N_2868);
nor U3041 (N_3041,N_2870,N_2938);
or U3042 (N_3042,N_2876,N_2928);
and U3043 (N_3043,N_2910,N_2843);
or U3044 (N_3044,N_2911,N_2993);
or U3045 (N_3045,N_2838,N_2828);
nand U3046 (N_3046,N_2831,N_2982);
nand U3047 (N_3047,N_2959,N_2944);
and U3048 (N_3048,N_2899,N_2933);
and U3049 (N_3049,N_2978,N_2896);
and U3050 (N_3050,N_2907,N_2812);
nand U3051 (N_3051,N_2857,N_2964);
nor U3052 (N_3052,N_2817,N_2926);
and U3053 (N_3053,N_2931,N_2810);
nand U3054 (N_3054,N_2832,N_2999);
nand U3055 (N_3055,N_2965,N_2945);
or U3056 (N_3056,N_2818,N_2919);
nor U3057 (N_3057,N_2845,N_2815);
or U3058 (N_3058,N_2969,N_2839);
nor U3059 (N_3059,N_2883,N_2846);
nor U3060 (N_3060,N_2992,N_2858);
or U3061 (N_3061,N_2935,N_2988);
and U3062 (N_3062,N_2898,N_2984);
and U3063 (N_3063,N_2864,N_2897);
nor U3064 (N_3064,N_2801,N_2872);
and U3065 (N_3065,N_2852,N_2904);
and U3066 (N_3066,N_2861,N_2821);
nand U3067 (N_3067,N_2996,N_2914);
nor U3068 (N_3068,N_2829,N_2925);
or U3069 (N_3069,N_2924,N_2967);
nor U3070 (N_3070,N_2976,N_2877);
nand U3071 (N_3071,N_2942,N_2947);
and U3072 (N_3072,N_2836,N_2807);
and U3073 (N_3073,N_2917,N_2983);
or U3074 (N_3074,N_2844,N_2968);
nor U3075 (N_3075,N_2889,N_2826);
or U3076 (N_3076,N_2987,N_2822);
or U3077 (N_3077,N_2909,N_2940);
nand U3078 (N_3078,N_2878,N_2905);
or U3079 (N_3079,N_2952,N_2954);
or U3080 (N_3080,N_2875,N_2866);
nand U3081 (N_3081,N_2980,N_2956);
or U3082 (N_3082,N_2986,N_2939);
nor U3083 (N_3083,N_2881,N_2851);
and U3084 (N_3084,N_2932,N_2916);
nor U3085 (N_3085,N_2847,N_2921);
or U3086 (N_3086,N_2855,N_2837);
and U3087 (N_3087,N_2915,N_2941);
nor U3088 (N_3088,N_2908,N_2860);
nor U3089 (N_3089,N_2888,N_2950);
nor U3090 (N_3090,N_2842,N_2827);
nand U3091 (N_3091,N_2962,N_2854);
and U3092 (N_3092,N_2853,N_2979);
nor U3093 (N_3093,N_2823,N_2985);
or U3094 (N_3094,N_2848,N_2834);
nand U3095 (N_3095,N_2811,N_2972);
or U3096 (N_3096,N_2884,N_2900);
nand U3097 (N_3097,N_2882,N_2970);
and U3098 (N_3098,N_2850,N_2893);
nor U3099 (N_3099,N_2835,N_2830);
or U3100 (N_3100,N_2958,N_2889);
or U3101 (N_3101,N_2847,N_2930);
or U3102 (N_3102,N_2984,N_2936);
nand U3103 (N_3103,N_2925,N_2930);
nor U3104 (N_3104,N_2876,N_2955);
nand U3105 (N_3105,N_2999,N_2959);
nand U3106 (N_3106,N_2922,N_2969);
xor U3107 (N_3107,N_2947,N_2913);
or U3108 (N_3108,N_2806,N_2922);
nor U3109 (N_3109,N_2930,N_2845);
and U3110 (N_3110,N_2943,N_2841);
nor U3111 (N_3111,N_2999,N_2903);
nor U3112 (N_3112,N_2881,N_2836);
nor U3113 (N_3113,N_2846,N_2816);
nor U3114 (N_3114,N_2914,N_2881);
nor U3115 (N_3115,N_2879,N_2828);
nor U3116 (N_3116,N_2881,N_2886);
nor U3117 (N_3117,N_2991,N_2884);
nor U3118 (N_3118,N_2935,N_2884);
nand U3119 (N_3119,N_2950,N_2928);
and U3120 (N_3120,N_2802,N_2926);
nand U3121 (N_3121,N_2975,N_2890);
or U3122 (N_3122,N_2808,N_2929);
xnor U3123 (N_3123,N_2892,N_2876);
nand U3124 (N_3124,N_2936,N_2962);
and U3125 (N_3125,N_2805,N_2965);
nor U3126 (N_3126,N_2924,N_2977);
nor U3127 (N_3127,N_2863,N_2870);
or U3128 (N_3128,N_2945,N_2835);
nand U3129 (N_3129,N_2965,N_2816);
xor U3130 (N_3130,N_2985,N_2975);
nor U3131 (N_3131,N_2831,N_2839);
and U3132 (N_3132,N_2909,N_2912);
nor U3133 (N_3133,N_2881,N_2925);
nor U3134 (N_3134,N_2947,N_2923);
and U3135 (N_3135,N_2844,N_2802);
nor U3136 (N_3136,N_2991,N_2971);
nor U3137 (N_3137,N_2932,N_2948);
and U3138 (N_3138,N_2939,N_2833);
and U3139 (N_3139,N_2954,N_2947);
or U3140 (N_3140,N_2857,N_2996);
nor U3141 (N_3141,N_2995,N_2912);
and U3142 (N_3142,N_2916,N_2909);
nand U3143 (N_3143,N_2864,N_2938);
and U3144 (N_3144,N_2821,N_2988);
nand U3145 (N_3145,N_2877,N_2845);
nand U3146 (N_3146,N_2991,N_2833);
and U3147 (N_3147,N_2821,N_2932);
and U3148 (N_3148,N_2952,N_2977);
nand U3149 (N_3149,N_2949,N_2805);
and U3150 (N_3150,N_2850,N_2937);
or U3151 (N_3151,N_2884,N_2993);
nand U3152 (N_3152,N_2874,N_2844);
or U3153 (N_3153,N_2820,N_2956);
nand U3154 (N_3154,N_2946,N_2807);
nor U3155 (N_3155,N_2928,N_2902);
nand U3156 (N_3156,N_2939,N_2881);
nand U3157 (N_3157,N_2819,N_2975);
and U3158 (N_3158,N_2830,N_2869);
or U3159 (N_3159,N_2803,N_2851);
nand U3160 (N_3160,N_2871,N_2870);
nand U3161 (N_3161,N_2918,N_2986);
and U3162 (N_3162,N_2828,N_2823);
and U3163 (N_3163,N_2905,N_2931);
nor U3164 (N_3164,N_2881,N_2932);
and U3165 (N_3165,N_2890,N_2838);
nand U3166 (N_3166,N_2851,N_2902);
nor U3167 (N_3167,N_2876,N_2815);
or U3168 (N_3168,N_2928,N_2870);
or U3169 (N_3169,N_2941,N_2889);
or U3170 (N_3170,N_2923,N_2968);
and U3171 (N_3171,N_2956,N_2982);
nor U3172 (N_3172,N_2967,N_2949);
or U3173 (N_3173,N_2811,N_2808);
nor U3174 (N_3174,N_2959,N_2912);
and U3175 (N_3175,N_2918,N_2840);
and U3176 (N_3176,N_2871,N_2812);
nor U3177 (N_3177,N_2904,N_2921);
or U3178 (N_3178,N_2954,N_2991);
and U3179 (N_3179,N_2883,N_2955);
or U3180 (N_3180,N_2869,N_2832);
or U3181 (N_3181,N_2915,N_2942);
and U3182 (N_3182,N_2874,N_2832);
and U3183 (N_3183,N_2817,N_2997);
nand U3184 (N_3184,N_2869,N_2871);
or U3185 (N_3185,N_2997,N_2938);
nor U3186 (N_3186,N_2811,N_2906);
and U3187 (N_3187,N_2893,N_2871);
and U3188 (N_3188,N_2925,N_2886);
nand U3189 (N_3189,N_2860,N_2923);
and U3190 (N_3190,N_2898,N_2922);
and U3191 (N_3191,N_2910,N_2955);
nand U3192 (N_3192,N_2938,N_2847);
and U3193 (N_3193,N_2904,N_2955);
nor U3194 (N_3194,N_2866,N_2879);
xor U3195 (N_3195,N_2975,N_2991);
nor U3196 (N_3196,N_2825,N_2859);
xor U3197 (N_3197,N_2830,N_2921);
nand U3198 (N_3198,N_2837,N_2868);
nor U3199 (N_3199,N_2814,N_2896);
nor U3200 (N_3200,N_3188,N_3198);
nor U3201 (N_3201,N_3050,N_3175);
nor U3202 (N_3202,N_3085,N_3015);
nor U3203 (N_3203,N_3096,N_3089);
nand U3204 (N_3204,N_3160,N_3146);
nand U3205 (N_3205,N_3046,N_3019);
or U3206 (N_3206,N_3101,N_3058);
and U3207 (N_3207,N_3075,N_3162);
and U3208 (N_3208,N_3167,N_3077);
or U3209 (N_3209,N_3071,N_3095);
or U3210 (N_3210,N_3025,N_3147);
nor U3211 (N_3211,N_3117,N_3044);
nor U3212 (N_3212,N_3183,N_3136);
and U3213 (N_3213,N_3047,N_3082);
or U3214 (N_3214,N_3007,N_3010);
or U3215 (N_3215,N_3110,N_3139);
and U3216 (N_3216,N_3114,N_3187);
and U3217 (N_3217,N_3121,N_3184);
and U3218 (N_3218,N_3126,N_3115);
nand U3219 (N_3219,N_3111,N_3173);
nand U3220 (N_3220,N_3185,N_3151);
and U3221 (N_3221,N_3169,N_3144);
and U3222 (N_3222,N_3065,N_3178);
and U3223 (N_3223,N_3195,N_3098);
and U3224 (N_3224,N_3141,N_3135);
or U3225 (N_3225,N_3153,N_3033);
or U3226 (N_3226,N_3070,N_3100);
or U3227 (N_3227,N_3036,N_3061);
nor U3228 (N_3228,N_3016,N_3009);
or U3229 (N_3229,N_3097,N_3055);
or U3230 (N_3230,N_3013,N_3042);
nand U3231 (N_3231,N_3152,N_3023);
and U3232 (N_3232,N_3022,N_3049);
or U3233 (N_3233,N_3155,N_3193);
nor U3234 (N_3234,N_3052,N_3130);
nand U3235 (N_3235,N_3053,N_3005);
nand U3236 (N_3236,N_3028,N_3035);
nand U3237 (N_3237,N_3069,N_3103);
and U3238 (N_3238,N_3051,N_3179);
and U3239 (N_3239,N_3094,N_3026);
nor U3240 (N_3240,N_3054,N_3003);
nand U3241 (N_3241,N_3149,N_3143);
nand U3242 (N_3242,N_3087,N_3090);
nor U3243 (N_3243,N_3181,N_3004);
nor U3244 (N_3244,N_3020,N_3186);
or U3245 (N_3245,N_3084,N_3159);
nand U3246 (N_3246,N_3060,N_3102);
nand U3247 (N_3247,N_3129,N_3012);
nor U3248 (N_3248,N_3000,N_3040);
nand U3249 (N_3249,N_3158,N_3164);
or U3250 (N_3250,N_3199,N_3088);
and U3251 (N_3251,N_3166,N_3133);
and U3252 (N_3252,N_3001,N_3108);
nand U3253 (N_3253,N_3029,N_3145);
nand U3254 (N_3254,N_3074,N_3018);
and U3255 (N_3255,N_3079,N_3017);
xor U3256 (N_3256,N_3083,N_3031);
nand U3257 (N_3257,N_3172,N_3154);
nor U3258 (N_3258,N_3045,N_3076);
nand U3259 (N_3259,N_3197,N_3128);
nor U3260 (N_3260,N_3113,N_3099);
nor U3261 (N_3261,N_3123,N_3125);
xnor U3262 (N_3262,N_3057,N_3170);
nor U3263 (N_3263,N_3072,N_3073);
nor U3264 (N_3264,N_3038,N_3171);
nand U3265 (N_3265,N_3156,N_3106);
or U3266 (N_3266,N_3177,N_3081);
nand U3267 (N_3267,N_3092,N_3067);
nand U3268 (N_3268,N_3180,N_3161);
nand U3269 (N_3269,N_3093,N_3137);
and U3270 (N_3270,N_3006,N_3043);
nand U3271 (N_3271,N_3191,N_3041);
and U3272 (N_3272,N_3086,N_3119);
and U3273 (N_3273,N_3030,N_3068);
and U3274 (N_3274,N_3064,N_3066);
or U3275 (N_3275,N_3062,N_3091);
nand U3276 (N_3276,N_3002,N_3032);
nor U3277 (N_3277,N_3142,N_3027);
nand U3278 (N_3278,N_3112,N_3021);
or U3279 (N_3279,N_3132,N_3104);
or U3280 (N_3280,N_3124,N_3138);
or U3281 (N_3281,N_3011,N_3182);
and U3282 (N_3282,N_3120,N_3163);
nand U3283 (N_3283,N_3148,N_3039);
or U3284 (N_3284,N_3048,N_3078);
nand U3285 (N_3285,N_3194,N_3118);
and U3286 (N_3286,N_3105,N_3190);
nor U3287 (N_3287,N_3034,N_3157);
or U3288 (N_3288,N_3174,N_3014);
and U3289 (N_3289,N_3196,N_3122);
or U3290 (N_3290,N_3189,N_3134);
or U3291 (N_3291,N_3037,N_3109);
nor U3292 (N_3292,N_3165,N_3107);
nand U3293 (N_3293,N_3008,N_3056);
nor U3294 (N_3294,N_3192,N_3080);
nor U3295 (N_3295,N_3131,N_3127);
and U3296 (N_3296,N_3063,N_3140);
nor U3297 (N_3297,N_3150,N_3116);
nor U3298 (N_3298,N_3059,N_3176);
nor U3299 (N_3299,N_3168,N_3024);
nand U3300 (N_3300,N_3073,N_3043);
and U3301 (N_3301,N_3106,N_3001);
or U3302 (N_3302,N_3150,N_3092);
or U3303 (N_3303,N_3119,N_3024);
or U3304 (N_3304,N_3143,N_3167);
and U3305 (N_3305,N_3060,N_3188);
nor U3306 (N_3306,N_3127,N_3182);
or U3307 (N_3307,N_3045,N_3035);
or U3308 (N_3308,N_3153,N_3049);
or U3309 (N_3309,N_3075,N_3105);
and U3310 (N_3310,N_3078,N_3173);
and U3311 (N_3311,N_3161,N_3022);
nor U3312 (N_3312,N_3004,N_3074);
nand U3313 (N_3313,N_3162,N_3154);
nor U3314 (N_3314,N_3060,N_3112);
nand U3315 (N_3315,N_3079,N_3108);
nand U3316 (N_3316,N_3193,N_3069);
nand U3317 (N_3317,N_3183,N_3150);
xnor U3318 (N_3318,N_3060,N_3097);
and U3319 (N_3319,N_3080,N_3082);
nand U3320 (N_3320,N_3131,N_3134);
nand U3321 (N_3321,N_3106,N_3165);
nor U3322 (N_3322,N_3004,N_3150);
or U3323 (N_3323,N_3110,N_3146);
nor U3324 (N_3324,N_3091,N_3122);
or U3325 (N_3325,N_3146,N_3106);
nor U3326 (N_3326,N_3177,N_3073);
nand U3327 (N_3327,N_3043,N_3138);
and U3328 (N_3328,N_3089,N_3013);
or U3329 (N_3329,N_3063,N_3182);
or U3330 (N_3330,N_3188,N_3067);
xor U3331 (N_3331,N_3088,N_3044);
nor U3332 (N_3332,N_3124,N_3054);
and U3333 (N_3333,N_3165,N_3098);
and U3334 (N_3334,N_3124,N_3010);
and U3335 (N_3335,N_3147,N_3032);
and U3336 (N_3336,N_3068,N_3019);
nand U3337 (N_3337,N_3064,N_3045);
or U3338 (N_3338,N_3163,N_3103);
nor U3339 (N_3339,N_3155,N_3103);
and U3340 (N_3340,N_3174,N_3156);
or U3341 (N_3341,N_3005,N_3027);
and U3342 (N_3342,N_3027,N_3056);
and U3343 (N_3343,N_3024,N_3013);
or U3344 (N_3344,N_3101,N_3135);
nor U3345 (N_3345,N_3101,N_3036);
nand U3346 (N_3346,N_3185,N_3052);
or U3347 (N_3347,N_3189,N_3155);
or U3348 (N_3348,N_3064,N_3138);
nand U3349 (N_3349,N_3094,N_3056);
and U3350 (N_3350,N_3053,N_3165);
nor U3351 (N_3351,N_3175,N_3059);
nor U3352 (N_3352,N_3027,N_3020);
nand U3353 (N_3353,N_3010,N_3067);
nor U3354 (N_3354,N_3017,N_3178);
or U3355 (N_3355,N_3067,N_3032);
nand U3356 (N_3356,N_3161,N_3068);
nor U3357 (N_3357,N_3173,N_3087);
nand U3358 (N_3358,N_3197,N_3165);
nor U3359 (N_3359,N_3170,N_3161);
nand U3360 (N_3360,N_3082,N_3186);
nand U3361 (N_3361,N_3058,N_3182);
nand U3362 (N_3362,N_3031,N_3133);
or U3363 (N_3363,N_3144,N_3109);
nor U3364 (N_3364,N_3125,N_3177);
nor U3365 (N_3365,N_3063,N_3132);
or U3366 (N_3366,N_3175,N_3081);
or U3367 (N_3367,N_3051,N_3151);
or U3368 (N_3368,N_3156,N_3135);
or U3369 (N_3369,N_3051,N_3123);
nand U3370 (N_3370,N_3179,N_3146);
and U3371 (N_3371,N_3193,N_3093);
nand U3372 (N_3372,N_3199,N_3007);
or U3373 (N_3373,N_3195,N_3150);
nor U3374 (N_3374,N_3041,N_3186);
and U3375 (N_3375,N_3088,N_3195);
and U3376 (N_3376,N_3009,N_3078);
nor U3377 (N_3377,N_3034,N_3171);
or U3378 (N_3378,N_3144,N_3082);
nand U3379 (N_3379,N_3172,N_3008);
nand U3380 (N_3380,N_3035,N_3177);
nand U3381 (N_3381,N_3007,N_3185);
or U3382 (N_3382,N_3090,N_3080);
or U3383 (N_3383,N_3094,N_3121);
nor U3384 (N_3384,N_3111,N_3081);
and U3385 (N_3385,N_3054,N_3020);
nor U3386 (N_3386,N_3038,N_3169);
or U3387 (N_3387,N_3047,N_3154);
and U3388 (N_3388,N_3158,N_3058);
or U3389 (N_3389,N_3160,N_3136);
nand U3390 (N_3390,N_3118,N_3149);
and U3391 (N_3391,N_3069,N_3081);
nor U3392 (N_3392,N_3052,N_3177);
nor U3393 (N_3393,N_3061,N_3100);
or U3394 (N_3394,N_3173,N_3029);
and U3395 (N_3395,N_3142,N_3198);
or U3396 (N_3396,N_3107,N_3064);
xor U3397 (N_3397,N_3038,N_3179);
or U3398 (N_3398,N_3054,N_3070);
or U3399 (N_3399,N_3094,N_3068);
nand U3400 (N_3400,N_3264,N_3307);
and U3401 (N_3401,N_3296,N_3277);
and U3402 (N_3402,N_3208,N_3287);
or U3403 (N_3403,N_3293,N_3203);
nor U3404 (N_3404,N_3285,N_3230);
nand U3405 (N_3405,N_3399,N_3303);
and U3406 (N_3406,N_3333,N_3266);
or U3407 (N_3407,N_3314,N_3334);
nor U3408 (N_3408,N_3269,N_3377);
and U3409 (N_3409,N_3283,N_3309);
and U3410 (N_3410,N_3376,N_3388);
nor U3411 (N_3411,N_3379,N_3321);
xnor U3412 (N_3412,N_3366,N_3268);
and U3413 (N_3413,N_3289,N_3292);
nand U3414 (N_3414,N_3360,N_3370);
or U3415 (N_3415,N_3343,N_3326);
and U3416 (N_3416,N_3319,N_3346);
or U3417 (N_3417,N_3240,N_3336);
or U3418 (N_3418,N_3340,N_3337);
nand U3419 (N_3419,N_3391,N_3227);
and U3420 (N_3420,N_3349,N_3272);
nand U3421 (N_3421,N_3342,N_3284);
or U3422 (N_3422,N_3276,N_3217);
or U3423 (N_3423,N_3235,N_3271);
or U3424 (N_3424,N_3219,N_3223);
nor U3425 (N_3425,N_3298,N_3282);
and U3426 (N_3426,N_3384,N_3251);
nand U3427 (N_3427,N_3244,N_3200);
nand U3428 (N_3428,N_3254,N_3329);
or U3429 (N_3429,N_3380,N_3369);
and U3430 (N_3430,N_3318,N_3338);
nand U3431 (N_3431,N_3241,N_3233);
nand U3432 (N_3432,N_3361,N_3280);
nand U3433 (N_3433,N_3308,N_3353);
nor U3434 (N_3434,N_3339,N_3239);
and U3435 (N_3435,N_3218,N_3205);
and U3436 (N_3436,N_3225,N_3273);
nor U3437 (N_3437,N_3204,N_3215);
and U3438 (N_3438,N_3226,N_3363);
nand U3439 (N_3439,N_3274,N_3359);
nor U3440 (N_3440,N_3324,N_3221);
nand U3441 (N_3441,N_3371,N_3356);
nor U3442 (N_3442,N_3220,N_3236);
and U3443 (N_3443,N_3259,N_3348);
or U3444 (N_3444,N_3228,N_3216);
nor U3445 (N_3445,N_3253,N_3263);
nor U3446 (N_3446,N_3290,N_3312);
or U3447 (N_3447,N_3232,N_3238);
nor U3448 (N_3448,N_3352,N_3341);
nand U3449 (N_3449,N_3301,N_3270);
nand U3450 (N_3450,N_3202,N_3330);
or U3451 (N_3451,N_3316,N_3247);
and U3452 (N_3452,N_3327,N_3392);
nand U3453 (N_3453,N_3389,N_3306);
and U3454 (N_3454,N_3210,N_3397);
nand U3455 (N_3455,N_3257,N_3393);
nand U3456 (N_3456,N_3390,N_3364);
nand U3457 (N_3457,N_3212,N_3351);
nor U3458 (N_3458,N_3386,N_3354);
and U3459 (N_3459,N_3286,N_3288);
or U3460 (N_3460,N_3211,N_3345);
nor U3461 (N_3461,N_3382,N_3234);
nor U3462 (N_3462,N_3237,N_3299);
and U3463 (N_3463,N_3350,N_3315);
nor U3464 (N_3464,N_3331,N_3249);
nor U3465 (N_3465,N_3291,N_3302);
nand U3466 (N_3466,N_3378,N_3385);
and U3467 (N_3467,N_3248,N_3347);
nand U3468 (N_3468,N_3267,N_3305);
or U3469 (N_3469,N_3367,N_3335);
or U3470 (N_3470,N_3256,N_3242);
and U3471 (N_3471,N_3313,N_3245);
nor U3472 (N_3472,N_3278,N_3322);
nand U3473 (N_3473,N_3320,N_3317);
or U3474 (N_3474,N_3325,N_3281);
nor U3475 (N_3475,N_3323,N_3252);
nor U3476 (N_3476,N_3365,N_3243);
and U3477 (N_3477,N_3209,N_3229);
nor U3478 (N_3478,N_3300,N_3368);
nand U3479 (N_3479,N_3311,N_3265);
or U3480 (N_3480,N_3374,N_3213);
nor U3481 (N_3481,N_3255,N_3260);
and U3482 (N_3482,N_3258,N_3355);
or U3483 (N_3483,N_3373,N_3395);
and U3484 (N_3484,N_3297,N_3295);
and U3485 (N_3485,N_3328,N_3332);
nor U3486 (N_3486,N_3396,N_3304);
and U3487 (N_3487,N_3357,N_3214);
and U3488 (N_3488,N_3279,N_3250);
nor U3489 (N_3489,N_3381,N_3398);
or U3490 (N_3490,N_3358,N_3275);
and U3491 (N_3491,N_3262,N_3201);
nand U3492 (N_3492,N_3383,N_3310);
nand U3493 (N_3493,N_3222,N_3261);
and U3494 (N_3494,N_3207,N_3344);
or U3495 (N_3495,N_3372,N_3294);
xor U3496 (N_3496,N_3206,N_3387);
and U3497 (N_3497,N_3375,N_3231);
nand U3498 (N_3498,N_3246,N_3394);
nand U3499 (N_3499,N_3362,N_3224);
or U3500 (N_3500,N_3212,N_3203);
xnor U3501 (N_3501,N_3321,N_3387);
or U3502 (N_3502,N_3248,N_3299);
nor U3503 (N_3503,N_3348,N_3254);
nand U3504 (N_3504,N_3296,N_3212);
nor U3505 (N_3505,N_3265,N_3232);
or U3506 (N_3506,N_3330,N_3260);
or U3507 (N_3507,N_3289,N_3357);
nand U3508 (N_3508,N_3214,N_3375);
and U3509 (N_3509,N_3371,N_3342);
xnor U3510 (N_3510,N_3203,N_3298);
or U3511 (N_3511,N_3394,N_3386);
nand U3512 (N_3512,N_3220,N_3370);
and U3513 (N_3513,N_3274,N_3254);
and U3514 (N_3514,N_3374,N_3256);
xor U3515 (N_3515,N_3305,N_3292);
nor U3516 (N_3516,N_3299,N_3378);
and U3517 (N_3517,N_3217,N_3257);
and U3518 (N_3518,N_3202,N_3252);
and U3519 (N_3519,N_3227,N_3377);
and U3520 (N_3520,N_3294,N_3391);
and U3521 (N_3521,N_3256,N_3296);
or U3522 (N_3522,N_3267,N_3383);
nor U3523 (N_3523,N_3228,N_3270);
or U3524 (N_3524,N_3277,N_3267);
nand U3525 (N_3525,N_3306,N_3322);
nand U3526 (N_3526,N_3317,N_3253);
nor U3527 (N_3527,N_3327,N_3398);
and U3528 (N_3528,N_3293,N_3305);
nand U3529 (N_3529,N_3306,N_3354);
or U3530 (N_3530,N_3377,N_3389);
nor U3531 (N_3531,N_3303,N_3396);
and U3532 (N_3532,N_3246,N_3358);
nand U3533 (N_3533,N_3203,N_3325);
nor U3534 (N_3534,N_3364,N_3235);
and U3535 (N_3535,N_3272,N_3388);
or U3536 (N_3536,N_3399,N_3254);
nand U3537 (N_3537,N_3208,N_3313);
nor U3538 (N_3538,N_3276,N_3235);
nor U3539 (N_3539,N_3281,N_3257);
nor U3540 (N_3540,N_3215,N_3274);
and U3541 (N_3541,N_3208,N_3320);
nor U3542 (N_3542,N_3200,N_3323);
nand U3543 (N_3543,N_3295,N_3327);
nor U3544 (N_3544,N_3264,N_3379);
nor U3545 (N_3545,N_3282,N_3334);
nor U3546 (N_3546,N_3356,N_3265);
and U3547 (N_3547,N_3335,N_3256);
or U3548 (N_3548,N_3359,N_3242);
nor U3549 (N_3549,N_3297,N_3310);
or U3550 (N_3550,N_3220,N_3336);
or U3551 (N_3551,N_3337,N_3206);
and U3552 (N_3552,N_3357,N_3253);
or U3553 (N_3553,N_3309,N_3375);
and U3554 (N_3554,N_3381,N_3269);
nand U3555 (N_3555,N_3389,N_3341);
nor U3556 (N_3556,N_3248,N_3301);
and U3557 (N_3557,N_3337,N_3346);
or U3558 (N_3558,N_3376,N_3206);
and U3559 (N_3559,N_3231,N_3213);
or U3560 (N_3560,N_3315,N_3225);
and U3561 (N_3561,N_3320,N_3332);
xor U3562 (N_3562,N_3367,N_3304);
or U3563 (N_3563,N_3262,N_3269);
nor U3564 (N_3564,N_3382,N_3220);
nand U3565 (N_3565,N_3391,N_3201);
nor U3566 (N_3566,N_3340,N_3278);
and U3567 (N_3567,N_3394,N_3349);
nor U3568 (N_3568,N_3285,N_3379);
nor U3569 (N_3569,N_3252,N_3316);
nand U3570 (N_3570,N_3227,N_3238);
nor U3571 (N_3571,N_3318,N_3297);
or U3572 (N_3572,N_3390,N_3357);
nand U3573 (N_3573,N_3300,N_3232);
or U3574 (N_3574,N_3306,N_3273);
nor U3575 (N_3575,N_3379,N_3224);
nor U3576 (N_3576,N_3232,N_3239);
nand U3577 (N_3577,N_3330,N_3243);
and U3578 (N_3578,N_3373,N_3376);
and U3579 (N_3579,N_3343,N_3247);
nor U3580 (N_3580,N_3365,N_3389);
nand U3581 (N_3581,N_3270,N_3202);
nand U3582 (N_3582,N_3220,N_3292);
nand U3583 (N_3583,N_3383,N_3300);
nor U3584 (N_3584,N_3240,N_3218);
nor U3585 (N_3585,N_3218,N_3353);
or U3586 (N_3586,N_3246,N_3247);
nor U3587 (N_3587,N_3222,N_3319);
and U3588 (N_3588,N_3314,N_3322);
nor U3589 (N_3589,N_3331,N_3366);
nand U3590 (N_3590,N_3368,N_3249);
nor U3591 (N_3591,N_3285,N_3294);
nand U3592 (N_3592,N_3320,N_3233);
or U3593 (N_3593,N_3397,N_3220);
or U3594 (N_3594,N_3244,N_3292);
nor U3595 (N_3595,N_3393,N_3379);
nor U3596 (N_3596,N_3297,N_3344);
nor U3597 (N_3597,N_3248,N_3249);
xnor U3598 (N_3598,N_3294,N_3286);
and U3599 (N_3599,N_3254,N_3368);
and U3600 (N_3600,N_3494,N_3580);
and U3601 (N_3601,N_3453,N_3406);
or U3602 (N_3602,N_3487,N_3426);
xnor U3603 (N_3603,N_3522,N_3536);
nor U3604 (N_3604,N_3405,N_3549);
and U3605 (N_3605,N_3596,N_3563);
and U3606 (N_3606,N_3553,N_3440);
nand U3607 (N_3607,N_3532,N_3485);
nand U3608 (N_3608,N_3471,N_3562);
nor U3609 (N_3609,N_3530,N_3495);
nor U3610 (N_3610,N_3551,N_3548);
or U3611 (N_3611,N_3497,N_3476);
and U3612 (N_3612,N_3493,N_3430);
nand U3613 (N_3613,N_3537,N_3540);
and U3614 (N_3614,N_3436,N_3462);
or U3615 (N_3615,N_3459,N_3467);
or U3616 (N_3616,N_3427,N_3445);
and U3617 (N_3617,N_3525,N_3458);
or U3618 (N_3618,N_3531,N_3552);
and U3619 (N_3619,N_3435,N_3450);
nand U3620 (N_3620,N_3533,N_3577);
or U3621 (N_3621,N_3508,N_3564);
nor U3622 (N_3622,N_3446,N_3439);
or U3623 (N_3623,N_3401,N_3403);
and U3624 (N_3624,N_3469,N_3437);
nor U3625 (N_3625,N_3490,N_3557);
nand U3626 (N_3626,N_3418,N_3466);
and U3627 (N_3627,N_3500,N_3491);
nor U3628 (N_3628,N_3443,N_3586);
nor U3629 (N_3629,N_3472,N_3432);
nor U3630 (N_3630,N_3504,N_3511);
or U3631 (N_3631,N_3544,N_3507);
nor U3632 (N_3632,N_3464,N_3543);
or U3633 (N_3633,N_3416,N_3528);
and U3634 (N_3634,N_3569,N_3502);
and U3635 (N_3635,N_3468,N_3474);
nand U3636 (N_3636,N_3428,N_3519);
or U3637 (N_3637,N_3415,N_3576);
nand U3638 (N_3638,N_3589,N_3411);
nor U3639 (N_3639,N_3566,N_3409);
nand U3640 (N_3640,N_3425,N_3587);
nor U3641 (N_3641,N_3441,N_3524);
and U3642 (N_3642,N_3595,N_3575);
or U3643 (N_3643,N_3514,N_3588);
nand U3644 (N_3644,N_3534,N_3527);
and U3645 (N_3645,N_3599,N_3579);
or U3646 (N_3646,N_3594,N_3456);
xor U3647 (N_3647,N_3565,N_3410);
nand U3648 (N_3648,N_3499,N_3463);
or U3649 (N_3649,N_3518,N_3545);
and U3650 (N_3650,N_3582,N_3482);
and U3651 (N_3651,N_3556,N_3400);
and U3652 (N_3652,N_3455,N_3479);
nor U3653 (N_3653,N_3470,N_3510);
nand U3654 (N_3654,N_3402,N_3521);
nand U3655 (N_3655,N_3578,N_3422);
nor U3656 (N_3656,N_3509,N_3442);
and U3657 (N_3657,N_3558,N_3496);
nand U3658 (N_3658,N_3567,N_3478);
and U3659 (N_3659,N_3583,N_3429);
nor U3660 (N_3660,N_3423,N_3572);
nor U3661 (N_3661,N_3505,N_3488);
or U3662 (N_3662,N_3561,N_3535);
and U3663 (N_3663,N_3503,N_3452);
nand U3664 (N_3664,N_3475,N_3420);
nor U3665 (N_3665,N_3581,N_3438);
nand U3666 (N_3666,N_3571,N_3538);
xor U3667 (N_3667,N_3513,N_3486);
nor U3668 (N_3668,N_3451,N_3570);
or U3669 (N_3669,N_3407,N_3591);
nand U3670 (N_3670,N_3520,N_3431);
and U3671 (N_3671,N_3444,N_3554);
nand U3672 (N_3672,N_3529,N_3477);
and U3673 (N_3673,N_3483,N_3526);
or U3674 (N_3674,N_3419,N_3457);
nand U3675 (N_3675,N_3568,N_3414);
nand U3676 (N_3676,N_3559,N_3593);
and U3677 (N_3677,N_3584,N_3461);
or U3678 (N_3678,N_3449,N_3448);
nor U3679 (N_3679,N_3421,N_3460);
nor U3680 (N_3680,N_3447,N_3542);
nor U3681 (N_3681,N_3516,N_3515);
or U3682 (N_3682,N_3404,N_3417);
or U3683 (N_3683,N_3501,N_3547);
or U3684 (N_3684,N_3424,N_3413);
and U3685 (N_3685,N_3517,N_3434);
nor U3686 (N_3686,N_3433,N_3484);
nand U3687 (N_3687,N_3489,N_3539);
xor U3688 (N_3688,N_3573,N_3481);
nand U3689 (N_3689,N_3492,N_3585);
nor U3690 (N_3690,N_3473,N_3408);
nand U3691 (N_3691,N_3541,N_3546);
nor U3692 (N_3692,N_3597,N_3498);
and U3693 (N_3693,N_3506,N_3523);
nor U3694 (N_3694,N_3574,N_3560);
nand U3695 (N_3695,N_3598,N_3592);
nand U3696 (N_3696,N_3550,N_3480);
or U3697 (N_3697,N_3512,N_3412);
or U3698 (N_3698,N_3590,N_3555);
nor U3699 (N_3699,N_3465,N_3454);
nand U3700 (N_3700,N_3552,N_3468);
and U3701 (N_3701,N_3463,N_3438);
or U3702 (N_3702,N_3567,N_3586);
nand U3703 (N_3703,N_3482,N_3512);
and U3704 (N_3704,N_3523,N_3571);
or U3705 (N_3705,N_3594,N_3505);
and U3706 (N_3706,N_3416,N_3453);
nor U3707 (N_3707,N_3530,N_3597);
nor U3708 (N_3708,N_3440,N_3505);
nor U3709 (N_3709,N_3548,N_3400);
or U3710 (N_3710,N_3565,N_3522);
nor U3711 (N_3711,N_3507,N_3528);
and U3712 (N_3712,N_3448,N_3569);
and U3713 (N_3713,N_3566,N_3406);
nor U3714 (N_3714,N_3410,N_3542);
and U3715 (N_3715,N_3417,N_3429);
and U3716 (N_3716,N_3568,N_3492);
or U3717 (N_3717,N_3508,N_3529);
nand U3718 (N_3718,N_3428,N_3515);
nor U3719 (N_3719,N_3421,N_3461);
xnor U3720 (N_3720,N_3411,N_3586);
or U3721 (N_3721,N_3436,N_3480);
xor U3722 (N_3722,N_3565,N_3556);
nor U3723 (N_3723,N_3440,N_3558);
nor U3724 (N_3724,N_3558,N_3467);
nor U3725 (N_3725,N_3515,N_3429);
xor U3726 (N_3726,N_3593,N_3539);
nand U3727 (N_3727,N_3547,N_3430);
xor U3728 (N_3728,N_3523,N_3583);
or U3729 (N_3729,N_3447,N_3489);
nand U3730 (N_3730,N_3532,N_3401);
nor U3731 (N_3731,N_3552,N_3550);
nor U3732 (N_3732,N_3587,N_3538);
or U3733 (N_3733,N_3563,N_3591);
nand U3734 (N_3734,N_3509,N_3422);
nand U3735 (N_3735,N_3587,N_3466);
and U3736 (N_3736,N_3501,N_3491);
nor U3737 (N_3737,N_3459,N_3422);
nor U3738 (N_3738,N_3524,N_3584);
nand U3739 (N_3739,N_3512,N_3458);
and U3740 (N_3740,N_3504,N_3435);
and U3741 (N_3741,N_3534,N_3404);
or U3742 (N_3742,N_3555,N_3453);
nand U3743 (N_3743,N_3539,N_3468);
and U3744 (N_3744,N_3407,N_3483);
nor U3745 (N_3745,N_3435,N_3420);
nand U3746 (N_3746,N_3576,N_3420);
or U3747 (N_3747,N_3484,N_3566);
nor U3748 (N_3748,N_3486,N_3410);
nor U3749 (N_3749,N_3492,N_3402);
or U3750 (N_3750,N_3593,N_3554);
nor U3751 (N_3751,N_3408,N_3470);
and U3752 (N_3752,N_3463,N_3507);
or U3753 (N_3753,N_3442,N_3583);
nand U3754 (N_3754,N_3588,N_3410);
nor U3755 (N_3755,N_3579,N_3460);
nand U3756 (N_3756,N_3406,N_3572);
nand U3757 (N_3757,N_3583,N_3557);
and U3758 (N_3758,N_3426,N_3477);
nor U3759 (N_3759,N_3451,N_3589);
and U3760 (N_3760,N_3569,N_3480);
or U3761 (N_3761,N_3551,N_3502);
and U3762 (N_3762,N_3476,N_3501);
or U3763 (N_3763,N_3424,N_3570);
nor U3764 (N_3764,N_3411,N_3500);
and U3765 (N_3765,N_3460,N_3451);
nand U3766 (N_3766,N_3400,N_3422);
nand U3767 (N_3767,N_3535,N_3503);
or U3768 (N_3768,N_3518,N_3419);
nand U3769 (N_3769,N_3542,N_3577);
nor U3770 (N_3770,N_3466,N_3480);
nor U3771 (N_3771,N_3573,N_3526);
nor U3772 (N_3772,N_3535,N_3416);
nor U3773 (N_3773,N_3494,N_3447);
nor U3774 (N_3774,N_3554,N_3565);
and U3775 (N_3775,N_3427,N_3547);
and U3776 (N_3776,N_3465,N_3573);
nor U3777 (N_3777,N_3558,N_3450);
or U3778 (N_3778,N_3441,N_3566);
or U3779 (N_3779,N_3412,N_3458);
nor U3780 (N_3780,N_3459,N_3597);
and U3781 (N_3781,N_3589,N_3573);
nand U3782 (N_3782,N_3501,N_3495);
or U3783 (N_3783,N_3406,N_3514);
nand U3784 (N_3784,N_3426,N_3484);
and U3785 (N_3785,N_3596,N_3512);
and U3786 (N_3786,N_3403,N_3556);
and U3787 (N_3787,N_3588,N_3518);
or U3788 (N_3788,N_3542,N_3527);
or U3789 (N_3789,N_3527,N_3554);
and U3790 (N_3790,N_3474,N_3507);
or U3791 (N_3791,N_3484,N_3565);
nor U3792 (N_3792,N_3489,N_3481);
and U3793 (N_3793,N_3583,N_3500);
or U3794 (N_3794,N_3433,N_3492);
nand U3795 (N_3795,N_3497,N_3463);
or U3796 (N_3796,N_3506,N_3495);
or U3797 (N_3797,N_3465,N_3414);
nand U3798 (N_3798,N_3487,N_3492);
nand U3799 (N_3799,N_3426,N_3444);
and U3800 (N_3800,N_3775,N_3625);
or U3801 (N_3801,N_3765,N_3647);
nor U3802 (N_3802,N_3727,N_3706);
xor U3803 (N_3803,N_3788,N_3690);
nand U3804 (N_3804,N_3646,N_3671);
and U3805 (N_3805,N_3792,N_3728);
nand U3806 (N_3806,N_3740,N_3779);
nand U3807 (N_3807,N_3620,N_3632);
nor U3808 (N_3808,N_3636,N_3637);
and U3809 (N_3809,N_3794,N_3767);
nor U3810 (N_3810,N_3617,N_3757);
and U3811 (N_3811,N_3601,N_3675);
nor U3812 (N_3812,N_3692,N_3662);
or U3813 (N_3813,N_3603,N_3708);
nand U3814 (N_3814,N_3630,N_3752);
nor U3815 (N_3815,N_3658,N_3715);
or U3816 (N_3816,N_3796,N_3781);
and U3817 (N_3817,N_3687,N_3633);
nand U3818 (N_3818,N_3761,N_3750);
and U3819 (N_3819,N_3677,N_3688);
or U3820 (N_3820,N_3741,N_3745);
nor U3821 (N_3821,N_3681,N_3602);
nand U3822 (N_3822,N_3669,N_3700);
and U3823 (N_3823,N_3771,N_3672);
and U3824 (N_3824,N_3698,N_3668);
nand U3825 (N_3825,N_3734,N_3654);
and U3826 (N_3826,N_3748,N_3753);
nor U3827 (N_3827,N_3642,N_3695);
or U3828 (N_3828,N_3665,N_3712);
or U3829 (N_3829,N_3782,N_3713);
nand U3830 (N_3830,N_3684,N_3718);
nand U3831 (N_3831,N_3680,N_3749);
nor U3832 (N_3832,N_3678,N_3778);
or U3833 (N_3833,N_3789,N_3600);
and U3834 (N_3834,N_3766,N_3650);
nand U3835 (N_3835,N_3631,N_3691);
or U3836 (N_3836,N_3670,N_3793);
nor U3837 (N_3837,N_3635,N_3655);
nor U3838 (N_3838,N_3615,N_3787);
nor U3839 (N_3839,N_3685,N_3686);
xor U3840 (N_3840,N_3723,N_3652);
or U3841 (N_3841,N_3744,N_3614);
or U3842 (N_3842,N_3747,N_3661);
nand U3843 (N_3843,N_3711,N_3697);
and U3844 (N_3844,N_3674,N_3693);
or U3845 (N_3845,N_3649,N_3657);
nor U3846 (N_3846,N_3759,N_3772);
or U3847 (N_3847,N_3730,N_3724);
and U3848 (N_3848,N_3703,N_3737);
nor U3849 (N_3849,N_3699,N_3610);
nand U3850 (N_3850,N_3755,N_3716);
or U3851 (N_3851,N_3758,N_3795);
nand U3852 (N_3852,N_3702,N_3664);
nor U3853 (N_3853,N_3621,N_3648);
nand U3854 (N_3854,N_3770,N_3790);
xnor U3855 (N_3855,N_3644,N_3607);
nor U3856 (N_3856,N_3624,N_3729);
or U3857 (N_3857,N_3682,N_3619);
and U3858 (N_3858,N_3705,N_3764);
nor U3859 (N_3859,N_3777,N_3645);
nor U3860 (N_3860,N_3673,N_3616);
and U3861 (N_3861,N_3738,N_3791);
or U3862 (N_3862,N_3634,N_3656);
xor U3863 (N_3863,N_3714,N_3627);
or U3864 (N_3864,N_3701,N_3612);
nor U3865 (N_3865,N_3784,N_3608);
nand U3866 (N_3866,N_3743,N_3722);
nor U3867 (N_3867,N_3604,N_3719);
or U3868 (N_3868,N_3696,N_3694);
nand U3869 (N_3869,N_3731,N_3639);
nand U3870 (N_3870,N_3643,N_3735);
and U3871 (N_3871,N_3683,N_3783);
nand U3872 (N_3872,N_3663,N_3609);
nand U3873 (N_3873,N_3689,N_3638);
or U3874 (N_3874,N_3679,N_3739);
nand U3875 (N_3875,N_3797,N_3799);
nor U3876 (N_3876,N_3732,N_3676);
or U3877 (N_3877,N_3760,N_3726);
and U3878 (N_3878,N_3742,N_3756);
xor U3879 (N_3879,N_3736,N_3660);
nor U3880 (N_3880,N_3763,N_3628);
or U3881 (N_3881,N_3720,N_3667);
nor U3882 (N_3882,N_3733,N_3623);
nor U3883 (N_3883,N_3629,N_3653);
or U3884 (N_3884,N_3709,N_3768);
nor U3885 (N_3885,N_3710,N_3776);
or U3886 (N_3886,N_3611,N_3751);
and U3887 (N_3887,N_3798,N_3773);
nor U3888 (N_3888,N_3746,N_3659);
and U3889 (N_3889,N_3606,N_3754);
or U3890 (N_3890,N_3651,N_3641);
nand U3891 (N_3891,N_3640,N_3725);
nand U3892 (N_3892,N_3780,N_3769);
nor U3893 (N_3893,N_3762,N_3626);
nor U3894 (N_3894,N_3785,N_3605);
nand U3895 (N_3895,N_3622,N_3666);
nor U3896 (N_3896,N_3721,N_3613);
nand U3897 (N_3897,N_3707,N_3704);
and U3898 (N_3898,N_3618,N_3786);
nand U3899 (N_3899,N_3717,N_3774);
nor U3900 (N_3900,N_3648,N_3759);
and U3901 (N_3901,N_3772,N_3782);
nand U3902 (N_3902,N_3797,N_3661);
and U3903 (N_3903,N_3746,N_3733);
and U3904 (N_3904,N_3600,N_3673);
and U3905 (N_3905,N_3762,N_3787);
nor U3906 (N_3906,N_3745,N_3746);
nor U3907 (N_3907,N_3601,N_3784);
nor U3908 (N_3908,N_3628,N_3726);
nor U3909 (N_3909,N_3790,N_3736);
nor U3910 (N_3910,N_3716,N_3774);
xor U3911 (N_3911,N_3603,N_3648);
nand U3912 (N_3912,N_3604,N_3691);
nand U3913 (N_3913,N_3781,N_3706);
xor U3914 (N_3914,N_3605,N_3758);
nor U3915 (N_3915,N_3640,N_3610);
and U3916 (N_3916,N_3660,N_3669);
xnor U3917 (N_3917,N_3678,N_3768);
and U3918 (N_3918,N_3699,N_3608);
nor U3919 (N_3919,N_3645,N_3788);
and U3920 (N_3920,N_3726,N_3791);
nand U3921 (N_3921,N_3760,N_3629);
and U3922 (N_3922,N_3604,N_3660);
or U3923 (N_3923,N_3681,N_3754);
nor U3924 (N_3924,N_3631,N_3604);
nor U3925 (N_3925,N_3775,N_3655);
and U3926 (N_3926,N_3738,N_3665);
nor U3927 (N_3927,N_3719,N_3693);
or U3928 (N_3928,N_3726,N_3756);
nor U3929 (N_3929,N_3677,N_3772);
nor U3930 (N_3930,N_3699,N_3636);
or U3931 (N_3931,N_3673,N_3779);
and U3932 (N_3932,N_3723,N_3610);
nand U3933 (N_3933,N_3752,N_3664);
or U3934 (N_3934,N_3644,N_3675);
and U3935 (N_3935,N_3731,N_3784);
nand U3936 (N_3936,N_3760,N_3736);
xor U3937 (N_3937,N_3784,N_3713);
or U3938 (N_3938,N_3677,N_3694);
nor U3939 (N_3939,N_3736,N_3626);
nor U3940 (N_3940,N_3657,N_3704);
and U3941 (N_3941,N_3754,N_3761);
and U3942 (N_3942,N_3602,N_3778);
or U3943 (N_3943,N_3693,N_3726);
nor U3944 (N_3944,N_3790,N_3607);
nand U3945 (N_3945,N_3733,N_3769);
nor U3946 (N_3946,N_3777,N_3753);
nand U3947 (N_3947,N_3644,N_3774);
or U3948 (N_3948,N_3614,N_3622);
and U3949 (N_3949,N_3683,N_3612);
and U3950 (N_3950,N_3729,N_3612);
nor U3951 (N_3951,N_3774,N_3714);
and U3952 (N_3952,N_3786,N_3743);
nor U3953 (N_3953,N_3785,N_3658);
or U3954 (N_3954,N_3605,N_3711);
and U3955 (N_3955,N_3763,N_3794);
or U3956 (N_3956,N_3731,N_3729);
nor U3957 (N_3957,N_3726,N_3601);
or U3958 (N_3958,N_3731,N_3615);
nor U3959 (N_3959,N_3626,N_3621);
nor U3960 (N_3960,N_3660,N_3702);
or U3961 (N_3961,N_3665,N_3612);
nand U3962 (N_3962,N_3787,N_3660);
nor U3963 (N_3963,N_3657,N_3661);
and U3964 (N_3964,N_3702,N_3721);
nor U3965 (N_3965,N_3731,N_3777);
nand U3966 (N_3966,N_3715,N_3607);
and U3967 (N_3967,N_3618,N_3799);
nand U3968 (N_3968,N_3661,N_3677);
nor U3969 (N_3969,N_3661,N_3606);
and U3970 (N_3970,N_3635,N_3658);
and U3971 (N_3971,N_3600,N_3770);
and U3972 (N_3972,N_3689,N_3712);
or U3973 (N_3973,N_3701,N_3795);
nor U3974 (N_3974,N_3636,N_3627);
nand U3975 (N_3975,N_3790,N_3606);
or U3976 (N_3976,N_3639,N_3608);
nand U3977 (N_3977,N_3792,N_3717);
or U3978 (N_3978,N_3631,N_3644);
and U3979 (N_3979,N_3743,N_3666);
nand U3980 (N_3980,N_3684,N_3753);
nand U3981 (N_3981,N_3761,N_3649);
or U3982 (N_3982,N_3740,N_3704);
or U3983 (N_3983,N_3694,N_3785);
or U3984 (N_3984,N_3640,N_3723);
nor U3985 (N_3985,N_3660,N_3746);
or U3986 (N_3986,N_3729,N_3709);
or U3987 (N_3987,N_3796,N_3658);
or U3988 (N_3988,N_3787,N_3782);
nor U3989 (N_3989,N_3615,N_3753);
or U3990 (N_3990,N_3648,N_3787);
nor U3991 (N_3991,N_3626,N_3768);
and U3992 (N_3992,N_3695,N_3603);
nor U3993 (N_3993,N_3644,N_3660);
nor U3994 (N_3994,N_3687,N_3699);
or U3995 (N_3995,N_3616,N_3755);
or U3996 (N_3996,N_3648,N_3748);
nand U3997 (N_3997,N_3793,N_3640);
or U3998 (N_3998,N_3742,N_3630);
nand U3999 (N_3999,N_3762,N_3601);
and U4000 (N_4000,N_3907,N_3936);
and U4001 (N_4001,N_3854,N_3906);
nor U4002 (N_4002,N_3988,N_3821);
nand U4003 (N_4003,N_3981,N_3855);
and U4004 (N_4004,N_3862,N_3928);
nand U4005 (N_4005,N_3958,N_3895);
and U4006 (N_4006,N_3800,N_3972);
nor U4007 (N_4007,N_3995,N_3980);
or U4008 (N_4008,N_3851,N_3898);
nand U4009 (N_4009,N_3813,N_3835);
nand U4010 (N_4010,N_3804,N_3865);
nand U4011 (N_4011,N_3923,N_3999);
or U4012 (N_4012,N_3987,N_3953);
nand U4013 (N_4013,N_3829,N_3998);
and U4014 (N_4014,N_3979,N_3856);
and U4015 (N_4015,N_3849,N_3875);
nor U4016 (N_4016,N_3834,N_3863);
or U4017 (N_4017,N_3910,N_3963);
or U4018 (N_4018,N_3899,N_3846);
nor U4019 (N_4019,N_3913,N_3891);
and U4020 (N_4020,N_3926,N_3909);
nand U4021 (N_4021,N_3884,N_3803);
and U4022 (N_4022,N_3845,N_3997);
nand U4023 (N_4023,N_3935,N_3982);
nand U4024 (N_4024,N_3925,N_3828);
nand U4025 (N_4025,N_3993,N_3954);
or U4026 (N_4026,N_3857,N_3830);
or U4027 (N_4027,N_3970,N_3808);
and U4028 (N_4028,N_3894,N_3843);
nor U4029 (N_4029,N_3806,N_3927);
nor U4030 (N_4030,N_3989,N_3918);
or U4031 (N_4031,N_3818,N_3990);
or U4032 (N_4032,N_3973,N_3827);
and U4033 (N_4033,N_3893,N_3915);
and U4034 (N_4034,N_3902,N_3873);
or U4035 (N_4035,N_3879,N_3940);
nand U4036 (N_4036,N_3815,N_3967);
nor U4037 (N_4037,N_3921,N_3876);
or U4038 (N_4038,N_3964,N_3872);
nor U4039 (N_4039,N_3831,N_3809);
nor U4040 (N_4040,N_3807,N_3971);
and U4041 (N_4041,N_3817,N_3945);
nor U4042 (N_4042,N_3937,N_3819);
nand U4043 (N_4043,N_3908,N_3983);
and U4044 (N_4044,N_3939,N_3892);
or U4045 (N_4045,N_3962,N_3832);
and U4046 (N_4046,N_3933,N_3942);
nand U4047 (N_4047,N_3969,N_3801);
and U4048 (N_4048,N_3931,N_3991);
nand U4049 (N_4049,N_3886,N_3950);
or U4050 (N_4050,N_3920,N_3816);
nor U4051 (N_4051,N_3974,N_3844);
and U4052 (N_4052,N_3957,N_3841);
and U4053 (N_4053,N_3978,N_3839);
nand U4054 (N_4054,N_3955,N_3826);
xor U4055 (N_4055,N_3805,N_3824);
nand U4056 (N_4056,N_3912,N_3883);
xor U4057 (N_4057,N_3919,N_3948);
and U4058 (N_4058,N_3889,N_3896);
nand U4059 (N_4059,N_3853,N_3871);
nor U4060 (N_4060,N_3901,N_3985);
or U4061 (N_4061,N_3952,N_3882);
nor U4062 (N_4062,N_3848,N_3840);
or U4063 (N_4063,N_3823,N_3992);
nor U4064 (N_4064,N_3975,N_3866);
or U4065 (N_4065,N_3837,N_3924);
nand U4066 (N_4066,N_3994,N_3966);
and U4067 (N_4067,N_3944,N_3885);
and U4068 (N_4068,N_3880,N_3802);
nand U4069 (N_4069,N_3977,N_3838);
nand U4070 (N_4070,N_3864,N_3938);
nor U4071 (N_4071,N_3850,N_3934);
nor U4072 (N_4072,N_3914,N_3874);
and U4073 (N_4073,N_3916,N_3897);
nand U4074 (N_4074,N_3956,N_3947);
nor U4075 (N_4075,N_3903,N_3986);
or U4076 (N_4076,N_3984,N_3941);
nor U4077 (N_4077,N_3904,N_3820);
nor U4078 (N_4078,N_3951,N_3881);
or U4079 (N_4079,N_3949,N_3946);
nand U4080 (N_4080,N_3825,N_3911);
or U4081 (N_4081,N_3961,N_3890);
nand U4082 (N_4082,N_3888,N_3968);
nor U4083 (N_4083,N_3965,N_3878);
nor U4084 (N_4084,N_3868,N_3929);
nor U4085 (N_4085,N_3867,N_3976);
or U4086 (N_4086,N_3858,N_3836);
or U4087 (N_4087,N_3811,N_3842);
and U4088 (N_4088,N_3930,N_3900);
nand U4089 (N_4089,N_3861,N_3932);
and U4090 (N_4090,N_3870,N_3960);
or U4091 (N_4091,N_3905,N_3922);
and U4092 (N_4092,N_3814,N_3833);
and U4093 (N_4093,N_3943,N_3859);
or U4094 (N_4094,N_3810,N_3852);
nor U4095 (N_4095,N_3812,N_3860);
nor U4096 (N_4096,N_3869,N_3917);
nand U4097 (N_4097,N_3887,N_3959);
and U4098 (N_4098,N_3847,N_3996);
or U4099 (N_4099,N_3822,N_3877);
nor U4100 (N_4100,N_3996,N_3914);
nand U4101 (N_4101,N_3807,N_3816);
nor U4102 (N_4102,N_3893,N_3923);
and U4103 (N_4103,N_3846,N_3928);
nor U4104 (N_4104,N_3826,N_3961);
and U4105 (N_4105,N_3944,N_3825);
or U4106 (N_4106,N_3913,N_3966);
nor U4107 (N_4107,N_3975,N_3920);
or U4108 (N_4108,N_3962,N_3961);
nor U4109 (N_4109,N_3874,N_3833);
or U4110 (N_4110,N_3825,N_3876);
nand U4111 (N_4111,N_3838,N_3836);
and U4112 (N_4112,N_3912,N_3973);
or U4113 (N_4113,N_3973,N_3964);
nor U4114 (N_4114,N_3980,N_3807);
xnor U4115 (N_4115,N_3842,N_3952);
nand U4116 (N_4116,N_3983,N_3937);
nand U4117 (N_4117,N_3998,N_3871);
nand U4118 (N_4118,N_3970,N_3968);
and U4119 (N_4119,N_3958,N_3884);
and U4120 (N_4120,N_3853,N_3801);
nor U4121 (N_4121,N_3885,N_3818);
or U4122 (N_4122,N_3923,N_3944);
and U4123 (N_4123,N_3849,N_3990);
or U4124 (N_4124,N_3871,N_3876);
or U4125 (N_4125,N_3833,N_3834);
or U4126 (N_4126,N_3917,N_3891);
or U4127 (N_4127,N_3909,N_3918);
or U4128 (N_4128,N_3809,N_3897);
or U4129 (N_4129,N_3855,N_3825);
nor U4130 (N_4130,N_3994,N_3805);
and U4131 (N_4131,N_3988,N_3987);
nand U4132 (N_4132,N_3918,N_3936);
or U4133 (N_4133,N_3977,N_3942);
and U4134 (N_4134,N_3849,N_3802);
nand U4135 (N_4135,N_3915,N_3854);
and U4136 (N_4136,N_3937,N_3888);
and U4137 (N_4137,N_3932,N_3813);
nor U4138 (N_4138,N_3841,N_3917);
or U4139 (N_4139,N_3823,N_3800);
or U4140 (N_4140,N_3889,N_3884);
nand U4141 (N_4141,N_3951,N_3891);
nand U4142 (N_4142,N_3855,N_3826);
or U4143 (N_4143,N_3975,N_3869);
or U4144 (N_4144,N_3980,N_3930);
and U4145 (N_4145,N_3987,N_3860);
and U4146 (N_4146,N_3853,N_3835);
and U4147 (N_4147,N_3888,N_3872);
or U4148 (N_4148,N_3848,N_3995);
nand U4149 (N_4149,N_3871,N_3847);
nand U4150 (N_4150,N_3832,N_3903);
and U4151 (N_4151,N_3975,N_3865);
nand U4152 (N_4152,N_3843,N_3940);
or U4153 (N_4153,N_3961,N_3818);
and U4154 (N_4154,N_3894,N_3823);
and U4155 (N_4155,N_3994,N_3940);
nor U4156 (N_4156,N_3997,N_3969);
nand U4157 (N_4157,N_3920,N_3979);
and U4158 (N_4158,N_3876,N_3820);
nor U4159 (N_4159,N_3819,N_3978);
and U4160 (N_4160,N_3989,N_3923);
nand U4161 (N_4161,N_3892,N_3826);
or U4162 (N_4162,N_3811,N_3983);
and U4163 (N_4163,N_3855,N_3999);
or U4164 (N_4164,N_3966,N_3818);
nand U4165 (N_4165,N_3848,N_3885);
nand U4166 (N_4166,N_3933,N_3820);
nor U4167 (N_4167,N_3936,N_3944);
nor U4168 (N_4168,N_3800,N_3988);
nor U4169 (N_4169,N_3802,N_3991);
nand U4170 (N_4170,N_3918,N_3924);
nand U4171 (N_4171,N_3817,N_3919);
nand U4172 (N_4172,N_3956,N_3853);
nor U4173 (N_4173,N_3981,N_3897);
nor U4174 (N_4174,N_3846,N_3947);
or U4175 (N_4175,N_3891,N_3832);
and U4176 (N_4176,N_3875,N_3872);
nor U4177 (N_4177,N_3860,N_3993);
nor U4178 (N_4178,N_3943,N_3921);
and U4179 (N_4179,N_3829,N_3800);
and U4180 (N_4180,N_3866,N_3869);
nand U4181 (N_4181,N_3889,N_3914);
and U4182 (N_4182,N_3995,N_3810);
and U4183 (N_4183,N_3851,N_3848);
or U4184 (N_4184,N_3890,N_3904);
nand U4185 (N_4185,N_3802,N_3967);
nor U4186 (N_4186,N_3997,N_3880);
and U4187 (N_4187,N_3930,N_3891);
xor U4188 (N_4188,N_3970,N_3925);
or U4189 (N_4189,N_3886,N_3866);
and U4190 (N_4190,N_3975,N_3911);
nor U4191 (N_4191,N_3897,N_3900);
and U4192 (N_4192,N_3896,N_3846);
and U4193 (N_4193,N_3961,N_3936);
nor U4194 (N_4194,N_3865,N_3964);
or U4195 (N_4195,N_3966,N_3929);
nor U4196 (N_4196,N_3897,N_3803);
or U4197 (N_4197,N_3978,N_3954);
nand U4198 (N_4198,N_3857,N_3815);
nand U4199 (N_4199,N_3835,N_3817);
nand U4200 (N_4200,N_4137,N_4138);
nand U4201 (N_4201,N_4139,N_4005);
or U4202 (N_4202,N_4140,N_4081);
or U4203 (N_4203,N_4177,N_4032);
and U4204 (N_4204,N_4169,N_4050);
and U4205 (N_4205,N_4194,N_4049);
nor U4206 (N_4206,N_4001,N_4136);
nor U4207 (N_4207,N_4092,N_4073);
nand U4208 (N_4208,N_4190,N_4184);
and U4209 (N_4209,N_4052,N_4007);
or U4210 (N_4210,N_4074,N_4173);
or U4211 (N_4211,N_4146,N_4198);
nand U4212 (N_4212,N_4183,N_4028);
nand U4213 (N_4213,N_4004,N_4153);
nor U4214 (N_4214,N_4199,N_4134);
or U4215 (N_4215,N_4022,N_4017);
nand U4216 (N_4216,N_4095,N_4068);
nand U4217 (N_4217,N_4106,N_4055);
and U4218 (N_4218,N_4192,N_4082);
nor U4219 (N_4219,N_4122,N_4119);
nand U4220 (N_4220,N_4030,N_4152);
or U4221 (N_4221,N_4008,N_4167);
nor U4222 (N_4222,N_4179,N_4035);
nor U4223 (N_4223,N_4096,N_4103);
nand U4224 (N_4224,N_4080,N_4175);
and U4225 (N_4225,N_4135,N_4161);
nor U4226 (N_4226,N_4130,N_4056);
or U4227 (N_4227,N_4129,N_4051);
and U4228 (N_4228,N_4057,N_4172);
nor U4229 (N_4229,N_4189,N_4133);
xor U4230 (N_4230,N_4011,N_4012);
or U4231 (N_4231,N_4141,N_4157);
and U4232 (N_4232,N_4180,N_4076);
or U4233 (N_4233,N_4039,N_4085);
nand U4234 (N_4234,N_4072,N_4009);
nand U4235 (N_4235,N_4164,N_4037);
nand U4236 (N_4236,N_4115,N_4053);
and U4237 (N_4237,N_4046,N_4124);
or U4238 (N_4238,N_4196,N_4016);
nand U4239 (N_4239,N_4086,N_4174);
and U4240 (N_4240,N_4041,N_4015);
nand U4241 (N_4241,N_4187,N_4063);
or U4242 (N_4242,N_4117,N_4099);
nand U4243 (N_4243,N_4029,N_4166);
and U4244 (N_4244,N_4059,N_4088);
and U4245 (N_4245,N_4123,N_4128);
and U4246 (N_4246,N_4091,N_4186);
or U4247 (N_4247,N_4062,N_4010);
or U4248 (N_4248,N_4165,N_4145);
and U4249 (N_4249,N_4150,N_4078);
xnor U4250 (N_4250,N_4038,N_4105);
and U4251 (N_4251,N_4191,N_4127);
nand U4252 (N_4252,N_4014,N_4060);
nand U4253 (N_4253,N_4098,N_4197);
or U4254 (N_4254,N_4090,N_4025);
and U4255 (N_4255,N_4147,N_4104);
nand U4256 (N_4256,N_4188,N_4125);
or U4257 (N_4257,N_4048,N_4000);
or U4258 (N_4258,N_4026,N_4185);
and U4259 (N_4259,N_4101,N_4084);
nor U4260 (N_4260,N_4043,N_4158);
and U4261 (N_4261,N_4019,N_4002);
and U4262 (N_4262,N_4155,N_4097);
nand U4263 (N_4263,N_4181,N_4064);
nand U4264 (N_4264,N_4176,N_4083);
nand U4265 (N_4265,N_4054,N_4077);
nor U4266 (N_4266,N_4061,N_4148);
nand U4267 (N_4267,N_4089,N_4065);
and U4268 (N_4268,N_4071,N_4151);
or U4269 (N_4269,N_4149,N_4110);
and U4270 (N_4270,N_4003,N_4093);
or U4271 (N_4271,N_4034,N_4079);
nand U4272 (N_4272,N_4144,N_4036);
nand U4273 (N_4273,N_4031,N_4075);
and U4274 (N_4274,N_4058,N_4126);
nor U4275 (N_4275,N_4163,N_4113);
or U4276 (N_4276,N_4021,N_4070);
nor U4277 (N_4277,N_4023,N_4044);
or U4278 (N_4278,N_4154,N_4024);
and U4279 (N_4279,N_4171,N_4162);
nand U4280 (N_4280,N_4178,N_4118);
or U4281 (N_4281,N_4170,N_4112);
nand U4282 (N_4282,N_4067,N_4018);
or U4283 (N_4283,N_4168,N_4040);
or U4284 (N_4284,N_4020,N_4143);
nand U4285 (N_4285,N_4042,N_4111);
or U4286 (N_4286,N_4156,N_4132);
nand U4287 (N_4287,N_4116,N_4109);
nor U4288 (N_4288,N_4094,N_4159);
and U4289 (N_4289,N_4108,N_4182);
nand U4290 (N_4290,N_4006,N_4114);
nand U4291 (N_4291,N_4033,N_4047);
nand U4292 (N_4292,N_4193,N_4107);
or U4293 (N_4293,N_4027,N_4013);
and U4294 (N_4294,N_4120,N_4131);
nor U4295 (N_4295,N_4102,N_4045);
nand U4296 (N_4296,N_4195,N_4069);
or U4297 (N_4297,N_4142,N_4066);
or U4298 (N_4298,N_4087,N_4160);
and U4299 (N_4299,N_4100,N_4121);
and U4300 (N_4300,N_4042,N_4112);
nor U4301 (N_4301,N_4065,N_4083);
nand U4302 (N_4302,N_4042,N_4066);
or U4303 (N_4303,N_4021,N_4129);
nand U4304 (N_4304,N_4040,N_4103);
nor U4305 (N_4305,N_4099,N_4058);
nor U4306 (N_4306,N_4072,N_4015);
and U4307 (N_4307,N_4089,N_4154);
and U4308 (N_4308,N_4154,N_4050);
nor U4309 (N_4309,N_4023,N_4130);
or U4310 (N_4310,N_4124,N_4188);
nor U4311 (N_4311,N_4054,N_4176);
nand U4312 (N_4312,N_4104,N_4117);
nand U4313 (N_4313,N_4179,N_4175);
or U4314 (N_4314,N_4196,N_4148);
or U4315 (N_4315,N_4136,N_4169);
nor U4316 (N_4316,N_4004,N_4189);
nor U4317 (N_4317,N_4167,N_4189);
and U4318 (N_4318,N_4066,N_4161);
nor U4319 (N_4319,N_4196,N_4105);
and U4320 (N_4320,N_4182,N_4077);
nor U4321 (N_4321,N_4193,N_4078);
or U4322 (N_4322,N_4087,N_4177);
nand U4323 (N_4323,N_4132,N_4074);
or U4324 (N_4324,N_4148,N_4142);
and U4325 (N_4325,N_4153,N_4115);
and U4326 (N_4326,N_4107,N_4124);
nand U4327 (N_4327,N_4079,N_4009);
and U4328 (N_4328,N_4104,N_4016);
and U4329 (N_4329,N_4115,N_4087);
or U4330 (N_4330,N_4102,N_4189);
nand U4331 (N_4331,N_4088,N_4100);
or U4332 (N_4332,N_4122,N_4113);
nand U4333 (N_4333,N_4040,N_4146);
nor U4334 (N_4334,N_4141,N_4039);
nand U4335 (N_4335,N_4074,N_4037);
nor U4336 (N_4336,N_4049,N_4179);
xor U4337 (N_4337,N_4017,N_4039);
nand U4338 (N_4338,N_4179,N_4025);
nor U4339 (N_4339,N_4177,N_4010);
or U4340 (N_4340,N_4082,N_4041);
xnor U4341 (N_4341,N_4087,N_4050);
or U4342 (N_4342,N_4109,N_4013);
nand U4343 (N_4343,N_4191,N_4074);
nand U4344 (N_4344,N_4108,N_4021);
nand U4345 (N_4345,N_4194,N_4131);
nand U4346 (N_4346,N_4002,N_4011);
and U4347 (N_4347,N_4100,N_4011);
nor U4348 (N_4348,N_4023,N_4051);
or U4349 (N_4349,N_4101,N_4053);
or U4350 (N_4350,N_4094,N_4197);
nand U4351 (N_4351,N_4095,N_4007);
nand U4352 (N_4352,N_4116,N_4191);
nand U4353 (N_4353,N_4156,N_4141);
nand U4354 (N_4354,N_4198,N_4035);
nand U4355 (N_4355,N_4084,N_4061);
and U4356 (N_4356,N_4136,N_4066);
nor U4357 (N_4357,N_4042,N_4089);
nand U4358 (N_4358,N_4071,N_4021);
or U4359 (N_4359,N_4198,N_4084);
or U4360 (N_4360,N_4183,N_4135);
and U4361 (N_4361,N_4042,N_4110);
nand U4362 (N_4362,N_4013,N_4127);
and U4363 (N_4363,N_4098,N_4157);
nor U4364 (N_4364,N_4006,N_4040);
and U4365 (N_4365,N_4089,N_4050);
and U4366 (N_4366,N_4170,N_4048);
and U4367 (N_4367,N_4196,N_4083);
nand U4368 (N_4368,N_4151,N_4078);
and U4369 (N_4369,N_4058,N_4111);
xor U4370 (N_4370,N_4189,N_4157);
nand U4371 (N_4371,N_4015,N_4061);
nand U4372 (N_4372,N_4176,N_4193);
nand U4373 (N_4373,N_4163,N_4009);
and U4374 (N_4374,N_4110,N_4185);
nor U4375 (N_4375,N_4137,N_4115);
xor U4376 (N_4376,N_4065,N_4104);
and U4377 (N_4377,N_4187,N_4068);
nor U4378 (N_4378,N_4066,N_4126);
nor U4379 (N_4379,N_4194,N_4192);
and U4380 (N_4380,N_4125,N_4007);
and U4381 (N_4381,N_4068,N_4133);
or U4382 (N_4382,N_4138,N_4157);
and U4383 (N_4383,N_4108,N_4187);
nand U4384 (N_4384,N_4123,N_4197);
nand U4385 (N_4385,N_4052,N_4150);
nor U4386 (N_4386,N_4098,N_4033);
nand U4387 (N_4387,N_4043,N_4000);
nor U4388 (N_4388,N_4037,N_4158);
nor U4389 (N_4389,N_4085,N_4113);
or U4390 (N_4390,N_4108,N_4014);
or U4391 (N_4391,N_4144,N_4072);
and U4392 (N_4392,N_4039,N_4006);
or U4393 (N_4393,N_4068,N_4193);
and U4394 (N_4394,N_4164,N_4074);
nand U4395 (N_4395,N_4163,N_4195);
and U4396 (N_4396,N_4135,N_4163);
xnor U4397 (N_4397,N_4154,N_4150);
nor U4398 (N_4398,N_4130,N_4038);
xor U4399 (N_4399,N_4025,N_4141);
xnor U4400 (N_4400,N_4354,N_4316);
nand U4401 (N_4401,N_4337,N_4391);
nand U4402 (N_4402,N_4234,N_4304);
nand U4403 (N_4403,N_4207,N_4346);
xnor U4404 (N_4404,N_4351,N_4232);
nand U4405 (N_4405,N_4375,N_4238);
and U4406 (N_4406,N_4208,N_4327);
or U4407 (N_4407,N_4203,N_4211);
nand U4408 (N_4408,N_4221,N_4274);
nor U4409 (N_4409,N_4385,N_4204);
or U4410 (N_4410,N_4300,N_4284);
nor U4411 (N_4411,N_4256,N_4380);
and U4412 (N_4412,N_4396,N_4215);
and U4413 (N_4413,N_4226,N_4254);
or U4414 (N_4414,N_4287,N_4271);
nor U4415 (N_4415,N_4214,N_4311);
nand U4416 (N_4416,N_4323,N_4383);
nand U4417 (N_4417,N_4326,N_4286);
or U4418 (N_4418,N_4305,N_4376);
and U4419 (N_4419,N_4355,N_4338);
and U4420 (N_4420,N_4301,N_4366);
and U4421 (N_4421,N_4367,N_4394);
nand U4422 (N_4422,N_4235,N_4297);
or U4423 (N_4423,N_4225,N_4374);
nor U4424 (N_4424,N_4223,N_4349);
nor U4425 (N_4425,N_4369,N_4229);
and U4426 (N_4426,N_4381,N_4213);
or U4427 (N_4427,N_4281,N_4210);
nor U4428 (N_4428,N_4263,N_4291);
or U4429 (N_4429,N_4359,N_4247);
and U4430 (N_4430,N_4280,N_4200);
nor U4431 (N_4431,N_4233,N_4264);
nor U4432 (N_4432,N_4277,N_4331);
and U4433 (N_4433,N_4228,N_4253);
nand U4434 (N_4434,N_4379,N_4219);
nor U4435 (N_4435,N_4356,N_4248);
xnor U4436 (N_4436,N_4290,N_4333);
nand U4437 (N_4437,N_4392,N_4384);
or U4438 (N_4438,N_4236,N_4307);
or U4439 (N_4439,N_4260,N_4372);
and U4440 (N_4440,N_4244,N_4205);
or U4441 (N_4441,N_4257,N_4231);
and U4442 (N_4442,N_4272,N_4270);
xnor U4443 (N_4443,N_4313,N_4388);
or U4444 (N_4444,N_4298,N_4212);
nand U4445 (N_4445,N_4251,N_4397);
or U4446 (N_4446,N_4340,N_4320);
and U4447 (N_4447,N_4329,N_4288);
nor U4448 (N_4448,N_4368,N_4275);
and U4449 (N_4449,N_4365,N_4216);
or U4450 (N_4450,N_4353,N_4330);
and U4451 (N_4451,N_4360,N_4227);
xor U4452 (N_4452,N_4268,N_4373);
xor U4453 (N_4453,N_4312,N_4357);
nor U4454 (N_4454,N_4308,N_4319);
or U4455 (N_4455,N_4362,N_4266);
or U4456 (N_4456,N_4398,N_4371);
nand U4457 (N_4457,N_4240,N_4255);
or U4458 (N_4458,N_4339,N_4387);
nand U4459 (N_4459,N_4309,N_4334);
or U4460 (N_4460,N_4241,N_4395);
and U4461 (N_4461,N_4341,N_4344);
nand U4462 (N_4462,N_4222,N_4265);
and U4463 (N_4463,N_4273,N_4269);
nor U4464 (N_4464,N_4336,N_4378);
nand U4465 (N_4465,N_4243,N_4306);
and U4466 (N_4466,N_4328,N_4347);
nand U4467 (N_4467,N_4246,N_4296);
and U4468 (N_4468,N_4345,N_4399);
nand U4469 (N_4469,N_4217,N_4314);
nand U4470 (N_4470,N_4202,N_4237);
and U4471 (N_4471,N_4324,N_4292);
nor U4472 (N_4472,N_4335,N_4332);
or U4473 (N_4473,N_4201,N_4317);
xnor U4474 (N_4474,N_4364,N_4325);
and U4475 (N_4475,N_4343,N_4230);
nor U4476 (N_4476,N_4262,N_4245);
nor U4477 (N_4477,N_4276,N_4294);
xnor U4478 (N_4478,N_4318,N_4249);
nor U4479 (N_4479,N_4224,N_4239);
nor U4480 (N_4480,N_4315,N_4370);
nor U4481 (N_4481,N_4377,N_4220);
and U4482 (N_4482,N_4390,N_4389);
xor U4483 (N_4483,N_4358,N_4252);
xor U4484 (N_4484,N_4206,N_4302);
and U4485 (N_4485,N_4348,N_4386);
nor U4486 (N_4486,N_4283,N_4250);
and U4487 (N_4487,N_4299,N_4382);
or U4488 (N_4488,N_4278,N_4261);
nor U4489 (N_4489,N_4352,N_4218);
nor U4490 (N_4490,N_4289,N_4393);
nand U4491 (N_4491,N_4295,N_4267);
nand U4492 (N_4492,N_4259,N_4321);
nor U4493 (N_4493,N_4322,N_4285);
or U4494 (N_4494,N_4361,N_4303);
and U4495 (N_4495,N_4242,N_4342);
xor U4496 (N_4496,N_4350,N_4282);
nand U4497 (N_4497,N_4279,N_4258);
nor U4498 (N_4498,N_4310,N_4363);
nand U4499 (N_4499,N_4209,N_4293);
nor U4500 (N_4500,N_4282,N_4212);
or U4501 (N_4501,N_4316,N_4200);
nand U4502 (N_4502,N_4274,N_4392);
and U4503 (N_4503,N_4213,N_4292);
nand U4504 (N_4504,N_4240,N_4256);
nor U4505 (N_4505,N_4299,N_4222);
nand U4506 (N_4506,N_4282,N_4231);
or U4507 (N_4507,N_4335,N_4340);
nand U4508 (N_4508,N_4399,N_4272);
and U4509 (N_4509,N_4353,N_4298);
xor U4510 (N_4510,N_4294,N_4366);
and U4511 (N_4511,N_4275,N_4339);
and U4512 (N_4512,N_4293,N_4301);
or U4513 (N_4513,N_4260,N_4349);
or U4514 (N_4514,N_4355,N_4337);
or U4515 (N_4515,N_4236,N_4399);
nor U4516 (N_4516,N_4251,N_4245);
nor U4517 (N_4517,N_4220,N_4239);
nor U4518 (N_4518,N_4243,N_4377);
and U4519 (N_4519,N_4257,N_4363);
nor U4520 (N_4520,N_4339,N_4303);
nor U4521 (N_4521,N_4288,N_4342);
and U4522 (N_4522,N_4277,N_4361);
nand U4523 (N_4523,N_4314,N_4278);
nand U4524 (N_4524,N_4377,N_4265);
nor U4525 (N_4525,N_4232,N_4220);
nand U4526 (N_4526,N_4264,N_4287);
and U4527 (N_4527,N_4250,N_4262);
or U4528 (N_4528,N_4216,N_4369);
and U4529 (N_4529,N_4291,N_4236);
nand U4530 (N_4530,N_4305,N_4282);
nor U4531 (N_4531,N_4210,N_4226);
and U4532 (N_4532,N_4335,N_4290);
nand U4533 (N_4533,N_4297,N_4313);
nor U4534 (N_4534,N_4207,N_4200);
nand U4535 (N_4535,N_4340,N_4321);
nand U4536 (N_4536,N_4283,N_4264);
and U4537 (N_4537,N_4373,N_4270);
nand U4538 (N_4538,N_4320,N_4252);
or U4539 (N_4539,N_4362,N_4392);
nor U4540 (N_4540,N_4324,N_4229);
and U4541 (N_4541,N_4311,N_4239);
nand U4542 (N_4542,N_4223,N_4242);
and U4543 (N_4543,N_4370,N_4327);
nor U4544 (N_4544,N_4265,N_4218);
nor U4545 (N_4545,N_4263,N_4296);
and U4546 (N_4546,N_4317,N_4334);
or U4547 (N_4547,N_4300,N_4204);
nand U4548 (N_4548,N_4206,N_4338);
or U4549 (N_4549,N_4318,N_4264);
and U4550 (N_4550,N_4280,N_4375);
nand U4551 (N_4551,N_4232,N_4396);
and U4552 (N_4552,N_4363,N_4324);
nand U4553 (N_4553,N_4300,N_4327);
nand U4554 (N_4554,N_4327,N_4254);
nor U4555 (N_4555,N_4310,N_4279);
or U4556 (N_4556,N_4293,N_4281);
nand U4557 (N_4557,N_4288,N_4332);
or U4558 (N_4558,N_4328,N_4343);
nand U4559 (N_4559,N_4355,N_4273);
nor U4560 (N_4560,N_4347,N_4312);
and U4561 (N_4561,N_4273,N_4279);
or U4562 (N_4562,N_4263,N_4286);
and U4563 (N_4563,N_4331,N_4367);
nor U4564 (N_4564,N_4292,N_4233);
and U4565 (N_4565,N_4220,N_4234);
nand U4566 (N_4566,N_4304,N_4315);
nand U4567 (N_4567,N_4351,N_4343);
or U4568 (N_4568,N_4292,N_4226);
or U4569 (N_4569,N_4397,N_4265);
or U4570 (N_4570,N_4225,N_4251);
or U4571 (N_4571,N_4352,N_4289);
nand U4572 (N_4572,N_4363,N_4238);
nand U4573 (N_4573,N_4377,N_4371);
or U4574 (N_4574,N_4351,N_4302);
or U4575 (N_4575,N_4264,N_4302);
or U4576 (N_4576,N_4215,N_4229);
and U4577 (N_4577,N_4324,N_4376);
nor U4578 (N_4578,N_4262,N_4361);
nand U4579 (N_4579,N_4278,N_4299);
nor U4580 (N_4580,N_4237,N_4291);
or U4581 (N_4581,N_4250,N_4364);
nor U4582 (N_4582,N_4248,N_4297);
and U4583 (N_4583,N_4352,N_4330);
nor U4584 (N_4584,N_4210,N_4304);
and U4585 (N_4585,N_4341,N_4267);
nor U4586 (N_4586,N_4282,N_4204);
and U4587 (N_4587,N_4362,N_4395);
nand U4588 (N_4588,N_4351,N_4368);
and U4589 (N_4589,N_4259,N_4392);
nand U4590 (N_4590,N_4234,N_4253);
or U4591 (N_4591,N_4234,N_4303);
nor U4592 (N_4592,N_4216,N_4212);
nor U4593 (N_4593,N_4292,N_4274);
and U4594 (N_4594,N_4342,N_4276);
nor U4595 (N_4595,N_4212,N_4245);
nand U4596 (N_4596,N_4309,N_4212);
nand U4597 (N_4597,N_4214,N_4336);
or U4598 (N_4598,N_4324,N_4247);
nor U4599 (N_4599,N_4391,N_4380);
nand U4600 (N_4600,N_4430,N_4481);
and U4601 (N_4601,N_4547,N_4543);
nor U4602 (N_4602,N_4446,N_4420);
nor U4603 (N_4603,N_4521,N_4524);
and U4604 (N_4604,N_4525,N_4549);
nor U4605 (N_4605,N_4472,N_4477);
nor U4606 (N_4606,N_4432,N_4480);
nor U4607 (N_4607,N_4449,N_4577);
nand U4608 (N_4608,N_4519,N_4502);
nand U4609 (N_4609,N_4450,N_4506);
or U4610 (N_4610,N_4542,N_4422);
nand U4611 (N_4611,N_4455,N_4591);
nor U4612 (N_4612,N_4579,N_4435);
nand U4613 (N_4613,N_4469,N_4434);
and U4614 (N_4614,N_4575,N_4567);
and U4615 (N_4615,N_4518,N_4517);
and U4616 (N_4616,N_4423,N_4565);
nand U4617 (N_4617,N_4511,N_4488);
and U4618 (N_4618,N_4428,N_4414);
nand U4619 (N_4619,N_4556,N_4476);
or U4620 (N_4620,N_4569,N_4410);
nor U4621 (N_4621,N_4587,N_4408);
and U4622 (N_4622,N_4558,N_4509);
nand U4623 (N_4623,N_4534,N_4593);
and U4624 (N_4624,N_4571,N_4453);
nand U4625 (N_4625,N_4454,N_4496);
and U4626 (N_4626,N_4424,N_4487);
nand U4627 (N_4627,N_4599,N_4507);
or U4628 (N_4628,N_4537,N_4528);
xor U4629 (N_4629,N_4568,N_4574);
nand U4630 (N_4630,N_4595,N_4463);
nand U4631 (N_4631,N_4526,N_4401);
nand U4632 (N_4632,N_4425,N_4426);
xnor U4633 (N_4633,N_4572,N_4527);
nor U4634 (N_4634,N_4514,N_4516);
and U4635 (N_4635,N_4531,N_4419);
nand U4636 (N_4636,N_4465,N_4484);
or U4637 (N_4637,N_4586,N_4532);
or U4638 (N_4638,N_4562,N_4437);
nor U4639 (N_4639,N_4457,N_4548);
and U4640 (N_4640,N_4535,N_4443);
xnor U4641 (N_4641,N_4486,N_4529);
or U4642 (N_4642,N_4545,N_4467);
or U4643 (N_4643,N_4444,N_4564);
nand U4644 (N_4644,N_4536,N_4493);
nor U4645 (N_4645,N_4539,N_4459);
or U4646 (N_4646,N_4466,N_4566);
and U4647 (N_4647,N_4563,N_4471);
and U4648 (N_4648,N_4584,N_4489);
or U4649 (N_4649,N_4560,N_4462);
or U4650 (N_4650,N_4581,N_4540);
and U4651 (N_4651,N_4473,N_4598);
nor U4652 (N_4652,N_4411,N_4533);
nand U4653 (N_4653,N_4482,N_4407);
nand U4654 (N_4654,N_4438,N_4427);
and U4655 (N_4655,N_4485,N_4510);
nand U4656 (N_4656,N_4541,N_4594);
or U4657 (N_4657,N_4580,N_4403);
nor U4658 (N_4658,N_4504,N_4523);
or U4659 (N_4659,N_4479,N_4447);
nor U4660 (N_4660,N_4530,N_4499);
nor U4661 (N_4661,N_4400,N_4413);
nor U4662 (N_4662,N_4458,N_4436);
xnor U4663 (N_4663,N_4559,N_4503);
or U4664 (N_4664,N_4554,N_4590);
or U4665 (N_4665,N_4583,N_4557);
nand U4666 (N_4666,N_4470,N_4513);
and U4667 (N_4667,N_4576,N_4573);
or U4668 (N_4668,N_4440,N_4417);
or U4669 (N_4669,N_4418,N_4448);
nor U4670 (N_4670,N_4585,N_4442);
nor U4671 (N_4671,N_4452,N_4464);
nor U4672 (N_4672,N_4468,N_4597);
nor U4673 (N_4673,N_4490,N_4546);
or U4674 (N_4674,N_4544,N_4421);
xor U4675 (N_4675,N_4588,N_4416);
xnor U4676 (N_4676,N_4409,N_4550);
or U4677 (N_4677,N_4555,N_4498);
and U4678 (N_4678,N_4495,N_4404);
and U4679 (N_4679,N_4515,N_4494);
and U4680 (N_4680,N_4483,N_4439);
nand U4681 (N_4681,N_4478,N_4592);
nor U4682 (N_4682,N_4441,N_4492);
and U4683 (N_4683,N_4500,N_4508);
nand U4684 (N_4684,N_4412,N_4429);
nand U4685 (N_4685,N_4551,N_4538);
and U4686 (N_4686,N_4456,N_4501);
or U4687 (N_4687,N_4553,N_4596);
nor U4688 (N_4688,N_4451,N_4461);
nor U4689 (N_4689,N_4497,N_4570);
nor U4690 (N_4690,N_4460,N_4582);
nand U4691 (N_4691,N_4578,N_4405);
xnor U4692 (N_4692,N_4402,N_4512);
and U4693 (N_4693,N_4491,N_4474);
xnor U4694 (N_4694,N_4561,N_4406);
and U4695 (N_4695,N_4505,N_4520);
nand U4696 (N_4696,N_4475,N_4431);
and U4697 (N_4697,N_4589,N_4445);
xor U4698 (N_4698,N_4552,N_4522);
and U4699 (N_4699,N_4433,N_4415);
nor U4700 (N_4700,N_4436,N_4466);
or U4701 (N_4701,N_4564,N_4530);
nand U4702 (N_4702,N_4487,N_4493);
nor U4703 (N_4703,N_4433,N_4594);
nand U4704 (N_4704,N_4442,N_4402);
nor U4705 (N_4705,N_4402,N_4415);
nor U4706 (N_4706,N_4549,N_4514);
nor U4707 (N_4707,N_4407,N_4550);
nor U4708 (N_4708,N_4434,N_4446);
nand U4709 (N_4709,N_4422,N_4590);
and U4710 (N_4710,N_4488,N_4404);
nand U4711 (N_4711,N_4596,N_4462);
and U4712 (N_4712,N_4518,N_4410);
nor U4713 (N_4713,N_4415,N_4443);
nor U4714 (N_4714,N_4522,N_4473);
nor U4715 (N_4715,N_4573,N_4535);
nor U4716 (N_4716,N_4435,N_4415);
or U4717 (N_4717,N_4442,N_4444);
or U4718 (N_4718,N_4441,N_4407);
nand U4719 (N_4719,N_4413,N_4477);
nand U4720 (N_4720,N_4525,N_4431);
nor U4721 (N_4721,N_4431,N_4540);
and U4722 (N_4722,N_4560,N_4484);
nor U4723 (N_4723,N_4580,N_4458);
nor U4724 (N_4724,N_4573,N_4413);
nor U4725 (N_4725,N_4546,N_4424);
or U4726 (N_4726,N_4572,N_4478);
or U4727 (N_4727,N_4494,N_4459);
nand U4728 (N_4728,N_4427,N_4509);
nand U4729 (N_4729,N_4472,N_4424);
or U4730 (N_4730,N_4597,N_4410);
or U4731 (N_4731,N_4515,N_4408);
and U4732 (N_4732,N_4536,N_4585);
nand U4733 (N_4733,N_4489,N_4576);
or U4734 (N_4734,N_4412,N_4584);
and U4735 (N_4735,N_4590,N_4523);
xnor U4736 (N_4736,N_4546,N_4547);
nor U4737 (N_4737,N_4537,N_4505);
nor U4738 (N_4738,N_4447,N_4521);
nor U4739 (N_4739,N_4432,N_4555);
and U4740 (N_4740,N_4496,N_4519);
nand U4741 (N_4741,N_4428,N_4565);
nand U4742 (N_4742,N_4406,N_4583);
nand U4743 (N_4743,N_4495,N_4434);
nor U4744 (N_4744,N_4547,N_4514);
nor U4745 (N_4745,N_4536,N_4444);
nor U4746 (N_4746,N_4534,N_4500);
or U4747 (N_4747,N_4415,N_4525);
and U4748 (N_4748,N_4437,N_4496);
nor U4749 (N_4749,N_4480,N_4592);
and U4750 (N_4750,N_4440,N_4573);
nor U4751 (N_4751,N_4587,N_4580);
nand U4752 (N_4752,N_4523,N_4423);
or U4753 (N_4753,N_4550,N_4526);
and U4754 (N_4754,N_4563,N_4545);
nor U4755 (N_4755,N_4578,N_4469);
or U4756 (N_4756,N_4576,N_4565);
nand U4757 (N_4757,N_4517,N_4451);
nor U4758 (N_4758,N_4426,N_4590);
and U4759 (N_4759,N_4549,N_4571);
and U4760 (N_4760,N_4595,N_4521);
nand U4761 (N_4761,N_4577,N_4451);
or U4762 (N_4762,N_4569,N_4454);
nor U4763 (N_4763,N_4448,N_4451);
and U4764 (N_4764,N_4595,N_4508);
nor U4765 (N_4765,N_4584,N_4598);
nand U4766 (N_4766,N_4439,N_4592);
or U4767 (N_4767,N_4545,N_4472);
or U4768 (N_4768,N_4576,N_4512);
nand U4769 (N_4769,N_4415,N_4473);
and U4770 (N_4770,N_4514,N_4586);
nor U4771 (N_4771,N_4554,N_4569);
and U4772 (N_4772,N_4522,N_4485);
nand U4773 (N_4773,N_4572,N_4406);
nand U4774 (N_4774,N_4474,N_4414);
nor U4775 (N_4775,N_4468,N_4502);
or U4776 (N_4776,N_4533,N_4570);
and U4777 (N_4777,N_4503,N_4500);
and U4778 (N_4778,N_4456,N_4483);
or U4779 (N_4779,N_4570,N_4581);
nand U4780 (N_4780,N_4547,N_4510);
and U4781 (N_4781,N_4424,N_4448);
nand U4782 (N_4782,N_4473,N_4553);
or U4783 (N_4783,N_4462,N_4400);
and U4784 (N_4784,N_4408,N_4433);
nand U4785 (N_4785,N_4511,N_4522);
nor U4786 (N_4786,N_4491,N_4511);
nor U4787 (N_4787,N_4402,N_4434);
nand U4788 (N_4788,N_4450,N_4420);
xor U4789 (N_4789,N_4411,N_4465);
or U4790 (N_4790,N_4593,N_4473);
nand U4791 (N_4791,N_4582,N_4545);
nor U4792 (N_4792,N_4427,N_4518);
nor U4793 (N_4793,N_4442,N_4550);
or U4794 (N_4794,N_4441,N_4424);
and U4795 (N_4795,N_4450,N_4454);
nand U4796 (N_4796,N_4407,N_4505);
nor U4797 (N_4797,N_4442,N_4594);
nand U4798 (N_4798,N_4569,N_4470);
nor U4799 (N_4799,N_4593,N_4503);
nand U4800 (N_4800,N_4777,N_4768);
nand U4801 (N_4801,N_4741,N_4729);
or U4802 (N_4802,N_4669,N_4720);
or U4803 (N_4803,N_4775,N_4666);
nand U4804 (N_4804,N_4726,N_4750);
xnor U4805 (N_4805,N_4665,N_4641);
nand U4806 (N_4806,N_4639,N_4752);
nor U4807 (N_4807,N_4761,N_4604);
nand U4808 (N_4808,N_4748,N_4769);
nor U4809 (N_4809,N_4677,N_4609);
and U4810 (N_4810,N_4773,N_4684);
and U4811 (N_4811,N_4793,N_4631);
nor U4812 (N_4812,N_4658,N_4643);
and U4813 (N_4813,N_4724,N_4765);
and U4814 (N_4814,N_4617,N_4790);
nand U4815 (N_4815,N_4664,N_4696);
nor U4816 (N_4816,N_4651,N_4672);
or U4817 (N_4817,N_4667,N_4632);
nor U4818 (N_4818,N_4700,N_4787);
and U4819 (N_4819,N_4685,N_4689);
nor U4820 (N_4820,N_4759,N_4762);
nor U4821 (N_4821,N_4786,N_4753);
nand U4822 (N_4822,N_4783,N_4742);
and U4823 (N_4823,N_4723,N_4784);
or U4824 (N_4824,N_4661,N_4659);
or U4825 (N_4825,N_4771,N_4674);
nand U4826 (N_4826,N_4745,N_4738);
and U4827 (N_4827,N_4757,N_4733);
nor U4828 (N_4828,N_4780,N_4764);
or U4829 (N_4829,N_4737,N_4613);
and U4830 (N_4830,N_4755,N_4697);
nor U4831 (N_4831,N_4678,N_4722);
nand U4832 (N_4832,N_4797,N_4714);
nor U4833 (N_4833,N_4623,N_4660);
xor U4834 (N_4834,N_4705,N_4735);
and U4835 (N_4835,N_4608,N_4727);
nor U4836 (N_4836,N_4616,N_4730);
or U4837 (N_4837,N_4682,N_4634);
nor U4838 (N_4838,N_4698,N_4652);
nor U4839 (N_4839,N_4712,N_4781);
nand U4840 (N_4840,N_4703,N_4734);
and U4841 (N_4841,N_4754,N_4646);
nor U4842 (N_4842,N_4789,N_4645);
nor U4843 (N_4843,N_4717,N_4680);
nand U4844 (N_4844,N_4721,N_4638);
and U4845 (N_4845,N_4602,N_4650);
nor U4846 (N_4846,N_4642,N_4605);
nand U4847 (N_4847,N_4760,N_4791);
or U4848 (N_4848,N_4725,N_4635);
and U4849 (N_4849,N_4654,N_4649);
or U4850 (N_4850,N_4612,N_4636);
or U4851 (N_4851,N_4624,N_4628);
nand U4852 (N_4852,N_4719,N_4653);
nor U4853 (N_4853,N_4692,N_4662);
nand U4854 (N_4854,N_4670,N_4776);
nand U4855 (N_4855,N_4648,N_4799);
xnor U4856 (N_4856,N_4770,N_4655);
nand U4857 (N_4857,N_4679,N_4763);
and U4858 (N_4858,N_4625,N_4621);
nand U4859 (N_4859,N_4600,N_4702);
nand U4860 (N_4860,N_4619,N_4676);
nand U4861 (N_4861,N_4728,N_4739);
or U4862 (N_4862,N_4701,N_4681);
or U4863 (N_4863,N_4746,N_4629);
nand U4864 (N_4864,N_4688,N_4663);
nor U4865 (N_4865,N_4690,N_4779);
nor U4866 (N_4866,N_4620,N_4610);
nor U4867 (N_4867,N_4626,N_4601);
nand U4868 (N_4868,N_4647,N_4673);
and U4869 (N_4869,N_4743,N_4756);
nor U4870 (N_4870,N_4668,N_4766);
and U4871 (N_4871,N_4644,N_4710);
and U4872 (N_4872,N_4603,N_4640);
and U4873 (N_4873,N_4686,N_4715);
or U4874 (N_4874,N_4788,N_4606);
and U4875 (N_4875,N_4618,N_4657);
nor U4876 (N_4876,N_4695,N_4731);
and U4877 (N_4877,N_4627,N_4633);
and U4878 (N_4878,N_4694,N_4785);
nor U4879 (N_4879,N_4706,N_4794);
or U4880 (N_4880,N_4751,N_4749);
nor U4881 (N_4881,N_4656,N_4758);
nor U4882 (N_4882,N_4713,N_4622);
nand U4883 (N_4883,N_4691,N_4614);
nor U4884 (N_4884,N_4607,N_4798);
or U4885 (N_4885,N_4687,N_4774);
nor U4886 (N_4886,N_4637,N_4683);
or U4887 (N_4887,N_4693,N_4708);
or U4888 (N_4888,N_4718,N_4615);
or U4889 (N_4889,N_4711,N_4671);
nand U4890 (N_4890,N_4778,N_4704);
xnor U4891 (N_4891,N_4611,N_4630);
and U4892 (N_4892,N_4792,N_4707);
xor U4893 (N_4893,N_4795,N_4716);
xnor U4894 (N_4894,N_4675,N_4772);
xor U4895 (N_4895,N_4740,N_4744);
and U4896 (N_4896,N_4767,N_4782);
nor U4897 (N_4897,N_4732,N_4736);
or U4898 (N_4898,N_4747,N_4709);
and U4899 (N_4899,N_4699,N_4796);
and U4900 (N_4900,N_4715,N_4779);
and U4901 (N_4901,N_4615,N_4751);
nor U4902 (N_4902,N_4748,N_4640);
and U4903 (N_4903,N_4626,N_4737);
and U4904 (N_4904,N_4772,N_4628);
or U4905 (N_4905,N_4772,N_4634);
and U4906 (N_4906,N_4783,N_4719);
and U4907 (N_4907,N_4754,N_4645);
or U4908 (N_4908,N_4644,N_4765);
and U4909 (N_4909,N_4734,N_4713);
or U4910 (N_4910,N_4646,N_4753);
nand U4911 (N_4911,N_4655,N_4753);
or U4912 (N_4912,N_4681,N_4653);
xor U4913 (N_4913,N_4776,N_4713);
or U4914 (N_4914,N_4770,N_4688);
nor U4915 (N_4915,N_4637,N_4723);
nor U4916 (N_4916,N_4659,N_4630);
or U4917 (N_4917,N_4658,N_4611);
or U4918 (N_4918,N_4704,N_4683);
xnor U4919 (N_4919,N_4612,N_4622);
xor U4920 (N_4920,N_4613,N_4722);
or U4921 (N_4921,N_4751,N_4602);
nand U4922 (N_4922,N_4673,N_4650);
or U4923 (N_4923,N_4717,N_4603);
and U4924 (N_4924,N_4676,N_4657);
or U4925 (N_4925,N_4677,N_4670);
xnor U4926 (N_4926,N_4753,N_4775);
nand U4927 (N_4927,N_4790,N_4663);
and U4928 (N_4928,N_4784,N_4794);
or U4929 (N_4929,N_4606,N_4643);
nor U4930 (N_4930,N_4607,N_4682);
and U4931 (N_4931,N_4771,N_4792);
and U4932 (N_4932,N_4725,N_4623);
and U4933 (N_4933,N_4661,N_4789);
and U4934 (N_4934,N_4749,N_4618);
or U4935 (N_4935,N_4625,N_4704);
or U4936 (N_4936,N_4619,N_4777);
or U4937 (N_4937,N_4683,N_4790);
nor U4938 (N_4938,N_4792,N_4702);
or U4939 (N_4939,N_4643,N_4621);
or U4940 (N_4940,N_4674,N_4609);
and U4941 (N_4941,N_4766,N_4785);
and U4942 (N_4942,N_4632,N_4763);
xnor U4943 (N_4943,N_4689,N_4767);
xor U4944 (N_4944,N_4780,N_4672);
nor U4945 (N_4945,N_4769,N_4790);
and U4946 (N_4946,N_4783,N_4674);
nand U4947 (N_4947,N_4768,N_4724);
nor U4948 (N_4948,N_4779,N_4777);
and U4949 (N_4949,N_4722,N_4662);
or U4950 (N_4950,N_4661,N_4664);
xor U4951 (N_4951,N_4640,N_4744);
nand U4952 (N_4952,N_4755,N_4745);
and U4953 (N_4953,N_4641,N_4623);
or U4954 (N_4954,N_4600,N_4754);
or U4955 (N_4955,N_4766,N_4757);
nand U4956 (N_4956,N_4623,N_4749);
nor U4957 (N_4957,N_4794,N_4704);
and U4958 (N_4958,N_4700,N_4630);
and U4959 (N_4959,N_4670,N_4743);
and U4960 (N_4960,N_4735,N_4740);
or U4961 (N_4961,N_4617,N_4728);
or U4962 (N_4962,N_4615,N_4671);
and U4963 (N_4963,N_4747,N_4748);
and U4964 (N_4964,N_4731,N_4793);
nor U4965 (N_4965,N_4753,N_4779);
or U4966 (N_4966,N_4684,N_4731);
nand U4967 (N_4967,N_4738,N_4627);
or U4968 (N_4968,N_4600,N_4788);
or U4969 (N_4969,N_4676,N_4649);
and U4970 (N_4970,N_4775,N_4729);
nor U4971 (N_4971,N_4618,N_4654);
nor U4972 (N_4972,N_4797,N_4762);
or U4973 (N_4973,N_4671,N_4782);
nor U4974 (N_4974,N_4641,N_4759);
and U4975 (N_4975,N_4742,N_4764);
and U4976 (N_4976,N_4695,N_4751);
and U4977 (N_4977,N_4641,N_4710);
nand U4978 (N_4978,N_4736,N_4643);
nor U4979 (N_4979,N_4677,N_4769);
nand U4980 (N_4980,N_4679,N_4761);
nand U4981 (N_4981,N_4770,N_4626);
xor U4982 (N_4982,N_4682,N_4797);
and U4983 (N_4983,N_4672,N_4609);
or U4984 (N_4984,N_4613,N_4781);
or U4985 (N_4985,N_4621,N_4697);
or U4986 (N_4986,N_4718,N_4659);
or U4987 (N_4987,N_4784,N_4796);
nand U4988 (N_4988,N_4777,N_4603);
and U4989 (N_4989,N_4683,N_4651);
and U4990 (N_4990,N_4732,N_4641);
nor U4991 (N_4991,N_4697,N_4612);
and U4992 (N_4992,N_4717,N_4763);
or U4993 (N_4993,N_4629,N_4768);
and U4994 (N_4994,N_4787,N_4797);
or U4995 (N_4995,N_4719,N_4710);
or U4996 (N_4996,N_4662,N_4700);
nand U4997 (N_4997,N_4601,N_4772);
nand U4998 (N_4998,N_4601,N_4711);
and U4999 (N_4999,N_4720,N_4665);
nand UO_0 (O_0,N_4822,N_4921);
nand UO_1 (O_1,N_4829,N_4900);
or UO_2 (O_2,N_4974,N_4809);
nand UO_3 (O_3,N_4848,N_4931);
and UO_4 (O_4,N_4924,N_4872);
nand UO_5 (O_5,N_4891,N_4912);
xor UO_6 (O_6,N_4847,N_4870);
and UO_7 (O_7,N_4975,N_4919);
or UO_8 (O_8,N_4856,N_4863);
nor UO_9 (O_9,N_4986,N_4853);
or UO_10 (O_10,N_4842,N_4917);
and UO_11 (O_11,N_4998,N_4945);
or UO_12 (O_12,N_4966,N_4994);
nor UO_13 (O_13,N_4845,N_4879);
or UO_14 (O_14,N_4837,N_4849);
xor UO_15 (O_15,N_4979,N_4904);
nor UO_16 (O_16,N_4988,N_4996);
nor UO_17 (O_17,N_4946,N_4898);
nor UO_18 (O_18,N_4852,N_4828);
or UO_19 (O_19,N_4936,N_4814);
or UO_20 (O_20,N_4937,N_4833);
and UO_21 (O_21,N_4869,N_4893);
xnor UO_22 (O_22,N_4867,N_4906);
and UO_23 (O_23,N_4816,N_4855);
and UO_24 (O_24,N_4942,N_4815);
or UO_25 (O_25,N_4982,N_4861);
and UO_26 (O_26,N_4883,N_4818);
and UO_27 (O_27,N_4830,N_4927);
nor UO_28 (O_28,N_4953,N_4968);
nand UO_29 (O_29,N_4955,N_4973);
and UO_30 (O_30,N_4956,N_4857);
nor UO_31 (O_31,N_4803,N_4985);
nand UO_32 (O_32,N_4808,N_4963);
nand UO_33 (O_33,N_4965,N_4826);
nor UO_34 (O_34,N_4925,N_4940);
nor UO_35 (O_35,N_4846,N_4922);
nor UO_36 (O_36,N_4881,N_4839);
or UO_37 (O_37,N_4920,N_4929);
or UO_38 (O_38,N_4962,N_4838);
or UO_39 (O_39,N_4810,N_4806);
nand UO_40 (O_40,N_4944,N_4913);
nand UO_41 (O_41,N_4844,N_4841);
or UO_42 (O_42,N_4882,N_4947);
and UO_43 (O_43,N_4878,N_4897);
nor UO_44 (O_44,N_4909,N_4908);
nand UO_45 (O_45,N_4888,N_4800);
nand UO_46 (O_46,N_4802,N_4880);
and UO_47 (O_47,N_4859,N_4840);
and UO_48 (O_48,N_4902,N_4943);
or UO_49 (O_49,N_4819,N_4801);
and UO_50 (O_50,N_4959,N_4860);
nand UO_51 (O_51,N_4989,N_4834);
nand UO_52 (O_52,N_4851,N_4907);
or UO_53 (O_53,N_4957,N_4886);
and UO_54 (O_54,N_4933,N_4875);
and UO_55 (O_55,N_4911,N_4884);
or UO_56 (O_56,N_4971,N_4941);
nand UO_57 (O_57,N_4915,N_4901);
or UO_58 (O_58,N_4843,N_4894);
and UO_59 (O_59,N_4916,N_4811);
or UO_60 (O_60,N_4961,N_4887);
or UO_61 (O_61,N_4821,N_4939);
or UO_62 (O_62,N_4923,N_4964);
nand UO_63 (O_63,N_4999,N_4934);
nand UO_64 (O_64,N_4899,N_4885);
xnor UO_65 (O_65,N_4954,N_4831);
nor UO_66 (O_66,N_4892,N_4984);
nor UO_67 (O_67,N_4823,N_4992);
xor UO_68 (O_68,N_4918,N_4864);
nand UO_69 (O_69,N_4895,N_4970);
or UO_70 (O_70,N_4871,N_4991);
and UO_71 (O_71,N_4952,N_4890);
and UO_72 (O_72,N_4812,N_4868);
nor UO_73 (O_73,N_4980,N_4896);
and UO_74 (O_74,N_4832,N_4951);
nand UO_75 (O_75,N_4873,N_4972);
and UO_76 (O_76,N_4854,N_4995);
and UO_77 (O_77,N_4835,N_4950);
nand UO_78 (O_78,N_4876,N_4866);
or UO_79 (O_79,N_4948,N_4928);
and UO_80 (O_80,N_4949,N_4807);
and UO_81 (O_81,N_4858,N_4820);
nor UO_82 (O_82,N_4889,N_4824);
nor UO_83 (O_83,N_4865,N_4827);
and UO_84 (O_84,N_4938,N_4805);
nor UO_85 (O_85,N_4977,N_4813);
nand UO_86 (O_86,N_4932,N_4969);
nand UO_87 (O_87,N_4983,N_4935);
nand UO_88 (O_88,N_4804,N_4910);
and UO_89 (O_89,N_4958,N_4905);
and UO_90 (O_90,N_4903,N_4850);
xor UO_91 (O_91,N_4926,N_4981);
nor UO_92 (O_92,N_4862,N_4987);
or UO_93 (O_93,N_4960,N_4978);
or UO_94 (O_94,N_4967,N_4817);
and UO_95 (O_95,N_4877,N_4874);
or UO_96 (O_96,N_4976,N_4825);
and UO_97 (O_97,N_4914,N_4990);
and UO_98 (O_98,N_4993,N_4930);
or UO_99 (O_99,N_4836,N_4997);
and UO_100 (O_100,N_4806,N_4851);
xnor UO_101 (O_101,N_4940,N_4895);
nor UO_102 (O_102,N_4840,N_4990);
nand UO_103 (O_103,N_4931,N_4936);
nor UO_104 (O_104,N_4942,N_4801);
nor UO_105 (O_105,N_4930,N_4962);
or UO_106 (O_106,N_4929,N_4854);
xnor UO_107 (O_107,N_4831,N_4967);
or UO_108 (O_108,N_4984,N_4942);
nand UO_109 (O_109,N_4915,N_4930);
nand UO_110 (O_110,N_4912,N_4942);
and UO_111 (O_111,N_4950,N_4957);
nor UO_112 (O_112,N_4875,N_4930);
or UO_113 (O_113,N_4859,N_4985);
or UO_114 (O_114,N_4936,N_4952);
and UO_115 (O_115,N_4987,N_4912);
nor UO_116 (O_116,N_4859,N_4862);
nand UO_117 (O_117,N_4995,N_4968);
and UO_118 (O_118,N_4981,N_4959);
and UO_119 (O_119,N_4827,N_4808);
nand UO_120 (O_120,N_4944,N_4980);
nand UO_121 (O_121,N_4864,N_4910);
and UO_122 (O_122,N_4943,N_4984);
and UO_123 (O_123,N_4966,N_4929);
or UO_124 (O_124,N_4815,N_4922);
or UO_125 (O_125,N_4859,N_4842);
nand UO_126 (O_126,N_4907,N_4848);
nand UO_127 (O_127,N_4986,N_4886);
nor UO_128 (O_128,N_4864,N_4862);
or UO_129 (O_129,N_4935,N_4861);
nand UO_130 (O_130,N_4831,N_4875);
and UO_131 (O_131,N_4925,N_4964);
or UO_132 (O_132,N_4858,N_4870);
and UO_133 (O_133,N_4853,N_4997);
and UO_134 (O_134,N_4868,N_4937);
and UO_135 (O_135,N_4962,N_4809);
nor UO_136 (O_136,N_4906,N_4975);
or UO_137 (O_137,N_4965,N_4991);
nor UO_138 (O_138,N_4832,N_4898);
or UO_139 (O_139,N_4810,N_4813);
and UO_140 (O_140,N_4810,N_4993);
xnor UO_141 (O_141,N_4984,N_4945);
or UO_142 (O_142,N_4913,N_4984);
or UO_143 (O_143,N_4906,N_4950);
or UO_144 (O_144,N_4805,N_4916);
nand UO_145 (O_145,N_4946,N_4942);
nand UO_146 (O_146,N_4811,N_4887);
or UO_147 (O_147,N_4905,N_4814);
or UO_148 (O_148,N_4905,N_4826);
xnor UO_149 (O_149,N_4896,N_4911);
and UO_150 (O_150,N_4927,N_4940);
and UO_151 (O_151,N_4897,N_4839);
nand UO_152 (O_152,N_4830,N_4883);
nand UO_153 (O_153,N_4876,N_4955);
and UO_154 (O_154,N_4908,N_4842);
or UO_155 (O_155,N_4871,N_4868);
or UO_156 (O_156,N_4800,N_4802);
nand UO_157 (O_157,N_4945,N_4921);
or UO_158 (O_158,N_4969,N_4949);
and UO_159 (O_159,N_4836,N_4885);
nand UO_160 (O_160,N_4882,N_4828);
nand UO_161 (O_161,N_4984,N_4801);
or UO_162 (O_162,N_4998,N_4922);
nand UO_163 (O_163,N_4913,N_4926);
nand UO_164 (O_164,N_4822,N_4944);
nor UO_165 (O_165,N_4979,N_4980);
xor UO_166 (O_166,N_4950,N_4980);
nand UO_167 (O_167,N_4861,N_4965);
and UO_168 (O_168,N_4956,N_4850);
nand UO_169 (O_169,N_4900,N_4918);
nand UO_170 (O_170,N_4871,N_4857);
and UO_171 (O_171,N_4959,N_4904);
nor UO_172 (O_172,N_4901,N_4889);
and UO_173 (O_173,N_4878,N_4991);
nor UO_174 (O_174,N_4870,N_4991);
and UO_175 (O_175,N_4921,N_4870);
and UO_176 (O_176,N_4867,N_4870);
xnor UO_177 (O_177,N_4993,N_4955);
and UO_178 (O_178,N_4898,N_4868);
nor UO_179 (O_179,N_4956,N_4900);
or UO_180 (O_180,N_4967,N_4883);
or UO_181 (O_181,N_4883,N_4911);
and UO_182 (O_182,N_4829,N_4982);
or UO_183 (O_183,N_4862,N_4991);
nand UO_184 (O_184,N_4904,N_4906);
and UO_185 (O_185,N_4897,N_4803);
nand UO_186 (O_186,N_4819,N_4855);
nand UO_187 (O_187,N_4933,N_4845);
nand UO_188 (O_188,N_4902,N_4992);
nand UO_189 (O_189,N_4820,N_4889);
nor UO_190 (O_190,N_4961,N_4963);
nand UO_191 (O_191,N_4987,N_4937);
nand UO_192 (O_192,N_4857,N_4932);
and UO_193 (O_193,N_4949,N_4955);
nor UO_194 (O_194,N_4815,N_4858);
nand UO_195 (O_195,N_4961,N_4870);
and UO_196 (O_196,N_4896,N_4960);
nand UO_197 (O_197,N_4849,N_4939);
or UO_198 (O_198,N_4915,N_4997);
or UO_199 (O_199,N_4845,N_4804);
nor UO_200 (O_200,N_4850,N_4826);
and UO_201 (O_201,N_4822,N_4935);
and UO_202 (O_202,N_4806,N_4972);
or UO_203 (O_203,N_4959,N_4953);
nand UO_204 (O_204,N_4951,N_4953);
or UO_205 (O_205,N_4813,N_4938);
nor UO_206 (O_206,N_4857,N_4931);
nor UO_207 (O_207,N_4980,N_4942);
nor UO_208 (O_208,N_4948,N_4874);
nand UO_209 (O_209,N_4811,N_4858);
nor UO_210 (O_210,N_4903,N_4930);
and UO_211 (O_211,N_4860,N_4988);
nand UO_212 (O_212,N_4876,N_4888);
nor UO_213 (O_213,N_4848,N_4915);
or UO_214 (O_214,N_4923,N_4970);
nor UO_215 (O_215,N_4858,N_4801);
nor UO_216 (O_216,N_4841,N_4904);
nand UO_217 (O_217,N_4868,N_4949);
nor UO_218 (O_218,N_4832,N_4812);
nor UO_219 (O_219,N_4841,N_4979);
or UO_220 (O_220,N_4968,N_4846);
and UO_221 (O_221,N_4862,N_4807);
nor UO_222 (O_222,N_4877,N_4962);
or UO_223 (O_223,N_4865,N_4927);
nor UO_224 (O_224,N_4953,N_4933);
nor UO_225 (O_225,N_4817,N_4906);
and UO_226 (O_226,N_4848,N_4961);
and UO_227 (O_227,N_4948,N_4915);
and UO_228 (O_228,N_4854,N_4858);
nand UO_229 (O_229,N_4861,N_4992);
xnor UO_230 (O_230,N_4868,N_4922);
and UO_231 (O_231,N_4902,N_4982);
nor UO_232 (O_232,N_4872,N_4833);
nand UO_233 (O_233,N_4886,N_4879);
or UO_234 (O_234,N_4987,N_4995);
or UO_235 (O_235,N_4942,N_4954);
nor UO_236 (O_236,N_4962,N_4835);
or UO_237 (O_237,N_4801,N_4845);
or UO_238 (O_238,N_4815,N_4872);
nor UO_239 (O_239,N_4870,N_4974);
nand UO_240 (O_240,N_4804,N_4829);
nor UO_241 (O_241,N_4933,N_4880);
nor UO_242 (O_242,N_4960,N_4985);
nand UO_243 (O_243,N_4871,N_4876);
and UO_244 (O_244,N_4916,N_4855);
nand UO_245 (O_245,N_4919,N_4864);
and UO_246 (O_246,N_4895,N_4834);
nand UO_247 (O_247,N_4832,N_4901);
or UO_248 (O_248,N_4865,N_4943);
nand UO_249 (O_249,N_4842,N_4872);
nand UO_250 (O_250,N_4903,N_4882);
nand UO_251 (O_251,N_4847,N_4852);
nor UO_252 (O_252,N_4980,N_4815);
nor UO_253 (O_253,N_4861,N_4995);
and UO_254 (O_254,N_4824,N_4953);
nand UO_255 (O_255,N_4931,N_4994);
nor UO_256 (O_256,N_4919,N_4868);
or UO_257 (O_257,N_4948,N_4843);
and UO_258 (O_258,N_4843,N_4854);
and UO_259 (O_259,N_4982,N_4927);
nor UO_260 (O_260,N_4850,N_4975);
and UO_261 (O_261,N_4925,N_4989);
nor UO_262 (O_262,N_4961,N_4899);
or UO_263 (O_263,N_4899,N_4915);
or UO_264 (O_264,N_4983,N_4987);
nand UO_265 (O_265,N_4966,N_4913);
or UO_266 (O_266,N_4907,N_4843);
nor UO_267 (O_267,N_4846,N_4970);
or UO_268 (O_268,N_4821,N_4967);
or UO_269 (O_269,N_4800,N_4957);
nor UO_270 (O_270,N_4933,N_4819);
and UO_271 (O_271,N_4913,N_4808);
nor UO_272 (O_272,N_4809,N_4944);
nand UO_273 (O_273,N_4877,N_4968);
nor UO_274 (O_274,N_4938,N_4810);
nor UO_275 (O_275,N_4817,N_4883);
or UO_276 (O_276,N_4918,N_4994);
or UO_277 (O_277,N_4833,N_4911);
or UO_278 (O_278,N_4824,N_4954);
and UO_279 (O_279,N_4831,N_4940);
and UO_280 (O_280,N_4980,N_4941);
and UO_281 (O_281,N_4839,N_4981);
or UO_282 (O_282,N_4906,N_4946);
nand UO_283 (O_283,N_4999,N_4899);
nand UO_284 (O_284,N_4869,N_4973);
nand UO_285 (O_285,N_4900,N_4891);
nor UO_286 (O_286,N_4936,N_4945);
nand UO_287 (O_287,N_4957,N_4804);
nor UO_288 (O_288,N_4951,N_4980);
and UO_289 (O_289,N_4991,N_4874);
nor UO_290 (O_290,N_4847,N_4993);
nand UO_291 (O_291,N_4861,N_4840);
or UO_292 (O_292,N_4812,N_4828);
and UO_293 (O_293,N_4935,N_4875);
nand UO_294 (O_294,N_4882,N_4942);
nand UO_295 (O_295,N_4865,N_4988);
nor UO_296 (O_296,N_4940,N_4997);
nand UO_297 (O_297,N_4994,N_4909);
or UO_298 (O_298,N_4983,N_4948);
or UO_299 (O_299,N_4933,N_4860);
and UO_300 (O_300,N_4899,N_4928);
nor UO_301 (O_301,N_4972,N_4903);
or UO_302 (O_302,N_4947,N_4875);
and UO_303 (O_303,N_4988,N_4842);
and UO_304 (O_304,N_4830,N_4914);
and UO_305 (O_305,N_4825,N_4950);
and UO_306 (O_306,N_4939,N_4867);
nor UO_307 (O_307,N_4976,N_4958);
and UO_308 (O_308,N_4837,N_4862);
nand UO_309 (O_309,N_4842,N_4857);
or UO_310 (O_310,N_4861,N_4901);
nand UO_311 (O_311,N_4826,N_4841);
and UO_312 (O_312,N_4849,N_4965);
or UO_313 (O_313,N_4975,N_4813);
nand UO_314 (O_314,N_4886,N_4934);
nor UO_315 (O_315,N_4852,N_4837);
nand UO_316 (O_316,N_4940,N_4859);
nand UO_317 (O_317,N_4822,N_4893);
and UO_318 (O_318,N_4810,N_4924);
or UO_319 (O_319,N_4950,N_4958);
or UO_320 (O_320,N_4911,N_4825);
or UO_321 (O_321,N_4806,N_4889);
nor UO_322 (O_322,N_4816,N_4923);
or UO_323 (O_323,N_4835,N_4919);
nor UO_324 (O_324,N_4899,N_4958);
and UO_325 (O_325,N_4839,N_4884);
or UO_326 (O_326,N_4879,N_4978);
xor UO_327 (O_327,N_4882,N_4816);
nor UO_328 (O_328,N_4957,N_4860);
and UO_329 (O_329,N_4931,N_4808);
nor UO_330 (O_330,N_4997,N_4928);
and UO_331 (O_331,N_4963,N_4838);
nor UO_332 (O_332,N_4830,N_4986);
xnor UO_333 (O_333,N_4875,N_4992);
or UO_334 (O_334,N_4836,N_4880);
and UO_335 (O_335,N_4870,N_4877);
and UO_336 (O_336,N_4911,N_4957);
or UO_337 (O_337,N_4981,N_4982);
nand UO_338 (O_338,N_4891,N_4996);
xnor UO_339 (O_339,N_4978,N_4976);
xnor UO_340 (O_340,N_4989,N_4861);
and UO_341 (O_341,N_4837,N_4802);
nand UO_342 (O_342,N_4807,N_4804);
xor UO_343 (O_343,N_4970,N_4853);
nor UO_344 (O_344,N_4904,N_4901);
nor UO_345 (O_345,N_4862,N_4971);
and UO_346 (O_346,N_4861,N_4986);
nor UO_347 (O_347,N_4999,N_4882);
xor UO_348 (O_348,N_4839,N_4988);
or UO_349 (O_349,N_4970,N_4829);
or UO_350 (O_350,N_4868,N_4872);
or UO_351 (O_351,N_4923,N_4881);
nor UO_352 (O_352,N_4934,N_4943);
xnor UO_353 (O_353,N_4921,N_4869);
and UO_354 (O_354,N_4992,N_4920);
or UO_355 (O_355,N_4808,N_4934);
nand UO_356 (O_356,N_4855,N_4912);
and UO_357 (O_357,N_4851,N_4871);
or UO_358 (O_358,N_4868,N_4893);
or UO_359 (O_359,N_4949,N_4855);
nor UO_360 (O_360,N_4837,N_4974);
or UO_361 (O_361,N_4921,N_4844);
nor UO_362 (O_362,N_4848,N_4801);
nand UO_363 (O_363,N_4940,N_4978);
nand UO_364 (O_364,N_4962,N_4924);
nor UO_365 (O_365,N_4986,N_4849);
nor UO_366 (O_366,N_4892,N_4815);
nor UO_367 (O_367,N_4957,N_4845);
or UO_368 (O_368,N_4947,N_4925);
xnor UO_369 (O_369,N_4821,N_4995);
or UO_370 (O_370,N_4843,N_4994);
nor UO_371 (O_371,N_4810,N_4928);
and UO_372 (O_372,N_4936,N_4803);
nand UO_373 (O_373,N_4838,N_4856);
and UO_374 (O_374,N_4916,N_4876);
nor UO_375 (O_375,N_4877,N_4914);
and UO_376 (O_376,N_4942,N_4956);
or UO_377 (O_377,N_4997,N_4920);
nor UO_378 (O_378,N_4857,N_4911);
and UO_379 (O_379,N_4945,N_4990);
or UO_380 (O_380,N_4864,N_4831);
nand UO_381 (O_381,N_4965,N_4814);
nor UO_382 (O_382,N_4912,N_4984);
or UO_383 (O_383,N_4975,N_4880);
nor UO_384 (O_384,N_4931,N_4938);
nor UO_385 (O_385,N_4944,N_4805);
nand UO_386 (O_386,N_4994,N_4849);
and UO_387 (O_387,N_4887,N_4817);
and UO_388 (O_388,N_4983,N_4883);
nand UO_389 (O_389,N_4985,N_4980);
and UO_390 (O_390,N_4810,N_4808);
nand UO_391 (O_391,N_4936,N_4916);
xnor UO_392 (O_392,N_4867,N_4922);
or UO_393 (O_393,N_4850,N_4936);
nor UO_394 (O_394,N_4873,N_4833);
and UO_395 (O_395,N_4962,N_4905);
or UO_396 (O_396,N_4852,N_4911);
and UO_397 (O_397,N_4823,N_4984);
or UO_398 (O_398,N_4886,N_4947);
xnor UO_399 (O_399,N_4801,N_4894);
and UO_400 (O_400,N_4818,N_4817);
nor UO_401 (O_401,N_4982,N_4833);
and UO_402 (O_402,N_4949,N_4988);
and UO_403 (O_403,N_4872,N_4916);
and UO_404 (O_404,N_4835,N_4873);
nor UO_405 (O_405,N_4953,N_4925);
and UO_406 (O_406,N_4872,N_4998);
nand UO_407 (O_407,N_4893,N_4976);
nand UO_408 (O_408,N_4905,N_4967);
and UO_409 (O_409,N_4979,N_4858);
and UO_410 (O_410,N_4852,N_4923);
nand UO_411 (O_411,N_4854,N_4998);
and UO_412 (O_412,N_4820,N_4976);
nand UO_413 (O_413,N_4904,N_4866);
nand UO_414 (O_414,N_4974,N_4862);
nand UO_415 (O_415,N_4855,N_4907);
nand UO_416 (O_416,N_4838,N_4843);
or UO_417 (O_417,N_4990,N_4978);
nand UO_418 (O_418,N_4931,N_4801);
and UO_419 (O_419,N_4806,N_4872);
nand UO_420 (O_420,N_4909,N_4945);
or UO_421 (O_421,N_4844,N_4962);
nand UO_422 (O_422,N_4859,N_4948);
and UO_423 (O_423,N_4809,N_4835);
nand UO_424 (O_424,N_4889,N_4800);
or UO_425 (O_425,N_4864,N_4933);
or UO_426 (O_426,N_4886,N_4919);
or UO_427 (O_427,N_4820,N_4945);
nand UO_428 (O_428,N_4882,N_4821);
or UO_429 (O_429,N_4926,N_4920);
and UO_430 (O_430,N_4956,N_4869);
and UO_431 (O_431,N_4846,N_4880);
nand UO_432 (O_432,N_4993,N_4833);
or UO_433 (O_433,N_4952,N_4874);
or UO_434 (O_434,N_4875,N_4944);
nand UO_435 (O_435,N_4894,N_4927);
and UO_436 (O_436,N_4925,N_4853);
and UO_437 (O_437,N_4925,N_4871);
nor UO_438 (O_438,N_4851,N_4834);
and UO_439 (O_439,N_4906,N_4961);
nand UO_440 (O_440,N_4869,N_4835);
and UO_441 (O_441,N_4856,N_4929);
and UO_442 (O_442,N_4927,N_4912);
nand UO_443 (O_443,N_4882,N_4817);
and UO_444 (O_444,N_4808,N_4969);
nor UO_445 (O_445,N_4908,N_4918);
nand UO_446 (O_446,N_4898,N_4875);
and UO_447 (O_447,N_4858,N_4899);
or UO_448 (O_448,N_4855,N_4946);
or UO_449 (O_449,N_4995,N_4807);
nand UO_450 (O_450,N_4895,N_4941);
and UO_451 (O_451,N_4879,N_4989);
and UO_452 (O_452,N_4942,N_4844);
nor UO_453 (O_453,N_4922,N_4904);
nor UO_454 (O_454,N_4969,N_4916);
and UO_455 (O_455,N_4836,N_4951);
or UO_456 (O_456,N_4845,N_4853);
or UO_457 (O_457,N_4869,N_4876);
and UO_458 (O_458,N_4897,N_4983);
nand UO_459 (O_459,N_4968,N_4876);
nor UO_460 (O_460,N_4969,N_4936);
nand UO_461 (O_461,N_4877,N_4903);
nand UO_462 (O_462,N_4853,N_4937);
nor UO_463 (O_463,N_4897,N_4829);
and UO_464 (O_464,N_4812,N_4934);
and UO_465 (O_465,N_4944,N_4974);
nor UO_466 (O_466,N_4900,N_4892);
and UO_467 (O_467,N_4909,N_4801);
nor UO_468 (O_468,N_4959,N_4855);
nor UO_469 (O_469,N_4888,N_4804);
nor UO_470 (O_470,N_4928,N_4945);
nand UO_471 (O_471,N_4810,N_4875);
nand UO_472 (O_472,N_4938,N_4800);
and UO_473 (O_473,N_4927,N_4881);
nor UO_474 (O_474,N_4975,N_4844);
or UO_475 (O_475,N_4829,N_4831);
nand UO_476 (O_476,N_4919,N_4903);
and UO_477 (O_477,N_4916,N_4974);
and UO_478 (O_478,N_4915,N_4827);
xor UO_479 (O_479,N_4894,N_4849);
nand UO_480 (O_480,N_4876,N_4867);
or UO_481 (O_481,N_4973,N_4905);
nor UO_482 (O_482,N_4923,N_4963);
nor UO_483 (O_483,N_4973,N_4946);
nand UO_484 (O_484,N_4807,N_4884);
nand UO_485 (O_485,N_4891,N_4863);
or UO_486 (O_486,N_4932,N_4821);
or UO_487 (O_487,N_4866,N_4961);
and UO_488 (O_488,N_4926,N_4908);
nor UO_489 (O_489,N_4860,N_4848);
nor UO_490 (O_490,N_4948,N_4854);
and UO_491 (O_491,N_4804,N_4980);
xnor UO_492 (O_492,N_4802,N_4886);
or UO_493 (O_493,N_4848,N_4993);
or UO_494 (O_494,N_4842,N_4886);
and UO_495 (O_495,N_4878,N_4882);
nor UO_496 (O_496,N_4856,N_4815);
or UO_497 (O_497,N_4816,N_4996);
or UO_498 (O_498,N_4892,N_4847);
or UO_499 (O_499,N_4814,N_4972);
and UO_500 (O_500,N_4800,N_4917);
and UO_501 (O_501,N_4870,N_4951);
nand UO_502 (O_502,N_4877,N_4858);
and UO_503 (O_503,N_4967,N_4979);
nand UO_504 (O_504,N_4855,N_4922);
nor UO_505 (O_505,N_4822,N_4818);
and UO_506 (O_506,N_4966,N_4955);
xor UO_507 (O_507,N_4906,N_4908);
and UO_508 (O_508,N_4882,N_4820);
and UO_509 (O_509,N_4934,N_4984);
nand UO_510 (O_510,N_4853,N_4875);
nor UO_511 (O_511,N_4835,N_4934);
and UO_512 (O_512,N_4997,N_4911);
nor UO_513 (O_513,N_4837,N_4985);
and UO_514 (O_514,N_4900,N_4883);
nor UO_515 (O_515,N_4899,N_4986);
or UO_516 (O_516,N_4910,N_4973);
nand UO_517 (O_517,N_4931,N_4828);
nor UO_518 (O_518,N_4826,N_4827);
and UO_519 (O_519,N_4836,N_4962);
nand UO_520 (O_520,N_4904,N_4974);
nand UO_521 (O_521,N_4870,N_4813);
nand UO_522 (O_522,N_4963,N_4904);
nor UO_523 (O_523,N_4871,N_4922);
or UO_524 (O_524,N_4828,N_4964);
and UO_525 (O_525,N_4928,N_4849);
nor UO_526 (O_526,N_4909,N_4937);
and UO_527 (O_527,N_4801,N_4817);
or UO_528 (O_528,N_4954,N_4968);
or UO_529 (O_529,N_4835,N_4831);
nor UO_530 (O_530,N_4968,N_4910);
and UO_531 (O_531,N_4956,N_4800);
or UO_532 (O_532,N_4963,N_4875);
nor UO_533 (O_533,N_4964,N_4836);
nand UO_534 (O_534,N_4895,N_4934);
nand UO_535 (O_535,N_4937,N_4875);
nor UO_536 (O_536,N_4818,N_4989);
nand UO_537 (O_537,N_4834,N_4813);
nand UO_538 (O_538,N_4989,N_4860);
nand UO_539 (O_539,N_4996,N_4944);
or UO_540 (O_540,N_4930,N_4860);
nor UO_541 (O_541,N_4861,N_4827);
xor UO_542 (O_542,N_4975,N_4807);
nor UO_543 (O_543,N_4967,N_4911);
nor UO_544 (O_544,N_4885,N_4817);
and UO_545 (O_545,N_4943,N_4831);
nand UO_546 (O_546,N_4891,N_4830);
or UO_547 (O_547,N_4810,N_4908);
nor UO_548 (O_548,N_4959,N_4956);
nand UO_549 (O_549,N_4851,N_4825);
or UO_550 (O_550,N_4857,N_4802);
nand UO_551 (O_551,N_4966,N_4914);
nor UO_552 (O_552,N_4975,N_4823);
xnor UO_553 (O_553,N_4980,N_4809);
nand UO_554 (O_554,N_4841,N_4886);
and UO_555 (O_555,N_4814,N_4973);
nand UO_556 (O_556,N_4884,N_4925);
nor UO_557 (O_557,N_4944,N_4854);
nand UO_558 (O_558,N_4819,N_4892);
nand UO_559 (O_559,N_4824,N_4838);
and UO_560 (O_560,N_4970,N_4847);
and UO_561 (O_561,N_4880,N_4934);
nor UO_562 (O_562,N_4966,N_4958);
nor UO_563 (O_563,N_4851,N_4922);
nor UO_564 (O_564,N_4970,N_4930);
or UO_565 (O_565,N_4999,N_4865);
and UO_566 (O_566,N_4968,N_4942);
nand UO_567 (O_567,N_4849,N_4991);
or UO_568 (O_568,N_4838,N_4991);
nand UO_569 (O_569,N_4934,N_4983);
nand UO_570 (O_570,N_4907,N_4826);
or UO_571 (O_571,N_4904,N_4927);
nor UO_572 (O_572,N_4885,N_4911);
or UO_573 (O_573,N_4853,N_4998);
or UO_574 (O_574,N_4831,N_4888);
nor UO_575 (O_575,N_4865,N_4921);
nor UO_576 (O_576,N_4865,N_4951);
or UO_577 (O_577,N_4905,N_4808);
nand UO_578 (O_578,N_4811,N_4995);
nor UO_579 (O_579,N_4910,N_4886);
and UO_580 (O_580,N_4825,N_4920);
and UO_581 (O_581,N_4883,N_4891);
nand UO_582 (O_582,N_4822,N_4922);
nor UO_583 (O_583,N_4825,N_4916);
nand UO_584 (O_584,N_4904,N_4892);
xor UO_585 (O_585,N_4841,N_4854);
nand UO_586 (O_586,N_4941,N_4968);
or UO_587 (O_587,N_4805,N_4966);
nor UO_588 (O_588,N_4862,N_4847);
nand UO_589 (O_589,N_4818,N_4813);
or UO_590 (O_590,N_4916,N_4931);
or UO_591 (O_591,N_4949,N_4930);
or UO_592 (O_592,N_4815,N_4866);
or UO_593 (O_593,N_4802,N_4902);
nand UO_594 (O_594,N_4906,N_4998);
or UO_595 (O_595,N_4837,N_4891);
and UO_596 (O_596,N_4903,N_4911);
xor UO_597 (O_597,N_4823,N_4858);
and UO_598 (O_598,N_4824,N_4844);
and UO_599 (O_599,N_4876,N_4919);
nor UO_600 (O_600,N_4936,N_4903);
or UO_601 (O_601,N_4959,N_4803);
nor UO_602 (O_602,N_4834,N_4875);
and UO_603 (O_603,N_4848,N_4983);
nor UO_604 (O_604,N_4953,N_4989);
or UO_605 (O_605,N_4983,N_4965);
nand UO_606 (O_606,N_4851,N_4998);
nor UO_607 (O_607,N_4803,N_4906);
and UO_608 (O_608,N_4845,N_4887);
nand UO_609 (O_609,N_4831,N_4916);
and UO_610 (O_610,N_4817,N_4859);
nand UO_611 (O_611,N_4961,N_4970);
nand UO_612 (O_612,N_4994,N_4883);
or UO_613 (O_613,N_4932,N_4986);
nand UO_614 (O_614,N_4800,N_4922);
nand UO_615 (O_615,N_4911,N_4951);
nor UO_616 (O_616,N_4925,N_4907);
or UO_617 (O_617,N_4997,N_4957);
and UO_618 (O_618,N_4939,N_4999);
and UO_619 (O_619,N_4962,N_4810);
and UO_620 (O_620,N_4853,N_4801);
or UO_621 (O_621,N_4894,N_4942);
or UO_622 (O_622,N_4911,N_4804);
or UO_623 (O_623,N_4867,N_4819);
nand UO_624 (O_624,N_4983,N_4830);
and UO_625 (O_625,N_4870,N_4940);
nor UO_626 (O_626,N_4882,N_4938);
and UO_627 (O_627,N_4996,N_4817);
or UO_628 (O_628,N_4927,N_4981);
nand UO_629 (O_629,N_4907,N_4956);
nor UO_630 (O_630,N_4841,N_4843);
nor UO_631 (O_631,N_4972,N_4981);
and UO_632 (O_632,N_4803,N_4805);
nand UO_633 (O_633,N_4873,N_4937);
nor UO_634 (O_634,N_4899,N_4808);
or UO_635 (O_635,N_4961,N_4998);
nand UO_636 (O_636,N_4816,N_4846);
and UO_637 (O_637,N_4872,N_4892);
xnor UO_638 (O_638,N_4919,N_4963);
and UO_639 (O_639,N_4847,N_4840);
nand UO_640 (O_640,N_4982,N_4949);
or UO_641 (O_641,N_4823,N_4910);
and UO_642 (O_642,N_4902,N_4899);
and UO_643 (O_643,N_4949,N_4829);
or UO_644 (O_644,N_4818,N_4843);
nor UO_645 (O_645,N_4908,N_4832);
and UO_646 (O_646,N_4865,N_4970);
nand UO_647 (O_647,N_4812,N_4908);
nor UO_648 (O_648,N_4835,N_4848);
nor UO_649 (O_649,N_4946,N_4922);
or UO_650 (O_650,N_4947,N_4867);
nor UO_651 (O_651,N_4819,N_4848);
or UO_652 (O_652,N_4912,N_4808);
xor UO_653 (O_653,N_4877,N_4900);
or UO_654 (O_654,N_4891,N_4940);
or UO_655 (O_655,N_4878,N_4989);
nor UO_656 (O_656,N_4990,N_4810);
nand UO_657 (O_657,N_4924,N_4949);
and UO_658 (O_658,N_4909,N_4842);
nand UO_659 (O_659,N_4848,N_4869);
nor UO_660 (O_660,N_4951,N_4959);
nand UO_661 (O_661,N_4996,N_4947);
or UO_662 (O_662,N_4939,N_4801);
and UO_663 (O_663,N_4906,N_4827);
and UO_664 (O_664,N_4972,N_4821);
and UO_665 (O_665,N_4969,N_4833);
nor UO_666 (O_666,N_4847,N_4994);
or UO_667 (O_667,N_4802,N_4993);
nor UO_668 (O_668,N_4982,N_4999);
nand UO_669 (O_669,N_4875,N_4838);
or UO_670 (O_670,N_4992,N_4954);
or UO_671 (O_671,N_4941,N_4997);
nand UO_672 (O_672,N_4851,N_4881);
nand UO_673 (O_673,N_4887,N_4926);
and UO_674 (O_674,N_4809,N_4867);
nor UO_675 (O_675,N_4905,N_4916);
or UO_676 (O_676,N_4907,N_4813);
nand UO_677 (O_677,N_4852,N_4867);
nor UO_678 (O_678,N_4929,N_4985);
nand UO_679 (O_679,N_4989,N_4913);
or UO_680 (O_680,N_4949,N_4922);
and UO_681 (O_681,N_4995,N_4824);
nand UO_682 (O_682,N_4854,N_4990);
nor UO_683 (O_683,N_4949,N_4843);
nand UO_684 (O_684,N_4900,N_4862);
and UO_685 (O_685,N_4800,N_4952);
or UO_686 (O_686,N_4996,N_4851);
nor UO_687 (O_687,N_4851,N_4993);
or UO_688 (O_688,N_4957,N_4977);
and UO_689 (O_689,N_4851,N_4818);
and UO_690 (O_690,N_4838,N_4880);
nor UO_691 (O_691,N_4860,N_4882);
nor UO_692 (O_692,N_4827,N_4978);
or UO_693 (O_693,N_4879,N_4946);
and UO_694 (O_694,N_4914,N_4823);
and UO_695 (O_695,N_4867,N_4861);
nand UO_696 (O_696,N_4840,N_4905);
nand UO_697 (O_697,N_4906,N_4881);
and UO_698 (O_698,N_4863,N_4805);
nor UO_699 (O_699,N_4993,N_4875);
and UO_700 (O_700,N_4865,N_4934);
and UO_701 (O_701,N_4948,N_4818);
or UO_702 (O_702,N_4801,N_4809);
and UO_703 (O_703,N_4964,N_4891);
nand UO_704 (O_704,N_4963,N_4962);
nand UO_705 (O_705,N_4912,N_4812);
nor UO_706 (O_706,N_4968,N_4946);
or UO_707 (O_707,N_4901,N_4801);
or UO_708 (O_708,N_4976,N_4972);
nand UO_709 (O_709,N_4929,N_4827);
nand UO_710 (O_710,N_4914,N_4928);
nor UO_711 (O_711,N_4972,N_4801);
nand UO_712 (O_712,N_4876,N_4808);
nor UO_713 (O_713,N_4961,N_4980);
and UO_714 (O_714,N_4942,N_4825);
and UO_715 (O_715,N_4816,N_4817);
xor UO_716 (O_716,N_4930,N_4873);
and UO_717 (O_717,N_4825,N_4981);
nor UO_718 (O_718,N_4878,N_4997);
nand UO_719 (O_719,N_4992,N_4972);
or UO_720 (O_720,N_4948,N_4893);
or UO_721 (O_721,N_4955,N_4883);
and UO_722 (O_722,N_4828,N_4905);
nand UO_723 (O_723,N_4969,N_4947);
or UO_724 (O_724,N_4866,N_4966);
nand UO_725 (O_725,N_4945,N_4891);
and UO_726 (O_726,N_4931,N_4836);
nand UO_727 (O_727,N_4902,N_4911);
nor UO_728 (O_728,N_4839,N_4852);
and UO_729 (O_729,N_4935,N_4924);
and UO_730 (O_730,N_4914,N_4980);
or UO_731 (O_731,N_4860,N_4869);
nand UO_732 (O_732,N_4874,N_4891);
nand UO_733 (O_733,N_4881,N_4853);
nor UO_734 (O_734,N_4956,N_4972);
nor UO_735 (O_735,N_4916,N_4972);
or UO_736 (O_736,N_4891,N_4974);
nor UO_737 (O_737,N_4838,N_4896);
or UO_738 (O_738,N_4890,N_4881);
nor UO_739 (O_739,N_4952,N_4888);
or UO_740 (O_740,N_4899,N_4936);
and UO_741 (O_741,N_4814,N_4844);
or UO_742 (O_742,N_4880,N_4853);
nand UO_743 (O_743,N_4809,N_4983);
nor UO_744 (O_744,N_4809,N_4829);
nand UO_745 (O_745,N_4890,N_4827);
or UO_746 (O_746,N_4940,N_4989);
and UO_747 (O_747,N_4981,N_4824);
and UO_748 (O_748,N_4977,N_4964);
or UO_749 (O_749,N_4826,N_4975);
and UO_750 (O_750,N_4844,N_4855);
nor UO_751 (O_751,N_4893,N_4806);
nand UO_752 (O_752,N_4858,N_4835);
nand UO_753 (O_753,N_4892,N_4851);
or UO_754 (O_754,N_4815,N_4857);
or UO_755 (O_755,N_4862,N_4989);
nand UO_756 (O_756,N_4928,N_4873);
nand UO_757 (O_757,N_4995,N_4823);
and UO_758 (O_758,N_4984,N_4835);
nor UO_759 (O_759,N_4878,N_4964);
or UO_760 (O_760,N_4917,N_4887);
and UO_761 (O_761,N_4995,N_4989);
or UO_762 (O_762,N_4857,N_4940);
nand UO_763 (O_763,N_4905,N_4857);
and UO_764 (O_764,N_4857,N_4895);
and UO_765 (O_765,N_4871,N_4895);
nand UO_766 (O_766,N_4803,N_4894);
nand UO_767 (O_767,N_4890,N_4926);
or UO_768 (O_768,N_4943,N_4896);
xor UO_769 (O_769,N_4811,N_4979);
nor UO_770 (O_770,N_4868,N_4874);
nand UO_771 (O_771,N_4814,N_4941);
xor UO_772 (O_772,N_4829,N_4858);
or UO_773 (O_773,N_4816,N_4967);
nor UO_774 (O_774,N_4896,N_4940);
and UO_775 (O_775,N_4972,N_4907);
or UO_776 (O_776,N_4930,N_4945);
nor UO_777 (O_777,N_4934,N_4988);
nor UO_778 (O_778,N_4925,N_4873);
or UO_779 (O_779,N_4861,N_4916);
and UO_780 (O_780,N_4852,N_4992);
and UO_781 (O_781,N_4858,N_4874);
nor UO_782 (O_782,N_4925,N_4856);
nor UO_783 (O_783,N_4813,N_4882);
xor UO_784 (O_784,N_4802,N_4865);
or UO_785 (O_785,N_4966,N_4932);
and UO_786 (O_786,N_4867,N_4917);
or UO_787 (O_787,N_4995,N_4808);
nor UO_788 (O_788,N_4963,N_4979);
and UO_789 (O_789,N_4991,N_4865);
nor UO_790 (O_790,N_4899,N_4895);
and UO_791 (O_791,N_4818,N_4953);
and UO_792 (O_792,N_4962,N_4943);
or UO_793 (O_793,N_4933,N_4993);
or UO_794 (O_794,N_4856,N_4923);
nand UO_795 (O_795,N_4860,N_4865);
or UO_796 (O_796,N_4822,N_4837);
nor UO_797 (O_797,N_4834,N_4945);
nand UO_798 (O_798,N_4905,N_4979);
or UO_799 (O_799,N_4944,N_4815);
and UO_800 (O_800,N_4902,N_4940);
nor UO_801 (O_801,N_4911,N_4930);
or UO_802 (O_802,N_4861,N_4860);
or UO_803 (O_803,N_4847,N_4991);
nand UO_804 (O_804,N_4869,N_4827);
xnor UO_805 (O_805,N_4984,N_4982);
nor UO_806 (O_806,N_4838,N_4893);
nor UO_807 (O_807,N_4895,N_4816);
or UO_808 (O_808,N_4878,N_4928);
and UO_809 (O_809,N_4982,N_4946);
or UO_810 (O_810,N_4825,N_4935);
and UO_811 (O_811,N_4911,N_4929);
nand UO_812 (O_812,N_4834,N_4881);
nor UO_813 (O_813,N_4903,N_4805);
or UO_814 (O_814,N_4958,N_4934);
nor UO_815 (O_815,N_4918,N_4956);
or UO_816 (O_816,N_4935,N_4872);
and UO_817 (O_817,N_4990,N_4943);
and UO_818 (O_818,N_4944,N_4935);
nor UO_819 (O_819,N_4925,N_4887);
nor UO_820 (O_820,N_4918,N_4946);
nand UO_821 (O_821,N_4946,N_4956);
nor UO_822 (O_822,N_4883,N_4997);
nor UO_823 (O_823,N_4829,N_4971);
or UO_824 (O_824,N_4915,N_4958);
nor UO_825 (O_825,N_4961,N_4957);
and UO_826 (O_826,N_4948,N_4996);
nor UO_827 (O_827,N_4971,N_4832);
nand UO_828 (O_828,N_4927,N_4802);
nand UO_829 (O_829,N_4902,N_4929);
xor UO_830 (O_830,N_4938,N_4919);
nand UO_831 (O_831,N_4895,N_4913);
nand UO_832 (O_832,N_4959,N_4901);
nor UO_833 (O_833,N_4951,N_4970);
nand UO_834 (O_834,N_4819,N_4950);
nand UO_835 (O_835,N_4838,N_4883);
and UO_836 (O_836,N_4928,N_4976);
or UO_837 (O_837,N_4828,N_4950);
nand UO_838 (O_838,N_4838,N_4884);
nor UO_839 (O_839,N_4832,N_4999);
nor UO_840 (O_840,N_4898,N_4855);
or UO_841 (O_841,N_4981,N_4934);
nor UO_842 (O_842,N_4853,N_4932);
nand UO_843 (O_843,N_4968,N_4976);
nand UO_844 (O_844,N_4926,N_4935);
or UO_845 (O_845,N_4967,N_4916);
and UO_846 (O_846,N_4917,N_4891);
or UO_847 (O_847,N_4937,N_4844);
or UO_848 (O_848,N_4975,N_4977);
nor UO_849 (O_849,N_4872,N_4951);
and UO_850 (O_850,N_4912,N_4892);
and UO_851 (O_851,N_4920,N_4942);
nor UO_852 (O_852,N_4948,N_4894);
and UO_853 (O_853,N_4816,N_4990);
xnor UO_854 (O_854,N_4895,N_4824);
nand UO_855 (O_855,N_4820,N_4954);
nor UO_856 (O_856,N_4837,N_4939);
or UO_857 (O_857,N_4851,N_4943);
nand UO_858 (O_858,N_4807,N_4925);
nand UO_859 (O_859,N_4865,N_4859);
nor UO_860 (O_860,N_4814,N_4893);
and UO_861 (O_861,N_4800,N_4824);
nand UO_862 (O_862,N_4939,N_4800);
and UO_863 (O_863,N_4836,N_4843);
or UO_864 (O_864,N_4922,N_4928);
nor UO_865 (O_865,N_4929,N_4899);
nor UO_866 (O_866,N_4887,N_4904);
and UO_867 (O_867,N_4913,N_4910);
and UO_868 (O_868,N_4859,N_4854);
and UO_869 (O_869,N_4864,N_4858);
and UO_870 (O_870,N_4839,N_4965);
and UO_871 (O_871,N_4947,N_4810);
and UO_872 (O_872,N_4895,N_4999);
nor UO_873 (O_873,N_4841,N_4950);
nor UO_874 (O_874,N_4857,N_4916);
nor UO_875 (O_875,N_4869,N_4867);
nor UO_876 (O_876,N_4986,N_4960);
nor UO_877 (O_877,N_4970,N_4892);
nor UO_878 (O_878,N_4850,N_4942);
nor UO_879 (O_879,N_4933,N_4843);
and UO_880 (O_880,N_4825,N_4901);
nand UO_881 (O_881,N_4830,N_4881);
and UO_882 (O_882,N_4809,N_4979);
and UO_883 (O_883,N_4932,N_4822);
or UO_884 (O_884,N_4996,N_4928);
or UO_885 (O_885,N_4857,N_4888);
or UO_886 (O_886,N_4933,N_4991);
nor UO_887 (O_887,N_4815,N_4842);
or UO_888 (O_888,N_4834,N_4986);
and UO_889 (O_889,N_4945,N_4810);
nor UO_890 (O_890,N_4879,N_4823);
and UO_891 (O_891,N_4806,N_4930);
nand UO_892 (O_892,N_4931,N_4978);
and UO_893 (O_893,N_4841,N_4842);
nand UO_894 (O_894,N_4883,N_4837);
nand UO_895 (O_895,N_4945,N_4971);
nor UO_896 (O_896,N_4975,N_4886);
and UO_897 (O_897,N_4877,N_4948);
and UO_898 (O_898,N_4845,N_4849);
and UO_899 (O_899,N_4854,N_4922);
or UO_900 (O_900,N_4854,N_4835);
or UO_901 (O_901,N_4995,N_4867);
and UO_902 (O_902,N_4901,N_4888);
nand UO_903 (O_903,N_4810,N_4953);
or UO_904 (O_904,N_4943,N_4840);
and UO_905 (O_905,N_4944,N_4925);
nor UO_906 (O_906,N_4983,N_4866);
nor UO_907 (O_907,N_4901,N_4940);
or UO_908 (O_908,N_4830,N_4908);
or UO_909 (O_909,N_4895,N_4836);
nand UO_910 (O_910,N_4839,N_4823);
and UO_911 (O_911,N_4952,N_4830);
or UO_912 (O_912,N_4904,N_4827);
and UO_913 (O_913,N_4987,N_4830);
and UO_914 (O_914,N_4919,N_4989);
and UO_915 (O_915,N_4814,N_4890);
nor UO_916 (O_916,N_4859,N_4993);
or UO_917 (O_917,N_4861,N_4896);
nand UO_918 (O_918,N_4853,N_4969);
or UO_919 (O_919,N_4870,N_4874);
nand UO_920 (O_920,N_4812,N_4961);
and UO_921 (O_921,N_4886,N_4887);
nor UO_922 (O_922,N_4831,N_4819);
and UO_923 (O_923,N_4955,N_4963);
or UO_924 (O_924,N_4900,N_4953);
nand UO_925 (O_925,N_4838,N_4895);
xnor UO_926 (O_926,N_4835,N_4966);
or UO_927 (O_927,N_4884,N_4852);
nor UO_928 (O_928,N_4913,N_4807);
nor UO_929 (O_929,N_4901,N_4993);
xnor UO_930 (O_930,N_4856,N_4811);
or UO_931 (O_931,N_4888,N_4980);
nor UO_932 (O_932,N_4879,N_4839);
nor UO_933 (O_933,N_4942,N_4983);
or UO_934 (O_934,N_4862,N_4803);
or UO_935 (O_935,N_4967,N_4896);
or UO_936 (O_936,N_4836,N_4918);
and UO_937 (O_937,N_4988,N_4819);
nor UO_938 (O_938,N_4891,N_4914);
or UO_939 (O_939,N_4896,N_4863);
or UO_940 (O_940,N_4816,N_4829);
or UO_941 (O_941,N_4851,N_4868);
and UO_942 (O_942,N_4899,N_4924);
nor UO_943 (O_943,N_4947,N_4944);
or UO_944 (O_944,N_4945,N_4956);
and UO_945 (O_945,N_4944,N_4973);
nor UO_946 (O_946,N_4912,N_4983);
or UO_947 (O_947,N_4837,N_4948);
nand UO_948 (O_948,N_4955,N_4812);
and UO_949 (O_949,N_4931,N_4823);
nand UO_950 (O_950,N_4828,N_4865);
nand UO_951 (O_951,N_4872,N_4810);
and UO_952 (O_952,N_4819,N_4973);
nand UO_953 (O_953,N_4857,N_4903);
nand UO_954 (O_954,N_4998,N_4985);
or UO_955 (O_955,N_4863,N_4969);
or UO_956 (O_956,N_4930,N_4978);
nand UO_957 (O_957,N_4886,N_4965);
nor UO_958 (O_958,N_4986,N_4809);
and UO_959 (O_959,N_4882,N_4968);
or UO_960 (O_960,N_4910,N_4856);
nor UO_961 (O_961,N_4891,N_4876);
nand UO_962 (O_962,N_4826,N_4818);
nand UO_963 (O_963,N_4922,N_4917);
or UO_964 (O_964,N_4975,N_4817);
and UO_965 (O_965,N_4805,N_4905);
and UO_966 (O_966,N_4903,N_4836);
nor UO_967 (O_967,N_4843,N_4977);
and UO_968 (O_968,N_4907,N_4942);
or UO_969 (O_969,N_4935,N_4906);
nor UO_970 (O_970,N_4862,N_4856);
and UO_971 (O_971,N_4902,N_4934);
and UO_972 (O_972,N_4887,N_4865);
nor UO_973 (O_973,N_4988,N_4826);
or UO_974 (O_974,N_4810,N_4912);
or UO_975 (O_975,N_4810,N_4959);
or UO_976 (O_976,N_4976,N_4962);
or UO_977 (O_977,N_4955,N_4981);
nor UO_978 (O_978,N_4903,N_4804);
nor UO_979 (O_979,N_4882,N_4975);
nand UO_980 (O_980,N_4967,N_4985);
and UO_981 (O_981,N_4955,N_4818);
and UO_982 (O_982,N_4841,N_4817);
nand UO_983 (O_983,N_4993,N_4964);
nor UO_984 (O_984,N_4800,N_4965);
or UO_985 (O_985,N_4851,N_4872);
nand UO_986 (O_986,N_4847,N_4947);
nor UO_987 (O_987,N_4814,N_4919);
nor UO_988 (O_988,N_4914,N_4894);
and UO_989 (O_989,N_4811,N_4876);
and UO_990 (O_990,N_4899,N_4848);
or UO_991 (O_991,N_4810,N_4865);
or UO_992 (O_992,N_4896,N_4955);
or UO_993 (O_993,N_4947,N_4898);
or UO_994 (O_994,N_4979,N_4953);
nor UO_995 (O_995,N_4919,N_4816);
or UO_996 (O_996,N_4964,N_4958);
and UO_997 (O_997,N_4915,N_4938);
xnor UO_998 (O_998,N_4958,N_4981);
or UO_999 (O_999,N_4970,N_4967);
endmodule