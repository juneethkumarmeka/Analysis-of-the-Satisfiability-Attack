module basic_500_3000_500_5_levels_5xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
and U0 (N_0,In_72,In_304);
or U1 (N_1,In_240,In_161);
or U2 (N_2,In_276,In_329);
nor U3 (N_3,In_208,In_33);
and U4 (N_4,In_20,In_222);
nand U5 (N_5,In_189,In_124);
nand U6 (N_6,In_285,In_256);
and U7 (N_7,In_365,In_363);
and U8 (N_8,In_235,In_19);
xor U9 (N_9,In_242,In_300);
nor U10 (N_10,In_482,In_224);
nor U11 (N_11,In_466,In_200);
or U12 (N_12,In_445,In_175);
xor U13 (N_13,In_491,In_112);
or U14 (N_14,In_23,In_195);
nor U15 (N_15,In_361,In_347);
nand U16 (N_16,In_486,In_31);
nand U17 (N_17,In_36,In_144);
xor U18 (N_18,In_54,In_318);
nand U19 (N_19,In_215,In_150);
and U20 (N_20,In_245,In_310);
nand U21 (N_21,In_132,In_472);
and U22 (N_22,In_226,In_1);
xor U23 (N_23,In_87,In_314);
and U24 (N_24,In_77,In_18);
and U25 (N_25,In_375,In_293);
and U26 (N_26,In_266,In_225);
or U27 (N_27,In_156,In_71);
or U28 (N_28,In_194,In_414);
nor U29 (N_29,In_191,In_349);
xnor U30 (N_30,In_313,In_163);
or U31 (N_31,In_320,In_452);
or U32 (N_32,In_86,In_436);
nor U33 (N_33,In_151,In_419);
nand U34 (N_34,In_32,In_0);
nor U35 (N_35,In_416,In_169);
and U36 (N_36,In_38,In_61);
nor U37 (N_37,In_427,In_186);
and U38 (N_38,In_400,In_387);
or U39 (N_39,In_442,In_223);
or U40 (N_40,In_483,In_360);
and U41 (N_41,In_115,In_160);
or U42 (N_42,In_253,In_37);
or U43 (N_43,In_475,In_214);
xor U44 (N_44,In_155,In_312);
nand U45 (N_45,In_455,In_460);
nor U46 (N_46,In_2,In_233);
or U47 (N_47,In_393,In_89);
or U48 (N_48,In_465,In_389);
nor U49 (N_49,In_342,In_481);
nand U50 (N_50,In_283,In_88);
and U51 (N_51,In_325,In_463);
or U52 (N_52,In_426,In_364);
nor U53 (N_53,In_410,In_492);
and U54 (N_54,In_374,In_476);
xor U55 (N_55,In_392,In_309);
or U56 (N_56,In_372,In_211);
nor U57 (N_57,In_243,In_430);
nor U58 (N_58,In_95,In_141);
xnor U59 (N_59,In_181,In_384);
nor U60 (N_60,In_143,In_92);
nor U61 (N_61,In_179,In_46);
and U62 (N_62,In_265,In_294);
and U63 (N_63,In_47,In_288);
xor U64 (N_64,In_129,In_403);
nand U65 (N_65,In_485,In_434);
and U66 (N_66,In_447,In_290);
nand U67 (N_67,In_284,In_353);
and U68 (N_68,In_27,In_296);
or U69 (N_69,In_127,In_108);
nand U70 (N_70,In_496,In_78);
nor U71 (N_71,In_74,In_148);
nor U72 (N_72,In_474,In_76);
or U73 (N_73,In_10,In_321);
nand U74 (N_74,In_450,In_12);
and U75 (N_75,In_324,In_136);
and U76 (N_76,In_187,In_261);
nor U77 (N_77,In_118,In_173);
nand U78 (N_78,In_66,In_446);
nand U79 (N_79,In_70,In_339);
xnor U80 (N_80,In_272,In_238);
nand U81 (N_81,In_107,In_84);
or U82 (N_82,In_332,In_103);
xnor U83 (N_83,In_139,In_221);
and U84 (N_84,In_282,In_281);
nor U85 (N_85,In_286,In_149);
or U86 (N_86,In_316,In_145);
xor U87 (N_87,In_473,In_184);
nor U88 (N_88,In_373,In_58);
nand U89 (N_89,In_159,In_16);
nand U90 (N_90,In_154,In_13);
xor U91 (N_91,In_75,In_448);
xor U92 (N_92,In_254,In_165);
xor U93 (N_93,In_96,In_303);
and U94 (N_94,In_461,In_362);
nand U95 (N_95,In_152,In_93);
nor U96 (N_96,In_390,In_62);
nor U97 (N_97,In_97,In_153);
xnor U98 (N_98,In_119,In_458);
nor U99 (N_99,In_326,In_269);
nor U100 (N_100,In_172,In_106);
or U101 (N_101,In_22,In_428);
nand U102 (N_102,In_415,In_30);
or U103 (N_103,In_57,In_134);
xor U104 (N_104,In_383,In_126);
or U105 (N_105,In_157,In_292);
nor U106 (N_106,In_228,In_6);
nand U107 (N_107,In_203,In_246);
xnor U108 (N_108,In_192,In_470);
nor U109 (N_109,In_82,In_91);
nor U110 (N_110,In_3,In_454);
nand U111 (N_111,In_83,In_80);
nand U112 (N_112,In_176,In_327);
xnor U113 (N_113,In_344,In_111);
and U114 (N_114,In_397,In_401);
or U115 (N_115,In_110,In_263);
and U116 (N_116,In_378,In_366);
or U117 (N_117,In_123,In_357);
and U118 (N_118,In_178,In_412);
and U119 (N_119,In_398,In_449);
nor U120 (N_120,In_291,In_217);
nand U121 (N_121,In_319,In_407);
nor U122 (N_122,In_333,In_437);
nand U123 (N_123,In_56,In_443);
or U124 (N_124,In_202,In_386);
or U125 (N_125,In_425,In_274);
and U126 (N_126,In_255,In_212);
nand U127 (N_127,In_370,In_188);
and U128 (N_128,In_494,In_498);
nor U129 (N_129,In_408,In_190);
and U130 (N_130,In_248,In_244);
nor U131 (N_131,In_51,In_69);
and U132 (N_132,In_423,In_346);
or U133 (N_133,In_354,In_17);
nand U134 (N_134,In_369,In_34);
nand U135 (N_135,In_8,In_334);
xor U136 (N_136,In_499,In_268);
or U137 (N_137,In_59,In_241);
nor U138 (N_138,In_424,In_236);
nor U139 (N_139,In_411,In_101);
nand U140 (N_140,In_478,In_413);
and U141 (N_141,In_338,In_125);
or U142 (N_142,In_488,In_120);
nand U143 (N_143,In_99,In_52);
nor U144 (N_144,In_230,In_198);
or U145 (N_145,In_121,In_402);
xnor U146 (N_146,In_444,In_468);
nor U147 (N_147,In_171,In_5);
xnor U148 (N_148,In_49,In_193);
nand U149 (N_149,In_182,In_297);
nor U150 (N_150,In_94,In_438);
or U151 (N_151,In_201,In_337);
and U152 (N_152,In_409,In_270);
and U153 (N_153,In_429,In_381);
xor U154 (N_154,In_260,In_133);
and U155 (N_155,In_180,In_376);
nand U156 (N_156,In_64,In_439);
nand U157 (N_157,In_469,In_41);
nand U158 (N_158,In_382,In_116);
nor U159 (N_159,In_128,In_250);
xor U160 (N_160,In_7,In_11);
or U161 (N_161,In_462,In_258);
nand U162 (N_162,In_307,In_495);
nor U163 (N_163,In_48,In_207);
and U164 (N_164,In_67,In_391);
xnor U165 (N_165,In_231,In_278);
or U166 (N_166,In_251,In_335);
and U167 (N_167,In_350,In_453);
and U168 (N_168,In_113,In_451);
nand U169 (N_169,In_218,In_493);
or U170 (N_170,In_237,In_287);
or U171 (N_171,In_90,In_114);
and U172 (N_172,In_205,In_177);
or U173 (N_173,In_50,In_273);
nand U174 (N_174,In_480,In_45);
or U175 (N_175,In_262,In_341);
and U176 (N_176,In_359,In_388);
or U177 (N_177,In_355,In_167);
and U178 (N_178,In_317,In_417);
and U179 (N_179,In_247,In_305);
xnor U180 (N_180,In_39,In_24);
nor U181 (N_181,In_239,In_396);
nand U182 (N_182,In_209,In_497);
nor U183 (N_183,In_323,In_25);
nand U184 (N_184,In_252,In_328);
nor U185 (N_185,In_422,In_348);
or U186 (N_186,In_371,In_102);
xor U187 (N_187,In_395,In_138);
or U188 (N_188,In_213,In_351);
nor U189 (N_189,In_441,In_131);
and U190 (N_190,In_234,In_477);
nand U191 (N_191,In_140,In_35);
nor U192 (N_192,In_220,In_279);
or U193 (N_193,In_68,In_368);
nor U194 (N_194,In_367,In_289);
xnor U195 (N_195,In_166,In_170);
or U196 (N_196,In_196,In_162);
and U197 (N_197,In_487,In_330);
or U198 (N_198,In_204,In_142);
nand U199 (N_199,In_264,In_104);
and U200 (N_200,In_26,In_277);
nand U201 (N_201,In_85,In_40);
and U202 (N_202,In_385,In_394);
or U203 (N_203,In_440,In_168);
nand U204 (N_204,In_405,In_60);
or U205 (N_205,In_421,In_356);
and U206 (N_206,In_122,In_216);
and U207 (N_207,In_479,In_280);
xor U208 (N_208,In_433,In_147);
and U209 (N_209,In_15,In_105);
or U210 (N_210,In_406,In_358);
and U211 (N_211,In_28,In_315);
xnor U212 (N_212,In_267,In_399);
or U213 (N_213,In_295,In_44);
nor U214 (N_214,In_467,In_4);
nand U215 (N_215,In_459,In_275);
and U216 (N_216,In_43,In_21);
nand U217 (N_217,In_206,In_302);
and U218 (N_218,In_489,In_457);
nand U219 (N_219,In_471,In_352);
and U220 (N_220,In_299,In_55);
nand U221 (N_221,In_301,In_298);
and U222 (N_222,In_183,In_229);
xnor U223 (N_223,In_29,In_185);
and U224 (N_224,In_199,In_232);
and U225 (N_225,In_63,In_484);
xor U226 (N_226,In_73,In_79);
or U227 (N_227,In_9,In_174);
and U228 (N_228,In_100,In_257);
or U229 (N_229,In_490,In_81);
nand U230 (N_230,In_331,In_117);
nand U231 (N_231,In_53,In_380);
nor U232 (N_232,In_432,In_271);
and U233 (N_233,In_137,In_130);
nor U234 (N_234,In_377,In_249);
nor U235 (N_235,In_210,In_308);
nor U236 (N_236,In_464,In_109);
and U237 (N_237,In_42,In_379);
or U238 (N_238,In_158,In_197);
and U239 (N_239,In_404,In_135);
xor U240 (N_240,In_345,In_227);
or U241 (N_241,In_259,In_420);
or U242 (N_242,In_311,In_340);
nor U243 (N_243,In_98,In_306);
or U244 (N_244,In_456,In_65);
nand U245 (N_245,In_418,In_164);
and U246 (N_246,In_336,In_146);
or U247 (N_247,In_322,In_219);
xor U248 (N_248,In_343,In_14);
nand U249 (N_249,In_431,In_435);
nand U250 (N_250,In_385,In_329);
nand U251 (N_251,In_321,In_289);
xor U252 (N_252,In_219,In_303);
or U253 (N_253,In_407,In_83);
and U254 (N_254,In_125,In_436);
nand U255 (N_255,In_442,In_46);
nor U256 (N_256,In_61,In_229);
nand U257 (N_257,In_387,In_468);
nor U258 (N_258,In_124,In_24);
or U259 (N_259,In_475,In_399);
and U260 (N_260,In_249,In_178);
nand U261 (N_261,In_241,In_193);
nor U262 (N_262,In_410,In_188);
xnor U263 (N_263,In_7,In_116);
nor U264 (N_264,In_306,In_316);
or U265 (N_265,In_79,In_206);
nand U266 (N_266,In_59,In_42);
or U267 (N_267,In_383,In_15);
and U268 (N_268,In_110,In_492);
nor U269 (N_269,In_363,In_53);
or U270 (N_270,In_392,In_284);
or U271 (N_271,In_373,In_439);
or U272 (N_272,In_268,In_449);
nor U273 (N_273,In_138,In_489);
nor U274 (N_274,In_374,In_159);
and U275 (N_275,In_161,In_468);
and U276 (N_276,In_483,In_27);
or U277 (N_277,In_365,In_132);
and U278 (N_278,In_240,In_481);
xor U279 (N_279,In_9,In_232);
or U280 (N_280,In_173,In_17);
nand U281 (N_281,In_361,In_11);
nor U282 (N_282,In_102,In_437);
nand U283 (N_283,In_409,In_250);
or U284 (N_284,In_415,In_8);
xnor U285 (N_285,In_123,In_111);
xor U286 (N_286,In_472,In_442);
xnor U287 (N_287,In_10,In_263);
nor U288 (N_288,In_251,In_108);
or U289 (N_289,In_464,In_235);
and U290 (N_290,In_82,In_164);
and U291 (N_291,In_18,In_491);
or U292 (N_292,In_419,In_249);
nand U293 (N_293,In_367,In_243);
nand U294 (N_294,In_252,In_313);
nand U295 (N_295,In_271,In_324);
nor U296 (N_296,In_346,In_15);
nand U297 (N_297,In_207,In_260);
nor U298 (N_298,In_289,In_264);
and U299 (N_299,In_374,In_44);
and U300 (N_300,In_354,In_292);
or U301 (N_301,In_118,In_255);
and U302 (N_302,In_435,In_199);
or U303 (N_303,In_137,In_224);
nor U304 (N_304,In_240,In_475);
nor U305 (N_305,In_193,In_52);
nand U306 (N_306,In_89,In_60);
nand U307 (N_307,In_491,In_366);
and U308 (N_308,In_222,In_384);
or U309 (N_309,In_177,In_139);
and U310 (N_310,In_307,In_463);
and U311 (N_311,In_226,In_205);
nor U312 (N_312,In_52,In_215);
or U313 (N_313,In_61,In_275);
nor U314 (N_314,In_467,In_354);
xor U315 (N_315,In_130,In_49);
nor U316 (N_316,In_376,In_431);
xor U317 (N_317,In_355,In_219);
xor U318 (N_318,In_193,In_454);
and U319 (N_319,In_93,In_22);
or U320 (N_320,In_67,In_101);
nand U321 (N_321,In_276,In_110);
nor U322 (N_322,In_176,In_302);
nor U323 (N_323,In_14,In_154);
and U324 (N_324,In_87,In_254);
xnor U325 (N_325,In_372,In_385);
or U326 (N_326,In_479,In_342);
nor U327 (N_327,In_105,In_471);
or U328 (N_328,In_86,In_186);
xnor U329 (N_329,In_315,In_470);
nand U330 (N_330,In_49,In_368);
nand U331 (N_331,In_43,In_196);
and U332 (N_332,In_250,In_100);
or U333 (N_333,In_385,In_125);
or U334 (N_334,In_123,In_352);
or U335 (N_335,In_53,In_247);
nor U336 (N_336,In_214,In_228);
xor U337 (N_337,In_159,In_49);
xnor U338 (N_338,In_124,In_180);
xor U339 (N_339,In_304,In_270);
nand U340 (N_340,In_463,In_383);
or U341 (N_341,In_138,In_485);
nor U342 (N_342,In_343,In_191);
nand U343 (N_343,In_469,In_204);
and U344 (N_344,In_290,In_432);
nand U345 (N_345,In_170,In_253);
xor U346 (N_346,In_469,In_18);
or U347 (N_347,In_159,In_443);
nor U348 (N_348,In_433,In_392);
or U349 (N_349,In_104,In_41);
or U350 (N_350,In_280,In_320);
nor U351 (N_351,In_216,In_451);
xnor U352 (N_352,In_373,In_486);
or U353 (N_353,In_204,In_201);
or U354 (N_354,In_232,In_163);
and U355 (N_355,In_106,In_385);
and U356 (N_356,In_353,In_46);
nor U357 (N_357,In_450,In_91);
nor U358 (N_358,In_95,In_436);
nand U359 (N_359,In_331,In_158);
nand U360 (N_360,In_150,In_483);
nand U361 (N_361,In_426,In_97);
or U362 (N_362,In_425,In_358);
or U363 (N_363,In_428,In_131);
nor U364 (N_364,In_223,In_302);
or U365 (N_365,In_58,In_352);
and U366 (N_366,In_348,In_28);
or U367 (N_367,In_418,In_392);
nand U368 (N_368,In_486,In_484);
and U369 (N_369,In_97,In_197);
or U370 (N_370,In_339,In_461);
or U371 (N_371,In_452,In_330);
nand U372 (N_372,In_371,In_209);
nor U373 (N_373,In_374,In_263);
xnor U374 (N_374,In_1,In_492);
or U375 (N_375,In_409,In_392);
nand U376 (N_376,In_211,In_200);
and U377 (N_377,In_278,In_369);
nand U378 (N_378,In_498,In_343);
or U379 (N_379,In_447,In_185);
or U380 (N_380,In_254,In_285);
and U381 (N_381,In_1,In_369);
nand U382 (N_382,In_12,In_255);
nor U383 (N_383,In_105,In_21);
or U384 (N_384,In_33,In_321);
and U385 (N_385,In_287,In_393);
nor U386 (N_386,In_381,In_33);
or U387 (N_387,In_289,In_434);
or U388 (N_388,In_114,In_7);
and U389 (N_389,In_436,In_443);
nor U390 (N_390,In_372,In_328);
nor U391 (N_391,In_452,In_286);
and U392 (N_392,In_126,In_490);
nand U393 (N_393,In_93,In_100);
and U394 (N_394,In_438,In_351);
or U395 (N_395,In_13,In_487);
nor U396 (N_396,In_27,In_124);
and U397 (N_397,In_190,In_428);
nor U398 (N_398,In_360,In_17);
nand U399 (N_399,In_272,In_322);
or U400 (N_400,In_314,In_101);
and U401 (N_401,In_298,In_391);
and U402 (N_402,In_319,In_51);
nand U403 (N_403,In_46,In_93);
and U404 (N_404,In_431,In_426);
or U405 (N_405,In_120,In_324);
nand U406 (N_406,In_219,In_426);
nand U407 (N_407,In_219,In_309);
nor U408 (N_408,In_321,In_498);
and U409 (N_409,In_64,In_218);
xnor U410 (N_410,In_134,In_469);
nor U411 (N_411,In_357,In_61);
and U412 (N_412,In_89,In_133);
nand U413 (N_413,In_305,In_164);
xnor U414 (N_414,In_12,In_207);
nor U415 (N_415,In_214,In_394);
nor U416 (N_416,In_118,In_77);
and U417 (N_417,In_119,In_378);
or U418 (N_418,In_396,In_401);
nand U419 (N_419,In_67,In_242);
nor U420 (N_420,In_225,In_119);
or U421 (N_421,In_297,In_299);
and U422 (N_422,In_375,In_117);
xor U423 (N_423,In_266,In_86);
and U424 (N_424,In_472,In_391);
or U425 (N_425,In_248,In_464);
or U426 (N_426,In_462,In_202);
and U427 (N_427,In_57,In_261);
nand U428 (N_428,In_110,In_488);
nor U429 (N_429,In_432,In_140);
nand U430 (N_430,In_45,In_481);
or U431 (N_431,In_58,In_114);
nand U432 (N_432,In_54,In_156);
nand U433 (N_433,In_229,In_17);
nand U434 (N_434,In_176,In_484);
nor U435 (N_435,In_497,In_177);
or U436 (N_436,In_409,In_249);
nor U437 (N_437,In_279,In_96);
or U438 (N_438,In_256,In_434);
and U439 (N_439,In_159,In_46);
xnor U440 (N_440,In_410,In_119);
nor U441 (N_441,In_198,In_73);
nand U442 (N_442,In_296,In_226);
or U443 (N_443,In_18,In_303);
or U444 (N_444,In_38,In_104);
xor U445 (N_445,In_132,In_373);
nor U446 (N_446,In_71,In_384);
nand U447 (N_447,In_402,In_78);
nand U448 (N_448,In_376,In_241);
nor U449 (N_449,In_244,In_411);
nand U450 (N_450,In_396,In_83);
nand U451 (N_451,In_406,In_166);
nor U452 (N_452,In_460,In_180);
and U453 (N_453,In_144,In_350);
or U454 (N_454,In_218,In_455);
nand U455 (N_455,In_370,In_423);
nor U456 (N_456,In_89,In_48);
or U457 (N_457,In_38,In_110);
nand U458 (N_458,In_178,In_201);
and U459 (N_459,In_45,In_288);
nand U460 (N_460,In_450,In_494);
or U461 (N_461,In_271,In_477);
nand U462 (N_462,In_437,In_159);
nor U463 (N_463,In_140,In_409);
and U464 (N_464,In_143,In_456);
or U465 (N_465,In_91,In_306);
nor U466 (N_466,In_175,In_438);
nor U467 (N_467,In_316,In_451);
and U468 (N_468,In_429,In_473);
or U469 (N_469,In_422,In_115);
nand U470 (N_470,In_473,In_312);
and U471 (N_471,In_118,In_288);
and U472 (N_472,In_493,In_128);
or U473 (N_473,In_282,In_376);
or U474 (N_474,In_336,In_245);
and U475 (N_475,In_413,In_177);
nor U476 (N_476,In_343,In_254);
nor U477 (N_477,In_129,In_364);
nor U478 (N_478,In_305,In_393);
xnor U479 (N_479,In_231,In_46);
nand U480 (N_480,In_98,In_139);
or U481 (N_481,In_423,In_218);
and U482 (N_482,In_70,In_116);
nand U483 (N_483,In_272,In_383);
nor U484 (N_484,In_405,In_36);
nor U485 (N_485,In_488,In_173);
nor U486 (N_486,In_17,In_85);
nand U487 (N_487,In_361,In_57);
and U488 (N_488,In_246,In_17);
or U489 (N_489,In_421,In_18);
and U490 (N_490,In_118,In_7);
xnor U491 (N_491,In_80,In_428);
or U492 (N_492,In_335,In_145);
or U493 (N_493,In_272,In_194);
or U494 (N_494,In_220,In_436);
or U495 (N_495,In_310,In_341);
nor U496 (N_496,In_153,In_335);
or U497 (N_497,In_441,In_142);
xor U498 (N_498,In_483,In_47);
or U499 (N_499,In_293,In_161);
or U500 (N_500,In_157,In_62);
nor U501 (N_501,In_284,In_148);
or U502 (N_502,In_319,In_178);
or U503 (N_503,In_110,In_268);
and U504 (N_504,In_107,In_471);
and U505 (N_505,In_197,In_201);
or U506 (N_506,In_376,In_469);
and U507 (N_507,In_100,In_66);
and U508 (N_508,In_399,In_72);
nand U509 (N_509,In_480,In_468);
nor U510 (N_510,In_383,In_283);
nand U511 (N_511,In_344,In_274);
nand U512 (N_512,In_279,In_264);
or U513 (N_513,In_155,In_217);
or U514 (N_514,In_347,In_401);
and U515 (N_515,In_108,In_244);
and U516 (N_516,In_313,In_415);
nor U517 (N_517,In_298,In_168);
or U518 (N_518,In_343,In_478);
and U519 (N_519,In_9,In_124);
nor U520 (N_520,In_339,In_59);
nor U521 (N_521,In_58,In_47);
nand U522 (N_522,In_143,In_237);
and U523 (N_523,In_417,In_26);
nand U524 (N_524,In_258,In_414);
and U525 (N_525,In_99,In_341);
nand U526 (N_526,In_386,In_372);
xor U527 (N_527,In_147,In_484);
and U528 (N_528,In_374,In_52);
or U529 (N_529,In_297,In_253);
nor U530 (N_530,In_288,In_46);
nand U531 (N_531,In_411,In_293);
nor U532 (N_532,In_443,In_232);
nor U533 (N_533,In_354,In_461);
nor U534 (N_534,In_221,In_28);
and U535 (N_535,In_66,In_445);
nand U536 (N_536,In_139,In_211);
nand U537 (N_537,In_358,In_492);
nand U538 (N_538,In_385,In_140);
and U539 (N_539,In_164,In_106);
xnor U540 (N_540,In_208,In_156);
or U541 (N_541,In_178,In_270);
nor U542 (N_542,In_125,In_380);
and U543 (N_543,In_41,In_20);
nand U544 (N_544,In_230,In_231);
nand U545 (N_545,In_171,In_196);
nand U546 (N_546,In_204,In_484);
and U547 (N_547,In_424,In_166);
xnor U548 (N_548,In_389,In_341);
nor U549 (N_549,In_352,In_458);
or U550 (N_550,In_251,In_492);
or U551 (N_551,In_115,In_132);
nand U552 (N_552,In_218,In_324);
nand U553 (N_553,In_446,In_428);
and U554 (N_554,In_276,In_315);
nor U555 (N_555,In_198,In_194);
nand U556 (N_556,In_191,In_229);
and U557 (N_557,In_364,In_434);
nand U558 (N_558,In_309,In_491);
nand U559 (N_559,In_417,In_173);
or U560 (N_560,In_371,In_369);
nand U561 (N_561,In_12,In_200);
nor U562 (N_562,In_431,In_437);
or U563 (N_563,In_416,In_260);
or U564 (N_564,In_472,In_445);
nor U565 (N_565,In_343,In_438);
nor U566 (N_566,In_237,In_404);
nor U567 (N_567,In_102,In_65);
nand U568 (N_568,In_212,In_104);
nor U569 (N_569,In_60,In_419);
and U570 (N_570,In_243,In_70);
and U571 (N_571,In_369,In_68);
or U572 (N_572,In_157,In_366);
nand U573 (N_573,In_318,In_200);
nand U574 (N_574,In_435,In_49);
and U575 (N_575,In_8,In_301);
nand U576 (N_576,In_444,In_467);
nor U577 (N_577,In_250,In_398);
nand U578 (N_578,In_309,In_124);
and U579 (N_579,In_443,In_293);
or U580 (N_580,In_179,In_24);
nor U581 (N_581,In_18,In_92);
or U582 (N_582,In_219,In_380);
nand U583 (N_583,In_397,In_315);
or U584 (N_584,In_109,In_278);
xor U585 (N_585,In_433,In_344);
and U586 (N_586,In_28,In_20);
or U587 (N_587,In_210,In_416);
nor U588 (N_588,In_466,In_416);
and U589 (N_589,In_350,In_58);
xor U590 (N_590,In_466,In_366);
nand U591 (N_591,In_403,In_292);
or U592 (N_592,In_88,In_67);
or U593 (N_593,In_361,In_491);
nand U594 (N_594,In_0,In_21);
nor U595 (N_595,In_431,In_379);
or U596 (N_596,In_487,In_436);
and U597 (N_597,In_387,In_399);
nand U598 (N_598,In_48,In_250);
nor U599 (N_599,In_72,In_230);
and U600 (N_600,N_475,N_47);
nor U601 (N_601,N_596,N_310);
nand U602 (N_602,N_559,N_248);
xnor U603 (N_603,N_593,N_374);
nor U604 (N_604,N_576,N_136);
nand U605 (N_605,N_105,N_404);
and U606 (N_606,N_480,N_431);
xor U607 (N_607,N_500,N_443);
and U608 (N_608,N_181,N_70);
or U609 (N_609,N_81,N_25);
nand U610 (N_610,N_53,N_71);
nor U611 (N_611,N_396,N_352);
and U612 (N_612,N_377,N_376);
nand U613 (N_613,N_472,N_92);
or U614 (N_614,N_27,N_38);
xor U615 (N_615,N_95,N_242);
nand U616 (N_616,N_183,N_291);
or U617 (N_617,N_501,N_348);
xnor U618 (N_618,N_8,N_147);
nor U619 (N_619,N_524,N_278);
nor U620 (N_620,N_196,N_355);
nor U621 (N_621,N_343,N_563);
and U622 (N_622,N_178,N_63);
and U623 (N_623,N_329,N_406);
and U624 (N_624,N_438,N_32);
and U625 (N_625,N_11,N_362);
nor U626 (N_626,N_201,N_499);
and U627 (N_627,N_36,N_79);
nand U628 (N_628,N_179,N_280);
and U629 (N_629,N_244,N_3);
and U630 (N_630,N_544,N_204);
nor U631 (N_631,N_307,N_508);
nand U632 (N_632,N_270,N_447);
xnor U633 (N_633,N_83,N_535);
or U634 (N_634,N_461,N_494);
nor U635 (N_635,N_65,N_262);
nand U636 (N_636,N_393,N_102);
xor U637 (N_637,N_314,N_211);
nor U638 (N_638,N_290,N_429);
nor U639 (N_639,N_209,N_552);
nor U640 (N_640,N_113,N_23);
or U641 (N_641,N_569,N_311);
nor U642 (N_642,N_582,N_5);
nor U643 (N_643,N_556,N_542);
nand U644 (N_644,N_571,N_579);
and U645 (N_645,N_149,N_325);
nand U646 (N_646,N_573,N_442);
and U647 (N_647,N_89,N_152);
nor U648 (N_648,N_111,N_331);
nand U649 (N_649,N_309,N_434);
nor U650 (N_650,N_564,N_586);
nor U651 (N_651,N_203,N_483);
nand U652 (N_652,N_52,N_509);
nand U653 (N_653,N_441,N_505);
nor U654 (N_654,N_220,N_567);
or U655 (N_655,N_444,N_91);
or U656 (N_656,N_534,N_546);
and U657 (N_657,N_421,N_344);
or U658 (N_658,N_96,N_504);
or U659 (N_659,N_14,N_24);
and U660 (N_660,N_550,N_0);
nor U661 (N_661,N_540,N_389);
or U662 (N_662,N_296,N_361);
or U663 (N_663,N_386,N_163);
nor U664 (N_664,N_265,N_455);
and U665 (N_665,N_492,N_510);
nand U666 (N_666,N_12,N_251);
and U667 (N_667,N_557,N_336);
xor U668 (N_668,N_46,N_541);
nor U669 (N_669,N_299,N_536);
or U670 (N_670,N_525,N_590);
nand U671 (N_671,N_380,N_597);
nand U672 (N_672,N_7,N_485);
and U673 (N_673,N_212,N_319);
nor U674 (N_674,N_587,N_538);
nand U675 (N_675,N_200,N_195);
or U676 (N_676,N_435,N_498);
or U677 (N_677,N_519,N_450);
nand U678 (N_678,N_22,N_130);
xor U679 (N_679,N_263,N_378);
and U680 (N_680,N_335,N_40);
or U681 (N_681,N_594,N_156);
nand U682 (N_682,N_295,N_10);
and U683 (N_683,N_543,N_381);
nand U684 (N_684,N_428,N_160);
or U685 (N_685,N_437,N_107);
nand U686 (N_686,N_529,N_155);
nor U687 (N_687,N_384,N_301);
nor U688 (N_688,N_315,N_80);
or U689 (N_689,N_109,N_60);
xnor U690 (N_690,N_229,N_144);
or U691 (N_691,N_560,N_74);
nand U692 (N_692,N_385,N_93);
nand U693 (N_693,N_253,N_207);
nand U694 (N_694,N_140,N_572);
nand U695 (N_695,N_148,N_375);
and U696 (N_696,N_436,N_240);
and U697 (N_697,N_390,N_527);
or U698 (N_698,N_566,N_82);
nor U699 (N_699,N_418,N_31);
nand U700 (N_700,N_121,N_45);
nor U701 (N_701,N_448,N_387);
nor U702 (N_702,N_139,N_339);
nand U703 (N_703,N_129,N_415);
nand U704 (N_704,N_119,N_231);
or U705 (N_705,N_164,N_513);
nand U706 (N_706,N_512,N_407);
nor U707 (N_707,N_128,N_249);
and U708 (N_708,N_427,N_324);
or U709 (N_709,N_146,N_454);
and U710 (N_710,N_135,N_106);
and U711 (N_711,N_250,N_49);
nand U712 (N_712,N_408,N_370);
nand U713 (N_713,N_167,N_59);
and U714 (N_714,N_16,N_267);
nor U715 (N_715,N_176,N_273);
or U716 (N_716,N_172,N_489);
and U717 (N_717,N_580,N_180);
and U718 (N_718,N_277,N_177);
xnor U719 (N_719,N_402,N_462);
and U720 (N_720,N_410,N_112);
and U721 (N_721,N_15,N_491);
and U722 (N_722,N_19,N_162);
or U723 (N_723,N_482,N_157);
nor U724 (N_724,N_574,N_116);
nor U725 (N_725,N_514,N_279);
xor U726 (N_726,N_161,N_391);
and U727 (N_727,N_39,N_218);
nand U728 (N_728,N_409,N_320);
and U729 (N_729,N_232,N_2);
and U730 (N_730,N_188,N_292);
nor U731 (N_731,N_479,N_284);
nand U732 (N_732,N_506,N_581);
or U733 (N_733,N_328,N_237);
and U734 (N_734,N_289,N_481);
nor U735 (N_735,N_61,N_252);
nor U736 (N_736,N_432,N_286);
and U737 (N_737,N_537,N_474);
nor U738 (N_738,N_312,N_187);
and U739 (N_739,N_397,N_145);
nand U740 (N_740,N_367,N_338);
nand U741 (N_741,N_532,N_227);
or U742 (N_742,N_401,N_118);
or U743 (N_743,N_453,N_424);
or U744 (N_744,N_342,N_142);
nor U745 (N_745,N_304,N_245);
nand U746 (N_746,N_236,N_360);
nor U747 (N_747,N_306,N_478);
and U748 (N_748,N_283,N_26);
nand U749 (N_749,N_383,N_354);
nand U750 (N_750,N_186,N_33);
nor U751 (N_751,N_457,N_568);
and U752 (N_752,N_558,N_28);
or U753 (N_753,N_426,N_549);
nand U754 (N_754,N_463,N_486);
nand U755 (N_755,N_271,N_206);
nor U756 (N_756,N_268,N_217);
and U757 (N_757,N_6,N_497);
and U758 (N_758,N_305,N_503);
or U759 (N_759,N_578,N_403);
nand U760 (N_760,N_507,N_589);
or U761 (N_761,N_465,N_371);
or U762 (N_762,N_423,N_123);
nand U763 (N_763,N_502,N_165);
or U764 (N_764,N_467,N_43);
or U765 (N_765,N_185,N_340);
xnor U766 (N_766,N_174,N_297);
nor U767 (N_767,N_205,N_517);
nand U768 (N_768,N_341,N_365);
nand U769 (N_769,N_484,N_224);
or U770 (N_770,N_228,N_565);
or U771 (N_771,N_334,N_21);
nor U772 (N_772,N_350,N_458);
or U773 (N_773,N_446,N_125);
nor U774 (N_774,N_30,N_477);
or U775 (N_775,N_235,N_199);
and U776 (N_776,N_9,N_238);
nor U777 (N_777,N_530,N_298);
and U778 (N_778,N_470,N_531);
or U779 (N_779,N_166,N_302);
nand U780 (N_780,N_54,N_192);
or U781 (N_781,N_141,N_583);
or U782 (N_782,N_98,N_269);
nor U783 (N_783,N_69,N_110);
nor U784 (N_784,N_372,N_216);
nor U785 (N_785,N_326,N_214);
nand U786 (N_786,N_158,N_193);
nor U787 (N_787,N_210,N_282);
and U788 (N_788,N_547,N_50);
and U789 (N_789,N_184,N_264);
or U790 (N_790,N_259,N_515);
and U791 (N_791,N_392,N_215);
nand U792 (N_792,N_511,N_570);
nand U793 (N_793,N_221,N_234);
nand U794 (N_794,N_420,N_132);
xor U795 (N_795,N_545,N_260);
or U796 (N_796,N_399,N_108);
xnor U797 (N_797,N_533,N_555);
or U798 (N_798,N_364,N_439);
and U799 (N_799,N_445,N_330);
nor U800 (N_800,N_133,N_41);
and U801 (N_801,N_34,N_285);
nand U802 (N_802,N_75,N_170);
and U803 (N_803,N_347,N_66);
and U804 (N_804,N_346,N_208);
and U805 (N_805,N_419,N_37);
and U806 (N_806,N_189,N_99);
and U807 (N_807,N_353,N_526);
nor U808 (N_808,N_359,N_175);
and U809 (N_809,N_395,N_363);
and U810 (N_810,N_449,N_337);
and U811 (N_811,N_464,N_78);
or U812 (N_812,N_122,N_276);
and U813 (N_813,N_520,N_86);
and U814 (N_814,N_323,N_433);
and U815 (N_815,N_57,N_588);
nor U816 (N_816,N_124,N_51);
nand U817 (N_817,N_169,N_76);
nor U818 (N_818,N_120,N_198);
nor U819 (N_819,N_230,N_261);
nor U820 (N_820,N_584,N_466);
nor U821 (N_821,N_197,N_171);
and U822 (N_822,N_523,N_321);
nor U823 (N_823,N_143,N_287);
or U824 (N_824,N_345,N_274);
nand U825 (N_825,N_190,N_562);
nand U826 (N_826,N_281,N_412);
nand U827 (N_827,N_168,N_247);
xnor U828 (N_828,N_368,N_68);
nor U829 (N_829,N_518,N_77);
nand U830 (N_830,N_351,N_539);
and U831 (N_831,N_317,N_411);
nand U832 (N_832,N_254,N_194);
nand U833 (N_833,N_90,N_528);
nand U834 (N_834,N_495,N_358);
nand U835 (N_835,N_48,N_476);
nand U836 (N_836,N_585,N_239);
or U837 (N_837,N_202,N_73);
nand U838 (N_838,N_382,N_42);
nand U839 (N_839,N_318,N_275);
xnor U840 (N_840,N_213,N_137);
nand U841 (N_841,N_561,N_488);
and U842 (N_842,N_131,N_219);
xor U843 (N_843,N_58,N_97);
or U844 (N_844,N_333,N_413);
or U845 (N_845,N_522,N_150);
nor U846 (N_846,N_496,N_551);
xor U847 (N_847,N_490,N_417);
and U848 (N_848,N_154,N_357);
or U849 (N_849,N_18,N_222);
nor U850 (N_850,N_379,N_266);
nor U851 (N_851,N_400,N_103);
and U852 (N_852,N_366,N_300);
nand U853 (N_853,N_226,N_598);
or U854 (N_854,N_575,N_1);
xor U855 (N_855,N_369,N_64);
nor U856 (N_856,N_332,N_13);
xnor U857 (N_857,N_256,N_398);
or U858 (N_858,N_592,N_294);
nor U859 (N_859,N_521,N_416);
or U860 (N_860,N_104,N_127);
and U861 (N_861,N_373,N_554);
or U862 (N_862,N_460,N_487);
or U863 (N_863,N_55,N_159);
or U864 (N_864,N_293,N_258);
nor U865 (N_865,N_303,N_272);
or U866 (N_866,N_422,N_468);
or U867 (N_867,N_313,N_233);
nor U868 (N_868,N_322,N_4);
and U869 (N_869,N_516,N_452);
or U870 (N_870,N_225,N_451);
xor U871 (N_871,N_591,N_138);
nand U872 (N_872,N_430,N_316);
or U873 (N_873,N_471,N_405);
and U874 (N_874,N_257,N_126);
nand U875 (N_875,N_115,N_29);
nand U876 (N_876,N_100,N_440);
and U877 (N_877,N_88,N_117);
nor U878 (N_878,N_553,N_548);
and U879 (N_879,N_151,N_425);
xnor U880 (N_880,N_493,N_85);
xnor U881 (N_881,N_17,N_599);
or U882 (N_882,N_473,N_577);
xnor U883 (N_883,N_72,N_191);
nand U884 (N_884,N_394,N_595);
nand U885 (N_885,N_327,N_182);
or U886 (N_886,N_44,N_56);
and U887 (N_887,N_241,N_20);
and U888 (N_888,N_414,N_246);
nor U889 (N_889,N_134,N_456);
xnor U890 (N_890,N_356,N_459);
or U891 (N_891,N_255,N_67);
and U892 (N_892,N_308,N_288);
nor U893 (N_893,N_243,N_173);
nor U894 (N_894,N_35,N_62);
nand U895 (N_895,N_84,N_94);
xnor U896 (N_896,N_349,N_223);
nand U897 (N_897,N_388,N_101);
nor U898 (N_898,N_469,N_114);
nand U899 (N_899,N_87,N_153);
nor U900 (N_900,N_253,N_188);
and U901 (N_901,N_202,N_482);
and U902 (N_902,N_445,N_64);
nor U903 (N_903,N_123,N_162);
or U904 (N_904,N_70,N_440);
or U905 (N_905,N_366,N_491);
nor U906 (N_906,N_400,N_489);
or U907 (N_907,N_529,N_231);
nand U908 (N_908,N_492,N_95);
and U909 (N_909,N_260,N_64);
nand U910 (N_910,N_329,N_224);
xnor U911 (N_911,N_250,N_587);
nand U912 (N_912,N_348,N_52);
or U913 (N_913,N_204,N_487);
or U914 (N_914,N_558,N_457);
xnor U915 (N_915,N_535,N_73);
and U916 (N_916,N_68,N_75);
xor U917 (N_917,N_216,N_317);
xor U918 (N_918,N_246,N_7);
or U919 (N_919,N_55,N_521);
and U920 (N_920,N_439,N_152);
nor U921 (N_921,N_332,N_207);
or U922 (N_922,N_13,N_157);
xor U923 (N_923,N_18,N_374);
xor U924 (N_924,N_103,N_371);
nand U925 (N_925,N_205,N_186);
nand U926 (N_926,N_447,N_246);
and U927 (N_927,N_459,N_81);
nand U928 (N_928,N_272,N_385);
or U929 (N_929,N_340,N_514);
nor U930 (N_930,N_168,N_130);
or U931 (N_931,N_297,N_372);
and U932 (N_932,N_589,N_309);
or U933 (N_933,N_336,N_265);
xnor U934 (N_934,N_385,N_501);
and U935 (N_935,N_197,N_370);
xnor U936 (N_936,N_429,N_263);
xnor U937 (N_937,N_577,N_5);
nor U938 (N_938,N_384,N_481);
xor U939 (N_939,N_212,N_468);
or U940 (N_940,N_411,N_366);
nor U941 (N_941,N_167,N_364);
and U942 (N_942,N_69,N_551);
or U943 (N_943,N_284,N_51);
nor U944 (N_944,N_115,N_99);
nand U945 (N_945,N_312,N_526);
or U946 (N_946,N_404,N_221);
or U947 (N_947,N_511,N_373);
nand U948 (N_948,N_452,N_263);
nand U949 (N_949,N_309,N_436);
nand U950 (N_950,N_564,N_369);
and U951 (N_951,N_104,N_110);
xnor U952 (N_952,N_409,N_265);
and U953 (N_953,N_296,N_466);
nand U954 (N_954,N_276,N_418);
xor U955 (N_955,N_305,N_477);
or U956 (N_956,N_319,N_520);
nor U957 (N_957,N_39,N_284);
or U958 (N_958,N_591,N_429);
xnor U959 (N_959,N_335,N_529);
nand U960 (N_960,N_140,N_354);
or U961 (N_961,N_294,N_170);
nand U962 (N_962,N_212,N_518);
or U963 (N_963,N_135,N_151);
nor U964 (N_964,N_525,N_540);
or U965 (N_965,N_514,N_244);
nand U966 (N_966,N_212,N_513);
or U967 (N_967,N_313,N_523);
and U968 (N_968,N_19,N_468);
nand U969 (N_969,N_271,N_204);
xor U970 (N_970,N_126,N_221);
or U971 (N_971,N_306,N_226);
and U972 (N_972,N_113,N_419);
and U973 (N_973,N_265,N_491);
nor U974 (N_974,N_101,N_456);
or U975 (N_975,N_8,N_181);
xor U976 (N_976,N_500,N_405);
nor U977 (N_977,N_78,N_424);
or U978 (N_978,N_442,N_366);
or U979 (N_979,N_374,N_32);
nand U980 (N_980,N_397,N_242);
xnor U981 (N_981,N_171,N_234);
and U982 (N_982,N_273,N_163);
and U983 (N_983,N_463,N_436);
or U984 (N_984,N_324,N_171);
and U985 (N_985,N_145,N_411);
nor U986 (N_986,N_26,N_101);
nand U987 (N_987,N_107,N_262);
nor U988 (N_988,N_580,N_107);
nand U989 (N_989,N_443,N_15);
xor U990 (N_990,N_167,N_263);
nor U991 (N_991,N_574,N_495);
and U992 (N_992,N_307,N_414);
and U993 (N_993,N_63,N_447);
and U994 (N_994,N_113,N_250);
nand U995 (N_995,N_3,N_129);
and U996 (N_996,N_478,N_333);
nor U997 (N_997,N_595,N_66);
nor U998 (N_998,N_23,N_350);
or U999 (N_999,N_177,N_560);
nand U1000 (N_1000,N_152,N_170);
nand U1001 (N_1001,N_576,N_558);
or U1002 (N_1002,N_355,N_188);
nand U1003 (N_1003,N_294,N_86);
and U1004 (N_1004,N_533,N_35);
and U1005 (N_1005,N_166,N_369);
or U1006 (N_1006,N_318,N_464);
nor U1007 (N_1007,N_575,N_505);
nand U1008 (N_1008,N_37,N_17);
nor U1009 (N_1009,N_577,N_137);
nor U1010 (N_1010,N_507,N_89);
nand U1011 (N_1011,N_153,N_132);
and U1012 (N_1012,N_298,N_158);
xor U1013 (N_1013,N_145,N_313);
or U1014 (N_1014,N_525,N_504);
or U1015 (N_1015,N_17,N_359);
nand U1016 (N_1016,N_485,N_19);
nand U1017 (N_1017,N_599,N_220);
and U1018 (N_1018,N_466,N_556);
and U1019 (N_1019,N_85,N_348);
or U1020 (N_1020,N_431,N_99);
and U1021 (N_1021,N_153,N_48);
or U1022 (N_1022,N_124,N_33);
nand U1023 (N_1023,N_62,N_254);
xor U1024 (N_1024,N_416,N_204);
nor U1025 (N_1025,N_473,N_85);
nand U1026 (N_1026,N_189,N_18);
nand U1027 (N_1027,N_46,N_533);
nand U1028 (N_1028,N_456,N_241);
nor U1029 (N_1029,N_523,N_373);
and U1030 (N_1030,N_263,N_227);
and U1031 (N_1031,N_365,N_515);
and U1032 (N_1032,N_504,N_139);
nand U1033 (N_1033,N_205,N_594);
and U1034 (N_1034,N_417,N_309);
and U1035 (N_1035,N_170,N_410);
nand U1036 (N_1036,N_428,N_453);
xnor U1037 (N_1037,N_586,N_323);
and U1038 (N_1038,N_494,N_518);
nand U1039 (N_1039,N_457,N_570);
xor U1040 (N_1040,N_317,N_236);
nor U1041 (N_1041,N_297,N_48);
and U1042 (N_1042,N_171,N_351);
or U1043 (N_1043,N_272,N_183);
and U1044 (N_1044,N_117,N_370);
nand U1045 (N_1045,N_23,N_76);
xor U1046 (N_1046,N_522,N_215);
nand U1047 (N_1047,N_350,N_553);
nand U1048 (N_1048,N_309,N_584);
nand U1049 (N_1049,N_238,N_592);
nand U1050 (N_1050,N_251,N_491);
xnor U1051 (N_1051,N_10,N_390);
nand U1052 (N_1052,N_3,N_329);
xor U1053 (N_1053,N_15,N_377);
and U1054 (N_1054,N_480,N_570);
nor U1055 (N_1055,N_397,N_297);
nand U1056 (N_1056,N_248,N_229);
or U1057 (N_1057,N_543,N_184);
or U1058 (N_1058,N_111,N_20);
nor U1059 (N_1059,N_207,N_584);
or U1060 (N_1060,N_150,N_272);
or U1061 (N_1061,N_230,N_302);
nor U1062 (N_1062,N_492,N_327);
or U1063 (N_1063,N_423,N_244);
and U1064 (N_1064,N_177,N_370);
nand U1065 (N_1065,N_19,N_553);
and U1066 (N_1066,N_312,N_73);
and U1067 (N_1067,N_304,N_405);
nor U1068 (N_1068,N_358,N_582);
nor U1069 (N_1069,N_265,N_128);
nor U1070 (N_1070,N_485,N_94);
nor U1071 (N_1071,N_562,N_18);
and U1072 (N_1072,N_1,N_133);
and U1073 (N_1073,N_137,N_292);
and U1074 (N_1074,N_144,N_376);
nand U1075 (N_1075,N_4,N_334);
nand U1076 (N_1076,N_101,N_465);
or U1077 (N_1077,N_94,N_316);
nor U1078 (N_1078,N_78,N_286);
or U1079 (N_1079,N_14,N_407);
xor U1080 (N_1080,N_475,N_311);
nand U1081 (N_1081,N_262,N_117);
and U1082 (N_1082,N_198,N_272);
or U1083 (N_1083,N_365,N_260);
nand U1084 (N_1084,N_585,N_572);
and U1085 (N_1085,N_92,N_559);
or U1086 (N_1086,N_260,N_281);
nand U1087 (N_1087,N_412,N_46);
xor U1088 (N_1088,N_81,N_466);
nand U1089 (N_1089,N_438,N_501);
nand U1090 (N_1090,N_231,N_7);
or U1091 (N_1091,N_134,N_131);
nand U1092 (N_1092,N_555,N_183);
and U1093 (N_1093,N_152,N_169);
and U1094 (N_1094,N_385,N_249);
and U1095 (N_1095,N_365,N_48);
nand U1096 (N_1096,N_560,N_595);
nor U1097 (N_1097,N_247,N_432);
nand U1098 (N_1098,N_593,N_424);
or U1099 (N_1099,N_545,N_399);
nand U1100 (N_1100,N_71,N_186);
or U1101 (N_1101,N_383,N_118);
xnor U1102 (N_1102,N_411,N_103);
nor U1103 (N_1103,N_498,N_363);
nor U1104 (N_1104,N_556,N_41);
nor U1105 (N_1105,N_424,N_328);
nor U1106 (N_1106,N_442,N_153);
nand U1107 (N_1107,N_514,N_35);
or U1108 (N_1108,N_134,N_566);
nor U1109 (N_1109,N_599,N_11);
nand U1110 (N_1110,N_249,N_599);
nor U1111 (N_1111,N_212,N_388);
or U1112 (N_1112,N_30,N_112);
and U1113 (N_1113,N_335,N_254);
and U1114 (N_1114,N_165,N_313);
and U1115 (N_1115,N_170,N_598);
nand U1116 (N_1116,N_63,N_548);
nand U1117 (N_1117,N_241,N_123);
nor U1118 (N_1118,N_48,N_138);
or U1119 (N_1119,N_523,N_480);
xnor U1120 (N_1120,N_467,N_501);
and U1121 (N_1121,N_397,N_286);
nor U1122 (N_1122,N_487,N_329);
nand U1123 (N_1123,N_445,N_270);
nand U1124 (N_1124,N_446,N_25);
nand U1125 (N_1125,N_506,N_299);
nand U1126 (N_1126,N_463,N_314);
and U1127 (N_1127,N_507,N_365);
nand U1128 (N_1128,N_240,N_128);
and U1129 (N_1129,N_208,N_14);
nor U1130 (N_1130,N_431,N_396);
nor U1131 (N_1131,N_277,N_361);
nor U1132 (N_1132,N_388,N_409);
nor U1133 (N_1133,N_96,N_331);
nor U1134 (N_1134,N_141,N_587);
and U1135 (N_1135,N_326,N_521);
nor U1136 (N_1136,N_568,N_168);
nand U1137 (N_1137,N_587,N_385);
nand U1138 (N_1138,N_67,N_343);
xor U1139 (N_1139,N_129,N_284);
or U1140 (N_1140,N_537,N_361);
nor U1141 (N_1141,N_112,N_229);
and U1142 (N_1142,N_186,N_580);
xnor U1143 (N_1143,N_58,N_436);
nor U1144 (N_1144,N_404,N_135);
and U1145 (N_1145,N_416,N_18);
or U1146 (N_1146,N_337,N_448);
nand U1147 (N_1147,N_248,N_456);
nand U1148 (N_1148,N_490,N_537);
nand U1149 (N_1149,N_203,N_346);
nand U1150 (N_1150,N_462,N_559);
and U1151 (N_1151,N_213,N_536);
nand U1152 (N_1152,N_575,N_328);
nor U1153 (N_1153,N_595,N_8);
or U1154 (N_1154,N_435,N_400);
or U1155 (N_1155,N_304,N_16);
nor U1156 (N_1156,N_538,N_100);
nor U1157 (N_1157,N_242,N_114);
nand U1158 (N_1158,N_135,N_318);
nor U1159 (N_1159,N_509,N_462);
or U1160 (N_1160,N_465,N_172);
or U1161 (N_1161,N_373,N_176);
xor U1162 (N_1162,N_75,N_503);
nand U1163 (N_1163,N_506,N_398);
and U1164 (N_1164,N_41,N_434);
nand U1165 (N_1165,N_491,N_272);
nand U1166 (N_1166,N_537,N_112);
or U1167 (N_1167,N_212,N_132);
and U1168 (N_1168,N_291,N_243);
and U1169 (N_1169,N_52,N_191);
nand U1170 (N_1170,N_332,N_565);
nand U1171 (N_1171,N_259,N_182);
and U1172 (N_1172,N_23,N_58);
nor U1173 (N_1173,N_450,N_576);
nor U1174 (N_1174,N_597,N_456);
or U1175 (N_1175,N_526,N_367);
and U1176 (N_1176,N_599,N_162);
and U1177 (N_1177,N_14,N_360);
xnor U1178 (N_1178,N_378,N_186);
and U1179 (N_1179,N_96,N_300);
and U1180 (N_1180,N_167,N_268);
or U1181 (N_1181,N_470,N_51);
or U1182 (N_1182,N_174,N_590);
nand U1183 (N_1183,N_173,N_89);
and U1184 (N_1184,N_111,N_506);
and U1185 (N_1185,N_479,N_229);
nor U1186 (N_1186,N_345,N_455);
and U1187 (N_1187,N_134,N_229);
or U1188 (N_1188,N_517,N_592);
nor U1189 (N_1189,N_474,N_438);
and U1190 (N_1190,N_327,N_532);
xnor U1191 (N_1191,N_502,N_520);
nand U1192 (N_1192,N_370,N_237);
nand U1193 (N_1193,N_225,N_359);
nor U1194 (N_1194,N_339,N_67);
or U1195 (N_1195,N_79,N_154);
nand U1196 (N_1196,N_530,N_555);
nand U1197 (N_1197,N_347,N_200);
nand U1198 (N_1198,N_4,N_97);
or U1199 (N_1199,N_408,N_585);
or U1200 (N_1200,N_1126,N_772);
nor U1201 (N_1201,N_863,N_804);
nor U1202 (N_1202,N_937,N_663);
or U1203 (N_1203,N_720,N_854);
and U1204 (N_1204,N_1112,N_820);
or U1205 (N_1205,N_717,N_1137);
xnor U1206 (N_1206,N_982,N_615);
or U1207 (N_1207,N_851,N_935);
nand U1208 (N_1208,N_1035,N_697);
or U1209 (N_1209,N_818,N_660);
and U1210 (N_1210,N_852,N_610);
or U1211 (N_1211,N_1109,N_791);
nor U1212 (N_1212,N_920,N_1075);
xor U1213 (N_1213,N_977,N_844);
or U1214 (N_1214,N_867,N_886);
and U1215 (N_1215,N_1133,N_666);
nor U1216 (N_1216,N_683,N_605);
or U1217 (N_1217,N_693,N_871);
and U1218 (N_1218,N_691,N_777);
nor U1219 (N_1219,N_698,N_1032);
and U1220 (N_1220,N_1163,N_827);
and U1221 (N_1221,N_946,N_1167);
or U1222 (N_1222,N_951,N_1192);
nor U1223 (N_1223,N_1123,N_744);
and U1224 (N_1224,N_923,N_799);
nand U1225 (N_1225,N_892,N_1073);
and U1226 (N_1226,N_896,N_828);
nor U1227 (N_1227,N_721,N_779);
nor U1228 (N_1228,N_736,N_908);
xor U1229 (N_1229,N_652,N_996);
nand U1230 (N_1230,N_753,N_1113);
nand U1231 (N_1231,N_927,N_943);
nand U1232 (N_1232,N_624,N_1168);
and U1233 (N_1233,N_1128,N_948);
nor U1234 (N_1234,N_1066,N_899);
and U1235 (N_1235,N_1037,N_1030);
and U1236 (N_1236,N_859,N_695);
nand U1237 (N_1237,N_1079,N_760);
nor U1238 (N_1238,N_606,N_797);
nand U1239 (N_1239,N_857,N_1040);
nand U1240 (N_1240,N_648,N_767);
or U1241 (N_1241,N_914,N_748);
xnor U1242 (N_1242,N_677,N_879);
or U1243 (N_1243,N_646,N_1161);
and U1244 (N_1244,N_862,N_809);
or U1245 (N_1245,N_990,N_637);
or U1246 (N_1246,N_706,N_626);
nor U1247 (N_1247,N_659,N_685);
and U1248 (N_1248,N_641,N_738);
nor U1249 (N_1249,N_814,N_623);
nand U1250 (N_1250,N_993,N_1012);
nand U1251 (N_1251,N_1063,N_1159);
xor U1252 (N_1252,N_1064,N_917);
or U1253 (N_1253,N_826,N_702);
and U1254 (N_1254,N_703,N_1180);
and U1255 (N_1255,N_1174,N_654);
or U1256 (N_1256,N_1067,N_1083);
and U1257 (N_1257,N_895,N_688);
nor U1258 (N_1258,N_672,N_1122);
xnor U1259 (N_1259,N_653,N_1042);
nor U1260 (N_1260,N_788,N_1096);
and U1261 (N_1261,N_671,N_620);
and U1262 (N_1262,N_785,N_942);
and U1263 (N_1263,N_1087,N_1149);
nand U1264 (N_1264,N_1018,N_836);
nand U1265 (N_1265,N_1028,N_1026);
nand U1266 (N_1266,N_764,N_1175);
or U1267 (N_1267,N_750,N_725);
or U1268 (N_1268,N_1015,N_1115);
nor U1269 (N_1269,N_658,N_740);
or U1270 (N_1270,N_1154,N_861);
nor U1271 (N_1271,N_1121,N_766);
nor U1272 (N_1272,N_1050,N_643);
xor U1273 (N_1273,N_971,N_656);
nor U1274 (N_1274,N_619,N_1024);
or U1275 (N_1275,N_898,N_819);
or U1276 (N_1276,N_1044,N_783);
nand U1277 (N_1277,N_746,N_841);
nor U1278 (N_1278,N_770,N_701);
nor U1279 (N_1279,N_934,N_612);
and U1280 (N_1280,N_1020,N_1006);
or U1281 (N_1281,N_604,N_711);
and U1282 (N_1282,N_911,N_773);
nor U1283 (N_1283,N_732,N_903);
and U1284 (N_1284,N_1136,N_860);
or U1285 (N_1285,N_918,N_930);
nor U1286 (N_1286,N_1094,N_1147);
and U1287 (N_1287,N_897,N_782);
nor U1288 (N_1288,N_800,N_616);
or U1289 (N_1289,N_1150,N_751);
nand U1290 (N_1290,N_823,N_668);
or U1291 (N_1291,N_1118,N_902);
or U1292 (N_1292,N_768,N_1106);
nor U1293 (N_1293,N_793,N_759);
xnor U1294 (N_1294,N_963,N_1068);
or U1295 (N_1295,N_661,N_1101);
xor U1296 (N_1296,N_792,N_1116);
and U1297 (N_1297,N_962,N_737);
nand U1298 (N_1298,N_1127,N_1141);
or U1299 (N_1299,N_667,N_815);
nor U1300 (N_1300,N_821,N_1186);
or U1301 (N_1301,N_1119,N_1196);
nand U1302 (N_1302,N_719,N_628);
nand U1303 (N_1303,N_651,N_912);
nand U1304 (N_1304,N_1190,N_954);
and U1305 (N_1305,N_1059,N_1130);
nor U1306 (N_1306,N_1048,N_1148);
and U1307 (N_1307,N_1074,N_713);
nor U1308 (N_1308,N_1086,N_869);
or U1309 (N_1309,N_795,N_1146);
or U1310 (N_1310,N_709,N_974);
or U1311 (N_1311,N_1003,N_617);
nand U1312 (N_1312,N_634,N_822);
nand U1313 (N_1313,N_925,N_994);
xnor U1314 (N_1314,N_728,N_1071);
and U1315 (N_1315,N_1093,N_1081);
nand U1316 (N_1316,N_1008,N_1041);
nor U1317 (N_1317,N_627,N_989);
nor U1318 (N_1318,N_931,N_1107);
and U1319 (N_1319,N_975,N_1102);
or U1320 (N_1320,N_1198,N_831);
nor U1321 (N_1321,N_998,N_763);
nor U1322 (N_1322,N_944,N_665);
and U1323 (N_1323,N_774,N_850);
nand U1324 (N_1324,N_647,N_621);
nand U1325 (N_1325,N_1043,N_858);
and U1326 (N_1326,N_1017,N_1090);
xor U1327 (N_1327,N_835,N_622);
nor U1328 (N_1328,N_889,N_716);
nor U1329 (N_1329,N_765,N_747);
nand U1330 (N_1330,N_1194,N_1053);
nor U1331 (N_1331,N_1124,N_781);
nor U1332 (N_1332,N_743,N_1185);
xor U1333 (N_1333,N_900,N_825);
or U1334 (N_1334,N_714,N_1010);
xor U1335 (N_1335,N_762,N_1111);
xnor U1336 (N_1336,N_676,N_838);
nand U1337 (N_1337,N_864,N_1135);
and U1338 (N_1338,N_1193,N_981);
or U1339 (N_1339,N_630,N_790);
nor U1340 (N_1340,N_674,N_1076);
or U1341 (N_1341,N_890,N_884);
and U1342 (N_1342,N_689,N_1001);
and U1343 (N_1343,N_915,N_1052);
nor U1344 (N_1344,N_1078,N_955);
or U1345 (N_1345,N_1069,N_893);
nand U1346 (N_1346,N_1016,N_947);
or U1347 (N_1347,N_887,N_832);
nand U1348 (N_1348,N_1179,N_1100);
or U1349 (N_1349,N_849,N_960);
nor U1350 (N_1350,N_855,N_1011);
xnor U1351 (N_1351,N_970,N_754);
and U1352 (N_1352,N_965,N_905);
nor U1353 (N_1353,N_649,N_1143);
nor U1354 (N_1354,N_1110,N_929);
nand U1355 (N_1355,N_1004,N_924);
or U1356 (N_1356,N_904,N_662);
nand U1357 (N_1357,N_913,N_723);
and U1358 (N_1358,N_1097,N_839);
nand U1359 (N_1359,N_878,N_1164);
and U1360 (N_1360,N_794,N_1065);
xnor U1361 (N_1361,N_873,N_1084);
nor U1362 (N_1362,N_1120,N_988);
nand U1363 (N_1363,N_876,N_976);
nand U1364 (N_1364,N_638,N_603);
or U1365 (N_1365,N_699,N_776);
and U1366 (N_1366,N_845,N_956);
or U1367 (N_1367,N_817,N_984);
nand U1368 (N_1368,N_1000,N_1153);
or U1369 (N_1369,N_999,N_805);
or U1370 (N_1370,N_938,N_964);
or U1371 (N_1371,N_611,N_629);
and U1372 (N_1372,N_803,N_967);
and U1373 (N_1373,N_694,N_690);
and U1374 (N_1374,N_885,N_1199);
nand U1375 (N_1375,N_847,N_881);
and U1376 (N_1376,N_731,N_1021);
nand U1377 (N_1377,N_966,N_1082);
nand U1378 (N_1378,N_812,N_882);
nor U1379 (N_1379,N_718,N_1061);
and U1380 (N_1380,N_866,N_761);
nand U1381 (N_1381,N_707,N_1165);
xnor U1382 (N_1382,N_940,N_921);
nor U1383 (N_1383,N_837,N_1013);
nand U1384 (N_1384,N_1144,N_843);
nand U1385 (N_1385,N_932,N_1023);
and U1386 (N_1386,N_1056,N_1181);
nand U1387 (N_1387,N_957,N_600);
nor U1388 (N_1388,N_686,N_1172);
or U1389 (N_1389,N_1027,N_687);
and U1390 (N_1390,N_644,N_657);
nor U1391 (N_1391,N_983,N_735);
or U1392 (N_1392,N_1139,N_1080);
xnor U1393 (N_1393,N_985,N_875);
nor U1394 (N_1394,N_1105,N_874);
and U1395 (N_1395,N_991,N_1054);
or U1396 (N_1396,N_916,N_1045);
or U1397 (N_1397,N_1095,N_883);
nor U1398 (N_1398,N_891,N_696);
and U1399 (N_1399,N_769,N_952);
nor U1400 (N_1400,N_953,N_992);
and U1401 (N_1401,N_1062,N_986);
nor U1402 (N_1402,N_910,N_1189);
xor U1403 (N_1403,N_1085,N_1142);
or U1404 (N_1404,N_880,N_901);
and U1405 (N_1405,N_1091,N_758);
nor U1406 (N_1406,N_1134,N_1009);
and U1407 (N_1407,N_1005,N_933);
and U1408 (N_1408,N_692,N_987);
nor U1409 (N_1409,N_1014,N_1019);
xor U1410 (N_1410,N_727,N_700);
or U1411 (N_1411,N_870,N_734);
and U1412 (N_1412,N_664,N_1131);
and U1413 (N_1413,N_877,N_848);
and U1414 (N_1414,N_907,N_1046);
xor U1415 (N_1415,N_950,N_1058);
nor U1416 (N_1416,N_1140,N_796);
and U1417 (N_1417,N_1157,N_1051);
nand U1418 (N_1418,N_1169,N_730);
nand U1419 (N_1419,N_1184,N_1156);
nand U1420 (N_1420,N_655,N_979);
nand U1421 (N_1421,N_1089,N_926);
or U1422 (N_1422,N_949,N_1070);
nor U1423 (N_1423,N_784,N_749);
or U1424 (N_1424,N_670,N_633);
or U1425 (N_1425,N_789,N_941);
and U1426 (N_1426,N_607,N_1171);
or U1427 (N_1427,N_787,N_1151);
nand U1428 (N_1428,N_798,N_724);
nand U1429 (N_1429,N_733,N_675);
or U1430 (N_1430,N_705,N_636);
or U1431 (N_1431,N_816,N_919);
nor U1432 (N_1432,N_1166,N_1155);
nor U1433 (N_1433,N_936,N_1177);
nor U1434 (N_1434,N_1117,N_1114);
and U1435 (N_1435,N_802,N_958);
nor U1436 (N_1436,N_906,N_807);
nor U1437 (N_1437,N_1092,N_980);
and U1438 (N_1438,N_856,N_1036);
and U1439 (N_1439,N_669,N_968);
xor U1440 (N_1440,N_1047,N_609);
nor U1441 (N_1441,N_1057,N_846);
nand U1442 (N_1442,N_1188,N_618);
or U1443 (N_1443,N_1049,N_715);
and U1444 (N_1444,N_1195,N_973);
and U1445 (N_1445,N_834,N_625);
nor U1446 (N_1446,N_729,N_757);
and U1447 (N_1447,N_972,N_1077);
and U1448 (N_1448,N_1055,N_1138);
nand U1449 (N_1449,N_673,N_639);
and U1450 (N_1450,N_997,N_1132);
or U1451 (N_1451,N_833,N_1125);
and U1452 (N_1452,N_808,N_1039);
nand U1453 (N_1453,N_631,N_1158);
and U1454 (N_1454,N_682,N_739);
nand U1455 (N_1455,N_745,N_704);
xor U1456 (N_1456,N_868,N_842);
nand U1457 (N_1457,N_1183,N_1170);
or U1458 (N_1458,N_756,N_632);
nand U1459 (N_1459,N_922,N_726);
and U1460 (N_1460,N_1007,N_1088);
nand U1461 (N_1461,N_1034,N_995);
and U1462 (N_1462,N_928,N_959);
nand U1463 (N_1463,N_1160,N_601);
nor U1464 (N_1464,N_1104,N_778);
nand U1465 (N_1465,N_909,N_613);
nand U1466 (N_1466,N_1103,N_1129);
xor U1467 (N_1467,N_1191,N_635);
or U1468 (N_1468,N_872,N_1176);
and U1469 (N_1469,N_645,N_780);
nor U1470 (N_1470,N_810,N_1025);
nand U1471 (N_1471,N_742,N_710);
and U1472 (N_1472,N_1033,N_978);
or U1473 (N_1473,N_1162,N_708);
or U1474 (N_1474,N_811,N_680);
nand U1475 (N_1475,N_853,N_1029);
nor U1476 (N_1476,N_829,N_684);
and U1477 (N_1477,N_786,N_840);
or U1478 (N_1478,N_1178,N_1152);
nor U1479 (N_1479,N_755,N_741);
xnor U1480 (N_1480,N_722,N_830);
and U1481 (N_1481,N_1098,N_771);
or U1482 (N_1482,N_801,N_1038);
nand U1483 (N_1483,N_961,N_1197);
nor U1484 (N_1484,N_1108,N_642);
nor U1485 (N_1485,N_1022,N_640);
nand U1486 (N_1486,N_678,N_1031);
and U1487 (N_1487,N_775,N_614);
nand U1488 (N_1488,N_1145,N_752);
nor U1489 (N_1489,N_712,N_939);
and U1490 (N_1490,N_824,N_650);
or U1491 (N_1491,N_1002,N_602);
nand U1492 (N_1492,N_1173,N_608);
nand U1493 (N_1493,N_888,N_969);
or U1494 (N_1494,N_679,N_1072);
xnor U1495 (N_1495,N_865,N_945);
and U1496 (N_1496,N_806,N_1060);
nor U1497 (N_1497,N_681,N_1099);
or U1498 (N_1498,N_813,N_1182);
nor U1499 (N_1499,N_894,N_1187);
nor U1500 (N_1500,N_1104,N_1012);
nand U1501 (N_1501,N_1179,N_1158);
nor U1502 (N_1502,N_976,N_840);
nand U1503 (N_1503,N_890,N_709);
or U1504 (N_1504,N_1173,N_1171);
or U1505 (N_1505,N_1125,N_941);
nor U1506 (N_1506,N_824,N_886);
and U1507 (N_1507,N_1084,N_1101);
and U1508 (N_1508,N_601,N_825);
nor U1509 (N_1509,N_898,N_989);
xor U1510 (N_1510,N_957,N_657);
and U1511 (N_1511,N_1170,N_860);
or U1512 (N_1512,N_630,N_1091);
xnor U1513 (N_1513,N_924,N_902);
xnor U1514 (N_1514,N_1038,N_807);
xnor U1515 (N_1515,N_713,N_1028);
nor U1516 (N_1516,N_731,N_916);
or U1517 (N_1517,N_1142,N_635);
and U1518 (N_1518,N_1195,N_1115);
or U1519 (N_1519,N_1094,N_966);
xor U1520 (N_1520,N_710,N_919);
nand U1521 (N_1521,N_1080,N_1173);
nor U1522 (N_1522,N_933,N_639);
nand U1523 (N_1523,N_1016,N_1079);
nand U1524 (N_1524,N_773,N_873);
and U1525 (N_1525,N_1137,N_732);
nand U1526 (N_1526,N_1056,N_1198);
nor U1527 (N_1527,N_631,N_925);
or U1528 (N_1528,N_721,N_895);
or U1529 (N_1529,N_977,N_711);
or U1530 (N_1530,N_813,N_1079);
nand U1531 (N_1531,N_739,N_862);
and U1532 (N_1532,N_652,N_822);
nor U1533 (N_1533,N_1004,N_1094);
or U1534 (N_1534,N_1157,N_1039);
and U1535 (N_1535,N_728,N_834);
xor U1536 (N_1536,N_788,N_643);
xnor U1537 (N_1537,N_1178,N_745);
and U1538 (N_1538,N_1094,N_896);
or U1539 (N_1539,N_1132,N_972);
or U1540 (N_1540,N_717,N_719);
nor U1541 (N_1541,N_762,N_616);
or U1542 (N_1542,N_1079,N_825);
or U1543 (N_1543,N_811,N_967);
nand U1544 (N_1544,N_1094,N_1182);
nand U1545 (N_1545,N_1009,N_993);
xnor U1546 (N_1546,N_686,N_1103);
or U1547 (N_1547,N_660,N_746);
xnor U1548 (N_1548,N_748,N_743);
nor U1549 (N_1549,N_786,N_697);
or U1550 (N_1550,N_1001,N_865);
or U1551 (N_1551,N_1157,N_676);
or U1552 (N_1552,N_809,N_963);
nor U1553 (N_1553,N_859,N_1166);
nand U1554 (N_1554,N_1198,N_819);
or U1555 (N_1555,N_894,N_1159);
xnor U1556 (N_1556,N_1104,N_613);
or U1557 (N_1557,N_1178,N_819);
and U1558 (N_1558,N_971,N_689);
nor U1559 (N_1559,N_1105,N_1196);
nand U1560 (N_1560,N_830,N_1193);
and U1561 (N_1561,N_948,N_1018);
or U1562 (N_1562,N_809,N_649);
or U1563 (N_1563,N_1067,N_1011);
nor U1564 (N_1564,N_817,N_739);
or U1565 (N_1565,N_990,N_969);
and U1566 (N_1566,N_911,N_1017);
and U1567 (N_1567,N_983,N_681);
xor U1568 (N_1568,N_1121,N_1039);
xor U1569 (N_1569,N_601,N_658);
and U1570 (N_1570,N_1051,N_1166);
and U1571 (N_1571,N_1053,N_1093);
nor U1572 (N_1572,N_926,N_1151);
and U1573 (N_1573,N_887,N_913);
nor U1574 (N_1574,N_1141,N_1002);
or U1575 (N_1575,N_1157,N_771);
xor U1576 (N_1576,N_799,N_1020);
and U1577 (N_1577,N_670,N_919);
nor U1578 (N_1578,N_979,N_908);
nand U1579 (N_1579,N_1032,N_949);
nand U1580 (N_1580,N_1092,N_1108);
or U1581 (N_1581,N_1027,N_1077);
nor U1582 (N_1582,N_1109,N_1188);
nor U1583 (N_1583,N_688,N_840);
nor U1584 (N_1584,N_1124,N_1044);
nand U1585 (N_1585,N_1155,N_1177);
or U1586 (N_1586,N_1156,N_767);
or U1587 (N_1587,N_650,N_984);
or U1588 (N_1588,N_697,N_727);
nand U1589 (N_1589,N_1076,N_764);
or U1590 (N_1590,N_1107,N_730);
and U1591 (N_1591,N_1144,N_1088);
nand U1592 (N_1592,N_731,N_923);
nand U1593 (N_1593,N_924,N_829);
and U1594 (N_1594,N_1085,N_911);
and U1595 (N_1595,N_1096,N_714);
or U1596 (N_1596,N_776,N_1046);
nand U1597 (N_1597,N_1130,N_800);
nand U1598 (N_1598,N_834,N_1059);
and U1599 (N_1599,N_901,N_661);
nand U1600 (N_1600,N_982,N_1089);
or U1601 (N_1601,N_880,N_649);
and U1602 (N_1602,N_975,N_662);
nand U1603 (N_1603,N_925,N_1150);
nand U1604 (N_1604,N_946,N_900);
nor U1605 (N_1605,N_795,N_790);
or U1606 (N_1606,N_770,N_847);
or U1607 (N_1607,N_931,N_610);
and U1608 (N_1608,N_1134,N_1158);
nand U1609 (N_1609,N_611,N_785);
nor U1610 (N_1610,N_1046,N_742);
or U1611 (N_1611,N_1128,N_974);
and U1612 (N_1612,N_803,N_681);
nor U1613 (N_1613,N_1014,N_864);
nand U1614 (N_1614,N_768,N_854);
or U1615 (N_1615,N_861,N_823);
xnor U1616 (N_1616,N_1162,N_949);
xnor U1617 (N_1617,N_710,N_688);
xnor U1618 (N_1618,N_699,N_1035);
nor U1619 (N_1619,N_1198,N_931);
nand U1620 (N_1620,N_746,N_607);
nand U1621 (N_1621,N_855,N_936);
nor U1622 (N_1622,N_1122,N_688);
xnor U1623 (N_1623,N_766,N_874);
nand U1624 (N_1624,N_746,N_722);
nand U1625 (N_1625,N_781,N_618);
nand U1626 (N_1626,N_1109,N_674);
nand U1627 (N_1627,N_874,N_1168);
nand U1628 (N_1628,N_642,N_1059);
nor U1629 (N_1629,N_869,N_636);
and U1630 (N_1630,N_759,N_1186);
and U1631 (N_1631,N_983,N_790);
nor U1632 (N_1632,N_853,N_927);
nor U1633 (N_1633,N_963,N_1145);
nand U1634 (N_1634,N_1106,N_1009);
and U1635 (N_1635,N_1013,N_816);
xnor U1636 (N_1636,N_990,N_674);
or U1637 (N_1637,N_1081,N_622);
or U1638 (N_1638,N_1151,N_920);
nor U1639 (N_1639,N_916,N_818);
nand U1640 (N_1640,N_646,N_1087);
nand U1641 (N_1641,N_721,N_1165);
nand U1642 (N_1642,N_1055,N_1123);
or U1643 (N_1643,N_828,N_946);
nand U1644 (N_1644,N_790,N_943);
nand U1645 (N_1645,N_871,N_969);
nor U1646 (N_1646,N_745,N_1042);
nor U1647 (N_1647,N_1195,N_633);
nor U1648 (N_1648,N_744,N_1085);
nand U1649 (N_1649,N_1126,N_835);
nand U1650 (N_1650,N_980,N_729);
nand U1651 (N_1651,N_769,N_1018);
nor U1652 (N_1652,N_1192,N_747);
or U1653 (N_1653,N_799,N_709);
nand U1654 (N_1654,N_682,N_928);
nor U1655 (N_1655,N_955,N_813);
or U1656 (N_1656,N_1054,N_903);
or U1657 (N_1657,N_808,N_613);
and U1658 (N_1658,N_1096,N_1057);
nor U1659 (N_1659,N_754,N_798);
nor U1660 (N_1660,N_721,N_828);
nor U1661 (N_1661,N_659,N_941);
and U1662 (N_1662,N_846,N_1178);
nand U1663 (N_1663,N_687,N_903);
or U1664 (N_1664,N_679,N_646);
and U1665 (N_1665,N_646,N_806);
xnor U1666 (N_1666,N_849,N_1016);
and U1667 (N_1667,N_671,N_666);
nor U1668 (N_1668,N_664,N_910);
nand U1669 (N_1669,N_723,N_772);
nor U1670 (N_1670,N_978,N_815);
or U1671 (N_1671,N_858,N_928);
or U1672 (N_1672,N_934,N_859);
or U1673 (N_1673,N_994,N_1084);
xnor U1674 (N_1674,N_808,N_620);
and U1675 (N_1675,N_1118,N_808);
nor U1676 (N_1676,N_1149,N_732);
and U1677 (N_1677,N_953,N_1101);
nor U1678 (N_1678,N_1123,N_868);
nand U1679 (N_1679,N_969,N_1176);
nor U1680 (N_1680,N_729,N_788);
or U1681 (N_1681,N_1039,N_1154);
nor U1682 (N_1682,N_770,N_707);
nand U1683 (N_1683,N_912,N_693);
nand U1684 (N_1684,N_1129,N_1154);
or U1685 (N_1685,N_846,N_921);
and U1686 (N_1686,N_951,N_1029);
and U1687 (N_1687,N_777,N_987);
or U1688 (N_1688,N_808,N_1090);
nor U1689 (N_1689,N_740,N_726);
xor U1690 (N_1690,N_1126,N_640);
and U1691 (N_1691,N_875,N_1135);
nand U1692 (N_1692,N_750,N_1041);
and U1693 (N_1693,N_668,N_1139);
nand U1694 (N_1694,N_970,N_888);
xnor U1695 (N_1695,N_920,N_1039);
or U1696 (N_1696,N_682,N_1089);
nor U1697 (N_1697,N_1024,N_837);
nor U1698 (N_1698,N_827,N_835);
or U1699 (N_1699,N_1023,N_930);
nand U1700 (N_1700,N_844,N_1100);
or U1701 (N_1701,N_1043,N_755);
nor U1702 (N_1702,N_699,N_989);
or U1703 (N_1703,N_1167,N_670);
nor U1704 (N_1704,N_1044,N_903);
and U1705 (N_1705,N_716,N_804);
and U1706 (N_1706,N_655,N_754);
and U1707 (N_1707,N_1171,N_960);
nand U1708 (N_1708,N_920,N_721);
nand U1709 (N_1709,N_737,N_915);
nor U1710 (N_1710,N_683,N_1158);
or U1711 (N_1711,N_965,N_995);
and U1712 (N_1712,N_790,N_846);
and U1713 (N_1713,N_885,N_620);
nor U1714 (N_1714,N_984,N_1111);
or U1715 (N_1715,N_634,N_601);
xor U1716 (N_1716,N_1146,N_627);
nand U1717 (N_1717,N_1022,N_1161);
or U1718 (N_1718,N_1078,N_965);
or U1719 (N_1719,N_1080,N_1157);
or U1720 (N_1720,N_849,N_1028);
or U1721 (N_1721,N_677,N_978);
xor U1722 (N_1722,N_638,N_680);
nand U1723 (N_1723,N_676,N_884);
or U1724 (N_1724,N_686,N_1087);
or U1725 (N_1725,N_711,N_1018);
nand U1726 (N_1726,N_744,N_704);
xor U1727 (N_1727,N_1063,N_1190);
and U1728 (N_1728,N_868,N_742);
nor U1729 (N_1729,N_958,N_881);
nand U1730 (N_1730,N_939,N_725);
or U1731 (N_1731,N_1180,N_732);
nor U1732 (N_1732,N_951,N_731);
nand U1733 (N_1733,N_1097,N_819);
xor U1734 (N_1734,N_638,N_1140);
or U1735 (N_1735,N_835,N_908);
or U1736 (N_1736,N_922,N_807);
and U1737 (N_1737,N_623,N_984);
nand U1738 (N_1738,N_891,N_624);
xnor U1739 (N_1739,N_1197,N_879);
nor U1740 (N_1740,N_944,N_1162);
xnor U1741 (N_1741,N_611,N_1054);
and U1742 (N_1742,N_1067,N_839);
and U1743 (N_1743,N_1089,N_798);
nand U1744 (N_1744,N_1047,N_936);
nand U1745 (N_1745,N_858,N_790);
nor U1746 (N_1746,N_737,N_937);
and U1747 (N_1747,N_1004,N_747);
xor U1748 (N_1748,N_1045,N_850);
or U1749 (N_1749,N_810,N_1093);
nand U1750 (N_1750,N_1159,N_931);
or U1751 (N_1751,N_965,N_1042);
nand U1752 (N_1752,N_603,N_756);
or U1753 (N_1753,N_939,N_1058);
or U1754 (N_1754,N_610,N_983);
or U1755 (N_1755,N_1122,N_680);
nor U1756 (N_1756,N_1070,N_618);
nor U1757 (N_1757,N_963,N_608);
nand U1758 (N_1758,N_1022,N_661);
or U1759 (N_1759,N_793,N_844);
nor U1760 (N_1760,N_736,N_857);
and U1761 (N_1761,N_687,N_1130);
nor U1762 (N_1762,N_1032,N_643);
and U1763 (N_1763,N_1023,N_1185);
or U1764 (N_1764,N_855,N_743);
or U1765 (N_1765,N_911,N_1069);
or U1766 (N_1766,N_1111,N_1137);
or U1767 (N_1767,N_1073,N_855);
and U1768 (N_1768,N_823,N_849);
nand U1769 (N_1769,N_892,N_1164);
or U1770 (N_1770,N_934,N_1191);
or U1771 (N_1771,N_1028,N_1085);
and U1772 (N_1772,N_1032,N_695);
and U1773 (N_1773,N_1042,N_679);
nor U1774 (N_1774,N_852,N_742);
xor U1775 (N_1775,N_731,N_817);
xor U1776 (N_1776,N_1176,N_635);
xor U1777 (N_1777,N_799,N_851);
nor U1778 (N_1778,N_726,N_975);
or U1779 (N_1779,N_1169,N_1008);
or U1780 (N_1780,N_819,N_1167);
or U1781 (N_1781,N_988,N_970);
xor U1782 (N_1782,N_1078,N_1053);
or U1783 (N_1783,N_908,N_728);
and U1784 (N_1784,N_814,N_1133);
nand U1785 (N_1785,N_608,N_731);
nand U1786 (N_1786,N_1154,N_712);
nor U1787 (N_1787,N_1047,N_921);
and U1788 (N_1788,N_693,N_634);
nor U1789 (N_1789,N_799,N_869);
or U1790 (N_1790,N_648,N_1132);
and U1791 (N_1791,N_610,N_1048);
or U1792 (N_1792,N_1142,N_1000);
nor U1793 (N_1793,N_650,N_947);
or U1794 (N_1794,N_1060,N_1138);
or U1795 (N_1795,N_777,N_674);
nand U1796 (N_1796,N_834,N_799);
nand U1797 (N_1797,N_1020,N_1046);
xor U1798 (N_1798,N_1039,N_681);
xor U1799 (N_1799,N_829,N_1199);
nor U1800 (N_1800,N_1633,N_1660);
and U1801 (N_1801,N_1708,N_1426);
and U1802 (N_1802,N_1254,N_1569);
xor U1803 (N_1803,N_1796,N_1518);
nand U1804 (N_1804,N_1514,N_1226);
or U1805 (N_1805,N_1447,N_1430);
or U1806 (N_1806,N_1616,N_1346);
and U1807 (N_1807,N_1448,N_1693);
nor U1808 (N_1808,N_1302,N_1663);
nand U1809 (N_1809,N_1428,N_1639);
nor U1810 (N_1810,N_1533,N_1535);
nor U1811 (N_1811,N_1750,N_1478);
and U1812 (N_1812,N_1532,N_1435);
and U1813 (N_1813,N_1352,N_1632);
and U1814 (N_1814,N_1722,N_1363);
and U1815 (N_1815,N_1218,N_1730);
and U1816 (N_1816,N_1592,N_1402);
xor U1817 (N_1817,N_1502,N_1701);
nand U1818 (N_1818,N_1513,N_1604);
xor U1819 (N_1819,N_1599,N_1798);
nand U1820 (N_1820,N_1232,N_1643);
nor U1821 (N_1821,N_1698,N_1765);
nor U1822 (N_1822,N_1760,N_1259);
or U1823 (N_1823,N_1622,N_1570);
or U1824 (N_1824,N_1574,N_1635);
nor U1825 (N_1825,N_1749,N_1705);
and U1826 (N_1826,N_1328,N_1648);
or U1827 (N_1827,N_1207,N_1624);
nand U1828 (N_1828,N_1679,N_1364);
nand U1829 (N_1829,N_1534,N_1271);
and U1830 (N_1830,N_1640,N_1618);
nand U1831 (N_1831,N_1290,N_1689);
xnor U1832 (N_1832,N_1313,N_1307);
nand U1833 (N_1833,N_1641,N_1475);
nor U1834 (N_1834,N_1751,N_1219);
and U1835 (N_1835,N_1748,N_1530);
and U1836 (N_1836,N_1595,N_1319);
and U1837 (N_1837,N_1339,N_1243);
nor U1838 (N_1838,N_1617,N_1706);
nand U1839 (N_1839,N_1281,N_1262);
and U1840 (N_1840,N_1436,N_1357);
or U1841 (N_1841,N_1270,N_1754);
nor U1842 (N_1842,N_1403,N_1332);
and U1843 (N_1843,N_1538,N_1345);
or U1844 (N_1844,N_1690,N_1309);
or U1845 (N_1845,N_1770,N_1761);
nand U1846 (N_1846,N_1227,N_1501);
and U1847 (N_1847,N_1318,N_1744);
nor U1848 (N_1848,N_1623,N_1598);
and U1849 (N_1849,N_1552,N_1284);
and U1850 (N_1850,N_1631,N_1713);
nor U1851 (N_1851,N_1253,N_1293);
nor U1852 (N_1852,N_1546,N_1509);
nor U1853 (N_1853,N_1659,N_1731);
and U1854 (N_1854,N_1782,N_1335);
and U1855 (N_1855,N_1238,N_1753);
nand U1856 (N_1856,N_1649,N_1220);
nor U1857 (N_1857,N_1579,N_1456);
and U1858 (N_1858,N_1490,N_1740);
and U1859 (N_1859,N_1555,N_1461);
or U1860 (N_1860,N_1576,N_1429);
xnor U1861 (N_1861,N_1497,N_1607);
and U1862 (N_1862,N_1463,N_1367);
nor U1863 (N_1863,N_1375,N_1386);
nand U1864 (N_1864,N_1645,N_1223);
nand U1865 (N_1865,N_1266,N_1383);
or U1866 (N_1866,N_1333,N_1491);
or U1867 (N_1867,N_1687,N_1504);
nor U1868 (N_1868,N_1344,N_1390);
nor U1869 (N_1869,N_1489,N_1756);
and U1870 (N_1870,N_1483,N_1746);
and U1871 (N_1871,N_1588,N_1331);
xnor U1872 (N_1872,N_1597,N_1771);
xor U1873 (N_1873,N_1289,N_1723);
and U1874 (N_1874,N_1303,N_1239);
nor U1875 (N_1875,N_1324,N_1288);
xnor U1876 (N_1876,N_1314,N_1421);
and U1877 (N_1877,N_1404,N_1629);
and U1878 (N_1878,N_1707,N_1712);
and U1879 (N_1879,N_1205,N_1443);
and U1880 (N_1880,N_1728,N_1469);
xnor U1881 (N_1881,N_1385,N_1638);
nor U1882 (N_1882,N_1374,N_1789);
and U1883 (N_1883,N_1371,N_1544);
nand U1884 (N_1884,N_1221,N_1755);
and U1885 (N_1885,N_1554,N_1373);
or U1886 (N_1886,N_1672,N_1353);
or U1887 (N_1887,N_1234,N_1279);
or U1888 (N_1888,N_1721,N_1260);
nand U1889 (N_1889,N_1591,N_1583);
or U1890 (N_1890,N_1275,N_1615);
nand U1891 (N_1891,N_1557,N_1778);
xnor U1892 (N_1892,N_1717,N_1425);
nor U1893 (N_1893,N_1337,N_1452);
or U1894 (N_1894,N_1681,N_1377);
or U1895 (N_1895,N_1274,N_1587);
nand U1896 (N_1896,N_1695,N_1568);
xnor U1897 (N_1897,N_1590,N_1556);
or U1898 (N_1898,N_1537,N_1764);
or U1899 (N_1899,N_1424,N_1272);
or U1900 (N_1900,N_1244,N_1773);
or U1901 (N_1901,N_1406,N_1358);
nor U1902 (N_1902,N_1342,N_1258);
nand U1903 (N_1903,N_1686,N_1738);
nor U1904 (N_1904,N_1348,N_1512);
and U1905 (N_1905,N_1376,N_1567);
or U1906 (N_1906,N_1321,N_1628);
or U1907 (N_1907,N_1246,N_1529);
nand U1908 (N_1908,N_1451,N_1264);
and U1909 (N_1909,N_1439,N_1602);
nor U1910 (N_1910,N_1212,N_1308);
nor U1911 (N_1911,N_1545,N_1393);
nor U1912 (N_1912,N_1236,N_1735);
nor U1913 (N_1913,N_1336,N_1691);
nand U1914 (N_1914,N_1206,N_1547);
or U1915 (N_1915,N_1630,N_1474);
nor U1916 (N_1916,N_1745,N_1669);
xor U1917 (N_1917,N_1280,N_1453);
nand U1918 (N_1918,N_1522,N_1454);
nand U1919 (N_1919,N_1397,N_1481);
or U1920 (N_1920,N_1601,N_1411);
xor U1921 (N_1921,N_1634,N_1528);
nor U1922 (N_1922,N_1656,N_1479);
or U1923 (N_1923,N_1763,N_1379);
and U1924 (N_1924,N_1255,N_1295);
or U1925 (N_1925,N_1322,N_1694);
or U1926 (N_1926,N_1580,N_1543);
or U1927 (N_1927,N_1500,N_1593);
and U1928 (N_1928,N_1487,N_1305);
nand U1929 (N_1929,N_1651,N_1596);
nand U1930 (N_1930,N_1298,N_1384);
or U1931 (N_1931,N_1667,N_1269);
nand U1932 (N_1932,N_1285,N_1503);
nand U1933 (N_1933,N_1432,N_1304);
or U1934 (N_1934,N_1654,N_1495);
or U1935 (N_1935,N_1440,N_1642);
nand U1936 (N_1936,N_1678,N_1445);
and U1937 (N_1937,N_1215,N_1431);
or U1938 (N_1938,N_1531,N_1499);
or U1939 (N_1939,N_1680,N_1664);
and U1940 (N_1940,N_1417,N_1767);
or U1941 (N_1941,N_1296,N_1739);
nand U1942 (N_1942,N_1449,N_1733);
xor U1943 (N_1943,N_1551,N_1351);
or U1944 (N_1944,N_1450,N_1210);
nand U1945 (N_1945,N_1525,N_1742);
nor U1946 (N_1946,N_1395,N_1389);
nand U1947 (N_1947,N_1784,N_1603);
or U1948 (N_1948,N_1225,N_1564);
nor U1949 (N_1949,N_1584,N_1419);
nor U1950 (N_1950,N_1540,N_1625);
nor U1951 (N_1951,N_1340,N_1407);
nand U1952 (N_1952,N_1409,N_1658);
nor U1953 (N_1953,N_1412,N_1359);
nand U1954 (N_1954,N_1216,N_1762);
or U1955 (N_1955,N_1790,N_1711);
nand U1956 (N_1956,N_1380,N_1571);
or U1957 (N_1957,N_1410,N_1741);
or U1958 (N_1958,N_1550,N_1392);
or U1959 (N_1959,N_1573,N_1369);
nand U1960 (N_1960,N_1473,N_1378);
or U1961 (N_1961,N_1621,N_1200);
or U1962 (N_1962,N_1263,N_1420);
nor U1963 (N_1963,N_1326,N_1278);
nor U1964 (N_1964,N_1787,N_1520);
and U1965 (N_1965,N_1671,N_1785);
xor U1966 (N_1966,N_1476,N_1413);
nor U1967 (N_1967,N_1725,N_1605);
nor U1968 (N_1968,N_1471,N_1776);
and U1969 (N_1969,N_1780,N_1468);
and U1970 (N_1970,N_1675,N_1460);
nor U1971 (N_1971,N_1416,N_1470);
nor U1972 (N_1972,N_1619,N_1283);
or U1973 (N_1973,N_1684,N_1791);
nand U1974 (N_1974,N_1526,N_1727);
or U1975 (N_1975,N_1758,N_1677);
nand U1976 (N_1976,N_1405,N_1323);
and U1977 (N_1977,N_1523,N_1610);
nand U1978 (N_1978,N_1674,N_1644);
nand U1979 (N_1979,N_1650,N_1614);
or U1980 (N_1980,N_1267,N_1788);
nand U1981 (N_1981,N_1797,N_1747);
nor U1982 (N_1982,N_1703,N_1437);
or U1983 (N_1983,N_1646,N_1779);
nand U1984 (N_1984,N_1310,N_1466);
nand U1985 (N_1985,N_1366,N_1472);
nand U1986 (N_1986,N_1710,N_1311);
nor U1987 (N_1987,N_1381,N_1370);
nand U1988 (N_1988,N_1287,N_1536);
xor U1989 (N_1989,N_1291,N_1222);
xor U1990 (N_1990,N_1657,N_1743);
nor U1991 (N_1991,N_1732,N_1434);
and U1992 (N_1992,N_1231,N_1620);
or U1993 (N_1993,N_1297,N_1203);
nor U1994 (N_1994,N_1714,N_1697);
and U1995 (N_1995,N_1565,N_1613);
nand U1996 (N_1996,N_1507,N_1415);
and U1997 (N_1997,N_1382,N_1508);
nand U1998 (N_1998,N_1757,N_1237);
nor U1999 (N_1999,N_1521,N_1338);
or U2000 (N_2000,N_1549,N_1582);
nand U2001 (N_2001,N_1465,N_1516);
nand U2002 (N_2002,N_1682,N_1427);
nand U2003 (N_2003,N_1360,N_1317);
nand U2004 (N_2004,N_1581,N_1505);
nor U2005 (N_2005,N_1217,N_1242);
nand U2006 (N_2006,N_1702,N_1792);
or U2007 (N_2007,N_1488,N_1396);
nor U2008 (N_2008,N_1372,N_1606);
nand U2009 (N_2009,N_1294,N_1665);
nor U2010 (N_2010,N_1752,N_1408);
nand U2011 (N_2011,N_1301,N_1330);
and U2012 (N_2012,N_1209,N_1441);
nand U2013 (N_2013,N_1299,N_1709);
or U2014 (N_2014,N_1315,N_1229);
nor U2015 (N_2015,N_1585,N_1252);
xnor U2016 (N_2016,N_1438,N_1388);
or U2017 (N_2017,N_1230,N_1341);
nand U2018 (N_2018,N_1729,N_1241);
nor U2019 (N_2019,N_1485,N_1716);
and U2020 (N_2020,N_1208,N_1647);
nor U2021 (N_2021,N_1464,N_1213);
xor U2022 (N_2022,N_1524,N_1398);
xor U2023 (N_2023,N_1320,N_1626);
and U2024 (N_2024,N_1467,N_1423);
or U2025 (N_2025,N_1548,N_1484);
or U2026 (N_2026,N_1662,N_1661);
or U2027 (N_2027,N_1575,N_1777);
or U2028 (N_2028,N_1276,N_1277);
nand U2029 (N_2029,N_1799,N_1566);
xor U2030 (N_2030,N_1480,N_1349);
and U2031 (N_2031,N_1772,N_1561);
or U2032 (N_2032,N_1211,N_1493);
or U2033 (N_2033,N_1462,N_1586);
and U2034 (N_2034,N_1256,N_1245);
or U2035 (N_2035,N_1433,N_1204);
and U2036 (N_2036,N_1399,N_1655);
and U2037 (N_2037,N_1612,N_1257);
or U2038 (N_2038,N_1233,N_1685);
and U2039 (N_2039,N_1235,N_1327);
and U2040 (N_2040,N_1692,N_1636);
and U2041 (N_2041,N_1362,N_1737);
xor U2042 (N_2042,N_1442,N_1673);
nor U2043 (N_2043,N_1676,N_1446);
nand U2044 (N_2044,N_1578,N_1734);
nand U2045 (N_2045,N_1356,N_1240);
or U2046 (N_2046,N_1214,N_1292);
or U2047 (N_2047,N_1696,N_1558);
and U2048 (N_2048,N_1572,N_1609);
nand U2049 (N_2049,N_1781,N_1251);
nand U2050 (N_2050,N_1719,N_1774);
or U2051 (N_2051,N_1511,N_1482);
nor U2052 (N_2052,N_1300,N_1224);
or U2053 (N_2053,N_1265,N_1365);
xor U2054 (N_2054,N_1510,N_1498);
or U2055 (N_2055,N_1343,N_1683);
and U2056 (N_2056,N_1492,N_1539);
or U2057 (N_2057,N_1391,N_1594);
or U2058 (N_2058,N_1248,N_1250);
nor U2059 (N_2059,N_1334,N_1249);
or U2060 (N_2060,N_1387,N_1312);
nor U2061 (N_2061,N_1228,N_1559);
and U2062 (N_2062,N_1541,N_1766);
nand U2063 (N_2063,N_1361,N_1736);
or U2064 (N_2064,N_1795,N_1724);
nand U2065 (N_2065,N_1589,N_1459);
nor U2066 (N_2066,N_1793,N_1794);
xor U2067 (N_2067,N_1394,N_1458);
and U2068 (N_2068,N_1611,N_1354);
xnor U2069 (N_2069,N_1652,N_1247);
nand U2070 (N_2070,N_1726,N_1422);
and U2071 (N_2071,N_1704,N_1477);
or U2072 (N_2072,N_1608,N_1718);
or U2073 (N_2073,N_1786,N_1496);
and U2074 (N_2074,N_1515,N_1688);
nor U2075 (N_2075,N_1316,N_1368);
nand U2076 (N_2076,N_1519,N_1273);
xor U2077 (N_2077,N_1261,N_1282);
or U2078 (N_2078,N_1783,N_1670);
nor U2079 (N_2079,N_1563,N_1699);
and U2080 (N_2080,N_1202,N_1201);
nand U2081 (N_2081,N_1637,N_1418);
nor U2082 (N_2082,N_1700,N_1325);
nor U2083 (N_2083,N_1268,N_1494);
and U2084 (N_2084,N_1715,N_1666);
nand U2085 (N_2085,N_1355,N_1553);
nand U2086 (N_2086,N_1306,N_1560);
and U2087 (N_2087,N_1347,N_1720);
xor U2088 (N_2088,N_1775,N_1506);
xnor U2089 (N_2089,N_1350,N_1400);
nand U2090 (N_2090,N_1457,N_1759);
nand U2091 (N_2091,N_1562,N_1455);
and U2092 (N_2092,N_1668,N_1401);
or U2093 (N_2093,N_1329,N_1444);
or U2094 (N_2094,N_1527,N_1414);
xnor U2095 (N_2095,N_1769,N_1542);
and U2096 (N_2096,N_1768,N_1627);
or U2097 (N_2097,N_1286,N_1486);
xor U2098 (N_2098,N_1577,N_1653);
and U2099 (N_2099,N_1517,N_1600);
or U2100 (N_2100,N_1329,N_1622);
and U2101 (N_2101,N_1378,N_1292);
nor U2102 (N_2102,N_1274,N_1593);
and U2103 (N_2103,N_1314,N_1726);
nor U2104 (N_2104,N_1461,N_1733);
xnor U2105 (N_2105,N_1769,N_1618);
nand U2106 (N_2106,N_1418,N_1781);
nand U2107 (N_2107,N_1311,N_1650);
nand U2108 (N_2108,N_1553,N_1204);
or U2109 (N_2109,N_1704,N_1237);
nand U2110 (N_2110,N_1664,N_1268);
or U2111 (N_2111,N_1714,N_1234);
nor U2112 (N_2112,N_1742,N_1416);
and U2113 (N_2113,N_1291,N_1635);
or U2114 (N_2114,N_1545,N_1546);
nor U2115 (N_2115,N_1539,N_1705);
and U2116 (N_2116,N_1467,N_1514);
nor U2117 (N_2117,N_1580,N_1492);
nand U2118 (N_2118,N_1238,N_1692);
xor U2119 (N_2119,N_1427,N_1758);
nor U2120 (N_2120,N_1604,N_1387);
or U2121 (N_2121,N_1247,N_1444);
and U2122 (N_2122,N_1462,N_1559);
nand U2123 (N_2123,N_1705,N_1403);
or U2124 (N_2124,N_1567,N_1794);
and U2125 (N_2125,N_1253,N_1522);
or U2126 (N_2126,N_1238,N_1583);
and U2127 (N_2127,N_1384,N_1599);
nor U2128 (N_2128,N_1754,N_1371);
xor U2129 (N_2129,N_1350,N_1273);
nand U2130 (N_2130,N_1260,N_1645);
nand U2131 (N_2131,N_1303,N_1365);
or U2132 (N_2132,N_1613,N_1454);
nand U2133 (N_2133,N_1424,N_1660);
xor U2134 (N_2134,N_1417,N_1418);
xnor U2135 (N_2135,N_1699,N_1459);
xnor U2136 (N_2136,N_1773,N_1640);
and U2137 (N_2137,N_1265,N_1444);
or U2138 (N_2138,N_1374,N_1353);
and U2139 (N_2139,N_1753,N_1440);
nor U2140 (N_2140,N_1722,N_1302);
or U2141 (N_2141,N_1385,N_1434);
nand U2142 (N_2142,N_1500,N_1762);
and U2143 (N_2143,N_1340,N_1672);
nor U2144 (N_2144,N_1689,N_1719);
or U2145 (N_2145,N_1226,N_1200);
nand U2146 (N_2146,N_1404,N_1745);
nor U2147 (N_2147,N_1472,N_1495);
nand U2148 (N_2148,N_1542,N_1304);
or U2149 (N_2149,N_1629,N_1785);
xor U2150 (N_2150,N_1411,N_1551);
nor U2151 (N_2151,N_1252,N_1299);
nand U2152 (N_2152,N_1794,N_1676);
and U2153 (N_2153,N_1602,N_1573);
and U2154 (N_2154,N_1792,N_1503);
and U2155 (N_2155,N_1552,N_1568);
or U2156 (N_2156,N_1590,N_1310);
or U2157 (N_2157,N_1460,N_1464);
xor U2158 (N_2158,N_1563,N_1477);
nor U2159 (N_2159,N_1250,N_1724);
or U2160 (N_2160,N_1371,N_1783);
nor U2161 (N_2161,N_1514,N_1258);
nor U2162 (N_2162,N_1457,N_1453);
nor U2163 (N_2163,N_1254,N_1411);
nand U2164 (N_2164,N_1228,N_1710);
nand U2165 (N_2165,N_1711,N_1703);
or U2166 (N_2166,N_1400,N_1724);
nand U2167 (N_2167,N_1351,N_1414);
or U2168 (N_2168,N_1528,N_1559);
nand U2169 (N_2169,N_1447,N_1468);
or U2170 (N_2170,N_1302,N_1743);
or U2171 (N_2171,N_1678,N_1268);
nand U2172 (N_2172,N_1613,N_1510);
or U2173 (N_2173,N_1296,N_1209);
xor U2174 (N_2174,N_1374,N_1544);
and U2175 (N_2175,N_1743,N_1371);
or U2176 (N_2176,N_1294,N_1798);
xor U2177 (N_2177,N_1696,N_1782);
nand U2178 (N_2178,N_1769,N_1249);
and U2179 (N_2179,N_1580,N_1790);
nand U2180 (N_2180,N_1443,N_1418);
and U2181 (N_2181,N_1651,N_1447);
nand U2182 (N_2182,N_1407,N_1544);
nand U2183 (N_2183,N_1646,N_1381);
nand U2184 (N_2184,N_1355,N_1358);
and U2185 (N_2185,N_1763,N_1271);
xnor U2186 (N_2186,N_1211,N_1553);
and U2187 (N_2187,N_1556,N_1661);
nor U2188 (N_2188,N_1465,N_1549);
or U2189 (N_2189,N_1672,N_1620);
nand U2190 (N_2190,N_1573,N_1638);
nand U2191 (N_2191,N_1442,N_1591);
or U2192 (N_2192,N_1715,N_1357);
or U2193 (N_2193,N_1392,N_1697);
and U2194 (N_2194,N_1703,N_1754);
or U2195 (N_2195,N_1791,N_1257);
nor U2196 (N_2196,N_1210,N_1256);
xnor U2197 (N_2197,N_1317,N_1625);
nand U2198 (N_2198,N_1652,N_1591);
nand U2199 (N_2199,N_1598,N_1721);
nor U2200 (N_2200,N_1522,N_1438);
nand U2201 (N_2201,N_1551,N_1676);
or U2202 (N_2202,N_1629,N_1560);
and U2203 (N_2203,N_1522,N_1728);
or U2204 (N_2204,N_1518,N_1265);
nand U2205 (N_2205,N_1278,N_1761);
or U2206 (N_2206,N_1508,N_1326);
and U2207 (N_2207,N_1403,N_1490);
or U2208 (N_2208,N_1300,N_1470);
nand U2209 (N_2209,N_1558,N_1541);
nand U2210 (N_2210,N_1231,N_1488);
nand U2211 (N_2211,N_1698,N_1408);
and U2212 (N_2212,N_1649,N_1363);
nand U2213 (N_2213,N_1282,N_1252);
nand U2214 (N_2214,N_1535,N_1563);
nor U2215 (N_2215,N_1415,N_1384);
xnor U2216 (N_2216,N_1271,N_1747);
nand U2217 (N_2217,N_1548,N_1790);
and U2218 (N_2218,N_1764,N_1478);
nor U2219 (N_2219,N_1619,N_1280);
xor U2220 (N_2220,N_1629,N_1634);
nand U2221 (N_2221,N_1593,N_1618);
nand U2222 (N_2222,N_1357,N_1372);
or U2223 (N_2223,N_1689,N_1582);
nor U2224 (N_2224,N_1546,N_1317);
nor U2225 (N_2225,N_1291,N_1496);
or U2226 (N_2226,N_1344,N_1793);
or U2227 (N_2227,N_1647,N_1623);
or U2228 (N_2228,N_1312,N_1318);
xor U2229 (N_2229,N_1549,N_1783);
and U2230 (N_2230,N_1619,N_1319);
nand U2231 (N_2231,N_1304,N_1680);
nand U2232 (N_2232,N_1484,N_1235);
and U2233 (N_2233,N_1775,N_1353);
and U2234 (N_2234,N_1787,N_1630);
xnor U2235 (N_2235,N_1598,N_1570);
and U2236 (N_2236,N_1267,N_1655);
nand U2237 (N_2237,N_1286,N_1511);
and U2238 (N_2238,N_1287,N_1628);
and U2239 (N_2239,N_1598,N_1250);
nand U2240 (N_2240,N_1587,N_1595);
or U2241 (N_2241,N_1658,N_1743);
nor U2242 (N_2242,N_1585,N_1629);
nor U2243 (N_2243,N_1246,N_1218);
and U2244 (N_2244,N_1654,N_1571);
nor U2245 (N_2245,N_1609,N_1251);
or U2246 (N_2246,N_1792,N_1542);
nand U2247 (N_2247,N_1568,N_1798);
nand U2248 (N_2248,N_1256,N_1714);
or U2249 (N_2249,N_1504,N_1491);
nor U2250 (N_2250,N_1703,N_1265);
and U2251 (N_2251,N_1615,N_1736);
nand U2252 (N_2252,N_1774,N_1540);
and U2253 (N_2253,N_1705,N_1508);
and U2254 (N_2254,N_1550,N_1470);
and U2255 (N_2255,N_1693,N_1518);
nand U2256 (N_2256,N_1411,N_1488);
and U2257 (N_2257,N_1737,N_1343);
or U2258 (N_2258,N_1251,N_1350);
nor U2259 (N_2259,N_1720,N_1391);
nor U2260 (N_2260,N_1790,N_1438);
nand U2261 (N_2261,N_1241,N_1749);
nor U2262 (N_2262,N_1642,N_1491);
nand U2263 (N_2263,N_1305,N_1313);
xor U2264 (N_2264,N_1791,N_1419);
nand U2265 (N_2265,N_1279,N_1585);
nor U2266 (N_2266,N_1627,N_1260);
and U2267 (N_2267,N_1233,N_1218);
or U2268 (N_2268,N_1278,N_1604);
or U2269 (N_2269,N_1295,N_1718);
or U2270 (N_2270,N_1473,N_1667);
or U2271 (N_2271,N_1701,N_1568);
and U2272 (N_2272,N_1364,N_1684);
or U2273 (N_2273,N_1309,N_1554);
nor U2274 (N_2274,N_1252,N_1512);
nor U2275 (N_2275,N_1587,N_1772);
nor U2276 (N_2276,N_1605,N_1573);
nand U2277 (N_2277,N_1511,N_1455);
xnor U2278 (N_2278,N_1421,N_1712);
nand U2279 (N_2279,N_1735,N_1391);
and U2280 (N_2280,N_1417,N_1612);
nor U2281 (N_2281,N_1240,N_1780);
nor U2282 (N_2282,N_1245,N_1551);
nand U2283 (N_2283,N_1407,N_1354);
or U2284 (N_2284,N_1228,N_1658);
nand U2285 (N_2285,N_1651,N_1677);
nor U2286 (N_2286,N_1264,N_1789);
and U2287 (N_2287,N_1250,N_1703);
nor U2288 (N_2288,N_1721,N_1793);
nor U2289 (N_2289,N_1551,N_1693);
or U2290 (N_2290,N_1315,N_1246);
nand U2291 (N_2291,N_1688,N_1218);
nand U2292 (N_2292,N_1404,N_1609);
nand U2293 (N_2293,N_1641,N_1341);
and U2294 (N_2294,N_1360,N_1576);
nor U2295 (N_2295,N_1316,N_1285);
and U2296 (N_2296,N_1650,N_1526);
nand U2297 (N_2297,N_1774,N_1507);
xor U2298 (N_2298,N_1253,N_1441);
and U2299 (N_2299,N_1346,N_1600);
xnor U2300 (N_2300,N_1623,N_1573);
xor U2301 (N_2301,N_1501,N_1686);
xnor U2302 (N_2302,N_1449,N_1290);
nand U2303 (N_2303,N_1627,N_1671);
or U2304 (N_2304,N_1729,N_1475);
nor U2305 (N_2305,N_1542,N_1289);
and U2306 (N_2306,N_1427,N_1680);
or U2307 (N_2307,N_1267,N_1581);
nand U2308 (N_2308,N_1344,N_1675);
nand U2309 (N_2309,N_1575,N_1220);
nor U2310 (N_2310,N_1726,N_1678);
and U2311 (N_2311,N_1412,N_1581);
and U2312 (N_2312,N_1481,N_1424);
nor U2313 (N_2313,N_1713,N_1563);
or U2314 (N_2314,N_1378,N_1641);
xor U2315 (N_2315,N_1204,N_1426);
nand U2316 (N_2316,N_1213,N_1266);
nand U2317 (N_2317,N_1405,N_1644);
and U2318 (N_2318,N_1759,N_1551);
nor U2319 (N_2319,N_1306,N_1645);
nand U2320 (N_2320,N_1790,N_1613);
or U2321 (N_2321,N_1601,N_1720);
nor U2322 (N_2322,N_1202,N_1450);
xor U2323 (N_2323,N_1570,N_1233);
or U2324 (N_2324,N_1244,N_1324);
and U2325 (N_2325,N_1229,N_1705);
nand U2326 (N_2326,N_1424,N_1244);
nor U2327 (N_2327,N_1496,N_1414);
or U2328 (N_2328,N_1485,N_1703);
or U2329 (N_2329,N_1540,N_1289);
nand U2330 (N_2330,N_1507,N_1647);
or U2331 (N_2331,N_1650,N_1253);
or U2332 (N_2332,N_1521,N_1481);
nand U2333 (N_2333,N_1374,N_1604);
and U2334 (N_2334,N_1735,N_1411);
and U2335 (N_2335,N_1305,N_1317);
or U2336 (N_2336,N_1406,N_1438);
or U2337 (N_2337,N_1466,N_1519);
nand U2338 (N_2338,N_1696,N_1748);
and U2339 (N_2339,N_1505,N_1383);
nor U2340 (N_2340,N_1488,N_1323);
or U2341 (N_2341,N_1575,N_1280);
and U2342 (N_2342,N_1315,N_1597);
or U2343 (N_2343,N_1630,N_1355);
nand U2344 (N_2344,N_1617,N_1344);
xor U2345 (N_2345,N_1451,N_1392);
or U2346 (N_2346,N_1263,N_1701);
nor U2347 (N_2347,N_1301,N_1777);
nand U2348 (N_2348,N_1669,N_1640);
nand U2349 (N_2349,N_1208,N_1576);
and U2350 (N_2350,N_1545,N_1240);
nor U2351 (N_2351,N_1595,N_1323);
and U2352 (N_2352,N_1779,N_1732);
and U2353 (N_2353,N_1346,N_1313);
nand U2354 (N_2354,N_1418,N_1560);
nand U2355 (N_2355,N_1520,N_1762);
or U2356 (N_2356,N_1275,N_1320);
or U2357 (N_2357,N_1504,N_1325);
nand U2358 (N_2358,N_1206,N_1648);
and U2359 (N_2359,N_1493,N_1227);
or U2360 (N_2360,N_1250,N_1448);
or U2361 (N_2361,N_1693,N_1592);
nor U2362 (N_2362,N_1674,N_1371);
xnor U2363 (N_2363,N_1371,N_1540);
nor U2364 (N_2364,N_1387,N_1221);
or U2365 (N_2365,N_1647,N_1309);
or U2366 (N_2366,N_1602,N_1433);
nor U2367 (N_2367,N_1291,N_1577);
and U2368 (N_2368,N_1677,N_1467);
and U2369 (N_2369,N_1505,N_1594);
and U2370 (N_2370,N_1340,N_1674);
nor U2371 (N_2371,N_1492,N_1466);
xnor U2372 (N_2372,N_1628,N_1275);
or U2373 (N_2373,N_1412,N_1563);
and U2374 (N_2374,N_1200,N_1453);
and U2375 (N_2375,N_1744,N_1380);
nor U2376 (N_2376,N_1736,N_1552);
and U2377 (N_2377,N_1597,N_1677);
and U2378 (N_2378,N_1283,N_1502);
nand U2379 (N_2379,N_1240,N_1360);
nor U2380 (N_2380,N_1349,N_1446);
xor U2381 (N_2381,N_1343,N_1698);
xnor U2382 (N_2382,N_1377,N_1477);
and U2383 (N_2383,N_1649,N_1657);
nand U2384 (N_2384,N_1256,N_1773);
or U2385 (N_2385,N_1763,N_1453);
nand U2386 (N_2386,N_1796,N_1474);
nand U2387 (N_2387,N_1372,N_1404);
xor U2388 (N_2388,N_1227,N_1435);
or U2389 (N_2389,N_1260,N_1629);
and U2390 (N_2390,N_1523,N_1699);
nand U2391 (N_2391,N_1675,N_1530);
nor U2392 (N_2392,N_1508,N_1577);
nor U2393 (N_2393,N_1347,N_1636);
nor U2394 (N_2394,N_1671,N_1502);
nand U2395 (N_2395,N_1741,N_1625);
and U2396 (N_2396,N_1760,N_1349);
nor U2397 (N_2397,N_1460,N_1376);
xnor U2398 (N_2398,N_1742,N_1567);
nor U2399 (N_2399,N_1598,N_1443);
or U2400 (N_2400,N_2250,N_1842);
nand U2401 (N_2401,N_1943,N_2278);
nand U2402 (N_2402,N_2169,N_2343);
nor U2403 (N_2403,N_2310,N_2206);
nor U2404 (N_2404,N_1925,N_2370);
nand U2405 (N_2405,N_2255,N_2109);
xnor U2406 (N_2406,N_2339,N_2311);
nand U2407 (N_2407,N_2285,N_1900);
or U2408 (N_2408,N_1879,N_1852);
and U2409 (N_2409,N_2092,N_1805);
and U2410 (N_2410,N_2194,N_2047);
nor U2411 (N_2411,N_1888,N_2275);
or U2412 (N_2412,N_1839,N_1807);
nand U2413 (N_2413,N_2234,N_2007);
and U2414 (N_2414,N_2034,N_2006);
and U2415 (N_2415,N_1959,N_2241);
nand U2416 (N_2416,N_2280,N_1941);
and U2417 (N_2417,N_2238,N_2178);
or U2418 (N_2418,N_2113,N_2367);
and U2419 (N_2419,N_1902,N_2071);
nor U2420 (N_2420,N_1808,N_2333);
nor U2421 (N_2421,N_1944,N_1806);
or U2422 (N_2422,N_2216,N_2145);
nand U2423 (N_2423,N_2325,N_2028);
and U2424 (N_2424,N_2291,N_2322);
or U2425 (N_2425,N_1969,N_2381);
nand U2426 (N_2426,N_2271,N_2055);
and U2427 (N_2427,N_2033,N_1967);
xnor U2428 (N_2428,N_1955,N_1843);
nor U2429 (N_2429,N_1878,N_1980);
and U2430 (N_2430,N_2363,N_2116);
nand U2431 (N_2431,N_1846,N_2282);
and U2432 (N_2432,N_2096,N_1896);
or U2433 (N_2433,N_2170,N_2215);
nor U2434 (N_2434,N_2098,N_2171);
and U2435 (N_2435,N_2036,N_1913);
and U2436 (N_2436,N_2064,N_2375);
nor U2437 (N_2437,N_2091,N_2154);
nor U2438 (N_2438,N_2199,N_2252);
nand U2439 (N_2439,N_2393,N_2382);
nand U2440 (N_2440,N_2023,N_2131);
nand U2441 (N_2441,N_2203,N_2321);
or U2442 (N_2442,N_2352,N_2383);
and U2443 (N_2443,N_2051,N_1811);
nor U2444 (N_2444,N_2144,N_2164);
nor U2445 (N_2445,N_2121,N_2002);
and U2446 (N_2446,N_2021,N_1826);
nor U2447 (N_2447,N_2218,N_1869);
nand U2448 (N_2448,N_1911,N_1928);
and U2449 (N_2449,N_2386,N_1887);
xnor U2450 (N_2450,N_2157,N_2069);
xnor U2451 (N_2451,N_1834,N_2084);
nor U2452 (N_2452,N_2156,N_2118);
or U2453 (N_2453,N_2079,N_2384);
xnor U2454 (N_2454,N_2320,N_2112);
nor U2455 (N_2455,N_2229,N_2290);
xnor U2456 (N_2456,N_2102,N_1990);
and U2457 (N_2457,N_2026,N_1853);
xnor U2458 (N_2458,N_2014,N_2262);
and U2459 (N_2459,N_1978,N_2004);
or U2460 (N_2460,N_2293,N_2183);
nand U2461 (N_2461,N_2269,N_2168);
xnor U2462 (N_2462,N_1858,N_1817);
or U2463 (N_2463,N_2334,N_2346);
nand U2464 (N_2464,N_1857,N_1872);
and U2465 (N_2465,N_2289,N_1971);
and U2466 (N_2466,N_1833,N_2000);
xor U2467 (N_2467,N_1828,N_1939);
xor U2468 (N_2468,N_2101,N_2374);
and U2469 (N_2469,N_1931,N_2324);
or U2470 (N_2470,N_1821,N_2056);
or U2471 (N_2471,N_2366,N_2158);
nor U2472 (N_2472,N_1914,N_1988);
or U2473 (N_2473,N_2176,N_2314);
or U2474 (N_2474,N_2240,N_1835);
nand U2475 (N_2475,N_2249,N_2057);
and U2476 (N_2476,N_2394,N_1915);
nand U2477 (N_2477,N_2181,N_2015);
nor U2478 (N_2478,N_2080,N_1844);
nor U2479 (N_2479,N_2088,N_2326);
nor U2480 (N_2480,N_2224,N_2013);
or U2481 (N_2481,N_2053,N_1832);
nand U2482 (N_2482,N_2122,N_2354);
and U2483 (N_2483,N_2242,N_2342);
nand U2484 (N_2484,N_2070,N_1917);
or U2485 (N_2485,N_1877,N_1875);
and U2486 (N_2486,N_1940,N_2274);
and U2487 (N_2487,N_1950,N_2040);
or U2488 (N_2488,N_2368,N_2175);
nor U2489 (N_2489,N_2348,N_2010);
xnor U2490 (N_2490,N_2086,N_2319);
nor U2491 (N_2491,N_2305,N_2042);
or U2492 (N_2492,N_1934,N_2373);
xor U2493 (N_2493,N_2141,N_2344);
xor U2494 (N_2494,N_2152,N_2085);
nand U2495 (N_2495,N_1983,N_1937);
nand U2496 (N_2496,N_2295,N_1957);
or U2497 (N_2497,N_1822,N_1809);
or U2498 (N_2498,N_2254,N_1840);
xor U2499 (N_2499,N_1927,N_1863);
xor U2500 (N_2500,N_2286,N_1836);
nand U2501 (N_2501,N_1970,N_1948);
nor U2502 (N_2502,N_2035,N_2193);
nand U2503 (N_2503,N_2399,N_2349);
and U2504 (N_2504,N_2020,N_1901);
nand U2505 (N_2505,N_2336,N_2068);
nand U2506 (N_2506,N_2331,N_2073);
nand U2507 (N_2507,N_1945,N_2153);
nor U2508 (N_2508,N_2233,N_1964);
nor U2509 (N_2509,N_2162,N_2037);
xnor U2510 (N_2510,N_1906,N_2202);
xnor U2511 (N_2511,N_2287,N_2371);
and U2512 (N_2512,N_2253,N_1841);
xnor U2513 (N_2513,N_2220,N_1803);
nand U2514 (N_2514,N_2385,N_2298);
nand U2515 (N_2515,N_2396,N_2221);
or U2516 (N_2516,N_1890,N_2207);
nor U2517 (N_2517,N_2312,N_2256);
nand U2518 (N_2518,N_2043,N_1947);
and U2519 (N_2519,N_1989,N_1831);
nor U2520 (N_2520,N_1953,N_1968);
nor U2521 (N_2521,N_1992,N_2188);
and U2522 (N_2522,N_1800,N_1812);
and U2523 (N_2523,N_1856,N_2066);
nand U2524 (N_2524,N_2140,N_2243);
nand U2525 (N_2525,N_1997,N_1973);
nor U2526 (N_2526,N_1825,N_2059);
and U2527 (N_2527,N_2378,N_2222);
and U2528 (N_2528,N_2192,N_2302);
or U2529 (N_2529,N_2273,N_2327);
nor U2530 (N_2530,N_2095,N_2226);
xor U2531 (N_2531,N_2029,N_2044);
nor U2532 (N_2532,N_2230,N_2317);
nor U2533 (N_2533,N_1966,N_2315);
nand U2534 (N_2534,N_1854,N_1999);
xor U2535 (N_2535,N_1910,N_2306);
nor U2536 (N_2536,N_1895,N_1884);
nand U2537 (N_2537,N_2045,N_2197);
nand U2538 (N_2538,N_1975,N_2318);
nand U2539 (N_2539,N_2265,N_1838);
nor U2540 (N_2540,N_2329,N_2398);
and U2541 (N_2541,N_2263,N_1848);
or U2542 (N_2542,N_2087,N_2227);
nand U2543 (N_2543,N_2397,N_2372);
xor U2544 (N_2544,N_1982,N_2143);
and U2545 (N_2545,N_2089,N_1918);
xnor U2546 (N_2546,N_2281,N_2106);
nand U2547 (N_2547,N_2150,N_2313);
or U2548 (N_2548,N_2038,N_1804);
or U2549 (N_2549,N_2135,N_1951);
nor U2550 (N_2550,N_2046,N_2142);
nor U2551 (N_2551,N_1837,N_2090);
nor U2552 (N_2552,N_2261,N_1880);
and U2553 (N_2553,N_2165,N_2332);
nand U2554 (N_2554,N_2097,N_2294);
nand U2555 (N_2555,N_2389,N_1889);
xor U2556 (N_2556,N_2134,N_2030);
or U2557 (N_2557,N_2107,N_2167);
nor U2558 (N_2558,N_2210,N_1851);
or U2559 (N_2559,N_1904,N_2304);
nand U2560 (N_2560,N_1985,N_1933);
xnor U2561 (N_2561,N_2223,N_2205);
and U2562 (N_2562,N_1824,N_1823);
nand U2563 (N_2563,N_2187,N_2151);
or U2564 (N_2564,N_2105,N_1886);
and U2565 (N_2565,N_1962,N_2211);
nand U2566 (N_2566,N_1958,N_1829);
or U2567 (N_2567,N_2180,N_2099);
nand U2568 (N_2568,N_1802,N_2369);
and U2569 (N_2569,N_1867,N_2377);
and U2570 (N_2570,N_1998,N_2024);
or U2571 (N_2571,N_2075,N_2054);
nor U2572 (N_2572,N_2387,N_1907);
and U2573 (N_2573,N_1952,N_2364);
and U2574 (N_2574,N_2359,N_1882);
nand U2575 (N_2575,N_2232,N_1814);
or U2576 (N_2576,N_2127,N_2365);
nand U2577 (N_2577,N_2048,N_2076);
or U2578 (N_2578,N_1898,N_1894);
nand U2579 (N_2579,N_2228,N_2128);
and U2580 (N_2580,N_2061,N_2357);
and U2581 (N_2581,N_1908,N_1827);
or U2582 (N_2582,N_2132,N_2001);
or U2583 (N_2583,N_2063,N_2246);
or U2584 (N_2584,N_1965,N_2270);
xor U2585 (N_2585,N_1899,N_1946);
nand U2586 (N_2586,N_2077,N_2258);
nand U2587 (N_2587,N_2173,N_2355);
or U2588 (N_2588,N_1954,N_2245);
or U2589 (N_2589,N_2277,N_1949);
and U2590 (N_2590,N_2161,N_2082);
or U2591 (N_2591,N_1986,N_2303);
nand U2592 (N_2592,N_2138,N_2209);
and U2593 (N_2593,N_2148,N_2239);
nor U2594 (N_2594,N_2005,N_1942);
and U2595 (N_2595,N_2078,N_2016);
and U2596 (N_2596,N_1864,N_2264);
or U2597 (N_2597,N_2388,N_1850);
nand U2598 (N_2598,N_2231,N_1815);
xnor U2599 (N_2599,N_2266,N_2247);
and U2600 (N_2600,N_1859,N_2012);
or U2601 (N_2601,N_1926,N_2074);
nor U2602 (N_2602,N_2114,N_1974);
nand U2603 (N_2603,N_1972,N_2031);
nand U2604 (N_2604,N_2213,N_1921);
nor U2605 (N_2605,N_1868,N_2185);
or U2606 (N_2606,N_1938,N_2126);
xnor U2607 (N_2607,N_1881,N_2177);
and U2608 (N_2608,N_2201,N_1893);
or U2609 (N_2609,N_1916,N_1984);
and U2610 (N_2610,N_2330,N_1874);
or U2611 (N_2611,N_2083,N_1987);
nor U2612 (N_2612,N_1995,N_2050);
nor U2613 (N_2613,N_2119,N_2019);
or U2614 (N_2614,N_2186,N_1905);
or U2615 (N_2615,N_2117,N_2093);
nand U2616 (N_2616,N_1861,N_1930);
and U2617 (N_2617,N_2251,N_1993);
and U2618 (N_2618,N_2353,N_2395);
nand U2619 (N_2619,N_2166,N_2284);
and U2620 (N_2620,N_2125,N_2335);
xor U2621 (N_2621,N_2149,N_1845);
nor U2622 (N_2622,N_2267,N_2139);
or U2623 (N_2623,N_1891,N_2276);
and U2624 (N_2624,N_2316,N_1924);
and U2625 (N_2625,N_1847,N_2376);
and U2626 (N_2626,N_2137,N_1996);
or U2627 (N_2627,N_2308,N_2337);
nor U2628 (N_2628,N_1923,N_2296);
xnor U2629 (N_2629,N_2356,N_1885);
or U2630 (N_2630,N_1963,N_2350);
or U2631 (N_2631,N_2214,N_1909);
nand U2632 (N_2632,N_2360,N_1830);
or U2633 (N_2633,N_2191,N_1979);
and U2634 (N_2634,N_2184,N_2288);
nor U2635 (N_2635,N_2300,N_2103);
or U2636 (N_2636,N_1849,N_2159);
and U2637 (N_2637,N_2268,N_2236);
and U2638 (N_2638,N_2379,N_2120);
or U2639 (N_2639,N_2338,N_2248);
and U2640 (N_2640,N_2060,N_2146);
nor U2641 (N_2641,N_1871,N_1855);
nor U2642 (N_2642,N_2062,N_2260);
nor U2643 (N_2643,N_2237,N_1865);
nor U2644 (N_2644,N_1897,N_1816);
or U2645 (N_2645,N_2341,N_1801);
or U2646 (N_2646,N_2208,N_2008);
nor U2647 (N_2647,N_2225,N_2217);
nand U2648 (N_2648,N_2307,N_2292);
and U2649 (N_2649,N_2133,N_2259);
or U2650 (N_2650,N_2130,N_1876);
nor U2651 (N_2651,N_2147,N_2041);
nor U2652 (N_2652,N_2198,N_2163);
nor U2653 (N_2653,N_1883,N_2011);
and U2654 (N_2654,N_2039,N_1920);
or U2655 (N_2655,N_1935,N_1862);
nand U2656 (N_2656,N_1819,N_2257);
nand U2657 (N_2657,N_1903,N_2340);
or U2658 (N_2658,N_2328,N_2174);
nor U2659 (N_2659,N_2160,N_2017);
nand U2660 (N_2660,N_2190,N_1932);
nor U2661 (N_2661,N_2018,N_2380);
or U2662 (N_2662,N_2392,N_2182);
nand U2663 (N_2663,N_2179,N_2081);
nor U2664 (N_2664,N_2189,N_2200);
nand U2665 (N_2665,N_2009,N_2052);
nand U2666 (N_2666,N_2111,N_1873);
and U2667 (N_2667,N_2358,N_2049);
or U2668 (N_2668,N_2309,N_2058);
xor U2669 (N_2669,N_2003,N_1994);
and U2670 (N_2670,N_2235,N_2272);
nor U2671 (N_2671,N_2136,N_2065);
nand U2672 (N_2672,N_2124,N_1976);
and U2673 (N_2673,N_1818,N_2100);
xnor U2674 (N_2674,N_1866,N_1870);
xor U2675 (N_2675,N_2195,N_1960);
nand U2676 (N_2676,N_1922,N_2362);
nand U2677 (N_2677,N_2155,N_2022);
and U2678 (N_2678,N_1820,N_2351);
or U2679 (N_2679,N_1936,N_2361);
nor U2680 (N_2680,N_1892,N_2067);
or U2681 (N_2681,N_2204,N_2094);
or U2682 (N_2682,N_2032,N_1860);
or U2683 (N_2683,N_2212,N_2115);
xnor U2684 (N_2684,N_1991,N_2391);
nor U2685 (N_2685,N_1961,N_1956);
nand U2686 (N_2686,N_2108,N_2283);
or U2687 (N_2687,N_2301,N_2110);
nor U2688 (N_2688,N_2345,N_2323);
and U2689 (N_2689,N_2172,N_2299);
nor U2690 (N_2690,N_1929,N_2347);
nor U2691 (N_2691,N_2244,N_1912);
nand U2692 (N_2692,N_2025,N_2297);
xor U2693 (N_2693,N_1810,N_1919);
and U2694 (N_2694,N_2279,N_1813);
or U2695 (N_2695,N_2123,N_2219);
or U2696 (N_2696,N_2129,N_2390);
xnor U2697 (N_2697,N_2196,N_2072);
or U2698 (N_2698,N_2104,N_1977);
nor U2699 (N_2699,N_2027,N_1981);
nor U2700 (N_2700,N_1985,N_2089);
nand U2701 (N_2701,N_2075,N_1803);
and U2702 (N_2702,N_2121,N_2046);
and U2703 (N_2703,N_2039,N_2388);
nor U2704 (N_2704,N_1849,N_2318);
and U2705 (N_2705,N_2058,N_2027);
nor U2706 (N_2706,N_1879,N_2091);
nor U2707 (N_2707,N_2116,N_2203);
nand U2708 (N_2708,N_2399,N_1904);
xor U2709 (N_2709,N_2202,N_2107);
and U2710 (N_2710,N_2189,N_2290);
or U2711 (N_2711,N_2133,N_2364);
xnor U2712 (N_2712,N_2006,N_1920);
nand U2713 (N_2713,N_2360,N_2239);
and U2714 (N_2714,N_2151,N_1845);
xnor U2715 (N_2715,N_2299,N_2062);
nand U2716 (N_2716,N_1851,N_2245);
or U2717 (N_2717,N_2050,N_2293);
or U2718 (N_2718,N_2284,N_2193);
and U2719 (N_2719,N_1997,N_2201);
or U2720 (N_2720,N_1924,N_2041);
nor U2721 (N_2721,N_2017,N_2023);
nor U2722 (N_2722,N_1941,N_2178);
and U2723 (N_2723,N_2393,N_2326);
and U2724 (N_2724,N_2069,N_2293);
nor U2725 (N_2725,N_1925,N_2198);
or U2726 (N_2726,N_2118,N_1955);
nand U2727 (N_2727,N_2266,N_2111);
and U2728 (N_2728,N_2394,N_2269);
and U2729 (N_2729,N_2383,N_2103);
and U2730 (N_2730,N_2122,N_1914);
or U2731 (N_2731,N_1945,N_2232);
nor U2732 (N_2732,N_2130,N_1837);
and U2733 (N_2733,N_2029,N_2387);
and U2734 (N_2734,N_2289,N_2290);
or U2735 (N_2735,N_2105,N_1979);
or U2736 (N_2736,N_2005,N_2073);
and U2737 (N_2737,N_1813,N_2298);
nor U2738 (N_2738,N_2226,N_2051);
and U2739 (N_2739,N_2074,N_1951);
nand U2740 (N_2740,N_2156,N_2250);
nand U2741 (N_2741,N_2346,N_2086);
or U2742 (N_2742,N_2194,N_2013);
nand U2743 (N_2743,N_1986,N_1816);
nor U2744 (N_2744,N_2098,N_2052);
nand U2745 (N_2745,N_2351,N_2202);
and U2746 (N_2746,N_1869,N_2249);
and U2747 (N_2747,N_2050,N_1865);
and U2748 (N_2748,N_1964,N_1917);
and U2749 (N_2749,N_2093,N_2030);
and U2750 (N_2750,N_1902,N_1994);
xor U2751 (N_2751,N_2021,N_2159);
or U2752 (N_2752,N_2097,N_1856);
and U2753 (N_2753,N_2062,N_2084);
or U2754 (N_2754,N_1995,N_2180);
nand U2755 (N_2755,N_2213,N_2081);
nand U2756 (N_2756,N_1896,N_2150);
nand U2757 (N_2757,N_2398,N_2271);
and U2758 (N_2758,N_2331,N_2103);
and U2759 (N_2759,N_2116,N_2112);
or U2760 (N_2760,N_2193,N_1842);
nor U2761 (N_2761,N_2062,N_1813);
or U2762 (N_2762,N_1923,N_2311);
and U2763 (N_2763,N_1835,N_2046);
nand U2764 (N_2764,N_2335,N_1971);
nand U2765 (N_2765,N_1978,N_2156);
and U2766 (N_2766,N_2169,N_2114);
and U2767 (N_2767,N_1907,N_2286);
and U2768 (N_2768,N_2133,N_1914);
nor U2769 (N_2769,N_1879,N_2162);
nand U2770 (N_2770,N_2222,N_2390);
nand U2771 (N_2771,N_1894,N_1889);
nor U2772 (N_2772,N_1864,N_1969);
xnor U2773 (N_2773,N_1915,N_2304);
nor U2774 (N_2774,N_2367,N_1976);
nor U2775 (N_2775,N_2300,N_1810);
nand U2776 (N_2776,N_2349,N_1853);
xor U2777 (N_2777,N_2283,N_2266);
or U2778 (N_2778,N_2164,N_2207);
xor U2779 (N_2779,N_1890,N_2099);
or U2780 (N_2780,N_2228,N_1932);
xor U2781 (N_2781,N_2015,N_2185);
nand U2782 (N_2782,N_1878,N_1948);
and U2783 (N_2783,N_2289,N_1967);
nand U2784 (N_2784,N_1866,N_2217);
or U2785 (N_2785,N_2276,N_2309);
and U2786 (N_2786,N_1881,N_2166);
xor U2787 (N_2787,N_2180,N_2245);
nor U2788 (N_2788,N_2081,N_2182);
xor U2789 (N_2789,N_1825,N_2150);
nor U2790 (N_2790,N_2310,N_2284);
nor U2791 (N_2791,N_1974,N_2284);
nor U2792 (N_2792,N_1960,N_2114);
and U2793 (N_2793,N_1899,N_1853);
xnor U2794 (N_2794,N_2195,N_1833);
nand U2795 (N_2795,N_2059,N_2259);
and U2796 (N_2796,N_1926,N_2035);
nor U2797 (N_2797,N_1815,N_2271);
nor U2798 (N_2798,N_1897,N_2276);
and U2799 (N_2799,N_2082,N_2135);
or U2800 (N_2800,N_1978,N_2012);
or U2801 (N_2801,N_2292,N_2195);
or U2802 (N_2802,N_2166,N_1933);
and U2803 (N_2803,N_2118,N_1947);
nand U2804 (N_2804,N_1971,N_2221);
nor U2805 (N_2805,N_2049,N_2264);
nor U2806 (N_2806,N_2222,N_2384);
and U2807 (N_2807,N_2367,N_2148);
and U2808 (N_2808,N_2379,N_1891);
or U2809 (N_2809,N_2181,N_2348);
nand U2810 (N_2810,N_1850,N_2016);
nor U2811 (N_2811,N_2263,N_2242);
and U2812 (N_2812,N_2383,N_2021);
xor U2813 (N_2813,N_1961,N_1805);
nor U2814 (N_2814,N_2034,N_2327);
nand U2815 (N_2815,N_2104,N_2307);
nand U2816 (N_2816,N_2132,N_2051);
nand U2817 (N_2817,N_2319,N_2350);
nand U2818 (N_2818,N_2063,N_2312);
nand U2819 (N_2819,N_2345,N_2365);
and U2820 (N_2820,N_2197,N_1838);
or U2821 (N_2821,N_1851,N_1841);
or U2822 (N_2822,N_1951,N_1986);
xnor U2823 (N_2823,N_2232,N_2349);
nand U2824 (N_2824,N_2108,N_1879);
or U2825 (N_2825,N_2383,N_2311);
and U2826 (N_2826,N_2128,N_2074);
nand U2827 (N_2827,N_2253,N_2147);
and U2828 (N_2828,N_1807,N_1835);
nand U2829 (N_2829,N_1874,N_1958);
or U2830 (N_2830,N_1937,N_2061);
nand U2831 (N_2831,N_2016,N_2248);
nand U2832 (N_2832,N_1860,N_2351);
or U2833 (N_2833,N_2033,N_1868);
nand U2834 (N_2834,N_2024,N_2131);
nand U2835 (N_2835,N_1807,N_2030);
nand U2836 (N_2836,N_2353,N_2289);
nand U2837 (N_2837,N_2073,N_2276);
nand U2838 (N_2838,N_2185,N_1854);
nand U2839 (N_2839,N_2106,N_2242);
nor U2840 (N_2840,N_2149,N_1871);
nand U2841 (N_2841,N_2038,N_1848);
or U2842 (N_2842,N_2220,N_2147);
and U2843 (N_2843,N_2022,N_2074);
nand U2844 (N_2844,N_2366,N_2283);
nand U2845 (N_2845,N_1880,N_2354);
and U2846 (N_2846,N_2135,N_1820);
or U2847 (N_2847,N_1980,N_2010);
or U2848 (N_2848,N_2345,N_1852);
or U2849 (N_2849,N_2298,N_2223);
or U2850 (N_2850,N_2252,N_2049);
nor U2851 (N_2851,N_1908,N_1853);
or U2852 (N_2852,N_2309,N_2056);
nor U2853 (N_2853,N_1843,N_2371);
nor U2854 (N_2854,N_2027,N_1934);
and U2855 (N_2855,N_2005,N_1839);
nor U2856 (N_2856,N_2364,N_1956);
nand U2857 (N_2857,N_1831,N_2254);
nand U2858 (N_2858,N_2319,N_1859);
nor U2859 (N_2859,N_2170,N_1913);
nor U2860 (N_2860,N_2039,N_2325);
xor U2861 (N_2861,N_2207,N_2057);
and U2862 (N_2862,N_1881,N_2368);
or U2863 (N_2863,N_2064,N_2392);
or U2864 (N_2864,N_2288,N_2246);
and U2865 (N_2865,N_1847,N_2377);
or U2866 (N_2866,N_1907,N_2344);
nor U2867 (N_2867,N_2139,N_1810);
or U2868 (N_2868,N_1951,N_1801);
and U2869 (N_2869,N_2203,N_2271);
or U2870 (N_2870,N_2144,N_2372);
nand U2871 (N_2871,N_2099,N_2171);
or U2872 (N_2872,N_2379,N_2184);
nor U2873 (N_2873,N_2003,N_1893);
xnor U2874 (N_2874,N_2364,N_2340);
xnor U2875 (N_2875,N_2308,N_2033);
or U2876 (N_2876,N_2226,N_2222);
and U2877 (N_2877,N_2180,N_2214);
nand U2878 (N_2878,N_2359,N_2216);
and U2879 (N_2879,N_2132,N_2097);
and U2880 (N_2880,N_1820,N_2271);
xnor U2881 (N_2881,N_2046,N_2249);
nand U2882 (N_2882,N_2236,N_1901);
nand U2883 (N_2883,N_2377,N_2392);
nor U2884 (N_2884,N_2059,N_2010);
nand U2885 (N_2885,N_2046,N_2199);
nor U2886 (N_2886,N_2128,N_2080);
nor U2887 (N_2887,N_1878,N_1952);
xor U2888 (N_2888,N_2060,N_2359);
nor U2889 (N_2889,N_2323,N_2229);
nand U2890 (N_2890,N_2372,N_1871);
nand U2891 (N_2891,N_1814,N_2216);
and U2892 (N_2892,N_2288,N_2321);
nand U2893 (N_2893,N_2351,N_2339);
nor U2894 (N_2894,N_1940,N_1948);
and U2895 (N_2895,N_2178,N_1944);
xnor U2896 (N_2896,N_2124,N_1856);
nand U2897 (N_2897,N_2068,N_1928);
and U2898 (N_2898,N_1849,N_2040);
and U2899 (N_2899,N_1917,N_2296);
and U2900 (N_2900,N_2214,N_2163);
nor U2901 (N_2901,N_2109,N_2339);
nor U2902 (N_2902,N_2338,N_2399);
and U2903 (N_2903,N_1929,N_2374);
xnor U2904 (N_2904,N_2247,N_2059);
and U2905 (N_2905,N_1964,N_2211);
or U2906 (N_2906,N_2256,N_1904);
nor U2907 (N_2907,N_2329,N_1843);
nand U2908 (N_2908,N_2393,N_2276);
or U2909 (N_2909,N_2388,N_1940);
nand U2910 (N_2910,N_2193,N_1979);
nor U2911 (N_2911,N_2350,N_2397);
and U2912 (N_2912,N_2058,N_2288);
xor U2913 (N_2913,N_2136,N_1821);
nor U2914 (N_2914,N_1920,N_2217);
or U2915 (N_2915,N_2391,N_2261);
nand U2916 (N_2916,N_2052,N_1871);
and U2917 (N_2917,N_2210,N_2038);
or U2918 (N_2918,N_2051,N_2277);
and U2919 (N_2919,N_2373,N_1971);
and U2920 (N_2920,N_2192,N_1845);
nand U2921 (N_2921,N_2332,N_2380);
or U2922 (N_2922,N_1828,N_1851);
or U2923 (N_2923,N_1908,N_2336);
or U2924 (N_2924,N_2274,N_2145);
nor U2925 (N_2925,N_2035,N_2350);
nor U2926 (N_2926,N_2051,N_1940);
nor U2927 (N_2927,N_2260,N_2357);
nand U2928 (N_2928,N_2284,N_2120);
nand U2929 (N_2929,N_2039,N_2117);
or U2930 (N_2930,N_2184,N_2306);
nor U2931 (N_2931,N_2248,N_1961);
or U2932 (N_2932,N_1943,N_2092);
or U2933 (N_2933,N_1987,N_2227);
and U2934 (N_2934,N_1830,N_2208);
nor U2935 (N_2935,N_2239,N_1851);
or U2936 (N_2936,N_2152,N_1811);
and U2937 (N_2937,N_2012,N_2387);
nand U2938 (N_2938,N_2042,N_1953);
or U2939 (N_2939,N_2012,N_1903);
nor U2940 (N_2940,N_2191,N_1969);
nand U2941 (N_2941,N_1933,N_2223);
nand U2942 (N_2942,N_2243,N_1888);
and U2943 (N_2943,N_2341,N_1968);
nand U2944 (N_2944,N_2391,N_2018);
nand U2945 (N_2945,N_2044,N_1909);
nand U2946 (N_2946,N_2068,N_2005);
nor U2947 (N_2947,N_2131,N_1951);
nor U2948 (N_2948,N_2330,N_2333);
or U2949 (N_2949,N_2023,N_1937);
nor U2950 (N_2950,N_1849,N_2127);
or U2951 (N_2951,N_1858,N_2390);
and U2952 (N_2952,N_2257,N_2334);
nand U2953 (N_2953,N_2022,N_2305);
nand U2954 (N_2954,N_2161,N_2110);
or U2955 (N_2955,N_2057,N_2155);
nor U2956 (N_2956,N_1917,N_1978);
and U2957 (N_2957,N_2055,N_2004);
nand U2958 (N_2958,N_1844,N_1894);
xnor U2959 (N_2959,N_2073,N_1947);
nand U2960 (N_2960,N_1869,N_1827);
and U2961 (N_2961,N_2238,N_1928);
nand U2962 (N_2962,N_1817,N_2230);
xor U2963 (N_2963,N_2183,N_1815);
and U2964 (N_2964,N_2030,N_2195);
and U2965 (N_2965,N_2364,N_1862);
or U2966 (N_2966,N_2107,N_2274);
and U2967 (N_2967,N_2223,N_2014);
and U2968 (N_2968,N_1980,N_2017);
nand U2969 (N_2969,N_1936,N_2304);
and U2970 (N_2970,N_2053,N_2347);
or U2971 (N_2971,N_1936,N_1844);
and U2972 (N_2972,N_2319,N_2006);
and U2973 (N_2973,N_1829,N_1864);
and U2974 (N_2974,N_1953,N_1857);
or U2975 (N_2975,N_2275,N_1966);
xnor U2976 (N_2976,N_1927,N_1900);
nor U2977 (N_2977,N_2093,N_2304);
xnor U2978 (N_2978,N_1907,N_2108);
and U2979 (N_2979,N_1989,N_1990);
nor U2980 (N_2980,N_2053,N_2144);
or U2981 (N_2981,N_1989,N_1854);
nand U2982 (N_2982,N_2313,N_2281);
nand U2983 (N_2983,N_2050,N_2209);
nand U2984 (N_2984,N_2114,N_1889);
nor U2985 (N_2985,N_2384,N_1978);
nor U2986 (N_2986,N_2392,N_1928);
and U2987 (N_2987,N_2397,N_2057);
nor U2988 (N_2988,N_2014,N_2001);
and U2989 (N_2989,N_2371,N_2031);
or U2990 (N_2990,N_1918,N_2333);
nor U2991 (N_2991,N_2081,N_2133);
nand U2992 (N_2992,N_1986,N_1940);
nor U2993 (N_2993,N_2318,N_2003);
xnor U2994 (N_2994,N_1899,N_2099);
and U2995 (N_2995,N_2338,N_1843);
or U2996 (N_2996,N_1940,N_2284);
and U2997 (N_2997,N_1840,N_2288);
or U2998 (N_2998,N_2297,N_2005);
nand U2999 (N_2999,N_1898,N_2210);
or UO_0 (O_0,N_2401,N_2599);
nand UO_1 (O_1,N_2406,N_2976);
and UO_2 (O_2,N_2596,N_2736);
nor UO_3 (O_3,N_2886,N_2862);
xnor UO_4 (O_4,N_2907,N_2423);
or UO_5 (O_5,N_2825,N_2992);
or UO_6 (O_6,N_2601,N_2660);
nor UO_7 (O_7,N_2796,N_2834);
and UO_8 (O_8,N_2570,N_2598);
or UO_9 (O_9,N_2893,N_2866);
nand UO_10 (O_10,N_2711,N_2823);
nand UO_11 (O_11,N_2538,N_2637);
or UO_12 (O_12,N_2575,N_2560);
nand UO_13 (O_13,N_2470,N_2433);
or UO_14 (O_14,N_2721,N_2475);
or UO_15 (O_15,N_2665,N_2629);
nor UO_16 (O_16,N_2627,N_2857);
or UO_17 (O_17,N_2841,N_2618);
nor UO_18 (O_18,N_2714,N_2718);
or UO_19 (O_19,N_2811,N_2690);
nand UO_20 (O_20,N_2858,N_2938);
nand UO_21 (O_21,N_2684,N_2940);
or UO_22 (O_22,N_2543,N_2682);
and UO_23 (O_23,N_2648,N_2790);
nor UO_24 (O_24,N_2557,N_2924);
nor UO_25 (O_25,N_2549,N_2454);
and UO_26 (O_26,N_2988,N_2849);
nor UO_27 (O_27,N_2888,N_2697);
and UO_28 (O_28,N_2656,N_2735);
or UO_29 (O_29,N_2683,N_2402);
nor UO_30 (O_30,N_2854,N_2771);
nand UO_31 (O_31,N_2593,N_2466);
nor UO_32 (O_32,N_2434,N_2542);
or UO_33 (O_33,N_2978,N_2931);
nor UO_34 (O_34,N_2800,N_2605);
nor UO_35 (O_35,N_2837,N_2567);
nor UO_36 (O_36,N_2960,N_2489);
and UO_37 (O_37,N_2701,N_2577);
nand UO_38 (O_38,N_2407,N_2864);
nor UO_39 (O_39,N_2508,N_2657);
xnor UO_40 (O_40,N_2578,N_2505);
nor UO_41 (O_41,N_2977,N_2915);
nor UO_42 (O_42,N_2498,N_2625);
or UO_43 (O_43,N_2524,N_2797);
nand UO_44 (O_44,N_2957,N_2713);
xor UO_45 (O_45,N_2677,N_2985);
and UO_46 (O_46,N_2614,N_2899);
xnor UO_47 (O_47,N_2617,N_2659);
and UO_48 (O_48,N_2744,N_2699);
xnor UO_49 (O_49,N_2843,N_2941);
nand UO_50 (O_50,N_2467,N_2485);
nand UO_51 (O_51,N_2817,N_2490);
nor UO_52 (O_52,N_2999,N_2424);
nand UO_53 (O_53,N_2952,N_2463);
or UO_54 (O_54,N_2753,N_2496);
or UO_55 (O_55,N_2820,N_2936);
or UO_56 (O_56,N_2780,N_2603);
or UO_57 (O_57,N_2891,N_2511);
nand UO_58 (O_58,N_2726,N_2668);
and UO_59 (O_59,N_2922,N_2669);
or UO_60 (O_60,N_2628,N_2422);
nand UO_61 (O_61,N_2623,N_2491);
nand UO_62 (O_62,N_2465,N_2851);
nor UO_63 (O_63,N_2492,N_2951);
nand UO_64 (O_64,N_2569,N_2692);
and UO_65 (O_65,N_2415,N_2550);
xor UO_66 (O_66,N_2788,N_2484);
nand UO_67 (O_67,N_2476,N_2822);
and UO_68 (O_68,N_2453,N_2462);
nor UO_69 (O_69,N_2408,N_2760);
or UO_70 (O_70,N_2742,N_2672);
or UO_71 (O_71,N_2876,N_2782);
or UO_72 (O_72,N_2717,N_2517);
and UO_73 (O_73,N_2725,N_2446);
or UO_74 (O_74,N_2739,N_2624);
xnor UO_75 (O_75,N_2981,N_2680);
and UO_76 (O_76,N_2416,N_2501);
or UO_77 (O_77,N_2932,N_2982);
and UO_78 (O_78,N_2762,N_2527);
nand UO_79 (O_79,N_2432,N_2715);
or UO_80 (O_80,N_2793,N_2970);
or UO_81 (O_81,N_2582,N_2808);
nand UO_82 (O_82,N_2873,N_2676);
and UO_83 (O_83,N_2486,N_2634);
or UO_84 (O_84,N_2927,N_2861);
nor UO_85 (O_85,N_2445,N_2691);
nor UO_86 (O_86,N_2644,N_2472);
or UO_87 (O_87,N_2609,N_2795);
nor UO_88 (O_88,N_2607,N_2908);
nor UO_89 (O_89,N_2968,N_2944);
and UO_90 (O_90,N_2564,N_2450);
xor UO_91 (O_91,N_2852,N_2794);
nor UO_92 (O_92,N_2548,N_2559);
or UO_93 (O_93,N_2473,N_2438);
nand UO_94 (O_94,N_2556,N_2917);
nand UO_95 (O_95,N_2612,N_2651);
and UO_96 (O_96,N_2881,N_2426);
and UO_97 (O_97,N_2905,N_2955);
or UO_98 (O_98,N_2942,N_2643);
nand UO_99 (O_99,N_2757,N_2555);
xor UO_100 (O_100,N_2980,N_2929);
nor UO_101 (O_101,N_2919,N_2580);
and UO_102 (O_102,N_2477,N_2497);
or UO_103 (O_103,N_2810,N_2914);
nand UO_104 (O_104,N_2845,N_2483);
or UO_105 (O_105,N_2500,N_2838);
or UO_106 (O_106,N_2877,N_2509);
nand UO_107 (O_107,N_2709,N_2778);
and UO_108 (O_108,N_2935,N_2719);
and UO_109 (O_109,N_2414,N_2452);
or UO_110 (O_110,N_2667,N_2602);
or UO_111 (O_111,N_2829,N_2541);
xnor UO_112 (O_112,N_2819,N_2534);
or UO_113 (O_113,N_2839,N_2769);
or UO_114 (O_114,N_2963,N_2703);
nand UO_115 (O_115,N_2996,N_2522);
or UO_116 (O_116,N_2840,N_2403);
and UO_117 (O_117,N_2400,N_2722);
or UO_118 (O_118,N_2633,N_2748);
or UO_119 (O_119,N_2673,N_2730);
and UO_120 (O_120,N_2558,N_2913);
and UO_121 (O_121,N_2895,N_2989);
or UO_122 (O_122,N_2975,N_2587);
and UO_123 (O_123,N_2640,N_2658);
nor UO_124 (O_124,N_2869,N_2745);
nand UO_125 (O_125,N_2740,N_2911);
nor UO_126 (O_126,N_2494,N_2595);
xnor UO_127 (O_127,N_2777,N_2551);
and UO_128 (O_128,N_2439,N_2576);
nand UO_129 (O_129,N_2809,N_2733);
or UO_130 (O_130,N_2768,N_2776);
or UO_131 (O_131,N_2724,N_2997);
xor UO_132 (O_132,N_2998,N_2889);
nand UO_133 (O_133,N_2850,N_2431);
nor UO_134 (O_134,N_2824,N_2689);
nor UO_135 (O_135,N_2826,N_2622);
and UO_136 (O_136,N_2664,N_2874);
or UO_137 (O_137,N_2912,N_2883);
nand UO_138 (O_138,N_2801,N_2920);
nor UO_139 (O_139,N_2743,N_2546);
and UO_140 (O_140,N_2784,N_2554);
nor UO_141 (O_141,N_2831,N_2562);
and UO_142 (O_142,N_2507,N_2661);
nor UO_143 (O_143,N_2758,N_2678);
or UO_144 (O_144,N_2458,N_2959);
nand UO_145 (O_145,N_2503,N_2860);
or UO_146 (O_146,N_2965,N_2815);
nor UO_147 (O_147,N_2571,N_2616);
and UO_148 (O_148,N_2934,N_2832);
nand UO_149 (O_149,N_2581,N_2608);
nand UO_150 (O_150,N_2774,N_2783);
nor UO_151 (O_151,N_2983,N_2887);
or UO_152 (O_152,N_2933,N_2592);
nor UO_153 (O_153,N_2412,N_2589);
or UO_154 (O_154,N_2687,N_2526);
nor UO_155 (O_155,N_2991,N_2420);
or UO_156 (O_156,N_2510,N_2513);
nand UO_157 (O_157,N_2947,N_2974);
and UO_158 (O_158,N_2767,N_2481);
nor UO_159 (O_159,N_2544,N_2856);
nor UO_160 (O_160,N_2499,N_2478);
xnor UO_161 (O_161,N_2844,N_2708);
and UO_162 (O_162,N_2532,N_2421);
nand UO_163 (O_163,N_2530,N_2611);
nor UO_164 (O_164,N_2720,N_2405);
or UO_165 (O_165,N_2537,N_2950);
and UO_166 (O_166,N_2652,N_2704);
or UO_167 (O_167,N_2946,N_2447);
nor UO_168 (O_168,N_2994,N_2653);
nand UO_169 (O_169,N_2504,N_2435);
or UO_170 (O_170,N_2961,N_2766);
nor UO_171 (O_171,N_2645,N_2518);
nor UO_172 (O_172,N_2727,N_2655);
or UO_173 (O_173,N_2828,N_2654);
nand UO_174 (O_174,N_2547,N_2419);
or UO_175 (O_175,N_2741,N_2943);
nand UO_176 (O_176,N_2460,N_2646);
or UO_177 (O_177,N_2441,N_2909);
nand UO_178 (O_178,N_2469,N_2910);
nor UO_179 (O_179,N_2506,N_2619);
or UO_180 (O_180,N_2479,N_2973);
xor UO_181 (O_181,N_2681,N_2679);
nor UO_182 (O_182,N_2563,N_2417);
or UO_183 (O_183,N_2901,N_2898);
nor UO_184 (O_184,N_2696,N_2896);
or UO_185 (O_185,N_2818,N_2647);
or UO_186 (O_186,N_2568,N_2761);
or UO_187 (O_187,N_2523,N_2902);
or UO_188 (O_188,N_2429,N_2807);
nor UO_189 (O_189,N_2954,N_2516);
or UO_190 (O_190,N_2512,N_2536);
and UO_191 (O_191,N_2613,N_2842);
xnor UO_192 (O_192,N_2533,N_2410);
nand UO_193 (O_193,N_2773,N_2700);
and UO_194 (O_194,N_2754,N_2586);
nor UO_195 (O_195,N_2666,N_2662);
nand UO_196 (O_196,N_2775,N_2882);
nor UO_197 (O_197,N_2585,N_2953);
nor UO_198 (O_198,N_2449,N_2867);
and UO_199 (O_199,N_2833,N_2962);
xor UO_200 (O_200,N_2791,N_2675);
or UO_201 (O_201,N_2650,N_2710);
nand UO_202 (O_202,N_2765,N_2620);
nor UO_203 (O_203,N_2847,N_2409);
nand UO_204 (O_204,N_2474,N_2671);
nand UO_205 (O_205,N_2900,N_2930);
nand UO_206 (O_206,N_2535,N_2734);
nor UO_207 (O_207,N_2885,N_2425);
or UO_208 (O_208,N_2565,N_2836);
nand UO_209 (O_209,N_2764,N_2418);
and UO_210 (O_210,N_2884,N_2604);
nor UO_211 (O_211,N_2615,N_2923);
and UO_212 (O_212,N_2816,N_2835);
nor UO_213 (O_213,N_2487,N_2814);
nor UO_214 (O_214,N_2798,N_2545);
nand UO_215 (O_215,N_2584,N_2488);
and UO_216 (O_216,N_2566,N_2440);
nor UO_217 (O_217,N_2482,N_2956);
or UO_218 (O_218,N_2493,N_2597);
nand UO_219 (O_219,N_2430,N_2695);
xnor UO_220 (O_220,N_2804,N_2972);
xor UO_221 (O_221,N_2827,N_2686);
xor UO_222 (O_222,N_2610,N_2728);
xnor UO_223 (O_223,N_2789,N_2442);
and UO_224 (O_224,N_2649,N_2949);
nand UO_225 (O_225,N_2868,N_2853);
and UO_226 (O_226,N_2456,N_2865);
and UO_227 (O_227,N_2529,N_2875);
nand UO_228 (O_228,N_2879,N_2631);
nand UO_229 (O_229,N_2404,N_2448);
nor UO_230 (O_230,N_2747,N_2706);
or UO_231 (O_231,N_2626,N_2755);
or UO_232 (O_232,N_2751,N_2903);
xor UO_233 (O_233,N_2759,N_2786);
and UO_234 (O_234,N_2471,N_2572);
or UO_235 (O_235,N_2579,N_2663);
nand UO_236 (O_236,N_2756,N_2806);
xor UO_237 (O_237,N_2750,N_2848);
or UO_238 (O_238,N_2594,N_2738);
nor UO_239 (O_239,N_2561,N_2880);
xnor UO_240 (O_240,N_2480,N_2606);
or UO_241 (O_241,N_2995,N_2525);
and UO_242 (O_242,N_2921,N_2641);
and UO_243 (O_243,N_2459,N_2772);
nand UO_244 (O_244,N_2846,N_2892);
xnor UO_245 (O_245,N_2515,N_2531);
nand UO_246 (O_246,N_2457,N_2732);
or UO_247 (O_247,N_2937,N_2785);
and UO_248 (O_248,N_2670,N_2763);
or UO_249 (O_249,N_2906,N_2871);
xnor UO_250 (O_250,N_2749,N_2698);
nand UO_251 (O_251,N_2813,N_2519);
or UO_252 (O_252,N_2642,N_2779);
xor UO_253 (O_253,N_2792,N_2945);
nor UO_254 (O_254,N_2712,N_2591);
and UO_255 (O_255,N_2705,N_2444);
nand UO_256 (O_256,N_2674,N_2693);
nand UO_257 (O_257,N_2918,N_2894);
and UO_258 (O_258,N_2729,N_2926);
or UO_259 (O_259,N_2639,N_2967);
nand UO_260 (O_260,N_2455,N_2993);
or UO_261 (O_261,N_2573,N_2702);
nand UO_262 (O_262,N_2521,N_2636);
or UO_263 (O_263,N_2990,N_2514);
or UO_264 (O_264,N_2413,N_2958);
nand UO_265 (O_265,N_2694,N_2539);
or UO_266 (O_266,N_2437,N_2855);
nand UO_267 (O_267,N_2781,N_2590);
and UO_268 (O_268,N_2979,N_2799);
nand UO_269 (O_269,N_2632,N_2969);
or UO_270 (O_270,N_2685,N_2803);
and UO_271 (O_271,N_2987,N_2746);
or UO_272 (O_272,N_2428,N_2731);
and UO_273 (O_273,N_2688,N_2986);
nor UO_274 (O_274,N_2872,N_2737);
xor UO_275 (O_275,N_2443,N_2984);
or UO_276 (O_276,N_2964,N_2635);
xnor UO_277 (O_277,N_2925,N_2904);
nand UO_278 (O_278,N_2502,N_2520);
xnor UO_279 (O_279,N_2630,N_2821);
or UO_280 (O_280,N_2805,N_2723);
and UO_281 (O_281,N_2752,N_2890);
nor UO_282 (O_282,N_2812,N_2948);
and UO_283 (O_283,N_2528,N_2583);
and UO_284 (O_284,N_2830,N_2787);
nor UO_285 (O_285,N_2588,N_2707);
or UO_286 (O_286,N_2928,N_2574);
and UO_287 (O_287,N_2552,N_2770);
and UO_288 (O_288,N_2600,N_2971);
and UO_289 (O_289,N_2863,N_2553);
nor UO_290 (O_290,N_2966,N_2461);
nor UO_291 (O_291,N_2427,N_2916);
nand UO_292 (O_292,N_2411,N_2878);
nor UO_293 (O_293,N_2939,N_2464);
nand UO_294 (O_294,N_2468,N_2451);
and UO_295 (O_295,N_2621,N_2870);
nor UO_296 (O_296,N_2859,N_2540);
or UO_297 (O_297,N_2716,N_2495);
and UO_298 (O_298,N_2638,N_2436);
and UO_299 (O_299,N_2802,N_2897);
nor UO_300 (O_300,N_2700,N_2937);
or UO_301 (O_301,N_2625,N_2945);
and UO_302 (O_302,N_2753,N_2608);
nand UO_303 (O_303,N_2762,N_2565);
nor UO_304 (O_304,N_2779,N_2580);
and UO_305 (O_305,N_2704,N_2628);
or UO_306 (O_306,N_2607,N_2602);
nand UO_307 (O_307,N_2767,N_2821);
or UO_308 (O_308,N_2941,N_2678);
nand UO_309 (O_309,N_2739,N_2913);
nor UO_310 (O_310,N_2879,N_2706);
nor UO_311 (O_311,N_2669,N_2451);
and UO_312 (O_312,N_2726,N_2546);
nor UO_313 (O_313,N_2404,N_2669);
or UO_314 (O_314,N_2644,N_2594);
nor UO_315 (O_315,N_2789,N_2485);
nand UO_316 (O_316,N_2415,N_2695);
or UO_317 (O_317,N_2641,N_2816);
or UO_318 (O_318,N_2544,N_2812);
or UO_319 (O_319,N_2948,N_2843);
nand UO_320 (O_320,N_2941,N_2793);
nor UO_321 (O_321,N_2999,N_2627);
or UO_322 (O_322,N_2848,N_2825);
nor UO_323 (O_323,N_2527,N_2934);
nor UO_324 (O_324,N_2934,N_2473);
nand UO_325 (O_325,N_2430,N_2936);
and UO_326 (O_326,N_2700,N_2466);
and UO_327 (O_327,N_2942,N_2879);
nand UO_328 (O_328,N_2491,N_2588);
nand UO_329 (O_329,N_2757,N_2762);
nand UO_330 (O_330,N_2542,N_2617);
nand UO_331 (O_331,N_2420,N_2496);
nand UO_332 (O_332,N_2843,N_2662);
nand UO_333 (O_333,N_2826,N_2959);
and UO_334 (O_334,N_2962,N_2587);
or UO_335 (O_335,N_2414,N_2883);
nor UO_336 (O_336,N_2872,N_2458);
and UO_337 (O_337,N_2948,N_2680);
nor UO_338 (O_338,N_2413,N_2646);
or UO_339 (O_339,N_2827,N_2573);
and UO_340 (O_340,N_2767,N_2783);
nand UO_341 (O_341,N_2523,N_2819);
xor UO_342 (O_342,N_2794,N_2486);
nor UO_343 (O_343,N_2647,N_2511);
nand UO_344 (O_344,N_2740,N_2629);
or UO_345 (O_345,N_2994,N_2811);
nand UO_346 (O_346,N_2620,N_2723);
or UO_347 (O_347,N_2430,N_2424);
nand UO_348 (O_348,N_2595,N_2464);
and UO_349 (O_349,N_2467,N_2591);
and UO_350 (O_350,N_2599,N_2418);
nand UO_351 (O_351,N_2836,N_2955);
or UO_352 (O_352,N_2678,N_2656);
or UO_353 (O_353,N_2983,N_2993);
or UO_354 (O_354,N_2452,N_2489);
nor UO_355 (O_355,N_2947,N_2486);
or UO_356 (O_356,N_2743,N_2822);
or UO_357 (O_357,N_2881,N_2938);
nand UO_358 (O_358,N_2903,N_2660);
or UO_359 (O_359,N_2417,N_2982);
nor UO_360 (O_360,N_2603,N_2799);
or UO_361 (O_361,N_2732,N_2631);
nand UO_362 (O_362,N_2583,N_2885);
and UO_363 (O_363,N_2652,N_2726);
nand UO_364 (O_364,N_2692,N_2656);
and UO_365 (O_365,N_2642,N_2433);
or UO_366 (O_366,N_2640,N_2665);
and UO_367 (O_367,N_2574,N_2843);
and UO_368 (O_368,N_2897,N_2972);
nand UO_369 (O_369,N_2999,N_2630);
nand UO_370 (O_370,N_2591,N_2578);
and UO_371 (O_371,N_2934,N_2946);
and UO_372 (O_372,N_2626,N_2806);
or UO_373 (O_373,N_2962,N_2746);
nor UO_374 (O_374,N_2851,N_2652);
or UO_375 (O_375,N_2408,N_2639);
and UO_376 (O_376,N_2419,N_2527);
or UO_377 (O_377,N_2413,N_2545);
or UO_378 (O_378,N_2711,N_2857);
nand UO_379 (O_379,N_2799,N_2558);
and UO_380 (O_380,N_2419,N_2890);
nand UO_381 (O_381,N_2477,N_2570);
xnor UO_382 (O_382,N_2474,N_2967);
nand UO_383 (O_383,N_2430,N_2917);
and UO_384 (O_384,N_2988,N_2513);
or UO_385 (O_385,N_2824,N_2549);
nand UO_386 (O_386,N_2750,N_2832);
or UO_387 (O_387,N_2612,N_2483);
nand UO_388 (O_388,N_2642,N_2660);
nand UO_389 (O_389,N_2934,N_2674);
or UO_390 (O_390,N_2412,N_2863);
nand UO_391 (O_391,N_2505,N_2426);
nand UO_392 (O_392,N_2599,N_2798);
and UO_393 (O_393,N_2567,N_2984);
or UO_394 (O_394,N_2507,N_2490);
xnor UO_395 (O_395,N_2697,N_2934);
and UO_396 (O_396,N_2422,N_2955);
nor UO_397 (O_397,N_2973,N_2456);
and UO_398 (O_398,N_2944,N_2532);
xnor UO_399 (O_399,N_2799,N_2601);
or UO_400 (O_400,N_2407,N_2610);
xor UO_401 (O_401,N_2672,N_2694);
and UO_402 (O_402,N_2604,N_2636);
or UO_403 (O_403,N_2659,N_2652);
and UO_404 (O_404,N_2471,N_2850);
nor UO_405 (O_405,N_2683,N_2772);
or UO_406 (O_406,N_2495,N_2836);
nand UO_407 (O_407,N_2659,N_2685);
and UO_408 (O_408,N_2953,N_2490);
nor UO_409 (O_409,N_2515,N_2625);
or UO_410 (O_410,N_2427,N_2437);
nand UO_411 (O_411,N_2434,N_2581);
nand UO_412 (O_412,N_2655,N_2431);
nor UO_413 (O_413,N_2962,N_2597);
nand UO_414 (O_414,N_2771,N_2710);
and UO_415 (O_415,N_2952,N_2456);
or UO_416 (O_416,N_2686,N_2646);
or UO_417 (O_417,N_2736,N_2841);
xnor UO_418 (O_418,N_2817,N_2442);
nand UO_419 (O_419,N_2542,N_2607);
and UO_420 (O_420,N_2552,N_2951);
or UO_421 (O_421,N_2604,N_2852);
nor UO_422 (O_422,N_2784,N_2401);
or UO_423 (O_423,N_2800,N_2827);
and UO_424 (O_424,N_2419,N_2647);
nand UO_425 (O_425,N_2780,N_2629);
and UO_426 (O_426,N_2942,N_2834);
nand UO_427 (O_427,N_2859,N_2518);
nand UO_428 (O_428,N_2608,N_2476);
and UO_429 (O_429,N_2420,N_2592);
nor UO_430 (O_430,N_2568,N_2540);
nor UO_431 (O_431,N_2577,N_2571);
xor UO_432 (O_432,N_2413,N_2961);
nor UO_433 (O_433,N_2962,N_2464);
nor UO_434 (O_434,N_2635,N_2467);
nor UO_435 (O_435,N_2551,N_2617);
or UO_436 (O_436,N_2756,N_2644);
and UO_437 (O_437,N_2519,N_2794);
or UO_438 (O_438,N_2689,N_2792);
nor UO_439 (O_439,N_2423,N_2631);
and UO_440 (O_440,N_2700,N_2682);
or UO_441 (O_441,N_2855,N_2635);
xnor UO_442 (O_442,N_2428,N_2801);
and UO_443 (O_443,N_2521,N_2473);
nor UO_444 (O_444,N_2444,N_2841);
and UO_445 (O_445,N_2488,N_2917);
and UO_446 (O_446,N_2723,N_2755);
or UO_447 (O_447,N_2425,N_2454);
xnor UO_448 (O_448,N_2709,N_2918);
xor UO_449 (O_449,N_2840,N_2982);
xnor UO_450 (O_450,N_2553,N_2745);
xor UO_451 (O_451,N_2547,N_2641);
and UO_452 (O_452,N_2795,N_2723);
nor UO_453 (O_453,N_2586,N_2950);
or UO_454 (O_454,N_2515,N_2698);
xor UO_455 (O_455,N_2487,N_2526);
or UO_456 (O_456,N_2702,N_2706);
nand UO_457 (O_457,N_2668,N_2961);
nor UO_458 (O_458,N_2734,N_2755);
xor UO_459 (O_459,N_2741,N_2624);
and UO_460 (O_460,N_2477,N_2981);
nand UO_461 (O_461,N_2519,N_2689);
or UO_462 (O_462,N_2589,N_2860);
or UO_463 (O_463,N_2462,N_2936);
nor UO_464 (O_464,N_2532,N_2524);
nor UO_465 (O_465,N_2528,N_2428);
nand UO_466 (O_466,N_2609,N_2874);
or UO_467 (O_467,N_2419,N_2950);
nand UO_468 (O_468,N_2830,N_2797);
and UO_469 (O_469,N_2645,N_2755);
nor UO_470 (O_470,N_2688,N_2450);
or UO_471 (O_471,N_2706,N_2699);
or UO_472 (O_472,N_2685,N_2518);
or UO_473 (O_473,N_2423,N_2411);
and UO_474 (O_474,N_2810,N_2882);
or UO_475 (O_475,N_2716,N_2570);
nor UO_476 (O_476,N_2787,N_2789);
xnor UO_477 (O_477,N_2855,N_2462);
and UO_478 (O_478,N_2790,N_2777);
xnor UO_479 (O_479,N_2878,N_2780);
nand UO_480 (O_480,N_2852,N_2456);
and UO_481 (O_481,N_2932,N_2479);
and UO_482 (O_482,N_2580,N_2648);
xnor UO_483 (O_483,N_2422,N_2977);
nor UO_484 (O_484,N_2818,N_2820);
or UO_485 (O_485,N_2954,N_2490);
or UO_486 (O_486,N_2451,N_2701);
nand UO_487 (O_487,N_2744,N_2585);
and UO_488 (O_488,N_2734,N_2775);
nand UO_489 (O_489,N_2793,N_2920);
nor UO_490 (O_490,N_2686,N_2622);
xor UO_491 (O_491,N_2973,N_2962);
nand UO_492 (O_492,N_2431,N_2570);
nor UO_493 (O_493,N_2669,N_2499);
nor UO_494 (O_494,N_2792,N_2464);
nor UO_495 (O_495,N_2762,N_2621);
nand UO_496 (O_496,N_2989,N_2607);
and UO_497 (O_497,N_2597,N_2596);
xnor UO_498 (O_498,N_2719,N_2894);
or UO_499 (O_499,N_2883,N_2685);
endmodule