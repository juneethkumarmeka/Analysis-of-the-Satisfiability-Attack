module basic_750_5000_1000_10_levels_10xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
nand U0 (N_0,In_408,In_423);
xor U1 (N_1,In_726,In_529);
nor U2 (N_2,In_561,In_500);
or U3 (N_3,In_679,In_442);
nand U4 (N_4,In_344,In_448);
and U5 (N_5,In_247,In_656);
nand U6 (N_6,In_40,In_749);
nor U7 (N_7,In_601,In_8);
nor U8 (N_8,In_721,In_740);
or U9 (N_9,In_392,In_107);
and U10 (N_10,In_20,In_515);
xnor U11 (N_11,In_146,In_616);
and U12 (N_12,In_108,In_145);
or U13 (N_13,In_307,In_670);
xor U14 (N_14,In_263,In_715);
nor U15 (N_15,In_122,In_433);
nor U16 (N_16,In_245,In_175);
nor U17 (N_17,In_511,In_608);
or U18 (N_18,In_243,In_476);
nor U19 (N_19,In_171,In_128);
xnor U20 (N_20,In_673,In_468);
nor U21 (N_21,In_270,In_135);
xnor U22 (N_22,In_334,In_86);
nand U23 (N_23,In_99,In_388);
nand U24 (N_24,In_420,In_300);
nand U25 (N_25,In_507,In_514);
xor U26 (N_26,In_488,In_183);
and U27 (N_27,In_505,In_301);
nand U28 (N_28,In_267,In_340);
and U29 (N_29,In_692,In_662);
or U30 (N_30,In_131,In_729);
nor U31 (N_31,In_123,In_155);
nand U32 (N_32,In_125,In_304);
nor U33 (N_33,In_173,In_78);
and U34 (N_34,In_238,In_547);
nor U35 (N_35,In_521,In_264);
nor U36 (N_36,In_716,In_34);
nor U37 (N_37,In_646,In_533);
xnor U38 (N_38,In_432,In_397);
nand U39 (N_39,In_704,In_479);
or U40 (N_40,In_728,In_580);
nand U41 (N_41,In_203,In_280);
or U42 (N_42,In_115,In_421);
nor U43 (N_43,In_193,In_395);
xnor U44 (N_44,In_284,In_396);
or U45 (N_45,In_355,In_711);
nor U46 (N_46,In_456,In_528);
and U47 (N_47,In_356,In_551);
nor U48 (N_48,In_502,In_672);
nor U49 (N_49,In_731,In_589);
and U50 (N_50,In_346,In_309);
or U51 (N_51,In_303,In_718);
nand U52 (N_52,In_540,In_567);
or U53 (N_53,In_15,In_215);
and U54 (N_54,In_75,In_541);
nand U55 (N_55,In_28,In_165);
xnor U56 (N_56,In_478,In_332);
or U57 (N_57,In_473,In_480);
xor U58 (N_58,In_363,In_273);
and U59 (N_59,In_229,In_156);
nand U60 (N_60,In_235,In_415);
and U61 (N_61,In_322,In_172);
xor U62 (N_62,In_216,In_629);
nor U63 (N_63,In_26,In_170);
and U64 (N_64,In_268,In_538);
nand U65 (N_65,In_292,In_253);
nor U66 (N_66,In_546,In_79);
or U67 (N_67,In_720,In_22);
nand U68 (N_68,In_364,In_96);
nor U69 (N_69,In_369,In_321);
and U70 (N_70,In_584,In_689);
and U71 (N_71,In_407,In_298);
xnor U72 (N_72,In_744,In_236);
xnor U73 (N_73,In_633,In_38);
xor U74 (N_74,In_299,In_76);
or U75 (N_75,In_176,In_709);
or U76 (N_76,In_545,In_517);
nand U77 (N_77,In_95,In_565);
and U78 (N_78,In_427,In_699);
nand U79 (N_79,In_470,In_387);
xor U80 (N_80,In_100,In_635);
xor U81 (N_81,In_204,In_587);
nand U82 (N_82,In_296,In_308);
nor U83 (N_83,In_80,In_652);
and U84 (N_84,In_83,In_378);
xnor U85 (N_85,In_668,In_320);
nor U86 (N_86,In_487,In_101);
xor U87 (N_87,In_437,In_714);
xor U88 (N_88,In_39,In_526);
nand U89 (N_89,In_249,In_47);
xnor U90 (N_90,In_82,In_534);
xnor U91 (N_91,In_458,In_119);
or U92 (N_92,In_312,In_191);
nor U93 (N_93,In_518,In_581);
nor U94 (N_94,In_681,In_106);
nor U95 (N_95,In_375,In_530);
nand U96 (N_96,In_196,In_252);
xnor U97 (N_97,In_461,In_688);
or U98 (N_98,In_341,In_390);
nor U99 (N_99,In_742,In_178);
nor U100 (N_100,In_683,In_462);
xnor U101 (N_101,In_293,In_331);
xnor U102 (N_102,In_443,In_35);
nor U103 (N_103,In_638,In_140);
and U104 (N_104,In_221,In_294);
nor U105 (N_105,In_282,In_66);
nand U106 (N_106,In_531,In_464);
xnor U107 (N_107,In_117,In_207);
or U108 (N_108,In_289,In_536);
nor U109 (N_109,In_241,In_647);
nand U110 (N_110,In_37,In_359);
xor U111 (N_111,In_642,In_677);
nand U112 (N_112,In_436,In_724);
xor U113 (N_113,In_674,In_149);
or U114 (N_114,In_212,In_2);
and U115 (N_115,In_305,In_297);
or U116 (N_116,In_326,In_648);
nor U117 (N_117,In_351,In_329);
and U118 (N_118,In_316,In_110);
xor U119 (N_119,In_445,In_112);
and U120 (N_120,In_434,In_10);
nand U121 (N_121,In_475,In_85);
xor U122 (N_122,In_560,In_625);
or U123 (N_123,In_315,In_105);
or U124 (N_124,In_276,In_350);
xor U125 (N_125,In_65,In_46);
nor U126 (N_126,In_266,In_136);
and U127 (N_127,In_684,In_357);
nand U128 (N_128,In_61,In_671);
xor U129 (N_129,In_365,In_482);
nor U130 (N_130,In_653,In_572);
xnor U131 (N_131,In_596,In_348);
and U132 (N_132,In_13,In_497);
nand U133 (N_133,In_93,In_201);
nand U134 (N_134,In_57,In_570);
nor U135 (N_135,In_218,In_412);
nor U136 (N_136,In_248,In_272);
xnor U137 (N_137,In_746,In_472);
xor U138 (N_138,In_250,In_559);
or U139 (N_139,In_738,In_379);
and U140 (N_140,In_523,In_457);
nor U141 (N_141,In_60,In_55);
xnor U142 (N_142,In_535,In_664);
or U143 (N_143,In_91,In_217);
nand U144 (N_144,In_634,In_202);
nand U145 (N_145,In_354,In_383);
nor U146 (N_146,In_532,In_694);
or U147 (N_147,In_513,In_114);
nand U148 (N_148,In_69,In_134);
nand U149 (N_149,In_640,In_499);
or U150 (N_150,In_695,In_59);
xor U151 (N_151,In_180,In_706);
and U152 (N_152,In_366,In_444);
nand U153 (N_153,In_143,In_385);
xnor U154 (N_154,In_230,In_328);
nand U155 (N_155,In_199,In_277);
and U156 (N_156,In_418,In_295);
nand U157 (N_157,In_279,In_370);
nand U158 (N_158,In_748,In_324);
nand U159 (N_159,In_111,In_51);
xnor U160 (N_160,In_113,In_214);
xnor U161 (N_161,In_409,In_345);
nand U162 (N_162,In_747,In_104);
or U163 (N_163,In_474,In_419);
or U164 (N_164,In_678,In_519);
nor U165 (N_165,In_211,In_636);
nor U166 (N_166,In_225,In_283);
nand U167 (N_167,In_522,In_158);
xnor U168 (N_168,In_624,In_441);
nand U169 (N_169,In_281,In_555);
or U170 (N_170,In_0,In_439);
nor U171 (N_171,In_362,In_144);
or U172 (N_172,In_43,In_594);
and U173 (N_173,In_597,In_542);
xnor U174 (N_174,In_730,In_219);
and U175 (N_175,In_380,In_353);
or U176 (N_176,In_583,In_325);
nor U177 (N_177,In_360,In_228);
or U178 (N_178,In_440,In_454);
xor U179 (N_179,In_210,In_72);
or U180 (N_180,In_349,In_36);
nor U181 (N_181,In_5,In_130);
xnor U182 (N_182,In_84,In_705);
nor U183 (N_183,In_242,In_571);
nand U184 (N_184,In_722,In_81);
or U185 (N_185,In_147,In_639);
and U186 (N_186,In_246,In_148);
and U187 (N_187,In_550,In_620);
or U188 (N_188,In_285,In_516);
nor U189 (N_189,In_31,In_422);
or U190 (N_190,In_399,In_707);
nor U191 (N_191,In_150,In_451);
nand U192 (N_192,In_339,In_413);
nor U193 (N_193,In_233,In_598);
or U194 (N_194,In_77,In_102);
xnor U195 (N_195,In_259,In_727);
or U196 (N_196,In_599,In_736);
nor U197 (N_197,In_493,In_1);
or U198 (N_198,In_665,In_605);
nand U199 (N_199,In_645,In_743);
xor U200 (N_200,In_557,In_382);
nor U201 (N_201,In_563,In_401);
or U202 (N_202,In_12,In_501);
or U203 (N_203,In_368,In_74);
nor U204 (N_204,In_361,In_492);
nor U205 (N_205,In_261,In_595);
or U206 (N_206,In_719,In_381);
nand U207 (N_207,In_209,In_92);
nand U208 (N_208,In_256,In_447);
xnor U209 (N_209,In_391,In_179);
nor U210 (N_210,In_693,In_735);
nand U211 (N_211,In_509,In_188);
or U212 (N_212,In_628,In_438);
and U213 (N_213,In_591,In_450);
or U214 (N_214,In_67,In_386);
nor U215 (N_215,In_459,In_260);
and U216 (N_216,In_568,In_71);
nor U217 (N_217,In_659,In_287);
and U218 (N_218,In_161,In_64);
and U219 (N_219,In_154,In_405);
or U220 (N_220,In_137,In_600);
and U221 (N_221,In_734,In_231);
xor U222 (N_222,In_612,In_213);
and U223 (N_223,In_335,In_9);
xnor U224 (N_224,In_337,In_142);
nor U225 (N_225,In_342,In_373);
xnor U226 (N_226,In_330,In_520);
nand U227 (N_227,In_489,In_288);
nand U228 (N_228,In_63,In_495);
xnor U229 (N_229,In_42,In_573);
nor U230 (N_230,In_30,In_6);
and U231 (N_231,In_669,In_611);
nand U232 (N_232,In_604,In_377);
or U233 (N_233,In_262,In_187);
nor U234 (N_234,In_741,In_661);
xor U235 (N_235,In_314,In_127);
and U236 (N_236,In_192,In_269);
nand U237 (N_237,In_562,In_244);
xnor U238 (N_238,In_319,In_622);
and U239 (N_239,In_52,In_524);
nor U240 (N_240,In_506,In_197);
and U241 (N_241,In_343,In_313);
nor U242 (N_242,In_49,In_306);
nand U243 (N_243,In_675,In_712);
xor U244 (N_244,In_537,In_333);
nor U245 (N_245,In_358,In_132);
or U246 (N_246,In_603,In_525);
nand U247 (N_247,In_11,In_318);
or U248 (N_248,In_124,In_402);
nand U249 (N_249,In_737,In_632);
xnor U250 (N_250,In_686,In_310);
and U251 (N_251,In_157,In_393);
nor U252 (N_252,In_163,In_558);
nor U253 (N_253,In_696,In_637);
and U254 (N_254,In_70,In_129);
nand U255 (N_255,In_103,In_29);
nand U256 (N_256,In_655,In_94);
nor U257 (N_257,In_713,In_471);
or U258 (N_258,In_374,In_549);
nor U259 (N_259,In_732,In_650);
nor U260 (N_260,In_160,In_430);
xor U261 (N_261,In_208,In_574);
and U262 (N_262,In_685,In_17);
nor U263 (N_263,In_630,In_676);
nor U264 (N_264,In_543,In_739);
nor U265 (N_265,In_254,In_278);
or U266 (N_266,In_658,In_651);
and U267 (N_267,In_631,In_190);
nor U268 (N_268,In_575,In_702);
or U269 (N_269,In_429,In_317);
xor U270 (N_270,In_186,In_623);
nor U271 (N_271,In_607,In_496);
nor U272 (N_272,In_126,In_16);
and U273 (N_273,In_234,In_494);
or U274 (N_274,In_613,In_490);
nor U275 (N_275,In_617,In_311);
and U276 (N_276,In_657,In_552);
nand U277 (N_277,In_224,In_428);
nor U278 (N_278,In_152,In_690);
or U279 (N_279,In_586,In_181);
or U280 (N_280,In_120,In_486);
nand U281 (N_281,In_166,In_411);
or U282 (N_282,In_621,In_404);
xnor U283 (N_283,In_45,In_138);
nand U284 (N_284,In_226,In_578);
or U285 (N_285,In_703,In_141);
nor U286 (N_286,In_153,In_302);
xor U287 (N_287,In_484,In_227);
nor U288 (N_288,In_723,In_687);
or U289 (N_289,In_697,In_431);
nor U290 (N_290,In_660,In_21);
xnor U291 (N_291,In_453,In_467);
or U292 (N_292,In_376,In_347);
nor U293 (N_293,In_426,In_90);
xnor U294 (N_294,In_7,In_44);
nor U295 (N_295,In_465,In_371);
or U296 (N_296,In_336,In_643);
and U297 (N_297,In_372,In_185);
and U298 (N_298,In_483,In_508);
nor U299 (N_299,In_58,In_3);
nand U300 (N_300,In_414,In_592);
xnor U301 (N_301,In_491,In_286);
nand U302 (N_302,In_290,In_352);
or U303 (N_303,In_485,In_708);
nand U304 (N_304,In_539,In_733);
xnor U305 (N_305,In_425,In_403);
or U306 (N_306,In_159,In_498);
and U307 (N_307,In_162,In_663);
xnor U308 (N_308,In_416,In_327);
nand U309 (N_309,In_118,In_466);
xnor U310 (N_310,In_554,In_452);
or U311 (N_311,In_88,In_579);
xor U312 (N_312,In_548,In_576);
nor U313 (N_313,In_133,In_627);
nand U314 (N_314,In_590,In_577);
and U315 (N_315,In_54,In_121);
or U316 (N_316,In_569,In_460);
and U317 (N_317,In_184,In_24);
xor U318 (N_318,In_553,In_644);
or U319 (N_319,In_14,In_109);
xor U320 (N_320,In_73,In_198);
nand U321 (N_321,In_504,In_626);
xor U322 (N_322,In_18,In_503);
and U323 (N_323,In_691,In_206);
or U324 (N_324,In_164,In_641);
and U325 (N_325,In_588,In_338);
and U326 (N_326,In_700,In_602);
and U327 (N_327,In_53,In_222);
xnor U328 (N_328,In_556,In_609);
xnor U329 (N_329,In_139,In_182);
nor U330 (N_330,In_367,In_510);
nor U331 (N_331,In_582,In_400);
or U332 (N_332,In_610,In_606);
xnor U333 (N_333,In_151,In_389);
or U334 (N_334,In_512,In_27);
and U335 (N_335,In_255,In_56);
nor U336 (N_336,In_544,In_654);
or U337 (N_337,In_48,In_62);
nand U338 (N_338,In_614,In_619);
and U339 (N_339,In_237,In_98);
and U340 (N_340,In_469,In_50);
nand U341 (N_341,In_449,In_195);
and U342 (N_342,In_265,In_32);
nor U343 (N_343,In_223,In_168);
or U344 (N_344,In_116,In_701);
nand U345 (N_345,In_698,In_417);
nand U346 (N_346,In_25,In_717);
nor U347 (N_347,In_240,In_323);
nand U348 (N_348,In_258,In_205);
or U349 (N_349,In_682,In_232);
xnor U350 (N_350,In_194,In_384);
or U351 (N_351,In_566,In_167);
and U352 (N_352,In_23,In_477);
nand U353 (N_353,In_406,In_463);
nor U354 (N_354,In_33,In_618);
or U355 (N_355,In_585,In_275);
xor U356 (N_356,In_41,In_169);
nor U357 (N_357,In_271,In_725);
and U358 (N_358,In_177,In_87);
nor U359 (N_359,In_680,In_615);
nor U360 (N_360,In_446,In_189);
or U361 (N_361,In_291,In_410);
and U362 (N_362,In_220,In_593);
xor U363 (N_363,In_251,In_481);
xnor U364 (N_364,In_174,In_398);
xnor U365 (N_365,In_667,In_200);
nand U366 (N_366,In_666,In_394);
xnor U367 (N_367,In_455,In_4);
and U368 (N_368,In_239,In_564);
xnor U369 (N_369,In_527,In_274);
or U370 (N_370,In_710,In_745);
nor U371 (N_371,In_257,In_649);
nand U372 (N_372,In_19,In_424);
xor U373 (N_373,In_68,In_97);
nand U374 (N_374,In_89,In_435);
xor U375 (N_375,In_68,In_220);
and U376 (N_376,In_628,In_549);
and U377 (N_377,In_713,In_269);
and U378 (N_378,In_78,In_744);
xnor U379 (N_379,In_446,In_416);
or U380 (N_380,In_691,In_392);
xnor U381 (N_381,In_501,In_411);
nand U382 (N_382,In_166,In_187);
nand U383 (N_383,In_28,In_185);
or U384 (N_384,In_356,In_170);
xnor U385 (N_385,In_544,In_45);
nand U386 (N_386,In_645,In_152);
nor U387 (N_387,In_676,In_729);
and U388 (N_388,In_203,In_714);
nand U389 (N_389,In_57,In_447);
nand U390 (N_390,In_709,In_562);
xor U391 (N_391,In_235,In_370);
nand U392 (N_392,In_44,In_484);
and U393 (N_393,In_598,In_354);
nor U394 (N_394,In_284,In_90);
nor U395 (N_395,In_155,In_234);
and U396 (N_396,In_344,In_94);
nand U397 (N_397,In_123,In_551);
nor U398 (N_398,In_340,In_452);
nor U399 (N_399,In_601,In_547);
nand U400 (N_400,In_131,In_128);
nand U401 (N_401,In_335,In_309);
or U402 (N_402,In_77,In_544);
nor U403 (N_403,In_123,In_682);
xor U404 (N_404,In_250,In_737);
nor U405 (N_405,In_456,In_92);
or U406 (N_406,In_260,In_408);
xor U407 (N_407,In_353,In_437);
and U408 (N_408,In_524,In_358);
nand U409 (N_409,In_124,In_663);
xnor U410 (N_410,In_336,In_394);
xnor U411 (N_411,In_686,In_347);
nand U412 (N_412,In_595,In_459);
nand U413 (N_413,In_339,In_213);
nor U414 (N_414,In_670,In_190);
nand U415 (N_415,In_152,In_587);
and U416 (N_416,In_589,In_329);
and U417 (N_417,In_239,In_289);
and U418 (N_418,In_427,In_310);
nand U419 (N_419,In_362,In_40);
nand U420 (N_420,In_731,In_11);
xor U421 (N_421,In_385,In_106);
or U422 (N_422,In_100,In_685);
or U423 (N_423,In_209,In_93);
nand U424 (N_424,In_459,In_32);
or U425 (N_425,In_663,In_578);
and U426 (N_426,In_72,In_273);
xor U427 (N_427,In_80,In_320);
xnor U428 (N_428,In_495,In_15);
nor U429 (N_429,In_310,In_581);
nand U430 (N_430,In_563,In_543);
xor U431 (N_431,In_561,In_679);
and U432 (N_432,In_385,In_269);
and U433 (N_433,In_547,In_650);
and U434 (N_434,In_334,In_149);
nand U435 (N_435,In_21,In_690);
or U436 (N_436,In_51,In_245);
or U437 (N_437,In_303,In_613);
or U438 (N_438,In_736,In_253);
or U439 (N_439,In_501,In_729);
nand U440 (N_440,In_350,In_325);
nor U441 (N_441,In_299,In_186);
nor U442 (N_442,In_557,In_216);
or U443 (N_443,In_409,In_741);
and U444 (N_444,In_539,In_148);
nor U445 (N_445,In_412,In_500);
nor U446 (N_446,In_0,In_592);
xor U447 (N_447,In_311,In_265);
and U448 (N_448,In_147,In_43);
xor U449 (N_449,In_122,In_644);
and U450 (N_450,In_375,In_607);
and U451 (N_451,In_192,In_216);
and U452 (N_452,In_665,In_708);
or U453 (N_453,In_681,In_747);
xnor U454 (N_454,In_165,In_423);
xnor U455 (N_455,In_400,In_61);
and U456 (N_456,In_570,In_279);
and U457 (N_457,In_168,In_314);
or U458 (N_458,In_201,In_297);
xor U459 (N_459,In_744,In_459);
nor U460 (N_460,In_484,In_205);
xor U461 (N_461,In_705,In_109);
nor U462 (N_462,In_641,In_500);
nor U463 (N_463,In_54,In_531);
and U464 (N_464,In_63,In_631);
nand U465 (N_465,In_6,In_742);
or U466 (N_466,In_631,In_349);
and U467 (N_467,In_641,In_544);
nor U468 (N_468,In_696,In_484);
and U469 (N_469,In_337,In_71);
xor U470 (N_470,In_231,In_104);
or U471 (N_471,In_71,In_550);
or U472 (N_472,In_345,In_650);
nor U473 (N_473,In_277,In_265);
nand U474 (N_474,In_469,In_626);
or U475 (N_475,In_515,In_480);
nor U476 (N_476,In_743,In_372);
nand U477 (N_477,In_618,In_268);
or U478 (N_478,In_118,In_741);
nor U479 (N_479,In_165,In_686);
xor U480 (N_480,In_495,In_624);
nand U481 (N_481,In_274,In_294);
nor U482 (N_482,In_103,In_319);
nor U483 (N_483,In_303,In_382);
nor U484 (N_484,In_681,In_144);
xor U485 (N_485,In_691,In_310);
and U486 (N_486,In_34,In_227);
or U487 (N_487,In_195,In_385);
nand U488 (N_488,In_583,In_12);
nand U489 (N_489,In_737,In_41);
or U490 (N_490,In_179,In_101);
and U491 (N_491,In_632,In_509);
nand U492 (N_492,In_726,In_456);
xor U493 (N_493,In_535,In_472);
nor U494 (N_494,In_458,In_165);
nand U495 (N_495,In_327,In_357);
and U496 (N_496,In_396,In_143);
nor U497 (N_497,In_492,In_609);
xor U498 (N_498,In_72,In_689);
and U499 (N_499,In_668,In_511);
nor U500 (N_500,N_417,N_494);
nor U501 (N_501,N_278,N_482);
xnor U502 (N_502,N_246,N_327);
or U503 (N_503,N_203,N_132);
nand U504 (N_504,N_336,N_234);
xnor U505 (N_505,N_75,N_484);
or U506 (N_506,N_253,N_287);
nand U507 (N_507,N_56,N_331);
nand U508 (N_508,N_399,N_83);
and U509 (N_509,N_88,N_361);
and U510 (N_510,N_163,N_76);
and U511 (N_511,N_230,N_215);
nor U512 (N_512,N_47,N_479);
nor U513 (N_513,N_60,N_339);
and U514 (N_514,N_323,N_174);
or U515 (N_515,N_410,N_413);
and U516 (N_516,N_297,N_492);
nor U517 (N_517,N_267,N_443);
nor U518 (N_518,N_370,N_344);
nand U519 (N_519,N_292,N_342);
nor U520 (N_520,N_462,N_309);
xnor U521 (N_521,N_397,N_69);
and U522 (N_522,N_487,N_362);
or U523 (N_523,N_464,N_70);
nand U524 (N_524,N_224,N_57);
xor U525 (N_525,N_185,N_142);
nor U526 (N_526,N_85,N_383);
nand U527 (N_527,N_145,N_369);
nand U528 (N_528,N_212,N_178);
xor U529 (N_529,N_66,N_28);
nor U530 (N_530,N_472,N_67);
and U531 (N_531,N_176,N_294);
and U532 (N_532,N_241,N_460);
or U533 (N_533,N_293,N_468);
or U534 (N_534,N_221,N_123);
and U535 (N_535,N_202,N_415);
nor U536 (N_536,N_391,N_190);
nor U537 (N_537,N_177,N_282);
nand U538 (N_538,N_473,N_52);
xnor U539 (N_539,N_108,N_244);
xor U540 (N_540,N_120,N_433);
xnor U541 (N_541,N_245,N_73);
xnor U542 (N_542,N_251,N_262);
and U543 (N_543,N_305,N_430);
nor U544 (N_544,N_191,N_345);
and U545 (N_545,N_124,N_161);
xnor U546 (N_546,N_50,N_384);
and U547 (N_547,N_208,N_197);
nand U548 (N_548,N_450,N_420);
nand U549 (N_549,N_377,N_49);
or U550 (N_550,N_189,N_233);
and U551 (N_551,N_381,N_222);
xor U552 (N_552,N_480,N_419);
nand U553 (N_553,N_112,N_330);
nand U554 (N_554,N_214,N_493);
and U555 (N_555,N_303,N_153);
and U556 (N_556,N_280,N_78);
xor U557 (N_557,N_31,N_347);
or U558 (N_558,N_187,N_119);
nor U559 (N_559,N_395,N_11);
nand U560 (N_560,N_9,N_439);
nor U561 (N_561,N_401,N_429);
nand U562 (N_562,N_40,N_160);
and U563 (N_563,N_220,N_201);
nand U564 (N_564,N_98,N_18);
xnor U565 (N_565,N_48,N_352);
or U566 (N_566,N_90,N_459);
and U567 (N_567,N_216,N_170);
or U568 (N_568,N_348,N_0);
nor U569 (N_569,N_407,N_263);
nand U570 (N_570,N_276,N_194);
and U571 (N_571,N_68,N_326);
or U572 (N_572,N_360,N_475);
nand U573 (N_573,N_269,N_324);
nand U574 (N_574,N_89,N_325);
nand U575 (N_575,N_34,N_416);
or U576 (N_576,N_300,N_42);
nand U577 (N_577,N_77,N_490);
nor U578 (N_578,N_219,N_72);
and U579 (N_579,N_62,N_288);
xnor U580 (N_580,N_449,N_350);
or U581 (N_581,N_435,N_489);
nand U582 (N_582,N_496,N_321);
or U583 (N_583,N_165,N_126);
xor U584 (N_584,N_301,N_143);
xor U585 (N_585,N_110,N_10);
xnor U586 (N_586,N_211,N_334);
and U587 (N_587,N_408,N_129);
xnor U588 (N_588,N_226,N_118);
nand U589 (N_589,N_95,N_146);
nor U590 (N_590,N_104,N_147);
or U591 (N_591,N_355,N_235);
and U592 (N_592,N_242,N_109);
xor U593 (N_593,N_273,N_284);
xor U594 (N_594,N_225,N_228);
and U595 (N_595,N_389,N_250);
and U596 (N_596,N_29,N_15);
xnor U597 (N_597,N_44,N_354);
and U598 (N_598,N_368,N_398);
nand U599 (N_599,N_283,N_38);
xor U600 (N_600,N_434,N_266);
xor U601 (N_601,N_247,N_396);
nand U602 (N_602,N_116,N_27);
nor U603 (N_603,N_101,N_454);
and U604 (N_604,N_356,N_337);
xnor U605 (N_605,N_128,N_30);
nand U606 (N_606,N_469,N_181);
xor U607 (N_607,N_12,N_257);
or U608 (N_608,N_55,N_311);
xor U609 (N_609,N_335,N_364);
and U610 (N_610,N_373,N_418);
or U611 (N_611,N_313,N_382);
and U612 (N_612,N_259,N_387);
nand U613 (N_613,N_385,N_173);
or U614 (N_614,N_80,N_23);
xor U615 (N_615,N_409,N_199);
or U616 (N_616,N_107,N_366);
nand U617 (N_617,N_150,N_299);
or U618 (N_618,N_476,N_317);
and U619 (N_619,N_111,N_394);
or U620 (N_620,N_333,N_148);
nor U621 (N_621,N_205,N_22);
xor U622 (N_622,N_236,N_471);
and U623 (N_623,N_87,N_427);
and U624 (N_624,N_268,N_204);
and U625 (N_625,N_314,N_281);
and U626 (N_626,N_65,N_100);
and U627 (N_627,N_96,N_239);
and U628 (N_628,N_367,N_358);
and U629 (N_629,N_180,N_285);
nor U630 (N_630,N_451,N_254);
nand U631 (N_631,N_54,N_441);
nand U632 (N_632,N_351,N_25);
nor U633 (N_633,N_179,N_315);
xnor U634 (N_634,N_156,N_372);
nand U635 (N_635,N_264,N_32);
nor U636 (N_636,N_117,N_470);
and U637 (N_637,N_209,N_298);
nor U638 (N_638,N_414,N_453);
and U639 (N_639,N_63,N_491);
xnor U640 (N_640,N_444,N_155);
nand U641 (N_641,N_33,N_388);
or U642 (N_642,N_227,N_171);
nor U643 (N_643,N_320,N_138);
or U644 (N_644,N_376,N_229);
or U645 (N_645,N_94,N_162);
or U646 (N_646,N_478,N_3);
xor U647 (N_647,N_74,N_270);
and U648 (N_648,N_167,N_19);
xor U649 (N_649,N_5,N_455);
xor U650 (N_650,N_477,N_402);
nor U651 (N_651,N_458,N_465);
or U652 (N_652,N_91,N_374);
or U653 (N_653,N_252,N_188);
and U654 (N_654,N_426,N_349);
nand U655 (N_655,N_483,N_137);
and U656 (N_656,N_41,N_379);
xor U657 (N_657,N_498,N_277);
and U658 (N_658,N_79,N_248);
nor U659 (N_659,N_316,N_58);
and U660 (N_660,N_103,N_365);
and U661 (N_661,N_403,N_461);
or U662 (N_662,N_265,N_196);
or U663 (N_663,N_121,N_279);
xor U664 (N_664,N_158,N_442);
and U665 (N_665,N_343,N_412);
xnor U666 (N_666,N_405,N_206);
nand U667 (N_667,N_424,N_291);
or U668 (N_668,N_275,N_428);
nand U669 (N_669,N_114,N_411);
xor U670 (N_670,N_237,N_456);
nand U671 (N_671,N_115,N_390);
nor U672 (N_672,N_488,N_7);
nor U673 (N_673,N_271,N_122);
xor U674 (N_674,N_463,N_231);
or U675 (N_675,N_125,N_332);
nor U676 (N_676,N_71,N_141);
or U677 (N_677,N_312,N_217);
nor U678 (N_678,N_8,N_436);
nor U679 (N_679,N_166,N_406);
xnor U680 (N_680,N_393,N_329);
nand U681 (N_681,N_290,N_422);
or U682 (N_682,N_218,N_159);
and U683 (N_683,N_249,N_431);
nor U684 (N_684,N_2,N_274);
xnor U685 (N_685,N_380,N_136);
nor U686 (N_686,N_447,N_183);
or U687 (N_687,N_485,N_82);
nand U688 (N_688,N_497,N_13);
xnor U689 (N_689,N_37,N_131);
xnor U690 (N_690,N_474,N_175);
nand U691 (N_691,N_113,N_21);
xor U692 (N_692,N_446,N_322);
and U693 (N_693,N_260,N_371);
nand U694 (N_694,N_39,N_296);
or U695 (N_695,N_445,N_93);
xnor U696 (N_696,N_168,N_289);
nand U697 (N_697,N_164,N_17);
xor U698 (N_698,N_213,N_400);
or U699 (N_699,N_328,N_363);
nor U700 (N_700,N_423,N_357);
or U701 (N_701,N_154,N_255);
nor U702 (N_702,N_36,N_139);
xnor U703 (N_703,N_61,N_272);
nand U704 (N_704,N_448,N_20);
xor U705 (N_705,N_157,N_238);
or U706 (N_706,N_1,N_210);
nand U707 (N_707,N_35,N_24);
and U708 (N_708,N_64,N_192);
or U709 (N_709,N_14,N_425);
xnor U710 (N_710,N_140,N_457);
nand U711 (N_711,N_346,N_134);
nor U712 (N_712,N_46,N_319);
and U713 (N_713,N_184,N_452);
or U714 (N_714,N_102,N_149);
xnor U715 (N_715,N_133,N_169);
nor U716 (N_716,N_375,N_404);
xnor U717 (N_717,N_304,N_438);
or U718 (N_718,N_302,N_386);
nor U719 (N_719,N_198,N_135);
or U720 (N_720,N_440,N_378);
nand U721 (N_721,N_51,N_261);
and U722 (N_722,N_340,N_295);
and U723 (N_723,N_243,N_338);
nor U724 (N_724,N_43,N_392);
and U725 (N_725,N_341,N_467);
and U726 (N_726,N_240,N_437);
xnor U727 (N_727,N_59,N_105);
and U728 (N_728,N_152,N_256);
nor U729 (N_729,N_353,N_481);
nor U730 (N_730,N_144,N_499);
xnor U731 (N_731,N_84,N_307);
nand U732 (N_732,N_232,N_306);
xor U733 (N_733,N_359,N_92);
or U734 (N_734,N_130,N_16);
and U735 (N_735,N_421,N_6);
xnor U736 (N_736,N_106,N_186);
xor U737 (N_737,N_223,N_486);
nor U738 (N_738,N_182,N_172);
and U739 (N_739,N_308,N_310);
nand U740 (N_740,N_495,N_45);
nor U741 (N_741,N_53,N_127);
xnor U742 (N_742,N_466,N_81);
nand U743 (N_743,N_258,N_195);
or U744 (N_744,N_86,N_97);
nand U745 (N_745,N_318,N_99);
nand U746 (N_746,N_200,N_193);
and U747 (N_747,N_432,N_4);
and U748 (N_748,N_286,N_151);
nor U749 (N_749,N_207,N_26);
or U750 (N_750,N_58,N_326);
nor U751 (N_751,N_268,N_389);
or U752 (N_752,N_440,N_202);
nand U753 (N_753,N_213,N_228);
or U754 (N_754,N_383,N_457);
nand U755 (N_755,N_105,N_439);
nand U756 (N_756,N_36,N_173);
and U757 (N_757,N_236,N_168);
or U758 (N_758,N_182,N_304);
xor U759 (N_759,N_343,N_217);
and U760 (N_760,N_414,N_182);
or U761 (N_761,N_299,N_400);
nand U762 (N_762,N_314,N_483);
nand U763 (N_763,N_283,N_72);
nor U764 (N_764,N_443,N_366);
xor U765 (N_765,N_23,N_168);
nor U766 (N_766,N_71,N_102);
or U767 (N_767,N_439,N_251);
or U768 (N_768,N_324,N_144);
and U769 (N_769,N_92,N_202);
nor U770 (N_770,N_415,N_491);
and U771 (N_771,N_50,N_174);
nand U772 (N_772,N_486,N_409);
nor U773 (N_773,N_219,N_7);
and U774 (N_774,N_64,N_315);
and U775 (N_775,N_216,N_485);
nor U776 (N_776,N_445,N_269);
xnor U777 (N_777,N_99,N_9);
nand U778 (N_778,N_279,N_310);
xnor U779 (N_779,N_176,N_287);
nor U780 (N_780,N_145,N_67);
and U781 (N_781,N_484,N_259);
nor U782 (N_782,N_346,N_385);
xor U783 (N_783,N_298,N_204);
xor U784 (N_784,N_21,N_472);
nand U785 (N_785,N_136,N_47);
nand U786 (N_786,N_359,N_188);
xnor U787 (N_787,N_147,N_201);
nor U788 (N_788,N_258,N_309);
and U789 (N_789,N_74,N_386);
nand U790 (N_790,N_449,N_469);
xor U791 (N_791,N_86,N_298);
xor U792 (N_792,N_437,N_31);
nand U793 (N_793,N_315,N_305);
nand U794 (N_794,N_160,N_352);
or U795 (N_795,N_472,N_271);
or U796 (N_796,N_452,N_212);
nor U797 (N_797,N_28,N_285);
or U798 (N_798,N_461,N_413);
xnor U799 (N_799,N_334,N_50);
xnor U800 (N_800,N_283,N_62);
xnor U801 (N_801,N_161,N_397);
nand U802 (N_802,N_83,N_455);
xor U803 (N_803,N_61,N_252);
nor U804 (N_804,N_197,N_124);
nand U805 (N_805,N_134,N_2);
nor U806 (N_806,N_229,N_21);
nand U807 (N_807,N_443,N_97);
and U808 (N_808,N_464,N_172);
or U809 (N_809,N_468,N_68);
or U810 (N_810,N_342,N_424);
and U811 (N_811,N_281,N_336);
xor U812 (N_812,N_454,N_165);
nor U813 (N_813,N_71,N_72);
and U814 (N_814,N_145,N_313);
nor U815 (N_815,N_122,N_24);
or U816 (N_816,N_53,N_415);
or U817 (N_817,N_470,N_254);
xnor U818 (N_818,N_251,N_444);
nor U819 (N_819,N_446,N_416);
nand U820 (N_820,N_469,N_21);
or U821 (N_821,N_121,N_327);
nor U822 (N_822,N_302,N_120);
or U823 (N_823,N_65,N_494);
nor U824 (N_824,N_382,N_293);
nand U825 (N_825,N_479,N_233);
and U826 (N_826,N_345,N_436);
or U827 (N_827,N_404,N_418);
nor U828 (N_828,N_166,N_44);
nand U829 (N_829,N_11,N_120);
nor U830 (N_830,N_40,N_476);
nand U831 (N_831,N_23,N_199);
xor U832 (N_832,N_499,N_157);
nor U833 (N_833,N_133,N_17);
and U834 (N_834,N_423,N_70);
nand U835 (N_835,N_16,N_247);
and U836 (N_836,N_416,N_268);
nor U837 (N_837,N_34,N_321);
nand U838 (N_838,N_116,N_268);
xor U839 (N_839,N_261,N_452);
nor U840 (N_840,N_184,N_178);
nor U841 (N_841,N_238,N_222);
or U842 (N_842,N_340,N_439);
or U843 (N_843,N_280,N_249);
nand U844 (N_844,N_351,N_284);
nand U845 (N_845,N_226,N_394);
and U846 (N_846,N_467,N_322);
xor U847 (N_847,N_319,N_277);
nor U848 (N_848,N_451,N_354);
xor U849 (N_849,N_231,N_312);
xor U850 (N_850,N_23,N_277);
xor U851 (N_851,N_122,N_211);
nand U852 (N_852,N_335,N_108);
nor U853 (N_853,N_120,N_314);
xor U854 (N_854,N_221,N_27);
xor U855 (N_855,N_362,N_243);
and U856 (N_856,N_219,N_426);
or U857 (N_857,N_282,N_221);
or U858 (N_858,N_135,N_326);
nor U859 (N_859,N_381,N_125);
nand U860 (N_860,N_335,N_153);
nor U861 (N_861,N_125,N_361);
and U862 (N_862,N_159,N_223);
or U863 (N_863,N_140,N_435);
and U864 (N_864,N_480,N_481);
nor U865 (N_865,N_1,N_496);
nand U866 (N_866,N_481,N_451);
xnor U867 (N_867,N_170,N_489);
nand U868 (N_868,N_8,N_219);
xnor U869 (N_869,N_473,N_264);
or U870 (N_870,N_332,N_350);
or U871 (N_871,N_233,N_210);
nand U872 (N_872,N_125,N_160);
nand U873 (N_873,N_124,N_456);
nand U874 (N_874,N_299,N_286);
or U875 (N_875,N_357,N_440);
or U876 (N_876,N_128,N_318);
and U877 (N_877,N_10,N_186);
nand U878 (N_878,N_443,N_484);
nor U879 (N_879,N_304,N_448);
and U880 (N_880,N_478,N_197);
nor U881 (N_881,N_345,N_80);
and U882 (N_882,N_397,N_460);
nor U883 (N_883,N_438,N_403);
and U884 (N_884,N_470,N_286);
and U885 (N_885,N_147,N_289);
and U886 (N_886,N_194,N_176);
nor U887 (N_887,N_314,N_187);
nor U888 (N_888,N_232,N_285);
xnor U889 (N_889,N_105,N_88);
or U890 (N_890,N_5,N_424);
nor U891 (N_891,N_267,N_63);
nand U892 (N_892,N_27,N_319);
nand U893 (N_893,N_323,N_116);
or U894 (N_894,N_240,N_120);
nor U895 (N_895,N_494,N_467);
nor U896 (N_896,N_451,N_223);
nor U897 (N_897,N_393,N_413);
nor U898 (N_898,N_201,N_479);
and U899 (N_899,N_458,N_227);
nor U900 (N_900,N_170,N_132);
xnor U901 (N_901,N_155,N_358);
nor U902 (N_902,N_228,N_352);
and U903 (N_903,N_248,N_294);
nor U904 (N_904,N_471,N_492);
and U905 (N_905,N_493,N_59);
and U906 (N_906,N_411,N_464);
or U907 (N_907,N_317,N_70);
and U908 (N_908,N_456,N_196);
and U909 (N_909,N_258,N_216);
nor U910 (N_910,N_368,N_325);
and U911 (N_911,N_367,N_172);
nor U912 (N_912,N_246,N_110);
or U913 (N_913,N_350,N_165);
and U914 (N_914,N_52,N_217);
nand U915 (N_915,N_213,N_122);
and U916 (N_916,N_415,N_92);
and U917 (N_917,N_95,N_117);
or U918 (N_918,N_472,N_259);
and U919 (N_919,N_439,N_92);
nand U920 (N_920,N_380,N_211);
or U921 (N_921,N_274,N_220);
or U922 (N_922,N_62,N_193);
and U923 (N_923,N_88,N_157);
nand U924 (N_924,N_103,N_187);
nor U925 (N_925,N_332,N_171);
nand U926 (N_926,N_12,N_298);
nand U927 (N_927,N_266,N_335);
nand U928 (N_928,N_284,N_197);
nand U929 (N_929,N_272,N_406);
and U930 (N_930,N_293,N_404);
or U931 (N_931,N_435,N_243);
nand U932 (N_932,N_192,N_419);
xor U933 (N_933,N_209,N_176);
xor U934 (N_934,N_372,N_474);
or U935 (N_935,N_39,N_371);
or U936 (N_936,N_266,N_24);
nor U937 (N_937,N_454,N_201);
xor U938 (N_938,N_136,N_173);
and U939 (N_939,N_390,N_480);
nand U940 (N_940,N_449,N_156);
and U941 (N_941,N_118,N_242);
xor U942 (N_942,N_20,N_495);
or U943 (N_943,N_461,N_496);
or U944 (N_944,N_240,N_334);
and U945 (N_945,N_148,N_385);
and U946 (N_946,N_145,N_359);
xor U947 (N_947,N_356,N_150);
xnor U948 (N_948,N_376,N_426);
and U949 (N_949,N_426,N_216);
and U950 (N_950,N_41,N_399);
nand U951 (N_951,N_390,N_338);
or U952 (N_952,N_237,N_69);
or U953 (N_953,N_18,N_248);
nor U954 (N_954,N_108,N_120);
nand U955 (N_955,N_350,N_3);
xor U956 (N_956,N_410,N_344);
nor U957 (N_957,N_460,N_167);
and U958 (N_958,N_406,N_395);
xnor U959 (N_959,N_303,N_293);
and U960 (N_960,N_94,N_156);
or U961 (N_961,N_23,N_482);
and U962 (N_962,N_479,N_252);
xnor U963 (N_963,N_80,N_319);
and U964 (N_964,N_408,N_222);
nor U965 (N_965,N_421,N_412);
and U966 (N_966,N_367,N_424);
nor U967 (N_967,N_198,N_54);
or U968 (N_968,N_437,N_353);
or U969 (N_969,N_231,N_386);
and U970 (N_970,N_6,N_273);
nor U971 (N_971,N_340,N_213);
nor U972 (N_972,N_325,N_353);
or U973 (N_973,N_372,N_242);
nor U974 (N_974,N_92,N_219);
nor U975 (N_975,N_427,N_349);
or U976 (N_976,N_85,N_195);
xor U977 (N_977,N_6,N_407);
or U978 (N_978,N_483,N_3);
nor U979 (N_979,N_352,N_13);
xor U980 (N_980,N_352,N_300);
xnor U981 (N_981,N_491,N_47);
nor U982 (N_982,N_154,N_477);
and U983 (N_983,N_472,N_423);
nor U984 (N_984,N_427,N_476);
nor U985 (N_985,N_169,N_443);
or U986 (N_986,N_469,N_34);
nand U987 (N_987,N_194,N_430);
or U988 (N_988,N_66,N_463);
nand U989 (N_989,N_413,N_287);
or U990 (N_990,N_187,N_11);
or U991 (N_991,N_322,N_498);
nor U992 (N_992,N_94,N_330);
or U993 (N_993,N_425,N_190);
xnor U994 (N_994,N_68,N_120);
nor U995 (N_995,N_312,N_133);
nor U996 (N_996,N_108,N_394);
nand U997 (N_997,N_222,N_142);
nand U998 (N_998,N_475,N_279);
nand U999 (N_999,N_101,N_316);
xor U1000 (N_1000,N_796,N_649);
xnor U1001 (N_1001,N_933,N_571);
or U1002 (N_1002,N_801,N_524);
and U1003 (N_1003,N_505,N_899);
and U1004 (N_1004,N_566,N_851);
or U1005 (N_1005,N_529,N_836);
nand U1006 (N_1006,N_884,N_690);
xnor U1007 (N_1007,N_647,N_810);
xnor U1008 (N_1008,N_693,N_778);
or U1009 (N_1009,N_597,N_931);
or U1010 (N_1010,N_754,N_717);
or U1011 (N_1011,N_946,N_808);
or U1012 (N_1012,N_681,N_977);
nor U1013 (N_1013,N_695,N_722);
nor U1014 (N_1014,N_903,N_557);
nand U1015 (N_1015,N_603,N_767);
or U1016 (N_1016,N_518,N_615);
and U1017 (N_1017,N_763,N_503);
nor U1018 (N_1018,N_756,N_687);
or U1019 (N_1019,N_830,N_611);
or U1020 (N_1020,N_626,N_959);
and U1021 (N_1021,N_636,N_525);
and U1022 (N_1022,N_547,N_844);
nand U1023 (N_1023,N_817,N_932);
nor U1024 (N_1024,N_834,N_877);
or U1025 (N_1025,N_981,N_545);
nand U1026 (N_1026,N_755,N_820);
nor U1027 (N_1027,N_869,N_749);
nand U1028 (N_1028,N_800,N_502);
nand U1029 (N_1029,N_881,N_898);
nand U1030 (N_1030,N_913,N_821);
nand U1031 (N_1031,N_573,N_788);
nand U1032 (N_1032,N_961,N_720);
and U1033 (N_1033,N_856,N_744);
nor U1034 (N_1034,N_882,N_811);
or U1035 (N_1035,N_991,N_731);
nand U1036 (N_1036,N_960,N_923);
and U1037 (N_1037,N_515,N_747);
or U1038 (N_1038,N_674,N_567);
or U1039 (N_1039,N_848,N_516);
nor U1040 (N_1040,N_842,N_945);
and U1041 (N_1041,N_528,N_766);
nor U1042 (N_1042,N_535,N_713);
nand U1043 (N_1043,N_812,N_908);
nand U1044 (N_1044,N_694,N_617);
xnor U1045 (N_1045,N_803,N_875);
xor U1046 (N_1046,N_580,N_829);
or U1047 (N_1047,N_601,N_520);
or U1048 (N_1048,N_828,N_854);
and U1049 (N_1049,N_980,N_789);
nand U1050 (N_1050,N_813,N_986);
nand U1051 (N_1051,N_537,N_760);
xnor U1052 (N_1052,N_950,N_994);
nand U1053 (N_1053,N_770,N_582);
xnor U1054 (N_1054,N_637,N_833);
xnor U1055 (N_1055,N_809,N_857);
nor U1056 (N_1056,N_584,N_939);
nor U1057 (N_1057,N_643,N_609);
nor U1058 (N_1058,N_952,N_546);
or U1059 (N_1059,N_753,N_879);
or U1060 (N_1060,N_562,N_688);
nand U1061 (N_1061,N_581,N_886);
xor U1062 (N_1062,N_995,N_565);
or U1063 (N_1063,N_534,N_672);
and U1064 (N_1064,N_937,N_924);
xnor U1065 (N_1065,N_954,N_594);
or U1066 (N_1066,N_948,N_559);
and U1067 (N_1067,N_521,N_673);
and U1068 (N_1068,N_867,N_911);
or U1069 (N_1069,N_530,N_662);
nand U1070 (N_1070,N_832,N_506);
xor U1071 (N_1071,N_648,N_987);
and U1072 (N_1072,N_577,N_839);
nand U1073 (N_1073,N_705,N_940);
xor U1074 (N_1074,N_508,N_587);
nand U1075 (N_1075,N_791,N_942);
nand U1076 (N_1076,N_659,N_783);
or U1077 (N_1077,N_676,N_989);
nor U1078 (N_1078,N_777,N_707);
xnor U1079 (N_1079,N_905,N_831);
nor U1080 (N_1080,N_644,N_576);
and U1081 (N_1081,N_645,N_727);
or U1082 (N_1082,N_764,N_919);
nor U1083 (N_1083,N_975,N_876);
nor U1084 (N_1084,N_752,N_852);
xor U1085 (N_1085,N_759,N_918);
and U1086 (N_1086,N_733,N_703);
nor U1087 (N_1087,N_982,N_550);
nand U1088 (N_1088,N_901,N_742);
or U1089 (N_1089,N_976,N_893);
or U1090 (N_1090,N_910,N_596);
nor U1091 (N_1091,N_679,N_929);
or U1092 (N_1092,N_664,N_953);
and U1093 (N_1093,N_974,N_885);
nand U1094 (N_1094,N_962,N_552);
xor U1095 (N_1095,N_712,N_883);
nor U1096 (N_1096,N_988,N_838);
nor U1097 (N_1097,N_650,N_651);
xnor U1098 (N_1098,N_627,N_790);
and U1099 (N_1099,N_914,N_668);
and U1100 (N_1100,N_678,N_523);
or U1101 (N_1101,N_549,N_787);
or U1102 (N_1102,N_775,N_589);
xnor U1103 (N_1103,N_973,N_804);
nand U1104 (N_1104,N_978,N_631);
nand U1105 (N_1105,N_697,N_938);
nor U1106 (N_1106,N_585,N_504);
and U1107 (N_1107,N_769,N_640);
or U1108 (N_1108,N_861,N_511);
nand U1109 (N_1109,N_999,N_880);
xnor U1110 (N_1110,N_564,N_837);
and U1111 (N_1111,N_887,N_781);
nand U1112 (N_1112,N_927,N_512);
xnor U1113 (N_1113,N_997,N_554);
or U1114 (N_1114,N_806,N_658);
or U1115 (N_1115,N_802,N_963);
nor U1116 (N_1116,N_639,N_930);
and U1117 (N_1117,N_873,N_711);
and U1118 (N_1118,N_538,N_616);
and U1119 (N_1119,N_814,N_827);
nor U1120 (N_1120,N_993,N_934);
nand U1121 (N_1121,N_598,N_865);
xnor U1122 (N_1122,N_620,N_665);
nor U1123 (N_1123,N_638,N_655);
nand U1124 (N_1124,N_556,N_500);
and U1125 (N_1125,N_907,N_970);
and U1126 (N_1126,N_536,N_772);
xor U1127 (N_1127,N_900,N_702);
and U1128 (N_1128,N_710,N_670);
nand U1129 (N_1129,N_544,N_728);
nand U1130 (N_1130,N_642,N_773);
nand U1131 (N_1131,N_669,N_780);
xnor U1132 (N_1132,N_872,N_849);
and U1133 (N_1133,N_714,N_721);
or U1134 (N_1134,N_941,N_758);
nand U1135 (N_1135,N_855,N_998);
or U1136 (N_1136,N_917,N_894);
nand U1137 (N_1137,N_588,N_915);
and U1138 (N_1138,N_983,N_569);
and U1139 (N_1139,N_606,N_685);
xor U1140 (N_1140,N_540,N_969);
xnor U1141 (N_1141,N_850,N_956);
nor U1142 (N_1142,N_807,N_586);
nor U1143 (N_1143,N_716,N_654);
nand U1144 (N_1144,N_936,N_951);
xnor U1145 (N_1145,N_684,N_990);
nor U1146 (N_1146,N_660,N_926);
nand U1147 (N_1147,N_698,N_671);
nor U1148 (N_1148,N_682,N_633);
xor U1149 (N_1149,N_735,N_708);
nand U1150 (N_1150,N_677,N_964);
and U1151 (N_1151,N_602,N_514);
xnor U1152 (N_1152,N_561,N_785);
and U1153 (N_1153,N_641,N_966);
nand U1154 (N_1154,N_771,N_551);
and U1155 (N_1155,N_526,N_510);
xor U1156 (N_1156,N_570,N_859);
and U1157 (N_1157,N_751,N_965);
nand U1158 (N_1158,N_696,N_578);
and U1159 (N_1159,N_745,N_605);
nor U1160 (N_1160,N_740,N_958);
nor U1161 (N_1161,N_661,N_748);
nand U1162 (N_1162,N_864,N_870);
and U1163 (N_1163,N_574,N_621);
nor U1164 (N_1164,N_675,N_794);
and U1165 (N_1165,N_835,N_853);
or U1166 (N_1166,N_701,N_909);
and U1167 (N_1167,N_610,N_736);
and U1168 (N_1168,N_619,N_624);
xnor U1169 (N_1169,N_968,N_683);
nand U1170 (N_1170,N_663,N_513);
xnor U1171 (N_1171,N_704,N_723);
and U1172 (N_1172,N_501,N_608);
nor U1173 (N_1173,N_522,N_579);
xnor U1174 (N_1174,N_706,N_955);
nor U1175 (N_1175,N_823,N_743);
xor U1176 (N_1176,N_692,N_762);
or U1177 (N_1177,N_667,N_891);
nor U1178 (N_1178,N_622,N_607);
nor U1179 (N_1179,N_846,N_825);
nand U1180 (N_1180,N_985,N_739);
nor U1181 (N_1181,N_623,N_774);
or U1182 (N_1182,N_657,N_847);
and U1183 (N_1183,N_614,N_819);
nand U1184 (N_1184,N_779,N_984);
nand U1185 (N_1185,N_737,N_730);
and U1186 (N_1186,N_822,N_527);
or U1187 (N_1187,N_878,N_591);
or U1188 (N_1188,N_784,N_972);
nor U1189 (N_1189,N_724,N_583);
nor U1190 (N_1190,N_533,N_904);
nor U1191 (N_1191,N_996,N_943);
nand U1192 (N_1192,N_746,N_572);
xor U1193 (N_1193,N_888,N_815);
xor U1194 (N_1194,N_845,N_653);
nand U1195 (N_1195,N_890,N_792);
nor U1196 (N_1196,N_531,N_532);
or U1197 (N_1197,N_971,N_656);
or U1198 (N_1198,N_889,N_863);
or U1199 (N_1199,N_841,N_866);
xor U1200 (N_1200,N_874,N_592);
xor U1201 (N_1201,N_519,N_797);
nand U1202 (N_1202,N_560,N_738);
or U1203 (N_1203,N_793,N_595);
nor U1204 (N_1204,N_840,N_912);
or U1205 (N_1205,N_613,N_539);
nor U1206 (N_1206,N_699,N_700);
xor U1207 (N_1207,N_776,N_593);
xor U1208 (N_1208,N_947,N_761);
and U1209 (N_1209,N_858,N_563);
nor U1210 (N_1210,N_921,N_741);
and U1211 (N_1211,N_786,N_646);
and U1212 (N_1212,N_862,N_928);
nand U1213 (N_1213,N_612,N_604);
nand U1214 (N_1214,N_553,N_826);
xnor U1215 (N_1215,N_542,N_719);
and U1216 (N_1216,N_600,N_892);
nand U1217 (N_1217,N_944,N_732);
or U1218 (N_1218,N_726,N_689);
and U1219 (N_1219,N_799,N_920);
and U1220 (N_1220,N_805,N_906);
xnor U1221 (N_1221,N_568,N_635);
and U1222 (N_1222,N_925,N_590);
and U1223 (N_1223,N_843,N_630);
xnor U1224 (N_1224,N_686,N_543);
nor U1225 (N_1225,N_718,N_725);
xnor U1226 (N_1226,N_750,N_967);
and U1227 (N_1227,N_795,N_628);
and U1228 (N_1228,N_871,N_757);
or U1229 (N_1229,N_902,N_895);
xnor U1230 (N_1230,N_715,N_558);
nand U1231 (N_1231,N_632,N_691);
nand U1232 (N_1232,N_625,N_957);
or U1233 (N_1233,N_666,N_765);
xnor U1234 (N_1234,N_541,N_798);
and U1235 (N_1235,N_868,N_507);
xnor U1236 (N_1236,N_734,N_916);
nor U1237 (N_1237,N_816,N_860);
nand U1238 (N_1238,N_935,N_922);
and U1239 (N_1239,N_629,N_729);
and U1240 (N_1240,N_634,N_509);
nor U1241 (N_1241,N_709,N_896);
xor U1242 (N_1242,N_652,N_979);
nor U1243 (N_1243,N_517,N_680);
and U1244 (N_1244,N_618,N_897);
or U1245 (N_1245,N_824,N_992);
and U1246 (N_1246,N_575,N_782);
or U1247 (N_1247,N_949,N_548);
nor U1248 (N_1248,N_818,N_555);
nand U1249 (N_1249,N_768,N_599);
xor U1250 (N_1250,N_987,N_766);
nor U1251 (N_1251,N_752,N_570);
nor U1252 (N_1252,N_645,N_974);
or U1253 (N_1253,N_519,N_658);
nor U1254 (N_1254,N_690,N_772);
xnor U1255 (N_1255,N_886,N_608);
xor U1256 (N_1256,N_940,N_532);
nor U1257 (N_1257,N_625,N_711);
or U1258 (N_1258,N_968,N_850);
nand U1259 (N_1259,N_734,N_865);
nor U1260 (N_1260,N_586,N_789);
and U1261 (N_1261,N_865,N_592);
and U1262 (N_1262,N_685,N_735);
or U1263 (N_1263,N_567,N_986);
nand U1264 (N_1264,N_858,N_648);
and U1265 (N_1265,N_949,N_607);
xor U1266 (N_1266,N_770,N_562);
nand U1267 (N_1267,N_636,N_713);
or U1268 (N_1268,N_744,N_700);
or U1269 (N_1269,N_711,N_890);
nor U1270 (N_1270,N_968,N_933);
or U1271 (N_1271,N_543,N_716);
or U1272 (N_1272,N_681,N_553);
and U1273 (N_1273,N_685,N_991);
or U1274 (N_1274,N_598,N_687);
and U1275 (N_1275,N_570,N_733);
nand U1276 (N_1276,N_969,N_626);
nand U1277 (N_1277,N_624,N_696);
or U1278 (N_1278,N_843,N_858);
nand U1279 (N_1279,N_627,N_638);
and U1280 (N_1280,N_512,N_929);
xnor U1281 (N_1281,N_870,N_939);
or U1282 (N_1282,N_987,N_649);
nor U1283 (N_1283,N_530,N_887);
nand U1284 (N_1284,N_721,N_693);
or U1285 (N_1285,N_582,N_839);
and U1286 (N_1286,N_508,N_530);
or U1287 (N_1287,N_852,N_815);
nand U1288 (N_1288,N_734,N_535);
xor U1289 (N_1289,N_585,N_807);
or U1290 (N_1290,N_692,N_815);
or U1291 (N_1291,N_643,N_893);
xor U1292 (N_1292,N_718,N_944);
nand U1293 (N_1293,N_570,N_897);
nor U1294 (N_1294,N_957,N_765);
and U1295 (N_1295,N_566,N_994);
nor U1296 (N_1296,N_763,N_722);
xnor U1297 (N_1297,N_855,N_961);
nor U1298 (N_1298,N_545,N_503);
xnor U1299 (N_1299,N_634,N_891);
or U1300 (N_1300,N_599,N_651);
nand U1301 (N_1301,N_729,N_559);
or U1302 (N_1302,N_523,N_749);
nand U1303 (N_1303,N_942,N_764);
nor U1304 (N_1304,N_941,N_996);
nor U1305 (N_1305,N_872,N_583);
xor U1306 (N_1306,N_834,N_711);
xnor U1307 (N_1307,N_939,N_972);
or U1308 (N_1308,N_732,N_565);
or U1309 (N_1309,N_540,N_509);
nand U1310 (N_1310,N_779,N_875);
or U1311 (N_1311,N_565,N_989);
or U1312 (N_1312,N_502,N_684);
nand U1313 (N_1313,N_725,N_647);
and U1314 (N_1314,N_633,N_584);
nor U1315 (N_1315,N_501,N_520);
and U1316 (N_1316,N_766,N_640);
and U1317 (N_1317,N_716,N_987);
nor U1318 (N_1318,N_836,N_928);
nand U1319 (N_1319,N_812,N_736);
and U1320 (N_1320,N_579,N_707);
and U1321 (N_1321,N_622,N_554);
and U1322 (N_1322,N_552,N_879);
nor U1323 (N_1323,N_647,N_957);
and U1324 (N_1324,N_594,N_585);
nor U1325 (N_1325,N_617,N_964);
xnor U1326 (N_1326,N_635,N_507);
xnor U1327 (N_1327,N_550,N_965);
nand U1328 (N_1328,N_794,N_548);
xnor U1329 (N_1329,N_639,N_569);
and U1330 (N_1330,N_736,N_900);
and U1331 (N_1331,N_602,N_654);
and U1332 (N_1332,N_537,N_609);
nor U1333 (N_1333,N_566,N_922);
xor U1334 (N_1334,N_912,N_915);
and U1335 (N_1335,N_613,N_542);
or U1336 (N_1336,N_709,N_879);
xor U1337 (N_1337,N_759,N_656);
xor U1338 (N_1338,N_928,N_731);
and U1339 (N_1339,N_853,N_752);
xnor U1340 (N_1340,N_603,N_789);
nand U1341 (N_1341,N_916,N_703);
nand U1342 (N_1342,N_660,N_741);
nand U1343 (N_1343,N_519,N_695);
or U1344 (N_1344,N_605,N_561);
and U1345 (N_1345,N_699,N_979);
nand U1346 (N_1346,N_660,N_958);
xnor U1347 (N_1347,N_852,N_983);
xnor U1348 (N_1348,N_505,N_883);
nor U1349 (N_1349,N_656,N_529);
xor U1350 (N_1350,N_548,N_931);
or U1351 (N_1351,N_514,N_909);
xnor U1352 (N_1352,N_504,N_917);
nand U1353 (N_1353,N_554,N_951);
and U1354 (N_1354,N_680,N_762);
or U1355 (N_1355,N_517,N_913);
or U1356 (N_1356,N_607,N_965);
and U1357 (N_1357,N_927,N_935);
nor U1358 (N_1358,N_645,N_897);
or U1359 (N_1359,N_919,N_901);
or U1360 (N_1360,N_768,N_832);
nor U1361 (N_1361,N_620,N_972);
and U1362 (N_1362,N_773,N_526);
nor U1363 (N_1363,N_677,N_774);
and U1364 (N_1364,N_539,N_916);
and U1365 (N_1365,N_569,N_613);
nand U1366 (N_1366,N_914,N_993);
or U1367 (N_1367,N_952,N_691);
nor U1368 (N_1368,N_940,N_691);
or U1369 (N_1369,N_561,N_672);
nor U1370 (N_1370,N_699,N_901);
nand U1371 (N_1371,N_532,N_947);
nor U1372 (N_1372,N_509,N_940);
or U1373 (N_1373,N_859,N_898);
or U1374 (N_1374,N_830,N_981);
xor U1375 (N_1375,N_613,N_507);
or U1376 (N_1376,N_666,N_994);
nand U1377 (N_1377,N_594,N_578);
nand U1378 (N_1378,N_740,N_556);
xnor U1379 (N_1379,N_787,N_839);
nand U1380 (N_1380,N_951,N_690);
nand U1381 (N_1381,N_551,N_954);
and U1382 (N_1382,N_588,N_532);
xor U1383 (N_1383,N_748,N_814);
nand U1384 (N_1384,N_795,N_766);
or U1385 (N_1385,N_543,N_728);
and U1386 (N_1386,N_812,N_934);
xor U1387 (N_1387,N_736,N_870);
or U1388 (N_1388,N_981,N_648);
xor U1389 (N_1389,N_947,N_720);
nor U1390 (N_1390,N_990,N_687);
xnor U1391 (N_1391,N_752,N_787);
or U1392 (N_1392,N_827,N_983);
and U1393 (N_1393,N_752,N_726);
or U1394 (N_1394,N_851,N_751);
and U1395 (N_1395,N_663,N_827);
nand U1396 (N_1396,N_628,N_742);
or U1397 (N_1397,N_585,N_550);
or U1398 (N_1398,N_603,N_562);
or U1399 (N_1399,N_899,N_654);
or U1400 (N_1400,N_766,N_868);
nand U1401 (N_1401,N_577,N_804);
xor U1402 (N_1402,N_552,N_728);
or U1403 (N_1403,N_979,N_822);
nand U1404 (N_1404,N_974,N_713);
or U1405 (N_1405,N_652,N_852);
xnor U1406 (N_1406,N_579,N_580);
xor U1407 (N_1407,N_808,N_631);
and U1408 (N_1408,N_639,N_670);
and U1409 (N_1409,N_686,N_748);
nand U1410 (N_1410,N_940,N_558);
and U1411 (N_1411,N_760,N_953);
nand U1412 (N_1412,N_555,N_562);
or U1413 (N_1413,N_903,N_552);
nor U1414 (N_1414,N_677,N_806);
and U1415 (N_1415,N_805,N_880);
xor U1416 (N_1416,N_954,N_922);
or U1417 (N_1417,N_655,N_634);
or U1418 (N_1418,N_972,N_960);
nand U1419 (N_1419,N_822,N_959);
or U1420 (N_1420,N_585,N_926);
nand U1421 (N_1421,N_999,N_879);
or U1422 (N_1422,N_518,N_795);
and U1423 (N_1423,N_923,N_597);
or U1424 (N_1424,N_649,N_601);
nor U1425 (N_1425,N_890,N_574);
and U1426 (N_1426,N_535,N_978);
and U1427 (N_1427,N_923,N_958);
nor U1428 (N_1428,N_854,N_981);
xor U1429 (N_1429,N_780,N_970);
nand U1430 (N_1430,N_802,N_763);
xnor U1431 (N_1431,N_669,N_579);
xnor U1432 (N_1432,N_919,N_889);
nor U1433 (N_1433,N_899,N_701);
and U1434 (N_1434,N_740,N_575);
and U1435 (N_1435,N_553,N_953);
and U1436 (N_1436,N_635,N_682);
xnor U1437 (N_1437,N_602,N_763);
and U1438 (N_1438,N_541,N_614);
and U1439 (N_1439,N_557,N_563);
xnor U1440 (N_1440,N_900,N_884);
nor U1441 (N_1441,N_952,N_791);
or U1442 (N_1442,N_950,N_614);
nor U1443 (N_1443,N_619,N_729);
nand U1444 (N_1444,N_949,N_596);
nand U1445 (N_1445,N_540,N_980);
nand U1446 (N_1446,N_935,N_628);
xnor U1447 (N_1447,N_988,N_896);
nor U1448 (N_1448,N_850,N_878);
nor U1449 (N_1449,N_722,N_687);
xnor U1450 (N_1450,N_741,N_770);
and U1451 (N_1451,N_659,N_936);
xnor U1452 (N_1452,N_732,N_558);
and U1453 (N_1453,N_739,N_746);
nand U1454 (N_1454,N_713,N_978);
nand U1455 (N_1455,N_824,N_675);
or U1456 (N_1456,N_584,N_721);
xor U1457 (N_1457,N_639,N_528);
nand U1458 (N_1458,N_787,N_631);
and U1459 (N_1459,N_844,N_503);
nand U1460 (N_1460,N_735,N_818);
nor U1461 (N_1461,N_824,N_601);
and U1462 (N_1462,N_789,N_614);
nand U1463 (N_1463,N_833,N_756);
or U1464 (N_1464,N_534,N_647);
xnor U1465 (N_1465,N_953,N_759);
nor U1466 (N_1466,N_867,N_577);
or U1467 (N_1467,N_740,N_637);
nand U1468 (N_1468,N_769,N_677);
nor U1469 (N_1469,N_875,N_651);
xnor U1470 (N_1470,N_881,N_702);
xor U1471 (N_1471,N_526,N_797);
and U1472 (N_1472,N_837,N_509);
and U1473 (N_1473,N_996,N_869);
and U1474 (N_1474,N_654,N_569);
or U1475 (N_1475,N_656,N_685);
nor U1476 (N_1476,N_766,N_681);
nor U1477 (N_1477,N_538,N_950);
xnor U1478 (N_1478,N_974,N_887);
nor U1479 (N_1479,N_980,N_838);
and U1480 (N_1480,N_891,N_666);
nor U1481 (N_1481,N_997,N_758);
nor U1482 (N_1482,N_594,N_971);
and U1483 (N_1483,N_847,N_683);
xor U1484 (N_1484,N_668,N_970);
or U1485 (N_1485,N_771,N_895);
nand U1486 (N_1486,N_736,N_878);
xor U1487 (N_1487,N_776,N_772);
or U1488 (N_1488,N_752,N_705);
or U1489 (N_1489,N_792,N_607);
nor U1490 (N_1490,N_826,N_872);
or U1491 (N_1491,N_789,N_920);
nor U1492 (N_1492,N_598,N_591);
nand U1493 (N_1493,N_860,N_748);
nand U1494 (N_1494,N_604,N_894);
xor U1495 (N_1495,N_643,N_788);
nand U1496 (N_1496,N_617,N_587);
xnor U1497 (N_1497,N_821,N_993);
or U1498 (N_1498,N_702,N_646);
xor U1499 (N_1499,N_941,N_519);
nand U1500 (N_1500,N_1259,N_1442);
nor U1501 (N_1501,N_1429,N_1353);
xor U1502 (N_1502,N_1072,N_1204);
nand U1503 (N_1503,N_1375,N_1203);
or U1504 (N_1504,N_1291,N_1330);
nand U1505 (N_1505,N_1369,N_1066);
or U1506 (N_1506,N_1361,N_1298);
or U1507 (N_1507,N_1338,N_1016);
nand U1508 (N_1508,N_1217,N_1230);
and U1509 (N_1509,N_1491,N_1385);
nand U1510 (N_1510,N_1024,N_1282);
and U1511 (N_1511,N_1246,N_1269);
or U1512 (N_1512,N_1003,N_1460);
or U1513 (N_1513,N_1015,N_1453);
nor U1514 (N_1514,N_1391,N_1010);
xnor U1515 (N_1515,N_1322,N_1105);
nor U1516 (N_1516,N_1107,N_1023);
nand U1517 (N_1517,N_1243,N_1323);
nor U1518 (N_1518,N_1043,N_1120);
or U1519 (N_1519,N_1441,N_1304);
nor U1520 (N_1520,N_1063,N_1077);
xor U1521 (N_1521,N_1394,N_1042);
xnor U1522 (N_1522,N_1214,N_1069);
or U1523 (N_1523,N_1218,N_1038);
nor U1524 (N_1524,N_1168,N_1412);
nor U1525 (N_1525,N_1183,N_1008);
nor U1526 (N_1526,N_1290,N_1134);
and U1527 (N_1527,N_1302,N_1007);
nor U1528 (N_1528,N_1462,N_1054);
or U1529 (N_1529,N_1033,N_1399);
nor U1530 (N_1530,N_1404,N_1374);
and U1531 (N_1531,N_1199,N_1157);
nor U1532 (N_1532,N_1414,N_1393);
and U1533 (N_1533,N_1045,N_1017);
or U1534 (N_1534,N_1140,N_1146);
nor U1535 (N_1535,N_1201,N_1459);
or U1536 (N_1536,N_1119,N_1215);
xor U1537 (N_1537,N_1294,N_1407);
nand U1538 (N_1538,N_1079,N_1430);
xnor U1539 (N_1539,N_1071,N_1397);
xnor U1540 (N_1540,N_1138,N_1306);
nand U1541 (N_1541,N_1152,N_1165);
xnor U1542 (N_1542,N_1435,N_1187);
or U1543 (N_1543,N_1360,N_1233);
xnor U1544 (N_1544,N_1293,N_1278);
or U1545 (N_1545,N_1347,N_1177);
nand U1546 (N_1546,N_1145,N_1110);
or U1547 (N_1547,N_1113,N_1026);
and U1548 (N_1548,N_1261,N_1185);
and U1549 (N_1549,N_1115,N_1193);
or U1550 (N_1550,N_1317,N_1175);
or U1551 (N_1551,N_1167,N_1213);
xnor U1552 (N_1552,N_1224,N_1277);
nor U1553 (N_1553,N_1482,N_1139);
or U1554 (N_1554,N_1315,N_1061);
nor U1555 (N_1555,N_1100,N_1422);
xnor U1556 (N_1556,N_1206,N_1104);
nand U1557 (N_1557,N_1471,N_1457);
xnor U1558 (N_1558,N_1254,N_1197);
nand U1559 (N_1559,N_1458,N_1235);
xor U1560 (N_1560,N_1301,N_1283);
nand U1561 (N_1561,N_1494,N_1247);
and U1562 (N_1562,N_1228,N_1162);
nand U1563 (N_1563,N_1195,N_1159);
nand U1564 (N_1564,N_1031,N_1091);
xnor U1565 (N_1565,N_1226,N_1078);
or U1566 (N_1566,N_1256,N_1194);
xnor U1567 (N_1567,N_1234,N_1281);
and U1568 (N_1568,N_1189,N_1192);
xnor U1569 (N_1569,N_1271,N_1171);
or U1570 (N_1570,N_1319,N_1497);
or U1571 (N_1571,N_1112,N_1173);
xnor U1572 (N_1572,N_1099,N_1341);
and U1573 (N_1573,N_1083,N_1350);
nor U1574 (N_1574,N_1439,N_1220);
or U1575 (N_1575,N_1499,N_1337);
and U1576 (N_1576,N_1287,N_1020);
and U1577 (N_1577,N_1464,N_1028);
or U1578 (N_1578,N_1292,N_1143);
xor U1579 (N_1579,N_1116,N_1202);
or U1580 (N_1580,N_1036,N_1046);
xor U1581 (N_1581,N_1090,N_1479);
nor U1582 (N_1582,N_1285,N_1465);
and U1583 (N_1583,N_1216,N_1095);
nor U1584 (N_1584,N_1027,N_1032);
nor U1585 (N_1585,N_1076,N_1073);
and U1586 (N_1586,N_1390,N_1142);
or U1587 (N_1587,N_1279,N_1419);
nor U1588 (N_1588,N_1000,N_1128);
xnor U1589 (N_1589,N_1005,N_1211);
or U1590 (N_1590,N_1280,N_1408);
xor U1591 (N_1591,N_1400,N_1469);
or U1592 (N_1592,N_1372,N_1082);
and U1593 (N_1593,N_1468,N_1300);
or U1594 (N_1594,N_1014,N_1483);
nand U1595 (N_1595,N_1373,N_1056);
nand U1596 (N_1596,N_1365,N_1263);
nand U1597 (N_1597,N_1198,N_1359);
nor U1598 (N_1598,N_1316,N_1172);
or U1599 (N_1599,N_1244,N_1225);
or U1600 (N_1600,N_1371,N_1018);
nand U1601 (N_1601,N_1455,N_1364);
or U1602 (N_1602,N_1219,N_1339);
or U1603 (N_1603,N_1039,N_1013);
nand U1604 (N_1604,N_1266,N_1133);
nand U1605 (N_1605,N_1321,N_1378);
nor U1606 (N_1606,N_1452,N_1093);
nor U1607 (N_1607,N_1002,N_1239);
nor U1608 (N_1608,N_1448,N_1310);
or U1609 (N_1609,N_1411,N_1086);
xor U1610 (N_1610,N_1074,N_1344);
and U1611 (N_1611,N_1409,N_1444);
and U1612 (N_1612,N_1262,N_1490);
nor U1613 (N_1613,N_1102,N_1208);
or U1614 (N_1614,N_1387,N_1147);
nand U1615 (N_1615,N_1154,N_1432);
nand U1616 (N_1616,N_1236,N_1470);
xnor U1617 (N_1617,N_1467,N_1421);
nand U1618 (N_1618,N_1067,N_1047);
xnor U1619 (N_1619,N_1416,N_1149);
or U1620 (N_1620,N_1351,N_1498);
nand U1621 (N_1621,N_1440,N_1305);
nor U1622 (N_1622,N_1477,N_1135);
nor U1623 (N_1623,N_1342,N_1264);
nor U1624 (N_1624,N_1260,N_1106);
nand U1625 (N_1625,N_1044,N_1200);
nor U1626 (N_1626,N_1284,N_1388);
nor U1627 (N_1627,N_1308,N_1403);
nand U1628 (N_1628,N_1144,N_1486);
xnor U1629 (N_1629,N_1380,N_1158);
and U1630 (N_1630,N_1318,N_1487);
nand U1631 (N_1631,N_1463,N_1205);
nor U1632 (N_1632,N_1049,N_1265);
xnor U1633 (N_1633,N_1025,N_1191);
nor U1634 (N_1634,N_1473,N_1155);
and U1635 (N_1635,N_1386,N_1249);
nand U1636 (N_1636,N_1227,N_1484);
nor U1637 (N_1637,N_1131,N_1237);
and U1638 (N_1638,N_1097,N_1210);
and U1639 (N_1639,N_1309,N_1212);
or U1640 (N_1640,N_1349,N_1059);
and U1641 (N_1641,N_1126,N_1184);
and U1642 (N_1642,N_1370,N_1030);
nor U1643 (N_1643,N_1474,N_1222);
nor U1644 (N_1644,N_1022,N_1009);
and U1645 (N_1645,N_1425,N_1492);
nor U1646 (N_1646,N_1050,N_1480);
and U1647 (N_1647,N_1103,N_1011);
xnor U1648 (N_1648,N_1313,N_1232);
and U1649 (N_1649,N_1229,N_1488);
nand U1650 (N_1650,N_1129,N_1141);
nand U1651 (N_1651,N_1314,N_1475);
nand U1652 (N_1652,N_1405,N_1345);
nand U1653 (N_1653,N_1118,N_1352);
or U1654 (N_1654,N_1446,N_1270);
and U1655 (N_1655,N_1132,N_1245);
nand U1656 (N_1656,N_1150,N_1325);
xor U1657 (N_1657,N_1163,N_1180);
or U1658 (N_1658,N_1121,N_1250);
xor U1659 (N_1659,N_1253,N_1257);
xnor U1660 (N_1660,N_1384,N_1311);
xor U1661 (N_1661,N_1242,N_1058);
nor U1662 (N_1662,N_1004,N_1109);
nand U1663 (N_1663,N_1445,N_1252);
nor U1664 (N_1664,N_1431,N_1274);
or U1665 (N_1665,N_1355,N_1286);
or U1666 (N_1666,N_1427,N_1334);
and U1667 (N_1667,N_1481,N_1117);
nor U1668 (N_1668,N_1124,N_1153);
xor U1669 (N_1669,N_1438,N_1413);
and U1670 (N_1670,N_1096,N_1437);
and U1671 (N_1671,N_1389,N_1493);
nand U1672 (N_1672,N_1434,N_1087);
nor U1673 (N_1673,N_1357,N_1248);
nor U1674 (N_1674,N_1272,N_1251);
and U1675 (N_1675,N_1207,N_1148);
and U1676 (N_1676,N_1057,N_1346);
nor U1677 (N_1677,N_1426,N_1041);
nand U1678 (N_1678,N_1295,N_1402);
nand U1679 (N_1679,N_1098,N_1307);
xnor U1680 (N_1680,N_1053,N_1333);
xnor U1681 (N_1681,N_1088,N_1169);
xor U1682 (N_1682,N_1006,N_1123);
nand U1683 (N_1683,N_1454,N_1258);
nor U1684 (N_1684,N_1415,N_1223);
nand U1685 (N_1685,N_1379,N_1417);
xnor U1686 (N_1686,N_1101,N_1085);
and U1687 (N_1687,N_1052,N_1156);
nor U1688 (N_1688,N_1179,N_1303);
and U1689 (N_1689,N_1450,N_1383);
or U1690 (N_1690,N_1130,N_1190);
and U1691 (N_1691,N_1151,N_1297);
nand U1692 (N_1692,N_1329,N_1186);
and U1693 (N_1693,N_1108,N_1070);
or U1694 (N_1694,N_1332,N_1398);
nor U1695 (N_1695,N_1166,N_1476);
xnor U1696 (N_1696,N_1288,N_1040);
and U1697 (N_1697,N_1368,N_1181);
xor U1698 (N_1698,N_1080,N_1164);
and U1699 (N_1699,N_1034,N_1068);
nand U1700 (N_1700,N_1392,N_1094);
and U1701 (N_1701,N_1451,N_1075);
or U1702 (N_1702,N_1362,N_1489);
or U1703 (N_1703,N_1433,N_1021);
or U1704 (N_1704,N_1268,N_1299);
nor U1705 (N_1705,N_1424,N_1472);
nand U1706 (N_1706,N_1447,N_1340);
nor U1707 (N_1707,N_1478,N_1221);
and U1708 (N_1708,N_1161,N_1401);
or U1709 (N_1709,N_1160,N_1037);
and U1710 (N_1710,N_1276,N_1324);
xor U1711 (N_1711,N_1019,N_1035);
or U1712 (N_1712,N_1320,N_1381);
nand U1713 (N_1713,N_1188,N_1328);
nor U1714 (N_1714,N_1289,N_1273);
nor U1715 (N_1715,N_1443,N_1348);
and U1716 (N_1716,N_1182,N_1326);
nand U1717 (N_1717,N_1048,N_1327);
nand U1718 (N_1718,N_1137,N_1111);
xnor U1719 (N_1719,N_1240,N_1127);
and U1720 (N_1720,N_1051,N_1255);
or U1721 (N_1721,N_1029,N_1354);
xor U1722 (N_1722,N_1065,N_1238);
xnor U1723 (N_1723,N_1196,N_1062);
nand U1724 (N_1724,N_1428,N_1376);
xor U1725 (N_1725,N_1363,N_1125);
and U1726 (N_1726,N_1122,N_1377);
nand U1727 (N_1727,N_1296,N_1012);
or U1728 (N_1728,N_1343,N_1174);
and U1729 (N_1729,N_1367,N_1060);
or U1730 (N_1730,N_1001,N_1136);
nand U1731 (N_1731,N_1495,N_1395);
nand U1732 (N_1732,N_1064,N_1089);
nand U1733 (N_1733,N_1176,N_1335);
nor U1734 (N_1734,N_1356,N_1275);
and U1735 (N_1735,N_1055,N_1178);
nand U1736 (N_1736,N_1092,N_1170);
or U1737 (N_1737,N_1466,N_1114);
nand U1738 (N_1738,N_1312,N_1406);
or U1739 (N_1739,N_1081,N_1241);
nor U1740 (N_1740,N_1436,N_1231);
xor U1741 (N_1741,N_1461,N_1267);
nand U1742 (N_1742,N_1420,N_1209);
nand U1743 (N_1743,N_1456,N_1418);
xnor U1744 (N_1744,N_1485,N_1358);
nand U1745 (N_1745,N_1084,N_1366);
xnor U1746 (N_1746,N_1396,N_1382);
nor U1747 (N_1747,N_1449,N_1410);
or U1748 (N_1748,N_1336,N_1423);
and U1749 (N_1749,N_1331,N_1496);
xor U1750 (N_1750,N_1436,N_1093);
nor U1751 (N_1751,N_1404,N_1305);
nand U1752 (N_1752,N_1176,N_1458);
nand U1753 (N_1753,N_1490,N_1396);
nand U1754 (N_1754,N_1434,N_1449);
or U1755 (N_1755,N_1271,N_1066);
nor U1756 (N_1756,N_1184,N_1121);
xor U1757 (N_1757,N_1031,N_1087);
nor U1758 (N_1758,N_1455,N_1143);
nand U1759 (N_1759,N_1403,N_1139);
nor U1760 (N_1760,N_1401,N_1187);
and U1761 (N_1761,N_1471,N_1406);
nor U1762 (N_1762,N_1010,N_1346);
nor U1763 (N_1763,N_1114,N_1051);
nand U1764 (N_1764,N_1131,N_1005);
and U1765 (N_1765,N_1207,N_1177);
and U1766 (N_1766,N_1217,N_1341);
or U1767 (N_1767,N_1034,N_1232);
and U1768 (N_1768,N_1403,N_1011);
nor U1769 (N_1769,N_1109,N_1369);
nand U1770 (N_1770,N_1487,N_1353);
nor U1771 (N_1771,N_1298,N_1065);
nand U1772 (N_1772,N_1387,N_1117);
or U1773 (N_1773,N_1227,N_1091);
xor U1774 (N_1774,N_1431,N_1282);
and U1775 (N_1775,N_1498,N_1106);
xor U1776 (N_1776,N_1357,N_1258);
nand U1777 (N_1777,N_1148,N_1471);
or U1778 (N_1778,N_1074,N_1027);
and U1779 (N_1779,N_1301,N_1420);
nand U1780 (N_1780,N_1099,N_1023);
nand U1781 (N_1781,N_1144,N_1291);
nor U1782 (N_1782,N_1018,N_1196);
nor U1783 (N_1783,N_1387,N_1139);
nand U1784 (N_1784,N_1029,N_1240);
nand U1785 (N_1785,N_1234,N_1162);
xor U1786 (N_1786,N_1322,N_1469);
nand U1787 (N_1787,N_1104,N_1178);
nor U1788 (N_1788,N_1326,N_1003);
nand U1789 (N_1789,N_1465,N_1088);
nand U1790 (N_1790,N_1253,N_1052);
nor U1791 (N_1791,N_1453,N_1444);
and U1792 (N_1792,N_1348,N_1341);
or U1793 (N_1793,N_1471,N_1001);
and U1794 (N_1794,N_1361,N_1469);
or U1795 (N_1795,N_1236,N_1490);
xnor U1796 (N_1796,N_1432,N_1169);
or U1797 (N_1797,N_1017,N_1038);
and U1798 (N_1798,N_1182,N_1141);
or U1799 (N_1799,N_1334,N_1264);
nand U1800 (N_1800,N_1169,N_1240);
nor U1801 (N_1801,N_1057,N_1117);
xnor U1802 (N_1802,N_1248,N_1464);
or U1803 (N_1803,N_1225,N_1289);
nor U1804 (N_1804,N_1433,N_1324);
nor U1805 (N_1805,N_1194,N_1163);
and U1806 (N_1806,N_1394,N_1323);
nor U1807 (N_1807,N_1105,N_1481);
and U1808 (N_1808,N_1223,N_1224);
nand U1809 (N_1809,N_1184,N_1026);
xnor U1810 (N_1810,N_1099,N_1168);
nand U1811 (N_1811,N_1390,N_1164);
and U1812 (N_1812,N_1181,N_1021);
nor U1813 (N_1813,N_1069,N_1126);
and U1814 (N_1814,N_1389,N_1423);
nand U1815 (N_1815,N_1356,N_1063);
nand U1816 (N_1816,N_1013,N_1462);
and U1817 (N_1817,N_1059,N_1271);
nand U1818 (N_1818,N_1119,N_1310);
or U1819 (N_1819,N_1392,N_1491);
xnor U1820 (N_1820,N_1390,N_1346);
and U1821 (N_1821,N_1065,N_1240);
and U1822 (N_1822,N_1204,N_1468);
and U1823 (N_1823,N_1494,N_1483);
or U1824 (N_1824,N_1251,N_1404);
nand U1825 (N_1825,N_1134,N_1160);
and U1826 (N_1826,N_1386,N_1333);
xor U1827 (N_1827,N_1140,N_1241);
nor U1828 (N_1828,N_1446,N_1491);
and U1829 (N_1829,N_1416,N_1199);
xor U1830 (N_1830,N_1177,N_1362);
and U1831 (N_1831,N_1441,N_1062);
or U1832 (N_1832,N_1243,N_1044);
nor U1833 (N_1833,N_1438,N_1237);
nor U1834 (N_1834,N_1414,N_1312);
and U1835 (N_1835,N_1384,N_1163);
nand U1836 (N_1836,N_1048,N_1007);
or U1837 (N_1837,N_1251,N_1484);
nand U1838 (N_1838,N_1154,N_1362);
xnor U1839 (N_1839,N_1332,N_1248);
xor U1840 (N_1840,N_1366,N_1483);
nand U1841 (N_1841,N_1145,N_1080);
nand U1842 (N_1842,N_1063,N_1115);
or U1843 (N_1843,N_1005,N_1188);
or U1844 (N_1844,N_1173,N_1365);
xor U1845 (N_1845,N_1085,N_1113);
and U1846 (N_1846,N_1299,N_1043);
xnor U1847 (N_1847,N_1169,N_1118);
or U1848 (N_1848,N_1133,N_1433);
and U1849 (N_1849,N_1087,N_1452);
and U1850 (N_1850,N_1213,N_1443);
nor U1851 (N_1851,N_1329,N_1059);
and U1852 (N_1852,N_1330,N_1252);
xnor U1853 (N_1853,N_1390,N_1458);
or U1854 (N_1854,N_1185,N_1244);
nor U1855 (N_1855,N_1348,N_1257);
or U1856 (N_1856,N_1231,N_1113);
or U1857 (N_1857,N_1350,N_1141);
or U1858 (N_1858,N_1034,N_1400);
and U1859 (N_1859,N_1422,N_1415);
or U1860 (N_1860,N_1361,N_1197);
and U1861 (N_1861,N_1057,N_1378);
xor U1862 (N_1862,N_1185,N_1466);
or U1863 (N_1863,N_1460,N_1396);
xnor U1864 (N_1864,N_1167,N_1236);
xnor U1865 (N_1865,N_1497,N_1175);
nor U1866 (N_1866,N_1343,N_1378);
nand U1867 (N_1867,N_1223,N_1484);
or U1868 (N_1868,N_1257,N_1447);
and U1869 (N_1869,N_1227,N_1426);
or U1870 (N_1870,N_1156,N_1451);
nand U1871 (N_1871,N_1433,N_1017);
or U1872 (N_1872,N_1067,N_1465);
or U1873 (N_1873,N_1191,N_1248);
or U1874 (N_1874,N_1224,N_1418);
nand U1875 (N_1875,N_1377,N_1029);
xor U1876 (N_1876,N_1287,N_1355);
or U1877 (N_1877,N_1141,N_1069);
nor U1878 (N_1878,N_1020,N_1027);
xor U1879 (N_1879,N_1084,N_1133);
or U1880 (N_1880,N_1024,N_1007);
xor U1881 (N_1881,N_1006,N_1141);
and U1882 (N_1882,N_1129,N_1373);
nor U1883 (N_1883,N_1072,N_1124);
nand U1884 (N_1884,N_1029,N_1203);
xor U1885 (N_1885,N_1360,N_1060);
and U1886 (N_1886,N_1061,N_1160);
or U1887 (N_1887,N_1291,N_1135);
nand U1888 (N_1888,N_1258,N_1409);
nand U1889 (N_1889,N_1408,N_1066);
or U1890 (N_1890,N_1179,N_1289);
nand U1891 (N_1891,N_1169,N_1008);
nand U1892 (N_1892,N_1002,N_1159);
nand U1893 (N_1893,N_1205,N_1008);
nand U1894 (N_1894,N_1053,N_1473);
nor U1895 (N_1895,N_1253,N_1273);
and U1896 (N_1896,N_1152,N_1276);
and U1897 (N_1897,N_1486,N_1155);
xor U1898 (N_1898,N_1342,N_1272);
or U1899 (N_1899,N_1243,N_1085);
nor U1900 (N_1900,N_1035,N_1253);
or U1901 (N_1901,N_1058,N_1231);
and U1902 (N_1902,N_1414,N_1015);
nor U1903 (N_1903,N_1420,N_1491);
nor U1904 (N_1904,N_1417,N_1168);
nand U1905 (N_1905,N_1357,N_1090);
nor U1906 (N_1906,N_1400,N_1051);
nand U1907 (N_1907,N_1090,N_1331);
and U1908 (N_1908,N_1024,N_1452);
or U1909 (N_1909,N_1051,N_1005);
and U1910 (N_1910,N_1123,N_1423);
nand U1911 (N_1911,N_1391,N_1226);
nand U1912 (N_1912,N_1464,N_1202);
and U1913 (N_1913,N_1312,N_1103);
and U1914 (N_1914,N_1321,N_1009);
and U1915 (N_1915,N_1217,N_1385);
or U1916 (N_1916,N_1374,N_1350);
and U1917 (N_1917,N_1472,N_1018);
nor U1918 (N_1918,N_1437,N_1441);
xor U1919 (N_1919,N_1303,N_1050);
nand U1920 (N_1920,N_1205,N_1200);
xor U1921 (N_1921,N_1141,N_1274);
xnor U1922 (N_1922,N_1251,N_1057);
or U1923 (N_1923,N_1183,N_1478);
or U1924 (N_1924,N_1013,N_1223);
or U1925 (N_1925,N_1477,N_1125);
or U1926 (N_1926,N_1443,N_1166);
nand U1927 (N_1927,N_1375,N_1302);
nand U1928 (N_1928,N_1360,N_1196);
nand U1929 (N_1929,N_1021,N_1224);
nand U1930 (N_1930,N_1358,N_1354);
nor U1931 (N_1931,N_1113,N_1239);
or U1932 (N_1932,N_1314,N_1019);
nor U1933 (N_1933,N_1205,N_1346);
nor U1934 (N_1934,N_1295,N_1160);
xnor U1935 (N_1935,N_1448,N_1100);
nand U1936 (N_1936,N_1114,N_1475);
nor U1937 (N_1937,N_1396,N_1165);
and U1938 (N_1938,N_1194,N_1181);
xor U1939 (N_1939,N_1100,N_1151);
or U1940 (N_1940,N_1213,N_1066);
xnor U1941 (N_1941,N_1456,N_1490);
nand U1942 (N_1942,N_1098,N_1426);
nand U1943 (N_1943,N_1311,N_1342);
xnor U1944 (N_1944,N_1479,N_1281);
nand U1945 (N_1945,N_1301,N_1191);
xor U1946 (N_1946,N_1137,N_1333);
nor U1947 (N_1947,N_1231,N_1483);
and U1948 (N_1948,N_1327,N_1272);
nand U1949 (N_1949,N_1044,N_1469);
nor U1950 (N_1950,N_1305,N_1150);
nand U1951 (N_1951,N_1090,N_1125);
xor U1952 (N_1952,N_1023,N_1313);
nor U1953 (N_1953,N_1475,N_1216);
or U1954 (N_1954,N_1151,N_1189);
nand U1955 (N_1955,N_1176,N_1216);
xnor U1956 (N_1956,N_1305,N_1387);
nand U1957 (N_1957,N_1408,N_1418);
or U1958 (N_1958,N_1226,N_1049);
nand U1959 (N_1959,N_1404,N_1209);
nand U1960 (N_1960,N_1149,N_1054);
xor U1961 (N_1961,N_1223,N_1377);
xnor U1962 (N_1962,N_1320,N_1353);
and U1963 (N_1963,N_1191,N_1348);
nor U1964 (N_1964,N_1010,N_1191);
xor U1965 (N_1965,N_1076,N_1349);
nand U1966 (N_1966,N_1113,N_1017);
or U1967 (N_1967,N_1058,N_1205);
xor U1968 (N_1968,N_1350,N_1359);
nand U1969 (N_1969,N_1101,N_1347);
xor U1970 (N_1970,N_1023,N_1251);
nor U1971 (N_1971,N_1464,N_1145);
and U1972 (N_1972,N_1015,N_1405);
or U1973 (N_1973,N_1227,N_1293);
xor U1974 (N_1974,N_1460,N_1487);
nand U1975 (N_1975,N_1402,N_1290);
nor U1976 (N_1976,N_1336,N_1117);
nand U1977 (N_1977,N_1415,N_1385);
xor U1978 (N_1978,N_1194,N_1106);
nand U1979 (N_1979,N_1498,N_1307);
nand U1980 (N_1980,N_1093,N_1108);
nor U1981 (N_1981,N_1000,N_1313);
xor U1982 (N_1982,N_1373,N_1069);
or U1983 (N_1983,N_1427,N_1165);
nand U1984 (N_1984,N_1474,N_1457);
or U1985 (N_1985,N_1202,N_1231);
nand U1986 (N_1986,N_1019,N_1444);
nand U1987 (N_1987,N_1217,N_1286);
xnor U1988 (N_1988,N_1434,N_1148);
xor U1989 (N_1989,N_1365,N_1363);
or U1990 (N_1990,N_1443,N_1180);
or U1991 (N_1991,N_1165,N_1177);
nand U1992 (N_1992,N_1277,N_1059);
nor U1993 (N_1993,N_1079,N_1280);
nor U1994 (N_1994,N_1197,N_1113);
nor U1995 (N_1995,N_1220,N_1227);
nand U1996 (N_1996,N_1382,N_1418);
and U1997 (N_1997,N_1436,N_1363);
nor U1998 (N_1998,N_1010,N_1477);
xnor U1999 (N_1999,N_1103,N_1110);
xor U2000 (N_2000,N_1925,N_1613);
xnor U2001 (N_2001,N_1568,N_1816);
nor U2002 (N_2002,N_1625,N_1840);
or U2003 (N_2003,N_1602,N_1616);
and U2004 (N_2004,N_1888,N_1710);
nor U2005 (N_2005,N_1525,N_1776);
nand U2006 (N_2006,N_1974,N_1968);
xnor U2007 (N_2007,N_1993,N_1695);
xnor U2008 (N_2008,N_1886,N_1813);
nor U2009 (N_2009,N_1735,N_1846);
nor U2010 (N_2010,N_1637,N_1989);
nor U2011 (N_2011,N_1782,N_1608);
nand U2012 (N_2012,N_1933,N_1825);
and U2013 (N_2013,N_1644,N_1648);
and U2014 (N_2014,N_1547,N_1551);
nand U2015 (N_2015,N_1538,N_1550);
and U2016 (N_2016,N_1949,N_1716);
or U2017 (N_2017,N_1717,N_1959);
nand U2018 (N_2018,N_1666,N_1961);
and U2019 (N_2019,N_1722,N_1788);
or U2020 (N_2020,N_1733,N_1509);
nand U2021 (N_2021,N_1573,N_1867);
nand U2022 (N_2022,N_1820,N_1905);
or U2023 (N_2023,N_1859,N_1750);
nand U2024 (N_2024,N_1576,N_1789);
xor U2025 (N_2025,N_1896,N_1621);
nor U2026 (N_2026,N_1661,N_1752);
and U2027 (N_2027,N_1996,N_1786);
or U2028 (N_2028,N_1600,N_1708);
xor U2029 (N_2029,N_1712,N_1690);
or U2030 (N_2030,N_1811,N_1552);
nand U2031 (N_2031,N_1895,N_1909);
or U2032 (N_2032,N_1502,N_1998);
and U2033 (N_2033,N_1728,N_1580);
nand U2034 (N_2034,N_1595,N_1609);
nand U2035 (N_2035,N_1512,N_1983);
or U2036 (N_2036,N_1734,N_1913);
nand U2037 (N_2037,N_1622,N_1539);
nand U2038 (N_2038,N_1962,N_1907);
nor U2039 (N_2039,N_1588,N_1884);
nand U2040 (N_2040,N_1534,N_1848);
or U2041 (N_2041,N_1599,N_1639);
xnor U2042 (N_2042,N_1725,N_1723);
and U2043 (N_2043,N_1957,N_1770);
xnor U2044 (N_2044,N_1756,N_1947);
or U2045 (N_2045,N_1822,N_1563);
nor U2046 (N_2046,N_1633,N_1543);
nand U2047 (N_2047,N_1901,N_1745);
xnor U2048 (N_2048,N_1932,N_1624);
nand U2049 (N_2049,N_1900,N_1919);
or U2050 (N_2050,N_1743,N_1650);
xor U2051 (N_2051,N_1673,N_1596);
nor U2052 (N_2052,N_1986,N_1781);
xnor U2053 (N_2053,N_1829,N_1706);
nand U2054 (N_2054,N_1652,N_1686);
nand U2055 (N_2055,N_1977,N_1808);
or U2056 (N_2056,N_1631,N_1852);
and U2057 (N_2057,N_1724,N_1775);
or U2058 (N_2058,N_1773,N_1793);
nand U2059 (N_2059,N_1649,N_1641);
xor U2060 (N_2060,N_1700,N_1975);
nor U2061 (N_2061,N_1893,N_1954);
and U2062 (N_2062,N_1918,N_1851);
and U2063 (N_2063,N_1567,N_1948);
and U2064 (N_2064,N_1601,N_1774);
nor U2065 (N_2065,N_1861,N_1713);
xnor U2066 (N_2066,N_1562,N_1772);
or U2067 (N_2067,N_1916,N_1777);
xor U2068 (N_2068,N_1912,N_1730);
or U2069 (N_2069,N_1967,N_1855);
xor U2070 (N_2070,N_1844,N_1979);
nand U2071 (N_2071,N_1672,N_1583);
or U2072 (N_2072,N_1603,N_1703);
xnor U2073 (N_2073,N_1529,N_1956);
nand U2074 (N_2074,N_1934,N_1875);
and U2075 (N_2075,N_1768,N_1759);
nand U2076 (N_2076,N_1620,N_1535);
xnor U2077 (N_2077,N_1513,N_1879);
nor U2078 (N_2078,N_1647,N_1541);
xor U2079 (N_2079,N_1718,N_1950);
nand U2080 (N_2080,N_1507,N_1936);
nor U2081 (N_2081,N_1678,N_1565);
nor U2082 (N_2082,N_1809,N_1584);
or U2083 (N_2083,N_1553,N_1696);
nor U2084 (N_2084,N_1737,N_1658);
or U2085 (N_2085,N_1878,N_1744);
and U2086 (N_2086,N_1662,N_1917);
xor U2087 (N_2087,N_1854,N_1812);
nor U2088 (N_2088,N_1510,N_1575);
or U2089 (N_2089,N_1694,N_1924);
nor U2090 (N_2090,N_1794,N_1972);
and U2091 (N_2091,N_1942,N_1570);
or U2092 (N_2092,N_1693,N_1530);
or U2093 (N_2093,N_1902,N_1869);
nor U2094 (N_2094,N_1978,N_1528);
xnor U2095 (N_2095,N_1532,N_1747);
nor U2096 (N_2096,N_1832,N_1892);
and U2097 (N_2097,N_1691,N_1798);
or U2098 (N_2098,N_1640,N_1858);
nand U2099 (N_2099,N_1517,N_1864);
nand U2100 (N_2100,N_1629,N_1843);
and U2101 (N_2101,N_1610,N_1739);
or U2102 (N_2102,N_1771,N_1515);
nand U2103 (N_2103,N_1623,N_1762);
nand U2104 (N_2104,N_1542,N_1738);
nand U2105 (N_2105,N_1800,N_1540);
nor U2106 (N_2106,N_1699,N_1757);
nor U2107 (N_2107,N_1780,N_1741);
or U2108 (N_2108,N_1654,N_1577);
nor U2109 (N_2109,N_1849,N_1635);
or U2110 (N_2110,N_1943,N_1559);
xor U2111 (N_2111,N_1819,N_1638);
and U2112 (N_2112,N_1958,N_1589);
nand U2113 (N_2113,N_1945,N_1676);
xor U2114 (N_2114,N_1834,N_1830);
or U2115 (N_2115,N_1862,N_1585);
nor U2116 (N_2116,N_1536,N_1561);
xnor U2117 (N_2117,N_1802,N_1668);
nor U2118 (N_2118,N_1898,N_1882);
nor U2119 (N_2119,N_1702,N_1579);
xor U2120 (N_2120,N_1597,N_1779);
and U2121 (N_2121,N_1921,N_1765);
nand U2122 (N_2122,N_1874,N_1522);
nand U2123 (N_2123,N_1763,N_1985);
nor U2124 (N_2124,N_1594,N_1806);
nand U2125 (N_2125,N_1791,N_1796);
and U2126 (N_2126,N_1749,N_1894);
or U2127 (N_2127,N_1951,N_1500);
xor U2128 (N_2128,N_1887,N_1731);
nand U2129 (N_2129,N_1607,N_1824);
nor U2130 (N_2130,N_1646,N_1904);
and U2131 (N_2131,N_1938,N_1685);
or U2132 (N_2132,N_1946,N_1684);
nand U2133 (N_2133,N_1995,N_1508);
and U2134 (N_2134,N_1593,N_1870);
or U2135 (N_2135,N_1994,N_1598);
nand U2136 (N_2136,N_1838,N_1628);
nor U2137 (N_2137,N_1922,N_1660);
nand U2138 (N_2138,N_1758,N_1826);
nand U2139 (N_2139,N_1842,N_1836);
nor U2140 (N_2140,N_1908,N_1634);
or U2141 (N_2141,N_1677,N_1885);
xnor U2142 (N_2142,N_1714,N_1755);
xor U2143 (N_2143,N_1665,N_1671);
xor U2144 (N_2144,N_1555,N_1564);
xnor U2145 (N_2145,N_1980,N_1619);
or U2146 (N_2146,N_1963,N_1630);
nand U2147 (N_2147,N_1581,N_1784);
or U2148 (N_2148,N_1973,N_1911);
nand U2149 (N_2149,N_1939,N_1632);
nand U2150 (N_2150,N_1732,N_1805);
xor U2151 (N_2151,N_1729,N_1627);
or U2152 (N_2152,N_1503,N_1823);
and U2153 (N_2153,N_1997,N_1828);
xor U2154 (N_2154,N_1523,N_1545);
or U2155 (N_2155,N_1860,N_1531);
or U2156 (N_2156,N_1674,N_1767);
or U2157 (N_2157,N_1516,N_1653);
or U2158 (N_2158,N_1636,N_1518);
and U2159 (N_2159,N_1866,N_1655);
xnor U2160 (N_2160,N_1711,N_1664);
xnor U2161 (N_2161,N_1971,N_1548);
and U2162 (N_2162,N_1814,N_1792);
and U2163 (N_2163,N_1651,N_1833);
and U2164 (N_2164,N_1872,N_1574);
or U2165 (N_2165,N_1719,N_1520);
nand U2166 (N_2166,N_1537,N_1856);
and U2167 (N_2167,N_1992,N_1558);
nand U2168 (N_2168,N_1604,N_1546);
nand U2169 (N_2169,N_1982,N_1835);
or U2170 (N_2170,N_1766,N_1605);
and U2171 (N_2171,N_1906,N_1783);
nand U2172 (N_2172,N_1929,N_1586);
or U2173 (N_2173,N_1795,N_1505);
nor U2174 (N_2174,N_1871,N_1821);
nor U2175 (N_2175,N_1940,N_1847);
or U2176 (N_2176,N_1850,N_1964);
and U2177 (N_2177,N_1790,N_1560);
nand U2178 (N_2178,N_1764,N_1663);
nor U2179 (N_2179,N_1999,N_1506);
and U2180 (N_2180,N_1720,N_1591);
nor U2181 (N_2181,N_1659,N_1556);
nand U2182 (N_2182,N_1526,N_1587);
nor U2183 (N_2183,N_1751,N_1903);
and U2184 (N_2184,N_1797,N_1923);
and U2185 (N_2185,N_1927,N_1746);
and U2186 (N_2186,N_1953,N_1504);
or U2187 (N_2187,N_1910,N_1952);
and U2188 (N_2188,N_1827,N_1914);
nor U2189 (N_2189,N_1928,N_1801);
nand U2190 (N_2190,N_1873,N_1617);
or U2191 (N_2191,N_1692,N_1645);
xor U2192 (N_2192,N_1527,N_1667);
xnor U2193 (N_2193,N_1804,N_1753);
xor U2194 (N_2194,N_1606,N_1614);
and U2195 (N_2195,N_1987,N_1742);
xor U2196 (N_2196,N_1981,N_1853);
xor U2197 (N_2197,N_1626,N_1698);
and U2198 (N_2198,N_1721,N_1960);
and U2199 (N_2199,N_1704,N_1857);
nor U2200 (N_2200,N_1841,N_1931);
nor U2201 (N_2201,N_1937,N_1831);
or U2202 (N_2202,N_1524,N_1807);
and U2203 (N_2203,N_1955,N_1889);
nand U2204 (N_2204,N_1803,N_1760);
nand U2205 (N_2205,N_1761,N_1839);
nand U2206 (N_2206,N_1754,N_1683);
or U2207 (N_2207,N_1680,N_1817);
and U2208 (N_2208,N_1521,N_1554);
nor U2209 (N_2209,N_1920,N_1881);
xnor U2210 (N_2210,N_1566,N_1578);
or U2211 (N_2211,N_1709,N_1787);
nor U2212 (N_2212,N_1689,N_1736);
or U2213 (N_2213,N_1815,N_1615);
nor U2214 (N_2214,N_1681,N_1514);
xor U2215 (N_2215,N_1880,N_1966);
xnor U2216 (N_2216,N_1557,N_1670);
nand U2217 (N_2217,N_1687,N_1890);
or U2218 (N_2218,N_1590,N_1915);
and U2219 (N_2219,N_1544,N_1656);
xnor U2220 (N_2220,N_1675,N_1533);
xnor U2221 (N_2221,N_1643,N_1969);
nand U2222 (N_2222,N_1810,N_1642);
xor U2223 (N_2223,N_1818,N_1705);
nor U2224 (N_2224,N_1863,N_1941);
and U2225 (N_2225,N_1549,N_1868);
xnor U2226 (N_2226,N_1519,N_1592);
or U2227 (N_2227,N_1740,N_1727);
or U2228 (N_2228,N_1865,N_1679);
nand U2229 (N_2229,N_1688,N_1891);
xnor U2230 (N_2230,N_1769,N_1926);
nor U2231 (N_2231,N_1612,N_1707);
nor U2232 (N_2232,N_1582,N_1572);
nand U2233 (N_2233,N_1697,N_1991);
or U2234 (N_2234,N_1976,N_1984);
nor U2235 (N_2235,N_1930,N_1715);
or U2236 (N_2236,N_1799,N_1944);
nand U2237 (N_2237,N_1845,N_1748);
nor U2238 (N_2238,N_1837,N_1611);
or U2239 (N_2239,N_1569,N_1657);
nor U2240 (N_2240,N_1571,N_1988);
nand U2241 (N_2241,N_1876,N_1970);
nand U2242 (N_2242,N_1669,N_1877);
and U2243 (N_2243,N_1785,N_1618);
xnor U2244 (N_2244,N_1501,N_1899);
nor U2245 (N_2245,N_1897,N_1965);
nand U2246 (N_2246,N_1511,N_1883);
nor U2247 (N_2247,N_1935,N_1778);
nand U2248 (N_2248,N_1726,N_1990);
nor U2249 (N_2249,N_1682,N_1701);
or U2250 (N_2250,N_1775,N_1730);
or U2251 (N_2251,N_1852,N_1742);
and U2252 (N_2252,N_1815,N_1622);
and U2253 (N_2253,N_1982,N_1605);
nor U2254 (N_2254,N_1589,N_1888);
nor U2255 (N_2255,N_1845,N_1551);
and U2256 (N_2256,N_1858,N_1866);
nor U2257 (N_2257,N_1523,N_1873);
xor U2258 (N_2258,N_1814,N_1640);
and U2259 (N_2259,N_1895,N_1879);
and U2260 (N_2260,N_1619,N_1503);
nand U2261 (N_2261,N_1547,N_1686);
or U2262 (N_2262,N_1726,N_1674);
xor U2263 (N_2263,N_1983,N_1558);
and U2264 (N_2264,N_1940,N_1955);
nor U2265 (N_2265,N_1994,N_1809);
and U2266 (N_2266,N_1531,N_1672);
nand U2267 (N_2267,N_1719,N_1752);
nor U2268 (N_2268,N_1891,N_1717);
xnor U2269 (N_2269,N_1804,N_1999);
or U2270 (N_2270,N_1881,N_1934);
or U2271 (N_2271,N_1990,N_1894);
xor U2272 (N_2272,N_1957,N_1523);
nor U2273 (N_2273,N_1853,N_1608);
nor U2274 (N_2274,N_1702,N_1694);
nand U2275 (N_2275,N_1707,N_1885);
and U2276 (N_2276,N_1630,N_1937);
nand U2277 (N_2277,N_1948,N_1831);
nor U2278 (N_2278,N_1714,N_1603);
nand U2279 (N_2279,N_1652,N_1684);
xnor U2280 (N_2280,N_1716,N_1539);
and U2281 (N_2281,N_1617,N_1877);
and U2282 (N_2282,N_1681,N_1555);
and U2283 (N_2283,N_1944,N_1724);
or U2284 (N_2284,N_1992,N_1956);
nand U2285 (N_2285,N_1641,N_1682);
nand U2286 (N_2286,N_1599,N_1767);
or U2287 (N_2287,N_1914,N_1865);
xnor U2288 (N_2288,N_1952,N_1552);
nand U2289 (N_2289,N_1835,N_1766);
and U2290 (N_2290,N_1637,N_1611);
nand U2291 (N_2291,N_1766,N_1646);
and U2292 (N_2292,N_1539,N_1791);
nand U2293 (N_2293,N_1727,N_1551);
nand U2294 (N_2294,N_1774,N_1542);
xor U2295 (N_2295,N_1657,N_1505);
xor U2296 (N_2296,N_1792,N_1828);
or U2297 (N_2297,N_1972,N_1645);
or U2298 (N_2298,N_1935,N_1618);
xor U2299 (N_2299,N_1605,N_1764);
or U2300 (N_2300,N_1585,N_1641);
or U2301 (N_2301,N_1837,N_1566);
nand U2302 (N_2302,N_1592,N_1619);
and U2303 (N_2303,N_1535,N_1692);
xor U2304 (N_2304,N_1581,N_1717);
nor U2305 (N_2305,N_1853,N_1923);
nor U2306 (N_2306,N_1789,N_1625);
nand U2307 (N_2307,N_1878,N_1711);
and U2308 (N_2308,N_1679,N_1665);
nand U2309 (N_2309,N_1870,N_1760);
nand U2310 (N_2310,N_1908,N_1892);
and U2311 (N_2311,N_1871,N_1646);
and U2312 (N_2312,N_1603,N_1724);
xor U2313 (N_2313,N_1967,N_1949);
xor U2314 (N_2314,N_1629,N_1979);
nor U2315 (N_2315,N_1512,N_1565);
xor U2316 (N_2316,N_1529,N_1843);
nor U2317 (N_2317,N_1882,N_1811);
nand U2318 (N_2318,N_1923,N_1920);
and U2319 (N_2319,N_1640,N_1831);
or U2320 (N_2320,N_1759,N_1554);
or U2321 (N_2321,N_1611,N_1871);
or U2322 (N_2322,N_1968,N_1506);
or U2323 (N_2323,N_1745,N_1948);
and U2324 (N_2324,N_1972,N_1639);
and U2325 (N_2325,N_1586,N_1766);
xnor U2326 (N_2326,N_1627,N_1988);
nand U2327 (N_2327,N_1682,N_1676);
nor U2328 (N_2328,N_1850,N_1974);
and U2329 (N_2329,N_1937,N_1985);
and U2330 (N_2330,N_1783,N_1682);
or U2331 (N_2331,N_1680,N_1826);
or U2332 (N_2332,N_1938,N_1930);
nor U2333 (N_2333,N_1596,N_1862);
or U2334 (N_2334,N_1777,N_1576);
nor U2335 (N_2335,N_1516,N_1666);
xor U2336 (N_2336,N_1848,N_1542);
or U2337 (N_2337,N_1571,N_1780);
xnor U2338 (N_2338,N_1686,N_1781);
and U2339 (N_2339,N_1763,N_1827);
nor U2340 (N_2340,N_1902,N_1642);
nor U2341 (N_2341,N_1701,N_1861);
or U2342 (N_2342,N_1544,N_1698);
xnor U2343 (N_2343,N_1817,N_1921);
nor U2344 (N_2344,N_1842,N_1662);
nor U2345 (N_2345,N_1768,N_1901);
nor U2346 (N_2346,N_1830,N_1558);
and U2347 (N_2347,N_1948,N_1687);
nor U2348 (N_2348,N_1835,N_1557);
xnor U2349 (N_2349,N_1645,N_1958);
nand U2350 (N_2350,N_1904,N_1853);
and U2351 (N_2351,N_1962,N_1544);
and U2352 (N_2352,N_1648,N_1959);
xor U2353 (N_2353,N_1889,N_1615);
nor U2354 (N_2354,N_1514,N_1968);
xnor U2355 (N_2355,N_1732,N_1839);
nand U2356 (N_2356,N_1763,N_1593);
or U2357 (N_2357,N_1781,N_1768);
and U2358 (N_2358,N_1860,N_1868);
and U2359 (N_2359,N_1619,N_1516);
nand U2360 (N_2360,N_1752,N_1538);
nand U2361 (N_2361,N_1721,N_1850);
nor U2362 (N_2362,N_1953,N_1583);
nor U2363 (N_2363,N_1829,N_1691);
xnor U2364 (N_2364,N_1695,N_1720);
xnor U2365 (N_2365,N_1842,N_1851);
nand U2366 (N_2366,N_1519,N_1517);
nand U2367 (N_2367,N_1521,N_1766);
nor U2368 (N_2368,N_1652,N_1888);
nand U2369 (N_2369,N_1507,N_1765);
nor U2370 (N_2370,N_1853,N_1605);
xnor U2371 (N_2371,N_1877,N_1874);
xor U2372 (N_2372,N_1597,N_1891);
nand U2373 (N_2373,N_1562,N_1524);
and U2374 (N_2374,N_1579,N_1699);
or U2375 (N_2375,N_1773,N_1807);
and U2376 (N_2376,N_1939,N_1727);
xnor U2377 (N_2377,N_1664,N_1962);
or U2378 (N_2378,N_1581,N_1708);
nor U2379 (N_2379,N_1658,N_1532);
nor U2380 (N_2380,N_1503,N_1590);
nor U2381 (N_2381,N_1955,N_1736);
xnor U2382 (N_2382,N_1827,N_1787);
nand U2383 (N_2383,N_1841,N_1855);
nand U2384 (N_2384,N_1529,N_1687);
or U2385 (N_2385,N_1570,N_1784);
nand U2386 (N_2386,N_1926,N_1777);
xnor U2387 (N_2387,N_1809,N_1654);
nand U2388 (N_2388,N_1991,N_1646);
xnor U2389 (N_2389,N_1976,N_1595);
or U2390 (N_2390,N_1707,N_1656);
nor U2391 (N_2391,N_1600,N_1919);
or U2392 (N_2392,N_1522,N_1811);
nand U2393 (N_2393,N_1517,N_1620);
nand U2394 (N_2394,N_1683,N_1795);
nor U2395 (N_2395,N_1728,N_1818);
nand U2396 (N_2396,N_1671,N_1870);
or U2397 (N_2397,N_1646,N_1730);
nor U2398 (N_2398,N_1955,N_1705);
or U2399 (N_2399,N_1532,N_1768);
nor U2400 (N_2400,N_1647,N_1805);
xor U2401 (N_2401,N_1757,N_1513);
nand U2402 (N_2402,N_1501,N_1520);
and U2403 (N_2403,N_1596,N_1603);
or U2404 (N_2404,N_1816,N_1991);
nand U2405 (N_2405,N_1925,N_1700);
nand U2406 (N_2406,N_1756,N_1633);
xnor U2407 (N_2407,N_1672,N_1955);
or U2408 (N_2408,N_1848,N_1932);
and U2409 (N_2409,N_1599,N_1641);
nand U2410 (N_2410,N_1625,N_1533);
and U2411 (N_2411,N_1964,N_1989);
and U2412 (N_2412,N_1827,N_1519);
nor U2413 (N_2413,N_1749,N_1773);
xnor U2414 (N_2414,N_1973,N_1859);
nor U2415 (N_2415,N_1711,N_1930);
or U2416 (N_2416,N_1804,N_1962);
or U2417 (N_2417,N_1938,N_1794);
nand U2418 (N_2418,N_1721,N_1869);
and U2419 (N_2419,N_1681,N_1799);
nor U2420 (N_2420,N_1728,N_1876);
or U2421 (N_2421,N_1882,N_1533);
and U2422 (N_2422,N_1848,N_1861);
nor U2423 (N_2423,N_1930,N_1885);
and U2424 (N_2424,N_1819,N_1573);
and U2425 (N_2425,N_1987,N_1663);
and U2426 (N_2426,N_1811,N_1701);
nor U2427 (N_2427,N_1738,N_1729);
nand U2428 (N_2428,N_1538,N_1938);
nand U2429 (N_2429,N_1890,N_1598);
nand U2430 (N_2430,N_1948,N_1909);
nand U2431 (N_2431,N_1891,N_1522);
and U2432 (N_2432,N_1921,N_1998);
nand U2433 (N_2433,N_1619,N_1751);
or U2434 (N_2434,N_1939,N_1677);
and U2435 (N_2435,N_1789,N_1857);
and U2436 (N_2436,N_1975,N_1758);
and U2437 (N_2437,N_1788,N_1525);
nand U2438 (N_2438,N_1924,N_1530);
nand U2439 (N_2439,N_1918,N_1802);
xor U2440 (N_2440,N_1597,N_1928);
nor U2441 (N_2441,N_1593,N_1740);
nor U2442 (N_2442,N_1629,N_1620);
nand U2443 (N_2443,N_1572,N_1600);
or U2444 (N_2444,N_1846,N_1525);
nor U2445 (N_2445,N_1950,N_1885);
nor U2446 (N_2446,N_1954,N_1905);
nor U2447 (N_2447,N_1699,N_1829);
and U2448 (N_2448,N_1562,N_1897);
nand U2449 (N_2449,N_1831,N_1527);
and U2450 (N_2450,N_1564,N_1728);
nor U2451 (N_2451,N_1928,N_1952);
xor U2452 (N_2452,N_1748,N_1673);
and U2453 (N_2453,N_1897,N_1507);
nand U2454 (N_2454,N_1814,N_1783);
and U2455 (N_2455,N_1525,N_1886);
nor U2456 (N_2456,N_1668,N_1855);
and U2457 (N_2457,N_1597,N_1842);
or U2458 (N_2458,N_1865,N_1661);
xor U2459 (N_2459,N_1863,N_1535);
nor U2460 (N_2460,N_1882,N_1951);
nor U2461 (N_2461,N_1925,N_1987);
xor U2462 (N_2462,N_1963,N_1960);
nand U2463 (N_2463,N_1584,N_1567);
nor U2464 (N_2464,N_1894,N_1836);
and U2465 (N_2465,N_1522,N_1929);
nor U2466 (N_2466,N_1588,N_1617);
nor U2467 (N_2467,N_1669,N_1774);
nand U2468 (N_2468,N_1613,N_1952);
nor U2469 (N_2469,N_1811,N_1574);
or U2470 (N_2470,N_1727,N_1875);
nand U2471 (N_2471,N_1889,N_1991);
and U2472 (N_2472,N_1841,N_1929);
nand U2473 (N_2473,N_1894,N_1679);
and U2474 (N_2474,N_1786,N_1839);
nand U2475 (N_2475,N_1509,N_1650);
xnor U2476 (N_2476,N_1919,N_1538);
nand U2477 (N_2477,N_1770,N_1786);
nand U2478 (N_2478,N_1579,N_1551);
and U2479 (N_2479,N_1750,N_1975);
nor U2480 (N_2480,N_1576,N_1843);
nor U2481 (N_2481,N_1848,N_1607);
xor U2482 (N_2482,N_1563,N_1805);
nand U2483 (N_2483,N_1939,N_1608);
nor U2484 (N_2484,N_1913,N_1639);
nand U2485 (N_2485,N_1548,N_1709);
nor U2486 (N_2486,N_1795,N_1684);
nor U2487 (N_2487,N_1531,N_1718);
and U2488 (N_2488,N_1624,N_1578);
or U2489 (N_2489,N_1883,N_1890);
and U2490 (N_2490,N_1652,N_1672);
or U2491 (N_2491,N_1824,N_1776);
and U2492 (N_2492,N_1771,N_1622);
and U2493 (N_2493,N_1646,N_1843);
or U2494 (N_2494,N_1745,N_1840);
xnor U2495 (N_2495,N_1609,N_1998);
or U2496 (N_2496,N_1815,N_1981);
nand U2497 (N_2497,N_1703,N_1901);
nand U2498 (N_2498,N_1542,N_1759);
nand U2499 (N_2499,N_1988,N_1827);
nand U2500 (N_2500,N_2414,N_2022);
and U2501 (N_2501,N_2427,N_2063);
nor U2502 (N_2502,N_2230,N_2431);
nor U2503 (N_2503,N_2157,N_2192);
nand U2504 (N_2504,N_2327,N_2398);
nand U2505 (N_2505,N_2301,N_2426);
nor U2506 (N_2506,N_2008,N_2288);
and U2507 (N_2507,N_2122,N_2121);
nand U2508 (N_2508,N_2281,N_2010);
or U2509 (N_2509,N_2170,N_2331);
and U2510 (N_2510,N_2056,N_2433);
or U2511 (N_2511,N_2064,N_2209);
or U2512 (N_2512,N_2393,N_2378);
and U2513 (N_2513,N_2241,N_2137);
nor U2514 (N_2514,N_2496,N_2035);
and U2515 (N_2515,N_2435,N_2268);
nor U2516 (N_2516,N_2345,N_2227);
nor U2517 (N_2517,N_2340,N_2462);
nand U2518 (N_2518,N_2445,N_2082);
nor U2519 (N_2519,N_2317,N_2114);
and U2520 (N_2520,N_2175,N_2286);
and U2521 (N_2521,N_2313,N_2015);
nand U2522 (N_2522,N_2150,N_2220);
xor U2523 (N_2523,N_2385,N_2436);
nand U2524 (N_2524,N_2441,N_2362);
and U2525 (N_2525,N_2029,N_2402);
and U2526 (N_2526,N_2389,N_2079);
xor U2527 (N_2527,N_2390,N_2388);
or U2528 (N_2528,N_2457,N_2172);
xnor U2529 (N_2529,N_2018,N_2471);
nor U2530 (N_2530,N_2005,N_2207);
or U2531 (N_2531,N_2463,N_2203);
and U2532 (N_2532,N_2120,N_2167);
or U2533 (N_2533,N_2208,N_2105);
and U2534 (N_2534,N_2376,N_2382);
xor U2535 (N_2535,N_2012,N_2131);
nand U2536 (N_2536,N_2284,N_2375);
and U2537 (N_2537,N_2406,N_2236);
nor U2538 (N_2538,N_2109,N_2159);
nor U2539 (N_2539,N_2239,N_2069);
nand U2540 (N_2540,N_2332,N_2279);
nor U2541 (N_2541,N_2196,N_2135);
and U2542 (N_2542,N_2380,N_2201);
and U2543 (N_2543,N_2271,N_2016);
or U2544 (N_2544,N_2118,N_2326);
nand U2545 (N_2545,N_2296,N_2106);
and U2546 (N_2546,N_2273,N_2335);
and U2547 (N_2547,N_2403,N_2358);
or U2548 (N_2548,N_2257,N_2229);
nor U2549 (N_2549,N_2161,N_2000);
or U2550 (N_2550,N_2495,N_2409);
nand U2551 (N_2551,N_2030,N_2184);
and U2552 (N_2552,N_2259,N_2142);
or U2553 (N_2553,N_2133,N_2071);
or U2554 (N_2554,N_2339,N_2193);
nand U2555 (N_2555,N_2162,N_2097);
or U2556 (N_2556,N_2085,N_2197);
nand U2557 (N_2557,N_2072,N_2421);
nor U2558 (N_2558,N_2488,N_2165);
nand U2559 (N_2559,N_2396,N_2434);
nor U2560 (N_2560,N_2334,N_2060);
and U2561 (N_2561,N_2026,N_2404);
or U2562 (N_2562,N_2101,N_2136);
nand U2563 (N_2563,N_2039,N_2231);
xnor U2564 (N_2564,N_2386,N_2492);
or U2565 (N_2565,N_2232,N_2074);
nor U2566 (N_2566,N_2164,N_2468);
nand U2567 (N_2567,N_2348,N_2399);
nand U2568 (N_2568,N_2212,N_2206);
nor U2569 (N_2569,N_2045,N_2202);
and U2570 (N_2570,N_2054,N_2213);
nor U2571 (N_2571,N_2081,N_2337);
and U2572 (N_2572,N_2077,N_2116);
and U2573 (N_2573,N_2475,N_2185);
nand U2574 (N_2574,N_2112,N_2473);
nor U2575 (N_2575,N_2467,N_2068);
and U2576 (N_2576,N_2065,N_2325);
and U2577 (N_2577,N_2117,N_2315);
nor U2578 (N_2578,N_2028,N_2311);
and U2579 (N_2579,N_2243,N_2310);
nand U2580 (N_2580,N_2373,N_2480);
or U2581 (N_2581,N_2351,N_2255);
nand U2582 (N_2582,N_2154,N_2489);
and U2583 (N_2583,N_2478,N_2225);
xnor U2584 (N_2584,N_2132,N_2372);
or U2585 (N_2585,N_2145,N_2044);
and U2586 (N_2586,N_2347,N_2002);
or U2587 (N_2587,N_2297,N_2490);
and U2588 (N_2588,N_2275,N_2219);
nor U2589 (N_2589,N_2407,N_2439);
nand U2590 (N_2590,N_2186,N_2452);
and U2591 (N_2591,N_2174,N_2391);
or U2592 (N_2592,N_2429,N_2417);
nand U2593 (N_2593,N_2305,N_2100);
and U2594 (N_2594,N_2400,N_2446);
and U2595 (N_2595,N_2080,N_2456);
xnor U2596 (N_2596,N_2156,N_2108);
nor U2597 (N_2597,N_2289,N_2138);
nor U2598 (N_2598,N_2277,N_2148);
or U2599 (N_2599,N_2422,N_2413);
xnor U2600 (N_2600,N_2126,N_2265);
nand U2601 (N_2601,N_2214,N_2019);
or U2602 (N_2602,N_2405,N_2075);
and U2603 (N_2603,N_2171,N_2093);
and U2604 (N_2604,N_2067,N_2425);
or U2605 (N_2605,N_2048,N_2307);
or U2606 (N_2606,N_2484,N_2123);
nor U2607 (N_2607,N_2254,N_2034);
xnor U2608 (N_2608,N_2053,N_2070);
nor U2609 (N_2609,N_2447,N_2240);
or U2610 (N_2610,N_2416,N_2444);
nand U2611 (N_2611,N_2418,N_2023);
or U2612 (N_2612,N_2188,N_2182);
or U2613 (N_2613,N_2483,N_2367);
nand U2614 (N_2614,N_2247,N_2383);
and U2615 (N_2615,N_2004,N_2139);
nand U2616 (N_2616,N_2049,N_2180);
nor U2617 (N_2617,N_2344,N_2249);
nand U2618 (N_2618,N_2218,N_2341);
or U2619 (N_2619,N_2274,N_2051);
nand U2620 (N_2620,N_2179,N_2124);
nor U2621 (N_2621,N_2168,N_2204);
nand U2622 (N_2622,N_2001,N_2256);
nor U2623 (N_2623,N_2497,N_2371);
or U2624 (N_2624,N_2059,N_2459);
nand U2625 (N_2625,N_2011,N_2454);
nand U2626 (N_2626,N_2353,N_2440);
nor U2627 (N_2627,N_2235,N_2266);
or U2628 (N_2628,N_2298,N_2430);
xor U2629 (N_2629,N_2368,N_2485);
nand U2630 (N_2630,N_2037,N_2195);
nor U2631 (N_2631,N_2083,N_2263);
nand U2632 (N_2632,N_2091,N_2248);
nand U2633 (N_2633,N_2094,N_2264);
or U2634 (N_2634,N_2365,N_2061);
and U2635 (N_2635,N_2163,N_2205);
nand U2636 (N_2636,N_2267,N_2377);
nand U2637 (N_2637,N_2328,N_2013);
nand U2638 (N_2638,N_2095,N_2487);
xnor U2639 (N_2639,N_2190,N_2181);
or U2640 (N_2640,N_2115,N_2448);
xnor U2641 (N_2641,N_2009,N_2363);
and U2642 (N_2642,N_2465,N_2153);
xnor U2643 (N_2643,N_2309,N_2217);
and U2644 (N_2644,N_2144,N_2324);
xnor U2645 (N_2645,N_2158,N_2366);
or U2646 (N_2646,N_2477,N_2222);
nor U2647 (N_2647,N_2323,N_2338);
xor U2648 (N_2648,N_2253,N_2166);
nor U2649 (N_2649,N_2451,N_2042);
nor U2650 (N_2650,N_2415,N_2278);
nand U2651 (N_2651,N_2107,N_2486);
nand U2652 (N_2652,N_2215,N_2043);
or U2653 (N_2653,N_2211,N_2238);
nand U2654 (N_2654,N_2125,N_2149);
nand U2655 (N_2655,N_2287,N_2140);
and U2656 (N_2656,N_2329,N_2453);
xnor U2657 (N_2657,N_2224,N_2272);
and U2658 (N_2658,N_2423,N_2152);
nor U2659 (N_2659,N_2088,N_2482);
and U2660 (N_2660,N_2320,N_2352);
nand U2661 (N_2661,N_2354,N_2499);
xnor U2662 (N_2662,N_2177,N_2031);
xor U2663 (N_2663,N_2096,N_2223);
nor U2664 (N_2664,N_2038,N_2343);
xor U2665 (N_2665,N_2410,N_2021);
and U2666 (N_2666,N_2104,N_2099);
and U2667 (N_2667,N_2442,N_2269);
or U2668 (N_2668,N_2319,N_2199);
or U2669 (N_2669,N_2007,N_2312);
nand U2670 (N_2670,N_2460,N_2127);
nor U2671 (N_2671,N_2342,N_2251);
nand U2672 (N_2672,N_2017,N_2474);
and U2673 (N_2673,N_2089,N_2191);
or U2674 (N_2674,N_2160,N_2027);
and U2675 (N_2675,N_2472,N_2349);
nor U2676 (N_2676,N_2151,N_2040);
nor U2677 (N_2677,N_2291,N_2078);
nor U2678 (N_2678,N_2146,N_2392);
nor U2679 (N_2679,N_2336,N_2194);
and U2680 (N_2680,N_2314,N_2073);
and U2681 (N_2681,N_2420,N_2176);
nor U2682 (N_2682,N_2102,N_2246);
nand U2683 (N_2683,N_2419,N_2303);
nand U2684 (N_2684,N_2424,N_2062);
nor U2685 (N_2685,N_2262,N_2355);
xor U2686 (N_2686,N_2090,N_2379);
and U2687 (N_2687,N_2491,N_2350);
nand U2688 (N_2688,N_2464,N_2234);
xor U2689 (N_2689,N_2050,N_2134);
and U2690 (N_2690,N_2129,N_2086);
xnor U2691 (N_2691,N_2438,N_2466);
xnor U2692 (N_2692,N_2250,N_2357);
xnor U2693 (N_2693,N_2066,N_2110);
nand U2694 (N_2694,N_2258,N_2128);
or U2695 (N_2695,N_2047,N_2443);
nand U2696 (N_2696,N_2198,N_2111);
nand U2697 (N_2697,N_2221,N_2178);
nor U2698 (N_2698,N_2183,N_2155);
and U2699 (N_2699,N_2458,N_2014);
and U2700 (N_2700,N_2322,N_2387);
and U2701 (N_2701,N_2479,N_2057);
and U2702 (N_2702,N_2189,N_2020);
nand U2703 (N_2703,N_2370,N_2302);
nand U2704 (N_2704,N_2098,N_2260);
xor U2705 (N_2705,N_2469,N_2033);
nor U2706 (N_2706,N_2316,N_2076);
or U2707 (N_2707,N_2003,N_2300);
nor U2708 (N_2708,N_2113,N_2280);
nor U2709 (N_2709,N_2493,N_2346);
or U2710 (N_2710,N_2295,N_2270);
or U2711 (N_2711,N_2226,N_2103);
or U2712 (N_2712,N_2032,N_2130);
xnor U2713 (N_2713,N_2200,N_2356);
nand U2714 (N_2714,N_2321,N_2361);
xnor U2715 (N_2715,N_2308,N_2237);
or U2716 (N_2716,N_2292,N_2006);
nor U2717 (N_2717,N_2318,N_2494);
nand U2718 (N_2718,N_2481,N_2384);
nor U2719 (N_2719,N_2092,N_2055);
or U2720 (N_2720,N_2364,N_2046);
nor U2721 (N_2721,N_2374,N_2058);
nor U2722 (N_2722,N_2242,N_2359);
xor U2723 (N_2723,N_2283,N_2169);
nor U2724 (N_2724,N_2087,N_2408);
or U2725 (N_2725,N_2245,N_2395);
or U2726 (N_2726,N_2330,N_2381);
and U2727 (N_2727,N_2276,N_2401);
nand U2728 (N_2728,N_2285,N_2084);
nor U2729 (N_2729,N_2228,N_2411);
nor U2730 (N_2730,N_2450,N_2306);
nor U2731 (N_2731,N_2173,N_2024);
and U2732 (N_2732,N_2476,N_2147);
or U2733 (N_2733,N_2244,N_2333);
nor U2734 (N_2734,N_2428,N_2282);
or U2735 (N_2735,N_2461,N_2432);
nor U2736 (N_2736,N_2119,N_2455);
nor U2737 (N_2737,N_2052,N_2437);
or U2738 (N_2738,N_2397,N_2210);
nand U2739 (N_2739,N_2369,N_2025);
xnor U2740 (N_2740,N_2041,N_2293);
nor U2741 (N_2741,N_2449,N_2394);
nand U2742 (N_2742,N_2233,N_2187);
xnor U2743 (N_2743,N_2290,N_2143);
nor U2744 (N_2744,N_2141,N_2498);
nor U2745 (N_2745,N_2261,N_2299);
nor U2746 (N_2746,N_2360,N_2216);
nor U2747 (N_2747,N_2036,N_2304);
and U2748 (N_2748,N_2252,N_2294);
xor U2749 (N_2749,N_2412,N_2470);
or U2750 (N_2750,N_2168,N_2303);
or U2751 (N_2751,N_2154,N_2160);
nor U2752 (N_2752,N_2114,N_2435);
xnor U2753 (N_2753,N_2034,N_2052);
or U2754 (N_2754,N_2436,N_2270);
or U2755 (N_2755,N_2198,N_2351);
xor U2756 (N_2756,N_2473,N_2125);
nor U2757 (N_2757,N_2060,N_2269);
nand U2758 (N_2758,N_2009,N_2257);
and U2759 (N_2759,N_2428,N_2114);
nor U2760 (N_2760,N_2098,N_2117);
xor U2761 (N_2761,N_2321,N_2294);
or U2762 (N_2762,N_2064,N_2011);
or U2763 (N_2763,N_2310,N_2084);
nor U2764 (N_2764,N_2363,N_2440);
xnor U2765 (N_2765,N_2435,N_2322);
xor U2766 (N_2766,N_2111,N_2306);
nand U2767 (N_2767,N_2029,N_2488);
nor U2768 (N_2768,N_2406,N_2456);
nand U2769 (N_2769,N_2335,N_2417);
nor U2770 (N_2770,N_2030,N_2043);
nor U2771 (N_2771,N_2171,N_2431);
nand U2772 (N_2772,N_2341,N_2059);
and U2773 (N_2773,N_2461,N_2333);
xor U2774 (N_2774,N_2183,N_2271);
nor U2775 (N_2775,N_2073,N_2167);
and U2776 (N_2776,N_2345,N_2091);
nor U2777 (N_2777,N_2307,N_2178);
nand U2778 (N_2778,N_2382,N_2055);
or U2779 (N_2779,N_2330,N_2053);
or U2780 (N_2780,N_2058,N_2437);
nor U2781 (N_2781,N_2493,N_2497);
nand U2782 (N_2782,N_2459,N_2375);
nand U2783 (N_2783,N_2041,N_2485);
and U2784 (N_2784,N_2218,N_2038);
nand U2785 (N_2785,N_2190,N_2330);
or U2786 (N_2786,N_2106,N_2175);
nand U2787 (N_2787,N_2057,N_2082);
nand U2788 (N_2788,N_2396,N_2214);
or U2789 (N_2789,N_2152,N_2049);
nor U2790 (N_2790,N_2110,N_2335);
nand U2791 (N_2791,N_2178,N_2183);
nor U2792 (N_2792,N_2146,N_2213);
or U2793 (N_2793,N_2263,N_2259);
and U2794 (N_2794,N_2026,N_2476);
and U2795 (N_2795,N_2334,N_2127);
nand U2796 (N_2796,N_2448,N_2349);
nand U2797 (N_2797,N_2126,N_2215);
or U2798 (N_2798,N_2227,N_2324);
nand U2799 (N_2799,N_2095,N_2227);
xor U2800 (N_2800,N_2416,N_2022);
or U2801 (N_2801,N_2004,N_2383);
xnor U2802 (N_2802,N_2183,N_2462);
or U2803 (N_2803,N_2087,N_2399);
or U2804 (N_2804,N_2267,N_2023);
or U2805 (N_2805,N_2344,N_2400);
xnor U2806 (N_2806,N_2002,N_2486);
nor U2807 (N_2807,N_2463,N_2047);
and U2808 (N_2808,N_2427,N_2154);
or U2809 (N_2809,N_2330,N_2010);
nand U2810 (N_2810,N_2260,N_2160);
xnor U2811 (N_2811,N_2460,N_2325);
nand U2812 (N_2812,N_2000,N_2431);
or U2813 (N_2813,N_2238,N_2265);
nor U2814 (N_2814,N_2069,N_2022);
nor U2815 (N_2815,N_2031,N_2244);
nor U2816 (N_2816,N_2392,N_2026);
nor U2817 (N_2817,N_2368,N_2204);
xor U2818 (N_2818,N_2070,N_2351);
and U2819 (N_2819,N_2120,N_2060);
and U2820 (N_2820,N_2147,N_2015);
nand U2821 (N_2821,N_2359,N_2494);
xnor U2822 (N_2822,N_2207,N_2123);
nor U2823 (N_2823,N_2211,N_2372);
or U2824 (N_2824,N_2328,N_2122);
nor U2825 (N_2825,N_2195,N_2396);
or U2826 (N_2826,N_2038,N_2010);
or U2827 (N_2827,N_2388,N_2476);
and U2828 (N_2828,N_2266,N_2009);
nor U2829 (N_2829,N_2010,N_2144);
nor U2830 (N_2830,N_2335,N_2132);
or U2831 (N_2831,N_2278,N_2034);
nor U2832 (N_2832,N_2435,N_2311);
or U2833 (N_2833,N_2128,N_2046);
nor U2834 (N_2834,N_2459,N_2001);
and U2835 (N_2835,N_2234,N_2272);
xnor U2836 (N_2836,N_2238,N_2456);
or U2837 (N_2837,N_2259,N_2336);
and U2838 (N_2838,N_2203,N_2106);
nor U2839 (N_2839,N_2077,N_2261);
nand U2840 (N_2840,N_2303,N_2169);
nand U2841 (N_2841,N_2051,N_2220);
nor U2842 (N_2842,N_2350,N_2119);
or U2843 (N_2843,N_2349,N_2436);
xor U2844 (N_2844,N_2185,N_2472);
and U2845 (N_2845,N_2116,N_2001);
xnor U2846 (N_2846,N_2458,N_2088);
nor U2847 (N_2847,N_2446,N_2307);
nor U2848 (N_2848,N_2497,N_2107);
and U2849 (N_2849,N_2125,N_2081);
nand U2850 (N_2850,N_2017,N_2311);
xnor U2851 (N_2851,N_2289,N_2239);
nand U2852 (N_2852,N_2086,N_2327);
or U2853 (N_2853,N_2191,N_2430);
xor U2854 (N_2854,N_2115,N_2279);
xnor U2855 (N_2855,N_2280,N_2110);
xor U2856 (N_2856,N_2178,N_2127);
or U2857 (N_2857,N_2420,N_2364);
and U2858 (N_2858,N_2049,N_2315);
nor U2859 (N_2859,N_2096,N_2190);
or U2860 (N_2860,N_2357,N_2143);
xnor U2861 (N_2861,N_2003,N_2470);
nor U2862 (N_2862,N_2403,N_2164);
xnor U2863 (N_2863,N_2180,N_2068);
nor U2864 (N_2864,N_2176,N_2034);
nor U2865 (N_2865,N_2139,N_2345);
or U2866 (N_2866,N_2096,N_2236);
and U2867 (N_2867,N_2006,N_2456);
and U2868 (N_2868,N_2325,N_2183);
nor U2869 (N_2869,N_2304,N_2350);
or U2870 (N_2870,N_2263,N_2454);
nand U2871 (N_2871,N_2093,N_2417);
nand U2872 (N_2872,N_2493,N_2176);
nor U2873 (N_2873,N_2068,N_2166);
nand U2874 (N_2874,N_2311,N_2155);
xor U2875 (N_2875,N_2292,N_2171);
and U2876 (N_2876,N_2059,N_2414);
and U2877 (N_2877,N_2018,N_2114);
nand U2878 (N_2878,N_2110,N_2303);
xnor U2879 (N_2879,N_2410,N_2224);
nand U2880 (N_2880,N_2089,N_2193);
and U2881 (N_2881,N_2172,N_2438);
xnor U2882 (N_2882,N_2302,N_2460);
and U2883 (N_2883,N_2299,N_2202);
and U2884 (N_2884,N_2096,N_2277);
nor U2885 (N_2885,N_2099,N_2218);
or U2886 (N_2886,N_2362,N_2164);
nor U2887 (N_2887,N_2258,N_2006);
nor U2888 (N_2888,N_2020,N_2062);
xnor U2889 (N_2889,N_2176,N_2139);
nand U2890 (N_2890,N_2017,N_2313);
and U2891 (N_2891,N_2005,N_2433);
and U2892 (N_2892,N_2325,N_2269);
nand U2893 (N_2893,N_2221,N_2385);
and U2894 (N_2894,N_2047,N_2150);
xnor U2895 (N_2895,N_2004,N_2169);
and U2896 (N_2896,N_2431,N_2269);
nand U2897 (N_2897,N_2027,N_2176);
nand U2898 (N_2898,N_2085,N_2143);
or U2899 (N_2899,N_2141,N_2364);
xor U2900 (N_2900,N_2346,N_2397);
and U2901 (N_2901,N_2428,N_2437);
xor U2902 (N_2902,N_2183,N_2058);
and U2903 (N_2903,N_2021,N_2063);
nand U2904 (N_2904,N_2174,N_2224);
or U2905 (N_2905,N_2461,N_2268);
nand U2906 (N_2906,N_2475,N_2477);
or U2907 (N_2907,N_2131,N_2113);
nor U2908 (N_2908,N_2474,N_2119);
nand U2909 (N_2909,N_2057,N_2410);
nor U2910 (N_2910,N_2198,N_2377);
and U2911 (N_2911,N_2127,N_2351);
nor U2912 (N_2912,N_2027,N_2464);
nor U2913 (N_2913,N_2105,N_2039);
nor U2914 (N_2914,N_2300,N_2139);
xnor U2915 (N_2915,N_2013,N_2025);
xor U2916 (N_2916,N_2060,N_2314);
xnor U2917 (N_2917,N_2290,N_2287);
or U2918 (N_2918,N_2433,N_2290);
or U2919 (N_2919,N_2212,N_2094);
xor U2920 (N_2920,N_2019,N_2150);
or U2921 (N_2921,N_2024,N_2140);
nor U2922 (N_2922,N_2062,N_2327);
nand U2923 (N_2923,N_2103,N_2188);
and U2924 (N_2924,N_2031,N_2218);
and U2925 (N_2925,N_2124,N_2109);
nand U2926 (N_2926,N_2296,N_2426);
and U2927 (N_2927,N_2136,N_2254);
xor U2928 (N_2928,N_2200,N_2495);
nor U2929 (N_2929,N_2464,N_2314);
nor U2930 (N_2930,N_2365,N_2089);
and U2931 (N_2931,N_2028,N_2265);
or U2932 (N_2932,N_2468,N_2490);
or U2933 (N_2933,N_2351,N_2197);
nand U2934 (N_2934,N_2258,N_2380);
xnor U2935 (N_2935,N_2086,N_2110);
nor U2936 (N_2936,N_2026,N_2372);
nand U2937 (N_2937,N_2119,N_2335);
nand U2938 (N_2938,N_2161,N_2256);
nand U2939 (N_2939,N_2163,N_2290);
or U2940 (N_2940,N_2313,N_2276);
nand U2941 (N_2941,N_2122,N_2472);
nor U2942 (N_2942,N_2155,N_2020);
nand U2943 (N_2943,N_2315,N_2475);
nor U2944 (N_2944,N_2122,N_2172);
nand U2945 (N_2945,N_2084,N_2165);
and U2946 (N_2946,N_2113,N_2437);
and U2947 (N_2947,N_2280,N_2481);
and U2948 (N_2948,N_2181,N_2369);
nand U2949 (N_2949,N_2077,N_2194);
and U2950 (N_2950,N_2253,N_2073);
and U2951 (N_2951,N_2428,N_2419);
or U2952 (N_2952,N_2225,N_2454);
nand U2953 (N_2953,N_2398,N_2339);
xor U2954 (N_2954,N_2241,N_2196);
and U2955 (N_2955,N_2323,N_2412);
xor U2956 (N_2956,N_2296,N_2440);
nor U2957 (N_2957,N_2265,N_2088);
nor U2958 (N_2958,N_2303,N_2022);
xor U2959 (N_2959,N_2225,N_2253);
nor U2960 (N_2960,N_2178,N_2430);
nor U2961 (N_2961,N_2095,N_2166);
nor U2962 (N_2962,N_2068,N_2223);
or U2963 (N_2963,N_2440,N_2359);
xor U2964 (N_2964,N_2291,N_2103);
and U2965 (N_2965,N_2387,N_2284);
nand U2966 (N_2966,N_2348,N_2477);
or U2967 (N_2967,N_2103,N_2228);
nor U2968 (N_2968,N_2394,N_2161);
and U2969 (N_2969,N_2302,N_2355);
nor U2970 (N_2970,N_2011,N_2453);
nand U2971 (N_2971,N_2116,N_2462);
or U2972 (N_2972,N_2300,N_2009);
nor U2973 (N_2973,N_2144,N_2017);
nand U2974 (N_2974,N_2134,N_2200);
or U2975 (N_2975,N_2226,N_2082);
xnor U2976 (N_2976,N_2042,N_2480);
and U2977 (N_2977,N_2434,N_2121);
nand U2978 (N_2978,N_2185,N_2254);
and U2979 (N_2979,N_2326,N_2159);
nor U2980 (N_2980,N_2381,N_2135);
xnor U2981 (N_2981,N_2171,N_2014);
nor U2982 (N_2982,N_2355,N_2015);
nor U2983 (N_2983,N_2309,N_2279);
nor U2984 (N_2984,N_2447,N_2140);
nor U2985 (N_2985,N_2328,N_2398);
or U2986 (N_2986,N_2231,N_2077);
or U2987 (N_2987,N_2341,N_2464);
and U2988 (N_2988,N_2102,N_2005);
nor U2989 (N_2989,N_2097,N_2302);
nand U2990 (N_2990,N_2431,N_2328);
xor U2991 (N_2991,N_2086,N_2252);
nand U2992 (N_2992,N_2354,N_2025);
and U2993 (N_2993,N_2459,N_2435);
nand U2994 (N_2994,N_2297,N_2192);
or U2995 (N_2995,N_2012,N_2112);
nor U2996 (N_2996,N_2164,N_2344);
nand U2997 (N_2997,N_2114,N_2130);
or U2998 (N_2998,N_2219,N_2446);
nor U2999 (N_2999,N_2441,N_2196);
nand U3000 (N_3000,N_2946,N_2724);
nand U3001 (N_3001,N_2607,N_2961);
nor U3002 (N_3002,N_2694,N_2606);
nand U3003 (N_3003,N_2516,N_2797);
and U3004 (N_3004,N_2661,N_2662);
nand U3005 (N_3005,N_2774,N_2522);
and U3006 (N_3006,N_2783,N_2872);
and U3007 (N_3007,N_2583,N_2752);
or U3008 (N_3008,N_2560,N_2845);
or U3009 (N_3009,N_2574,N_2646);
nor U3010 (N_3010,N_2943,N_2954);
and U3011 (N_3011,N_2543,N_2830);
nor U3012 (N_3012,N_2802,N_2926);
and U3013 (N_3013,N_2894,N_2692);
xor U3014 (N_3014,N_2799,N_2586);
nand U3015 (N_3015,N_2791,N_2908);
nor U3016 (N_3016,N_2949,N_2902);
xor U3017 (N_3017,N_2892,N_2742);
xnor U3018 (N_3018,N_2660,N_2823);
and U3019 (N_3019,N_2681,N_2804);
or U3020 (N_3020,N_2618,N_2502);
nand U3021 (N_3021,N_2716,N_2906);
xor U3022 (N_3022,N_2856,N_2763);
nand U3023 (N_3023,N_2666,N_2665);
or U3024 (N_3024,N_2937,N_2948);
nor U3025 (N_3025,N_2966,N_2539);
nand U3026 (N_3026,N_2995,N_2792);
xnor U3027 (N_3027,N_2918,N_2766);
xor U3028 (N_3028,N_2858,N_2729);
nor U3029 (N_3029,N_2749,N_2537);
nor U3030 (N_3030,N_2726,N_2691);
xnor U3031 (N_3031,N_2655,N_2865);
nand U3032 (N_3032,N_2754,N_2788);
xor U3033 (N_3033,N_2887,N_2520);
and U3034 (N_3034,N_2934,N_2773);
xnor U3035 (N_3035,N_2873,N_2963);
and U3036 (N_3036,N_2815,N_2523);
and U3037 (N_3037,N_2953,N_2593);
nor U3038 (N_3038,N_2955,N_2693);
nor U3039 (N_3039,N_2893,N_2811);
or U3040 (N_3040,N_2862,N_2825);
or U3041 (N_3041,N_2798,N_2772);
xor U3042 (N_3042,N_2542,N_2679);
nand U3043 (N_3043,N_2617,N_2989);
nor U3044 (N_3044,N_2612,N_2891);
nor U3045 (N_3045,N_2707,N_2972);
nand U3046 (N_3046,N_2636,N_2680);
and U3047 (N_3047,N_2981,N_2965);
and U3048 (N_3048,N_2806,N_2909);
and U3049 (N_3049,N_2718,N_2736);
or U3050 (N_3050,N_2820,N_2577);
nand U3051 (N_3051,N_2647,N_2581);
or U3052 (N_3052,N_2822,N_2855);
nand U3053 (N_3053,N_2505,N_2985);
or U3054 (N_3054,N_2641,N_2904);
nand U3055 (N_3055,N_2915,N_2905);
xnor U3056 (N_3056,N_2675,N_2594);
xnor U3057 (N_3057,N_2973,N_2554);
nor U3058 (N_3058,N_2785,N_2698);
or U3059 (N_3059,N_2920,N_2957);
and U3060 (N_3060,N_2673,N_2575);
nor U3061 (N_3061,N_2923,N_2750);
or U3062 (N_3062,N_2587,N_2759);
xnor U3063 (N_3063,N_2927,N_2870);
nand U3064 (N_3064,N_2551,N_2640);
nor U3065 (N_3065,N_2595,N_2987);
and U3066 (N_3066,N_2755,N_2760);
or U3067 (N_3067,N_2863,N_2980);
nand U3068 (N_3068,N_2968,N_2991);
nand U3069 (N_3069,N_2510,N_2525);
and U3070 (N_3070,N_2992,N_2877);
nand U3071 (N_3071,N_2951,N_2964);
and U3072 (N_3072,N_2999,N_2690);
and U3073 (N_3073,N_2765,N_2795);
nor U3074 (N_3074,N_2901,N_2545);
nor U3075 (N_3075,N_2580,N_2710);
nand U3076 (N_3076,N_2851,N_2935);
xnor U3077 (N_3077,N_2850,N_2881);
nand U3078 (N_3078,N_2979,N_2816);
nor U3079 (N_3079,N_2558,N_2883);
and U3080 (N_3080,N_2814,N_2743);
nand U3081 (N_3081,N_2534,N_2559);
xor U3082 (N_3082,N_2631,N_2501);
or U3083 (N_3083,N_2805,N_2711);
or U3084 (N_3084,N_2609,N_2764);
xor U3085 (N_3085,N_2713,N_2531);
and U3086 (N_3086,N_2738,N_2977);
and U3087 (N_3087,N_2960,N_2996);
nand U3088 (N_3088,N_2614,N_2727);
or U3089 (N_3089,N_2890,N_2967);
and U3090 (N_3090,N_2793,N_2526);
or U3091 (N_3091,N_2770,N_2982);
and U3092 (N_3092,N_2590,N_2530);
xnor U3093 (N_3093,N_2599,N_2637);
and U3094 (N_3094,N_2549,N_2807);
nor U3095 (N_3095,N_2834,N_2635);
nand U3096 (N_3096,N_2723,N_2734);
nand U3097 (N_3097,N_2553,N_2817);
nand U3098 (N_3098,N_2848,N_2997);
xnor U3099 (N_3099,N_2677,N_2767);
and U3100 (N_3100,N_2527,N_2653);
nor U3101 (N_3101,N_2535,N_2676);
or U3102 (N_3102,N_2952,N_2518);
and U3103 (N_3103,N_2717,N_2928);
nor U3104 (N_3104,N_2888,N_2550);
nor U3105 (N_3105,N_2623,N_2566);
and U3106 (N_3106,N_2777,N_2719);
xor U3107 (N_3107,N_2567,N_2757);
nand U3108 (N_3108,N_2541,N_2866);
xnor U3109 (N_3109,N_2878,N_2624);
nor U3110 (N_3110,N_2591,N_2896);
nand U3111 (N_3111,N_2859,N_2688);
and U3112 (N_3112,N_2740,N_2514);
nand U3113 (N_3113,N_2990,N_2974);
or U3114 (N_3114,N_2976,N_2503);
xor U3115 (N_3115,N_2652,N_2854);
xnor U3116 (N_3116,N_2867,N_2782);
nor U3117 (N_3117,N_2720,N_2648);
and U3118 (N_3118,N_2962,N_2644);
and U3119 (N_3119,N_2722,N_2536);
or U3120 (N_3120,N_2784,N_2538);
and U3121 (N_3121,N_2628,N_2658);
nand U3122 (N_3122,N_2731,N_2544);
nor U3123 (N_3123,N_2900,N_2689);
and U3124 (N_3124,N_2512,N_2875);
nand U3125 (N_3125,N_2695,N_2843);
nand U3126 (N_3126,N_2939,N_2708);
and U3127 (N_3127,N_2746,N_2769);
nor U3128 (N_3128,N_2564,N_2801);
nor U3129 (N_3129,N_2500,N_2728);
and U3130 (N_3130,N_2584,N_2771);
and U3131 (N_3131,N_2778,N_2921);
nor U3132 (N_3132,N_2839,N_2576);
xnor U3133 (N_3133,N_2956,N_2751);
nor U3134 (N_3134,N_2712,N_2657);
or U3135 (N_3135,N_2916,N_2971);
and U3136 (N_3136,N_2936,N_2533);
xor U3137 (N_3137,N_2944,N_2899);
nor U3138 (N_3138,N_2903,N_2611);
xnor U3139 (N_3139,N_2781,N_2803);
xor U3140 (N_3140,N_2630,N_2813);
nor U3141 (N_3141,N_2786,N_2715);
and U3142 (N_3142,N_2563,N_2886);
and U3143 (N_3143,N_2827,N_2546);
nand U3144 (N_3144,N_2589,N_2914);
xnor U3145 (N_3145,N_2958,N_2998);
and U3146 (N_3146,N_2733,N_2568);
and U3147 (N_3147,N_2620,N_2669);
or U3148 (N_3148,N_2622,N_2730);
nand U3149 (N_3149,N_2632,N_2600);
or U3150 (N_3150,N_2959,N_2790);
nor U3151 (N_3151,N_2598,N_2950);
or U3152 (N_3152,N_2508,N_2868);
and U3153 (N_3153,N_2701,N_2643);
and U3154 (N_3154,N_2838,N_2529);
nand U3155 (N_3155,N_2664,N_2604);
and U3156 (N_3156,N_2696,N_2672);
or U3157 (N_3157,N_2684,N_2621);
nor U3158 (N_3158,N_2744,N_2513);
xnor U3159 (N_3159,N_2809,N_2940);
nor U3160 (N_3160,N_2524,N_2861);
xnor U3161 (N_3161,N_2678,N_2638);
and U3162 (N_3162,N_2613,N_2569);
xnor U3163 (N_3163,N_2933,N_2919);
and U3164 (N_3164,N_2970,N_2945);
or U3165 (N_3165,N_2619,N_2789);
and U3166 (N_3166,N_2645,N_2649);
xor U3167 (N_3167,N_2706,N_2885);
or U3168 (N_3168,N_2685,N_2924);
and U3169 (N_3169,N_2704,N_2555);
nand U3170 (N_3170,N_2853,N_2847);
and U3171 (N_3171,N_2651,N_2504);
and U3172 (N_3172,N_2860,N_2884);
xnor U3173 (N_3173,N_2849,N_2938);
and U3174 (N_3174,N_2824,N_2983);
nor U3175 (N_3175,N_2633,N_2882);
nand U3176 (N_3176,N_2929,N_2829);
xnor U3177 (N_3177,N_2776,N_2922);
nand U3178 (N_3178,N_2913,N_2988);
nor U3179 (N_3179,N_2747,N_2852);
nand U3180 (N_3180,N_2548,N_2532);
nor U3181 (N_3181,N_2605,N_2656);
nand U3182 (N_3182,N_2602,N_2697);
nor U3183 (N_3183,N_2596,N_2753);
nor U3184 (N_3184,N_2984,N_2917);
nand U3185 (N_3185,N_2654,N_2840);
and U3186 (N_3186,N_2519,N_2842);
or U3187 (N_3187,N_2642,N_2570);
xnor U3188 (N_3188,N_2898,N_2857);
xor U3189 (N_3189,N_2650,N_2846);
nor U3190 (N_3190,N_2741,N_2528);
or U3191 (N_3191,N_2779,N_2756);
and U3192 (N_3192,N_2699,N_2796);
and U3193 (N_3193,N_2841,N_2725);
xnor U3194 (N_3194,N_2969,N_2907);
nand U3195 (N_3195,N_2674,N_2748);
nor U3196 (N_3196,N_2876,N_2941);
xor U3197 (N_3197,N_2597,N_2561);
and U3198 (N_3198,N_2703,N_2592);
and U3199 (N_3199,N_2578,N_2603);
nor U3200 (N_3200,N_2932,N_2844);
and U3201 (N_3201,N_2615,N_2818);
xnor U3202 (N_3202,N_2687,N_2702);
and U3203 (N_3203,N_2836,N_2511);
xnor U3204 (N_3204,N_2761,N_2625);
nor U3205 (N_3205,N_2683,N_2874);
and U3206 (N_3206,N_2700,N_2745);
nand U3207 (N_3207,N_2616,N_2509);
nor U3208 (N_3208,N_2831,N_2864);
xor U3209 (N_3209,N_2629,N_2947);
xnor U3210 (N_3210,N_2735,N_2552);
or U3211 (N_3211,N_2714,N_2925);
nand U3212 (N_3212,N_2762,N_2709);
and U3213 (N_3213,N_2506,N_2572);
and U3214 (N_3214,N_2837,N_2768);
nor U3215 (N_3215,N_2889,N_2871);
and U3216 (N_3216,N_2540,N_2556);
and U3217 (N_3217,N_2670,N_2880);
xnor U3218 (N_3218,N_2808,N_2810);
and U3219 (N_3219,N_2721,N_2758);
nor U3220 (N_3220,N_2910,N_2780);
xor U3221 (N_3221,N_2671,N_2812);
nor U3222 (N_3222,N_2521,N_2562);
nand U3223 (N_3223,N_2821,N_2517);
nand U3224 (N_3224,N_2663,N_2942);
nand U3225 (N_3225,N_2557,N_2579);
or U3226 (N_3226,N_2634,N_2828);
nor U3227 (N_3227,N_2739,N_2667);
or U3228 (N_3228,N_2705,N_2737);
or U3229 (N_3229,N_2930,N_2978);
nand U3230 (N_3230,N_2895,N_2826);
and U3231 (N_3231,N_2787,N_2912);
xor U3232 (N_3232,N_2627,N_2668);
nor U3233 (N_3233,N_2775,N_2639);
or U3234 (N_3234,N_2835,N_2682);
and U3235 (N_3235,N_2832,N_2507);
and U3236 (N_3236,N_2794,N_2897);
or U3237 (N_3237,N_2975,N_2879);
nand U3238 (N_3238,N_2911,N_2732);
xnor U3239 (N_3239,N_2588,N_2986);
nor U3240 (N_3240,N_2573,N_2571);
nor U3241 (N_3241,N_2931,N_2659);
xor U3242 (N_3242,N_2608,N_2833);
xor U3243 (N_3243,N_2601,N_2582);
xnor U3244 (N_3244,N_2585,N_2800);
and U3245 (N_3245,N_2515,N_2565);
nor U3246 (N_3246,N_2686,N_2994);
nand U3247 (N_3247,N_2869,N_2547);
nor U3248 (N_3248,N_2626,N_2993);
xnor U3249 (N_3249,N_2610,N_2819);
xnor U3250 (N_3250,N_2684,N_2843);
and U3251 (N_3251,N_2557,N_2616);
and U3252 (N_3252,N_2764,N_2737);
xnor U3253 (N_3253,N_2513,N_2895);
and U3254 (N_3254,N_2901,N_2624);
or U3255 (N_3255,N_2596,N_2927);
nand U3256 (N_3256,N_2698,N_2996);
nand U3257 (N_3257,N_2746,N_2610);
or U3258 (N_3258,N_2771,N_2596);
or U3259 (N_3259,N_2707,N_2847);
xor U3260 (N_3260,N_2844,N_2752);
xor U3261 (N_3261,N_2577,N_2713);
and U3262 (N_3262,N_2632,N_2614);
or U3263 (N_3263,N_2592,N_2584);
nor U3264 (N_3264,N_2794,N_2798);
nor U3265 (N_3265,N_2520,N_2781);
nor U3266 (N_3266,N_2608,N_2823);
nor U3267 (N_3267,N_2934,N_2745);
xor U3268 (N_3268,N_2824,N_2613);
nand U3269 (N_3269,N_2650,N_2967);
xnor U3270 (N_3270,N_2573,N_2720);
and U3271 (N_3271,N_2571,N_2958);
and U3272 (N_3272,N_2802,N_2922);
xnor U3273 (N_3273,N_2505,N_2646);
nor U3274 (N_3274,N_2690,N_2579);
or U3275 (N_3275,N_2536,N_2797);
nor U3276 (N_3276,N_2500,N_2971);
nor U3277 (N_3277,N_2687,N_2895);
nand U3278 (N_3278,N_2657,N_2621);
nand U3279 (N_3279,N_2606,N_2702);
and U3280 (N_3280,N_2536,N_2598);
nand U3281 (N_3281,N_2503,N_2973);
or U3282 (N_3282,N_2606,N_2773);
nand U3283 (N_3283,N_2655,N_2644);
nor U3284 (N_3284,N_2582,N_2578);
and U3285 (N_3285,N_2681,N_2665);
nor U3286 (N_3286,N_2565,N_2669);
nand U3287 (N_3287,N_2983,N_2556);
and U3288 (N_3288,N_2666,N_2805);
and U3289 (N_3289,N_2705,N_2601);
and U3290 (N_3290,N_2879,N_2983);
nor U3291 (N_3291,N_2966,N_2826);
or U3292 (N_3292,N_2811,N_2673);
or U3293 (N_3293,N_2982,N_2753);
xnor U3294 (N_3294,N_2836,N_2732);
nor U3295 (N_3295,N_2755,N_2813);
nand U3296 (N_3296,N_2764,N_2600);
nand U3297 (N_3297,N_2786,N_2630);
and U3298 (N_3298,N_2837,N_2832);
or U3299 (N_3299,N_2727,N_2628);
or U3300 (N_3300,N_2620,N_2853);
and U3301 (N_3301,N_2577,N_2654);
nand U3302 (N_3302,N_2915,N_2896);
and U3303 (N_3303,N_2511,N_2667);
nand U3304 (N_3304,N_2575,N_2730);
nand U3305 (N_3305,N_2754,N_2606);
and U3306 (N_3306,N_2605,N_2941);
or U3307 (N_3307,N_2735,N_2952);
nand U3308 (N_3308,N_2974,N_2783);
or U3309 (N_3309,N_2957,N_2515);
or U3310 (N_3310,N_2673,N_2996);
xor U3311 (N_3311,N_2506,N_2699);
and U3312 (N_3312,N_2827,N_2764);
or U3313 (N_3313,N_2795,N_2884);
nor U3314 (N_3314,N_2568,N_2849);
xor U3315 (N_3315,N_2680,N_2801);
nor U3316 (N_3316,N_2573,N_2714);
xnor U3317 (N_3317,N_2754,N_2899);
and U3318 (N_3318,N_2607,N_2654);
or U3319 (N_3319,N_2662,N_2549);
nor U3320 (N_3320,N_2811,N_2902);
or U3321 (N_3321,N_2990,N_2670);
and U3322 (N_3322,N_2545,N_2568);
nor U3323 (N_3323,N_2584,N_2637);
or U3324 (N_3324,N_2901,N_2916);
and U3325 (N_3325,N_2780,N_2754);
nor U3326 (N_3326,N_2540,N_2802);
nand U3327 (N_3327,N_2525,N_2870);
and U3328 (N_3328,N_2802,N_2899);
or U3329 (N_3329,N_2611,N_2841);
or U3330 (N_3330,N_2885,N_2655);
and U3331 (N_3331,N_2705,N_2590);
and U3332 (N_3332,N_2739,N_2625);
xor U3333 (N_3333,N_2548,N_2668);
nor U3334 (N_3334,N_2748,N_2551);
or U3335 (N_3335,N_2878,N_2742);
xor U3336 (N_3336,N_2851,N_2879);
or U3337 (N_3337,N_2913,N_2651);
nand U3338 (N_3338,N_2990,N_2864);
and U3339 (N_3339,N_2775,N_2958);
xnor U3340 (N_3340,N_2846,N_2635);
nand U3341 (N_3341,N_2896,N_2776);
and U3342 (N_3342,N_2808,N_2770);
xnor U3343 (N_3343,N_2917,N_2559);
nand U3344 (N_3344,N_2604,N_2563);
and U3345 (N_3345,N_2593,N_2724);
nor U3346 (N_3346,N_2715,N_2555);
or U3347 (N_3347,N_2738,N_2518);
or U3348 (N_3348,N_2929,N_2968);
nand U3349 (N_3349,N_2832,N_2763);
xor U3350 (N_3350,N_2602,N_2818);
nand U3351 (N_3351,N_2649,N_2595);
and U3352 (N_3352,N_2577,N_2780);
and U3353 (N_3353,N_2768,N_2730);
or U3354 (N_3354,N_2973,N_2864);
xnor U3355 (N_3355,N_2894,N_2964);
nand U3356 (N_3356,N_2849,N_2964);
nor U3357 (N_3357,N_2747,N_2523);
or U3358 (N_3358,N_2787,N_2743);
nand U3359 (N_3359,N_2668,N_2590);
nand U3360 (N_3360,N_2795,N_2784);
or U3361 (N_3361,N_2655,N_2523);
nand U3362 (N_3362,N_2963,N_2901);
and U3363 (N_3363,N_2769,N_2694);
xnor U3364 (N_3364,N_2865,N_2763);
or U3365 (N_3365,N_2543,N_2790);
and U3366 (N_3366,N_2714,N_2817);
xor U3367 (N_3367,N_2609,N_2923);
xnor U3368 (N_3368,N_2826,N_2670);
or U3369 (N_3369,N_2563,N_2624);
nor U3370 (N_3370,N_2576,N_2695);
nand U3371 (N_3371,N_2539,N_2663);
nand U3372 (N_3372,N_2762,N_2641);
or U3373 (N_3373,N_2843,N_2538);
xor U3374 (N_3374,N_2749,N_2798);
or U3375 (N_3375,N_2535,N_2684);
nor U3376 (N_3376,N_2884,N_2964);
and U3377 (N_3377,N_2689,N_2845);
nand U3378 (N_3378,N_2570,N_2986);
xnor U3379 (N_3379,N_2673,N_2823);
nor U3380 (N_3380,N_2985,N_2852);
nand U3381 (N_3381,N_2636,N_2865);
xnor U3382 (N_3382,N_2575,N_2591);
nand U3383 (N_3383,N_2981,N_2826);
and U3384 (N_3384,N_2696,N_2615);
xor U3385 (N_3385,N_2704,N_2808);
nand U3386 (N_3386,N_2932,N_2641);
and U3387 (N_3387,N_2666,N_2842);
nor U3388 (N_3388,N_2808,N_2729);
nand U3389 (N_3389,N_2771,N_2652);
xnor U3390 (N_3390,N_2916,N_2668);
nor U3391 (N_3391,N_2569,N_2797);
or U3392 (N_3392,N_2801,N_2950);
and U3393 (N_3393,N_2742,N_2515);
xnor U3394 (N_3394,N_2770,N_2788);
xnor U3395 (N_3395,N_2653,N_2762);
or U3396 (N_3396,N_2783,N_2786);
and U3397 (N_3397,N_2959,N_2786);
and U3398 (N_3398,N_2530,N_2933);
nand U3399 (N_3399,N_2847,N_2983);
or U3400 (N_3400,N_2573,N_2598);
xor U3401 (N_3401,N_2635,N_2977);
nand U3402 (N_3402,N_2639,N_2506);
or U3403 (N_3403,N_2805,N_2949);
xor U3404 (N_3404,N_2899,N_2780);
xor U3405 (N_3405,N_2704,N_2537);
xnor U3406 (N_3406,N_2646,N_2880);
xor U3407 (N_3407,N_2773,N_2576);
nand U3408 (N_3408,N_2888,N_2505);
nand U3409 (N_3409,N_2528,N_2641);
or U3410 (N_3410,N_2846,N_2536);
nand U3411 (N_3411,N_2501,N_2711);
or U3412 (N_3412,N_2832,N_2729);
nor U3413 (N_3413,N_2600,N_2935);
nor U3414 (N_3414,N_2628,N_2927);
nand U3415 (N_3415,N_2617,N_2528);
nor U3416 (N_3416,N_2752,N_2578);
and U3417 (N_3417,N_2965,N_2800);
nor U3418 (N_3418,N_2828,N_2742);
xnor U3419 (N_3419,N_2666,N_2906);
or U3420 (N_3420,N_2502,N_2576);
nand U3421 (N_3421,N_2778,N_2659);
or U3422 (N_3422,N_2808,N_2699);
or U3423 (N_3423,N_2661,N_2830);
or U3424 (N_3424,N_2963,N_2533);
nor U3425 (N_3425,N_2959,N_2810);
nor U3426 (N_3426,N_2921,N_2818);
and U3427 (N_3427,N_2633,N_2917);
or U3428 (N_3428,N_2505,N_2567);
nor U3429 (N_3429,N_2907,N_2666);
and U3430 (N_3430,N_2802,N_2569);
xor U3431 (N_3431,N_2998,N_2888);
nand U3432 (N_3432,N_2706,N_2603);
nor U3433 (N_3433,N_2536,N_2637);
nand U3434 (N_3434,N_2894,N_2530);
and U3435 (N_3435,N_2885,N_2724);
nand U3436 (N_3436,N_2810,N_2767);
nor U3437 (N_3437,N_2726,N_2993);
nand U3438 (N_3438,N_2864,N_2860);
nor U3439 (N_3439,N_2837,N_2621);
or U3440 (N_3440,N_2632,N_2730);
or U3441 (N_3441,N_2546,N_2981);
xnor U3442 (N_3442,N_2703,N_2996);
nand U3443 (N_3443,N_2530,N_2551);
or U3444 (N_3444,N_2627,N_2557);
or U3445 (N_3445,N_2870,N_2526);
nor U3446 (N_3446,N_2707,N_2768);
nand U3447 (N_3447,N_2538,N_2742);
nand U3448 (N_3448,N_2509,N_2676);
nand U3449 (N_3449,N_2573,N_2682);
or U3450 (N_3450,N_2670,N_2997);
nor U3451 (N_3451,N_2658,N_2900);
nand U3452 (N_3452,N_2823,N_2610);
nand U3453 (N_3453,N_2536,N_2625);
xor U3454 (N_3454,N_2899,N_2963);
nand U3455 (N_3455,N_2844,N_2877);
and U3456 (N_3456,N_2554,N_2803);
nor U3457 (N_3457,N_2996,N_2992);
nand U3458 (N_3458,N_2766,N_2980);
xor U3459 (N_3459,N_2930,N_2786);
or U3460 (N_3460,N_2736,N_2984);
or U3461 (N_3461,N_2950,N_2606);
xor U3462 (N_3462,N_2628,N_2828);
or U3463 (N_3463,N_2580,N_2581);
xnor U3464 (N_3464,N_2667,N_2606);
or U3465 (N_3465,N_2965,N_2523);
and U3466 (N_3466,N_2650,N_2826);
xnor U3467 (N_3467,N_2796,N_2759);
xor U3468 (N_3468,N_2584,N_2653);
nor U3469 (N_3469,N_2899,N_2810);
or U3470 (N_3470,N_2884,N_2607);
xnor U3471 (N_3471,N_2839,N_2926);
nor U3472 (N_3472,N_2954,N_2949);
or U3473 (N_3473,N_2795,N_2704);
and U3474 (N_3474,N_2704,N_2857);
nand U3475 (N_3475,N_2554,N_2760);
nand U3476 (N_3476,N_2707,N_2907);
or U3477 (N_3477,N_2510,N_2552);
xor U3478 (N_3478,N_2526,N_2813);
xnor U3479 (N_3479,N_2997,N_2986);
nand U3480 (N_3480,N_2580,N_2528);
or U3481 (N_3481,N_2924,N_2823);
xnor U3482 (N_3482,N_2976,N_2605);
nor U3483 (N_3483,N_2919,N_2670);
and U3484 (N_3484,N_2573,N_2905);
and U3485 (N_3485,N_2638,N_2691);
or U3486 (N_3486,N_2516,N_2852);
or U3487 (N_3487,N_2731,N_2998);
nand U3488 (N_3488,N_2711,N_2763);
xnor U3489 (N_3489,N_2609,N_2643);
xor U3490 (N_3490,N_2912,N_2589);
xor U3491 (N_3491,N_2958,N_2888);
nor U3492 (N_3492,N_2863,N_2616);
nand U3493 (N_3493,N_2685,N_2984);
or U3494 (N_3494,N_2829,N_2936);
and U3495 (N_3495,N_2666,N_2733);
and U3496 (N_3496,N_2702,N_2569);
nand U3497 (N_3497,N_2507,N_2795);
nor U3498 (N_3498,N_2719,N_2511);
xor U3499 (N_3499,N_2649,N_2769);
xnor U3500 (N_3500,N_3364,N_3374);
and U3501 (N_3501,N_3164,N_3330);
or U3502 (N_3502,N_3196,N_3241);
and U3503 (N_3503,N_3087,N_3111);
nand U3504 (N_3504,N_3098,N_3336);
nor U3505 (N_3505,N_3022,N_3274);
nand U3506 (N_3506,N_3074,N_3486);
nor U3507 (N_3507,N_3232,N_3358);
and U3508 (N_3508,N_3207,N_3032);
or U3509 (N_3509,N_3134,N_3491);
and U3510 (N_3510,N_3346,N_3165);
nand U3511 (N_3511,N_3193,N_3200);
nor U3512 (N_3512,N_3266,N_3126);
xor U3513 (N_3513,N_3009,N_3019);
nor U3514 (N_3514,N_3179,N_3391);
xor U3515 (N_3515,N_3464,N_3063);
or U3516 (N_3516,N_3268,N_3349);
and U3517 (N_3517,N_3414,N_3122);
and U3518 (N_3518,N_3112,N_3413);
xnor U3519 (N_3519,N_3119,N_3154);
xor U3520 (N_3520,N_3146,N_3497);
xor U3521 (N_3521,N_3451,N_3214);
xnor U3522 (N_3522,N_3075,N_3331);
nor U3523 (N_3523,N_3192,N_3294);
nor U3524 (N_3524,N_3013,N_3357);
nand U3525 (N_3525,N_3435,N_3334);
xnor U3526 (N_3526,N_3166,N_3162);
and U3527 (N_3527,N_3276,N_3113);
nand U3528 (N_3528,N_3024,N_3416);
or U3529 (N_3529,N_3237,N_3229);
nor U3530 (N_3530,N_3141,N_3296);
nor U3531 (N_3531,N_3107,N_3121);
and U3532 (N_3532,N_3204,N_3406);
nand U3533 (N_3533,N_3463,N_3493);
and U3534 (N_3534,N_3050,N_3350);
xnor U3535 (N_3535,N_3286,N_3040);
and U3536 (N_3536,N_3030,N_3360);
and U3537 (N_3537,N_3039,N_3475);
xor U3538 (N_3538,N_3084,N_3324);
nor U3539 (N_3539,N_3446,N_3295);
nor U3540 (N_3540,N_3407,N_3459);
nor U3541 (N_3541,N_3086,N_3395);
nand U3542 (N_3542,N_3474,N_3454);
xnor U3543 (N_3543,N_3436,N_3227);
nand U3544 (N_3544,N_3333,N_3014);
xnor U3545 (N_3545,N_3223,N_3428);
and U3546 (N_3546,N_3473,N_3423);
xor U3547 (N_3547,N_3230,N_3297);
nand U3548 (N_3548,N_3021,N_3219);
and U3549 (N_3549,N_3400,N_3234);
and U3550 (N_3550,N_3410,N_3145);
nor U3551 (N_3551,N_3258,N_3368);
xor U3552 (N_3552,N_3314,N_3054);
and U3553 (N_3553,N_3303,N_3338);
nand U3554 (N_3554,N_3081,N_3218);
xnor U3555 (N_3555,N_3137,N_3280);
nand U3556 (N_3556,N_3148,N_3259);
nor U3557 (N_3557,N_3199,N_3016);
nor U3558 (N_3558,N_3217,N_3434);
nor U3559 (N_3559,N_3092,N_3181);
nor U3560 (N_3560,N_3102,N_3109);
and U3561 (N_3561,N_3184,N_3382);
xnor U3562 (N_3562,N_3356,N_3370);
xnor U3563 (N_3563,N_3028,N_3305);
nor U3564 (N_3564,N_3208,N_3139);
nor U3565 (N_3565,N_3341,N_3490);
nor U3566 (N_3566,N_3495,N_3002);
nor U3567 (N_3567,N_3460,N_3053);
nor U3568 (N_3568,N_3328,N_3124);
nor U3569 (N_3569,N_3147,N_3479);
and U3570 (N_3570,N_3467,N_3004);
xnor U3571 (N_3571,N_3441,N_3047);
nor U3572 (N_3572,N_3096,N_3094);
and U3573 (N_3573,N_3290,N_3045);
nor U3574 (N_3574,N_3292,N_3299);
nor U3575 (N_3575,N_3221,N_3369);
xnor U3576 (N_3576,N_3345,N_3335);
nand U3577 (N_3577,N_3225,N_3197);
xnor U3578 (N_3578,N_3455,N_3373);
or U3579 (N_3579,N_3427,N_3038);
xnor U3580 (N_3580,N_3052,N_3355);
and U3581 (N_3581,N_3307,N_3452);
nand U3582 (N_3582,N_3066,N_3059);
nor U3583 (N_3583,N_3253,N_3178);
nor U3584 (N_3584,N_3317,N_3321);
and U3585 (N_3585,N_3211,N_3097);
nand U3586 (N_3586,N_3329,N_3320);
nor U3587 (N_3587,N_3070,N_3056);
nand U3588 (N_3588,N_3449,N_3213);
xor U3589 (N_3589,N_3309,N_3342);
xnor U3590 (N_3590,N_3037,N_3313);
xor U3591 (N_3591,N_3142,N_3186);
or U3592 (N_3592,N_3363,N_3224);
xor U3593 (N_3593,N_3120,N_3488);
nand U3594 (N_3594,N_3131,N_3017);
nor U3595 (N_3595,N_3380,N_3287);
xnor U3596 (N_3596,N_3362,N_3083);
xnor U3597 (N_3597,N_3477,N_3472);
xor U3598 (N_3598,N_3239,N_3228);
xnor U3599 (N_3599,N_3215,N_3171);
or U3600 (N_3600,N_3301,N_3461);
nand U3601 (N_3601,N_3319,N_3149);
xnor U3602 (N_3602,N_3457,N_3035);
or U3603 (N_3603,N_3379,N_3023);
nor U3604 (N_3604,N_3422,N_3409);
nand U3605 (N_3605,N_3240,N_3143);
xnor U3606 (N_3606,N_3318,N_3298);
nand U3607 (N_3607,N_3302,N_3062);
nand U3608 (N_3608,N_3496,N_3348);
xor U3609 (N_3609,N_3114,N_3392);
and U3610 (N_3610,N_3402,N_3271);
and U3611 (N_3611,N_3068,N_3169);
xor U3612 (N_3612,N_3442,N_3006);
xor U3613 (N_3613,N_3291,N_3123);
and U3614 (N_3614,N_3125,N_3383);
nand U3615 (N_3615,N_3426,N_3099);
or U3616 (N_3616,N_3265,N_3351);
nand U3617 (N_3617,N_3417,N_3150);
nand U3618 (N_3618,N_3007,N_3285);
nand U3619 (N_3619,N_3182,N_3160);
or U3620 (N_3620,N_3262,N_3484);
nand U3621 (N_3621,N_3337,N_3419);
or U3622 (N_3622,N_3263,N_3327);
or U3623 (N_3623,N_3482,N_3401);
and U3624 (N_3624,N_3140,N_3310);
nor U3625 (N_3625,N_3060,N_3105);
nor U3626 (N_3626,N_3172,N_3385);
or U3627 (N_3627,N_3210,N_3470);
xor U3628 (N_3628,N_3177,N_3389);
or U3629 (N_3629,N_3088,N_3072);
nor U3630 (N_3630,N_3079,N_3300);
or U3631 (N_3631,N_3010,N_3055);
xor U3632 (N_3632,N_3101,N_3384);
or U3633 (N_3633,N_3151,N_3026);
and U3634 (N_3634,N_3311,N_3043);
and U3635 (N_3635,N_3085,N_3403);
and U3636 (N_3636,N_3163,N_3250);
xnor U3637 (N_3637,N_3202,N_3339);
nand U3638 (N_3638,N_3306,N_3308);
nor U3639 (N_3639,N_3278,N_3432);
or U3640 (N_3640,N_3387,N_3071);
xor U3641 (N_3641,N_3439,N_3194);
and U3642 (N_3642,N_3458,N_3418);
and U3643 (N_3643,N_3051,N_3251);
or U3644 (N_3644,N_3393,N_3190);
and U3645 (N_3645,N_3279,N_3245);
nor U3646 (N_3646,N_3003,N_3275);
nor U3647 (N_3647,N_3222,N_3233);
xnor U3648 (N_3648,N_3077,N_3424);
nor U3649 (N_3649,N_3367,N_3246);
nand U3650 (N_3650,N_3359,N_3116);
xor U3651 (N_3651,N_3069,N_3332);
xnor U3652 (N_3652,N_3089,N_3156);
nand U3653 (N_3653,N_3153,N_3018);
nand U3654 (N_3654,N_3248,N_3483);
xor U3655 (N_3655,N_3343,N_3000);
and U3656 (N_3656,N_3183,N_3170);
xor U3657 (N_3657,N_3421,N_3191);
xor U3658 (N_3658,N_3205,N_3159);
nand U3659 (N_3659,N_3261,N_3462);
nand U3660 (N_3660,N_3133,N_3354);
or U3661 (N_3661,N_3315,N_3173);
and U3662 (N_3662,N_3492,N_3443);
nor U3663 (N_3663,N_3106,N_3008);
nor U3664 (N_3664,N_3438,N_3242);
and U3665 (N_3665,N_3236,N_3431);
xnor U3666 (N_3666,N_3203,N_3238);
and U3667 (N_3667,N_3381,N_3041);
nand U3668 (N_3668,N_3277,N_3243);
and U3669 (N_3669,N_3257,N_3188);
or U3670 (N_3670,N_3130,N_3256);
or U3671 (N_3671,N_3175,N_3405);
or U3672 (N_3672,N_3386,N_3174);
nor U3673 (N_3673,N_3005,N_3450);
and U3674 (N_3674,N_3076,N_3378);
xor U3675 (N_3675,N_3100,N_3377);
nand U3676 (N_3676,N_3167,N_3244);
nor U3677 (N_3677,N_3352,N_3394);
or U3678 (N_3678,N_3375,N_3272);
nor U3679 (N_3679,N_3110,N_3020);
or U3680 (N_3680,N_3091,N_3411);
xnor U3681 (N_3681,N_3058,N_3104);
nand U3682 (N_3682,N_3117,N_3231);
nor U3683 (N_3683,N_3361,N_3161);
nand U3684 (N_3684,N_3412,N_3185);
or U3685 (N_3685,N_3046,N_3408);
nor U3686 (N_3686,N_3304,N_3042);
and U3687 (N_3687,N_3015,N_3398);
and U3688 (N_3688,N_3235,N_3080);
or U3689 (N_3689,N_3078,N_3399);
or U3690 (N_3690,N_3425,N_3440);
nand U3691 (N_3691,N_3201,N_3312);
xnor U3692 (N_3692,N_3048,N_3049);
or U3693 (N_3693,N_3437,N_3136);
nand U3694 (N_3694,N_3034,N_3273);
or U3695 (N_3695,N_3453,N_3444);
nand U3696 (N_3696,N_3390,N_3445);
nor U3697 (N_3697,N_3415,N_3388);
nor U3698 (N_3698,N_3064,N_3353);
xnor U3699 (N_3699,N_3476,N_3430);
nor U3700 (N_3700,N_3264,N_3397);
nor U3701 (N_3701,N_3469,N_3249);
or U3702 (N_3702,N_3095,N_3176);
xor U3703 (N_3703,N_3220,N_3031);
xnor U3704 (N_3704,N_3025,N_3340);
and U3705 (N_3705,N_3326,N_3465);
or U3706 (N_3706,N_3157,N_3061);
and U3707 (N_3707,N_3322,N_3288);
or U3708 (N_3708,N_3158,N_3344);
xor U3709 (N_3709,N_3429,N_3082);
and U3710 (N_3710,N_3489,N_3471);
nand U3711 (N_3711,N_3293,N_3135);
or U3712 (N_3712,N_3138,N_3216);
or U3713 (N_3713,N_3093,N_3487);
xnor U3714 (N_3714,N_3283,N_3044);
xor U3715 (N_3715,N_3494,N_3067);
xnor U3716 (N_3716,N_3254,N_3212);
nand U3717 (N_3717,N_3270,N_3090);
and U3718 (N_3718,N_3115,N_3209);
nand U3719 (N_3719,N_3168,N_3001);
nor U3720 (N_3720,N_3057,N_3485);
nand U3721 (N_3721,N_3448,N_3481);
or U3722 (N_3722,N_3396,N_3012);
xor U3723 (N_3723,N_3247,N_3189);
or U3724 (N_3724,N_3198,N_3255);
nand U3725 (N_3725,N_3118,N_3128);
and U3726 (N_3726,N_3281,N_3371);
nand U3727 (N_3727,N_3466,N_3404);
and U3728 (N_3728,N_3260,N_3108);
nor U3729 (N_3729,N_3132,N_3468);
nor U3730 (N_3730,N_3187,N_3456);
nand U3731 (N_3731,N_3289,N_3129);
or U3732 (N_3732,N_3027,N_3029);
or U3733 (N_3733,N_3447,N_3366);
nand U3734 (N_3734,N_3252,N_3365);
or U3735 (N_3735,N_3267,N_3376);
nand U3736 (N_3736,N_3282,N_3073);
and U3737 (N_3737,N_3325,N_3323);
nand U3738 (N_3738,N_3269,N_3103);
or U3739 (N_3739,N_3226,N_3152);
or U3740 (N_3740,N_3011,N_3284);
or U3741 (N_3741,N_3127,N_3480);
nor U3742 (N_3742,N_3433,N_3316);
nand U3743 (N_3743,N_3478,N_3180);
xor U3744 (N_3744,N_3498,N_3144);
or U3745 (N_3745,N_3155,N_3347);
xor U3746 (N_3746,N_3033,N_3065);
xnor U3747 (N_3747,N_3036,N_3420);
nand U3748 (N_3748,N_3206,N_3195);
nand U3749 (N_3749,N_3372,N_3499);
nor U3750 (N_3750,N_3230,N_3409);
or U3751 (N_3751,N_3358,N_3472);
and U3752 (N_3752,N_3161,N_3465);
nand U3753 (N_3753,N_3104,N_3088);
nand U3754 (N_3754,N_3322,N_3353);
or U3755 (N_3755,N_3353,N_3094);
or U3756 (N_3756,N_3403,N_3412);
xor U3757 (N_3757,N_3104,N_3426);
nand U3758 (N_3758,N_3412,N_3059);
or U3759 (N_3759,N_3413,N_3152);
xnor U3760 (N_3760,N_3383,N_3490);
and U3761 (N_3761,N_3022,N_3161);
or U3762 (N_3762,N_3365,N_3140);
nand U3763 (N_3763,N_3434,N_3067);
nor U3764 (N_3764,N_3375,N_3261);
and U3765 (N_3765,N_3216,N_3331);
xor U3766 (N_3766,N_3294,N_3389);
and U3767 (N_3767,N_3199,N_3343);
xor U3768 (N_3768,N_3018,N_3376);
nand U3769 (N_3769,N_3299,N_3240);
nand U3770 (N_3770,N_3279,N_3368);
or U3771 (N_3771,N_3126,N_3201);
and U3772 (N_3772,N_3290,N_3243);
or U3773 (N_3773,N_3208,N_3025);
and U3774 (N_3774,N_3356,N_3130);
nor U3775 (N_3775,N_3166,N_3003);
or U3776 (N_3776,N_3221,N_3391);
or U3777 (N_3777,N_3393,N_3303);
nor U3778 (N_3778,N_3057,N_3315);
and U3779 (N_3779,N_3360,N_3070);
nand U3780 (N_3780,N_3058,N_3340);
xnor U3781 (N_3781,N_3241,N_3256);
or U3782 (N_3782,N_3190,N_3450);
nand U3783 (N_3783,N_3306,N_3396);
or U3784 (N_3784,N_3383,N_3007);
and U3785 (N_3785,N_3118,N_3482);
nor U3786 (N_3786,N_3027,N_3378);
nand U3787 (N_3787,N_3302,N_3110);
or U3788 (N_3788,N_3083,N_3099);
or U3789 (N_3789,N_3375,N_3426);
or U3790 (N_3790,N_3372,N_3439);
nand U3791 (N_3791,N_3137,N_3335);
nor U3792 (N_3792,N_3214,N_3391);
nand U3793 (N_3793,N_3171,N_3274);
or U3794 (N_3794,N_3180,N_3344);
nand U3795 (N_3795,N_3378,N_3322);
and U3796 (N_3796,N_3395,N_3309);
nand U3797 (N_3797,N_3121,N_3455);
xor U3798 (N_3798,N_3159,N_3495);
or U3799 (N_3799,N_3433,N_3449);
and U3800 (N_3800,N_3368,N_3013);
xnor U3801 (N_3801,N_3493,N_3189);
and U3802 (N_3802,N_3297,N_3098);
and U3803 (N_3803,N_3322,N_3196);
and U3804 (N_3804,N_3136,N_3292);
nand U3805 (N_3805,N_3348,N_3273);
or U3806 (N_3806,N_3232,N_3097);
nand U3807 (N_3807,N_3169,N_3473);
nand U3808 (N_3808,N_3087,N_3179);
or U3809 (N_3809,N_3078,N_3294);
and U3810 (N_3810,N_3042,N_3206);
xnor U3811 (N_3811,N_3326,N_3232);
and U3812 (N_3812,N_3245,N_3498);
or U3813 (N_3813,N_3255,N_3309);
xnor U3814 (N_3814,N_3423,N_3463);
and U3815 (N_3815,N_3312,N_3265);
nand U3816 (N_3816,N_3156,N_3188);
or U3817 (N_3817,N_3033,N_3425);
nor U3818 (N_3818,N_3036,N_3448);
nand U3819 (N_3819,N_3220,N_3455);
nor U3820 (N_3820,N_3492,N_3288);
nor U3821 (N_3821,N_3237,N_3408);
or U3822 (N_3822,N_3070,N_3247);
xor U3823 (N_3823,N_3124,N_3239);
or U3824 (N_3824,N_3312,N_3376);
nand U3825 (N_3825,N_3066,N_3365);
or U3826 (N_3826,N_3434,N_3252);
nor U3827 (N_3827,N_3021,N_3326);
nand U3828 (N_3828,N_3350,N_3418);
nor U3829 (N_3829,N_3033,N_3223);
nor U3830 (N_3830,N_3108,N_3076);
xor U3831 (N_3831,N_3113,N_3226);
nand U3832 (N_3832,N_3078,N_3498);
and U3833 (N_3833,N_3253,N_3361);
nand U3834 (N_3834,N_3294,N_3473);
nor U3835 (N_3835,N_3494,N_3155);
and U3836 (N_3836,N_3054,N_3082);
nand U3837 (N_3837,N_3206,N_3389);
nand U3838 (N_3838,N_3412,N_3426);
nand U3839 (N_3839,N_3312,N_3069);
or U3840 (N_3840,N_3374,N_3140);
and U3841 (N_3841,N_3237,N_3104);
or U3842 (N_3842,N_3015,N_3037);
nand U3843 (N_3843,N_3441,N_3380);
xor U3844 (N_3844,N_3008,N_3036);
and U3845 (N_3845,N_3301,N_3452);
nor U3846 (N_3846,N_3336,N_3323);
xnor U3847 (N_3847,N_3095,N_3161);
xor U3848 (N_3848,N_3093,N_3030);
and U3849 (N_3849,N_3423,N_3447);
nand U3850 (N_3850,N_3232,N_3387);
and U3851 (N_3851,N_3256,N_3109);
nor U3852 (N_3852,N_3325,N_3300);
nor U3853 (N_3853,N_3253,N_3096);
and U3854 (N_3854,N_3399,N_3089);
xor U3855 (N_3855,N_3348,N_3217);
nand U3856 (N_3856,N_3005,N_3247);
nand U3857 (N_3857,N_3168,N_3108);
xnor U3858 (N_3858,N_3237,N_3172);
nand U3859 (N_3859,N_3370,N_3093);
xor U3860 (N_3860,N_3125,N_3199);
or U3861 (N_3861,N_3196,N_3134);
xnor U3862 (N_3862,N_3423,N_3406);
nand U3863 (N_3863,N_3058,N_3103);
xnor U3864 (N_3864,N_3250,N_3325);
and U3865 (N_3865,N_3006,N_3389);
nor U3866 (N_3866,N_3055,N_3228);
or U3867 (N_3867,N_3018,N_3245);
xnor U3868 (N_3868,N_3009,N_3257);
nor U3869 (N_3869,N_3070,N_3067);
or U3870 (N_3870,N_3178,N_3015);
xor U3871 (N_3871,N_3197,N_3435);
xor U3872 (N_3872,N_3301,N_3446);
nor U3873 (N_3873,N_3267,N_3392);
and U3874 (N_3874,N_3100,N_3198);
and U3875 (N_3875,N_3364,N_3461);
xnor U3876 (N_3876,N_3346,N_3267);
xnor U3877 (N_3877,N_3202,N_3006);
or U3878 (N_3878,N_3073,N_3029);
nor U3879 (N_3879,N_3118,N_3071);
or U3880 (N_3880,N_3372,N_3058);
xor U3881 (N_3881,N_3473,N_3429);
nand U3882 (N_3882,N_3248,N_3262);
nor U3883 (N_3883,N_3415,N_3323);
nand U3884 (N_3884,N_3443,N_3106);
or U3885 (N_3885,N_3198,N_3022);
or U3886 (N_3886,N_3330,N_3236);
nand U3887 (N_3887,N_3371,N_3409);
nand U3888 (N_3888,N_3342,N_3297);
or U3889 (N_3889,N_3150,N_3315);
xor U3890 (N_3890,N_3118,N_3021);
and U3891 (N_3891,N_3247,N_3429);
xnor U3892 (N_3892,N_3081,N_3416);
nand U3893 (N_3893,N_3115,N_3360);
and U3894 (N_3894,N_3304,N_3181);
nor U3895 (N_3895,N_3385,N_3494);
nor U3896 (N_3896,N_3170,N_3199);
nand U3897 (N_3897,N_3499,N_3115);
and U3898 (N_3898,N_3253,N_3348);
xor U3899 (N_3899,N_3244,N_3329);
and U3900 (N_3900,N_3048,N_3103);
nor U3901 (N_3901,N_3485,N_3271);
nor U3902 (N_3902,N_3398,N_3051);
nand U3903 (N_3903,N_3414,N_3206);
xor U3904 (N_3904,N_3164,N_3235);
xor U3905 (N_3905,N_3260,N_3045);
xnor U3906 (N_3906,N_3333,N_3382);
nor U3907 (N_3907,N_3336,N_3012);
and U3908 (N_3908,N_3253,N_3353);
nor U3909 (N_3909,N_3056,N_3483);
and U3910 (N_3910,N_3356,N_3354);
xnor U3911 (N_3911,N_3361,N_3127);
xor U3912 (N_3912,N_3497,N_3367);
or U3913 (N_3913,N_3009,N_3466);
or U3914 (N_3914,N_3095,N_3172);
or U3915 (N_3915,N_3147,N_3245);
and U3916 (N_3916,N_3330,N_3424);
nand U3917 (N_3917,N_3492,N_3177);
nand U3918 (N_3918,N_3163,N_3275);
nand U3919 (N_3919,N_3444,N_3497);
nor U3920 (N_3920,N_3239,N_3332);
xor U3921 (N_3921,N_3134,N_3130);
nor U3922 (N_3922,N_3114,N_3385);
and U3923 (N_3923,N_3327,N_3273);
nand U3924 (N_3924,N_3301,N_3118);
nand U3925 (N_3925,N_3011,N_3066);
and U3926 (N_3926,N_3489,N_3286);
nand U3927 (N_3927,N_3381,N_3345);
and U3928 (N_3928,N_3442,N_3283);
nor U3929 (N_3929,N_3190,N_3230);
or U3930 (N_3930,N_3336,N_3321);
or U3931 (N_3931,N_3141,N_3173);
or U3932 (N_3932,N_3054,N_3002);
nand U3933 (N_3933,N_3346,N_3323);
or U3934 (N_3934,N_3084,N_3121);
xor U3935 (N_3935,N_3052,N_3472);
and U3936 (N_3936,N_3443,N_3132);
xor U3937 (N_3937,N_3248,N_3398);
nand U3938 (N_3938,N_3093,N_3451);
nor U3939 (N_3939,N_3406,N_3332);
or U3940 (N_3940,N_3441,N_3334);
nor U3941 (N_3941,N_3465,N_3156);
and U3942 (N_3942,N_3268,N_3369);
xor U3943 (N_3943,N_3300,N_3384);
nand U3944 (N_3944,N_3495,N_3287);
or U3945 (N_3945,N_3335,N_3393);
nand U3946 (N_3946,N_3130,N_3263);
nor U3947 (N_3947,N_3068,N_3273);
xor U3948 (N_3948,N_3107,N_3136);
nor U3949 (N_3949,N_3004,N_3291);
and U3950 (N_3950,N_3239,N_3378);
nand U3951 (N_3951,N_3373,N_3393);
xnor U3952 (N_3952,N_3431,N_3133);
and U3953 (N_3953,N_3404,N_3457);
nor U3954 (N_3954,N_3044,N_3279);
nand U3955 (N_3955,N_3407,N_3290);
nand U3956 (N_3956,N_3276,N_3129);
or U3957 (N_3957,N_3156,N_3371);
nor U3958 (N_3958,N_3308,N_3256);
and U3959 (N_3959,N_3280,N_3371);
nor U3960 (N_3960,N_3047,N_3162);
xnor U3961 (N_3961,N_3405,N_3427);
nor U3962 (N_3962,N_3215,N_3094);
nor U3963 (N_3963,N_3015,N_3418);
and U3964 (N_3964,N_3341,N_3194);
xnor U3965 (N_3965,N_3101,N_3122);
nor U3966 (N_3966,N_3310,N_3476);
xor U3967 (N_3967,N_3434,N_3388);
xnor U3968 (N_3968,N_3032,N_3133);
nor U3969 (N_3969,N_3273,N_3202);
or U3970 (N_3970,N_3252,N_3110);
or U3971 (N_3971,N_3396,N_3370);
xor U3972 (N_3972,N_3374,N_3125);
xnor U3973 (N_3973,N_3085,N_3151);
xnor U3974 (N_3974,N_3484,N_3410);
and U3975 (N_3975,N_3309,N_3169);
xnor U3976 (N_3976,N_3034,N_3021);
nand U3977 (N_3977,N_3462,N_3004);
nor U3978 (N_3978,N_3141,N_3054);
nor U3979 (N_3979,N_3476,N_3429);
xor U3980 (N_3980,N_3122,N_3396);
nor U3981 (N_3981,N_3074,N_3230);
and U3982 (N_3982,N_3315,N_3335);
and U3983 (N_3983,N_3491,N_3218);
nand U3984 (N_3984,N_3434,N_3166);
and U3985 (N_3985,N_3365,N_3185);
or U3986 (N_3986,N_3249,N_3376);
xor U3987 (N_3987,N_3267,N_3012);
xnor U3988 (N_3988,N_3367,N_3368);
xnor U3989 (N_3989,N_3072,N_3319);
nor U3990 (N_3990,N_3096,N_3341);
or U3991 (N_3991,N_3451,N_3253);
nand U3992 (N_3992,N_3028,N_3229);
nor U3993 (N_3993,N_3486,N_3301);
or U3994 (N_3994,N_3242,N_3173);
or U3995 (N_3995,N_3326,N_3369);
nand U3996 (N_3996,N_3014,N_3456);
and U3997 (N_3997,N_3001,N_3173);
or U3998 (N_3998,N_3407,N_3479);
nand U3999 (N_3999,N_3287,N_3058);
or U4000 (N_4000,N_3501,N_3948);
or U4001 (N_4001,N_3872,N_3694);
xnor U4002 (N_4002,N_3550,N_3805);
nand U4003 (N_4003,N_3749,N_3963);
nor U4004 (N_4004,N_3651,N_3785);
nor U4005 (N_4005,N_3896,N_3610);
nor U4006 (N_4006,N_3628,N_3953);
nand U4007 (N_4007,N_3995,N_3833);
nor U4008 (N_4008,N_3835,N_3546);
and U4009 (N_4009,N_3851,N_3516);
and U4010 (N_4010,N_3678,N_3685);
nand U4011 (N_4011,N_3912,N_3656);
nand U4012 (N_4012,N_3968,N_3765);
xor U4013 (N_4013,N_3727,N_3775);
and U4014 (N_4014,N_3604,N_3873);
nor U4015 (N_4015,N_3630,N_3665);
nor U4016 (N_4016,N_3574,N_3876);
nor U4017 (N_4017,N_3752,N_3527);
nor U4018 (N_4018,N_3682,N_3780);
nor U4019 (N_4019,N_3809,N_3684);
and U4020 (N_4020,N_3571,N_3850);
nor U4021 (N_4021,N_3657,N_3987);
xnor U4022 (N_4022,N_3523,N_3594);
nand U4023 (N_4023,N_3695,N_3741);
and U4024 (N_4024,N_3888,N_3794);
nor U4025 (N_4025,N_3900,N_3869);
xnor U4026 (N_4026,N_3577,N_3878);
or U4027 (N_4027,N_3757,N_3843);
nand U4028 (N_4028,N_3822,N_3629);
nand U4029 (N_4029,N_3999,N_3803);
nor U4030 (N_4030,N_3553,N_3773);
nand U4031 (N_4031,N_3790,N_3668);
nor U4032 (N_4032,N_3838,N_3725);
xor U4033 (N_4033,N_3856,N_3735);
nor U4034 (N_4034,N_3680,N_3811);
nor U4035 (N_4035,N_3880,N_3903);
nor U4036 (N_4036,N_3959,N_3631);
and U4037 (N_4037,N_3861,N_3864);
nand U4038 (N_4038,N_3638,N_3879);
or U4039 (N_4039,N_3881,N_3917);
xnor U4040 (N_4040,N_3992,N_3931);
xnor U4041 (N_4041,N_3793,N_3619);
and U4042 (N_4042,N_3672,N_3579);
nand U4043 (N_4043,N_3715,N_3890);
or U4044 (N_4044,N_3994,N_3905);
or U4045 (N_4045,N_3940,N_3556);
xor U4046 (N_4046,N_3731,N_3690);
and U4047 (N_4047,N_3918,N_3595);
or U4048 (N_4048,N_3598,N_3836);
and U4049 (N_4049,N_3744,N_3808);
nor U4050 (N_4050,N_3576,N_3691);
xnor U4051 (N_4051,N_3779,N_3892);
and U4052 (N_4052,N_3935,N_3828);
xnor U4053 (N_4053,N_3600,N_3841);
and U4054 (N_4054,N_3602,N_3711);
xor U4055 (N_4055,N_3804,N_3558);
nor U4056 (N_4056,N_3853,N_3966);
xor U4057 (N_4057,N_3519,N_3818);
or U4058 (N_4058,N_3789,N_3743);
nor U4059 (N_4059,N_3531,N_3732);
nor U4060 (N_4060,N_3875,N_3842);
nand U4061 (N_4061,N_3667,N_3588);
xnor U4062 (N_4062,N_3988,N_3518);
nand U4063 (N_4063,N_3693,N_3521);
xor U4064 (N_4064,N_3816,N_3946);
nand U4065 (N_4065,N_3502,N_3812);
nor U4066 (N_4066,N_3707,N_3884);
and U4067 (N_4067,N_3647,N_3777);
and U4068 (N_4068,N_3973,N_3740);
and U4069 (N_4069,N_3887,N_3754);
nand U4070 (N_4070,N_3768,N_3990);
nor U4071 (N_4071,N_3825,N_3541);
and U4072 (N_4072,N_3526,N_3854);
or U4073 (N_4073,N_3852,N_3616);
and U4074 (N_4074,N_3522,N_3700);
nand U4075 (N_4075,N_3986,N_3882);
nand U4076 (N_4076,N_3596,N_3955);
nor U4077 (N_4077,N_3625,N_3747);
and U4078 (N_4078,N_3923,N_3704);
or U4079 (N_4079,N_3671,N_3956);
and U4080 (N_4080,N_3593,N_3559);
nor U4081 (N_4081,N_3507,N_3834);
xor U4082 (N_4082,N_3796,N_3542);
nand U4083 (N_4083,N_3951,N_3589);
nand U4084 (N_4084,N_3952,N_3860);
nand U4085 (N_4085,N_3839,N_3958);
nor U4086 (N_4086,N_3899,N_3746);
and U4087 (N_4087,N_3549,N_3907);
nand U4088 (N_4088,N_3617,N_3670);
nand U4089 (N_4089,N_3554,N_3934);
xor U4090 (N_4090,N_3814,N_3837);
nor U4091 (N_4091,N_3911,N_3646);
xor U4092 (N_4092,N_3795,N_3883);
nand U4093 (N_4093,N_3538,N_3991);
or U4094 (N_4094,N_3632,N_3648);
nor U4095 (N_4095,N_3664,N_3904);
nand U4096 (N_4096,N_3915,N_3524);
nand U4097 (N_4097,N_3535,N_3705);
nand U4098 (N_4098,N_3967,N_3712);
xnor U4099 (N_4099,N_3797,N_3548);
or U4100 (N_4100,N_3784,N_3761);
nand U4101 (N_4101,N_3925,N_3529);
and U4102 (N_4102,N_3792,N_3969);
and U4103 (N_4103,N_3563,N_3960);
xor U4104 (N_4104,N_3800,N_3644);
nor U4105 (N_4105,N_3929,N_3573);
or U4106 (N_4106,N_3738,N_3511);
and U4107 (N_4107,N_3788,N_3688);
nor U4108 (N_4108,N_3945,N_3512);
and U4109 (N_4109,N_3654,N_3659);
nor U4110 (N_4110,N_3823,N_3802);
xnor U4111 (N_4111,N_3916,N_3720);
or U4112 (N_4112,N_3871,N_3620);
xor U4113 (N_4113,N_3846,N_3640);
or U4114 (N_4114,N_3635,N_3643);
or U4115 (N_4115,N_3555,N_3626);
nand U4116 (N_4116,N_3980,N_3742);
and U4117 (N_4117,N_3791,N_3655);
or U4118 (N_4118,N_3599,N_3772);
xor U4119 (N_4119,N_3893,N_3520);
and U4120 (N_4120,N_3636,N_3939);
xor U4121 (N_4121,N_3862,N_3806);
and U4122 (N_4122,N_3503,N_3639);
xnor U4123 (N_4123,N_3763,N_3957);
or U4124 (N_4124,N_3504,N_3962);
xnor U4125 (N_4125,N_3847,N_3611);
nor U4126 (N_4126,N_3983,N_3622);
xnor U4127 (N_4127,N_3745,N_3859);
and U4128 (N_4128,N_3820,N_3982);
or U4129 (N_4129,N_3845,N_3927);
or U4130 (N_4130,N_3545,N_3509);
nor U4131 (N_4131,N_3815,N_3702);
or U4132 (N_4132,N_3585,N_3714);
and U4133 (N_4133,N_3947,N_3783);
nand U4134 (N_4134,N_3551,N_3724);
nor U4135 (N_4135,N_3584,N_3965);
or U4136 (N_4136,N_3920,N_3674);
nor U4137 (N_4137,N_3798,N_3567);
nor U4138 (N_4138,N_3832,N_3698);
and U4139 (N_4139,N_3561,N_3943);
nor U4140 (N_4140,N_3606,N_3645);
or U4141 (N_4141,N_3889,N_3985);
nor U4142 (N_4142,N_3539,N_3621);
xnor U4143 (N_4143,N_3897,N_3591);
or U4144 (N_4144,N_3612,N_3762);
nor U4145 (N_4145,N_3544,N_3902);
xor U4146 (N_4146,N_3592,N_3716);
xor U4147 (N_4147,N_3649,N_3997);
and U4148 (N_4148,N_3569,N_3717);
and U4149 (N_4149,N_3696,N_3575);
nand U4150 (N_4150,N_3865,N_3572);
and U4151 (N_4151,N_3801,N_3613);
nand U4152 (N_4152,N_3863,N_3623);
and U4153 (N_4153,N_3901,N_3739);
xor U4154 (N_4154,N_3660,N_3689);
and U4155 (N_4155,N_3510,N_3683);
xor U4156 (N_4156,N_3528,N_3874);
nand U4157 (N_4157,N_3870,N_3508);
xor U4158 (N_4158,N_3505,N_3867);
nand U4159 (N_4159,N_3910,N_3857);
nand U4160 (N_4160,N_3827,N_3998);
or U4161 (N_4161,N_3937,N_3637);
and U4162 (N_4162,N_3760,N_3642);
or U4163 (N_4163,N_3517,N_3970);
xor U4164 (N_4164,N_3961,N_3941);
nand U4165 (N_4165,N_3663,N_3766);
nand U4166 (N_4166,N_3755,N_3580);
or U4167 (N_4167,N_3938,N_3774);
and U4168 (N_4168,N_3650,N_3891);
nor U4169 (N_4169,N_3547,N_3721);
and U4170 (N_4170,N_3676,N_3587);
nand U4171 (N_4171,N_3877,N_3679);
nor U4172 (N_4172,N_3566,N_3624);
xnor U4173 (N_4173,N_3767,N_3607);
or U4174 (N_4174,N_3618,N_3608);
and U4175 (N_4175,N_3787,N_3532);
xnor U4176 (N_4176,N_3949,N_3758);
or U4177 (N_4177,N_3954,N_3866);
nor U4178 (N_4178,N_3933,N_3984);
nor U4179 (N_4179,N_3964,N_3906);
xnor U4180 (N_4180,N_3719,N_3898);
nand U4181 (N_4181,N_3776,N_3681);
or U4182 (N_4182,N_3979,N_3615);
nor U4183 (N_4183,N_3855,N_3686);
xnor U4184 (N_4184,N_3936,N_3560);
nor U4185 (N_4185,N_3942,N_3653);
and U4186 (N_4186,N_3733,N_3971);
or U4187 (N_4187,N_3930,N_3848);
and U4188 (N_4188,N_3753,N_3540);
or U4189 (N_4189,N_3993,N_3652);
and U4190 (N_4190,N_3662,N_3661);
xor U4191 (N_4191,N_3978,N_3533);
and U4192 (N_4192,N_3976,N_3722);
and U4193 (N_4193,N_3819,N_3736);
nor U4194 (N_4194,N_3677,N_3675);
or U4195 (N_4195,N_3737,N_3759);
nor U4196 (N_4196,N_3778,N_3543);
xnor U4197 (N_4197,N_3534,N_3692);
nand U4198 (N_4198,N_3666,N_3868);
xor U4199 (N_4199,N_3603,N_3728);
nor U4200 (N_4200,N_3633,N_3515);
and U4201 (N_4201,N_3748,N_3530);
and U4202 (N_4202,N_3718,N_3981);
xor U4203 (N_4203,N_3919,N_3597);
and U4204 (N_4204,N_3886,N_3996);
nand U4205 (N_4205,N_3500,N_3977);
nor U4206 (N_4206,N_3706,N_3817);
nand U4207 (N_4207,N_3989,N_3909);
xor U4208 (N_4208,N_3770,N_3729);
or U4209 (N_4209,N_3926,N_3627);
nand U4210 (N_4210,N_3914,N_3756);
nor U4211 (N_4211,N_3703,N_3751);
nand U4212 (N_4212,N_3565,N_3582);
or U4213 (N_4213,N_3974,N_3726);
nor U4214 (N_4214,N_3568,N_3713);
xnor U4215 (N_4215,N_3641,N_3858);
or U4216 (N_4216,N_3932,N_3781);
xnor U4217 (N_4217,N_3849,N_3506);
nand U4218 (N_4218,N_3697,N_3699);
nand U4219 (N_4219,N_3924,N_3922);
xnor U4220 (N_4220,N_3583,N_3614);
or U4221 (N_4221,N_3764,N_3605);
xnor U4222 (N_4222,N_3821,N_3813);
xnor U4223 (N_4223,N_3710,N_3514);
xnor U4224 (N_4224,N_3885,N_3944);
or U4225 (N_4225,N_3552,N_3824);
and U4226 (N_4226,N_3921,N_3840);
nor U4227 (N_4227,N_3709,N_3830);
and U4228 (N_4228,N_3769,N_3972);
nor U4229 (N_4229,N_3826,N_3895);
or U4230 (N_4230,N_3590,N_3734);
xnor U4231 (N_4231,N_3687,N_3829);
or U4232 (N_4232,N_3525,N_3564);
xnor U4233 (N_4233,N_3908,N_3658);
and U4234 (N_4234,N_3750,N_3537);
nand U4235 (N_4235,N_3844,N_3581);
nand U4236 (N_4236,N_3786,N_3562);
nor U4237 (N_4237,N_3634,N_3701);
nand U4238 (N_4238,N_3782,N_3913);
nand U4239 (N_4239,N_3669,N_3723);
xor U4240 (N_4240,N_3578,N_3799);
nand U4241 (N_4241,N_3810,N_3975);
nand U4242 (N_4242,N_3708,N_3894);
xor U4243 (N_4243,N_3609,N_3570);
or U4244 (N_4244,N_3586,N_3928);
nand U4245 (N_4245,N_3950,N_3831);
or U4246 (N_4246,N_3536,N_3771);
or U4247 (N_4247,N_3673,N_3807);
nor U4248 (N_4248,N_3730,N_3557);
nand U4249 (N_4249,N_3513,N_3601);
or U4250 (N_4250,N_3798,N_3840);
nand U4251 (N_4251,N_3749,N_3973);
nand U4252 (N_4252,N_3855,N_3545);
and U4253 (N_4253,N_3929,N_3741);
and U4254 (N_4254,N_3947,N_3956);
nand U4255 (N_4255,N_3886,N_3677);
nor U4256 (N_4256,N_3902,N_3727);
nand U4257 (N_4257,N_3736,N_3599);
nor U4258 (N_4258,N_3500,N_3975);
xor U4259 (N_4259,N_3584,N_3731);
and U4260 (N_4260,N_3829,N_3782);
or U4261 (N_4261,N_3669,N_3757);
nor U4262 (N_4262,N_3677,N_3529);
nand U4263 (N_4263,N_3892,N_3999);
and U4264 (N_4264,N_3975,N_3768);
xnor U4265 (N_4265,N_3578,N_3961);
xnor U4266 (N_4266,N_3673,N_3832);
xor U4267 (N_4267,N_3948,N_3521);
or U4268 (N_4268,N_3642,N_3990);
nand U4269 (N_4269,N_3918,N_3924);
xnor U4270 (N_4270,N_3903,N_3813);
xor U4271 (N_4271,N_3962,N_3858);
nor U4272 (N_4272,N_3713,N_3957);
nand U4273 (N_4273,N_3835,N_3598);
nand U4274 (N_4274,N_3983,N_3649);
xor U4275 (N_4275,N_3864,N_3897);
nor U4276 (N_4276,N_3949,N_3942);
nand U4277 (N_4277,N_3962,N_3691);
and U4278 (N_4278,N_3885,N_3508);
or U4279 (N_4279,N_3846,N_3767);
nor U4280 (N_4280,N_3642,N_3998);
xnor U4281 (N_4281,N_3673,N_3702);
nand U4282 (N_4282,N_3914,N_3992);
nor U4283 (N_4283,N_3923,N_3569);
nor U4284 (N_4284,N_3671,N_3988);
xor U4285 (N_4285,N_3587,N_3920);
xor U4286 (N_4286,N_3971,N_3672);
and U4287 (N_4287,N_3863,N_3963);
xnor U4288 (N_4288,N_3688,N_3863);
nor U4289 (N_4289,N_3723,N_3502);
nand U4290 (N_4290,N_3745,N_3720);
xnor U4291 (N_4291,N_3507,N_3746);
nand U4292 (N_4292,N_3971,N_3885);
xnor U4293 (N_4293,N_3728,N_3597);
xor U4294 (N_4294,N_3835,N_3686);
nor U4295 (N_4295,N_3680,N_3748);
nand U4296 (N_4296,N_3717,N_3770);
xor U4297 (N_4297,N_3714,N_3591);
nor U4298 (N_4298,N_3869,N_3899);
nand U4299 (N_4299,N_3769,N_3977);
nand U4300 (N_4300,N_3601,N_3588);
nand U4301 (N_4301,N_3641,N_3601);
nor U4302 (N_4302,N_3757,N_3501);
nor U4303 (N_4303,N_3663,N_3974);
or U4304 (N_4304,N_3525,N_3663);
or U4305 (N_4305,N_3926,N_3978);
nor U4306 (N_4306,N_3889,N_3801);
xor U4307 (N_4307,N_3688,N_3964);
nand U4308 (N_4308,N_3740,N_3595);
and U4309 (N_4309,N_3959,N_3979);
and U4310 (N_4310,N_3910,N_3884);
and U4311 (N_4311,N_3690,N_3873);
xnor U4312 (N_4312,N_3854,N_3830);
nand U4313 (N_4313,N_3706,N_3584);
nor U4314 (N_4314,N_3836,N_3888);
or U4315 (N_4315,N_3780,N_3700);
nand U4316 (N_4316,N_3862,N_3920);
or U4317 (N_4317,N_3895,N_3630);
nor U4318 (N_4318,N_3753,N_3903);
nor U4319 (N_4319,N_3974,N_3658);
nor U4320 (N_4320,N_3975,N_3619);
and U4321 (N_4321,N_3687,N_3926);
and U4322 (N_4322,N_3734,N_3645);
nand U4323 (N_4323,N_3939,N_3988);
xor U4324 (N_4324,N_3640,N_3993);
nand U4325 (N_4325,N_3845,N_3533);
or U4326 (N_4326,N_3917,N_3798);
or U4327 (N_4327,N_3589,N_3502);
nand U4328 (N_4328,N_3558,N_3627);
nand U4329 (N_4329,N_3673,N_3548);
and U4330 (N_4330,N_3588,N_3914);
xnor U4331 (N_4331,N_3851,N_3652);
or U4332 (N_4332,N_3699,N_3920);
nor U4333 (N_4333,N_3912,N_3849);
xor U4334 (N_4334,N_3600,N_3509);
and U4335 (N_4335,N_3801,N_3947);
xor U4336 (N_4336,N_3792,N_3636);
or U4337 (N_4337,N_3966,N_3804);
xor U4338 (N_4338,N_3893,N_3505);
or U4339 (N_4339,N_3829,N_3732);
xnor U4340 (N_4340,N_3725,N_3966);
nor U4341 (N_4341,N_3971,N_3860);
nor U4342 (N_4342,N_3876,N_3618);
nand U4343 (N_4343,N_3787,N_3732);
and U4344 (N_4344,N_3896,N_3686);
xor U4345 (N_4345,N_3851,N_3767);
nand U4346 (N_4346,N_3739,N_3852);
nor U4347 (N_4347,N_3626,N_3595);
and U4348 (N_4348,N_3950,N_3719);
nor U4349 (N_4349,N_3529,N_3657);
nand U4350 (N_4350,N_3762,N_3841);
or U4351 (N_4351,N_3729,N_3885);
nor U4352 (N_4352,N_3849,N_3702);
nand U4353 (N_4353,N_3596,N_3601);
nand U4354 (N_4354,N_3593,N_3972);
or U4355 (N_4355,N_3930,N_3810);
nand U4356 (N_4356,N_3981,N_3922);
or U4357 (N_4357,N_3891,N_3976);
or U4358 (N_4358,N_3953,N_3688);
nor U4359 (N_4359,N_3640,N_3501);
and U4360 (N_4360,N_3787,N_3748);
xnor U4361 (N_4361,N_3997,N_3803);
and U4362 (N_4362,N_3674,N_3763);
nand U4363 (N_4363,N_3877,N_3704);
xnor U4364 (N_4364,N_3775,N_3585);
or U4365 (N_4365,N_3719,N_3800);
xor U4366 (N_4366,N_3961,N_3991);
and U4367 (N_4367,N_3799,N_3608);
and U4368 (N_4368,N_3525,N_3693);
nand U4369 (N_4369,N_3656,N_3580);
nor U4370 (N_4370,N_3735,N_3758);
nand U4371 (N_4371,N_3641,N_3864);
or U4372 (N_4372,N_3741,N_3921);
or U4373 (N_4373,N_3512,N_3898);
nand U4374 (N_4374,N_3714,N_3967);
and U4375 (N_4375,N_3551,N_3832);
nor U4376 (N_4376,N_3992,N_3835);
or U4377 (N_4377,N_3822,N_3764);
or U4378 (N_4378,N_3606,N_3921);
xor U4379 (N_4379,N_3657,N_3696);
nor U4380 (N_4380,N_3528,N_3633);
or U4381 (N_4381,N_3511,N_3882);
and U4382 (N_4382,N_3746,N_3559);
and U4383 (N_4383,N_3596,N_3981);
nor U4384 (N_4384,N_3662,N_3983);
and U4385 (N_4385,N_3656,N_3693);
xnor U4386 (N_4386,N_3841,N_3627);
nor U4387 (N_4387,N_3726,N_3605);
or U4388 (N_4388,N_3980,N_3942);
or U4389 (N_4389,N_3918,N_3945);
xor U4390 (N_4390,N_3517,N_3857);
nand U4391 (N_4391,N_3585,N_3547);
xnor U4392 (N_4392,N_3601,N_3811);
nor U4393 (N_4393,N_3820,N_3594);
nand U4394 (N_4394,N_3866,N_3992);
and U4395 (N_4395,N_3699,N_3872);
and U4396 (N_4396,N_3902,N_3752);
and U4397 (N_4397,N_3862,N_3930);
nor U4398 (N_4398,N_3724,N_3887);
and U4399 (N_4399,N_3786,N_3884);
or U4400 (N_4400,N_3748,N_3870);
nor U4401 (N_4401,N_3667,N_3706);
nand U4402 (N_4402,N_3887,N_3661);
or U4403 (N_4403,N_3748,N_3791);
and U4404 (N_4404,N_3849,N_3766);
nand U4405 (N_4405,N_3532,N_3666);
and U4406 (N_4406,N_3709,N_3595);
and U4407 (N_4407,N_3801,N_3535);
nand U4408 (N_4408,N_3721,N_3715);
or U4409 (N_4409,N_3967,N_3613);
or U4410 (N_4410,N_3986,N_3982);
nor U4411 (N_4411,N_3996,N_3979);
xnor U4412 (N_4412,N_3777,N_3527);
xnor U4413 (N_4413,N_3988,N_3729);
xor U4414 (N_4414,N_3615,N_3951);
or U4415 (N_4415,N_3910,N_3899);
or U4416 (N_4416,N_3619,N_3849);
or U4417 (N_4417,N_3733,N_3668);
nor U4418 (N_4418,N_3607,N_3985);
or U4419 (N_4419,N_3934,N_3930);
nor U4420 (N_4420,N_3741,N_3709);
xor U4421 (N_4421,N_3782,N_3996);
nor U4422 (N_4422,N_3564,N_3974);
nand U4423 (N_4423,N_3782,N_3824);
nand U4424 (N_4424,N_3938,N_3999);
and U4425 (N_4425,N_3909,N_3743);
xor U4426 (N_4426,N_3990,N_3773);
nor U4427 (N_4427,N_3836,N_3663);
and U4428 (N_4428,N_3920,N_3822);
and U4429 (N_4429,N_3777,N_3520);
and U4430 (N_4430,N_3761,N_3764);
nand U4431 (N_4431,N_3589,N_3870);
nor U4432 (N_4432,N_3573,N_3530);
xnor U4433 (N_4433,N_3703,N_3501);
xor U4434 (N_4434,N_3778,N_3852);
or U4435 (N_4435,N_3916,N_3565);
or U4436 (N_4436,N_3721,N_3699);
nor U4437 (N_4437,N_3652,N_3507);
xnor U4438 (N_4438,N_3779,N_3588);
and U4439 (N_4439,N_3812,N_3864);
or U4440 (N_4440,N_3820,N_3677);
or U4441 (N_4441,N_3536,N_3917);
and U4442 (N_4442,N_3880,N_3683);
nand U4443 (N_4443,N_3771,N_3515);
xnor U4444 (N_4444,N_3685,N_3645);
or U4445 (N_4445,N_3678,N_3753);
or U4446 (N_4446,N_3812,N_3979);
xor U4447 (N_4447,N_3727,N_3834);
nand U4448 (N_4448,N_3852,N_3889);
and U4449 (N_4449,N_3969,N_3602);
and U4450 (N_4450,N_3650,N_3589);
xnor U4451 (N_4451,N_3926,N_3593);
and U4452 (N_4452,N_3948,N_3747);
or U4453 (N_4453,N_3924,N_3675);
or U4454 (N_4454,N_3804,N_3958);
nand U4455 (N_4455,N_3585,N_3969);
nand U4456 (N_4456,N_3673,N_3681);
nand U4457 (N_4457,N_3810,N_3676);
nor U4458 (N_4458,N_3891,N_3705);
and U4459 (N_4459,N_3643,N_3554);
nand U4460 (N_4460,N_3855,N_3724);
xnor U4461 (N_4461,N_3580,N_3967);
or U4462 (N_4462,N_3536,N_3960);
nor U4463 (N_4463,N_3842,N_3622);
nor U4464 (N_4464,N_3914,N_3535);
nor U4465 (N_4465,N_3513,N_3857);
xor U4466 (N_4466,N_3555,N_3596);
or U4467 (N_4467,N_3541,N_3747);
nand U4468 (N_4468,N_3833,N_3929);
nor U4469 (N_4469,N_3899,N_3636);
nor U4470 (N_4470,N_3878,N_3600);
nand U4471 (N_4471,N_3708,N_3648);
nor U4472 (N_4472,N_3905,N_3722);
nor U4473 (N_4473,N_3843,N_3890);
xnor U4474 (N_4474,N_3765,N_3548);
and U4475 (N_4475,N_3983,N_3539);
nand U4476 (N_4476,N_3896,N_3693);
nor U4477 (N_4477,N_3508,N_3995);
xor U4478 (N_4478,N_3808,N_3900);
nor U4479 (N_4479,N_3765,N_3600);
and U4480 (N_4480,N_3926,N_3748);
or U4481 (N_4481,N_3573,N_3950);
or U4482 (N_4482,N_3892,N_3784);
nand U4483 (N_4483,N_3795,N_3914);
nor U4484 (N_4484,N_3693,N_3998);
nand U4485 (N_4485,N_3543,N_3668);
xnor U4486 (N_4486,N_3883,N_3860);
xnor U4487 (N_4487,N_3911,N_3661);
or U4488 (N_4488,N_3776,N_3911);
and U4489 (N_4489,N_3883,N_3662);
and U4490 (N_4490,N_3524,N_3672);
nand U4491 (N_4491,N_3735,N_3535);
nand U4492 (N_4492,N_3737,N_3763);
nand U4493 (N_4493,N_3524,N_3831);
xor U4494 (N_4494,N_3524,N_3640);
or U4495 (N_4495,N_3749,N_3793);
nand U4496 (N_4496,N_3937,N_3516);
xnor U4497 (N_4497,N_3669,N_3623);
or U4498 (N_4498,N_3668,N_3851);
xnor U4499 (N_4499,N_3785,N_3927);
xor U4500 (N_4500,N_4053,N_4241);
nand U4501 (N_4501,N_4339,N_4215);
xor U4502 (N_4502,N_4125,N_4432);
xor U4503 (N_4503,N_4165,N_4128);
or U4504 (N_4504,N_4462,N_4039);
nand U4505 (N_4505,N_4275,N_4299);
nand U4506 (N_4506,N_4461,N_4109);
and U4507 (N_4507,N_4146,N_4400);
nor U4508 (N_4508,N_4218,N_4315);
and U4509 (N_4509,N_4176,N_4269);
nand U4510 (N_4510,N_4348,N_4197);
or U4511 (N_4511,N_4494,N_4173);
xor U4512 (N_4512,N_4338,N_4119);
and U4513 (N_4513,N_4496,N_4464);
or U4514 (N_4514,N_4322,N_4105);
and U4515 (N_4515,N_4291,N_4435);
xor U4516 (N_4516,N_4442,N_4476);
and U4517 (N_4517,N_4074,N_4472);
nand U4518 (N_4518,N_4025,N_4304);
nand U4519 (N_4519,N_4305,N_4356);
and U4520 (N_4520,N_4045,N_4179);
nor U4521 (N_4521,N_4307,N_4018);
or U4522 (N_4522,N_4080,N_4183);
nor U4523 (N_4523,N_4365,N_4450);
nor U4524 (N_4524,N_4187,N_4216);
and U4525 (N_4525,N_4298,N_4444);
and U4526 (N_4526,N_4401,N_4290);
nand U4527 (N_4527,N_4376,N_4051);
xor U4528 (N_4528,N_4387,N_4182);
nor U4529 (N_4529,N_4482,N_4029);
nor U4530 (N_4530,N_4005,N_4085);
nand U4531 (N_4531,N_4204,N_4301);
nor U4532 (N_4532,N_4255,N_4424);
xnor U4533 (N_4533,N_4416,N_4200);
xnor U4534 (N_4534,N_4433,N_4309);
nor U4535 (N_4535,N_4156,N_4382);
nand U4536 (N_4536,N_4224,N_4420);
xor U4537 (N_4537,N_4266,N_4172);
nand U4538 (N_4538,N_4055,N_4280);
nor U4539 (N_4539,N_4478,N_4016);
nor U4540 (N_4540,N_4340,N_4064);
xor U4541 (N_4541,N_4415,N_4405);
nor U4542 (N_4542,N_4486,N_4363);
xnor U4543 (N_4543,N_4078,N_4288);
or U4544 (N_4544,N_4246,N_4075);
xor U4545 (N_4545,N_4271,N_4487);
or U4546 (N_4546,N_4161,N_4135);
xnor U4547 (N_4547,N_4122,N_4113);
xnor U4548 (N_4548,N_4419,N_4274);
and U4549 (N_4549,N_4004,N_4091);
xnor U4550 (N_4550,N_4093,N_4495);
xnor U4551 (N_4551,N_4023,N_4098);
nor U4552 (N_4552,N_4196,N_4333);
or U4553 (N_4553,N_4010,N_4422);
nand U4554 (N_4554,N_4430,N_4431);
or U4555 (N_4555,N_4465,N_4072);
xnor U4556 (N_4556,N_4469,N_4167);
xnor U4557 (N_4557,N_4151,N_4483);
and U4558 (N_4558,N_4263,N_4059);
nor U4559 (N_4559,N_4367,N_4492);
nand U4560 (N_4560,N_4355,N_4398);
or U4561 (N_4561,N_4017,N_4238);
xor U4562 (N_4562,N_4047,N_4297);
nor U4563 (N_4563,N_4272,N_4243);
or U4564 (N_4564,N_4493,N_4032);
nand U4565 (N_4565,N_4295,N_4049);
or U4566 (N_4566,N_4421,N_4330);
or U4567 (N_4567,N_4323,N_4068);
xnor U4568 (N_4568,N_4357,N_4199);
or U4569 (N_4569,N_4079,N_4184);
or U4570 (N_4570,N_4012,N_4067);
xor U4571 (N_4571,N_4203,N_4043);
nand U4572 (N_4572,N_4250,N_4396);
or U4573 (N_4573,N_4285,N_4436);
or U4574 (N_4574,N_4201,N_4477);
and U4575 (N_4575,N_4437,N_4115);
nand U4576 (N_4576,N_4058,N_4256);
or U4577 (N_4577,N_4024,N_4389);
or U4578 (N_4578,N_4137,N_4236);
and U4579 (N_4579,N_4453,N_4038);
nor U4580 (N_4580,N_4314,N_4484);
or U4581 (N_4581,N_4441,N_4221);
xnor U4582 (N_4582,N_4364,N_4268);
or U4583 (N_4583,N_4106,N_4087);
nor U4584 (N_4584,N_4403,N_4410);
nand U4585 (N_4585,N_4498,N_4481);
nand U4586 (N_4586,N_4136,N_4252);
or U4587 (N_4587,N_4379,N_4020);
xor U4588 (N_4588,N_4028,N_4220);
nand U4589 (N_4589,N_4014,N_4037);
nand U4590 (N_4590,N_4158,N_4011);
nor U4591 (N_4591,N_4157,N_4211);
nor U4592 (N_4592,N_4057,N_4287);
nor U4593 (N_4593,N_4192,N_4374);
or U4594 (N_4594,N_4378,N_4070);
xor U4595 (N_4595,N_4116,N_4104);
and U4596 (N_4596,N_4293,N_4066);
xnor U4597 (N_4597,N_4267,N_4448);
nand U4598 (N_4598,N_4359,N_4153);
xor U4599 (N_4599,N_4162,N_4111);
nor U4600 (N_4600,N_4097,N_4394);
nand U4601 (N_4601,N_4063,N_4342);
xnor U4602 (N_4602,N_4000,N_4407);
or U4603 (N_4603,N_4036,N_4463);
and U4604 (N_4604,N_4142,N_4491);
or U4605 (N_4605,N_4060,N_4245);
or U4606 (N_4606,N_4457,N_4308);
nor U4607 (N_4607,N_4344,N_4209);
and U4608 (N_4608,N_4230,N_4319);
nand U4609 (N_4609,N_4313,N_4311);
nand U4610 (N_4610,N_4145,N_4026);
xor U4611 (N_4611,N_4223,N_4351);
or U4612 (N_4612,N_4101,N_4380);
or U4613 (N_4613,N_4402,N_4099);
nor U4614 (N_4614,N_4121,N_4439);
and U4615 (N_4615,N_4373,N_4033);
nor U4616 (N_4616,N_4178,N_4316);
xor U4617 (N_4617,N_4390,N_4471);
xor U4618 (N_4618,N_4324,N_4454);
nand U4619 (N_4619,N_4320,N_4088);
nor U4620 (N_4620,N_4118,N_4412);
nor U4621 (N_4621,N_4131,N_4369);
xnor U4622 (N_4622,N_4082,N_4233);
nor U4623 (N_4623,N_4377,N_4191);
xor U4624 (N_4624,N_4027,N_4152);
or U4625 (N_4625,N_4445,N_4166);
xor U4626 (N_4626,N_4022,N_4260);
and U4627 (N_4627,N_4352,N_4207);
and U4628 (N_4628,N_4100,N_4044);
xnor U4629 (N_4629,N_4213,N_4132);
or U4630 (N_4630,N_4214,N_4334);
xnor U4631 (N_4631,N_4103,N_4321);
or U4632 (N_4632,N_4054,N_4076);
xnor U4633 (N_4633,N_4458,N_4225);
and U4634 (N_4634,N_4248,N_4107);
and U4635 (N_4635,N_4235,N_4001);
or U4636 (N_4636,N_4096,N_4434);
and U4637 (N_4637,N_4426,N_4035);
and U4638 (N_4638,N_4485,N_4185);
or U4639 (N_4639,N_4449,N_4084);
nor U4640 (N_4640,N_4126,N_4470);
or U4641 (N_4641,N_4460,N_4194);
nand U4642 (N_4642,N_4234,N_4041);
and U4643 (N_4643,N_4294,N_4466);
or U4644 (N_4644,N_4186,N_4386);
and U4645 (N_4645,N_4354,N_4081);
nand U4646 (N_4646,N_4117,N_4335);
nor U4647 (N_4647,N_4490,N_4325);
or U4648 (N_4648,N_4177,N_4007);
or U4649 (N_4649,N_4456,N_4264);
nor U4650 (N_4650,N_4127,N_4222);
xor U4651 (N_4651,N_4034,N_4008);
nor U4652 (N_4652,N_4284,N_4347);
nor U4653 (N_4653,N_4110,N_4447);
or U4654 (N_4654,N_4013,N_4312);
and U4655 (N_4655,N_4289,N_4489);
or U4656 (N_4656,N_4042,N_4019);
or U4657 (N_4657,N_4446,N_4242);
xnor U4658 (N_4658,N_4219,N_4229);
xor U4659 (N_4659,N_4071,N_4303);
nand U4660 (N_4660,N_4261,N_4208);
nand U4661 (N_4661,N_4408,N_4190);
nor U4662 (N_4662,N_4056,N_4069);
nor U4663 (N_4663,N_4180,N_4168);
xor U4664 (N_4664,N_4343,N_4046);
and U4665 (N_4665,N_4003,N_4452);
and U4666 (N_4666,N_4331,N_4112);
and U4667 (N_4667,N_4296,N_4278);
and U4668 (N_4668,N_4141,N_4370);
or U4669 (N_4669,N_4048,N_4292);
nor U4670 (N_4670,N_4360,N_4475);
nand U4671 (N_4671,N_4328,N_4336);
or U4672 (N_4672,N_4193,N_4232);
nand U4673 (N_4673,N_4383,N_4164);
or U4674 (N_4674,N_4362,N_4258);
nor U4675 (N_4675,N_4217,N_4413);
xor U4676 (N_4676,N_4002,N_4251);
nand U4677 (N_4677,N_4226,N_4247);
nor U4678 (N_4678,N_4423,N_4160);
or U4679 (N_4679,N_4329,N_4273);
nor U4680 (N_4680,N_4130,N_4050);
nand U4681 (N_4681,N_4406,N_4332);
and U4682 (N_4682,N_4253,N_4358);
nand U4683 (N_4683,N_4006,N_4140);
and U4684 (N_4684,N_4254,N_4170);
xor U4685 (N_4685,N_4497,N_4114);
nand U4686 (N_4686,N_4265,N_4205);
or U4687 (N_4687,N_4414,N_4094);
xor U4688 (N_4688,N_4231,N_4052);
or U4689 (N_4689,N_4030,N_4451);
or U4690 (N_4690,N_4404,N_4065);
xnor U4691 (N_4691,N_4326,N_4409);
nor U4692 (N_4692,N_4120,N_4061);
or U4693 (N_4693,N_4371,N_4108);
and U4694 (N_4694,N_4418,N_4455);
and U4695 (N_4695,N_4134,N_4189);
nor U4696 (N_4696,N_4089,N_4124);
and U4697 (N_4697,N_4353,N_4227);
nand U4698 (N_4698,N_4198,N_4474);
nor U4699 (N_4699,N_4195,N_4237);
or U4700 (N_4700,N_4210,N_4350);
nand U4701 (N_4701,N_4440,N_4427);
xnor U4702 (N_4702,N_4286,N_4399);
nor U4703 (N_4703,N_4073,N_4206);
and U4704 (N_4704,N_4300,N_4385);
nand U4705 (N_4705,N_4388,N_4015);
or U4706 (N_4706,N_4149,N_4171);
xnor U4707 (N_4707,N_4479,N_4163);
xor U4708 (N_4708,N_4083,N_4429);
nand U4709 (N_4709,N_4480,N_4090);
nor U4710 (N_4710,N_4174,N_4391);
or U4711 (N_4711,N_4129,N_4092);
nor U4712 (N_4712,N_4499,N_4438);
xor U4713 (N_4713,N_4147,N_4148);
and U4714 (N_4714,N_4346,N_4372);
and U4715 (N_4715,N_4468,N_4138);
nand U4716 (N_4716,N_4306,N_4488);
and U4717 (N_4717,N_4368,N_4086);
nor U4718 (N_4718,N_4302,N_4240);
and U4719 (N_4719,N_4181,N_4031);
nand U4720 (N_4720,N_4349,N_4366);
and U4721 (N_4721,N_4259,N_4212);
nand U4722 (N_4722,N_4262,N_4175);
nor U4723 (N_4723,N_4411,N_4062);
or U4724 (N_4724,N_4009,N_4425);
nor U4725 (N_4725,N_4159,N_4395);
nor U4726 (N_4726,N_4102,N_4384);
and U4727 (N_4727,N_4310,N_4276);
nor U4728 (N_4728,N_4417,N_4467);
nor U4729 (N_4729,N_4282,N_4393);
nand U4730 (N_4730,N_4202,N_4381);
or U4731 (N_4731,N_4443,N_4155);
or U4732 (N_4732,N_4397,N_4375);
or U4733 (N_4733,N_4459,N_4281);
nand U4734 (N_4734,N_4239,N_4283);
nand U4735 (N_4735,N_4040,N_4169);
nor U4736 (N_4736,N_4244,N_4277);
or U4737 (N_4737,N_4361,N_4228);
nor U4738 (N_4738,N_4317,N_4154);
and U4739 (N_4739,N_4188,N_4144);
xor U4740 (N_4740,N_4133,N_4139);
nand U4741 (N_4741,N_4123,N_4279);
nor U4742 (N_4742,N_4249,N_4257);
nor U4743 (N_4743,N_4428,N_4150);
nand U4744 (N_4744,N_4318,N_4341);
nor U4745 (N_4745,N_4143,N_4392);
nor U4746 (N_4746,N_4337,N_4473);
nor U4747 (N_4747,N_4077,N_4270);
xor U4748 (N_4748,N_4327,N_4345);
or U4749 (N_4749,N_4021,N_4095);
nor U4750 (N_4750,N_4250,N_4078);
or U4751 (N_4751,N_4245,N_4370);
xor U4752 (N_4752,N_4188,N_4090);
nor U4753 (N_4753,N_4316,N_4206);
xnor U4754 (N_4754,N_4081,N_4412);
nor U4755 (N_4755,N_4346,N_4134);
nand U4756 (N_4756,N_4132,N_4153);
or U4757 (N_4757,N_4498,N_4238);
or U4758 (N_4758,N_4388,N_4075);
nor U4759 (N_4759,N_4400,N_4419);
xor U4760 (N_4760,N_4294,N_4143);
and U4761 (N_4761,N_4408,N_4238);
or U4762 (N_4762,N_4187,N_4157);
and U4763 (N_4763,N_4279,N_4278);
and U4764 (N_4764,N_4233,N_4307);
nor U4765 (N_4765,N_4383,N_4480);
nand U4766 (N_4766,N_4173,N_4316);
nor U4767 (N_4767,N_4068,N_4403);
nand U4768 (N_4768,N_4096,N_4011);
nand U4769 (N_4769,N_4116,N_4457);
or U4770 (N_4770,N_4412,N_4259);
or U4771 (N_4771,N_4073,N_4221);
or U4772 (N_4772,N_4143,N_4190);
and U4773 (N_4773,N_4203,N_4053);
nor U4774 (N_4774,N_4206,N_4280);
or U4775 (N_4775,N_4039,N_4439);
and U4776 (N_4776,N_4226,N_4498);
nor U4777 (N_4777,N_4462,N_4270);
nor U4778 (N_4778,N_4059,N_4156);
nand U4779 (N_4779,N_4408,N_4323);
xnor U4780 (N_4780,N_4138,N_4318);
and U4781 (N_4781,N_4447,N_4390);
nor U4782 (N_4782,N_4114,N_4129);
and U4783 (N_4783,N_4273,N_4004);
nand U4784 (N_4784,N_4182,N_4218);
and U4785 (N_4785,N_4285,N_4406);
and U4786 (N_4786,N_4084,N_4144);
nor U4787 (N_4787,N_4053,N_4080);
nand U4788 (N_4788,N_4129,N_4415);
or U4789 (N_4789,N_4380,N_4008);
and U4790 (N_4790,N_4115,N_4319);
or U4791 (N_4791,N_4199,N_4374);
or U4792 (N_4792,N_4417,N_4058);
nor U4793 (N_4793,N_4114,N_4301);
xnor U4794 (N_4794,N_4258,N_4447);
or U4795 (N_4795,N_4159,N_4110);
and U4796 (N_4796,N_4042,N_4424);
or U4797 (N_4797,N_4074,N_4014);
nand U4798 (N_4798,N_4478,N_4005);
and U4799 (N_4799,N_4163,N_4331);
or U4800 (N_4800,N_4395,N_4482);
or U4801 (N_4801,N_4226,N_4156);
and U4802 (N_4802,N_4044,N_4180);
and U4803 (N_4803,N_4399,N_4113);
nor U4804 (N_4804,N_4024,N_4466);
nor U4805 (N_4805,N_4055,N_4352);
nand U4806 (N_4806,N_4009,N_4176);
xor U4807 (N_4807,N_4090,N_4396);
and U4808 (N_4808,N_4458,N_4466);
xnor U4809 (N_4809,N_4060,N_4209);
or U4810 (N_4810,N_4281,N_4422);
nor U4811 (N_4811,N_4438,N_4433);
and U4812 (N_4812,N_4110,N_4321);
xnor U4813 (N_4813,N_4310,N_4375);
nor U4814 (N_4814,N_4437,N_4464);
and U4815 (N_4815,N_4302,N_4121);
nand U4816 (N_4816,N_4419,N_4265);
and U4817 (N_4817,N_4422,N_4378);
nor U4818 (N_4818,N_4306,N_4360);
nand U4819 (N_4819,N_4124,N_4366);
or U4820 (N_4820,N_4197,N_4233);
nor U4821 (N_4821,N_4095,N_4332);
nor U4822 (N_4822,N_4073,N_4395);
xnor U4823 (N_4823,N_4308,N_4200);
xnor U4824 (N_4824,N_4170,N_4272);
xnor U4825 (N_4825,N_4384,N_4131);
or U4826 (N_4826,N_4215,N_4435);
and U4827 (N_4827,N_4184,N_4145);
and U4828 (N_4828,N_4423,N_4197);
or U4829 (N_4829,N_4067,N_4386);
nor U4830 (N_4830,N_4301,N_4165);
nand U4831 (N_4831,N_4414,N_4107);
and U4832 (N_4832,N_4350,N_4316);
or U4833 (N_4833,N_4228,N_4173);
and U4834 (N_4834,N_4250,N_4205);
xor U4835 (N_4835,N_4006,N_4310);
nand U4836 (N_4836,N_4449,N_4440);
or U4837 (N_4837,N_4103,N_4227);
nor U4838 (N_4838,N_4057,N_4096);
and U4839 (N_4839,N_4243,N_4131);
or U4840 (N_4840,N_4147,N_4107);
nand U4841 (N_4841,N_4119,N_4044);
and U4842 (N_4842,N_4441,N_4481);
or U4843 (N_4843,N_4227,N_4489);
and U4844 (N_4844,N_4200,N_4197);
nand U4845 (N_4845,N_4328,N_4485);
xor U4846 (N_4846,N_4066,N_4472);
nand U4847 (N_4847,N_4173,N_4297);
nor U4848 (N_4848,N_4228,N_4212);
or U4849 (N_4849,N_4366,N_4099);
nor U4850 (N_4850,N_4307,N_4075);
and U4851 (N_4851,N_4266,N_4129);
or U4852 (N_4852,N_4189,N_4037);
nor U4853 (N_4853,N_4427,N_4407);
or U4854 (N_4854,N_4499,N_4348);
and U4855 (N_4855,N_4051,N_4152);
or U4856 (N_4856,N_4174,N_4092);
nor U4857 (N_4857,N_4450,N_4379);
nor U4858 (N_4858,N_4120,N_4230);
or U4859 (N_4859,N_4055,N_4416);
xor U4860 (N_4860,N_4071,N_4411);
and U4861 (N_4861,N_4299,N_4189);
or U4862 (N_4862,N_4233,N_4128);
xor U4863 (N_4863,N_4036,N_4103);
nor U4864 (N_4864,N_4387,N_4367);
nand U4865 (N_4865,N_4383,N_4133);
and U4866 (N_4866,N_4402,N_4130);
nor U4867 (N_4867,N_4053,N_4160);
or U4868 (N_4868,N_4030,N_4299);
and U4869 (N_4869,N_4193,N_4050);
nand U4870 (N_4870,N_4367,N_4463);
and U4871 (N_4871,N_4043,N_4048);
xnor U4872 (N_4872,N_4427,N_4253);
xor U4873 (N_4873,N_4004,N_4431);
nor U4874 (N_4874,N_4164,N_4485);
nor U4875 (N_4875,N_4206,N_4020);
or U4876 (N_4876,N_4180,N_4321);
nor U4877 (N_4877,N_4311,N_4419);
nor U4878 (N_4878,N_4217,N_4405);
and U4879 (N_4879,N_4303,N_4001);
nand U4880 (N_4880,N_4339,N_4105);
nor U4881 (N_4881,N_4327,N_4376);
or U4882 (N_4882,N_4169,N_4267);
or U4883 (N_4883,N_4389,N_4379);
xnor U4884 (N_4884,N_4404,N_4036);
nand U4885 (N_4885,N_4303,N_4090);
and U4886 (N_4886,N_4310,N_4110);
nand U4887 (N_4887,N_4030,N_4057);
and U4888 (N_4888,N_4484,N_4313);
xor U4889 (N_4889,N_4310,N_4248);
xor U4890 (N_4890,N_4412,N_4398);
nand U4891 (N_4891,N_4364,N_4237);
and U4892 (N_4892,N_4361,N_4109);
nand U4893 (N_4893,N_4037,N_4179);
or U4894 (N_4894,N_4403,N_4003);
nor U4895 (N_4895,N_4107,N_4153);
nand U4896 (N_4896,N_4030,N_4463);
nand U4897 (N_4897,N_4041,N_4252);
nor U4898 (N_4898,N_4280,N_4444);
and U4899 (N_4899,N_4089,N_4264);
nor U4900 (N_4900,N_4131,N_4398);
xor U4901 (N_4901,N_4193,N_4282);
nand U4902 (N_4902,N_4341,N_4085);
nor U4903 (N_4903,N_4388,N_4361);
and U4904 (N_4904,N_4461,N_4154);
or U4905 (N_4905,N_4420,N_4255);
nor U4906 (N_4906,N_4057,N_4023);
or U4907 (N_4907,N_4289,N_4054);
xnor U4908 (N_4908,N_4127,N_4235);
nor U4909 (N_4909,N_4495,N_4244);
nor U4910 (N_4910,N_4227,N_4273);
nor U4911 (N_4911,N_4181,N_4422);
nor U4912 (N_4912,N_4108,N_4064);
nor U4913 (N_4913,N_4197,N_4187);
nor U4914 (N_4914,N_4441,N_4224);
nand U4915 (N_4915,N_4483,N_4217);
nor U4916 (N_4916,N_4208,N_4153);
and U4917 (N_4917,N_4327,N_4301);
nand U4918 (N_4918,N_4211,N_4332);
and U4919 (N_4919,N_4033,N_4275);
nand U4920 (N_4920,N_4429,N_4439);
or U4921 (N_4921,N_4012,N_4457);
xnor U4922 (N_4922,N_4095,N_4074);
or U4923 (N_4923,N_4238,N_4318);
nor U4924 (N_4924,N_4137,N_4132);
nand U4925 (N_4925,N_4155,N_4118);
or U4926 (N_4926,N_4499,N_4274);
xnor U4927 (N_4927,N_4000,N_4434);
nand U4928 (N_4928,N_4078,N_4424);
nand U4929 (N_4929,N_4285,N_4355);
nor U4930 (N_4930,N_4249,N_4101);
or U4931 (N_4931,N_4045,N_4219);
and U4932 (N_4932,N_4421,N_4369);
xor U4933 (N_4933,N_4348,N_4484);
and U4934 (N_4934,N_4065,N_4483);
or U4935 (N_4935,N_4480,N_4194);
nand U4936 (N_4936,N_4381,N_4200);
nor U4937 (N_4937,N_4498,N_4248);
and U4938 (N_4938,N_4294,N_4235);
and U4939 (N_4939,N_4022,N_4170);
xor U4940 (N_4940,N_4415,N_4411);
xor U4941 (N_4941,N_4140,N_4284);
nand U4942 (N_4942,N_4024,N_4035);
or U4943 (N_4943,N_4465,N_4489);
and U4944 (N_4944,N_4414,N_4157);
or U4945 (N_4945,N_4435,N_4000);
and U4946 (N_4946,N_4237,N_4259);
nand U4947 (N_4947,N_4079,N_4481);
and U4948 (N_4948,N_4095,N_4499);
xor U4949 (N_4949,N_4115,N_4482);
or U4950 (N_4950,N_4323,N_4340);
nand U4951 (N_4951,N_4227,N_4366);
xnor U4952 (N_4952,N_4333,N_4113);
or U4953 (N_4953,N_4303,N_4021);
nand U4954 (N_4954,N_4453,N_4138);
nor U4955 (N_4955,N_4377,N_4431);
nand U4956 (N_4956,N_4352,N_4329);
xnor U4957 (N_4957,N_4307,N_4407);
and U4958 (N_4958,N_4498,N_4069);
nor U4959 (N_4959,N_4347,N_4077);
and U4960 (N_4960,N_4180,N_4458);
or U4961 (N_4961,N_4141,N_4388);
or U4962 (N_4962,N_4270,N_4301);
xnor U4963 (N_4963,N_4165,N_4348);
and U4964 (N_4964,N_4396,N_4027);
or U4965 (N_4965,N_4041,N_4458);
nand U4966 (N_4966,N_4419,N_4289);
and U4967 (N_4967,N_4417,N_4224);
xor U4968 (N_4968,N_4424,N_4103);
or U4969 (N_4969,N_4105,N_4244);
and U4970 (N_4970,N_4479,N_4010);
and U4971 (N_4971,N_4379,N_4210);
nand U4972 (N_4972,N_4478,N_4248);
nor U4973 (N_4973,N_4025,N_4128);
nand U4974 (N_4974,N_4411,N_4119);
or U4975 (N_4975,N_4233,N_4202);
nand U4976 (N_4976,N_4404,N_4224);
and U4977 (N_4977,N_4432,N_4455);
xnor U4978 (N_4978,N_4328,N_4277);
xor U4979 (N_4979,N_4392,N_4107);
nor U4980 (N_4980,N_4320,N_4432);
nand U4981 (N_4981,N_4308,N_4310);
and U4982 (N_4982,N_4124,N_4129);
and U4983 (N_4983,N_4287,N_4106);
and U4984 (N_4984,N_4361,N_4459);
xnor U4985 (N_4985,N_4072,N_4067);
nand U4986 (N_4986,N_4165,N_4333);
or U4987 (N_4987,N_4468,N_4404);
nor U4988 (N_4988,N_4262,N_4277);
or U4989 (N_4989,N_4352,N_4480);
xor U4990 (N_4990,N_4411,N_4420);
and U4991 (N_4991,N_4167,N_4123);
or U4992 (N_4992,N_4236,N_4459);
or U4993 (N_4993,N_4075,N_4081);
xnor U4994 (N_4994,N_4159,N_4282);
and U4995 (N_4995,N_4341,N_4094);
nand U4996 (N_4996,N_4316,N_4359);
nand U4997 (N_4997,N_4379,N_4368);
nand U4998 (N_4998,N_4058,N_4066);
nand U4999 (N_4999,N_4332,N_4138);
xnor UO_0 (O_0,N_4559,N_4865);
nand UO_1 (O_1,N_4843,N_4632);
and UO_2 (O_2,N_4514,N_4675);
xor UO_3 (O_3,N_4872,N_4605);
and UO_4 (O_4,N_4700,N_4595);
and UO_5 (O_5,N_4538,N_4877);
nand UO_6 (O_6,N_4989,N_4859);
and UO_7 (O_7,N_4880,N_4755);
nand UO_8 (O_8,N_4724,N_4784);
or UO_9 (O_9,N_4682,N_4516);
xor UO_10 (O_10,N_4555,N_4931);
or UO_11 (O_11,N_4846,N_4671);
and UO_12 (O_12,N_4864,N_4888);
xor UO_13 (O_13,N_4968,N_4806);
nand UO_14 (O_14,N_4519,N_4789);
nor UO_15 (O_15,N_4933,N_4578);
or UO_16 (O_16,N_4556,N_4820);
nor UO_17 (O_17,N_4657,N_4857);
xor UO_18 (O_18,N_4739,N_4730);
or UO_19 (O_19,N_4916,N_4737);
nand UO_20 (O_20,N_4701,N_4860);
and UO_21 (O_21,N_4500,N_4629);
and UO_22 (O_22,N_4696,N_4898);
nor UO_23 (O_23,N_4855,N_4845);
and UO_24 (O_24,N_4823,N_4583);
nor UO_25 (O_25,N_4972,N_4527);
nand UO_26 (O_26,N_4508,N_4803);
xor UO_27 (O_27,N_4738,N_4644);
nor UO_28 (O_28,N_4734,N_4952);
nor UO_29 (O_29,N_4854,N_4853);
xor UO_30 (O_30,N_4997,N_4785);
nand UO_31 (O_31,N_4658,N_4711);
or UO_32 (O_32,N_4897,N_4908);
xor UO_33 (O_33,N_4746,N_4679);
xor UO_34 (O_34,N_4725,N_4546);
or UO_35 (O_35,N_4768,N_4866);
nor UO_36 (O_36,N_4673,N_4764);
and UO_37 (O_37,N_4541,N_4608);
nand UO_38 (O_38,N_4603,N_4732);
and UO_39 (O_39,N_4572,N_4506);
nand UO_40 (O_40,N_4532,N_4715);
nand UO_41 (O_41,N_4907,N_4534);
and UO_42 (O_42,N_4645,N_4920);
xnor UO_43 (O_43,N_4960,N_4777);
or UO_44 (O_44,N_4970,N_4975);
nand UO_45 (O_45,N_4837,N_4979);
xnor UO_46 (O_46,N_4856,N_4616);
nand UO_47 (O_47,N_4669,N_4827);
nor UO_48 (O_48,N_4905,N_4552);
or UO_49 (O_49,N_4874,N_4901);
xor UO_50 (O_50,N_4790,N_4526);
xnor UO_51 (O_51,N_4625,N_4835);
nor UO_52 (O_52,N_4766,N_4903);
and UO_53 (O_53,N_4973,N_4999);
and UO_54 (O_54,N_4798,N_4723);
nor UO_55 (O_55,N_4650,N_4709);
xor UO_56 (O_56,N_4512,N_4831);
and UO_57 (O_57,N_4930,N_4811);
nor UO_58 (O_58,N_4704,N_4513);
and UO_59 (O_59,N_4545,N_4763);
xor UO_60 (O_60,N_4653,N_4956);
nand UO_61 (O_61,N_4713,N_4560);
nor UO_62 (O_62,N_4627,N_4943);
and UO_63 (O_63,N_4733,N_4630);
nor UO_64 (O_64,N_4941,N_4996);
or UO_65 (O_65,N_4664,N_4776);
xnor UO_66 (O_66,N_4949,N_4988);
xnor UO_67 (O_67,N_4567,N_4980);
nand UO_68 (O_68,N_4707,N_4544);
and UO_69 (O_69,N_4576,N_4992);
xnor UO_70 (O_70,N_4942,N_4579);
or UO_71 (O_71,N_4502,N_4727);
and UO_72 (O_72,N_4944,N_4794);
and UO_73 (O_73,N_4935,N_4847);
nor UO_74 (O_74,N_4585,N_4986);
and UO_75 (O_75,N_4726,N_4805);
or UO_76 (O_76,N_4531,N_4976);
and UO_77 (O_77,N_4521,N_4965);
or UO_78 (O_78,N_4833,N_4587);
or UO_79 (O_79,N_4719,N_4743);
nor UO_80 (O_80,N_4774,N_4554);
xor UO_81 (O_81,N_4917,N_4800);
nand UO_82 (O_82,N_4926,N_4598);
xor UO_83 (O_83,N_4614,N_4957);
xnor UO_84 (O_84,N_4543,N_4720);
nor UO_85 (O_85,N_4735,N_4773);
nor UO_86 (O_86,N_4558,N_4981);
nor UO_87 (O_87,N_4934,N_4836);
and UO_88 (O_88,N_4987,N_4652);
and UO_89 (O_89,N_4580,N_4649);
or UO_90 (O_90,N_4588,N_4796);
or UO_91 (O_91,N_4540,N_4550);
or UO_92 (O_92,N_4690,N_4520);
nand UO_93 (O_93,N_4816,N_4721);
xnor UO_94 (O_94,N_4814,N_4818);
and UO_95 (O_95,N_4772,N_4563);
nor UO_96 (O_96,N_4691,N_4678);
and UO_97 (O_97,N_4535,N_4640);
nand UO_98 (O_98,N_4883,N_4716);
xor UO_99 (O_99,N_4852,N_4950);
xnor UO_100 (O_100,N_4828,N_4600);
nor UO_101 (O_101,N_4524,N_4659);
xnor UO_102 (O_102,N_4830,N_4984);
and UO_103 (O_103,N_4548,N_4677);
or UO_104 (O_104,N_4802,N_4870);
xor UO_105 (O_105,N_4757,N_4947);
xor UO_106 (O_106,N_4937,N_4517);
or UO_107 (O_107,N_4891,N_4611);
nor UO_108 (O_108,N_4710,N_4684);
xnor UO_109 (O_109,N_4876,N_4528);
or UO_110 (O_110,N_4536,N_4939);
nor UO_111 (O_111,N_4887,N_4919);
or UO_112 (O_112,N_4667,N_4672);
and UO_113 (O_113,N_4788,N_4889);
nand UO_114 (O_114,N_4680,N_4760);
and UO_115 (O_115,N_4615,N_4728);
xor UO_116 (O_116,N_4551,N_4523);
and UO_117 (O_117,N_4892,N_4714);
nand UO_118 (O_118,N_4601,N_4886);
and UO_119 (O_119,N_4791,N_4770);
or UO_120 (O_120,N_4745,N_4634);
nand UO_121 (O_121,N_4529,N_4838);
nor UO_122 (O_122,N_4861,N_4792);
xor UO_123 (O_123,N_4951,N_4620);
nand UO_124 (O_124,N_4923,N_4825);
nor UO_125 (O_125,N_4695,N_4656);
nand UO_126 (O_126,N_4851,N_4963);
nand UO_127 (O_127,N_4841,N_4844);
and UO_128 (O_128,N_4964,N_4638);
or UO_129 (O_129,N_4940,N_4573);
xor UO_130 (O_130,N_4626,N_4668);
nor UO_131 (O_131,N_4651,N_4596);
xor UO_132 (O_132,N_4624,N_4922);
and UO_133 (O_133,N_4869,N_4592);
xnor UO_134 (O_134,N_4740,N_4910);
nand UO_135 (O_135,N_4688,N_4879);
or UO_136 (O_136,N_4775,N_4708);
and UO_137 (O_137,N_4797,N_4685);
or UO_138 (O_138,N_4561,N_4863);
or UO_139 (O_139,N_4594,N_4894);
or UO_140 (O_140,N_4779,N_4842);
nand UO_141 (O_141,N_4602,N_4660);
and UO_142 (O_142,N_4966,N_4769);
and UO_143 (O_143,N_4821,N_4610);
or UO_144 (O_144,N_4881,N_4501);
xnor UO_145 (O_145,N_4961,N_4812);
or UO_146 (O_146,N_4982,N_4599);
xnor UO_147 (O_147,N_4718,N_4912);
or UO_148 (O_148,N_4515,N_4815);
and UO_149 (O_149,N_4974,N_4782);
xor UO_150 (O_150,N_4754,N_4813);
and UO_151 (O_151,N_4566,N_4758);
xor UO_152 (O_152,N_4547,N_4744);
nor UO_153 (O_153,N_4822,N_4537);
and UO_154 (O_154,N_4850,N_4778);
nand UO_155 (O_155,N_4875,N_4697);
and UO_156 (O_156,N_4993,N_4533);
xnor UO_157 (O_157,N_4712,N_4868);
and UO_158 (O_158,N_4575,N_4646);
and UO_159 (O_159,N_4932,N_4804);
nand UO_160 (O_160,N_4748,N_4848);
xor UO_161 (O_161,N_4826,N_4689);
nand UO_162 (O_162,N_4693,N_4642);
or UO_163 (O_163,N_4643,N_4783);
nor UO_164 (O_164,N_4510,N_4590);
nor UO_165 (O_165,N_4749,N_4895);
nor UO_166 (O_166,N_4702,N_4906);
nor UO_167 (O_167,N_4562,N_4666);
xnor UO_168 (O_168,N_4604,N_4589);
xnor UO_169 (O_169,N_4808,N_4581);
nor UO_170 (O_170,N_4871,N_4570);
nand UO_171 (O_171,N_4717,N_4765);
xnor UO_172 (O_172,N_4948,N_4687);
nand UO_173 (O_173,N_4810,N_4676);
nand UO_174 (O_174,N_4584,N_4703);
or UO_175 (O_175,N_4809,N_4882);
and UO_176 (O_176,N_4839,N_4606);
xnor UO_177 (O_177,N_4801,N_4539);
and UO_178 (O_178,N_4662,N_4913);
and UO_179 (O_179,N_4832,N_4557);
nand UO_180 (O_180,N_4681,N_4530);
xnor UO_181 (O_181,N_4819,N_4824);
and UO_182 (O_182,N_4998,N_4504);
or UO_183 (O_183,N_4674,N_4953);
xor UO_184 (O_184,N_4741,N_4522);
nand UO_185 (O_185,N_4571,N_4636);
xor UO_186 (O_186,N_4663,N_4705);
and UO_187 (O_187,N_4885,N_4577);
and UO_188 (O_188,N_4756,N_4762);
nor UO_189 (O_189,N_4647,N_4582);
or UO_190 (O_190,N_4736,N_4503);
and UO_191 (O_191,N_4661,N_4817);
and UO_192 (O_192,N_4747,N_4958);
or UO_193 (O_193,N_4752,N_4729);
xor UO_194 (O_194,N_4631,N_4623);
and UO_195 (O_195,N_4549,N_4962);
nand UO_196 (O_196,N_4786,N_4896);
or UO_197 (O_197,N_4890,N_4670);
and UO_198 (O_198,N_4635,N_4936);
or UO_199 (O_199,N_4665,N_4722);
nand UO_200 (O_200,N_4591,N_4927);
or UO_201 (O_201,N_4928,N_4751);
nor UO_202 (O_202,N_4639,N_4706);
nand UO_203 (O_203,N_4621,N_4946);
or UO_204 (O_204,N_4918,N_4893);
and UO_205 (O_205,N_4929,N_4593);
nand UO_206 (O_206,N_4904,N_4613);
xnor UO_207 (O_207,N_4654,N_4862);
nand UO_208 (O_208,N_4771,N_4699);
or UO_209 (O_209,N_4900,N_4759);
or UO_210 (O_210,N_4967,N_4925);
and UO_211 (O_211,N_4607,N_4955);
xor UO_212 (O_212,N_4641,N_4971);
or UO_213 (O_213,N_4750,N_4622);
and UO_214 (O_214,N_4692,N_4954);
and UO_215 (O_215,N_4921,N_4731);
nor UO_216 (O_216,N_4924,N_4990);
or UO_217 (O_217,N_4618,N_4867);
nand UO_218 (O_218,N_4915,N_4795);
and UO_219 (O_219,N_4909,N_4799);
and UO_220 (O_220,N_4609,N_4633);
nor UO_221 (O_221,N_4655,N_4780);
nand UO_222 (O_222,N_4509,N_4781);
and UO_223 (O_223,N_4518,N_4507);
nand UO_224 (O_224,N_4995,N_4565);
xor UO_225 (O_225,N_4568,N_4542);
nand UO_226 (O_226,N_4899,N_4648);
and UO_227 (O_227,N_4753,N_4694);
nand UO_228 (O_228,N_4793,N_4834);
nand UO_229 (O_229,N_4902,N_4698);
and UO_230 (O_230,N_4969,N_4840);
or UO_231 (O_231,N_4945,N_4938);
or UO_232 (O_232,N_4637,N_4617);
or UO_233 (O_233,N_4564,N_4991);
xor UO_234 (O_234,N_4829,N_4569);
xnor UO_235 (O_235,N_4985,N_4525);
xor UO_236 (O_236,N_4511,N_4873);
xnor UO_237 (O_237,N_4761,N_4612);
or UO_238 (O_238,N_4878,N_4914);
xor UO_239 (O_239,N_4686,N_4683);
and UO_240 (O_240,N_4505,N_4767);
nand UO_241 (O_241,N_4807,N_4849);
nor UO_242 (O_242,N_4978,N_4959);
xor UO_243 (O_243,N_4884,N_4586);
and UO_244 (O_244,N_4994,N_4977);
nor UO_245 (O_245,N_4742,N_4911);
nor UO_246 (O_246,N_4574,N_4983);
and UO_247 (O_247,N_4597,N_4628);
nand UO_248 (O_248,N_4619,N_4858);
and UO_249 (O_249,N_4787,N_4553);
and UO_250 (O_250,N_4540,N_4829);
or UO_251 (O_251,N_4981,N_4538);
nand UO_252 (O_252,N_4846,N_4739);
nand UO_253 (O_253,N_4810,N_4952);
and UO_254 (O_254,N_4931,N_4893);
nor UO_255 (O_255,N_4535,N_4753);
nor UO_256 (O_256,N_4837,N_4903);
nor UO_257 (O_257,N_4820,N_4513);
nand UO_258 (O_258,N_4603,N_4797);
nand UO_259 (O_259,N_4701,N_4841);
nor UO_260 (O_260,N_4864,N_4521);
nor UO_261 (O_261,N_4680,N_4807);
or UO_262 (O_262,N_4821,N_4578);
nand UO_263 (O_263,N_4514,N_4563);
nor UO_264 (O_264,N_4625,N_4560);
or UO_265 (O_265,N_4981,N_4886);
or UO_266 (O_266,N_4549,N_4582);
nand UO_267 (O_267,N_4987,N_4762);
or UO_268 (O_268,N_4849,N_4594);
nand UO_269 (O_269,N_4577,N_4631);
xor UO_270 (O_270,N_4643,N_4635);
and UO_271 (O_271,N_4941,N_4669);
or UO_272 (O_272,N_4760,N_4603);
nand UO_273 (O_273,N_4638,N_4713);
nor UO_274 (O_274,N_4884,N_4860);
or UO_275 (O_275,N_4603,N_4619);
and UO_276 (O_276,N_4650,N_4575);
and UO_277 (O_277,N_4701,N_4783);
xor UO_278 (O_278,N_4726,N_4872);
or UO_279 (O_279,N_4943,N_4559);
nand UO_280 (O_280,N_4633,N_4516);
and UO_281 (O_281,N_4519,N_4788);
and UO_282 (O_282,N_4794,N_4963);
or UO_283 (O_283,N_4765,N_4916);
nand UO_284 (O_284,N_4571,N_4813);
nand UO_285 (O_285,N_4669,N_4567);
nor UO_286 (O_286,N_4682,N_4505);
nand UO_287 (O_287,N_4616,N_4700);
or UO_288 (O_288,N_4524,N_4980);
or UO_289 (O_289,N_4772,N_4738);
xor UO_290 (O_290,N_4532,N_4639);
nand UO_291 (O_291,N_4990,N_4972);
and UO_292 (O_292,N_4983,N_4975);
nor UO_293 (O_293,N_4973,N_4767);
nand UO_294 (O_294,N_4949,N_4946);
nor UO_295 (O_295,N_4514,N_4852);
and UO_296 (O_296,N_4616,N_4816);
and UO_297 (O_297,N_4593,N_4615);
xnor UO_298 (O_298,N_4876,N_4760);
xor UO_299 (O_299,N_4926,N_4858);
nor UO_300 (O_300,N_4998,N_4506);
and UO_301 (O_301,N_4809,N_4648);
xnor UO_302 (O_302,N_4730,N_4917);
nor UO_303 (O_303,N_4752,N_4749);
and UO_304 (O_304,N_4631,N_4745);
nor UO_305 (O_305,N_4659,N_4700);
or UO_306 (O_306,N_4515,N_4559);
nand UO_307 (O_307,N_4741,N_4988);
or UO_308 (O_308,N_4775,N_4600);
nor UO_309 (O_309,N_4510,N_4589);
or UO_310 (O_310,N_4776,N_4803);
nand UO_311 (O_311,N_4883,N_4943);
xnor UO_312 (O_312,N_4551,N_4770);
xor UO_313 (O_313,N_4599,N_4830);
nand UO_314 (O_314,N_4519,N_4813);
xor UO_315 (O_315,N_4614,N_4762);
and UO_316 (O_316,N_4915,N_4933);
and UO_317 (O_317,N_4808,N_4989);
or UO_318 (O_318,N_4654,N_4503);
and UO_319 (O_319,N_4784,N_4638);
xor UO_320 (O_320,N_4902,N_4963);
nor UO_321 (O_321,N_4634,N_4781);
nand UO_322 (O_322,N_4913,N_4734);
or UO_323 (O_323,N_4887,N_4616);
nor UO_324 (O_324,N_4812,N_4784);
nor UO_325 (O_325,N_4702,N_4823);
nand UO_326 (O_326,N_4538,N_4813);
and UO_327 (O_327,N_4808,N_4957);
xnor UO_328 (O_328,N_4714,N_4549);
nand UO_329 (O_329,N_4907,N_4787);
nand UO_330 (O_330,N_4939,N_4856);
and UO_331 (O_331,N_4865,N_4897);
xor UO_332 (O_332,N_4996,N_4849);
or UO_333 (O_333,N_4928,N_4668);
nor UO_334 (O_334,N_4665,N_4694);
nand UO_335 (O_335,N_4686,N_4570);
nor UO_336 (O_336,N_4905,N_4626);
nor UO_337 (O_337,N_4761,N_4864);
nand UO_338 (O_338,N_4988,N_4709);
xnor UO_339 (O_339,N_4742,N_4840);
nand UO_340 (O_340,N_4503,N_4861);
and UO_341 (O_341,N_4609,N_4706);
and UO_342 (O_342,N_4850,N_4932);
nand UO_343 (O_343,N_4653,N_4869);
and UO_344 (O_344,N_4639,N_4726);
nand UO_345 (O_345,N_4852,N_4812);
nand UO_346 (O_346,N_4687,N_4941);
and UO_347 (O_347,N_4947,N_4817);
nand UO_348 (O_348,N_4856,N_4608);
and UO_349 (O_349,N_4819,N_4877);
and UO_350 (O_350,N_4632,N_4978);
and UO_351 (O_351,N_4854,N_4649);
nor UO_352 (O_352,N_4939,N_4726);
and UO_353 (O_353,N_4659,N_4651);
nor UO_354 (O_354,N_4558,N_4744);
xnor UO_355 (O_355,N_4928,N_4893);
and UO_356 (O_356,N_4759,N_4906);
or UO_357 (O_357,N_4839,N_4970);
xor UO_358 (O_358,N_4597,N_4810);
xnor UO_359 (O_359,N_4865,N_4674);
xnor UO_360 (O_360,N_4670,N_4537);
or UO_361 (O_361,N_4751,N_4913);
nor UO_362 (O_362,N_4945,N_4883);
nor UO_363 (O_363,N_4773,N_4698);
xor UO_364 (O_364,N_4703,N_4608);
and UO_365 (O_365,N_4991,N_4774);
nand UO_366 (O_366,N_4725,N_4882);
nor UO_367 (O_367,N_4655,N_4514);
or UO_368 (O_368,N_4830,N_4677);
nand UO_369 (O_369,N_4817,N_4785);
xor UO_370 (O_370,N_4944,N_4719);
or UO_371 (O_371,N_4662,N_4783);
nor UO_372 (O_372,N_4949,N_4599);
nand UO_373 (O_373,N_4509,N_4743);
nand UO_374 (O_374,N_4573,N_4506);
xnor UO_375 (O_375,N_4731,N_4564);
or UO_376 (O_376,N_4834,N_4983);
nor UO_377 (O_377,N_4567,N_4720);
and UO_378 (O_378,N_4889,N_4726);
nor UO_379 (O_379,N_4559,N_4899);
nor UO_380 (O_380,N_4745,N_4917);
and UO_381 (O_381,N_4777,N_4574);
or UO_382 (O_382,N_4851,N_4794);
and UO_383 (O_383,N_4777,N_4660);
nor UO_384 (O_384,N_4730,N_4942);
and UO_385 (O_385,N_4926,N_4979);
xor UO_386 (O_386,N_4767,N_4855);
xor UO_387 (O_387,N_4550,N_4932);
or UO_388 (O_388,N_4610,N_4931);
nand UO_389 (O_389,N_4672,N_4807);
and UO_390 (O_390,N_4605,N_4770);
or UO_391 (O_391,N_4773,N_4697);
or UO_392 (O_392,N_4827,N_4867);
xnor UO_393 (O_393,N_4531,N_4864);
nand UO_394 (O_394,N_4918,N_4894);
xor UO_395 (O_395,N_4968,N_4960);
nor UO_396 (O_396,N_4994,N_4944);
or UO_397 (O_397,N_4516,N_4792);
and UO_398 (O_398,N_4717,N_4924);
or UO_399 (O_399,N_4775,N_4529);
xor UO_400 (O_400,N_4549,N_4777);
xnor UO_401 (O_401,N_4551,N_4790);
nor UO_402 (O_402,N_4879,N_4880);
or UO_403 (O_403,N_4877,N_4765);
nor UO_404 (O_404,N_4917,N_4746);
nand UO_405 (O_405,N_4782,N_4980);
and UO_406 (O_406,N_4573,N_4552);
nor UO_407 (O_407,N_4951,N_4836);
or UO_408 (O_408,N_4752,N_4694);
and UO_409 (O_409,N_4569,N_4691);
and UO_410 (O_410,N_4938,N_4696);
or UO_411 (O_411,N_4778,N_4688);
or UO_412 (O_412,N_4605,N_4602);
or UO_413 (O_413,N_4771,N_4524);
xnor UO_414 (O_414,N_4994,N_4879);
xnor UO_415 (O_415,N_4768,N_4575);
nor UO_416 (O_416,N_4546,N_4637);
or UO_417 (O_417,N_4804,N_4622);
or UO_418 (O_418,N_4837,N_4723);
or UO_419 (O_419,N_4998,N_4627);
xor UO_420 (O_420,N_4747,N_4799);
xor UO_421 (O_421,N_4569,N_4692);
nand UO_422 (O_422,N_4792,N_4837);
nor UO_423 (O_423,N_4573,N_4831);
and UO_424 (O_424,N_4701,N_4541);
xnor UO_425 (O_425,N_4942,N_4953);
nand UO_426 (O_426,N_4577,N_4538);
or UO_427 (O_427,N_4754,N_4625);
nor UO_428 (O_428,N_4718,N_4776);
nand UO_429 (O_429,N_4918,N_4904);
or UO_430 (O_430,N_4768,N_4697);
nor UO_431 (O_431,N_4899,N_4900);
nand UO_432 (O_432,N_4555,N_4878);
xnor UO_433 (O_433,N_4806,N_4969);
or UO_434 (O_434,N_4910,N_4732);
xnor UO_435 (O_435,N_4559,N_4620);
and UO_436 (O_436,N_4553,N_4654);
nand UO_437 (O_437,N_4868,N_4677);
and UO_438 (O_438,N_4903,N_4663);
or UO_439 (O_439,N_4786,N_4680);
or UO_440 (O_440,N_4691,N_4959);
or UO_441 (O_441,N_4957,N_4806);
nor UO_442 (O_442,N_4969,N_4727);
nand UO_443 (O_443,N_4778,N_4971);
nor UO_444 (O_444,N_4733,N_4757);
nand UO_445 (O_445,N_4914,N_4853);
nand UO_446 (O_446,N_4943,N_4758);
nand UO_447 (O_447,N_4638,N_4772);
xor UO_448 (O_448,N_4986,N_4624);
nor UO_449 (O_449,N_4942,N_4875);
or UO_450 (O_450,N_4664,N_4968);
and UO_451 (O_451,N_4629,N_4509);
and UO_452 (O_452,N_4875,N_4543);
xnor UO_453 (O_453,N_4995,N_4562);
or UO_454 (O_454,N_4926,N_4830);
nand UO_455 (O_455,N_4895,N_4933);
and UO_456 (O_456,N_4644,N_4523);
or UO_457 (O_457,N_4555,N_4591);
nor UO_458 (O_458,N_4788,N_4962);
and UO_459 (O_459,N_4559,N_4609);
or UO_460 (O_460,N_4789,N_4509);
or UO_461 (O_461,N_4610,N_4995);
xor UO_462 (O_462,N_4823,N_4801);
and UO_463 (O_463,N_4843,N_4743);
xnor UO_464 (O_464,N_4532,N_4947);
nand UO_465 (O_465,N_4731,N_4963);
or UO_466 (O_466,N_4843,N_4996);
or UO_467 (O_467,N_4933,N_4616);
xnor UO_468 (O_468,N_4858,N_4862);
or UO_469 (O_469,N_4883,N_4863);
nand UO_470 (O_470,N_4813,N_4688);
xnor UO_471 (O_471,N_4650,N_4669);
xor UO_472 (O_472,N_4699,N_4984);
or UO_473 (O_473,N_4669,N_4559);
xnor UO_474 (O_474,N_4753,N_4647);
nand UO_475 (O_475,N_4943,N_4672);
and UO_476 (O_476,N_4978,N_4828);
nor UO_477 (O_477,N_4614,N_4500);
or UO_478 (O_478,N_4510,N_4653);
xnor UO_479 (O_479,N_4776,N_4628);
and UO_480 (O_480,N_4887,N_4622);
and UO_481 (O_481,N_4666,N_4662);
and UO_482 (O_482,N_4972,N_4883);
nand UO_483 (O_483,N_4546,N_4657);
xnor UO_484 (O_484,N_4902,N_4547);
nor UO_485 (O_485,N_4841,N_4934);
and UO_486 (O_486,N_4630,N_4783);
or UO_487 (O_487,N_4672,N_4792);
nand UO_488 (O_488,N_4678,N_4625);
xnor UO_489 (O_489,N_4900,N_4778);
nor UO_490 (O_490,N_4952,N_4688);
nor UO_491 (O_491,N_4614,N_4991);
nor UO_492 (O_492,N_4908,N_4793);
or UO_493 (O_493,N_4788,N_4852);
and UO_494 (O_494,N_4626,N_4694);
nand UO_495 (O_495,N_4553,N_4818);
xnor UO_496 (O_496,N_4860,N_4529);
and UO_497 (O_497,N_4637,N_4776);
nor UO_498 (O_498,N_4663,N_4682);
nor UO_499 (O_499,N_4539,N_4947);
and UO_500 (O_500,N_4733,N_4657);
and UO_501 (O_501,N_4938,N_4948);
nand UO_502 (O_502,N_4937,N_4616);
xor UO_503 (O_503,N_4864,N_4778);
and UO_504 (O_504,N_4960,N_4900);
xnor UO_505 (O_505,N_4552,N_4565);
nor UO_506 (O_506,N_4759,N_4894);
xor UO_507 (O_507,N_4984,N_4871);
nor UO_508 (O_508,N_4826,N_4724);
nand UO_509 (O_509,N_4882,N_4533);
nand UO_510 (O_510,N_4784,N_4772);
xor UO_511 (O_511,N_4856,N_4680);
and UO_512 (O_512,N_4660,N_4655);
nand UO_513 (O_513,N_4631,N_4744);
or UO_514 (O_514,N_4641,N_4731);
and UO_515 (O_515,N_4904,N_4562);
nand UO_516 (O_516,N_4677,N_4862);
xnor UO_517 (O_517,N_4875,N_4614);
or UO_518 (O_518,N_4624,N_4794);
or UO_519 (O_519,N_4547,N_4876);
nand UO_520 (O_520,N_4831,N_4841);
nand UO_521 (O_521,N_4521,N_4990);
or UO_522 (O_522,N_4721,N_4651);
nor UO_523 (O_523,N_4513,N_4666);
and UO_524 (O_524,N_4658,N_4548);
nor UO_525 (O_525,N_4533,N_4601);
nor UO_526 (O_526,N_4897,N_4989);
and UO_527 (O_527,N_4604,N_4769);
or UO_528 (O_528,N_4628,N_4742);
nand UO_529 (O_529,N_4592,N_4998);
nor UO_530 (O_530,N_4996,N_4719);
or UO_531 (O_531,N_4771,N_4928);
or UO_532 (O_532,N_4924,N_4541);
and UO_533 (O_533,N_4664,N_4517);
nor UO_534 (O_534,N_4705,N_4685);
or UO_535 (O_535,N_4837,N_4772);
and UO_536 (O_536,N_4771,N_4782);
nor UO_537 (O_537,N_4865,N_4677);
nand UO_538 (O_538,N_4760,N_4548);
or UO_539 (O_539,N_4878,N_4848);
nand UO_540 (O_540,N_4546,N_4565);
nand UO_541 (O_541,N_4550,N_4532);
xnor UO_542 (O_542,N_4581,N_4550);
xor UO_543 (O_543,N_4503,N_4966);
or UO_544 (O_544,N_4566,N_4501);
nor UO_545 (O_545,N_4821,N_4874);
nand UO_546 (O_546,N_4529,N_4722);
and UO_547 (O_547,N_4626,N_4660);
xor UO_548 (O_548,N_4573,N_4708);
nand UO_549 (O_549,N_4949,N_4764);
or UO_550 (O_550,N_4976,N_4664);
xnor UO_551 (O_551,N_4507,N_4617);
xor UO_552 (O_552,N_4796,N_4890);
or UO_553 (O_553,N_4524,N_4753);
nor UO_554 (O_554,N_4924,N_4881);
and UO_555 (O_555,N_4616,N_4605);
nor UO_556 (O_556,N_4977,N_4965);
xor UO_557 (O_557,N_4617,N_4746);
nand UO_558 (O_558,N_4620,N_4632);
nor UO_559 (O_559,N_4904,N_4882);
nor UO_560 (O_560,N_4983,N_4749);
or UO_561 (O_561,N_4756,N_4691);
or UO_562 (O_562,N_4766,N_4512);
nor UO_563 (O_563,N_4880,N_4587);
xnor UO_564 (O_564,N_4752,N_4662);
xor UO_565 (O_565,N_4741,N_4905);
nand UO_566 (O_566,N_4671,N_4798);
xor UO_567 (O_567,N_4600,N_4577);
or UO_568 (O_568,N_4611,N_4796);
nor UO_569 (O_569,N_4847,N_4828);
and UO_570 (O_570,N_4800,N_4971);
nor UO_571 (O_571,N_4982,N_4919);
or UO_572 (O_572,N_4901,N_4790);
xnor UO_573 (O_573,N_4519,N_4664);
xnor UO_574 (O_574,N_4941,N_4724);
nor UO_575 (O_575,N_4636,N_4868);
or UO_576 (O_576,N_4560,N_4836);
and UO_577 (O_577,N_4722,N_4565);
and UO_578 (O_578,N_4900,N_4631);
or UO_579 (O_579,N_4962,N_4728);
nand UO_580 (O_580,N_4761,N_4875);
nand UO_581 (O_581,N_4825,N_4680);
xnor UO_582 (O_582,N_4905,N_4972);
nor UO_583 (O_583,N_4897,N_4545);
nand UO_584 (O_584,N_4746,N_4812);
nand UO_585 (O_585,N_4637,N_4970);
nor UO_586 (O_586,N_4766,N_4595);
and UO_587 (O_587,N_4646,N_4905);
nand UO_588 (O_588,N_4580,N_4667);
nor UO_589 (O_589,N_4906,N_4620);
and UO_590 (O_590,N_4921,N_4504);
and UO_591 (O_591,N_4753,N_4754);
nand UO_592 (O_592,N_4508,N_4902);
or UO_593 (O_593,N_4746,N_4738);
nand UO_594 (O_594,N_4943,N_4660);
and UO_595 (O_595,N_4983,N_4752);
nand UO_596 (O_596,N_4931,N_4900);
or UO_597 (O_597,N_4668,N_4910);
nand UO_598 (O_598,N_4816,N_4799);
nor UO_599 (O_599,N_4568,N_4755);
nor UO_600 (O_600,N_4873,N_4844);
and UO_601 (O_601,N_4839,N_4507);
nor UO_602 (O_602,N_4808,N_4682);
and UO_603 (O_603,N_4991,N_4516);
or UO_604 (O_604,N_4614,N_4605);
nand UO_605 (O_605,N_4594,N_4978);
nor UO_606 (O_606,N_4545,N_4766);
nand UO_607 (O_607,N_4641,N_4847);
xnor UO_608 (O_608,N_4523,N_4716);
or UO_609 (O_609,N_4708,N_4711);
and UO_610 (O_610,N_4780,N_4916);
and UO_611 (O_611,N_4836,N_4807);
nor UO_612 (O_612,N_4700,N_4513);
nand UO_613 (O_613,N_4942,N_4917);
xor UO_614 (O_614,N_4703,N_4834);
xor UO_615 (O_615,N_4697,N_4954);
nand UO_616 (O_616,N_4921,N_4646);
nor UO_617 (O_617,N_4916,N_4588);
nand UO_618 (O_618,N_4813,N_4765);
xnor UO_619 (O_619,N_4902,N_4844);
nor UO_620 (O_620,N_4924,N_4527);
xor UO_621 (O_621,N_4736,N_4921);
nor UO_622 (O_622,N_4859,N_4882);
nor UO_623 (O_623,N_4908,N_4824);
and UO_624 (O_624,N_4571,N_4819);
nand UO_625 (O_625,N_4662,N_4606);
and UO_626 (O_626,N_4673,N_4555);
and UO_627 (O_627,N_4724,N_4675);
nand UO_628 (O_628,N_4906,N_4856);
nand UO_629 (O_629,N_4972,N_4957);
nor UO_630 (O_630,N_4745,N_4787);
and UO_631 (O_631,N_4741,N_4922);
and UO_632 (O_632,N_4555,N_4784);
xor UO_633 (O_633,N_4918,N_4722);
nand UO_634 (O_634,N_4710,N_4826);
or UO_635 (O_635,N_4894,N_4821);
and UO_636 (O_636,N_4580,N_4615);
nor UO_637 (O_637,N_4653,N_4665);
nand UO_638 (O_638,N_4550,N_4830);
or UO_639 (O_639,N_4600,N_4646);
and UO_640 (O_640,N_4885,N_4646);
xor UO_641 (O_641,N_4720,N_4878);
or UO_642 (O_642,N_4641,N_4540);
xnor UO_643 (O_643,N_4554,N_4564);
or UO_644 (O_644,N_4873,N_4672);
nor UO_645 (O_645,N_4859,N_4908);
nor UO_646 (O_646,N_4767,N_4646);
xor UO_647 (O_647,N_4501,N_4748);
nand UO_648 (O_648,N_4506,N_4653);
xor UO_649 (O_649,N_4712,N_4699);
xnor UO_650 (O_650,N_4989,N_4828);
nand UO_651 (O_651,N_4587,N_4692);
or UO_652 (O_652,N_4614,N_4587);
nor UO_653 (O_653,N_4876,N_4531);
nor UO_654 (O_654,N_4580,N_4674);
and UO_655 (O_655,N_4818,N_4769);
or UO_656 (O_656,N_4771,N_4534);
or UO_657 (O_657,N_4829,N_4926);
nor UO_658 (O_658,N_4593,N_4813);
and UO_659 (O_659,N_4891,N_4518);
or UO_660 (O_660,N_4864,N_4734);
nor UO_661 (O_661,N_4755,N_4693);
nor UO_662 (O_662,N_4581,N_4692);
xor UO_663 (O_663,N_4804,N_4544);
xnor UO_664 (O_664,N_4913,N_4896);
nor UO_665 (O_665,N_4948,N_4718);
xnor UO_666 (O_666,N_4879,N_4611);
or UO_667 (O_667,N_4904,N_4538);
nor UO_668 (O_668,N_4523,N_4620);
nand UO_669 (O_669,N_4556,N_4999);
or UO_670 (O_670,N_4999,N_4621);
or UO_671 (O_671,N_4501,N_4969);
nand UO_672 (O_672,N_4929,N_4864);
or UO_673 (O_673,N_4546,N_4780);
nor UO_674 (O_674,N_4651,N_4555);
nand UO_675 (O_675,N_4646,N_4680);
nand UO_676 (O_676,N_4932,N_4984);
nor UO_677 (O_677,N_4730,N_4802);
nor UO_678 (O_678,N_4844,N_4583);
nor UO_679 (O_679,N_4741,N_4646);
or UO_680 (O_680,N_4604,N_4796);
nand UO_681 (O_681,N_4691,N_4942);
nor UO_682 (O_682,N_4539,N_4898);
and UO_683 (O_683,N_4825,N_4697);
nand UO_684 (O_684,N_4663,N_4928);
nor UO_685 (O_685,N_4895,N_4680);
xor UO_686 (O_686,N_4869,N_4690);
nand UO_687 (O_687,N_4911,N_4549);
xor UO_688 (O_688,N_4585,N_4500);
or UO_689 (O_689,N_4914,N_4778);
or UO_690 (O_690,N_4945,N_4924);
nand UO_691 (O_691,N_4880,N_4692);
and UO_692 (O_692,N_4655,N_4538);
nand UO_693 (O_693,N_4865,N_4815);
xnor UO_694 (O_694,N_4857,N_4738);
xnor UO_695 (O_695,N_4999,N_4551);
xnor UO_696 (O_696,N_4706,N_4572);
nor UO_697 (O_697,N_4898,N_4893);
and UO_698 (O_698,N_4948,N_4567);
or UO_699 (O_699,N_4641,N_4557);
or UO_700 (O_700,N_4581,N_4665);
nand UO_701 (O_701,N_4823,N_4990);
and UO_702 (O_702,N_4510,N_4992);
xnor UO_703 (O_703,N_4573,N_4504);
xnor UO_704 (O_704,N_4822,N_4735);
xnor UO_705 (O_705,N_4829,N_4823);
nor UO_706 (O_706,N_4626,N_4888);
or UO_707 (O_707,N_4762,N_4635);
nand UO_708 (O_708,N_4835,N_4916);
nand UO_709 (O_709,N_4785,N_4680);
xnor UO_710 (O_710,N_4547,N_4597);
nor UO_711 (O_711,N_4826,N_4557);
xor UO_712 (O_712,N_4842,N_4871);
nor UO_713 (O_713,N_4652,N_4511);
xor UO_714 (O_714,N_4748,N_4638);
and UO_715 (O_715,N_4634,N_4581);
nor UO_716 (O_716,N_4722,N_4581);
and UO_717 (O_717,N_4697,N_4974);
xor UO_718 (O_718,N_4731,N_4961);
and UO_719 (O_719,N_4818,N_4820);
nand UO_720 (O_720,N_4818,N_4685);
or UO_721 (O_721,N_4788,N_4540);
nor UO_722 (O_722,N_4746,N_4858);
nor UO_723 (O_723,N_4911,N_4642);
and UO_724 (O_724,N_4695,N_4609);
nand UO_725 (O_725,N_4685,N_4741);
and UO_726 (O_726,N_4573,N_4602);
and UO_727 (O_727,N_4978,N_4555);
nand UO_728 (O_728,N_4655,N_4729);
nand UO_729 (O_729,N_4745,N_4741);
or UO_730 (O_730,N_4962,N_4938);
or UO_731 (O_731,N_4581,N_4844);
and UO_732 (O_732,N_4719,N_4565);
and UO_733 (O_733,N_4575,N_4649);
nor UO_734 (O_734,N_4660,N_4759);
and UO_735 (O_735,N_4524,N_4539);
xor UO_736 (O_736,N_4830,N_4634);
and UO_737 (O_737,N_4554,N_4702);
or UO_738 (O_738,N_4901,N_4706);
or UO_739 (O_739,N_4831,N_4661);
nand UO_740 (O_740,N_4766,N_4791);
and UO_741 (O_741,N_4691,N_4704);
or UO_742 (O_742,N_4670,N_4504);
nand UO_743 (O_743,N_4993,N_4963);
nor UO_744 (O_744,N_4814,N_4508);
nand UO_745 (O_745,N_4542,N_4843);
or UO_746 (O_746,N_4809,N_4875);
nor UO_747 (O_747,N_4807,N_4974);
or UO_748 (O_748,N_4608,N_4706);
nand UO_749 (O_749,N_4666,N_4763);
or UO_750 (O_750,N_4542,N_4948);
nor UO_751 (O_751,N_4582,N_4699);
and UO_752 (O_752,N_4611,N_4968);
xnor UO_753 (O_753,N_4587,N_4500);
and UO_754 (O_754,N_4804,N_4892);
nor UO_755 (O_755,N_4810,N_4948);
nor UO_756 (O_756,N_4607,N_4655);
xnor UO_757 (O_757,N_4848,N_4752);
nand UO_758 (O_758,N_4809,N_4797);
nor UO_759 (O_759,N_4722,N_4857);
nor UO_760 (O_760,N_4785,N_4760);
nand UO_761 (O_761,N_4500,N_4565);
xor UO_762 (O_762,N_4763,N_4816);
and UO_763 (O_763,N_4602,N_4680);
xor UO_764 (O_764,N_4539,N_4712);
xor UO_765 (O_765,N_4896,N_4833);
and UO_766 (O_766,N_4594,N_4778);
and UO_767 (O_767,N_4576,N_4737);
or UO_768 (O_768,N_4911,N_4561);
or UO_769 (O_769,N_4979,N_4620);
and UO_770 (O_770,N_4608,N_4869);
and UO_771 (O_771,N_4633,N_4893);
nand UO_772 (O_772,N_4611,N_4571);
and UO_773 (O_773,N_4959,N_4926);
and UO_774 (O_774,N_4750,N_4795);
nand UO_775 (O_775,N_4628,N_4600);
and UO_776 (O_776,N_4841,N_4609);
xnor UO_777 (O_777,N_4713,N_4581);
or UO_778 (O_778,N_4630,N_4681);
and UO_779 (O_779,N_4691,N_4651);
xnor UO_780 (O_780,N_4906,N_4983);
xor UO_781 (O_781,N_4937,N_4776);
nand UO_782 (O_782,N_4870,N_4971);
nand UO_783 (O_783,N_4833,N_4618);
nand UO_784 (O_784,N_4728,N_4842);
xor UO_785 (O_785,N_4765,N_4689);
or UO_786 (O_786,N_4878,N_4862);
nand UO_787 (O_787,N_4744,N_4707);
nor UO_788 (O_788,N_4959,N_4962);
and UO_789 (O_789,N_4835,N_4802);
xnor UO_790 (O_790,N_4729,N_4746);
or UO_791 (O_791,N_4643,N_4710);
or UO_792 (O_792,N_4853,N_4531);
nor UO_793 (O_793,N_4867,N_4903);
or UO_794 (O_794,N_4631,N_4835);
nor UO_795 (O_795,N_4672,N_4591);
and UO_796 (O_796,N_4573,N_4646);
nand UO_797 (O_797,N_4904,N_4631);
nor UO_798 (O_798,N_4971,N_4707);
nor UO_799 (O_799,N_4793,N_4755);
or UO_800 (O_800,N_4504,N_4754);
nor UO_801 (O_801,N_4907,N_4781);
nor UO_802 (O_802,N_4676,N_4962);
nor UO_803 (O_803,N_4701,N_4671);
xnor UO_804 (O_804,N_4671,N_4904);
or UO_805 (O_805,N_4718,N_4830);
nor UO_806 (O_806,N_4701,N_4871);
nor UO_807 (O_807,N_4732,N_4993);
and UO_808 (O_808,N_4655,N_4866);
nor UO_809 (O_809,N_4850,N_4802);
or UO_810 (O_810,N_4682,N_4528);
nand UO_811 (O_811,N_4630,N_4638);
nor UO_812 (O_812,N_4559,N_4758);
or UO_813 (O_813,N_4566,N_4516);
and UO_814 (O_814,N_4657,N_4984);
or UO_815 (O_815,N_4912,N_4557);
and UO_816 (O_816,N_4620,N_4613);
or UO_817 (O_817,N_4675,N_4912);
or UO_818 (O_818,N_4997,N_4719);
nor UO_819 (O_819,N_4860,N_4728);
nand UO_820 (O_820,N_4726,N_4640);
xor UO_821 (O_821,N_4847,N_4675);
or UO_822 (O_822,N_4987,N_4802);
and UO_823 (O_823,N_4873,N_4972);
or UO_824 (O_824,N_4695,N_4935);
nor UO_825 (O_825,N_4556,N_4872);
or UO_826 (O_826,N_4540,N_4672);
xor UO_827 (O_827,N_4774,N_4777);
and UO_828 (O_828,N_4712,N_4698);
or UO_829 (O_829,N_4834,N_4696);
and UO_830 (O_830,N_4745,N_4640);
or UO_831 (O_831,N_4507,N_4644);
or UO_832 (O_832,N_4874,N_4900);
or UO_833 (O_833,N_4698,N_4802);
nor UO_834 (O_834,N_4684,N_4738);
xor UO_835 (O_835,N_4523,N_4799);
xnor UO_836 (O_836,N_4630,N_4859);
nand UO_837 (O_837,N_4758,N_4951);
and UO_838 (O_838,N_4582,N_4503);
or UO_839 (O_839,N_4983,N_4974);
nand UO_840 (O_840,N_4851,N_4890);
nand UO_841 (O_841,N_4630,N_4811);
xor UO_842 (O_842,N_4729,N_4986);
and UO_843 (O_843,N_4718,N_4997);
and UO_844 (O_844,N_4836,N_4644);
nand UO_845 (O_845,N_4582,N_4670);
xor UO_846 (O_846,N_4671,N_4567);
or UO_847 (O_847,N_4580,N_4842);
and UO_848 (O_848,N_4843,N_4849);
and UO_849 (O_849,N_4625,N_4741);
nand UO_850 (O_850,N_4676,N_4577);
or UO_851 (O_851,N_4850,N_4861);
nand UO_852 (O_852,N_4882,N_4641);
xor UO_853 (O_853,N_4976,N_4909);
xnor UO_854 (O_854,N_4965,N_4518);
nand UO_855 (O_855,N_4509,N_4892);
nand UO_856 (O_856,N_4632,N_4596);
nor UO_857 (O_857,N_4514,N_4771);
nand UO_858 (O_858,N_4985,N_4901);
or UO_859 (O_859,N_4761,N_4548);
nand UO_860 (O_860,N_4890,N_4581);
nor UO_861 (O_861,N_4630,N_4906);
nand UO_862 (O_862,N_4832,N_4535);
nand UO_863 (O_863,N_4755,N_4961);
nor UO_864 (O_864,N_4589,N_4630);
nor UO_865 (O_865,N_4701,N_4589);
or UO_866 (O_866,N_4692,N_4673);
nand UO_867 (O_867,N_4953,N_4800);
xor UO_868 (O_868,N_4874,N_4936);
nand UO_869 (O_869,N_4636,N_4665);
nor UO_870 (O_870,N_4679,N_4623);
nor UO_871 (O_871,N_4658,N_4607);
and UO_872 (O_872,N_4962,N_4529);
nand UO_873 (O_873,N_4623,N_4787);
xor UO_874 (O_874,N_4694,N_4760);
nand UO_875 (O_875,N_4608,N_4579);
nor UO_876 (O_876,N_4999,N_4882);
xor UO_877 (O_877,N_4833,N_4577);
or UO_878 (O_878,N_4702,N_4562);
nor UO_879 (O_879,N_4639,N_4753);
and UO_880 (O_880,N_4751,N_4905);
or UO_881 (O_881,N_4694,N_4622);
and UO_882 (O_882,N_4809,N_4704);
nand UO_883 (O_883,N_4909,N_4896);
xnor UO_884 (O_884,N_4974,N_4562);
xnor UO_885 (O_885,N_4569,N_4798);
or UO_886 (O_886,N_4510,N_4935);
nor UO_887 (O_887,N_4523,N_4804);
or UO_888 (O_888,N_4747,N_4934);
or UO_889 (O_889,N_4993,N_4653);
nor UO_890 (O_890,N_4757,N_4832);
or UO_891 (O_891,N_4545,N_4770);
and UO_892 (O_892,N_4860,N_4932);
nor UO_893 (O_893,N_4799,N_4975);
xor UO_894 (O_894,N_4951,N_4529);
and UO_895 (O_895,N_4912,N_4616);
and UO_896 (O_896,N_4884,N_4753);
nand UO_897 (O_897,N_4581,N_4850);
xnor UO_898 (O_898,N_4628,N_4635);
or UO_899 (O_899,N_4766,N_4984);
or UO_900 (O_900,N_4954,N_4551);
nand UO_901 (O_901,N_4563,N_4730);
or UO_902 (O_902,N_4744,N_4799);
and UO_903 (O_903,N_4641,N_4651);
xor UO_904 (O_904,N_4618,N_4729);
or UO_905 (O_905,N_4531,N_4855);
xor UO_906 (O_906,N_4801,N_4576);
nor UO_907 (O_907,N_4956,N_4639);
or UO_908 (O_908,N_4598,N_4707);
xor UO_909 (O_909,N_4817,N_4960);
nand UO_910 (O_910,N_4597,N_4527);
and UO_911 (O_911,N_4817,N_4747);
nor UO_912 (O_912,N_4583,N_4552);
nor UO_913 (O_913,N_4728,N_4643);
nor UO_914 (O_914,N_4575,N_4691);
nor UO_915 (O_915,N_4815,N_4617);
and UO_916 (O_916,N_4907,N_4637);
nor UO_917 (O_917,N_4968,N_4834);
nor UO_918 (O_918,N_4996,N_4529);
xnor UO_919 (O_919,N_4507,N_4665);
nand UO_920 (O_920,N_4562,N_4759);
or UO_921 (O_921,N_4665,N_4654);
and UO_922 (O_922,N_4590,N_4521);
and UO_923 (O_923,N_4771,N_4849);
nand UO_924 (O_924,N_4636,N_4820);
or UO_925 (O_925,N_4869,N_4850);
xnor UO_926 (O_926,N_4644,N_4666);
nor UO_927 (O_927,N_4786,N_4646);
nor UO_928 (O_928,N_4818,N_4506);
and UO_929 (O_929,N_4955,N_4848);
nand UO_930 (O_930,N_4926,N_4983);
and UO_931 (O_931,N_4609,N_4928);
nor UO_932 (O_932,N_4544,N_4527);
or UO_933 (O_933,N_4907,N_4846);
or UO_934 (O_934,N_4823,N_4752);
or UO_935 (O_935,N_4824,N_4834);
and UO_936 (O_936,N_4955,N_4818);
nor UO_937 (O_937,N_4931,N_4640);
and UO_938 (O_938,N_4843,N_4627);
nand UO_939 (O_939,N_4605,N_4735);
nand UO_940 (O_940,N_4805,N_4527);
or UO_941 (O_941,N_4787,N_4886);
xor UO_942 (O_942,N_4756,N_4712);
xnor UO_943 (O_943,N_4652,N_4737);
nor UO_944 (O_944,N_4605,N_4718);
and UO_945 (O_945,N_4601,N_4779);
xor UO_946 (O_946,N_4588,N_4853);
xor UO_947 (O_947,N_4605,N_4540);
nor UO_948 (O_948,N_4768,N_4513);
and UO_949 (O_949,N_4847,N_4698);
nor UO_950 (O_950,N_4753,N_4954);
or UO_951 (O_951,N_4856,N_4932);
xnor UO_952 (O_952,N_4500,N_4895);
and UO_953 (O_953,N_4891,N_4570);
or UO_954 (O_954,N_4924,N_4654);
nand UO_955 (O_955,N_4516,N_4835);
or UO_956 (O_956,N_4518,N_4706);
nor UO_957 (O_957,N_4668,N_4979);
nand UO_958 (O_958,N_4625,N_4706);
nor UO_959 (O_959,N_4764,N_4842);
nand UO_960 (O_960,N_4720,N_4831);
and UO_961 (O_961,N_4591,N_4503);
or UO_962 (O_962,N_4913,N_4542);
or UO_963 (O_963,N_4762,N_4974);
or UO_964 (O_964,N_4526,N_4977);
nor UO_965 (O_965,N_4719,N_4894);
nor UO_966 (O_966,N_4910,N_4742);
nand UO_967 (O_967,N_4701,N_4849);
and UO_968 (O_968,N_4525,N_4662);
or UO_969 (O_969,N_4588,N_4965);
nand UO_970 (O_970,N_4818,N_4895);
xor UO_971 (O_971,N_4794,N_4749);
xor UO_972 (O_972,N_4693,N_4632);
xor UO_973 (O_973,N_4604,N_4682);
nor UO_974 (O_974,N_4762,N_4728);
and UO_975 (O_975,N_4669,N_4725);
and UO_976 (O_976,N_4542,N_4860);
xnor UO_977 (O_977,N_4830,N_4705);
nor UO_978 (O_978,N_4930,N_4574);
nand UO_979 (O_979,N_4998,N_4673);
xnor UO_980 (O_980,N_4851,N_4959);
and UO_981 (O_981,N_4824,N_4900);
xor UO_982 (O_982,N_4993,N_4778);
nand UO_983 (O_983,N_4527,N_4960);
nand UO_984 (O_984,N_4732,N_4672);
nor UO_985 (O_985,N_4971,N_4569);
xnor UO_986 (O_986,N_4686,N_4956);
or UO_987 (O_987,N_4760,N_4829);
and UO_988 (O_988,N_4804,N_4558);
xor UO_989 (O_989,N_4838,N_4678);
xor UO_990 (O_990,N_4682,N_4881);
nor UO_991 (O_991,N_4916,N_4912);
nor UO_992 (O_992,N_4552,N_4559);
nor UO_993 (O_993,N_4503,N_4542);
or UO_994 (O_994,N_4860,N_4930);
and UO_995 (O_995,N_4940,N_4521);
nand UO_996 (O_996,N_4556,N_4764);
and UO_997 (O_997,N_4511,N_4760);
xnor UO_998 (O_998,N_4841,N_4707);
nand UO_999 (O_999,N_4614,N_4811);
endmodule