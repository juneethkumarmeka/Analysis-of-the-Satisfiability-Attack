module basic_500_3000_500_30_levels_2xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_469,In_309);
nor U1 (N_1,In_45,In_389);
or U2 (N_2,In_166,In_449);
nand U3 (N_3,In_262,In_441);
nand U4 (N_4,In_12,In_418);
and U5 (N_5,In_326,In_303);
nor U6 (N_6,In_382,In_125);
nor U7 (N_7,In_398,In_76);
nor U8 (N_8,In_77,In_132);
nand U9 (N_9,In_481,In_457);
or U10 (N_10,In_150,In_133);
and U11 (N_11,In_446,In_58);
nor U12 (N_12,In_206,In_37);
nor U13 (N_13,In_71,In_474);
or U14 (N_14,In_270,In_95);
and U15 (N_15,In_113,In_250);
nand U16 (N_16,In_184,In_280);
nand U17 (N_17,In_232,In_185);
or U18 (N_18,In_152,In_233);
nor U19 (N_19,In_222,In_484);
or U20 (N_20,In_43,In_147);
nor U21 (N_21,In_117,In_290);
nand U22 (N_22,In_317,In_293);
nor U23 (N_23,In_458,In_301);
nor U24 (N_24,In_492,In_9);
nand U25 (N_25,In_41,In_489);
or U26 (N_26,In_494,In_91);
nand U27 (N_27,In_347,In_116);
xnor U28 (N_28,In_306,In_288);
or U29 (N_29,In_35,In_496);
and U30 (N_30,In_115,In_50);
nand U31 (N_31,In_221,In_148);
and U32 (N_32,In_238,In_213);
and U33 (N_33,In_159,In_413);
or U34 (N_34,In_248,In_64);
and U35 (N_35,In_102,In_103);
or U36 (N_36,In_209,In_371);
or U37 (N_37,In_465,In_427);
nor U38 (N_38,In_15,In_245);
or U39 (N_39,In_453,In_359);
or U40 (N_40,In_271,In_214);
or U41 (N_41,In_193,In_459);
nor U42 (N_42,In_257,In_331);
nor U43 (N_43,In_395,In_32);
nand U44 (N_44,In_447,In_190);
nor U45 (N_45,In_111,In_487);
nand U46 (N_46,In_131,In_188);
or U47 (N_47,In_439,In_333);
nand U48 (N_48,In_471,In_94);
nor U49 (N_49,In_33,In_176);
or U50 (N_50,In_160,In_315);
and U51 (N_51,In_320,In_414);
nand U52 (N_52,In_313,In_302);
or U53 (N_53,In_143,In_51);
and U54 (N_54,In_468,In_140);
nor U55 (N_55,In_251,In_341);
nand U56 (N_56,In_234,In_400);
nor U57 (N_57,In_377,In_443);
nand U58 (N_58,In_174,In_63);
and U59 (N_59,In_92,In_304);
nand U60 (N_60,In_155,In_365);
or U61 (N_61,In_224,In_460);
nand U62 (N_62,In_110,In_6);
nand U63 (N_63,In_67,In_139);
or U64 (N_64,In_380,In_287);
and U65 (N_65,In_401,In_119);
nor U66 (N_66,In_438,In_65);
xnor U67 (N_67,In_219,In_429);
or U68 (N_68,In_196,In_24);
and U69 (N_69,In_416,In_226);
nand U70 (N_70,In_210,In_467);
or U71 (N_71,In_450,In_114);
nor U72 (N_72,In_411,In_23);
and U73 (N_73,In_292,In_229);
nand U74 (N_74,In_370,In_483);
and U75 (N_75,In_73,In_87);
or U76 (N_76,In_191,In_476);
and U77 (N_77,In_274,In_410);
nand U78 (N_78,In_26,In_495);
or U79 (N_79,In_19,In_375);
or U80 (N_80,In_345,In_212);
nand U81 (N_81,In_454,In_109);
or U82 (N_82,In_249,In_85);
and U83 (N_83,In_104,In_408);
nor U84 (N_84,In_479,In_181);
nand U85 (N_85,In_175,In_129);
nand U86 (N_86,In_216,In_300);
nand U87 (N_87,In_311,In_38);
nor U88 (N_88,In_462,In_463);
nand U89 (N_89,In_8,In_156);
nor U90 (N_90,In_170,In_118);
xor U91 (N_91,In_217,In_151);
or U92 (N_92,In_225,In_373);
or U93 (N_93,In_440,In_349);
nor U94 (N_94,In_338,In_81);
nand U95 (N_95,In_464,In_430);
nor U96 (N_96,In_25,In_253);
xor U97 (N_97,In_261,In_165);
or U98 (N_98,In_218,In_357);
and U99 (N_99,In_491,In_407);
nor U100 (N_100,In_36,N_45);
and U101 (N_101,In_437,In_88);
nor U102 (N_102,In_436,N_26);
or U103 (N_103,In_265,N_50);
and U104 (N_104,In_172,In_5);
or U105 (N_105,In_74,N_27);
and U106 (N_106,N_83,In_296);
and U107 (N_107,In_242,In_391);
or U108 (N_108,N_89,In_305);
and U109 (N_109,In_383,In_272);
or U110 (N_110,In_426,In_402);
nand U111 (N_111,In_268,In_478);
and U112 (N_112,In_252,N_0);
nand U113 (N_113,In_40,In_381);
nand U114 (N_114,In_163,In_2);
and U115 (N_115,In_387,In_186);
and U116 (N_116,In_142,N_40);
nor U117 (N_117,N_24,In_455);
and U118 (N_118,In_100,N_87);
nand U119 (N_119,In_348,In_84);
nor U120 (N_120,N_66,In_211);
xor U121 (N_121,In_66,In_278);
nand U122 (N_122,In_86,N_55);
xnor U123 (N_123,N_79,In_161);
nand U124 (N_124,In_445,In_256);
nor U125 (N_125,In_195,In_145);
or U126 (N_126,N_22,In_497);
nor U127 (N_127,In_403,In_379);
nand U128 (N_128,In_158,In_204);
nand U129 (N_129,N_15,In_169);
nand U130 (N_130,N_49,In_361);
nand U131 (N_131,N_34,In_397);
and U132 (N_132,In_404,In_82);
nand U133 (N_133,In_28,In_0);
nand U134 (N_134,In_263,In_243);
nor U135 (N_135,N_63,In_281);
and U136 (N_136,In_10,In_98);
nor U137 (N_137,In_178,In_390);
or U138 (N_138,In_39,In_294);
or U139 (N_139,In_260,In_363);
nand U140 (N_140,In_126,In_275);
and U141 (N_141,N_69,In_336);
nor U142 (N_142,In_157,In_422);
xnor U143 (N_143,N_51,N_18);
nor U144 (N_144,In_324,In_374);
or U145 (N_145,In_419,In_202);
and U146 (N_146,In_255,In_13);
and U147 (N_147,In_69,In_187);
and U148 (N_148,In_325,In_442);
nor U149 (N_149,In_415,In_332);
or U150 (N_150,N_81,In_291);
nor U151 (N_151,In_197,N_37);
nor U152 (N_152,In_354,In_428);
and U153 (N_153,In_246,In_388);
and U154 (N_154,In_4,In_189);
and U155 (N_155,N_96,In_396);
or U156 (N_156,In_490,In_120);
and U157 (N_157,In_72,In_171);
or U158 (N_158,N_48,N_12);
xor U159 (N_159,N_20,N_28);
nand U160 (N_160,In_231,In_499);
nor U161 (N_161,In_282,N_90);
nand U162 (N_162,In_392,In_141);
xor U163 (N_163,N_13,N_4);
and U164 (N_164,N_6,In_48);
and U165 (N_165,In_298,N_8);
and U166 (N_166,In_208,In_97);
nand U167 (N_167,In_394,In_54);
and U168 (N_168,In_376,In_328);
nand U169 (N_169,N_77,N_57);
and U170 (N_170,In_399,In_179);
and U171 (N_171,In_137,In_486);
nor U172 (N_172,N_73,In_127);
nand U173 (N_173,In_29,In_488);
or U174 (N_174,In_386,In_482);
or U175 (N_175,In_475,In_17);
or U176 (N_176,In_96,In_277);
nor U177 (N_177,In_254,In_307);
or U178 (N_178,In_409,In_144);
nor U179 (N_179,N_32,In_107);
or U180 (N_180,N_72,In_14);
nand U181 (N_181,N_68,In_31);
nor U182 (N_182,In_472,In_283);
nand U183 (N_183,N_3,In_424);
nand U184 (N_184,In_167,In_205);
or U185 (N_185,In_378,N_25);
or U186 (N_186,In_228,In_11);
nand U187 (N_187,N_39,In_90);
nor U188 (N_188,In_337,N_61);
and U189 (N_189,In_89,In_55);
nor U190 (N_190,In_344,In_346);
and U191 (N_191,In_168,N_56);
or U192 (N_192,In_203,In_16);
nor U193 (N_193,In_61,N_47);
nand U194 (N_194,In_201,In_200);
nor U195 (N_195,In_227,In_123);
nand U196 (N_196,In_49,In_339);
or U197 (N_197,In_405,In_372);
nand U198 (N_198,In_106,In_417);
nand U199 (N_199,In_406,N_16);
xnor U200 (N_200,N_88,N_155);
nor U201 (N_201,In_319,N_186);
and U202 (N_202,In_192,N_84);
nor U203 (N_203,N_193,N_120);
or U204 (N_204,In_470,N_151);
nand U205 (N_205,In_273,In_180);
nand U206 (N_206,N_122,In_59);
or U207 (N_207,N_173,In_352);
or U208 (N_208,In_461,In_295);
nand U209 (N_209,In_30,In_78);
and U210 (N_210,N_54,In_485);
nor U211 (N_211,N_117,In_57);
nand U212 (N_212,N_38,N_108);
and U213 (N_213,N_182,N_97);
nand U214 (N_214,In_299,In_34);
or U215 (N_215,N_195,In_334);
or U216 (N_216,N_1,In_149);
nor U217 (N_217,In_70,N_17);
and U218 (N_218,N_94,In_435);
and U219 (N_219,N_181,N_78);
or U220 (N_220,N_110,In_289);
nor U221 (N_221,In_138,N_198);
or U222 (N_222,N_180,N_189);
xor U223 (N_223,In_360,In_244);
or U224 (N_224,In_369,N_152);
or U225 (N_225,In_385,In_285);
nand U226 (N_226,In_177,N_169);
nor U227 (N_227,N_146,In_101);
nor U228 (N_228,In_321,In_420);
or U229 (N_229,N_145,In_135);
and U230 (N_230,N_147,N_35);
and U231 (N_231,In_456,N_143);
xor U232 (N_232,N_76,N_53);
nand U233 (N_233,N_21,In_47);
or U234 (N_234,In_318,In_215);
and U235 (N_235,In_473,N_184);
and U236 (N_236,In_356,In_93);
or U237 (N_237,N_23,N_102);
nor U238 (N_238,N_41,In_79);
nor U239 (N_239,In_182,N_118);
nor U240 (N_240,N_9,N_163);
nand U241 (N_241,N_46,N_177);
and U242 (N_242,In_134,N_70);
nand U243 (N_243,N_123,In_60);
or U244 (N_244,N_149,N_139);
or U245 (N_245,N_159,In_42);
or U246 (N_246,N_119,In_362);
or U247 (N_247,N_105,In_237);
or U248 (N_248,In_266,N_175);
nor U249 (N_249,In_308,In_112);
nand U250 (N_250,N_140,N_199);
or U251 (N_251,N_80,N_134);
and U252 (N_252,In_432,In_183);
and U253 (N_253,In_122,In_162);
nor U254 (N_254,In_75,In_284);
and U255 (N_255,N_116,N_125);
or U256 (N_256,In_53,In_46);
or U257 (N_257,N_101,In_153);
and U258 (N_258,N_95,N_104);
nand U259 (N_259,N_59,N_67);
nor U260 (N_260,N_167,N_86);
and U261 (N_261,In_198,N_142);
and U262 (N_262,In_342,In_366);
and U263 (N_263,N_52,N_115);
nor U264 (N_264,In_279,In_247);
or U265 (N_265,In_56,In_27);
nand U266 (N_266,In_316,In_310);
or U267 (N_267,In_80,N_127);
or U268 (N_268,In_146,In_358);
or U269 (N_269,In_164,N_153);
nor U270 (N_270,In_433,N_10);
nor U271 (N_271,N_141,N_31);
nor U272 (N_272,In_276,N_64);
or U273 (N_273,N_99,In_444);
or U274 (N_274,In_421,In_18);
or U275 (N_275,N_168,In_314);
and U276 (N_276,N_36,In_21);
and U277 (N_277,N_7,N_190);
nand U278 (N_278,N_107,N_157);
xnor U279 (N_279,In_384,In_173);
nand U280 (N_280,N_44,N_136);
and U281 (N_281,N_188,In_393);
nand U282 (N_282,N_130,N_92);
nor U283 (N_283,In_312,In_351);
and U284 (N_284,N_161,N_58);
nor U285 (N_285,N_62,N_196);
nor U286 (N_286,N_128,In_269);
nand U287 (N_287,N_106,N_100);
or U288 (N_288,N_93,In_136);
nand U289 (N_289,N_187,N_98);
nor U290 (N_290,In_452,N_138);
and U291 (N_291,In_322,N_109);
or U292 (N_292,N_126,N_150);
xor U293 (N_293,N_185,N_103);
xor U294 (N_294,N_124,N_132);
nor U295 (N_295,N_170,In_340);
or U296 (N_296,N_82,In_236);
and U297 (N_297,N_19,In_286);
nor U298 (N_298,In_194,N_75);
nand U299 (N_299,In_68,In_207);
or U300 (N_300,N_156,N_158);
or U301 (N_301,N_165,N_204);
nor U302 (N_302,N_203,N_220);
nand U303 (N_303,In_367,N_11);
nor U304 (N_304,In_220,N_240);
and U305 (N_305,N_239,N_292);
xnor U306 (N_306,N_164,N_231);
or U307 (N_307,N_278,N_283);
or U308 (N_308,In_124,N_275);
nand U309 (N_309,N_297,N_246);
or U310 (N_310,N_191,In_199);
and U311 (N_311,In_498,N_285);
nand U312 (N_312,In_99,N_284);
and U313 (N_313,In_105,N_176);
nor U314 (N_314,In_128,In_259);
and U315 (N_315,In_466,N_29);
or U316 (N_316,N_248,N_250);
nand U317 (N_317,N_74,N_295);
nor U318 (N_318,N_296,In_240);
or U319 (N_319,N_282,N_257);
nor U320 (N_320,N_260,N_227);
and U321 (N_321,N_215,N_251);
nand U322 (N_322,In_258,N_294);
or U323 (N_323,N_254,N_154);
and U324 (N_324,In_297,In_323);
nor U325 (N_325,In_108,N_207);
and U326 (N_326,N_270,N_226);
nand U327 (N_327,N_194,N_111);
nor U328 (N_328,N_233,In_7);
nor U329 (N_329,N_243,N_205);
and U330 (N_330,N_249,N_213);
or U331 (N_331,N_113,N_162);
nor U332 (N_332,In_368,In_353);
nand U333 (N_333,N_277,In_52);
nand U334 (N_334,N_280,N_148);
or U335 (N_335,In_1,In_83);
nand U336 (N_336,N_252,In_121);
nand U337 (N_337,N_131,N_121);
nor U338 (N_338,N_179,N_267);
nand U339 (N_339,N_133,In_335);
nand U340 (N_340,N_230,In_62);
nand U341 (N_341,N_172,N_241);
and U342 (N_342,In_241,N_30);
nand U343 (N_343,In_477,N_228);
nor U344 (N_344,In_327,N_291);
nor U345 (N_345,In_44,In_451);
or U346 (N_346,N_247,N_229);
or U347 (N_347,N_258,N_236);
and U348 (N_348,N_279,N_268);
nand U349 (N_349,N_289,N_299);
or U350 (N_350,N_221,N_264);
or U351 (N_351,N_212,In_230);
or U352 (N_352,In_329,N_71);
or U353 (N_353,In_355,N_206);
nor U354 (N_354,N_201,N_2);
nand U355 (N_355,N_224,In_235);
nand U356 (N_356,N_276,N_286);
nand U357 (N_357,N_166,N_253);
nand U358 (N_358,In_412,N_298);
nand U359 (N_359,N_262,N_200);
and U360 (N_360,N_42,N_211);
nor U361 (N_361,In_22,N_214);
nand U362 (N_362,N_287,In_493);
nand U363 (N_363,N_225,In_350);
or U364 (N_364,N_43,N_245);
nor U365 (N_365,N_192,N_210);
nor U366 (N_366,N_114,N_174);
and U367 (N_367,In_448,N_255);
nor U368 (N_368,N_217,N_129);
nand U369 (N_369,In_154,N_263);
and U370 (N_370,N_216,N_272);
and U371 (N_371,N_171,N_242);
and U372 (N_372,N_290,N_274);
nor U373 (N_373,In_264,In_480);
and U374 (N_374,In_434,N_271);
and U375 (N_375,N_208,N_91);
nor U376 (N_376,In_239,In_223);
nor U377 (N_377,In_330,N_238);
and U378 (N_378,N_261,N_244);
and U379 (N_379,In_343,In_130);
nor U380 (N_380,N_269,N_265);
or U381 (N_381,In_364,In_425);
and U382 (N_382,N_234,N_85);
nand U383 (N_383,In_431,N_65);
nand U384 (N_384,N_5,N_222);
nor U385 (N_385,N_273,N_223);
and U386 (N_386,N_232,N_281);
nor U387 (N_387,N_178,N_293);
and U388 (N_388,N_266,N_135);
or U389 (N_389,N_144,N_288);
nor U390 (N_390,N_219,N_183);
nor U391 (N_391,In_3,N_33);
or U392 (N_392,In_267,In_20);
and U393 (N_393,N_218,N_112);
or U394 (N_394,N_235,N_160);
nand U395 (N_395,N_60,N_259);
nand U396 (N_396,In_423,N_137);
or U397 (N_397,N_202,N_237);
and U398 (N_398,N_209,N_14);
or U399 (N_399,N_197,N_256);
and U400 (N_400,N_314,N_380);
nor U401 (N_401,N_391,N_338);
or U402 (N_402,N_318,N_320);
or U403 (N_403,N_377,N_310);
and U404 (N_404,N_370,N_335);
or U405 (N_405,N_358,N_307);
xnor U406 (N_406,N_383,N_395);
nor U407 (N_407,N_331,N_366);
nor U408 (N_408,N_300,N_349);
nor U409 (N_409,N_305,N_390);
or U410 (N_410,N_302,N_352);
nor U411 (N_411,N_332,N_384);
or U412 (N_412,N_371,N_396);
nor U413 (N_413,N_319,N_367);
nand U414 (N_414,N_336,N_379);
nand U415 (N_415,N_378,N_317);
nor U416 (N_416,N_340,N_389);
or U417 (N_417,N_354,N_327);
nand U418 (N_418,N_372,N_392);
or U419 (N_419,N_334,N_313);
nor U420 (N_420,N_368,N_309);
nand U421 (N_421,N_343,N_394);
nand U422 (N_422,N_324,N_342);
or U423 (N_423,N_375,N_337);
nand U424 (N_424,N_382,N_308);
nand U425 (N_425,N_304,N_353);
or U426 (N_426,N_365,N_323);
or U427 (N_427,N_345,N_329);
and U428 (N_428,N_393,N_328);
nand U429 (N_429,N_325,N_388);
and U430 (N_430,N_350,N_315);
nor U431 (N_431,N_361,N_398);
and U432 (N_432,N_374,N_385);
nand U433 (N_433,N_333,N_397);
nand U434 (N_434,N_330,N_362);
nand U435 (N_435,N_360,N_387);
nand U436 (N_436,N_356,N_326);
nand U437 (N_437,N_321,N_376);
or U438 (N_438,N_339,N_364);
and U439 (N_439,N_301,N_369);
xnor U440 (N_440,N_306,N_363);
nand U441 (N_441,N_351,N_311);
nor U442 (N_442,N_346,N_303);
nor U443 (N_443,N_348,N_341);
or U444 (N_444,N_381,N_344);
and U445 (N_445,N_359,N_312);
nor U446 (N_446,N_355,N_347);
and U447 (N_447,N_322,N_386);
or U448 (N_448,N_316,N_357);
nor U449 (N_449,N_373,N_399);
nand U450 (N_450,N_339,N_354);
or U451 (N_451,N_338,N_335);
nand U452 (N_452,N_358,N_336);
nor U453 (N_453,N_330,N_396);
and U454 (N_454,N_311,N_375);
nand U455 (N_455,N_396,N_326);
and U456 (N_456,N_385,N_379);
nand U457 (N_457,N_353,N_355);
nand U458 (N_458,N_388,N_379);
or U459 (N_459,N_328,N_332);
and U460 (N_460,N_306,N_350);
or U461 (N_461,N_333,N_366);
xnor U462 (N_462,N_335,N_332);
nand U463 (N_463,N_367,N_399);
nand U464 (N_464,N_337,N_356);
nand U465 (N_465,N_359,N_316);
nor U466 (N_466,N_369,N_317);
or U467 (N_467,N_305,N_334);
nand U468 (N_468,N_307,N_384);
nor U469 (N_469,N_376,N_399);
nor U470 (N_470,N_300,N_301);
nor U471 (N_471,N_328,N_369);
and U472 (N_472,N_358,N_309);
nand U473 (N_473,N_397,N_312);
or U474 (N_474,N_369,N_339);
nor U475 (N_475,N_323,N_335);
and U476 (N_476,N_321,N_388);
or U477 (N_477,N_399,N_336);
nor U478 (N_478,N_308,N_390);
nand U479 (N_479,N_310,N_384);
nand U480 (N_480,N_313,N_328);
and U481 (N_481,N_377,N_300);
nor U482 (N_482,N_351,N_354);
nand U483 (N_483,N_342,N_359);
or U484 (N_484,N_371,N_355);
nand U485 (N_485,N_333,N_330);
and U486 (N_486,N_325,N_329);
nor U487 (N_487,N_387,N_355);
or U488 (N_488,N_370,N_389);
nand U489 (N_489,N_358,N_312);
and U490 (N_490,N_340,N_365);
nand U491 (N_491,N_341,N_317);
nand U492 (N_492,N_330,N_356);
and U493 (N_493,N_328,N_379);
nor U494 (N_494,N_320,N_322);
nor U495 (N_495,N_306,N_365);
or U496 (N_496,N_339,N_359);
or U497 (N_497,N_306,N_337);
or U498 (N_498,N_390,N_360);
nand U499 (N_499,N_320,N_314);
or U500 (N_500,N_498,N_434);
nand U501 (N_501,N_435,N_462);
nand U502 (N_502,N_448,N_432);
nand U503 (N_503,N_437,N_486);
and U504 (N_504,N_418,N_417);
and U505 (N_505,N_488,N_410);
or U506 (N_506,N_441,N_427);
and U507 (N_507,N_494,N_458);
or U508 (N_508,N_463,N_466);
or U509 (N_509,N_438,N_474);
or U510 (N_510,N_492,N_426);
nand U511 (N_511,N_467,N_482);
and U512 (N_512,N_496,N_453);
nand U513 (N_513,N_484,N_464);
nor U514 (N_514,N_450,N_440);
nand U515 (N_515,N_476,N_419);
and U516 (N_516,N_493,N_430);
and U517 (N_517,N_491,N_409);
nand U518 (N_518,N_414,N_444);
nor U519 (N_519,N_424,N_459);
nand U520 (N_520,N_469,N_460);
nand U521 (N_521,N_446,N_405);
nor U522 (N_522,N_451,N_449);
nor U523 (N_523,N_497,N_406);
nor U524 (N_524,N_431,N_468);
and U525 (N_525,N_415,N_421);
and U526 (N_526,N_407,N_411);
nand U527 (N_527,N_428,N_499);
or U528 (N_528,N_470,N_452);
nor U529 (N_529,N_472,N_423);
or U530 (N_530,N_412,N_439);
nand U531 (N_531,N_413,N_455);
nand U532 (N_532,N_456,N_429);
and U533 (N_533,N_425,N_457);
nor U534 (N_534,N_471,N_461);
nor U535 (N_535,N_436,N_442);
xor U536 (N_536,N_478,N_420);
nor U537 (N_537,N_408,N_403);
and U538 (N_538,N_402,N_495);
nor U539 (N_539,N_400,N_481);
and U540 (N_540,N_485,N_422);
nor U541 (N_541,N_404,N_433);
nor U542 (N_542,N_445,N_447);
nor U543 (N_543,N_443,N_465);
nor U544 (N_544,N_401,N_416);
and U545 (N_545,N_483,N_479);
nand U546 (N_546,N_489,N_477);
and U547 (N_547,N_480,N_454);
nand U548 (N_548,N_490,N_475);
and U549 (N_549,N_487,N_473);
nor U550 (N_550,N_492,N_461);
and U551 (N_551,N_455,N_408);
nand U552 (N_552,N_446,N_441);
nand U553 (N_553,N_457,N_426);
or U554 (N_554,N_434,N_463);
nand U555 (N_555,N_430,N_403);
nor U556 (N_556,N_415,N_495);
nor U557 (N_557,N_417,N_400);
and U558 (N_558,N_468,N_458);
nor U559 (N_559,N_453,N_460);
or U560 (N_560,N_436,N_452);
and U561 (N_561,N_464,N_476);
or U562 (N_562,N_400,N_436);
and U563 (N_563,N_470,N_423);
or U564 (N_564,N_439,N_447);
or U565 (N_565,N_497,N_491);
nor U566 (N_566,N_471,N_490);
nand U567 (N_567,N_489,N_466);
and U568 (N_568,N_429,N_486);
nor U569 (N_569,N_416,N_442);
or U570 (N_570,N_424,N_435);
and U571 (N_571,N_403,N_400);
nor U572 (N_572,N_490,N_428);
or U573 (N_573,N_400,N_407);
nor U574 (N_574,N_491,N_411);
or U575 (N_575,N_444,N_442);
and U576 (N_576,N_405,N_447);
nor U577 (N_577,N_447,N_414);
and U578 (N_578,N_495,N_445);
and U579 (N_579,N_409,N_417);
nand U580 (N_580,N_401,N_408);
nor U581 (N_581,N_467,N_472);
nand U582 (N_582,N_470,N_446);
or U583 (N_583,N_429,N_451);
nor U584 (N_584,N_460,N_482);
or U585 (N_585,N_453,N_441);
nor U586 (N_586,N_437,N_435);
nand U587 (N_587,N_496,N_419);
and U588 (N_588,N_481,N_441);
or U589 (N_589,N_415,N_406);
nand U590 (N_590,N_408,N_419);
nand U591 (N_591,N_436,N_411);
and U592 (N_592,N_458,N_456);
nand U593 (N_593,N_411,N_464);
nor U594 (N_594,N_421,N_472);
nor U595 (N_595,N_436,N_487);
nand U596 (N_596,N_458,N_485);
nand U597 (N_597,N_452,N_457);
nor U598 (N_598,N_441,N_480);
and U599 (N_599,N_417,N_450);
nand U600 (N_600,N_508,N_511);
nand U601 (N_601,N_523,N_565);
nor U602 (N_602,N_596,N_502);
or U603 (N_603,N_581,N_507);
nor U604 (N_604,N_526,N_589);
and U605 (N_605,N_543,N_572);
or U606 (N_606,N_591,N_549);
or U607 (N_607,N_592,N_524);
or U608 (N_608,N_500,N_527);
nand U609 (N_609,N_521,N_598);
nor U610 (N_610,N_571,N_537);
nand U611 (N_611,N_597,N_529);
and U612 (N_612,N_547,N_530);
nor U613 (N_613,N_552,N_557);
and U614 (N_614,N_566,N_564);
nor U615 (N_615,N_520,N_570);
nor U616 (N_616,N_593,N_568);
or U617 (N_617,N_539,N_545);
nand U618 (N_618,N_510,N_509);
and U619 (N_619,N_594,N_551);
nand U620 (N_620,N_567,N_588);
nand U621 (N_621,N_585,N_519);
or U622 (N_622,N_579,N_516);
nor U623 (N_623,N_569,N_501);
nor U624 (N_624,N_558,N_550);
or U625 (N_625,N_513,N_574);
and U626 (N_626,N_504,N_587);
or U627 (N_627,N_503,N_556);
and U628 (N_628,N_535,N_563);
and U629 (N_629,N_584,N_532);
and U630 (N_630,N_586,N_540);
and U631 (N_631,N_577,N_578);
nand U632 (N_632,N_560,N_522);
or U633 (N_633,N_512,N_534);
nor U634 (N_634,N_517,N_505);
and U635 (N_635,N_544,N_533);
and U636 (N_636,N_590,N_525);
nand U637 (N_637,N_599,N_555);
or U638 (N_638,N_515,N_541);
nor U639 (N_639,N_561,N_548);
and U640 (N_640,N_553,N_518);
nand U641 (N_641,N_583,N_506);
nor U642 (N_642,N_546,N_576);
and U643 (N_643,N_559,N_536);
nand U644 (N_644,N_531,N_542);
or U645 (N_645,N_573,N_538);
and U646 (N_646,N_580,N_582);
nand U647 (N_647,N_595,N_514);
nand U648 (N_648,N_575,N_554);
nand U649 (N_649,N_528,N_562);
xor U650 (N_650,N_595,N_504);
nand U651 (N_651,N_590,N_586);
and U652 (N_652,N_545,N_544);
nand U653 (N_653,N_583,N_517);
xor U654 (N_654,N_563,N_545);
and U655 (N_655,N_563,N_544);
nor U656 (N_656,N_526,N_533);
or U657 (N_657,N_539,N_506);
or U658 (N_658,N_544,N_516);
or U659 (N_659,N_503,N_590);
nand U660 (N_660,N_566,N_573);
nor U661 (N_661,N_583,N_579);
or U662 (N_662,N_533,N_504);
or U663 (N_663,N_596,N_523);
or U664 (N_664,N_519,N_551);
or U665 (N_665,N_583,N_531);
and U666 (N_666,N_508,N_591);
or U667 (N_667,N_507,N_503);
or U668 (N_668,N_540,N_579);
xor U669 (N_669,N_553,N_521);
nand U670 (N_670,N_505,N_529);
nor U671 (N_671,N_532,N_551);
nor U672 (N_672,N_543,N_567);
or U673 (N_673,N_510,N_517);
nand U674 (N_674,N_560,N_507);
or U675 (N_675,N_507,N_504);
nand U676 (N_676,N_524,N_593);
nor U677 (N_677,N_528,N_563);
nor U678 (N_678,N_568,N_598);
and U679 (N_679,N_508,N_532);
and U680 (N_680,N_516,N_529);
nor U681 (N_681,N_539,N_558);
and U682 (N_682,N_502,N_520);
and U683 (N_683,N_555,N_587);
nand U684 (N_684,N_558,N_537);
nand U685 (N_685,N_537,N_511);
or U686 (N_686,N_521,N_599);
or U687 (N_687,N_587,N_534);
and U688 (N_688,N_584,N_505);
and U689 (N_689,N_515,N_560);
nor U690 (N_690,N_509,N_593);
nor U691 (N_691,N_570,N_524);
nand U692 (N_692,N_537,N_559);
or U693 (N_693,N_578,N_584);
or U694 (N_694,N_596,N_539);
nand U695 (N_695,N_533,N_573);
and U696 (N_696,N_530,N_555);
or U697 (N_697,N_588,N_507);
or U698 (N_698,N_588,N_562);
or U699 (N_699,N_547,N_569);
nor U700 (N_700,N_679,N_653);
and U701 (N_701,N_633,N_692);
or U702 (N_702,N_689,N_662);
nand U703 (N_703,N_680,N_688);
and U704 (N_704,N_626,N_685);
or U705 (N_705,N_641,N_621);
nand U706 (N_706,N_619,N_652);
nand U707 (N_707,N_684,N_672);
nor U708 (N_708,N_644,N_620);
and U709 (N_709,N_697,N_664);
and U710 (N_710,N_670,N_624);
nor U711 (N_711,N_650,N_645);
nor U712 (N_712,N_658,N_681);
nand U713 (N_713,N_642,N_687);
nor U714 (N_714,N_659,N_606);
nand U715 (N_715,N_635,N_682);
nor U716 (N_716,N_676,N_647);
or U717 (N_717,N_600,N_637);
nand U718 (N_718,N_604,N_695);
nand U719 (N_719,N_661,N_625);
and U720 (N_720,N_615,N_691);
and U721 (N_721,N_675,N_643);
nand U722 (N_722,N_616,N_663);
or U723 (N_723,N_665,N_686);
xnor U724 (N_724,N_602,N_605);
or U725 (N_725,N_607,N_656);
and U726 (N_726,N_618,N_634);
nand U727 (N_727,N_690,N_636);
nand U728 (N_728,N_648,N_609);
or U729 (N_729,N_654,N_646);
nand U730 (N_730,N_627,N_628);
nand U731 (N_731,N_699,N_630);
and U732 (N_732,N_608,N_683);
nor U733 (N_733,N_603,N_601);
or U734 (N_734,N_667,N_666);
nor U735 (N_735,N_613,N_660);
and U736 (N_736,N_617,N_614);
nand U737 (N_737,N_696,N_649);
nor U738 (N_738,N_629,N_640);
nand U739 (N_739,N_673,N_694);
nand U740 (N_740,N_611,N_668);
nor U741 (N_741,N_631,N_677);
nor U742 (N_742,N_669,N_610);
nor U743 (N_743,N_622,N_678);
nand U744 (N_744,N_651,N_632);
and U745 (N_745,N_693,N_639);
nand U746 (N_746,N_698,N_638);
and U747 (N_747,N_657,N_623);
nor U748 (N_748,N_655,N_674);
nand U749 (N_749,N_671,N_612);
or U750 (N_750,N_691,N_621);
and U751 (N_751,N_633,N_683);
nand U752 (N_752,N_642,N_627);
or U753 (N_753,N_612,N_624);
and U754 (N_754,N_665,N_677);
nor U755 (N_755,N_672,N_669);
or U756 (N_756,N_606,N_692);
nand U757 (N_757,N_615,N_623);
and U758 (N_758,N_673,N_667);
nor U759 (N_759,N_674,N_633);
or U760 (N_760,N_656,N_642);
nand U761 (N_761,N_661,N_650);
nand U762 (N_762,N_608,N_657);
nor U763 (N_763,N_648,N_653);
or U764 (N_764,N_674,N_667);
or U765 (N_765,N_637,N_664);
nor U766 (N_766,N_602,N_645);
and U767 (N_767,N_618,N_679);
and U768 (N_768,N_674,N_658);
nand U769 (N_769,N_681,N_616);
nand U770 (N_770,N_669,N_674);
nor U771 (N_771,N_657,N_660);
and U772 (N_772,N_676,N_686);
and U773 (N_773,N_611,N_648);
xnor U774 (N_774,N_697,N_683);
or U775 (N_775,N_605,N_625);
nor U776 (N_776,N_694,N_663);
and U777 (N_777,N_625,N_628);
nor U778 (N_778,N_617,N_642);
nand U779 (N_779,N_620,N_693);
or U780 (N_780,N_628,N_647);
nand U781 (N_781,N_630,N_658);
nand U782 (N_782,N_604,N_621);
or U783 (N_783,N_666,N_605);
xor U784 (N_784,N_634,N_605);
and U785 (N_785,N_600,N_697);
or U786 (N_786,N_658,N_604);
or U787 (N_787,N_692,N_689);
nor U788 (N_788,N_669,N_699);
nand U789 (N_789,N_689,N_627);
nand U790 (N_790,N_644,N_675);
or U791 (N_791,N_661,N_633);
xnor U792 (N_792,N_625,N_639);
nand U793 (N_793,N_652,N_687);
or U794 (N_794,N_609,N_614);
nor U795 (N_795,N_613,N_646);
and U796 (N_796,N_692,N_605);
nand U797 (N_797,N_646,N_653);
nand U798 (N_798,N_661,N_689);
and U799 (N_799,N_614,N_695);
or U800 (N_800,N_746,N_753);
nand U801 (N_801,N_703,N_771);
nand U802 (N_802,N_745,N_760);
nand U803 (N_803,N_750,N_704);
and U804 (N_804,N_708,N_783);
nand U805 (N_805,N_780,N_735);
nand U806 (N_806,N_742,N_748);
or U807 (N_807,N_736,N_768);
or U808 (N_808,N_751,N_729);
nor U809 (N_809,N_749,N_782);
and U810 (N_810,N_796,N_716);
and U811 (N_811,N_710,N_776);
or U812 (N_812,N_781,N_763);
or U813 (N_813,N_743,N_784);
or U814 (N_814,N_707,N_758);
nand U815 (N_815,N_791,N_769);
nor U816 (N_816,N_793,N_731);
or U817 (N_817,N_792,N_701);
nand U818 (N_818,N_773,N_762);
and U819 (N_819,N_728,N_723);
or U820 (N_820,N_759,N_702);
and U821 (N_821,N_705,N_714);
nand U822 (N_822,N_789,N_717);
nand U823 (N_823,N_715,N_799);
or U824 (N_824,N_752,N_772);
and U825 (N_825,N_770,N_730);
and U826 (N_826,N_764,N_788);
or U827 (N_827,N_777,N_724);
and U828 (N_828,N_755,N_754);
or U829 (N_829,N_774,N_719);
xor U830 (N_830,N_794,N_718);
nor U831 (N_831,N_721,N_741);
nand U832 (N_832,N_727,N_720);
or U833 (N_833,N_725,N_787);
nand U834 (N_834,N_722,N_739);
nor U835 (N_835,N_790,N_775);
nand U836 (N_836,N_785,N_709);
nor U837 (N_837,N_711,N_737);
and U838 (N_838,N_744,N_786);
nand U839 (N_839,N_713,N_712);
or U840 (N_840,N_733,N_767);
and U841 (N_841,N_738,N_756);
nand U842 (N_842,N_766,N_706);
and U843 (N_843,N_765,N_747);
nand U844 (N_844,N_779,N_778);
nand U845 (N_845,N_732,N_734);
nor U846 (N_846,N_797,N_740);
and U847 (N_847,N_700,N_795);
nor U848 (N_848,N_761,N_798);
or U849 (N_849,N_726,N_757);
and U850 (N_850,N_731,N_734);
nor U851 (N_851,N_790,N_745);
or U852 (N_852,N_752,N_799);
nand U853 (N_853,N_745,N_756);
nand U854 (N_854,N_760,N_762);
nand U855 (N_855,N_747,N_799);
nand U856 (N_856,N_730,N_781);
and U857 (N_857,N_744,N_732);
nor U858 (N_858,N_792,N_752);
or U859 (N_859,N_767,N_715);
nor U860 (N_860,N_727,N_757);
nor U861 (N_861,N_765,N_750);
and U862 (N_862,N_748,N_706);
nor U863 (N_863,N_747,N_786);
nand U864 (N_864,N_705,N_725);
and U865 (N_865,N_769,N_716);
nand U866 (N_866,N_793,N_766);
and U867 (N_867,N_791,N_740);
nand U868 (N_868,N_796,N_750);
and U869 (N_869,N_742,N_735);
and U870 (N_870,N_753,N_796);
nand U871 (N_871,N_797,N_721);
and U872 (N_872,N_745,N_724);
nor U873 (N_873,N_724,N_791);
and U874 (N_874,N_773,N_747);
and U875 (N_875,N_713,N_736);
nand U876 (N_876,N_767,N_765);
or U877 (N_877,N_732,N_772);
and U878 (N_878,N_792,N_700);
nand U879 (N_879,N_754,N_797);
or U880 (N_880,N_710,N_745);
or U881 (N_881,N_734,N_784);
and U882 (N_882,N_721,N_758);
nor U883 (N_883,N_719,N_795);
or U884 (N_884,N_718,N_742);
nor U885 (N_885,N_759,N_750);
and U886 (N_886,N_758,N_756);
nand U887 (N_887,N_786,N_743);
nand U888 (N_888,N_770,N_798);
nand U889 (N_889,N_746,N_769);
and U890 (N_890,N_737,N_704);
and U891 (N_891,N_746,N_703);
nand U892 (N_892,N_794,N_778);
nor U893 (N_893,N_701,N_726);
or U894 (N_894,N_727,N_756);
and U895 (N_895,N_759,N_723);
nor U896 (N_896,N_723,N_797);
nand U897 (N_897,N_707,N_728);
nand U898 (N_898,N_782,N_746);
nor U899 (N_899,N_701,N_705);
nand U900 (N_900,N_831,N_853);
and U901 (N_901,N_882,N_892);
and U902 (N_902,N_893,N_861);
or U903 (N_903,N_802,N_800);
xnor U904 (N_904,N_847,N_801);
or U905 (N_905,N_829,N_874);
or U906 (N_906,N_811,N_870);
nor U907 (N_907,N_835,N_812);
or U908 (N_908,N_838,N_858);
and U909 (N_909,N_865,N_868);
and U910 (N_910,N_808,N_839);
xnor U911 (N_911,N_846,N_851);
and U912 (N_912,N_805,N_821);
and U913 (N_913,N_859,N_825);
nand U914 (N_914,N_849,N_857);
xnor U915 (N_915,N_819,N_872);
and U916 (N_916,N_852,N_817);
xnor U917 (N_917,N_814,N_813);
nor U918 (N_918,N_815,N_824);
and U919 (N_919,N_883,N_866);
nor U920 (N_920,N_889,N_885);
nand U921 (N_921,N_818,N_871);
or U922 (N_922,N_848,N_832);
nand U923 (N_923,N_803,N_879);
nor U924 (N_924,N_887,N_804);
nor U925 (N_925,N_862,N_816);
or U926 (N_926,N_855,N_807);
or U927 (N_927,N_834,N_833);
and U928 (N_928,N_844,N_899);
nand U929 (N_929,N_806,N_888);
and U930 (N_930,N_864,N_854);
nand U931 (N_931,N_809,N_869);
or U932 (N_932,N_827,N_896);
and U933 (N_933,N_897,N_826);
or U934 (N_934,N_845,N_856);
nand U935 (N_935,N_881,N_841);
and U936 (N_936,N_867,N_875);
and U937 (N_937,N_830,N_886);
or U938 (N_938,N_891,N_880);
and U939 (N_939,N_822,N_837);
nand U940 (N_940,N_877,N_842);
or U941 (N_941,N_828,N_850);
and U942 (N_942,N_810,N_876);
nand U943 (N_943,N_840,N_890);
nor U944 (N_944,N_878,N_836);
nand U945 (N_945,N_863,N_843);
or U946 (N_946,N_898,N_873);
and U947 (N_947,N_894,N_895);
nor U948 (N_948,N_823,N_884);
nor U949 (N_949,N_860,N_820);
and U950 (N_950,N_866,N_886);
nand U951 (N_951,N_875,N_889);
nor U952 (N_952,N_883,N_873);
nand U953 (N_953,N_897,N_896);
and U954 (N_954,N_804,N_812);
nand U955 (N_955,N_831,N_846);
and U956 (N_956,N_889,N_856);
nor U957 (N_957,N_811,N_845);
and U958 (N_958,N_831,N_868);
and U959 (N_959,N_881,N_807);
nor U960 (N_960,N_889,N_851);
nand U961 (N_961,N_819,N_888);
or U962 (N_962,N_882,N_833);
nor U963 (N_963,N_843,N_854);
or U964 (N_964,N_895,N_880);
nor U965 (N_965,N_860,N_891);
and U966 (N_966,N_815,N_896);
nor U967 (N_967,N_897,N_886);
and U968 (N_968,N_831,N_807);
xor U969 (N_969,N_840,N_878);
or U970 (N_970,N_852,N_869);
or U971 (N_971,N_802,N_849);
nand U972 (N_972,N_875,N_873);
nor U973 (N_973,N_874,N_838);
nor U974 (N_974,N_841,N_818);
and U975 (N_975,N_881,N_837);
xnor U976 (N_976,N_850,N_843);
and U977 (N_977,N_887,N_878);
and U978 (N_978,N_832,N_831);
nand U979 (N_979,N_850,N_852);
or U980 (N_980,N_879,N_880);
nand U981 (N_981,N_818,N_832);
nand U982 (N_982,N_848,N_840);
or U983 (N_983,N_891,N_844);
or U984 (N_984,N_897,N_840);
and U985 (N_985,N_842,N_828);
nor U986 (N_986,N_887,N_841);
nor U987 (N_987,N_850,N_829);
xnor U988 (N_988,N_876,N_840);
nand U989 (N_989,N_874,N_857);
nor U990 (N_990,N_831,N_841);
nor U991 (N_991,N_854,N_800);
or U992 (N_992,N_833,N_885);
nand U993 (N_993,N_832,N_876);
and U994 (N_994,N_830,N_891);
nand U995 (N_995,N_867,N_883);
nor U996 (N_996,N_877,N_869);
nor U997 (N_997,N_800,N_863);
nor U998 (N_998,N_893,N_806);
or U999 (N_999,N_836,N_885);
or U1000 (N_1000,N_941,N_926);
or U1001 (N_1001,N_977,N_948);
nor U1002 (N_1002,N_994,N_987);
nor U1003 (N_1003,N_903,N_920);
and U1004 (N_1004,N_908,N_947);
xor U1005 (N_1005,N_957,N_969);
or U1006 (N_1006,N_988,N_936);
nand U1007 (N_1007,N_966,N_995);
nor U1008 (N_1008,N_978,N_934);
nand U1009 (N_1009,N_963,N_980);
and U1010 (N_1010,N_958,N_912);
nor U1011 (N_1011,N_921,N_968);
nand U1012 (N_1012,N_946,N_923);
nand U1013 (N_1013,N_982,N_952);
nand U1014 (N_1014,N_949,N_983);
and U1015 (N_1015,N_956,N_916);
nand U1016 (N_1016,N_991,N_902);
or U1017 (N_1017,N_967,N_944);
or U1018 (N_1018,N_935,N_975);
nand U1019 (N_1019,N_917,N_922);
or U1020 (N_1020,N_954,N_915);
xnor U1021 (N_1021,N_986,N_945);
nor U1022 (N_1022,N_998,N_940);
or U1023 (N_1023,N_964,N_990);
xnor U1024 (N_1024,N_913,N_937);
nor U1025 (N_1025,N_971,N_943);
nor U1026 (N_1026,N_992,N_930);
nand U1027 (N_1027,N_996,N_953);
and U1028 (N_1028,N_906,N_972);
nor U1029 (N_1029,N_955,N_939);
nor U1030 (N_1030,N_959,N_927);
nor U1031 (N_1031,N_984,N_919);
nand U1032 (N_1032,N_904,N_909);
nand U1033 (N_1033,N_976,N_970);
nand U1034 (N_1034,N_900,N_938);
and U1035 (N_1035,N_989,N_911);
or U1036 (N_1036,N_961,N_932);
nand U1037 (N_1037,N_910,N_924);
nor U1038 (N_1038,N_985,N_997);
and U1039 (N_1039,N_965,N_999);
or U1040 (N_1040,N_942,N_931);
and U1041 (N_1041,N_914,N_929);
nor U1042 (N_1042,N_918,N_951);
or U1043 (N_1043,N_907,N_973);
xor U1044 (N_1044,N_901,N_981);
and U1045 (N_1045,N_979,N_974);
nor U1046 (N_1046,N_928,N_950);
nand U1047 (N_1047,N_925,N_960);
nor U1048 (N_1048,N_993,N_962);
or U1049 (N_1049,N_905,N_933);
nand U1050 (N_1050,N_956,N_978);
nand U1051 (N_1051,N_925,N_991);
or U1052 (N_1052,N_993,N_988);
and U1053 (N_1053,N_984,N_937);
or U1054 (N_1054,N_909,N_920);
or U1055 (N_1055,N_981,N_999);
or U1056 (N_1056,N_986,N_930);
and U1057 (N_1057,N_929,N_939);
or U1058 (N_1058,N_929,N_903);
and U1059 (N_1059,N_951,N_985);
nor U1060 (N_1060,N_913,N_975);
nor U1061 (N_1061,N_966,N_987);
xnor U1062 (N_1062,N_925,N_965);
nand U1063 (N_1063,N_986,N_908);
nand U1064 (N_1064,N_955,N_997);
nand U1065 (N_1065,N_942,N_995);
nor U1066 (N_1066,N_938,N_930);
nand U1067 (N_1067,N_987,N_997);
or U1068 (N_1068,N_913,N_938);
and U1069 (N_1069,N_993,N_927);
or U1070 (N_1070,N_934,N_972);
nand U1071 (N_1071,N_923,N_981);
nand U1072 (N_1072,N_967,N_901);
and U1073 (N_1073,N_996,N_901);
nor U1074 (N_1074,N_970,N_939);
or U1075 (N_1075,N_933,N_913);
nor U1076 (N_1076,N_932,N_979);
or U1077 (N_1077,N_939,N_935);
nand U1078 (N_1078,N_944,N_902);
nor U1079 (N_1079,N_952,N_929);
nor U1080 (N_1080,N_990,N_900);
nand U1081 (N_1081,N_948,N_970);
nor U1082 (N_1082,N_916,N_928);
and U1083 (N_1083,N_949,N_968);
nand U1084 (N_1084,N_981,N_938);
nor U1085 (N_1085,N_922,N_900);
or U1086 (N_1086,N_921,N_972);
xnor U1087 (N_1087,N_971,N_985);
nand U1088 (N_1088,N_901,N_984);
nand U1089 (N_1089,N_901,N_998);
nand U1090 (N_1090,N_989,N_996);
and U1091 (N_1091,N_997,N_984);
and U1092 (N_1092,N_976,N_979);
and U1093 (N_1093,N_930,N_988);
nand U1094 (N_1094,N_944,N_904);
or U1095 (N_1095,N_933,N_909);
and U1096 (N_1096,N_935,N_992);
nor U1097 (N_1097,N_969,N_915);
nand U1098 (N_1098,N_910,N_990);
nor U1099 (N_1099,N_994,N_970);
or U1100 (N_1100,N_1021,N_1038);
or U1101 (N_1101,N_1042,N_1003);
nor U1102 (N_1102,N_1037,N_1004);
and U1103 (N_1103,N_1055,N_1081);
xnor U1104 (N_1104,N_1091,N_1007);
and U1105 (N_1105,N_1056,N_1093);
nand U1106 (N_1106,N_1010,N_1043);
nor U1107 (N_1107,N_1031,N_1090);
or U1108 (N_1108,N_1029,N_1012);
nor U1109 (N_1109,N_1066,N_1008);
nand U1110 (N_1110,N_1089,N_1016);
nor U1111 (N_1111,N_1033,N_1046);
and U1112 (N_1112,N_1065,N_1079);
and U1113 (N_1113,N_1067,N_1092);
and U1114 (N_1114,N_1086,N_1098);
and U1115 (N_1115,N_1013,N_1022);
nand U1116 (N_1116,N_1099,N_1000);
nand U1117 (N_1117,N_1070,N_1096);
and U1118 (N_1118,N_1063,N_1001);
nor U1119 (N_1119,N_1040,N_1072);
and U1120 (N_1120,N_1014,N_1052);
and U1121 (N_1121,N_1084,N_1064);
and U1122 (N_1122,N_1094,N_1034);
nor U1123 (N_1123,N_1006,N_1026);
or U1124 (N_1124,N_1076,N_1039);
nor U1125 (N_1125,N_1061,N_1071);
or U1126 (N_1126,N_1095,N_1083);
nor U1127 (N_1127,N_1002,N_1009);
nand U1128 (N_1128,N_1053,N_1023);
xnor U1129 (N_1129,N_1097,N_1062);
nand U1130 (N_1130,N_1085,N_1032);
nand U1131 (N_1131,N_1011,N_1051);
or U1132 (N_1132,N_1028,N_1078);
or U1133 (N_1133,N_1088,N_1073);
nor U1134 (N_1134,N_1075,N_1036);
nand U1135 (N_1135,N_1019,N_1044);
and U1136 (N_1136,N_1060,N_1068);
or U1137 (N_1137,N_1030,N_1054);
or U1138 (N_1138,N_1047,N_1058);
nor U1139 (N_1139,N_1015,N_1048);
and U1140 (N_1140,N_1059,N_1027);
or U1141 (N_1141,N_1049,N_1024);
and U1142 (N_1142,N_1035,N_1069);
nand U1143 (N_1143,N_1005,N_1082);
nor U1144 (N_1144,N_1018,N_1050);
nor U1145 (N_1145,N_1080,N_1077);
nor U1146 (N_1146,N_1017,N_1074);
and U1147 (N_1147,N_1057,N_1045);
xor U1148 (N_1148,N_1041,N_1087);
nor U1149 (N_1149,N_1020,N_1025);
nor U1150 (N_1150,N_1092,N_1099);
nor U1151 (N_1151,N_1056,N_1010);
nor U1152 (N_1152,N_1062,N_1032);
nor U1153 (N_1153,N_1064,N_1081);
nor U1154 (N_1154,N_1052,N_1036);
and U1155 (N_1155,N_1077,N_1062);
and U1156 (N_1156,N_1062,N_1038);
or U1157 (N_1157,N_1098,N_1038);
nand U1158 (N_1158,N_1081,N_1038);
nand U1159 (N_1159,N_1037,N_1035);
nor U1160 (N_1160,N_1022,N_1019);
and U1161 (N_1161,N_1089,N_1008);
nor U1162 (N_1162,N_1012,N_1070);
nand U1163 (N_1163,N_1008,N_1096);
nand U1164 (N_1164,N_1008,N_1030);
or U1165 (N_1165,N_1098,N_1075);
and U1166 (N_1166,N_1075,N_1050);
and U1167 (N_1167,N_1062,N_1024);
nand U1168 (N_1168,N_1075,N_1041);
nand U1169 (N_1169,N_1025,N_1029);
nand U1170 (N_1170,N_1013,N_1050);
or U1171 (N_1171,N_1024,N_1021);
nor U1172 (N_1172,N_1051,N_1041);
nand U1173 (N_1173,N_1000,N_1013);
nor U1174 (N_1174,N_1070,N_1073);
or U1175 (N_1175,N_1028,N_1086);
or U1176 (N_1176,N_1053,N_1052);
or U1177 (N_1177,N_1088,N_1043);
and U1178 (N_1178,N_1099,N_1098);
nand U1179 (N_1179,N_1099,N_1081);
nand U1180 (N_1180,N_1069,N_1075);
and U1181 (N_1181,N_1003,N_1075);
or U1182 (N_1182,N_1073,N_1052);
nor U1183 (N_1183,N_1043,N_1056);
and U1184 (N_1184,N_1041,N_1030);
or U1185 (N_1185,N_1089,N_1096);
nand U1186 (N_1186,N_1019,N_1067);
nand U1187 (N_1187,N_1004,N_1032);
and U1188 (N_1188,N_1068,N_1029);
and U1189 (N_1189,N_1088,N_1096);
and U1190 (N_1190,N_1000,N_1017);
nand U1191 (N_1191,N_1019,N_1073);
and U1192 (N_1192,N_1042,N_1094);
and U1193 (N_1193,N_1013,N_1016);
and U1194 (N_1194,N_1011,N_1020);
or U1195 (N_1195,N_1012,N_1051);
and U1196 (N_1196,N_1025,N_1059);
or U1197 (N_1197,N_1010,N_1086);
nor U1198 (N_1198,N_1084,N_1053);
and U1199 (N_1199,N_1006,N_1070);
and U1200 (N_1200,N_1149,N_1125);
nand U1201 (N_1201,N_1169,N_1198);
nand U1202 (N_1202,N_1145,N_1153);
or U1203 (N_1203,N_1148,N_1136);
and U1204 (N_1204,N_1124,N_1191);
nor U1205 (N_1205,N_1105,N_1138);
and U1206 (N_1206,N_1199,N_1134);
or U1207 (N_1207,N_1143,N_1185);
nor U1208 (N_1208,N_1119,N_1158);
or U1209 (N_1209,N_1151,N_1128);
nor U1210 (N_1210,N_1144,N_1171);
xnor U1211 (N_1211,N_1176,N_1131);
nand U1212 (N_1212,N_1140,N_1123);
or U1213 (N_1213,N_1186,N_1107);
nor U1214 (N_1214,N_1192,N_1101);
nand U1215 (N_1215,N_1184,N_1103);
and U1216 (N_1216,N_1142,N_1115);
or U1217 (N_1217,N_1165,N_1155);
and U1218 (N_1218,N_1137,N_1196);
nor U1219 (N_1219,N_1100,N_1168);
or U1220 (N_1220,N_1116,N_1161);
and U1221 (N_1221,N_1154,N_1152);
nor U1222 (N_1222,N_1189,N_1164);
nor U1223 (N_1223,N_1114,N_1178);
or U1224 (N_1224,N_1156,N_1129);
nand U1225 (N_1225,N_1112,N_1159);
nand U1226 (N_1226,N_1170,N_1130);
nand U1227 (N_1227,N_1118,N_1150);
nand U1228 (N_1228,N_1126,N_1174);
nand U1229 (N_1229,N_1108,N_1187);
and U1230 (N_1230,N_1146,N_1180);
nand U1231 (N_1231,N_1188,N_1117);
or U1232 (N_1232,N_1121,N_1181);
and U1233 (N_1233,N_1147,N_1177);
nor U1234 (N_1234,N_1175,N_1193);
or U1235 (N_1235,N_1141,N_1157);
nor U1236 (N_1236,N_1194,N_1106);
nand U1237 (N_1237,N_1172,N_1163);
nand U1238 (N_1238,N_1197,N_1104);
or U1239 (N_1239,N_1162,N_1102);
xor U1240 (N_1240,N_1179,N_1111);
or U1241 (N_1241,N_1135,N_1109);
and U1242 (N_1242,N_1190,N_1167);
and U1243 (N_1243,N_1160,N_1120);
nor U1244 (N_1244,N_1113,N_1110);
or U1245 (N_1245,N_1139,N_1127);
and U1246 (N_1246,N_1166,N_1173);
or U1247 (N_1247,N_1133,N_1183);
nand U1248 (N_1248,N_1182,N_1195);
nand U1249 (N_1249,N_1132,N_1122);
nand U1250 (N_1250,N_1126,N_1196);
nor U1251 (N_1251,N_1157,N_1116);
and U1252 (N_1252,N_1158,N_1173);
or U1253 (N_1253,N_1164,N_1182);
or U1254 (N_1254,N_1133,N_1147);
and U1255 (N_1255,N_1198,N_1171);
nor U1256 (N_1256,N_1189,N_1185);
nand U1257 (N_1257,N_1179,N_1102);
or U1258 (N_1258,N_1167,N_1135);
nor U1259 (N_1259,N_1154,N_1125);
nor U1260 (N_1260,N_1168,N_1186);
and U1261 (N_1261,N_1151,N_1179);
nand U1262 (N_1262,N_1100,N_1159);
nor U1263 (N_1263,N_1192,N_1155);
and U1264 (N_1264,N_1133,N_1136);
and U1265 (N_1265,N_1121,N_1120);
or U1266 (N_1266,N_1170,N_1165);
and U1267 (N_1267,N_1102,N_1134);
xor U1268 (N_1268,N_1155,N_1177);
and U1269 (N_1269,N_1192,N_1196);
and U1270 (N_1270,N_1186,N_1129);
nand U1271 (N_1271,N_1123,N_1176);
or U1272 (N_1272,N_1173,N_1186);
or U1273 (N_1273,N_1188,N_1149);
nor U1274 (N_1274,N_1189,N_1152);
nor U1275 (N_1275,N_1140,N_1186);
and U1276 (N_1276,N_1131,N_1134);
and U1277 (N_1277,N_1146,N_1159);
nor U1278 (N_1278,N_1152,N_1119);
and U1279 (N_1279,N_1196,N_1101);
nand U1280 (N_1280,N_1141,N_1127);
or U1281 (N_1281,N_1183,N_1108);
nor U1282 (N_1282,N_1192,N_1179);
nand U1283 (N_1283,N_1151,N_1149);
or U1284 (N_1284,N_1152,N_1131);
nor U1285 (N_1285,N_1190,N_1197);
and U1286 (N_1286,N_1109,N_1174);
or U1287 (N_1287,N_1131,N_1137);
nand U1288 (N_1288,N_1172,N_1102);
and U1289 (N_1289,N_1111,N_1187);
or U1290 (N_1290,N_1110,N_1169);
or U1291 (N_1291,N_1124,N_1165);
and U1292 (N_1292,N_1172,N_1189);
nor U1293 (N_1293,N_1127,N_1142);
nor U1294 (N_1294,N_1180,N_1172);
or U1295 (N_1295,N_1126,N_1198);
and U1296 (N_1296,N_1189,N_1174);
nand U1297 (N_1297,N_1105,N_1149);
nand U1298 (N_1298,N_1172,N_1128);
and U1299 (N_1299,N_1101,N_1120);
or U1300 (N_1300,N_1239,N_1208);
and U1301 (N_1301,N_1221,N_1274);
nor U1302 (N_1302,N_1280,N_1237);
and U1303 (N_1303,N_1253,N_1298);
and U1304 (N_1304,N_1278,N_1273);
nand U1305 (N_1305,N_1236,N_1248);
nand U1306 (N_1306,N_1276,N_1207);
xor U1307 (N_1307,N_1257,N_1211);
nor U1308 (N_1308,N_1234,N_1202);
nand U1309 (N_1309,N_1260,N_1287);
nand U1310 (N_1310,N_1220,N_1281);
and U1311 (N_1311,N_1264,N_1204);
and U1312 (N_1312,N_1256,N_1200);
nor U1313 (N_1313,N_1284,N_1296);
and U1314 (N_1314,N_1210,N_1255);
nor U1315 (N_1315,N_1251,N_1222);
and U1316 (N_1316,N_1246,N_1252);
nor U1317 (N_1317,N_1244,N_1288);
xnor U1318 (N_1318,N_1268,N_1279);
xor U1319 (N_1319,N_1240,N_1265);
nand U1320 (N_1320,N_1242,N_1263);
or U1321 (N_1321,N_1247,N_1277);
nand U1322 (N_1322,N_1282,N_1230);
nor U1323 (N_1323,N_1275,N_1217);
nand U1324 (N_1324,N_1233,N_1269);
nor U1325 (N_1325,N_1201,N_1286);
nand U1326 (N_1326,N_1231,N_1245);
or U1327 (N_1327,N_1215,N_1243);
or U1328 (N_1328,N_1250,N_1214);
and U1329 (N_1329,N_1227,N_1267);
or U1330 (N_1330,N_1293,N_1238);
and U1331 (N_1331,N_1232,N_1218);
nor U1332 (N_1332,N_1297,N_1292);
or U1333 (N_1333,N_1225,N_1272);
nand U1334 (N_1334,N_1209,N_1219);
nor U1335 (N_1335,N_1270,N_1212);
or U1336 (N_1336,N_1203,N_1259);
or U1337 (N_1337,N_1205,N_1291);
nand U1338 (N_1338,N_1226,N_1285);
nand U1339 (N_1339,N_1266,N_1283);
nand U1340 (N_1340,N_1206,N_1229);
or U1341 (N_1341,N_1262,N_1290);
nor U1342 (N_1342,N_1241,N_1223);
nand U1343 (N_1343,N_1228,N_1294);
or U1344 (N_1344,N_1216,N_1224);
and U1345 (N_1345,N_1213,N_1258);
or U1346 (N_1346,N_1299,N_1289);
nor U1347 (N_1347,N_1235,N_1295);
nand U1348 (N_1348,N_1271,N_1249);
nand U1349 (N_1349,N_1261,N_1254);
or U1350 (N_1350,N_1230,N_1226);
xor U1351 (N_1351,N_1254,N_1204);
or U1352 (N_1352,N_1209,N_1218);
or U1353 (N_1353,N_1227,N_1217);
nor U1354 (N_1354,N_1289,N_1248);
nand U1355 (N_1355,N_1242,N_1285);
or U1356 (N_1356,N_1267,N_1287);
nand U1357 (N_1357,N_1228,N_1283);
nor U1358 (N_1358,N_1280,N_1250);
or U1359 (N_1359,N_1241,N_1277);
nor U1360 (N_1360,N_1245,N_1238);
nand U1361 (N_1361,N_1262,N_1230);
or U1362 (N_1362,N_1220,N_1225);
nand U1363 (N_1363,N_1207,N_1201);
nor U1364 (N_1364,N_1225,N_1242);
or U1365 (N_1365,N_1290,N_1263);
nor U1366 (N_1366,N_1202,N_1258);
and U1367 (N_1367,N_1248,N_1218);
and U1368 (N_1368,N_1208,N_1231);
or U1369 (N_1369,N_1234,N_1286);
or U1370 (N_1370,N_1291,N_1203);
and U1371 (N_1371,N_1252,N_1269);
or U1372 (N_1372,N_1283,N_1246);
nand U1373 (N_1373,N_1229,N_1261);
nor U1374 (N_1374,N_1219,N_1248);
and U1375 (N_1375,N_1219,N_1225);
and U1376 (N_1376,N_1221,N_1204);
nor U1377 (N_1377,N_1282,N_1220);
nand U1378 (N_1378,N_1213,N_1201);
nor U1379 (N_1379,N_1225,N_1237);
or U1380 (N_1380,N_1265,N_1266);
xnor U1381 (N_1381,N_1235,N_1245);
and U1382 (N_1382,N_1201,N_1218);
nor U1383 (N_1383,N_1253,N_1232);
and U1384 (N_1384,N_1221,N_1252);
and U1385 (N_1385,N_1284,N_1299);
nor U1386 (N_1386,N_1210,N_1251);
or U1387 (N_1387,N_1273,N_1223);
or U1388 (N_1388,N_1215,N_1228);
nand U1389 (N_1389,N_1270,N_1207);
nand U1390 (N_1390,N_1250,N_1230);
nand U1391 (N_1391,N_1250,N_1267);
and U1392 (N_1392,N_1261,N_1204);
or U1393 (N_1393,N_1289,N_1263);
nand U1394 (N_1394,N_1228,N_1238);
nand U1395 (N_1395,N_1206,N_1256);
or U1396 (N_1396,N_1280,N_1228);
or U1397 (N_1397,N_1222,N_1276);
and U1398 (N_1398,N_1200,N_1278);
nor U1399 (N_1399,N_1259,N_1260);
and U1400 (N_1400,N_1332,N_1384);
nand U1401 (N_1401,N_1395,N_1387);
or U1402 (N_1402,N_1367,N_1301);
nand U1403 (N_1403,N_1399,N_1361);
or U1404 (N_1404,N_1371,N_1325);
or U1405 (N_1405,N_1333,N_1372);
xnor U1406 (N_1406,N_1391,N_1343);
xnor U1407 (N_1407,N_1313,N_1357);
nor U1408 (N_1408,N_1340,N_1394);
nor U1409 (N_1409,N_1349,N_1386);
nand U1410 (N_1410,N_1393,N_1323);
nand U1411 (N_1411,N_1388,N_1354);
nor U1412 (N_1412,N_1348,N_1305);
nand U1413 (N_1413,N_1366,N_1315);
or U1414 (N_1414,N_1383,N_1328);
or U1415 (N_1415,N_1304,N_1363);
nor U1416 (N_1416,N_1318,N_1329);
xnor U1417 (N_1417,N_1317,N_1389);
or U1418 (N_1418,N_1345,N_1375);
or U1419 (N_1419,N_1339,N_1369);
nor U1420 (N_1420,N_1338,N_1309);
nor U1421 (N_1421,N_1310,N_1355);
nand U1422 (N_1422,N_1351,N_1359);
and U1423 (N_1423,N_1335,N_1336);
nand U1424 (N_1424,N_1327,N_1358);
nor U1425 (N_1425,N_1352,N_1306);
and U1426 (N_1426,N_1373,N_1365);
nor U1427 (N_1427,N_1346,N_1324);
nand U1428 (N_1428,N_1307,N_1385);
and U1429 (N_1429,N_1312,N_1379);
nor U1430 (N_1430,N_1350,N_1370);
or U1431 (N_1431,N_1374,N_1381);
or U1432 (N_1432,N_1356,N_1337);
nor U1433 (N_1433,N_1378,N_1334);
nand U1434 (N_1434,N_1321,N_1311);
nor U1435 (N_1435,N_1347,N_1302);
nand U1436 (N_1436,N_1303,N_1326);
nand U1437 (N_1437,N_1397,N_1368);
nor U1438 (N_1438,N_1396,N_1353);
nand U1439 (N_1439,N_1360,N_1390);
and U1440 (N_1440,N_1320,N_1308);
or U1441 (N_1441,N_1314,N_1319);
or U1442 (N_1442,N_1377,N_1344);
and U1443 (N_1443,N_1392,N_1300);
nand U1444 (N_1444,N_1380,N_1362);
and U1445 (N_1445,N_1322,N_1331);
nand U1446 (N_1446,N_1382,N_1398);
or U1447 (N_1447,N_1330,N_1342);
nor U1448 (N_1448,N_1364,N_1341);
nor U1449 (N_1449,N_1376,N_1316);
xor U1450 (N_1450,N_1332,N_1326);
or U1451 (N_1451,N_1327,N_1343);
or U1452 (N_1452,N_1395,N_1339);
nand U1453 (N_1453,N_1311,N_1326);
xnor U1454 (N_1454,N_1350,N_1399);
nand U1455 (N_1455,N_1313,N_1380);
nand U1456 (N_1456,N_1310,N_1337);
and U1457 (N_1457,N_1379,N_1351);
or U1458 (N_1458,N_1300,N_1315);
nor U1459 (N_1459,N_1356,N_1385);
and U1460 (N_1460,N_1360,N_1363);
nand U1461 (N_1461,N_1353,N_1354);
nand U1462 (N_1462,N_1396,N_1339);
nor U1463 (N_1463,N_1317,N_1328);
and U1464 (N_1464,N_1305,N_1351);
or U1465 (N_1465,N_1385,N_1300);
and U1466 (N_1466,N_1342,N_1329);
or U1467 (N_1467,N_1391,N_1368);
nand U1468 (N_1468,N_1322,N_1305);
or U1469 (N_1469,N_1336,N_1348);
or U1470 (N_1470,N_1351,N_1326);
or U1471 (N_1471,N_1308,N_1388);
or U1472 (N_1472,N_1367,N_1399);
and U1473 (N_1473,N_1318,N_1312);
nand U1474 (N_1474,N_1310,N_1349);
or U1475 (N_1475,N_1395,N_1318);
and U1476 (N_1476,N_1347,N_1318);
and U1477 (N_1477,N_1359,N_1337);
and U1478 (N_1478,N_1355,N_1399);
or U1479 (N_1479,N_1383,N_1325);
and U1480 (N_1480,N_1379,N_1311);
and U1481 (N_1481,N_1360,N_1336);
nand U1482 (N_1482,N_1325,N_1381);
and U1483 (N_1483,N_1335,N_1300);
nand U1484 (N_1484,N_1316,N_1346);
nand U1485 (N_1485,N_1351,N_1314);
nand U1486 (N_1486,N_1352,N_1345);
and U1487 (N_1487,N_1359,N_1383);
or U1488 (N_1488,N_1308,N_1391);
or U1489 (N_1489,N_1389,N_1355);
nor U1490 (N_1490,N_1300,N_1332);
or U1491 (N_1491,N_1357,N_1374);
xnor U1492 (N_1492,N_1310,N_1320);
nor U1493 (N_1493,N_1339,N_1343);
nor U1494 (N_1494,N_1318,N_1389);
or U1495 (N_1495,N_1365,N_1364);
nor U1496 (N_1496,N_1341,N_1383);
and U1497 (N_1497,N_1353,N_1333);
and U1498 (N_1498,N_1383,N_1377);
nand U1499 (N_1499,N_1360,N_1394);
or U1500 (N_1500,N_1404,N_1458);
xnor U1501 (N_1501,N_1405,N_1447);
nor U1502 (N_1502,N_1498,N_1409);
or U1503 (N_1503,N_1417,N_1430);
nand U1504 (N_1504,N_1472,N_1418);
or U1505 (N_1505,N_1401,N_1461);
and U1506 (N_1506,N_1457,N_1481);
and U1507 (N_1507,N_1471,N_1492);
nor U1508 (N_1508,N_1411,N_1440);
and U1509 (N_1509,N_1469,N_1466);
nand U1510 (N_1510,N_1412,N_1455);
nand U1511 (N_1511,N_1470,N_1419);
or U1512 (N_1512,N_1420,N_1479);
xor U1513 (N_1513,N_1446,N_1442);
or U1514 (N_1514,N_1487,N_1454);
xnor U1515 (N_1515,N_1443,N_1437);
nand U1516 (N_1516,N_1475,N_1436);
or U1517 (N_1517,N_1478,N_1493);
and U1518 (N_1518,N_1425,N_1482);
nand U1519 (N_1519,N_1459,N_1410);
and U1520 (N_1520,N_1415,N_1460);
nand U1521 (N_1521,N_1464,N_1465);
nor U1522 (N_1522,N_1413,N_1400);
nor U1523 (N_1523,N_1426,N_1473);
nand U1524 (N_1524,N_1421,N_1422);
and U1525 (N_1525,N_1445,N_1407);
xor U1526 (N_1526,N_1483,N_1485);
or U1527 (N_1527,N_1449,N_1428);
nand U1528 (N_1528,N_1423,N_1435);
nand U1529 (N_1529,N_1477,N_1489);
or U1530 (N_1530,N_1448,N_1462);
and U1531 (N_1531,N_1496,N_1402);
or U1532 (N_1532,N_1441,N_1414);
nor U1533 (N_1533,N_1408,N_1488);
nand U1534 (N_1534,N_1494,N_1429);
nand U1535 (N_1535,N_1403,N_1453);
nor U1536 (N_1536,N_1468,N_1439);
and U1537 (N_1537,N_1452,N_1480);
nor U1538 (N_1538,N_1427,N_1431);
or U1539 (N_1539,N_1438,N_1424);
nand U1540 (N_1540,N_1490,N_1406);
and U1541 (N_1541,N_1495,N_1467);
nand U1542 (N_1542,N_1433,N_1484);
nand U1543 (N_1543,N_1474,N_1486);
nand U1544 (N_1544,N_1476,N_1491);
and U1545 (N_1545,N_1456,N_1450);
nor U1546 (N_1546,N_1432,N_1416);
and U1547 (N_1547,N_1444,N_1499);
and U1548 (N_1548,N_1463,N_1434);
nand U1549 (N_1549,N_1497,N_1451);
and U1550 (N_1550,N_1418,N_1444);
or U1551 (N_1551,N_1485,N_1455);
or U1552 (N_1552,N_1464,N_1482);
nand U1553 (N_1553,N_1442,N_1410);
or U1554 (N_1554,N_1457,N_1490);
nand U1555 (N_1555,N_1494,N_1436);
and U1556 (N_1556,N_1461,N_1498);
nor U1557 (N_1557,N_1457,N_1436);
nor U1558 (N_1558,N_1455,N_1466);
nor U1559 (N_1559,N_1475,N_1490);
and U1560 (N_1560,N_1463,N_1406);
nor U1561 (N_1561,N_1493,N_1495);
and U1562 (N_1562,N_1472,N_1486);
or U1563 (N_1563,N_1465,N_1412);
nor U1564 (N_1564,N_1455,N_1471);
nand U1565 (N_1565,N_1428,N_1479);
nor U1566 (N_1566,N_1440,N_1486);
nand U1567 (N_1567,N_1469,N_1435);
nand U1568 (N_1568,N_1438,N_1487);
nand U1569 (N_1569,N_1492,N_1434);
and U1570 (N_1570,N_1434,N_1437);
or U1571 (N_1571,N_1479,N_1493);
and U1572 (N_1572,N_1410,N_1439);
nor U1573 (N_1573,N_1469,N_1437);
nand U1574 (N_1574,N_1450,N_1409);
nand U1575 (N_1575,N_1458,N_1439);
nor U1576 (N_1576,N_1488,N_1495);
nor U1577 (N_1577,N_1465,N_1468);
and U1578 (N_1578,N_1410,N_1402);
nand U1579 (N_1579,N_1428,N_1460);
or U1580 (N_1580,N_1410,N_1423);
or U1581 (N_1581,N_1469,N_1414);
nand U1582 (N_1582,N_1442,N_1491);
nand U1583 (N_1583,N_1449,N_1480);
or U1584 (N_1584,N_1484,N_1458);
nor U1585 (N_1585,N_1433,N_1405);
or U1586 (N_1586,N_1473,N_1446);
or U1587 (N_1587,N_1429,N_1434);
nand U1588 (N_1588,N_1435,N_1498);
nor U1589 (N_1589,N_1411,N_1431);
nor U1590 (N_1590,N_1492,N_1482);
or U1591 (N_1591,N_1493,N_1436);
nor U1592 (N_1592,N_1438,N_1493);
nor U1593 (N_1593,N_1451,N_1438);
xor U1594 (N_1594,N_1440,N_1443);
and U1595 (N_1595,N_1440,N_1445);
and U1596 (N_1596,N_1433,N_1456);
nand U1597 (N_1597,N_1462,N_1488);
and U1598 (N_1598,N_1438,N_1457);
or U1599 (N_1599,N_1485,N_1442);
nor U1600 (N_1600,N_1543,N_1540);
or U1601 (N_1601,N_1587,N_1511);
or U1602 (N_1602,N_1509,N_1575);
nor U1603 (N_1603,N_1542,N_1533);
or U1604 (N_1604,N_1565,N_1539);
nor U1605 (N_1605,N_1514,N_1558);
nand U1606 (N_1606,N_1552,N_1522);
nor U1607 (N_1607,N_1526,N_1554);
xnor U1608 (N_1608,N_1561,N_1524);
or U1609 (N_1609,N_1596,N_1536);
or U1610 (N_1610,N_1571,N_1574);
or U1611 (N_1611,N_1590,N_1503);
and U1612 (N_1612,N_1557,N_1553);
nand U1613 (N_1613,N_1528,N_1599);
nand U1614 (N_1614,N_1568,N_1521);
and U1615 (N_1615,N_1585,N_1500);
or U1616 (N_1616,N_1573,N_1597);
or U1617 (N_1617,N_1507,N_1576);
and U1618 (N_1618,N_1537,N_1506);
or U1619 (N_1619,N_1530,N_1551);
xnor U1620 (N_1620,N_1563,N_1549);
and U1621 (N_1621,N_1560,N_1529);
nor U1622 (N_1622,N_1535,N_1508);
nand U1623 (N_1623,N_1584,N_1593);
nor U1624 (N_1624,N_1566,N_1505);
or U1625 (N_1625,N_1502,N_1520);
or U1626 (N_1626,N_1517,N_1541);
or U1627 (N_1627,N_1501,N_1579);
nand U1628 (N_1628,N_1586,N_1578);
and U1629 (N_1629,N_1547,N_1531);
nor U1630 (N_1630,N_1512,N_1550);
xor U1631 (N_1631,N_1504,N_1555);
or U1632 (N_1632,N_1570,N_1591);
and U1633 (N_1633,N_1594,N_1545);
nor U1634 (N_1634,N_1523,N_1519);
or U1635 (N_1635,N_1562,N_1583);
or U1636 (N_1636,N_1513,N_1595);
or U1637 (N_1637,N_1580,N_1559);
or U1638 (N_1638,N_1569,N_1534);
nor U1639 (N_1639,N_1598,N_1572);
nor U1640 (N_1640,N_1518,N_1556);
nor U1641 (N_1641,N_1527,N_1510);
or U1642 (N_1642,N_1581,N_1525);
and U1643 (N_1643,N_1589,N_1567);
or U1644 (N_1644,N_1546,N_1592);
nor U1645 (N_1645,N_1516,N_1538);
or U1646 (N_1646,N_1588,N_1582);
or U1647 (N_1647,N_1548,N_1564);
nor U1648 (N_1648,N_1544,N_1577);
nand U1649 (N_1649,N_1515,N_1532);
nor U1650 (N_1650,N_1554,N_1518);
or U1651 (N_1651,N_1599,N_1519);
and U1652 (N_1652,N_1545,N_1502);
nor U1653 (N_1653,N_1503,N_1520);
nor U1654 (N_1654,N_1551,N_1565);
or U1655 (N_1655,N_1539,N_1509);
nand U1656 (N_1656,N_1557,N_1519);
nand U1657 (N_1657,N_1516,N_1542);
and U1658 (N_1658,N_1598,N_1563);
and U1659 (N_1659,N_1546,N_1575);
or U1660 (N_1660,N_1582,N_1581);
nor U1661 (N_1661,N_1577,N_1588);
nand U1662 (N_1662,N_1587,N_1528);
nor U1663 (N_1663,N_1527,N_1565);
or U1664 (N_1664,N_1515,N_1582);
nand U1665 (N_1665,N_1502,N_1556);
nand U1666 (N_1666,N_1581,N_1598);
and U1667 (N_1667,N_1533,N_1537);
nor U1668 (N_1668,N_1556,N_1581);
or U1669 (N_1669,N_1584,N_1515);
nor U1670 (N_1670,N_1570,N_1524);
and U1671 (N_1671,N_1506,N_1563);
nor U1672 (N_1672,N_1520,N_1523);
xor U1673 (N_1673,N_1510,N_1580);
and U1674 (N_1674,N_1547,N_1535);
or U1675 (N_1675,N_1523,N_1535);
nor U1676 (N_1676,N_1531,N_1523);
nand U1677 (N_1677,N_1528,N_1593);
nand U1678 (N_1678,N_1599,N_1512);
nand U1679 (N_1679,N_1584,N_1571);
or U1680 (N_1680,N_1539,N_1598);
nand U1681 (N_1681,N_1508,N_1566);
or U1682 (N_1682,N_1514,N_1511);
and U1683 (N_1683,N_1520,N_1553);
and U1684 (N_1684,N_1509,N_1527);
nand U1685 (N_1685,N_1502,N_1592);
and U1686 (N_1686,N_1538,N_1518);
nor U1687 (N_1687,N_1587,N_1546);
nand U1688 (N_1688,N_1597,N_1540);
or U1689 (N_1689,N_1534,N_1563);
nor U1690 (N_1690,N_1518,N_1576);
or U1691 (N_1691,N_1586,N_1592);
nand U1692 (N_1692,N_1569,N_1589);
nand U1693 (N_1693,N_1546,N_1571);
or U1694 (N_1694,N_1548,N_1572);
nor U1695 (N_1695,N_1537,N_1536);
or U1696 (N_1696,N_1570,N_1571);
or U1697 (N_1697,N_1590,N_1518);
or U1698 (N_1698,N_1513,N_1575);
or U1699 (N_1699,N_1544,N_1533);
nand U1700 (N_1700,N_1698,N_1682);
nand U1701 (N_1701,N_1612,N_1655);
and U1702 (N_1702,N_1684,N_1661);
or U1703 (N_1703,N_1624,N_1689);
nand U1704 (N_1704,N_1672,N_1690);
and U1705 (N_1705,N_1618,N_1608);
nor U1706 (N_1706,N_1605,N_1683);
nor U1707 (N_1707,N_1636,N_1637);
and U1708 (N_1708,N_1604,N_1693);
or U1709 (N_1709,N_1610,N_1635);
and U1710 (N_1710,N_1658,N_1695);
nor U1711 (N_1711,N_1613,N_1674);
and U1712 (N_1712,N_1609,N_1606);
nand U1713 (N_1713,N_1673,N_1660);
and U1714 (N_1714,N_1686,N_1666);
and U1715 (N_1715,N_1639,N_1669);
nand U1716 (N_1716,N_1650,N_1601);
or U1717 (N_1717,N_1617,N_1688);
or U1718 (N_1718,N_1694,N_1671);
and U1719 (N_1719,N_1629,N_1691);
or U1720 (N_1720,N_1657,N_1631);
nor U1721 (N_1721,N_1651,N_1692);
or U1722 (N_1722,N_1662,N_1600);
nor U1723 (N_1723,N_1640,N_1643);
and U1724 (N_1724,N_1628,N_1630);
nand U1725 (N_1725,N_1675,N_1696);
and U1726 (N_1726,N_1614,N_1648);
or U1727 (N_1727,N_1653,N_1645);
or U1728 (N_1728,N_1665,N_1647);
nand U1729 (N_1729,N_1616,N_1644);
or U1730 (N_1730,N_1641,N_1676);
nand U1731 (N_1731,N_1681,N_1620);
and U1732 (N_1732,N_1634,N_1633);
and U1733 (N_1733,N_1611,N_1642);
nand U1734 (N_1734,N_1621,N_1656);
and U1735 (N_1735,N_1670,N_1615);
nor U1736 (N_1736,N_1664,N_1627);
or U1737 (N_1737,N_1638,N_1649);
nand U1738 (N_1738,N_1646,N_1699);
and U1739 (N_1739,N_1632,N_1679);
nor U1740 (N_1740,N_1603,N_1622);
xor U1741 (N_1741,N_1685,N_1678);
or U1742 (N_1742,N_1663,N_1602);
and U1743 (N_1743,N_1626,N_1623);
nor U1744 (N_1744,N_1659,N_1668);
nand U1745 (N_1745,N_1619,N_1667);
nor U1746 (N_1746,N_1687,N_1677);
and U1747 (N_1747,N_1607,N_1697);
xnor U1748 (N_1748,N_1680,N_1652);
and U1749 (N_1749,N_1654,N_1625);
or U1750 (N_1750,N_1686,N_1672);
and U1751 (N_1751,N_1660,N_1608);
and U1752 (N_1752,N_1658,N_1634);
and U1753 (N_1753,N_1633,N_1665);
nor U1754 (N_1754,N_1629,N_1666);
and U1755 (N_1755,N_1690,N_1636);
xor U1756 (N_1756,N_1601,N_1685);
and U1757 (N_1757,N_1696,N_1644);
nor U1758 (N_1758,N_1674,N_1658);
nor U1759 (N_1759,N_1651,N_1610);
nand U1760 (N_1760,N_1686,N_1649);
nor U1761 (N_1761,N_1608,N_1641);
nand U1762 (N_1762,N_1678,N_1652);
nor U1763 (N_1763,N_1642,N_1682);
and U1764 (N_1764,N_1638,N_1661);
nor U1765 (N_1765,N_1641,N_1681);
or U1766 (N_1766,N_1670,N_1640);
and U1767 (N_1767,N_1688,N_1662);
and U1768 (N_1768,N_1664,N_1640);
or U1769 (N_1769,N_1600,N_1620);
nand U1770 (N_1770,N_1662,N_1642);
nor U1771 (N_1771,N_1650,N_1607);
xnor U1772 (N_1772,N_1610,N_1601);
nand U1773 (N_1773,N_1667,N_1696);
nor U1774 (N_1774,N_1659,N_1666);
nand U1775 (N_1775,N_1675,N_1694);
and U1776 (N_1776,N_1673,N_1602);
and U1777 (N_1777,N_1686,N_1635);
xnor U1778 (N_1778,N_1673,N_1654);
nor U1779 (N_1779,N_1601,N_1636);
and U1780 (N_1780,N_1697,N_1635);
and U1781 (N_1781,N_1681,N_1642);
nor U1782 (N_1782,N_1693,N_1606);
nand U1783 (N_1783,N_1606,N_1611);
nand U1784 (N_1784,N_1615,N_1645);
nand U1785 (N_1785,N_1619,N_1644);
or U1786 (N_1786,N_1606,N_1648);
or U1787 (N_1787,N_1642,N_1617);
nand U1788 (N_1788,N_1626,N_1638);
nor U1789 (N_1789,N_1668,N_1673);
nand U1790 (N_1790,N_1602,N_1670);
and U1791 (N_1791,N_1654,N_1641);
or U1792 (N_1792,N_1698,N_1695);
and U1793 (N_1793,N_1635,N_1682);
nand U1794 (N_1794,N_1654,N_1680);
and U1795 (N_1795,N_1637,N_1632);
and U1796 (N_1796,N_1654,N_1605);
or U1797 (N_1797,N_1657,N_1607);
and U1798 (N_1798,N_1699,N_1620);
nor U1799 (N_1799,N_1638,N_1633);
or U1800 (N_1800,N_1776,N_1747);
or U1801 (N_1801,N_1721,N_1781);
and U1802 (N_1802,N_1768,N_1741);
and U1803 (N_1803,N_1765,N_1739);
nor U1804 (N_1804,N_1718,N_1715);
or U1805 (N_1805,N_1756,N_1750);
and U1806 (N_1806,N_1792,N_1732);
nor U1807 (N_1807,N_1790,N_1773);
nor U1808 (N_1808,N_1772,N_1733);
nand U1809 (N_1809,N_1797,N_1703);
nand U1810 (N_1810,N_1714,N_1738);
nor U1811 (N_1811,N_1746,N_1785);
or U1812 (N_1812,N_1763,N_1745);
or U1813 (N_1813,N_1710,N_1751);
or U1814 (N_1814,N_1755,N_1722);
or U1815 (N_1815,N_1724,N_1701);
nor U1816 (N_1816,N_1786,N_1717);
and U1817 (N_1817,N_1766,N_1783);
nor U1818 (N_1818,N_1713,N_1711);
nor U1819 (N_1819,N_1725,N_1704);
nor U1820 (N_1820,N_1770,N_1708);
and U1821 (N_1821,N_1700,N_1705);
nor U1822 (N_1822,N_1779,N_1706);
nor U1823 (N_1823,N_1742,N_1769);
nand U1824 (N_1824,N_1794,N_1749);
nor U1825 (N_1825,N_1743,N_1729);
nor U1826 (N_1826,N_1753,N_1799);
or U1827 (N_1827,N_1788,N_1736);
or U1828 (N_1828,N_1760,N_1734);
nor U1829 (N_1829,N_1719,N_1754);
and U1830 (N_1830,N_1709,N_1767);
nand U1831 (N_1831,N_1791,N_1748);
and U1832 (N_1832,N_1730,N_1716);
and U1833 (N_1833,N_1771,N_1731);
nor U1834 (N_1834,N_1702,N_1744);
nor U1835 (N_1835,N_1778,N_1759);
nor U1836 (N_1836,N_1796,N_1780);
or U1837 (N_1837,N_1735,N_1723);
and U1838 (N_1838,N_1793,N_1774);
nand U1839 (N_1839,N_1795,N_1737);
or U1840 (N_1840,N_1712,N_1726);
or U1841 (N_1841,N_1728,N_1789);
nor U1842 (N_1842,N_1752,N_1777);
and U1843 (N_1843,N_1740,N_1761);
nor U1844 (N_1844,N_1707,N_1775);
nand U1845 (N_1845,N_1720,N_1758);
and U1846 (N_1846,N_1787,N_1762);
nor U1847 (N_1847,N_1757,N_1764);
nor U1848 (N_1848,N_1798,N_1727);
or U1849 (N_1849,N_1784,N_1782);
nor U1850 (N_1850,N_1745,N_1770);
and U1851 (N_1851,N_1747,N_1798);
nor U1852 (N_1852,N_1777,N_1708);
nor U1853 (N_1853,N_1790,N_1713);
or U1854 (N_1854,N_1714,N_1706);
nor U1855 (N_1855,N_1769,N_1757);
nand U1856 (N_1856,N_1730,N_1732);
nor U1857 (N_1857,N_1759,N_1726);
and U1858 (N_1858,N_1762,N_1724);
xnor U1859 (N_1859,N_1719,N_1784);
and U1860 (N_1860,N_1740,N_1784);
or U1861 (N_1861,N_1760,N_1780);
nand U1862 (N_1862,N_1791,N_1746);
nand U1863 (N_1863,N_1794,N_1741);
nand U1864 (N_1864,N_1736,N_1707);
nand U1865 (N_1865,N_1726,N_1725);
or U1866 (N_1866,N_1730,N_1748);
or U1867 (N_1867,N_1708,N_1761);
and U1868 (N_1868,N_1714,N_1777);
nand U1869 (N_1869,N_1711,N_1776);
or U1870 (N_1870,N_1734,N_1728);
or U1871 (N_1871,N_1716,N_1750);
xnor U1872 (N_1872,N_1786,N_1767);
or U1873 (N_1873,N_1715,N_1704);
nor U1874 (N_1874,N_1719,N_1710);
or U1875 (N_1875,N_1790,N_1732);
or U1876 (N_1876,N_1746,N_1739);
nor U1877 (N_1877,N_1765,N_1701);
nor U1878 (N_1878,N_1709,N_1794);
nand U1879 (N_1879,N_1793,N_1743);
or U1880 (N_1880,N_1787,N_1728);
or U1881 (N_1881,N_1792,N_1727);
nand U1882 (N_1882,N_1739,N_1799);
and U1883 (N_1883,N_1708,N_1756);
and U1884 (N_1884,N_1771,N_1701);
nor U1885 (N_1885,N_1759,N_1782);
or U1886 (N_1886,N_1753,N_1701);
nand U1887 (N_1887,N_1752,N_1754);
nor U1888 (N_1888,N_1772,N_1775);
or U1889 (N_1889,N_1717,N_1762);
nor U1890 (N_1890,N_1766,N_1734);
xnor U1891 (N_1891,N_1767,N_1782);
or U1892 (N_1892,N_1727,N_1743);
xnor U1893 (N_1893,N_1708,N_1784);
nand U1894 (N_1894,N_1710,N_1784);
or U1895 (N_1895,N_1709,N_1703);
nor U1896 (N_1896,N_1759,N_1728);
or U1897 (N_1897,N_1775,N_1726);
nor U1898 (N_1898,N_1770,N_1718);
nor U1899 (N_1899,N_1749,N_1747);
and U1900 (N_1900,N_1894,N_1822);
and U1901 (N_1901,N_1843,N_1806);
nand U1902 (N_1902,N_1891,N_1817);
and U1903 (N_1903,N_1872,N_1824);
nand U1904 (N_1904,N_1811,N_1852);
or U1905 (N_1905,N_1835,N_1854);
nor U1906 (N_1906,N_1881,N_1836);
and U1907 (N_1907,N_1897,N_1803);
xnor U1908 (N_1908,N_1880,N_1826);
nor U1909 (N_1909,N_1865,N_1884);
nor U1910 (N_1910,N_1812,N_1805);
or U1911 (N_1911,N_1885,N_1810);
or U1912 (N_1912,N_1873,N_1815);
nand U1913 (N_1913,N_1828,N_1899);
or U1914 (N_1914,N_1839,N_1847);
or U1915 (N_1915,N_1896,N_1819);
or U1916 (N_1916,N_1802,N_1820);
and U1917 (N_1917,N_1851,N_1849);
and U1918 (N_1918,N_1816,N_1800);
or U1919 (N_1919,N_1809,N_1878);
or U1920 (N_1920,N_1823,N_1832);
and U1921 (N_1921,N_1887,N_1818);
and U1922 (N_1922,N_1868,N_1845);
nor U1923 (N_1923,N_1883,N_1864);
nand U1924 (N_1924,N_1888,N_1814);
and U1925 (N_1925,N_1831,N_1876);
and U1926 (N_1926,N_1848,N_1829);
nor U1927 (N_1927,N_1858,N_1863);
and U1928 (N_1928,N_1877,N_1833);
or U1929 (N_1929,N_1862,N_1825);
nand U1930 (N_1930,N_1807,N_1861);
or U1931 (N_1931,N_1837,N_1859);
nor U1932 (N_1932,N_1892,N_1875);
nor U1933 (N_1933,N_1842,N_1838);
nand U1934 (N_1934,N_1840,N_1804);
nand U1935 (N_1935,N_1886,N_1853);
and U1936 (N_1936,N_1841,N_1866);
and U1937 (N_1937,N_1893,N_1856);
and U1938 (N_1938,N_1827,N_1813);
nand U1939 (N_1939,N_1898,N_1879);
and U1940 (N_1940,N_1882,N_1890);
or U1941 (N_1941,N_1830,N_1821);
or U1942 (N_1942,N_1889,N_1844);
nand U1943 (N_1943,N_1895,N_1850);
and U1944 (N_1944,N_1869,N_1857);
nor U1945 (N_1945,N_1808,N_1860);
nor U1946 (N_1946,N_1867,N_1855);
or U1947 (N_1947,N_1874,N_1870);
nor U1948 (N_1948,N_1871,N_1846);
nand U1949 (N_1949,N_1834,N_1801);
nand U1950 (N_1950,N_1864,N_1858);
and U1951 (N_1951,N_1839,N_1859);
nand U1952 (N_1952,N_1899,N_1888);
nor U1953 (N_1953,N_1815,N_1808);
nand U1954 (N_1954,N_1814,N_1884);
or U1955 (N_1955,N_1891,N_1873);
nor U1956 (N_1956,N_1875,N_1828);
nor U1957 (N_1957,N_1879,N_1827);
or U1958 (N_1958,N_1806,N_1842);
and U1959 (N_1959,N_1824,N_1807);
nand U1960 (N_1960,N_1898,N_1859);
or U1961 (N_1961,N_1845,N_1821);
and U1962 (N_1962,N_1862,N_1884);
or U1963 (N_1963,N_1804,N_1838);
nor U1964 (N_1964,N_1848,N_1803);
nor U1965 (N_1965,N_1881,N_1846);
nand U1966 (N_1966,N_1889,N_1883);
nor U1967 (N_1967,N_1884,N_1897);
and U1968 (N_1968,N_1801,N_1809);
nor U1969 (N_1969,N_1837,N_1847);
nor U1970 (N_1970,N_1832,N_1848);
or U1971 (N_1971,N_1878,N_1858);
and U1972 (N_1972,N_1864,N_1889);
and U1973 (N_1973,N_1849,N_1899);
or U1974 (N_1974,N_1809,N_1884);
nand U1975 (N_1975,N_1874,N_1876);
and U1976 (N_1976,N_1824,N_1874);
nor U1977 (N_1977,N_1825,N_1827);
nand U1978 (N_1978,N_1827,N_1886);
nand U1979 (N_1979,N_1857,N_1855);
or U1980 (N_1980,N_1868,N_1894);
and U1981 (N_1981,N_1833,N_1863);
and U1982 (N_1982,N_1844,N_1869);
and U1983 (N_1983,N_1819,N_1895);
nor U1984 (N_1984,N_1839,N_1894);
or U1985 (N_1985,N_1894,N_1812);
and U1986 (N_1986,N_1865,N_1859);
nand U1987 (N_1987,N_1846,N_1847);
nor U1988 (N_1988,N_1828,N_1893);
nand U1989 (N_1989,N_1893,N_1830);
and U1990 (N_1990,N_1822,N_1873);
xnor U1991 (N_1991,N_1820,N_1855);
nor U1992 (N_1992,N_1844,N_1873);
and U1993 (N_1993,N_1816,N_1832);
nor U1994 (N_1994,N_1823,N_1876);
nor U1995 (N_1995,N_1824,N_1877);
and U1996 (N_1996,N_1882,N_1832);
and U1997 (N_1997,N_1886,N_1849);
or U1998 (N_1998,N_1844,N_1849);
nor U1999 (N_1999,N_1827,N_1851);
nor U2000 (N_2000,N_1969,N_1983);
nand U2001 (N_2001,N_1981,N_1925);
or U2002 (N_2002,N_1948,N_1993);
or U2003 (N_2003,N_1960,N_1936);
nand U2004 (N_2004,N_1980,N_1963);
nor U2005 (N_2005,N_1997,N_1905);
nand U2006 (N_2006,N_1998,N_1911);
or U2007 (N_2007,N_1932,N_1924);
xnor U2008 (N_2008,N_1938,N_1907);
nor U2009 (N_2009,N_1937,N_1929);
nor U2010 (N_2010,N_1957,N_1962);
or U2011 (N_2011,N_1978,N_1972);
nand U2012 (N_2012,N_1914,N_1927);
nor U2013 (N_2013,N_1989,N_1946);
or U2014 (N_2014,N_1912,N_1943);
or U2015 (N_2015,N_1903,N_1994);
or U2016 (N_2016,N_1967,N_1922);
and U2017 (N_2017,N_1923,N_1906);
or U2018 (N_2018,N_1949,N_1951);
xor U2019 (N_2019,N_1992,N_1999);
nor U2020 (N_2020,N_1935,N_1956);
xnor U2021 (N_2021,N_1934,N_1970);
and U2022 (N_2022,N_1982,N_1995);
nor U2023 (N_2023,N_1910,N_1973);
or U2024 (N_2024,N_1909,N_1974);
nand U2025 (N_2025,N_1926,N_1954);
nor U2026 (N_2026,N_1940,N_1953);
or U2027 (N_2027,N_1966,N_1987);
and U2028 (N_2028,N_1955,N_1920);
or U2029 (N_2029,N_1996,N_1918);
and U2030 (N_2030,N_1976,N_1947);
and U2031 (N_2031,N_1950,N_1917);
nand U2032 (N_2032,N_1939,N_1916);
and U2033 (N_2033,N_1915,N_1933);
nor U2034 (N_2034,N_1986,N_1958);
nand U2035 (N_2035,N_1900,N_1941);
or U2036 (N_2036,N_1928,N_1919);
or U2037 (N_2037,N_1904,N_1988);
nor U2038 (N_2038,N_1931,N_1913);
nand U2039 (N_2039,N_1991,N_1942);
or U2040 (N_2040,N_1902,N_1975);
nand U2041 (N_2041,N_1944,N_1945);
nand U2042 (N_2042,N_1908,N_1971);
nand U2043 (N_2043,N_1990,N_1961);
nor U2044 (N_2044,N_1959,N_1921);
nand U2045 (N_2045,N_1968,N_1964);
nand U2046 (N_2046,N_1930,N_1977);
or U2047 (N_2047,N_1952,N_1985);
and U2048 (N_2048,N_1979,N_1965);
or U2049 (N_2049,N_1901,N_1984);
nor U2050 (N_2050,N_1951,N_1936);
nor U2051 (N_2051,N_1908,N_1914);
nand U2052 (N_2052,N_1978,N_1933);
or U2053 (N_2053,N_1951,N_1966);
or U2054 (N_2054,N_1967,N_1941);
nand U2055 (N_2055,N_1969,N_1973);
and U2056 (N_2056,N_1988,N_1915);
nand U2057 (N_2057,N_1906,N_1967);
and U2058 (N_2058,N_1909,N_1972);
and U2059 (N_2059,N_1967,N_1918);
and U2060 (N_2060,N_1915,N_1914);
and U2061 (N_2061,N_1902,N_1990);
nand U2062 (N_2062,N_1987,N_1925);
nand U2063 (N_2063,N_1943,N_1909);
and U2064 (N_2064,N_1970,N_1929);
or U2065 (N_2065,N_1960,N_1949);
and U2066 (N_2066,N_1906,N_1934);
and U2067 (N_2067,N_1942,N_1989);
nand U2068 (N_2068,N_1931,N_1953);
xnor U2069 (N_2069,N_1962,N_1913);
nor U2070 (N_2070,N_1945,N_1992);
and U2071 (N_2071,N_1935,N_1955);
or U2072 (N_2072,N_1995,N_1977);
or U2073 (N_2073,N_1902,N_1916);
or U2074 (N_2074,N_1954,N_1969);
or U2075 (N_2075,N_1918,N_1969);
nor U2076 (N_2076,N_1931,N_1938);
and U2077 (N_2077,N_1915,N_1930);
nor U2078 (N_2078,N_1941,N_1988);
nand U2079 (N_2079,N_1951,N_1903);
and U2080 (N_2080,N_1920,N_1994);
nand U2081 (N_2081,N_1950,N_1923);
and U2082 (N_2082,N_1955,N_1937);
and U2083 (N_2083,N_1993,N_1941);
and U2084 (N_2084,N_1918,N_1901);
or U2085 (N_2085,N_1972,N_1995);
and U2086 (N_2086,N_1910,N_1990);
and U2087 (N_2087,N_1990,N_1928);
nor U2088 (N_2088,N_1997,N_1991);
or U2089 (N_2089,N_1900,N_1931);
nand U2090 (N_2090,N_1962,N_1983);
nand U2091 (N_2091,N_1949,N_1921);
and U2092 (N_2092,N_1995,N_1955);
xor U2093 (N_2093,N_1984,N_1944);
or U2094 (N_2094,N_1919,N_1950);
xnor U2095 (N_2095,N_1913,N_1964);
or U2096 (N_2096,N_1997,N_1964);
or U2097 (N_2097,N_1937,N_1914);
and U2098 (N_2098,N_1938,N_1939);
nor U2099 (N_2099,N_1925,N_1995);
or U2100 (N_2100,N_2007,N_2040);
nor U2101 (N_2101,N_2064,N_2048);
nand U2102 (N_2102,N_2083,N_2094);
or U2103 (N_2103,N_2014,N_2049);
or U2104 (N_2104,N_2006,N_2051);
nand U2105 (N_2105,N_2059,N_2066);
and U2106 (N_2106,N_2052,N_2019);
or U2107 (N_2107,N_2032,N_2054);
xnor U2108 (N_2108,N_2025,N_2062);
and U2109 (N_2109,N_2043,N_2079);
and U2110 (N_2110,N_2009,N_2002);
nor U2111 (N_2111,N_2013,N_2057);
and U2112 (N_2112,N_2060,N_2071);
nor U2113 (N_2113,N_2078,N_2041);
nand U2114 (N_2114,N_2020,N_2090);
nand U2115 (N_2115,N_2005,N_2080);
nand U2116 (N_2116,N_2092,N_2017);
nand U2117 (N_2117,N_2055,N_2097);
nand U2118 (N_2118,N_2058,N_2023);
nand U2119 (N_2119,N_2028,N_2036);
nand U2120 (N_2120,N_2045,N_2076);
and U2121 (N_2121,N_2082,N_2075);
or U2122 (N_2122,N_2037,N_2016);
or U2123 (N_2123,N_2047,N_2022);
or U2124 (N_2124,N_2069,N_2018);
or U2125 (N_2125,N_2026,N_2004);
or U2126 (N_2126,N_2073,N_2030);
nand U2127 (N_2127,N_2012,N_2089);
nand U2128 (N_2128,N_2033,N_2096);
or U2129 (N_2129,N_2053,N_2087);
and U2130 (N_2130,N_2029,N_2093);
nor U2131 (N_2131,N_2063,N_2084);
or U2132 (N_2132,N_2015,N_2070);
and U2133 (N_2133,N_2098,N_2001);
or U2134 (N_2134,N_2067,N_2061);
nand U2135 (N_2135,N_2068,N_2081);
nor U2136 (N_2136,N_2024,N_2046);
nand U2137 (N_2137,N_2008,N_2050);
xor U2138 (N_2138,N_2044,N_2091);
and U2139 (N_2139,N_2074,N_2056);
nand U2140 (N_2140,N_2039,N_2035);
nand U2141 (N_2141,N_2003,N_2034);
and U2142 (N_2142,N_2086,N_2010);
and U2143 (N_2143,N_2031,N_2072);
or U2144 (N_2144,N_2027,N_2038);
nor U2145 (N_2145,N_2099,N_2021);
nor U2146 (N_2146,N_2042,N_2000);
and U2147 (N_2147,N_2095,N_2088);
nand U2148 (N_2148,N_2085,N_2011);
and U2149 (N_2149,N_2077,N_2065);
or U2150 (N_2150,N_2045,N_2061);
and U2151 (N_2151,N_2073,N_2037);
or U2152 (N_2152,N_2030,N_2033);
or U2153 (N_2153,N_2025,N_2072);
nor U2154 (N_2154,N_2046,N_2033);
or U2155 (N_2155,N_2096,N_2056);
and U2156 (N_2156,N_2087,N_2055);
nand U2157 (N_2157,N_2015,N_2057);
nor U2158 (N_2158,N_2001,N_2069);
xnor U2159 (N_2159,N_2074,N_2045);
and U2160 (N_2160,N_2053,N_2017);
nor U2161 (N_2161,N_2014,N_2029);
nor U2162 (N_2162,N_2014,N_2070);
and U2163 (N_2163,N_2013,N_2054);
or U2164 (N_2164,N_2041,N_2092);
nor U2165 (N_2165,N_2051,N_2010);
nor U2166 (N_2166,N_2069,N_2076);
or U2167 (N_2167,N_2072,N_2080);
and U2168 (N_2168,N_2080,N_2057);
nand U2169 (N_2169,N_2044,N_2072);
nand U2170 (N_2170,N_2042,N_2006);
or U2171 (N_2171,N_2077,N_2010);
nand U2172 (N_2172,N_2064,N_2006);
xnor U2173 (N_2173,N_2008,N_2055);
nand U2174 (N_2174,N_2093,N_2025);
or U2175 (N_2175,N_2060,N_2091);
nand U2176 (N_2176,N_2053,N_2093);
nand U2177 (N_2177,N_2056,N_2040);
or U2178 (N_2178,N_2002,N_2067);
and U2179 (N_2179,N_2072,N_2065);
or U2180 (N_2180,N_2065,N_2027);
or U2181 (N_2181,N_2029,N_2097);
nor U2182 (N_2182,N_2036,N_2060);
nand U2183 (N_2183,N_2014,N_2010);
xor U2184 (N_2184,N_2028,N_2082);
or U2185 (N_2185,N_2023,N_2059);
nand U2186 (N_2186,N_2090,N_2040);
and U2187 (N_2187,N_2017,N_2034);
or U2188 (N_2188,N_2046,N_2073);
and U2189 (N_2189,N_2041,N_2019);
nand U2190 (N_2190,N_2033,N_2079);
nand U2191 (N_2191,N_2003,N_2038);
nand U2192 (N_2192,N_2036,N_2098);
and U2193 (N_2193,N_2003,N_2076);
and U2194 (N_2194,N_2094,N_2013);
and U2195 (N_2195,N_2032,N_2093);
and U2196 (N_2196,N_2023,N_2010);
or U2197 (N_2197,N_2084,N_2058);
and U2198 (N_2198,N_2046,N_2098);
nand U2199 (N_2199,N_2072,N_2048);
and U2200 (N_2200,N_2134,N_2138);
and U2201 (N_2201,N_2131,N_2137);
or U2202 (N_2202,N_2194,N_2189);
nor U2203 (N_2203,N_2143,N_2171);
nor U2204 (N_2204,N_2151,N_2152);
nor U2205 (N_2205,N_2145,N_2181);
xor U2206 (N_2206,N_2106,N_2177);
and U2207 (N_2207,N_2182,N_2150);
nand U2208 (N_2208,N_2133,N_2179);
nor U2209 (N_2209,N_2193,N_2123);
and U2210 (N_2210,N_2117,N_2109);
and U2211 (N_2211,N_2139,N_2184);
and U2212 (N_2212,N_2136,N_2168);
and U2213 (N_2213,N_2164,N_2163);
nor U2214 (N_2214,N_2142,N_2119);
nor U2215 (N_2215,N_2128,N_2146);
nor U2216 (N_2216,N_2198,N_2159);
nand U2217 (N_2217,N_2147,N_2175);
and U2218 (N_2218,N_2118,N_2155);
or U2219 (N_2219,N_2108,N_2105);
nor U2220 (N_2220,N_2174,N_2183);
nor U2221 (N_2221,N_2122,N_2148);
nand U2222 (N_2222,N_2186,N_2104);
or U2223 (N_2223,N_2169,N_2141);
and U2224 (N_2224,N_2190,N_2129);
or U2225 (N_2225,N_2154,N_2172);
or U2226 (N_2226,N_2178,N_2107);
or U2227 (N_2227,N_2120,N_2170);
or U2228 (N_2228,N_2187,N_2153);
nand U2229 (N_2229,N_2127,N_2135);
and U2230 (N_2230,N_2158,N_2111);
nor U2231 (N_2231,N_2140,N_2110);
nor U2232 (N_2232,N_2114,N_2160);
nand U2233 (N_2233,N_2125,N_2102);
nand U2234 (N_2234,N_2176,N_2126);
nor U2235 (N_2235,N_2121,N_2132);
or U2236 (N_2236,N_2157,N_2191);
or U2237 (N_2237,N_2124,N_2166);
nor U2238 (N_2238,N_2196,N_2100);
nor U2239 (N_2239,N_2101,N_2167);
xnor U2240 (N_2240,N_2197,N_2185);
nor U2241 (N_2241,N_2162,N_2188);
nor U2242 (N_2242,N_2113,N_2115);
and U2243 (N_2243,N_2149,N_2180);
nand U2244 (N_2244,N_2116,N_2130);
and U2245 (N_2245,N_2103,N_2112);
or U2246 (N_2246,N_2156,N_2144);
nor U2247 (N_2247,N_2199,N_2195);
and U2248 (N_2248,N_2161,N_2173);
or U2249 (N_2249,N_2165,N_2192);
and U2250 (N_2250,N_2118,N_2190);
or U2251 (N_2251,N_2137,N_2112);
or U2252 (N_2252,N_2174,N_2130);
nor U2253 (N_2253,N_2153,N_2194);
nor U2254 (N_2254,N_2113,N_2145);
nor U2255 (N_2255,N_2141,N_2165);
and U2256 (N_2256,N_2133,N_2113);
nor U2257 (N_2257,N_2107,N_2171);
and U2258 (N_2258,N_2189,N_2102);
nor U2259 (N_2259,N_2132,N_2156);
or U2260 (N_2260,N_2137,N_2102);
nand U2261 (N_2261,N_2177,N_2139);
xor U2262 (N_2262,N_2179,N_2165);
nand U2263 (N_2263,N_2116,N_2148);
and U2264 (N_2264,N_2178,N_2183);
nor U2265 (N_2265,N_2185,N_2158);
nand U2266 (N_2266,N_2189,N_2160);
or U2267 (N_2267,N_2168,N_2112);
nor U2268 (N_2268,N_2102,N_2121);
nand U2269 (N_2269,N_2173,N_2183);
nor U2270 (N_2270,N_2192,N_2116);
nand U2271 (N_2271,N_2106,N_2168);
nor U2272 (N_2272,N_2127,N_2169);
nand U2273 (N_2273,N_2169,N_2122);
or U2274 (N_2274,N_2154,N_2174);
or U2275 (N_2275,N_2138,N_2101);
nor U2276 (N_2276,N_2106,N_2119);
nor U2277 (N_2277,N_2137,N_2198);
or U2278 (N_2278,N_2113,N_2128);
or U2279 (N_2279,N_2104,N_2150);
nand U2280 (N_2280,N_2109,N_2166);
nand U2281 (N_2281,N_2182,N_2131);
nor U2282 (N_2282,N_2169,N_2154);
nor U2283 (N_2283,N_2165,N_2199);
nor U2284 (N_2284,N_2135,N_2141);
or U2285 (N_2285,N_2197,N_2164);
or U2286 (N_2286,N_2165,N_2122);
and U2287 (N_2287,N_2113,N_2144);
and U2288 (N_2288,N_2138,N_2157);
nand U2289 (N_2289,N_2109,N_2103);
and U2290 (N_2290,N_2146,N_2123);
nand U2291 (N_2291,N_2110,N_2118);
nand U2292 (N_2292,N_2114,N_2161);
and U2293 (N_2293,N_2123,N_2130);
nand U2294 (N_2294,N_2123,N_2105);
nand U2295 (N_2295,N_2175,N_2199);
nand U2296 (N_2296,N_2103,N_2149);
xor U2297 (N_2297,N_2190,N_2198);
and U2298 (N_2298,N_2171,N_2194);
nor U2299 (N_2299,N_2117,N_2169);
nand U2300 (N_2300,N_2293,N_2298);
nor U2301 (N_2301,N_2241,N_2285);
nor U2302 (N_2302,N_2227,N_2295);
nor U2303 (N_2303,N_2296,N_2223);
or U2304 (N_2304,N_2265,N_2284);
and U2305 (N_2305,N_2280,N_2269);
and U2306 (N_2306,N_2250,N_2277);
nand U2307 (N_2307,N_2207,N_2274);
or U2308 (N_2308,N_2268,N_2264);
nor U2309 (N_2309,N_2239,N_2242);
nand U2310 (N_2310,N_2259,N_2234);
nand U2311 (N_2311,N_2292,N_2246);
xor U2312 (N_2312,N_2283,N_2263);
nand U2313 (N_2313,N_2238,N_2279);
nor U2314 (N_2314,N_2249,N_2218);
or U2315 (N_2315,N_2226,N_2244);
nand U2316 (N_2316,N_2270,N_2253);
or U2317 (N_2317,N_2212,N_2240);
nand U2318 (N_2318,N_2290,N_2267);
and U2319 (N_2319,N_2233,N_2282);
nor U2320 (N_2320,N_2230,N_2281);
or U2321 (N_2321,N_2257,N_2261);
nor U2322 (N_2322,N_2213,N_2215);
nand U2323 (N_2323,N_2245,N_2210);
nand U2324 (N_2324,N_2252,N_2299);
and U2325 (N_2325,N_2208,N_2237);
nand U2326 (N_2326,N_2222,N_2228);
and U2327 (N_2327,N_2201,N_2200);
or U2328 (N_2328,N_2225,N_2291);
or U2329 (N_2329,N_2254,N_2272);
or U2330 (N_2330,N_2273,N_2258);
or U2331 (N_2331,N_2266,N_2286);
and U2332 (N_2332,N_2243,N_2256);
nor U2333 (N_2333,N_2235,N_2219);
and U2334 (N_2334,N_2203,N_2275);
nor U2335 (N_2335,N_2232,N_2229);
nor U2336 (N_2336,N_2294,N_2216);
nand U2337 (N_2337,N_2271,N_2262);
nand U2338 (N_2338,N_2260,N_2289);
or U2339 (N_2339,N_2236,N_2247);
nor U2340 (N_2340,N_2217,N_2221);
or U2341 (N_2341,N_2206,N_2211);
and U2342 (N_2342,N_2251,N_2224);
nor U2343 (N_2343,N_2202,N_2204);
nor U2344 (N_2344,N_2209,N_2205);
nand U2345 (N_2345,N_2287,N_2214);
and U2346 (N_2346,N_2248,N_2255);
nor U2347 (N_2347,N_2278,N_2276);
or U2348 (N_2348,N_2231,N_2288);
nand U2349 (N_2349,N_2297,N_2220);
or U2350 (N_2350,N_2295,N_2254);
or U2351 (N_2351,N_2297,N_2231);
or U2352 (N_2352,N_2200,N_2281);
or U2353 (N_2353,N_2294,N_2235);
and U2354 (N_2354,N_2271,N_2247);
nand U2355 (N_2355,N_2256,N_2299);
nor U2356 (N_2356,N_2236,N_2280);
nand U2357 (N_2357,N_2203,N_2225);
nor U2358 (N_2358,N_2265,N_2226);
nor U2359 (N_2359,N_2213,N_2247);
or U2360 (N_2360,N_2224,N_2282);
and U2361 (N_2361,N_2286,N_2275);
nor U2362 (N_2362,N_2240,N_2261);
nand U2363 (N_2363,N_2217,N_2286);
and U2364 (N_2364,N_2226,N_2281);
nor U2365 (N_2365,N_2291,N_2222);
and U2366 (N_2366,N_2262,N_2220);
or U2367 (N_2367,N_2277,N_2246);
or U2368 (N_2368,N_2200,N_2240);
xor U2369 (N_2369,N_2213,N_2228);
and U2370 (N_2370,N_2268,N_2242);
nor U2371 (N_2371,N_2212,N_2236);
nand U2372 (N_2372,N_2282,N_2255);
or U2373 (N_2373,N_2279,N_2284);
nor U2374 (N_2374,N_2282,N_2278);
nor U2375 (N_2375,N_2295,N_2210);
or U2376 (N_2376,N_2248,N_2221);
nor U2377 (N_2377,N_2274,N_2206);
nand U2378 (N_2378,N_2246,N_2263);
and U2379 (N_2379,N_2218,N_2294);
nor U2380 (N_2380,N_2285,N_2255);
nor U2381 (N_2381,N_2296,N_2258);
nor U2382 (N_2382,N_2224,N_2252);
or U2383 (N_2383,N_2225,N_2246);
or U2384 (N_2384,N_2295,N_2235);
or U2385 (N_2385,N_2246,N_2251);
nand U2386 (N_2386,N_2283,N_2266);
or U2387 (N_2387,N_2293,N_2232);
and U2388 (N_2388,N_2238,N_2248);
nor U2389 (N_2389,N_2206,N_2258);
nor U2390 (N_2390,N_2267,N_2257);
and U2391 (N_2391,N_2253,N_2296);
or U2392 (N_2392,N_2271,N_2295);
nand U2393 (N_2393,N_2267,N_2202);
nor U2394 (N_2394,N_2224,N_2271);
and U2395 (N_2395,N_2273,N_2219);
or U2396 (N_2396,N_2222,N_2266);
nand U2397 (N_2397,N_2231,N_2238);
or U2398 (N_2398,N_2288,N_2236);
nand U2399 (N_2399,N_2201,N_2273);
xor U2400 (N_2400,N_2349,N_2352);
and U2401 (N_2401,N_2391,N_2394);
nand U2402 (N_2402,N_2329,N_2353);
nand U2403 (N_2403,N_2367,N_2354);
nor U2404 (N_2404,N_2381,N_2377);
or U2405 (N_2405,N_2386,N_2314);
and U2406 (N_2406,N_2310,N_2316);
nand U2407 (N_2407,N_2385,N_2340);
or U2408 (N_2408,N_2360,N_2372);
and U2409 (N_2409,N_2389,N_2382);
nor U2410 (N_2410,N_2309,N_2331);
and U2411 (N_2411,N_2319,N_2311);
nand U2412 (N_2412,N_2355,N_2374);
nor U2413 (N_2413,N_2344,N_2398);
nor U2414 (N_2414,N_2336,N_2363);
nor U2415 (N_2415,N_2312,N_2332);
nand U2416 (N_2416,N_2368,N_2393);
or U2417 (N_2417,N_2345,N_2350);
nor U2418 (N_2418,N_2392,N_2337);
nor U2419 (N_2419,N_2303,N_2395);
and U2420 (N_2420,N_2313,N_2357);
or U2421 (N_2421,N_2301,N_2343);
nor U2422 (N_2422,N_2317,N_2396);
nor U2423 (N_2423,N_2365,N_2308);
nor U2424 (N_2424,N_2384,N_2302);
and U2425 (N_2425,N_2306,N_2339);
or U2426 (N_2426,N_2348,N_2358);
and U2427 (N_2427,N_2346,N_2379);
nor U2428 (N_2428,N_2304,N_2338);
nand U2429 (N_2429,N_2333,N_2334);
nor U2430 (N_2430,N_2369,N_2300);
and U2431 (N_2431,N_2375,N_2335);
nand U2432 (N_2432,N_2373,N_2321);
nor U2433 (N_2433,N_2325,N_2362);
or U2434 (N_2434,N_2328,N_2370);
xor U2435 (N_2435,N_2342,N_2397);
or U2436 (N_2436,N_2341,N_2327);
nand U2437 (N_2437,N_2390,N_2318);
and U2438 (N_2438,N_2347,N_2330);
nand U2439 (N_2439,N_2364,N_2378);
nor U2440 (N_2440,N_2320,N_2376);
and U2441 (N_2441,N_2359,N_2399);
and U2442 (N_2442,N_2388,N_2322);
nor U2443 (N_2443,N_2361,N_2305);
nor U2444 (N_2444,N_2366,N_2380);
nor U2445 (N_2445,N_2371,N_2315);
nand U2446 (N_2446,N_2307,N_2324);
or U2447 (N_2447,N_2351,N_2323);
or U2448 (N_2448,N_2326,N_2387);
nor U2449 (N_2449,N_2356,N_2383);
and U2450 (N_2450,N_2346,N_2390);
and U2451 (N_2451,N_2381,N_2333);
or U2452 (N_2452,N_2321,N_2353);
and U2453 (N_2453,N_2383,N_2354);
and U2454 (N_2454,N_2301,N_2383);
and U2455 (N_2455,N_2370,N_2356);
or U2456 (N_2456,N_2308,N_2379);
nor U2457 (N_2457,N_2371,N_2353);
and U2458 (N_2458,N_2341,N_2371);
and U2459 (N_2459,N_2384,N_2361);
nor U2460 (N_2460,N_2328,N_2316);
nor U2461 (N_2461,N_2382,N_2320);
and U2462 (N_2462,N_2387,N_2309);
nor U2463 (N_2463,N_2378,N_2307);
and U2464 (N_2464,N_2388,N_2356);
nor U2465 (N_2465,N_2316,N_2305);
nand U2466 (N_2466,N_2315,N_2377);
and U2467 (N_2467,N_2386,N_2356);
nand U2468 (N_2468,N_2326,N_2343);
or U2469 (N_2469,N_2328,N_2337);
nand U2470 (N_2470,N_2350,N_2336);
and U2471 (N_2471,N_2318,N_2391);
and U2472 (N_2472,N_2396,N_2307);
xnor U2473 (N_2473,N_2353,N_2319);
nor U2474 (N_2474,N_2341,N_2394);
nor U2475 (N_2475,N_2347,N_2319);
nand U2476 (N_2476,N_2348,N_2376);
and U2477 (N_2477,N_2357,N_2343);
and U2478 (N_2478,N_2391,N_2348);
or U2479 (N_2479,N_2325,N_2356);
nand U2480 (N_2480,N_2347,N_2308);
nand U2481 (N_2481,N_2346,N_2338);
and U2482 (N_2482,N_2371,N_2350);
nand U2483 (N_2483,N_2374,N_2352);
nand U2484 (N_2484,N_2364,N_2376);
nand U2485 (N_2485,N_2312,N_2329);
nor U2486 (N_2486,N_2350,N_2365);
and U2487 (N_2487,N_2346,N_2380);
nor U2488 (N_2488,N_2384,N_2342);
nor U2489 (N_2489,N_2334,N_2347);
and U2490 (N_2490,N_2368,N_2310);
or U2491 (N_2491,N_2398,N_2384);
nor U2492 (N_2492,N_2359,N_2310);
nor U2493 (N_2493,N_2375,N_2377);
nor U2494 (N_2494,N_2302,N_2383);
or U2495 (N_2495,N_2374,N_2382);
nor U2496 (N_2496,N_2388,N_2321);
and U2497 (N_2497,N_2336,N_2380);
and U2498 (N_2498,N_2386,N_2363);
or U2499 (N_2499,N_2372,N_2344);
or U2500 (N_2500,N_2418,N_2407);
or U2501 (N_2501,N_2466,N_2441);
nand U2502 (N_2502,N_2435,N_2474);
nand U2503 (N_2503,N_2429,N_2477);
nor U2504 (N_2504,N_2412,N_2449);
or U2505 (N_2505,N_2454,N_2492);
nand U2506 (N_2506,N_2445,N_2462);
and U2507 (N_2507,N_2450,N_2434);
nand U2508 (N_2508,N_2497,N_2408);
nand U2509 (N_2509,N_2458,N_2444);
nand U2510 (N_2510,N_2425,N_2448);
and U2511 (N_2511,N_2410,N_2489);
xnor U2512 (N_2512,N_2485,N_2433);
nand U2513 (N_2513,N_2414,N_2438);
and U2514 (N_2514,N_2476,N_2487);
nand U2515 (N_2515,N_2424,N_2478);
xnor U2516 (N_2516,N_2459,N_2437);
and U2517 (N_2517,N_2480,N_2420);
and U2518 (N_2518,N_2453,N_2421);
nor U2519 (N_2519,N_2439,N_2427);
or U2520 (N_2520,N_2455,N_2402);
nand U2521 (N_2521,N_2482,N_2432);
xnor U2522 (N_2522,N_2481,N_2409);
or U2523 (N_2523,N_2401,N_2484);
nor U2524 (N_2524,N_2415,N_2457);
nor U2525 (N_2525,N_2488,N_2467);
nand U2526 (N_2526,N_2490,N_2486);
or U2527 (N_2527,N_2495,N_2447);
nand U2528 (N_2528,N_2442,N_2464);
nor U2529 (N_2529,N_2460,N_2436);
and U2530 (N_2530,N_2498,N_2494);
nor U2531 (N_2531,N_2468,N_2431);
or U2532 (N_2532,N_2419,N_2417);
nand U2533 (N_2533,N_2471,N_2400);
and U2534 (N_2534,N_2470,N_2404);
or U2535 (N_2535,N_2428,N_2496);
nand U2536 (N_2536,N_2423,N_2483);
nand U2537 (N_2537,N_2493,N_2456);
nand U2538 (N_2538,N_2403,N_2465);
or U2539 (N_2539,N_2440,N_2491);
nor U2540 (N_2540,N_2443,N_2446);
and U2541 (N_2541,N_2469,N_2411);
nand U2542 (N_2542,N_2473,N_2430);
nor U2543 (N_2543,N_2405,N_2426);
or U2544 (N_2544,N_2413,N_2452);
or U2545 (N_2545,N_2463,N_2422);
or U2546 (N_2546,N_2451,N_2416);
nand U2547 (N_2547,N_2461,N_2406);
nand U2548 (N_2548,N_2475,N_2472);
xnor U2549 (N_2549,N_2499,N_2479);
and U2550 (N_2550,N_2466,N_2495);
or U2551 (N_2551,N_2467,N_2457);
nor U2552 (N_2552,N_2401,N_2439);
nand U2553 (N_2553,N_2461,N_2430);
and U2554 (N_2554,N_2445,N_2441);
or U2555 (N_2555,N_2456,N_2460);
or U2556 (N_2556,N_2447,N_2492);
and U2557 (N_2557,N_2426,N_2438);
nor U2558 (N_2558,N_2452,N_2463);
and U2559 (N_2559,N_2427,N_2435);
nand U2560 (N_2560,N_2416,N_2423);
or U2561 (N_2561,N_2473,N_2477);
nor U2562 (N_2562,N_2498,N_2465);
nor U2563 (N_2563,N_2431,N_2498);
nand U2564 (N_2564,N_2488,N_2455);
nor U2565 (N_2565,N_2404,N_2475);
and U2566 (N_2566,N_2415,N_2435);
or U2567 (N_2567,N_2426,N_2476);
and U2568 (N_2568,N_2478,N_2422);
or U2569 (N_2569,N_2416,N_2444);
nand U2570 (N_2570,N_2496,N_2480);
nand U2571 (N_2571,N_2457,N_2470);
nor U2572 (N_2572,N_2411,N_2481);
nand U2573 (N_2573,N_2417,N_2400);
or U2574 (N_2574,N_2433,N_2455);
nor U2575 (N_2575,N_2465,N_2449);
or U2576 (N_2576,N_2414,N_2425);
and U2577 (N_2577,N_2465,N_2431);
and U2578 (N_2578,N_2458,N_2493);
and U2579 (N_2579,N_2448,N_2470);
nand U2580 (N_2580,N_2493,N_2417);
and U2581 (N_2581,N_2489,N_2447);
and U2582 (N_2582,N_2442,N_2444);
nand U2583 (N_2583,N_2441,N_2459);
nand U2584 (N_2584,N_2458,N_2439);
nand U2585 (N_2585,N_2439,N_2481);
nor U2586 (N_2586,N_2471,N_2411);
and U2587 (N_2587,N_2456,N_2407);
or U2588 (N_2588,N_2495,N_2461);
nand U2589 (N_2589,N_2469,N_2443);
and U2590 (N_2590,N_2462,N_2440);
nor U2591 (N_2591,N_2413,N_2498);
xnor U2592 (N_2592,N_2498,N_2469);
and U2593 (N_2593,N_2499,N_2469);
nor U2594 (N_2594,N_2492,N_2473);
nor U2595 (N_2595,N_2476,N_2472);
or U2596 (N_2596,N_2451,N_2439);
and U2597 (N_2597,N_2469,N_2448);
nor U2598 (N_2598,N_2405,N_2403);
or U2599 (N_2599,N_2479,N_2457);
nor U2600 (N_2600,N_2557,N_2577);
nor U2601 (N_2601,N_2553,N_2531);
nor U2602 (N_2602,N_2594,N_2595);
and U2603 (N_2603,N_2597,N_2546);
nor U2604 (N_2604,N_2504,N_2535);
and U2605 (N_2605,N_2506,N_2524);
nand U2606 (N_2606,N_2582,N_2566);
or U2607 (N_2607,N_2534,N_2563);
nor U2608 (N_2608,N_2585,N_2522);
nand U2609 (N_2609,N_2558,N_2575);
or U2610 (N_2610,N_2599,N_2526);
nor U2611 (N_2611,N_2552,N_2569);
nor U2612 (N_2612,N_2519,N_2516);
or U2613 (N_2613,N_2556,N_2521);
or U2614 (N_2614,N_2571,N_2573);
xor U2615 (N_2615,N_2503,N_2512);
and U2616 (N_2616,N_2505,N_2510);
nand U2617 (N_2617,N_2545,N_2513);
and U2618 (N_2618,N_2578,N_2529);
or U2619 (N_2619,N_2501,N_2525);
and U2620 (N_2620,N_2540,N_2561);
and U2621 (N_2621,N_2514,N_2502);
nor U2622 (N_2622,N_2507,N_2520);
nand U2623 (N_2623,N_2588,N_2517);
nor U2624 (N_2624,N_2565,N_2579);
nor U2625 (N_2625,N_2518,N_2500);
nor U2626 (N_2626,N_2593,N_2567);
nor U2627 (N_2627,N_2598,N_2544);
and U2628 (N_2628,N_2527,N_2564);
or U2629 (N_2629,N_2590,N_2554);
nor U2630 (N_2630,N_2562,N_2533);
or U2631 (N_2631,N_2509,N_2537);
nand U2632 (N_2632,N_2580,N_2574);
and U2633 (N_2633,N_2539,N_2592);
xor U2634 (N_2634,N_2584,N_2549);
nor U2635 (N_2635,N_2568,N_2591);
and U2636 (N_2636,N_2532,N_2589);
nand U2637 (N_2637,N_2581,N_2551);
nor U2638 (N_2638,N_2560,N_2511);
and U2639 (N_2639,N_2550,N_2538);
nand U2640 (N_2640,N_2523,N_2548);
nand U2641 (N_2641,N_2555,N_2572);
and U2642 (N_2642,N_2541,N_2508);
or U2643 (N_2643,N_2587,N_2543);
nand U2644 (N_2644,N_2559,N_2515);
and U2645 (N_2645,N_2586,N_2596);
nand U2646 (N_2646,N_2576,N_2542);
xnor U2647 (N_2647,N_2570,N_2530);
nor U2648 (N_2648,N_2547,N_2583);
nor U2649 (N_2649,N_2528,N_2536);
nor U2650 (N_2650,N_2514,N_2588);
nor U2651 (N_2651,N_2541,N_2563);
xor U2652 (N_2652,N_2580,N_2536);
nand U2653 (N_2653,N_2570,N_2548);
nand U2654 (N_2654,N_2502,N_2570);
nand U2655 (N_2655,N_2556,N_2536);
nor U2656 (N_2656,N_2544,N_2585);
nand U2657 (N_2657,N_2571,N_2522);
nand U2658 (N_2658,N_2544,N_2511);
nand U2659 (N_2659,N_2579,N_2529);
nor U2660 (N_2660,N_2540,N_2572);
or U2661 (N_2661,N_2585,N_2555);
nand U2662 (N_2662,N_2538,N_2575);
or U2663 (N_2663,N_2585,N_2579);
and U2664 (N_2664,N_2520,N_2552);
nor U2665 (N_2665,N_2511,N_2564);
and U2666 (N_2666,N_2541,N_2575);
or U2667 (N_2667,N_2549,N_2574);
nor U2668 (N_2668,N_2552,N_2500);
nand U2669 (N_2669,N_2506,N_2568);
or U2670 (N_2670,N_2598,N_2515);
and U2671 (N_2671,N_2501,N_2526);
and U2672 (N_2672,N_2517,N_2507);
or U2673 (N_2673,N_2574,N_2548);
nor U2674 (N_2674,N_2563,N_2593);
nor U2675 (N_2675,N_2569,N_2590);
and U2676 (N_2676,N_2560,N_2591);
nor U2677 (N_2677,N_2594,N_2507);
nor U2678 (N_2678,N_2587,N_2577);
nand U2679 (N_2679,N_2546,N_2596);
and U2680 (N_2680,N_2597,N_2534);
nand U2681 (N_2681,N_2568,N_2509);
or U2682 (N_2682,N_2565,N_2551);
or U2683 (N_2683,N_2569,N_2520);
or U2684 (N_2684,N_2580,N_2590);
nor U2685 (N_2685,N_2517,N_2570);
and U2686 (N_2686,N_2534,N_2555);
nor U2687 (N_2687,N_2558,N_2581);
and U2688 (N_2688,N_2563,N_2501);
nor U2689 (N_2689,N_2511,N_2508);
nor U2690 (N_2690,N_2537,N_2522);
nand U2691 (N_2691,N_2534,N_2537);
xor U2692 (N_2692,N_2558,N_2548);
and U2693 (N_2693,N_2587,N_2594);
or U2694 (N_2694,N_2531,N_2544);
nor U2695 (N_2695,N_2583,N_2570);
and U2696 (N_2696,N_2541,N_2587);
nor U2697 (N_2697,N_2579,N_2592);
or U2698 (N_2698,N_2583,N_2520);
nand U2699 (N_2699,N_2571,N_2555);
or U2700 (N_2700,N_2643,N_2653);
and U2701 (N_2701,N_2620,N_2609);
and U2702 (N_2702,N_2650,N_2663);
and U2703 (N_2703,N_2674,N_2625);
or U2704 (N_2704,N_2698,N_2681);
and U2705 (N_2705,N_2616,N_2676);
and U2706 (N_2706,N_2672,N_2668);
nor U2707 (N_2707,N_2659,N_2673);
nor U2708 (N_2708,N_2687,N_2656);
nor U2709 (N_2709,N_2636,N_2611);
and U2710 (N_2710,N_2604,N_2637);
nor U2711 (N_2711,N_2655,N_2610);
and U2712 (N_2712,N_2662,N_2683);
or U2713 (N_2713,N_2670,N_2621);
and U2714 (N_2714,N_2615,N_2608);
or U2715 (N_2715,N_2617,N_2646);
nand U2716 (N_2716,N_2622,N_2626);
or U2717 (N_2717,N_2657,N_2624);
or U2718 (N_2718,N_2614,N_2680);
nand U2719 (N_2719,N_2634,N_2660);
nor U2720 (N_2720,N_2664,N_2632);
and U2721 (N_2721,N_2684,N_2693);
and U2722 (N_2722,N_2629,N_2665);
nand U2723 (N_2723,N_2633,N_2623);
or U2724 (N_2724,N_2699,N_2627);
nor U2725 (N_2725,N_2640,N_2619);
nor U2726 (N_2726,N_2645,N_2658);
and U2727 (N_2727,N_2605,N_2631);
or U2728 (N_2728,N_2601,N_2677);
or U2729 (N_2729,N_2675,N_2661);
or U2730 (N_2730,N_2602,N_2613);
nand U2731 (N_2731,N_2692,N_2679);
nand U2732 (N_2732,N_2635,N_2651);
or U2733 (N_2733,N_2654,N_2689);
nor U2734 (N_2734,N_2638,N_2649);
or U2735 (N_2735,N_2686,N_2688);
and U2736 (N_2736,N_2666,N_2694);
or U2737 (N_2737,N_2682,N_2612);
and U2738 (N_2738,N_2606,N_2630);
nor U2739 (N_2739,N_2690,N_2642);
and U2740 (N_2740,N_2671,N_2691);
and U2741 (N_2741,N_2697,N_2600);
nor U2742 (N_2742,N_2685,N_2603);
and U2743 (N_2743,N_2647,N_2648);
nand U2744 (N_2744,N_2669,N_2667);
and U2745 (N_2745,N_2639,N_2695);
or U2746 (N_2746,N_2641,N_2607);
or U2747 (N_2747,N_2678,N_2644);
nor U2748 (N_2748,N_2652,N_2618);
nor U2749 (N_2749,N_2696,N_2628);
nand U2750 (N_2750,N_2638,N_2641);
and U2751 (N_2751,N_2693,N_2664);
and U2752 (N_2752,N_2636,N_2666);
nor U2753 (N_2753,N_2622,N_2694);
nand U2754 (N_2754,N_2687,N_2642);
and U2755 (N_2755,N_2683,N_2692);
nor U2756 (N_2756,N_2683,N_2632);
nand U2757 (N_2757,N_2669,N_2679);
nor U2758 (N_2758,N_2639,N_2605);
and U2759 (N_2759,N_2649,N_2629);
and U2760 (N_2760,N_2637,N_2676);
nand U2761 (N_2761,N_2682,N_2605);
or U2762 (N_2762,N_2628,N_2689);
and U2763 (N_2763,N_2617,N_2673);
and U2764 (N_2764,N_2666,N_2628);
nand U2765 (N_2765,N_2699,N_2670);
and U2766 (N_2766,N_2670,N_2643);
nor U2767 (N_2767,N_2624,N_2651);
nor U2768 (N_2768,N_2659,N_2687);
nand U2769 (N_2769,N_2658,N_2600);
or U2770 (N_2770,N_2635,N_2674);
xor U2771 (N_2771,N_2670,N_2606);
nor U2772 (N_2772,N_2622,N_2621);
or U2773 (N_2773,N_2620,N_2671);
nor U2774 (N_2774,N_2636,N_2606);
nor U2775 (N_2775,N_2675,N_2699);
and U2776 (N_2776,N_2646,N_2614);
nor U2777 (N_2777,N_2618,N_2614);
nor U2778 (N_2778,N_2683,N_2605);
nand U2779 (N_2779,N_2687,N_2650);
and U2780 (N_2780,N_2674,N_2667);
nand U2781 (N_2781,N_2676,N_2668);
nor U2782 (N_2782,N_2695,N_2677);
and U2783 (N_2783,N_2661,N_2609);
or U2784 (N_2784,N_2612,N_2653);
nor U2785 (N_2785,N_2645,N_2643);
nor U2786 (N_2786,N_2667,N_2637);
nor U2787 (N_2787,N_2619,N_2695);
nor U2788 (N_2788,N_2647,N_2606);
or U2789 (N_2789,N_2646,N_2622);
and U2790 (N_2790,N_2629,N_2646);
nand U2791 (N_2791,N_2671,N_2605);
and U2792 (N_2792,N_2688,N_2677);
or U2793 (N_2793,N_2647,N_2654);
and U2794 (N_2794,N_2634,N_2612);
and U2795 (N_2795,N_2672,N_2658);
and U2796 (N_2796,N_2689,N_2684);
nor U2797 (N_2797,N_2652,N_2690);
xor U2798 (N_2798,N_2686,N_2641);
nand U2799 (N_2799,N_2627,N_2647);
nor U2800 (N_2800,N_2714,N_2723);
or U2801 (N_2801,N_2739,N_2729);
and U2802 (N_2802,N_2716,N_2712);
and U2803 (N_2803,N_2749,N_2795);
or U2804 (N_2804,N_2721,N_2797);
and U2805 (N_2805,N_2762,N_2715);
and U2806 (N_2806,N_2759,N_2796);
and U2807 (N_2807,N_2746,N_2777);
nand U2808 (N_2808,N_2773,N_2700);
nor U2809 (N_2809,N_2748,N_2752);
and U2810 (N_2810,N_2707,N_2730);
or U2811 (N_2811,N_2760,N_2705);
nand U2812 (N_2812,N_2711,N_2744);
or U2813 (N_2813,N_2772,N_2787);
nor U2814 (N_2814,N_2740,N_2709);
or U2815 (N_2815,N_2734,N_2756);
or U2816 (N_2816,N_2780,N_2771);
and U2817 (N_2817,N_2754,N_2738);
and U2818 (N_2818,N_2733,N_2704);
nor U2819 (N_2819,N_2785,N_2783);
nand U2820 (N_2820,N_2793,N_2782);
and U2821 (N_2821,N_2718,N_2779);
nand U2822 (N_2822,N_2719,N_2727);
and U2823 (N_2823,N_2743,N_2732);
and U2824 (N_2824,N_2774,N_2728);
nor U2825 (N_2825,N_2725,N_2742);
or U2826 (N_2826,N_2717,N_2789);
and U2827 (N_2827,N_2781,N_2758);
and U2828 (N_2828,N_2726,N_2778);
xor U2829 (N_2829,N_2799,N_2794);
nand U2830 (N_2830,N_2706,N_2757);
and U2831 (N_2831,N_2790,N_2710);
nand U2832 (N_2832,N_2763,N_2765);
and U2833 (N_2833,N_2735,N_2753);
and U2834 (N_2834,N_2741,N_2702);
or U2835 (N_2835,N_2703,N_2770);
and U2836 (N_2836,N_2737,N_2768);
nor U2837 (N_2837,N_2755,N_2767);
or U2838 (N_2838,N_2708,N_2722);
nand U2839 (N_2839,N_2776,N_2764);
or U2840 (N_2840,N_2751,N_2775);
nor U2841 (N_2841,N_2750,N_2713);
nor U2842 (N_2842,N_2731,N_2724);
and U2843 (N_2843,N_2761,N_2745);
nor U2844 (N_2844,N_2747,N_2769);
nor U2845 (N_2845,N_2701,N_2788);
nand U2846 (N_2846,N_2786,N_2791);
nor U2847 (N_2847,N_2784,N_2736);
or U2848 (N_2848,N_2798,N_2720);
nor U2849 (N_2849,N_2766,N_2792);
nor U2850 (N_2850,N_2771,N_2795);
nand U2851 (N_2851,N_2710,N_2775);
and U2852 (N_2852,N_2710,N_2785);
or U2853 (N_2853,N_2703,N_2781);
and U2854 (N_2854,N_2752,N_2781);
or U2855 (N_2855,N_2790,N_2764);
nor U2856 (N_2856,N_2797,N_2743);
and U2857 (N_2857,N_2741,N_2780);
nand U2858 (N_2858,N_2709,N_2766);
nand U2859 (N_2859,N_2795,N_2748);
nand U2860 (N_2860,N_2717,N_2791);
or U2861 (N_2861,N_2723,N_2752);
and U2862 (N_2862,N_2712,N_2726);
or U2863 (N_2863,N_2781,N_2744);
nor U2864 (N_2864,N_2775,N_2798);
nor U2865 (N_2865,N_2770,N_2734);
and U2866 (N_2866,N_2716,N_2771);
nand U2867 (N_2867,N_2780,N_2764);
nand U2868 (N_2868,N_2731,N_2709);
nor U2869 (N_2869,N_2728,N_2776);
nor U2870 (N_2870,N_2765,N_2761);
nand U2871 (N_2871,N_2762,N_2725);
nor U2872 (N_2872,N_2725,N_2796);
nor U2873 (N_2873,N_2711,N_2736);
and U2874 (N_2874,N_2759,N_2784);
and U2875 (N_2875,N_2787,N_2719);
nand U2876 (N_2876,N_2727,N_2728);
and U2877 (N_2877,N_2740,N_2717);
or U2878 (N_2878,N_2716,N_2769);
nor U2879 (N_2879,N_2751,N_2710);
nand U2880 (N_2880,N_2799,N_2745);
nand U2881 (N_2881,N_2766,N_2706);
or U2882 (N_2882,N_2796,N_2779);
nand U2883 (N_2883,N_2784,N_2705);
and U2884 (N_2884,N_2736,N_2794);
nand U2885 (N_2885,N_2717,N_2734);
and U2886 (N_2886,N_2771,N_2728);
nand U2887 (N_2887,N_2718,N_2744);
and U2888 (N_2888,N_2745,N_2788);
or U2889 (N_2889,N_2784,N_2755);
and U2890 (N_2890,N_2701,N_2710);
nand U2891 (N_2891,N_2736,N_2739);
or U2892 (N_2892,N_2760,N_2736);
or U2893 (N_2893,N_2718,N_2773);
and U2894 (N_2894,N_2745,N_2736);
or U2895 (N_2895,N_2753,N_2705);
xnor U2896 (N_2896,N_2771,N_2787);
xor U2897 (N_2897,N_2720,N_2776);
nand U2898 (N_2898,N_2777,N_2702);
and U2899 (N_2899,N_2790,N_2783);
and U2900 (N_2900,N_2858,N_2899);
nand U2901 (N_2901,N_2801,N_2828);
nor U2902 (N_2902,N_2888,N_2823);
and U2903 (N_2903,N_2835,N_2873);
and U2904 (N_2904,N_2884,N_2876);
and U2905 (N_2905,N_2819,N_2879);
nor U2906 (N_2906,N_2824,N_2829);
nand U2907 (N_2907,N_2894,N_2870);
and U2908 (N_2908,N_2865,N_2874);
and U2909 (N_2909,N_2802,N_2882);
nand U2910 (N_2910,N_2843,N_2878);
xor U2911 (N_2911,N_2803,N_2834);
and U2912 (N_2912,N_2836,N_2827);
xor U2913 (N_2913,N_2848,N_2881);
and U2914 (N_2914,N_2825,N_2861);
nor U2915 (N_2915,N_2816,N_2862);
and U2916 (N_2916,N_2840,N_2859);
nor U2917 (N_2917,N_2847,N_2864);
nand U2918 (N_2918,N_2877,N_2849);
and U2919 (N_2919,N_2872,N_2892);
nand U2920 (N_2920,N_2813,N_2854);
xnor U2921 (N_2921,N_2885,N_2838);
or U2922 (N_2922,N_2866,N_2868);
nor U2923 (N_2923,N_2886,N_2889);
and U2924 (N_2924,N_2852,N_2810);
and U2925 (N_2925,N_2842,N_2815);
nand U2926 (N_2926,N_2821,N_2871);
or U2927 (N_2927,N_2818,N_2826);
nand U2928 (N_2928,N_2893,N_2806);
nand U2929 (N_2929,N_2833,N_2814);
and U2930 (N_2930,N_2841,N_2855);
nand U2931 (N_2931,N_2898,N_2822);
or U2932 (N_2932,N_2832,N_2896);
nor U2933 (N_2933,N_2867,N_2880);
nor U2934 (N_2934,N_2887,N_2839);
and U2935 (N_2935,N_2811,N_2807);
or U2936 (N_2936,N_2809,N_2897);
and U2937 (N_2937,N_2890,N_2820);
or U2938 (N_2938,N_2895,N_2812);
or U2939 (N_2939,N_2851,N_2845);
nand U2940 (N_2940,N_2856,N_2817);
nor U2941 (N_2941,N_2808,N_2805);
nor U2942 (N_2942,N_2863,N_2860);
nand U2943 (N_2943,N_2883,N_2857);
or U2944 (N_2944,N_2846,N_2804);
nand U2945 (N_2945,N_2891,N_2850);
nor U2946 (N_2946,N_2875,N_2831);
or U2947 (N_2947,N_2800,N_2844);
or U2948 (N_2948,N_2830,N_2853);
nor U2949 (N_2949,N_2837,N_2869);
or U2950 (N_2950,N_2865,N_2832);
and U2951 (N_2951,N_2819,N_2893);
nor U2952 (N_2952,N_2822,N_2892);
nor U2953 (N_2953,N_2844,N_2890);
or U2954 (N_2954,N_2873,N_2895);
nor U2955 (N_2955,N_2837,N_2800);
nand U2956 (N_2956,N_2869,N_2826);
and U2957 (N_2957,N_2895,N_2807);
and U2958 (N_2958,N_2816,N_2881);
nor U2959 (N_2959,N_2812,N_2889);
nand U2960 (N_2960,N_2873,N_2825);
or U2961 (N_2961,N_2814,N_2812);
and U2962 (N_2962,N_2824,N_2817);
nand U2963 (N_2963,N_2885,N_2898);
nor U2964 (N_2964,N_2887,N_2832);
or U2965 (N_2965,N_2848,N_2871);
and U2966 (N_2966,N_2829,N_2855);
nor U2967 (N_2967,N_2800,N_2885);
or U2968 (N_2968,N_2877,N_2866);
or U2969 (N_2969,N_2862,N_2809);
and U2970 (N_2970,N_2876,N_2826);
nor U2971 (N_2971,N_2808,N_2883);
or U2972 (N_2972,N_2854,N_2886);
nor U2973 (N_2973,N_2891,N_2857);
nor U2974 (N_2974,N_2895,N_2874);
or U2975 (N_2975,N_2833,N_2867);
nor U2976 (N_2976,N_2892,N_2817);
and U2977 (N_2977,N_2838,N_2828);
nand U2978 (N_2978,N_2893,N_2807);
nor U2979 (N_2979,N_2869,N_2839);
or U2980 (N_2980,N_2894,N_2831);
nor U2981 (N_2981,N_2853,N_2840);
or U2982 (N_2982,N_2813,N_2867);
nand U2983 (N_2983,N_2889,N_2870);
xnor U2984 (N_2984,N_2870,N_2884);
nand U2985 (N_2985,N_2831,N_2872);
or U2986 (N_2986,N_2846,N_2840);
and U2987 (N_2987,N_2891,N_2808);
and U2988 (N_2988,N_2877,N_2887);
nor U2989 (N_2989,N_2809,N_2874);
nor U2990 (N_2990,N_2830,N_2839);
nand U2991 (N_2991,N_2829,N_2853);
nand U2992 (N_2992,N_2810,N_2800);
nand U2993 (N_2993,N_2800,N_2865);
and U2994 (N_2994,N_2899,N_2849);
nand U2995 (N_2995,N_2876,N_2877);
nand U2996 (N_2996,N_2835,N_2839);
and U2997 (N_2997,N_2842,N_2807);
or U2998 (N_2998,N_2833,N_2826);
nor U2999 (N_2999,N_2859,N_2811);
nor UO_0 (O_0,N_2969,N_2936);
and UO_1 (O_1,N_2908,N_2945);
nand UO_2 (O_2,N_2998,N_2919);
and UO_3 (O_3,N_2978,N_2985);
xnor UO_4 (O_4,N_2902,N_2965);
or UO_5 (O_5,N_2983,N_2932);
or UO_6 (O_6,N_2967,N_2938);
nand UO_7 (O_7,N_2923,N_2929);
or UO_8 (O_8,N_2964,N_2909);
and UO_9 (O_9,N_2900,N_2982);
nor UO_10 (O_10,N_2995,N_2947);
and UO_11 (O_11,N_2941,N_2907);
nand UO_12 (O_12,N_2925,N_2970);
and UO_13 (O_13,N_2915,N_2974);
or UO_14 (O_14,N_2912,N_2956);
nand UO_15 (O_15,N_2904,N_2981);
or UO_16 (O_16,N_2901,N_2986);
nand UO_17 (O_17,N_2943,N_2950);
nand UO_18 (O_18,N_2952,N_2918);
nor UO_19 (O_19,N_2999,N_2922);
or UO_20 (O_20,N_2994,N_2931);
and UO_21 (O_21,N_2917,N_2975);
and UO_22 (O_22,N_2903,N_2976);
nor UO_23 (O_23,N_2988,N_2959);
or UO_24 (O_24,N_2928,N_2963);
nor UO_25 (O_25,N_2989,N_2991);
nand UO_26 (O_26,N_2926,N_2997);
and UO_27 (O_27,N_2937,N_2955);
nand UO_28 (O_28,N_2993,N_2992);
nor UO_29 (O_29,N_2961,N_2953);
and UO_30 (O_30,N_2984,N_2939);
nor UO_31 (O_31,N_2916,N_2971);
or UO_32 (O_32,N_2949,N_2973);
nor UO_33 (O_33,N_2948,N_2933);
and UO_34 (O_34,N_2987,N_2951);
nand UO_35 (O_35,N_2966,N_2972);
and UO_36 (O_36,N_2911,N_2957);
or UO_37 (O_37,N_2944,N_2960);
nor UO_38 (O_38,N_2921,N_2920);
nand UO_39 (O_39,N_2979,N_2924);
or UO_40 (O_40,N_2996,N_2914);
nor UO_41 (O_41,N_2930,N_2927);
nand UO_42 (O_42,N_2980,N_2910);
and UO_43 (O_43,N_2962,N_2935);
nand UO_44 (O_44,N_2906,N_2946);
and UO_45 (O_45,N_2905,N_2942);
nand UO_46 (O_46,N_2990,N_2958);
nor UO_47 (O_47,N_2913,N_2954);
or UO_48 (O_48,N_2934,N_2968);
or UO_49 (O_49,N_2940,N_2977);
and UO_50 (O_50,N_2968,N_2960);
and UO_51 (O_51,N_2949,N_2998);
and UO_52 (O_52,N_2981,N_2968);
nor UO_53 (O_53,N_2951,N_2930);
and UO_54 (O_54,N_2941,N_2951);
or UO_55 (O_55,N_2980,N_2909);
or UO_56 (O_56,N_2945,N_2900);
nand UO_57 (O_57,N_2993,N_2973);
and UO_58 (O_58,N_2937,N_2929);
or UO_59 (O_59,N_2935,N_2969);
and UO_60 (O_60,N_2922,N_2951);
nor UO_61 (O_61,N_2991,N_2965);
nand UO_62 (O_62,N_2964,N_2985);
or UO_63 (O_63,N_2901,N_2943);
or UO_64 (O_64,N_2994,N_2943);
nor UO_65 (O_65,N_2969,N_2911);
nand UO_66 (O_66,N_2952,N_2965);
or UO_67 (O_67,N_2985,N_2906);
nand UO_68 (O_68,N_2925,N_2900);
nor UO_69 (O_69,N_2957,N_2936);
or UO_70 (O_70,N_2911,N_2930);
nor UO_71 (O_71,N_2953,N_2965);
nand UO_72 (O_72,N_2984,N_2964);
or UO_73 (O_73,N_2997,N_2952);
or UO_74 (O_74,N_2921,N_2909);
nor UO_75 (O_75,N_2961,N_2952);
nand UO_76 (O_76,N_2955,N_2951);
nand UO_77 (O_77,N_2929,N_2936);
nor UO_78 (O_78,N_2964,N_2911);
or UO_79 (O_79,N_2999,N_2924);
and UO_80 (O_80,N_2999,N_2948);
and UO_81 (O_81,N_2944,N_2969);
or UO_82 (O_82,N_2979,N_2968);
and UO_83 (O_83,N_2978,N_2999);
nand UO_84 (O_84,N_2922,N_2984);
nor UO_85 (O_85,N_2995,N_2954);
nand UO_86 (O_86,N_2986,N_2956);
nand UO_87 (O_87,N_2906,N_2943);
or UO_88 (O_88,N_2939,N_2925);
and UO_89 (O_89,N_2981,N_2940);
and UO_90 (O_90,N_2997,N_2996);
nand UO_91 (O_91,N_2900,N_2938);
and UO_92 (O_92,N_2942,N_2952);
nand UO_93 (O_93,N_2938,N_2974);
or UO_94 (O_94,N_2913,N_2949);
nand UO_95 (O_95,N_2981,N_2938);
nor UO_96 (O_96,N_2927,N_2963);
or UO_97 (O_97,N_2939,N_2903);
nand UO_98 (O_98,N_2939,N_2904);
and UO_99 (O_99,N_2922,N_2938);
or UO_100 (O_100,N_2945,N_2957);
nand UO_101 (O_101,N_2996,N_2954);
and UO_102 (O_102,N_2938,N_2924);
nor UO_103 (O_103,N_2901,N_2976);
or UO_104 (O_104,N_2958,N_2944);
nand UO_105 (O_105,N_2956,N_2918);
nand UO_106 (O_106,N_2990,N_2913);
nor UO_107 (O_107,N_2933,N_2932);
and UO_108 (O_108,N_2930,N_2924);
nand UO_109 (O_109,N_2936,N_2914);
or UO_110 (O_110,N_2958,N_2978);
nand UO_111 (O_111,N_2951,N_2989);
or UO_112 (O_112,N_2946,N_2901);
nand UO_113 (O_113,N_2955,N_2967);
and UO_114 (O_114,N_2926,N_2933);
nor UO_115 (O_115,N_2912,N_2948);
nor UO_116 (O_116,N_2961,N_2975);
nand UO_117 (O_117,N_2969,N_2932);
or UO_118 (O_118,N_2915,N_2913);
or UO_119 (O_119,N_2937,N_2922);
nor UO_120 (O_120,N_2904,N_2921);
nand UO_121 (O_121,N_2994,N_2989);
nand UO_122 (O_122,N_2912,N_2941);
or UO_123 (O_123,N_2973,N_2957);
nor UO_124 (O_124,N_2980,N_2942);
nand UO_125 (O_125,N_2926,N_2978);
or UO_126 (O_126,N_2961,N_2978);
nand UO_127 (O_127,N_2946,N_2949);
and UO_128 (O_128,N_2956,N_2925);
xnor UO_129 (O_129,N_2985,N_2916);
nand UO_130 (O_130,N_2962,N_2964);
and UO_131 (O_131,N_2920,N_2942);
nor UO_132 (O_132,N_2914,N_2909);
nor UO_133 (O_133,N_2993,N_2999);
nand UO_134 (O_134,N_2903,N_2900);
nor UO_135 (O_135,N_2952,N_2978);
and UO_136 (O_136,N_2928,N_2930);
or UO_137 (O_137,N_2964,N_2976);
nand UO_138 (O_138,N_2998,N_2961);
or UO_139 (O_139,N_2954,N_2961);
or UO_140 (O_140,N_2973,N_2983);
nand UO_141 (O_141,N_2969,N_2919);
nand UO_142 (O_142,N_2994,N_2961);
and UO_143 (O_143,N_2997,N_2964);
or UO_144 (O_144,N_2944,N_2950);
or UO_145 (O_145,N_2971,N_2953);
nand UO_146 (O_146,N_2927,N_2957);
or UO_147 (O_147,N_2916,N_2926);
xnor UO_148 (O_148,N_2963,N_2932);
nand UO_149 (O_149,N_2970,N_2978);
and UO_150 (O_150,N_2995,N_2913);
nand UO_151 (O_151,N_2960,N_2934);
or UO_152 (O_152,N_2987,N_2986);
or UO_153 (O_153,N_2995,N_2965);
and UO_154 (O_154,N_2925,N_2923);
and UO_155 (O_155,N_2952,N_2928);
and UO_156 (O_156,N_2912,N_2954);
nand UO_157 (O_157,N_2972,N_2946);
nand UO_158 (O_158,N_2921,N_2924);
xnor UO_159 (O_159,N_2926,N_2923);
and UO_160 (O_160,N_2970,N_2952);
nor UO_161 (O_161,N_2921,N_2965);
nor UO_162 (O_162,N_2933,N_2970);
and UO_163 (O_163,N_2962,N_2937);
nand UO_164 (O_164,N_2942,N_2918);
and UO_165 (O_165,N_2928,N_2995);
nand UO_166 (O_166,N_2977,N_2917);
and UO_167 (O_167,N_2994,N_2946);
nor UO_168 (O_168,N_2933,N_2950);
or UO_169 (O_169,N_2915,N_2937);
and UO_170 (O_170,N_2931,N_2963);
nor UO_171 (O_171,N_2977,N_2952);
nor UO_172 (O_172,N_2944,N_2913);
and UO_173 (O_173,N_2967,N_2984);
or UO_174 (O_174,N_2938,N_2949);
and UO_175 (O_175,N_2962,N_2976);
nand UO_176 (O_176,N_2986,N_2942);
and UO_177 (O_177,N_2999,N_2960);
nor UO_178 (O_178,N_2920,N_2977);
or UO_179 (O_179,N_2935,N_2932);
nand UO_180 (O_180,N_2989,N_2910);
nor UO_181 (O_181,N_2963,N_2914);
nor UO_182 (O_182,N_2902,N_2991);
xnor UO_183 (O_183,N_2943,N_2937);
nand UO_184 (O_184,N_2903,N_2993);
and UO_185 (O_185,N_2999,N_2968);
and UO_186 (O_186,N_2924,N_2962);
or UO_187 (O_187,N_2998,N_2921);
or UO_188 (O_188,N_2903,N_2917);
nand UO_189 (O_189,N_2916,N_2941);
nor UO_190 (O_190,N_2940,N_2907);
or UO_191 (O_191,N_2981,N_2931);
nand UO_192 (O_192,N_2903,N_2906);
nand UO_193 (O_193,N_2980,N_2985);
or UO_194 (O_194,N_2981,N_2987);
or UO_195 (O_195,N_2992,N_2929);
nand UO_196 (O_196,N_2964,N_2965);
and UO_197 (O_197,N_2936,N_2951);
and UO_198 (O_198,N_2936,N_2984);
nor UO_199 (O_199,N_2993,N_2921);
and UO_200 (O_200,N_2922,N_2973);
nor UO_201 (O_201,N_2977,N_2950);
or UO_202 (O_202,N_2954,N_2916);
nor UO_203 (O_203,N_2988,N_2941);
and UO_204 (O_204,N_2928,N_2954);
nor UO_205 (O_205,N_2943,N_2992);
or UO_206 (O_206,N_2909,N_2997);
nand UO_207 (O_207,N_2988,N_2924);
nand UO_208 (O_208,N_2939,N_2924);
or UO_209 (O_209,N_2918,N_2902);
or UO_210 (O_210,N_2912,N_2979);
or UO_211 (O_211,N_2955,N_2954);
and UO_212 (O_212,N_2975,N_2947);
nand UO_213 (O_213,N_2949,N_2982);
nor UO_214 (O_214,N_2983,N_2997);
nand UO_215 (O_215,N_2954,N_2963);
nand UO_216 (O_216,N_2941,N_2930);
or UO_217 (O_217,N_2980,N_2984);
and UO_218 (O_218,N_2935,N_2912);
or UO_219 (O_219,N_2983,N_2982);
nand UO_220 (O_220,N_2904,N_2993);
xor UO_221 (O_221,N_2940,N_2965);
or UO_222 (O_222,N_2942,N_2922);
nand UO_223 (O_223,N_2904,N_2932);
or UO_224 (O_224,N_2968,N_2989);
and UO_225 (O_225,N_2923,N_2984);
or UO_226 (O_226,N_2985,N_2974);
and UO_227 (O_227,N_2995,N_2978);
or UO_228 (O_228,N_2929,N_2909);
or UO_229 (O_229,N_2966,N_2916);
nor UO_230 (O_230,N_2935,N_2948);
nor UO_231 (O_231,N_2927,N_2969);
nand UO_232 (O_232,N_2998,N_2955);
nand UO_233 (O_233,N_2956,N_2931);
nor UO_234 (O_234,N_2960,N_2940);
and UO_235 (O_235,N_2950,N_2903);
nand UO_236 (O_236,N_2997,N_2920);
nor UO_237 (O_237,N_2931,N_2923);
nand UO_238 (O_238,N_2946,N_2985);
nor UO_239 (O_239,N_2958,N_2966);
nand UO_240 (O_240,N_2952,N_2998);
or UO_241 (O_241,N_2997,N_2991);
nor UO_242 (O_242,N_2962,N_2956);
nand UO_243 (O_243,N_2944,N_2909);
xnor UO_244 (O_244,N_2904,N_2990);
nor UO_245 (O_245,N_2991,N_2933);
or UO_246 (O_246,N_2977,N_2985);
and UO_247 (O_247,N_2971,N_2956);
nand UO_248 (O_248,N_2985,N_2927);
or UO_249 (O_249,N_2926,N_2959);
and UO_250 (O_250,N_2991,N_2983);
and UO_251 (O_251,N_2907,N_2942);
nor UO_252 (O_252,N_2935,N_2992);
or UO_253 (O_253,N_2926,N_2910);
and UO_254 (O_254,N_2958,N_2979);
nor UO_255 (O_255,N_2915,N_2924);
nand UO_256 (O_256,N_2964,N_2914);
nand UO_257 (O_257,N_2955,N_2910);
nor UO_258 (O_258,N_2916,N_2927);
and UO_259 (O_259,N_2966,N_2921);
and UO_260 (O_260,N_2924,N_2989);
or UO_261 (O_261,N_2922,N_2931);
xor UO_262 (O_262,N_2923,N_2965);
nor UO_263 (O_263,N_2966,N_2940);
and UO_264 (O_264,N_2925,N_2943);
and UO_265 (O_265,N_2978,N_2992);
nor UO_266 (O_266,N_2906,N_2993);
nor UO_267 (O_267,N_2969,N_2989);
and UO_268 (O_268,N_2925,N_2901);
or UO_269 (O_269,N_2923,N_2971);
nand UO_270 (O_270,N_2964,N_2989);
or UO_271 (O_271,N_2954,N_2970);
or UO_272 (O_272,N_2907,N_2996);
or UO_273 (O_273,N_2903,N_2965);
nand UO_274 (O_274,N_2957,N_2976);
nor UO_275 (O_275,N_2929,N_2935);
nor UO_276 (O_276,N_2923,N_2934);
nor UO_277 (O_277,N_2914,N_2934);
or UO_278 (O_278,N_2971,N_2907);
and UO_279 (O_279,N_2927,N_2929);
or UO_280 (O_280,N_2917,N_2957);
and UO_281 (O_281,N_2939,N_2910);
nor UO_282 (O_282,N_2945,N_2928);
nand UO_283 (O_283,N_2920,N_2981);
nand UO_284 (O_284,N_2918,N_2924);
nor UO_285 (O_285,N_2928,N_2910);
or UO_286 (O_286,N_2910,N_2945);
and UO_287 (O_287,N_2962,N_2949);
or UO_288 (O_288,N_2933,N_2915);
nand UO_289 (O_289,N_2986,N_2945);
nor UO_290 (O_290,N_2966,N_2997);
nor UO_291 (O_291,N_2972,N_2982);
and UO_292 (O_292,N_2915,N_2998);
xor UO_293 (O_293,N_2922,N_2991);
xnor UO_294 (O_294,N_2905,N_2935);
or UO_295 (O_295,N_2950,N_2931);
nor UO_296 (O_296,N_2985,N_2932);
or UO_297 (O_297,N_2918,N_2990);
nand UO_298 (O_298,N_2998,N_2937);
and UO_299 (O_299,N_2944,N_2946);
or UO_300 (O_300,N_2914,N_2942);
and UO_301 (O_301,N_2940,N_2932);
nor UO_302 (O_302,N_2986,N_2973);
and UO_303 (O_303,N_2939,N_2901);
nand UO_304 (O_304,N_2974,N_2998);
nor UO_305 (O_305,N_2909,N_2989);
or UO_306 (O_306,N_2987,N_2982);
and UO_307 (O_307,N_2928,N_2973);
and UO_308 (O_308,N_2903,N_2926);
nor UO_309 (O_309,N_2925,N_2998);
nand UO_310 (O_310,N_2920,N_2937);
or UO_311 (O_311,N_2954,N_2978);
nor UO_312 (O_312,N_2983,N_2907);
nand UO_313 (O_313,N_2982,N_2933);
nor UO_314 (O_314,N_2974,N_2986);
nand UO_315 (O_315,N_2900,N_2936);
nor UO_316 (O_316,N_2935,N_2911);
and UO_317 (O_317,N_2907,N_2937);
nand UO_318 (O_318,N_2984,N_2930);
nor UO_319 (O_319,N_2951,N_2915);
nor UO_320 (O_320,N_2933,N_2937);
nor UO_321 (O_321,N_2943,N_2905);
or UO_322 (O_322,N_2976,N_2954);
and UO_323 (O_323,N_2936,N_2912);
or UO_324 (O_324,N_2919,N_2980);
or UO_325 (O_325,N_2947,N_2928);
nor UO_326 (O_326,N_2961,N_2976);
or UO_327 (O_327,N_2964,N_2991);
nand UO_328 (O_328,N_2982,N_2921);
and UO_329 (O_329,N_2992,N_2946);
nand UO_330 (O_330,N_2932,N_2988);
or UO_331 (O_331,N_2950,N_2930);
and UO_332 (O_332,N_2956,N_2945);
nor UO_333 (O_333,N_2967,N_2978);
or UO_334 (O_334,N_2988,N_2929);
nor UO_335 (O_335,N_2957,N_2974);
xnor UO_336 (O_336,N_2969,N_2926);
or UO_337 (O_337,N_2988,N_2911);
or UO_338 (O_338,N_2961,N_2980);
nor UO_339 (O_339,N_2924,N_2954);
nand UO_340 (O_340,N_2912,N_2981);
and UO_341 (O_341,N_2986,N_2967);
and UO_342 (O_342,N_2905,N_2996);
nand UO_343 (O_343,N_2997,N_2904);
and UO_344 (O_344,N_2961,N_2914);
or UO_345 (O_345,N_2999,N_2975);
xnor UO_346 (O_346,N_2918,N_2981);
nor UO_347 (O_347,N_2907,N_2946);
nor UO_348 (O_348,N_2988,N_2960);
nand UO_349 (O_349,N_2974,N_2926);
and UO_350 (O_350,N_2925,N_2960);
and UO_351 (O_351,N_2913,N_2910);
or UO_352 (O_352,N_2993,N_2971);
nor UO_353 (O_353,N_2949,N_2956);
and UO_354 (O_354,N_2986,N_2991);
and UO_355 (O_355,N_2993,N_2926);
nand UO_356 (O_356,N_2900,N_2960);
and UO_357 (O_357,N_2972,N_2916);
nand UO_358 (O_358,N_2992,N_2934);
and UO_359 (O_359,N_2976,N_2906);
nor UO_360 (O_360,N_2986,N_2931);
nand UO_361 (O_361,N_2954,N_2907);
nor UO_362 (O_362,N_2987,N_2992);
and UO_363 (O_363,N_2946,N_2922);
and UO_364 (O_364,N_2968,N_2909);
or UO_365 (O_365,N_2960,N_2939);
nand UO_366 (O_366,N_2902,N_2982);
nor UO_367 (O_367,N_2904,N_2980);
nor UO_368 (O_368,N_2955,N_2928);
nand UO_369 (O_369,N_2935,N_2900);
and UO_370 (O_370,N_2901,N_2929);
xor UO_371 (O_371,N_2947,N_2934);
and UO_372 (O_372,N_2947,N_2998);
nand UO_373 (O_373,N_2911,N_2934);
or UO_374 (O_374,N_2905,N_2973);
nand UO_375 (O_375,N_2935,N_2993);
nand UO_376 (O_376,N_2990,N_2924);
or UO_377 (O_377,N_2909,N_2971);
or UO_378 (O_378,N_2992,N_2953);
and UO_379 (O_379,N_2922,N_2976);
nand UO_380 (O_380,N_2967,N_2995);
nor UO_381 (O_381,N_2987,N_2947);
xnor UO_382 (O_382,N_2906,N_2930);
or UO_383 (O_383,N_2921,N_2951);
nand UO_384 (O_384,N_2906,N_2952);
and UO_385 (O_385,N_2970,N_2941);
nand UO_386 (O_386,N_2977,N_2986);
nand UO_387 (O_387,N_2909,N_2961);
and UO_388 (O_388,N_2925,N_2988);
nor UO_389 (O_389,N_2932,N_2972);
or UO_390 (O_390,N_2994,N_2920);
nor UO_391 (O_391,N_2993,N_2990);
nor UO_392 (O_392,N_2917,N_2938);
nand UO_393 (O_393,N_2941,N_2905);
or UO_394 (O_394,N_2998,N_2927);
nand UO_395 (O_395,N_2964,N_2906);
nand UO_396 (O_396,N_2933,N_2978);
nor UO_397 (O_397,N_2945,N_2950);
nor UO_398 (O_398,N_2932,N_2966);
or UO_399 (O_399,N_2982,N_2945);
nand UO_400 (O_400,N_2924,N_2970);
or UO_401 (O_401,N_2922,N_2987);
nand UO_402 (O_402,N_2915,N_2942);
and UO_403 (O_403,N_2994,N_2964);
nand UO_404 (O_404,N_2909,N_2928);
nor UO_405 (O_405,N_2902,N_2932);
or UO_406 (O_406,N_2937,N_2935);
nor UO_407 (O_407,N_2926,N_2983);
and UO_408 (O_408,N_2959,N_2965);
nor UO_409 (O_409,N_2943,N_2910);
and UO_410 (O_410,N_2952,N_2959);
nand UO_411 (O_411,N_2975,N_2985);
nand UO_412 (O_412,N_2933,N_2962);
or UO_413 (O_413,N_2986,N_2935);
and UO_414 (O_414,N_2983,N_2920);
nand UO_415 (O_415,N_2940,N_2998);
and UO_416 (O_416,N_2975,N_2969);
xor UO_417 (O_417,N_2951,N_2953);
and UO_418 (O_418,N_2972,N_2987);
nor UO_419 (O_419,N_2930,N_2905);
nand UO_420 (O_420,N_2936,N_2910);
nor UO_421 (O_421,N_2924,N_2953);
nor UO_422 (O_422,N_2920,N_2905);
nor UO_423 (O_423,N_2966,N_2934);
nand UO_424 (O_424,N_2968,N_2994);
nor UO_425 (O_425,N_2974,N_2956);
nand UO_426 (O_426,N_2959,N_2971);
and UO_427 (O_427,N_2909,N_2970);
nand UO_428 (O_428,N_2962,N_2910);
nor UO_429 (O_429,N_2982,N_2971);
and UO_430 (O_430,N_2928,N_2904);
or UO_431 (O_431,N_2962,N_2930);
or UO_432 (O_432,N_2945,N_2924);
or UO_433 (O_433,N_2950,N_2927);
nor UO_434 (O_434,N_2965,N_2922);
and UO_435 (O_435,N_2988,N_2970);
nor UO_436 (O_436,N_2906,N_2919);
nand UO_437 (O_437,N_2975,N_2981);
or UO_438 (O_438,N_2947,N_2993);
or UO_439 (O_439,N_2970,N_2945);
nand UO_440 (O_440,N_2922,N_2961);
nand UO_441 (O_441,N_2982,N_2939);
or UO_442 (O_442,N_2967,N_2908);
nor UO_443 (O_443,N_2942,N_2991);
and UO_444 (O_444,N_2900,N_2970);
nand UO_445 (O_445,N_2947,N_2923);
xnor UO_446 (O_446,N_2912,N_2908);
or UO_447 (O_447,N_2972,N_2964);
nor UO_448 (O_448,N_2933,N_2949);
nor UO_449 (O_449,N_2961,N_2991);
nand UO_450 (O_450,N_2987,N_2974);
and UO_451 (O_451,N_2960,N_2917);
and UO_452 (O_452,N_2966,N_2974);
and UO_453 (O_453,N_2918,N_2919);
or UO_454 (O_454,N_2919,N_2952);
or UO_455 (O_455,N_2910,N_2978);
nand UO_456 (O_456,N_2971,N_2974);
nor UO_457 (O_457,N_2902,N_2997);
nor UO_458 (O_458,N_2949,N_2942);
and UO_459 (O_459,N_2900,N_2992);
nor UO_460 (O_460,N_2913,N_2901);
nor UO_461 (O_461,N_2915,N_2902);
nand UO_462 (O_462,N_2935,N_2990);
or UO_463 (O_463,N_2916,N_2955);
and UO_464 (O_464,N_2934,N_2952);
nand UO_465 (O_465,N_2987,N_2904);
nand UO_466 (O_466,N_2900,N_2934);
nor UO_467 (O_467,N_2983,N_2992);
or UO_468 (O_468,N_2943,N_2931);
nor UO_469 (O_469,N_2978,N_2984);
or UO_470 (O_470,N_2994,N_2963);
or UO_471 (O_471,N_2937,N_2987);
nand UO_472 (O_472,N_2998,N_2953);
nand UO_473 (O_473,N_2999,N_2903);
nor UO_474 (O_474,N_2948,N_2969);
or UO_475 (O_475,N_2915,N_2922);
nor UO_476 (O_476,N_2979,N_2928);
xor UO_477 (O_477,N_2910,N_2958);
or UO_478 (O_478,N_2964,N_2903);
and UO_479 (O_479,N_2936,N_2959);
and UO_480 (O_480,N_2924,N_2920);
nand UO_481 (O_481,N_2943,N_2920);
nand UO_482 (O_482,N_2901,N_2930);
nor UO_483 (O_483,N_2923,N_2939);
nand UO_484 (O_484,N_2913,N_2919);
and UO_485 (O_485,N_2977,N_2964);
nand UO_486 (O_486,N_2969,N_2922);
nor UO_487 (O_487,N_2952,N_2966);
and UO_488 (O_488,N_2947,N_2990);
and UO_489 (O_489,N_2971,N_2906);
nand UO_490 (O_490,N_2985,N_2957);
nand UO_491 (O_491,N_2912,N_2930);
nand UO_492 (O_492,N_2973,N_2981);
or UO_493 (O_493,N_2971,N_2903);
nor UO_494 (O_494,N_2929,N_2999);
and UO_495 (O_495,N_2906,N_2941);
and UO_496 (O_496,N_2991,N_2921);
and UO_497 (O_497,N_2962,N_2934);
nor UO_498 (O_498,N_2903,N_2983);
nand UO_499 (O_499,N_2930,N_2989);
endmodule