module basic_500_3000_500_15_levels_10xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_419,In_447);
or U1 (N_1,In_73,In_369);
xnor U2 (N_2,In_8,In_498);
xor U3 (N_3,In_344,In_475);
nand U4 (N_4,In_381,In_249);
xnor U5 (N_5,In_286,In_185);
nor U6 (N_6,In_218,In_64);
nand U7 (N_7,In_171,In_164);
xor U8 (N_8,In_352,In_347);
and U9 (N_9,In_413,In_220);
or U10 (N_10,In_148,In_44);
xnor U11 (N_11,In_410,In_400);
and U12 (N_12,In_281,In_244);
nor U13 (N_13,In_277,In_82);
nand U14 (N_14,In_407,In_319);
or U15 (N_15,In_366,In_191);
nand U16 (N_16,In_241,In_97);
nand U17 (N_17,In_160,In_259);
nor U18 (N_18,In_140,In_132);
xnor U19 (N_19,In_386,In_485);
nor U20 (N_20,In_7,In_91);
nor U21 (N_21,In_405,In_494);
xnor U22 (N_22,In_284,In_60);
and U23 (N_23,In_77,In_204);
xnor U24 (N_24,In_302,In_263);
xor U25 (N_25,In_264,In_9);
and U26 (N_26,In_415,In_179);
or U27 (N_27,In_463,In_349);
or U28 (N_28,In_374,In_52);
nor U29 (N_29,In_247,In_432);
or U30 (N_30,In_20,In_226);
nor U31 (N_31,In_10,In_280);
nor U32 (N_32,In_454,In_106);
nand U33 (N_33,In_130,In_112);
or U34 (N_34,In_190,In_465);
and U35 (N_35,In_385,In_476);
nand U36 (N_36,In_467,In_293);
nor U37 (N_37,In_0,In_285);
nand U38 (N_38,In_1,In_239);
xnor U39 (N_39,In_201,In_92);
or U40 (N_40,In_438,In_43);
xnor U41 (N_41,In_442,In_208);
nand U42 (N_42,In_493,In_471);
and U43 (N_43,In_83,In_236);
nor U44 (N_44,In_240,In_306);
or U45 (N_45,In_428,In_154);
nand U46 (N_46,In_327,In_2);
or U47 (N_47,In_159,In_150);
xnor U48 (N_48,In_417,In_170);
and U49 (N_49,In_448,In_416);
xnor U50 (N_50,In_359,In_304);
nor U51 (N_51,In_300,In_470);
nand U52 (N_52,In_368,In_224);
or U53 (N_53,In_50,In_440);
nand U54 (N_54,In_151,In_118);
xor U55 (N_55,In_245,In_363);
nor U56 (N_56,In_328,In_392);
or U57 (N_57,In_353,In_215);
and U58 (N_58,In_375,In_153);
or U59 (N_59,In_488,In_315);
or U60 (N_60,In_129,In_325);
and U61 (N_61,In_358,In_174);
or U62 (N_62,In_289,In_48);
xor U63 (N_63,In_422,In_88);
or U64 (N_64,In_453,In_290);
xor U65 (N_65,In_287,In_324);
nor U66 (N_66,In_279,In_98);
and U67 (N_67,In_477,In_131);
xnor U68 (N_68,In_212,In_68);
and U69 (N_69,In_231,In_305);
or U70 (N_70,In_162,In_182);
or U71 (N_71,In_181,In_25);
nor U72 (N_72,In_458,In_108);
nor U73 (N_73,In_340,In_96);
nor U74 (N_74,In_398,In_312);
and U75 (N_75,In_156,In_478);
and U76 (N_76,In_188,In_23);
nor U77 (N_77,In_404,In_283);
nor U78 (N_78,In_409,In_371);
nand U79 (N_79,In_322,In_210);
nand U80 (N_80,In_85,In_394);
or U81 (N_81,In_391,In_141);
and U82 (N_82,In_142,In_298);
xor U83 (N_83,In_49,In_147);
nand U84 (N_84,In_46,In_89);
xor U85 (N_85,In_313,In_21);
or U86 (N_86,In_261,In_446);
or U87 (N_87,In_459,In_180);
xor U88 (N_88,In_119,In_127);
xor U89 (N_89,In_137,In_445);
nand U90 (N_90,In_491,In_403);
nor U91 (N_91,In_176,In_354);
and U92 (N_92,In_42,In_5);
nand U93 (N_93,In_219,In_361);
nor U94 (N_94,In_152,In_111);
xor U95 (N_95,In_232,In_32);
nor U96 (N_96,In_139,In_317);
and U97 (N_97,In_243,In_155);
and U98 (N_98,In_230,In_225);
or U99 (N_99,In_86,In_124);
or U100 (N_100,In_267,In_272);
xnor U101 (N_101,In_296,In_449);
xor U102 (N_102,In_310,In_339);
nor U103 (N_103,In_84,In_166);
or U104 (N_104,In_307,In_376);
nor U105 (N_105,In_406,In_135);
nand U106 (N_106,In_408,In_474);
and U107 (N_107,In_299,In_211);
nor U108 (N_108,In_456,In_58);
and U109 (N_109,In_496,In_274);
xnor U110 (N_110,In_341,In_37);
nor U111 (N_111,In_33,In_297);
xor U112 (N_112,In_79,In_273);
and U113 (N_113,In_499,In_269);
nand U114 (N_114,In_214,In_81);
nor U115 (N_115,In_402,In_158);
nand U116 (N_116,In_168,In_246);
nand U117 (N_117,In_431,In_275);
xnor U118 (N_118,In_288,In_87);
nor U119 (N_119,In_489,In_24);
nor U120 (N_120,In_198,In_426);
nand U121 (N_121,In_452,In_401);
nand U122 (N_122,In_175,In_423);
xnor U123 (N_123,In_40,In_473);
or U124 (N_124,In_104,In_378);
and U125 (N_125,In_26,In_45);
and U126 (N_126,In_462,In_16);
nor U127 (N_127,In_38,In_479);
nand U128 (N_128,In_451,In_66);
nand U129 (N_129,In_303,In_250);
and U130 (N_130,In_100,In_65);
and U131 (N_131,In_427,In_17);
nand U132 (N_132,In_257,In_469);
nor U133 (N_133,In_433,In_357);
or U134 (N_134,In_80,In_332);
xor U135 (N_135,In_12,In_348);
xnor U136 (N_136,In_107,In_487);
nand U137 (N_137,In_457,In_194);
nand U138 (N_138,In_429,In_276);
nor U139 (N_139,In_480,In_123);
nand U140 (N_140,In_377,In_125);
nand U141 (N_141,In_292,In_260);
or U142 (N_142,In_146,In_439);
nor U143 (N_143,In_425,In_157);
xnor U144 (N_144,In_63,In_203);
xor U145 (N_145,In_389,In_387);
nor U146 (N_146,In_196,In_268);
xor U147 (N_147,In_183,In_242);
or U148 (N_148,In_418,In_238);
and U149 (N_149,In_78,In_57);
nand U150 (N_150,In_109,In_390);
xnor U151 (N_151,In_397,In_128);
xor U152 (N_152,In_53,In_364);
nand U153 (N_153,In_253,In_421);
nand U154 (N_154,In_193,In_435);
or U155 (N_155,In_56,In_6);
xnor U156 (N_156,In_169,In_94);
and U157 (N_157,In_138,In_136);
nor U158 (N_158,In_420,In_436);
and U159 (N_159,In_497,In_481);
xnor U160 (N_160,In_309,In_346);
xor U161 (N_161,In_365,In_110);
nand U162 (N_162,In_206,In_270);
xor U163 (N_163,In_321,In_103);
xnor U164 (N_164,In_216,In_116);
nand U165 (N_165,In_223,In_76);
nand U166 (N_166,In_337,In_460);
or U167 (N_167,In_30,In_258);
nand U168 (N_168,In_101,In_102);
and U169 (N_169,In_330,In_39);
and U170 (N_170,In_149,In_75);
xor U171 (N_171,In_202,In_184);
nand U172 (N_172,In_70,In_134);
nor U173 (N_173,In_115,In_172);
and U174 (N_174,In_343,In_372);
nand U175 (N_175,In_27,In_29);
nor U176 (N_176,In_165,In_3);
nor U177 (N_177,In_120,In_11);
and U178 (N_178,In_61,In_388);
or U179 (N_179,In_14,In_59);
nor U180 (N_180,In_373,In_338);
xor U181 (N_181,In_395,In_237);
xnor U182 (N_182,In_67,In_495);
nor U183 (N_183,In_144,In_199);
or U184 (N_184,In_320,In_483);
xnor U185 (N_185,In_47,In_486);
nand U186 (N_186,In_444,In_200);
or U187 (N_187,In_318,In_329);
or U188 (N_188,In_173,In_351);
nand U189 (N_189,In_424,In_209);
nand U190 (N_190,In_95,In_314);
or U191 (N_191,In_468,In_187);
and U192 (N_192,In_221,In_163);
or U193 (N_193,In_19,In_31);
and U194 (N_194,In_434,In_331);
or U195 (N_195,In_370,In_455);
and U196 (N_196,In_255,In_117);
or U197 (N_197,In_256,In_430);
nor U198 (N_198,In_482,In_414);
xor U199 (N_199,In_71,In_143);
nor U200 (N_200,In_362,N_133);
nor U201 (N_201,In_35,In_396);
xnor U202 (N_202,In_99,In_192);
or U203 (N_203,N_41,N_89);
nor U204 (N_204,N_194,In_72);
xnor U205 (N_205,N_137,N_99);
or U206 (N_206,N_92,N_58);
or U207 (N_207,In_323,In_484);
and U208 (N_208,In_161,In_178);
nor U209 (N_209,In_380,N_109);
nor U210 (N_210,In_189,N_182);
nand U211 (N_211,In_252,In_251);
or U212 (N_212,N_197,N_118);
xor U213 (N_213,In_294,N_155);
and U214 (N_214,N_32,N_119);
nand U215 (N_215,N_104,In_254);
or U216 (N_216,N_56,N_112);
or U217 (N_217,N_144,N_108);
nor U218 (N_218,N_80,N_186);
and U219 (N_219,N_167,N_84);
or U220 (N_220,N_42,In_437);
xor U221 (N_221,N_25,N_37);
xor U222 (N_222,In_186,In_450);
nor U223 (N_223,N_9,In_126);
nor U224 (N_224,N_178,N_27);
and U225 (N_225,N_183,N_165);
xor U226 (N_226,In_205,In_443);
and U227 (N_227,N_181,N_132);
or U228 (N_228,N_71,N_184);
nor U229 (N_229,In_308,N_188);
nand U230 (N_230,N_111,In_41);
nand U231 (N_231,N_7,In_412);
nor U232 (N_232,N_115,N_45);
nand U233 (N_233,In_51,N_35);
and U234 (N_234,N_16,N_131);
nor U235 (N_235,N_64,N_19);
nor U236 (N_236,N_40,N_34);
or U237 (N_237,In_466,N_13);
or U238 (N_238,N_180,N_2);
xor U239 (N_239,N_91,N_107);
and U240 (N_240,N_76,N_10);
or U241 (N_241,N_1,In_383);
nor U242 (N_242,N_193,N_147);
nand U243 (N_243,In_233,In_336);
or U244 (N_244,N_46,In_360);
nand U245 (N_245,N_195,N_69);
nand U246 (N_246,N_113,In_114);
xor U247 (N_247,N_23,N_143);
and U248 (N_248,In_441,N_148);
and U249 (N_249,N_153,N_24);
nor U250 (N_250,N_114,N_11);
xor U251 (N_251,N_152,N_170);
xnor U252 (N_252,N_159,In_235);
nor U253 (N_253,In_228,N_161);
xor U254 (N_254,In_335,N_149);
xnor U255 (N_255,N_63,N_60);
and U256 (N_256,N_157,N_21);
nand U257 (N_257,In_34,N_123);
xor U258 (N_258,In_492,N_128);
xor U259 (N_259,In_464,N_52);
nor U260 (N_260,N_130,N_168);
xnor U261 (N_261,N_146,N_62);
or U262 (N_262,N_6,In_213);
or U263 (N_263,N_4,In_93);
and U264 (N_264,In_69,N_136);
nor U265 (N_265,In_248,N_65);
or U266 (N_266,In_326,In_121);
nor U267 (N_267,N_189,N_176);
or U268 (N_268,N_97,N_12);
and U269 (N_269,N_154,N_169);
or U270 (N_270,N_162,In_291);
or U271 (N_271,N_26,N_74);
and U272 (N_272,In_229,N_179);
or U273 (N_273,N_135,In_207);
nand U274 (N_274,In_22,In_282);
nand U275 (N_275,In_145,N_47);
or U276 (N_276,In_13,N_103);
or U277 (N_277,N_50,N_61);
nand U278 (N_278,N_185,N_14);
nand U279 (N_279,In_393,N_105);
and U280 (N_280,In_54,In_301);
xnor U281 (N_281,N_55,In_266);
and U282 (N_282,N_15,In_278);
nand U283 (N_283,N_5,N_124);
xor U284 (N_284,N_38,N_98);
nand U285 (N_285,In_167,N_49);
nor U286 (N_286,N_191,In_295);
and U287 (N_287,N_199,N_127);
and U288 (N_288,N_87,N_90);
xnor U289 (N_289,In_334,N_190);
nand U290 (N_290,N_134,In_262);
and U291 (N_291,In_265,In_399);
nand U292 (N_292,In_356,N_79);
xnor U293 (N_293,In_382,In_222);
and U294 (N_294,In_133,N_36);
or U295 (N_295,N_187,In_28);
xnor U296 (N_296,N_33,N_48);
or U297 (N_297,N_70,N_141);
nor U298 (N_298,In_74,In_367);
and U299 (N_299,N_151,N_142);
nor U300 (N_300,In_316,In_122);
and U301 (N_301,In_18,In_55);
xor U302 (N_302,N_120,N_140);
xor U303 (N_303,In_384,In_345);
nand U304 (N_304,N_57,N_43);
nor U305 (N_305,N_81,In_90);
or U306 (N_306,N_138,N_44);
nand U307 (N_307,N_125,N_39);
and U308 (N_308,N_59,N_67);
nand U309 (N_309,N_17,N_73);
xor U310 (N_310,N_102,N_116);
nand U311 (N_311,N_93,N_101);
nand U312 (N_312,N_0,N_121);
xor U313 (N_313,N_196,N_53);
xnor U314 (N_314,N_54,N_29);
or U315 (N_315,N_174,In_197);
nand U316 (N_316,N_198,N_171);
or U317 (N_317,N_72,In_62);
nor U318 (N_318,N_166,N_51);
and U319 (N_319,N_139,In_113);
nand U320 (N_320,N_160,N_8);
nor U321 (N_321,In_195,N_145);
or U322 (N_322,N_88,N_30);
nor U323 (N_323,N_164,N_158);
nand U324 (N_324,N_77,N_96);
and U325 (N_325,In_105,N_110);
nand U326 (N_326,N_68,In_36);
and U327 (N_327,N_75,N_66);
and U328 (N_328,N_95,N_94);
and U329 (N_329,In_271,N_163);
and U330 (N_330,N_20,N_106);
and U331 (N_331,N_22,N_156);
nor U332 (N_332,N_86,N_192);
or U333 (N_333,In_311,In_461);
and U334 (N_334,N_175,N_18);
nand U335 (N_335,In_490,N_117);
and U336 (N_336,In_4,N_129);
xor U337 (N_337,In_355,In_15);
or U338 (N_338,N_28,N_31);
nor U339 (N_339,In_177,In_411);
and U340 (N_340,N_100,N_85);
or U341 (N_341,In_342,In_350);
xor U342 (N_342,N_122,N_177);
nor U343 (N_343,N_172,N_3);
nor U344 (N_344,In_333,N_83);
or U345 (N_345,N_126,In_472);
and U346 (N_346,In_234,N_78);
and U347 (N_347,In_379,In_227);
xor U348 (N_348,N_82,In_217);
nand U349 (N_349,N_150,N_173);
xor U350 (N_350,N_121,N_168);
nand U351 (N_351,N_127,In_55);
nor U352 (N_352,In_362,In_207);
or U353 (N_353,N_91,N_153);
nand U354 (N_354,In_233,In_262);
nor U355 (N_355,In_333,In_36);
nand U356 (N_356,N_191,N_171);
and U357 (N_357,N_117,N_171);
and U358 (N_358,N_140,N_174);
or U359 (N_359,N_128,N_198);
xnor U360 (N_360,In_367,In_51);
nor U361 (N_361,N_63,N_12);
xnor U362 (N_362,In_235,In_282);
nand U363 (N_363,N_168,N_189);
xnor U364 (N_364,In_342,N_73);
or U365 (N_365,N_64,In_28);
or U366 (N_366,N_62,N_153);
or U367 (N_367,In_382,In_213);
nor U368 (N_368,N_151,N_0);
xnor U369 (N_369,N_138,N_121);
xor U370 (N_370,In_227,N_37);
nor U371 (N_371,N_39,In_192);
nor U372 (N_372,In_362,N_148);
xnor U373 (N_373,In_472,N_15);
and U374 (N_374,N_130,N_50);
or U375 (N_375,N_62,N_42);
nor U376 (N_376,In_72,In_360);
nor U377 (N_377,N_160,N_198);
xor U378 (N_378,N_20,N_123);
or U379 (N_379,In_294,N_19);
xor U380 (N_380,In_271,N_2);
or U381 (N_381,N_172,In_466);
nand U382 (N_382,N_198,N_185);
xnor U383 (N_383,In_262,N_168);
nor U384 (N_384,N_96,N_36);
and U385 (N_385,N_17,In_308);
and U386 (N_386,In_311,N_141);
nor U387 (N_387,In_217,N_198);
xnor U388 (N_388,In_161,N_104);
nor U389 (N_389,N_167,N_98);
nand U390 (N_390,In_301,In_490);
xnor U391 (N_391,N_82,N_103);
nand U392 (N_392,In_122,N_116);
nor U393 (N_393,N_67,N_91);
and U394 (N_394,In_295,In_15);
or U395 (N_395,In_308,In_412);
or U396 (N_396,N_76,N_138);
and U397 (N_397,N_42,In_195);
and U398 (N_398,In_356,N_125);
and U399 (N_399,N_1,N_69);
nor U400 (N_400,N_277,N_273);
xor U401 (N_401,N_336,N_296);
xor U402 (N_402,N_395,N_239);
xor U403 (N_403,N_321,N_348);
nand U404 (N_404,N_326,N_249);
nor U405 (N_405,N_286,N_298);
or U406 (N_406,N_381,N_283);
nand U407 (N_407,N_274,N_337);
xnor U408 (N_408,N_302,N_370);
and U409 (N_409,N_371,N_203);
xnor U410 (N_410,N_354,N_369);
and U411 (N_411,N_372,N_309);
or U412 (N_412,N_361,N_256);
and U413 (N_413,N_243,N_317);
nor U414 (N_414,N_234,N_271);
and U415 (N_415,N_366,N_291);
nor U416 (N_416,N_259,N_209);
nand U417 (N_417,N_299,N_233);
and U418 (N_418,N_315,N_282);
or U419 (N_419,N_264,N_327);
nand U420 (N_420,N_288,N_367);
or U421 (N_421,N_376,N_303);
xnor U422 (N_422,N_229,N_397);
xor U423 (N_423,N_211,N_386);
nor U424 (N_424,N_265,N_329);
xnor U425 (N_425,N_280,N_230);
and U426 (N_426,N_232,N_224);
xnor U427 (N_427,N_379,N_260);
nand U428 (N_428,N_295,N_284);
and U429 (N_429,N_385,N_287);
xor U430 (N_430,N_347,N_206);
nor U431 (N_431,N_279,N_208);
nor U432 (N_432,N_335,N_262);
nor U433 (N_433,N_306,N_364);
nor U434 (N_434,N_226,N_377);
and U435 (N_435,N_242,N_305);
nand U436 (N_436,N_251,N_345);
nor U437 (N_437,N_318,N_328);
xor U438 (N_438,N_268,N_263);
or U439 (N_439,N_236,N_300);
nor U440 (N_440,N_350,N_297);
nor U441 (N_441,N_355,N_320);
xor U442 (N_442,N_272,N_332);
nand U443 (N_443,N_235,N_219);
nand U444 (N_444,N_240,N_252);
xor U445 (N_445,N_257,N_352);
or U446 (N_446,N_330,N_338);
nor U447 (N_447,N_325,N_204);
nor U448 (N_448,N_289,N_270);
nor U449 (N_449,N_246,N_205);
nor U450 (N_450,N_313,N_258);
and U451 (N_451,N_393,N_213);
or U452 (N_452,N_275,N_356);
or U453 (N_453,N_293,N_222);
nand U454 (N_454,N_374,N_245);
nor U455 (N_455,N_387,N_241);
nor U456 (N_456,N_380,N_254);
and U457 (N_457,N_359,N_333);
nor U458 (N_458,N_216,N_394);
nand U459 (N_459,N_292,N_248);
and U460 (N_460,N_261,N_331);
nand U461 (N_461,N_382,N_343);
nand U462 (N_462,N_389,N_368);
and U463 (N_463,N_391,N_215);
and U464 (N_464,N_228,N_316);
nor U465 (N_465,N_384,N_398);
and U466 (N_466,N_324,N_323);
nand U467 (N_467,N_383,N_390);
nand U468 (N_468,N_304,N_221);
nor U469 (N_469,N_278,N_244);
xor U470 (N_470,N_250,N_267);
nor U471 (N_471,N_362,N_399);
nor U472 (N_472,N_238,N_231);
and U473 (N_473,N_255,N_351);
or U474 (N_474,N_217,N_357);
nand U475 (N_475,N_227,N_301);
and U476 (N_476,N_223,N_349);
nand U477 (N_477,N_334,N_311);
nand U478 (N_478,N_373,N_363);
nor U479 (N_479,N_225,N_378);
and U480 (N_480,N_207,N_269);
nor U481 (N_481,N_358,N_392);
xnor U482 (N_482,N_375,N_319);
nand U483 (N_483,N_308,N_285);
xnor U484 (N_484,N_200,N_237);
xor U485 (N_485,N_218,N_307);
and U486 (N_486,N_388,N_281);
nor U487 (N_487,N_266,N_365);
xor U488 (N_488,N_202,N_247);
nor U489 (N_489,N_201,N_346);
nand U490 (N_490,N_322,N_396);
nor U491 (N_491,N_210,N_353);
xor U492 (N_492,N_294,N_220);
xor U493 (N_493,N_290,N_314);
or U494 (N_494,N_339,N_310);
nand U495 (N_495,N_360,N_342);
nand U496 (N_496,N_341,N_214);
nor U497 (N_497,N_344,N_212);
xor U498 (N_498,N_340,N_276);
and U499 (N_499,N_253,N_312);
nor U500 (N_500,N_255,N_349);
nand U501 (N_501,N_227,N_293);
xnor U502 (N_502,N_358,N_317);
nand U503 (N_503,N_316,N_333);
nor U504 (N_504,N_365,N_236);
and U505 (N_505,N_333,N_350);
nand U506 (N_506,N_397,N_256);
xor U507 (N_507,N_365,N_346);
or U508 (N_508,N_312,N_388);
xor U509 (N_509,N_248,N_218);
and U510 (N_510,N_322,N_222);
and U511 (N_511,N_260,N_351);
nand U512 (N_512,N_351,N_206);
nand U513 (N_513,N_344,N_336);
nor U514 (N_514,N_267,N_200);
xor U515 (N_515,N_348,N_347);
nand U516 (N_516,N_301,N_262);
nand U517 (N_517,N_270,N_326);
xor U518 (N_518,N_253,N_354);
or U519 (N_519,N_349,N_230);
nand U520 (N_520,N_380,N_300);
nor U521 (N_521,N_372,N_318);
or U522 (N_522,N_266,N_393);
nand U523 (N_523,N_201,N_215);
xor U524 (N_524,N_335,N_372);
and U525 (N_525,N_320,N_240);
and U526 (N_526,N_226,N_310);
and U527 (N_527,N_288,N_237);
nand U528 (N_528,N_267,N_360);
and U529 (N_529,N_391,N_300);
nand U530 (N_530,N_356,N_218);
and U531 (N_531,N_338,N_214);
nand U532 (N_532,N_366,N_351);
and U533 (N_533,N_225,N_281);
or U534 (N_534,N_341,N_314);
or U535 (N_535,N_216,N_286);
nand U536 (N_536,N_299,N_399);
or U537 (N_537,N_216,N_218);
or U538 (N_538,N_281,N_234);
nand U539 (N_539,N_381,N_271);
nand U540 (N_540,N_303,N_215);
or U541 (N_541,N_277,N_247);
nor U542 (N_542,N_302,N_372);
nand U543 (N_543,N_277,N_296);
xor U544 (N_544,N_373,N_207);
and U545 (N_545,N_351,N_223);
nor U546 (N_546,N_243,N_316);
and U547 (N_547,N_364,N_386);
or U548 (N_548,N_250,N_202);
and U549 (N_549,N_388,N_393);
xnor U550 (N_550,N_281,N_209);
or U551 (N_551,N_301,N_384);
xnor U552 (N_552,N_380,N_377);
and U553 (N_553,N_299,N_251);
xor U554 (N_554,N_340,N_306);
nand U555 (N_555,N_263,N_209);
nand U556 (N_556,N_285,N_336);
xnor U557 (N_557,N_333,N_295);
or U558 (N_558,N_233,N_200);
xor U559 (N_559,N_354,N_322);
nor U560 (N_560,N_293,N_316);
or U561 (N_561,N_356,N_250);
nor U562 (N_562,N_387,N_257);
nor U563 (N_563,N_225,N_283);
or U564 (N_564,N_277,N_233);
nand U565 (N_565,N_271,N_345);
nor U566 (N_566,N_237,N_385);
xnor U567 (N_567,N_223,N_201);
nand U568 (N_568,N_232,N_226);
xor U569 (N_569,N_277,N_205);
nor U570 (N_570,N_356,N_389);
xor U571 (N_571,N_200,N_244);
and U572 (N_572,N_247,N_365);
nand U573 (N_573,N_238,N_385);
or U574 (N_574,N_324,N_271);
or U575 (N_575,N_289,N_292);
nor U576 (N_576,N_294,N_300);
nand U577 (N_577,N_205,N_226);
nor U578 (N_578,N_284,N_211);
nand U579 (N_579,N_354,N_348);
and U580 (N_580,N_272,N_366);
nand U581 (N_581,N_300,N_235);
nor U582 (N_582,N_377,N_234);
nor U583 (N_583,N_332,N_317);
nand U584 (N_584,N_343,N_221);
xor U585 (N_585,N_262,N_237);
xor U586 (N_586,N_387,N_325);
and U587 (N_587,N_328,N_300);
nor U588 (N_588,N_340,N_217);
nand U589 (N_589,N_366,N_263);
xnor U590 (N_590,N_272,N_249);
or U591 (N_591,N_281,N_384);
nand U592 (N_592,N_324,N_322);
xor U593 (N_593,N_309,N_369);
nor U594 (N_594,N_228,N_362);
nor U595 (N_595,N_269,N_306);
or U596 (N_596,N_390,N_391);
nand U597 (N_597,N_226,N_337);
or U598 (N_598,N_315,N_369);
or U599 (N_599,N_381,N_376);
xnor U600 (N_600,N_520,N_562);
xnor U601 (N_601,N_478,N_539);
or U602 (N_602,N_564,N_406);
or U603 (N_603,N_524,N_491);
or U604 (N_604,N_447,N_438);
and U605 (N_605,N_474,N_456);
or U606 (N_606,N_545,N_429);
xnor U607 (N_607,N_566,N_473);
and U608 (N_608,N_461,N_536);
nor U609 (N_609,N_567,N_578);
xnor U610 (N_610,N_479,N_581);
nand U611 (N_611,N_549,N_541);
and U612 (N_612,N_553,N_455);
or U613 (N_613,N_584,N_527);
nor U614 (N_614,N_445,N_498);
and U615 (N_615,N_501,N_522);
nand U616 (N_616,N_535,N_476);
and U617 (N_617,N_579,N_439);
nor U618 (N_618,N_568,N_440);
and U619 (N_619,N_526,N_471);
nand U620 (N_620,N_443,N_523);
xnor U621 (N_621,N_437,N_518);
or U622 (N_622,N_550,N_516);
and U623 (N_623,N_519,N_483);
or U624 (N_624,N_577,N_582);
nand U625 (N_625,N_414,N_413);
or U626 (N_626,N_555,N_446);
nand U627 (N_627,N_521,N_534);
nand U628 (N_628,N_420,N_515);
or U629 (N_629,N_411,N_513);
nor U630 (N_630,N_466,N_563);
nand U631 (N_631,N_401,N_454);
nand U632 (N_632,N_587,N_552);
nor U633 (N_633,N_595,N_505);
nor U634 (N_634,N_415,N_530);
and U635 (N_635,N_422,N_418);
nor U636 (N_636,N_484,N_481);
nand U637 (N_637,N_571,N_493);
and U638 (N_638,N_442,N_598);
xnor U639 (N_639,N_404,N_494);
or U640 (N_640,N_407,N_594);
or U641 (N_641,N_512,N_434);
and U642 (N_642,N_532,N_464);
nor U643 (N_643,N_589,N_528);
and U644 (N_644,N_585,N_435);
xor U645 (N_645,N_517,N_495);
or U646 (N_646,N_542,N_509);
nor U647 (N_647,N_569,N_427);
nand U648 (N_648,N_540,N_410);
nor U649 (N_649,N_458,N_499);
xnor U650 (N_650,N_432,N_490);
nor U651 (N_651,N_596,N_412);
and U652 (N_652,N_544,N_421);
xor U653 (N_653,N_428,N_425);
or U654 (N_654,N_575,N_580);
nor U655 (N_655,N_463,N_444);
and U656 (N_656,N_472,N_408);
nand U657 (N_657,N_405,N_590);
xor U658 (N_658,N_504,N_572);
nor U659 (N_659,N_573,N_460);
xnor U660 (N_660,N_486,N_469);
and U661 (N_661,N_475,N_487);
nor U662 (N_662,N_588,N_424);
and U663 (N_663,N_531,N_431);
and U664 (N_664,N_551,N_554);
nand U665 (N_665,N_548,N_565);
xor U666 (N_666,N_574,N_480);
nor U667 (N_667,N_506,N_496);
or U668 (N_668,N_462,N_488);
and U669 (N_669,N_537,N_583);
and U670 (N_670,N_529,N_525);
nand U671 (N_671,N_543,N_538);
or U672 (N_672,N_417,N_453);
and U673 (N_673,N_423,N_556);
or U674 (N_674,N_433,N_502);
xnor U675 (N_675,N_482,N_470);
nor U676 (N_676,N_508,N_465);
xnor U677 (N_677,N_403,N_511);
or U678 (N_678,N_409,N_570);
nor U679 (N_679,N_514,N_558);
or U680 (N_680,N_593,N_451);
nor U681 (N_681,N_500,N_485);
nand U682 (N_682,N_419,N_477);
nor U683 (N_683,N_467,N_599);
nand U684 (N_684,N_441,N_426);
nor U685 (N_685,N_492,N_557);
nor U686 (N_686,N_452,N_560);
and U687 (N_687,N_459,N_586);
and U688 (N_688,N_591,N_561);
xor U689 (N_689,N_546,N_597);
xor U690 (N_690,N_436,N_510);
or U691 (N_691,N_497,N_507);
and U692 (N_692,N_400,N_468);
xor U693 (N_693,N_448,N_449);
nand U694 (N_694,N_489,N_503);
nand U695 (N_695,N_533,N_592);
nor U696 (N_696,N_430,N_450);
nand U697 (N_697,N_416,N_402);
and U698 (N_698,N_559,N_457);
nand U699 (N_699,N_547,N_576);
xor U700 (N_700,N_525,N_436);
or U701 (N_701,N_460,N_428);
nand U702 (N_702,N_411,N_491);
and U703 (N_703,N_594,N_502);
xor U704 (N_704,N_500,N_425);
nor U705 (N_705,N_510,N_554);
nor U706 (N_706,N_583,N_558);
and U707 (N_707,N_415,N_576);
or U708 (N_708,N_415,N_541);
nor U709 (N_709,N_435,N_437);
nand U710 (N_710,N_517,N_503);
nor U711 (N_711,N_532,N_471);
or U712 (N_712,N_525,N_466);
xor U713 (N_713,N_513,N_540);
xor U714 (N_714,N_485,N_418);
or U715 (N_715,N_530,N_515);
or U716 (N_716,N_478,N_422);
nor U717 (N_717,N_525,N_515);
nor U718 (N_718,N_585,N_461);
and U719 (N_719,N_455,N_456);
nor U720 (N_720,N_460,N_517);
and U721 (N_721,N_580,N_554);
nand U722 (N_722,N_430,N_407);
nand U723 (N_723,N_496,N_522);
and U724 (N_724,N_598,N_403);
nor U725 (N_725,N_402,N_527);
xor U726 (N_726,N_408,N_474);
and U727 (N_727,N_555,N_533);
or U728 (N_728,N_594,N_467);
nor U729 (N_729,N_516,N_519);
nand U730 (N_730,N_588,N_565);
xnor U731 (N_731,N_590,N_420);
and U732 (N_732,N_423,N_506);
xor U733 (N_733,N_548,N_479);
nor U734 (N_734,N_452,N_475);
xnor U735 (N_735,N_459,N_468);
xnor U736 (N_736,N_574,N_522);
or U737 (N_737,N_565,N_427);
nor U738 (N_738,N_511,N_472);
and U739 (N_739,N_511,N_493);
nand U740 (N_740,N_455,N_551);
xor U741 (N_741,N_587,N_522);
nand U742 (N_742,N_412,N_473);
xor U743 (N_743,N_434,N_529);
nand U744 (N_744,N_543,N_429);
and U745 (N_745,N_482,N_590);
nor U746 (N_746,N_405,N_522);
xnor U747 (N_747,N_592,N_473);
xnor U748 (N_748,N_586,N_476);
and U749 (N_749,N_402,N_444);
xnor U750 (N_750,N_542,N_424);
nand U751 (N_751,N_580,N_589);
or U752 (N_752,N_534,N_593);
xnor U753 (N_753,N_546,N_537);
and U754 (N_754,N_553,N_505);
xnor U755 (N_755,N_442,N_409);
and U756 (N_756,N_470,N_562);
nor U757 (N_757,N_414,N_520);
or U758 (N_758,N_597,N_418);
and U759 (N_759,N_469,N_587);
nor U760 (N_760,N_556,N_538);
xnor U761 (N_761,N_556,N_501);
nand U762 (N_762,N_518,N_446);
or U763 (N_763,N_591,N_508);
nor U764 (N_764,N_468,N_535);
or U765 (N_765,N_451,N_561);
nand U766 (N_766,N_448,N_541);
and U767 (N_767,N_524,N_556);
or U768 (N_768,N_589,N_536);
nor U769 (N_769,N_456,N_526);
nor U770 (N_770,N_423,N_547);
nor U771 (N_771,N_591,N_457);
or U772 (N_772,N_496,N_404);
nor U773 (N_773,N_575,N_566);
nand U774 (N_774,N_517,N_535);
or U775 (N_775,N_418,N_437);
nor U776 (N_776,N_549,N_402);
or U777 (N_777,N_533,N_553);
or U778 (N_778,N_531,N_408);
nand U779 (N_779,N_433,N_521);
and U780 (N_780,N_531,N_481);
xnor U781 (N_781,N_511,N_457);
nor U782 (N_782,N_521,N_425);
nor U783 (N_783,N_430,N_424);
or U784 (N_784,N_582,N_445);
or U785 (N_785,N_494,N_433);
nor U786 (N_786,N_421,N_493);
xnor U787 (N_787,N_552,N_539);
xor U788 (N_788,N_429,N_484);
or U789 (N_789,N_556,N_464);
or U790 (N_790,N_521,N_528);
and U791 (N_791,N_482,N_501);
nor U792 (N_792,N_415,N_412);
and U793 (N_793,N_515,N_454);
or U794 (N_794,N_469,N_436);
nor U795 (N_795,N_423,N_486);
xor U796 (N_796,N_470,N_474);
nand U797 (N_797,N_583,N_528);
xor U798 (N_798,N_455,N_434);
or U799 (N_799,N_425,N_572);
nor U800 (N_800,N_752,N_794);
and U801 (N_801,N_707,N_725);
or U802 (N_802,N_740,N_691);
nor U803 (N_803,N_775,N_739);
nand U804 (N_804,N_641,N_728);
nor U805 (N_805,N_726,N_757);
nor U806 (N_806,N_665,N_733);
nand U807 (N_807,N_652,N_636);
xor U808 (N_808,N_784,N_699);
nor U809 (N_809,N_727,N_661);
nor U810 (N_810,N_756,N_700);
nand U811 (N_811,N_731,N_619);
xor U812 (N_812,N_714,N_702);
nand U813 (N_813,N_710,N_717);
or U814 (N_814,N_716,N_603);
nor U815 (N_815,N_704,N_643);
nor U816 (N_816,N_780,N_692);
nand U817 (N_817,N_631,N_747);
and U818 (N_818,N_654,N_608);
nor U819 (N_819,N_783,N_650);
nor U820 (N_820,N_778,N_790);
xor U821 (N_821,N_750,N_645);
or U822 (N_822,N_796,N_754);
nor U823 (N_823,N_737,N_697);
nor U824 (N_824,N_687,N_760);
xor U825 (N_825,N_708,N_604);
or U826 (N_826,N_635,N_673);
xor U827 (N_827,N_639,N_656);
nor U828 (N_828,N_690,N_625);
or U829 (N_829,N_615,N_749);
nand U830 (N_830,N_605,N_621);
xor U831 (N_831,N_715,N_669);
nor U832 (N_832,N_683,N_633);
or U833 (N_833,N_718,N_644);
and U834 (N_834,N_688,N_667);
or U835 (N_835,N_789,N_773);
or U836 (N_836,N_674,N_614);
nor U837 (N_837,N_632,N_616);
nand U838 (N_838,N_613,N_768);
or U839 (N_839,N_620,N_767);
and U840 (N_840,N_763,N_722);
nand U841 (N_841,N_666,N_751);
nand U842 (N_842,N_770,N_676);
and U843 (N_843,N_629,N_745);
or U844 (N_844,N_779,N_764);
or U845 (N_845,N_719,N_709);
xor U846 (N_846,N_762,N_606);
and U847 (N_847,N_686,N_617);
and U848 (N_848,N_677,N_637);
nor U849 (N_849,N_701,N_706);
xor U850 (N_850,N_729,N_774);
nor U851 (N_851,N_735,N_658);
and U852 (N_852,N_678,N_689);
xnor U853 (N_853,N_680,N_797);
or U854 (N_854,N_647,N_662);
xnor U855 (N_855,N_713,N_723);
nand U856 (N_856,N_798,N_732);
or U857 (N_857,N_782,N_685);
or U858 (N_858,N_761,N_787);
xor U859 (N_859,N_696,N_785);
or U860 (N_860,N_659,N_743);
nor U861 (N_861,N_651,N_623);
xnor U862 (N_862,N_628,N_765);
nor U863 (N_863,N_712,N_698);
nor U864 (N_864,N_653,N_720);
nand U865 (N_865,N_781,N_612);
and U866 (N_866,N_758,N_759);
xnor U867 (N_867,N_642,N_695);
nor U868 (N_868,N_655,N_791);
nand U869 (N_869,N_611,N_755);
nor U870 (N_870,N_772,N_694);
or U871 (N_871,N_646,N_601);
and U872 (N_872,N_624,N_771);
nor U873 (N_873,N_607,N_675);
or U874 (N_874,N_634,N_744);
and U875 (N_875,N_721,N_618);
or U876 (N_876,N_703,N_753);
nand U877 (N_877,N_600,N_610);
xnor U878 (N_878,N_711,N_681);
or U879 (N_879,N_640,N_630);
nand U880 (N_880,N_736,N_734);
nand U881 (N_881,N_668,N_799);
and U882 (N_882,N_730,N_657);
or U883 (N_883,N_742,N_648);
and U884 (N_884,N_638,N_788);
nand U885 (N_885,N_660,N_682);
nor U886 (N_886,N_684,N_724);
and U887 (N_887,N_609,N_664);
and U888 (N_888,N_776,N_670);
nand U889 (N_889,N_602,N_748);
nor U890 (N_890,N_741,N_693);
and U891 (N_891,N_769,N_746);
and U892 (N_892,N_649,N_627);
and U893 (N_893,N_738,N_792);
and U894 (N_894,N_777,N_679);
nor U895 (N_895,N_795,N_766);
xnor U896 (N_896,N_626,N_663);
nand U897 (N_897,N_786,N_705);
and U898 (N_898,N_793,N_672);
nor U899 (N_899,N_671,N_622);
nand U900 (N_900,N_733,N_668);
xor U901 (N_901,N_660,N_677);
and U902 (N_902,N_715,N_606);
nand U903 (N_903,N_607,N_742);
and U904 (N_904,N_603,N_630);
xnor U905 (N_905,N_691,N_796);
nor U906 (N_906,N_730,N_664);
and U907 (N_907,N_650,N_614);
nand U908 (N_908,N_750,N_711);
xor U909 (N_909,N_730,N_764);
or U910 (N_910,N_640,N_727);
xor U911 (N_911,N_740,N_788);
and U912 (N_912,N_706,N_620);
nor U913 (N_913,N_745,N_717);
nand U914 (N_914,N_731,N_782);
and U915 (N_915,N_633,N_753);
nor U916 (N_916,N_763,N_731);
xnor U917 (N_917,N_615,N_727);
xnor U918 (N_918,N_603,N_722);
nor U919 (N_919,N_688,N_691);
or U920 (N_920,N_704,N_661);
xnor U921 (N_921,N_683,N_661);
nand U922 (N_922,N_657,N_752);
xnor U923 (N_923,N_747,N_796);
nor U924 (N_924,N_611,N_783);
nor U925 (N_925,N_665,N_727);
xnor U926 (N_926,N_635,N_646);
nand U927 (N_927,N_778,N_612);
nor U928 (N_928,N_775,N_787);
or U929 (N_929,N_770,N_642);
xnor U930 (N_930,N_729,N_685);
or U931 (N_931,N_665,N_754);
and U932 (N_932,N_608,N_756);
nand U933 (N_933,N_618,N_655);
nor U934 (N_934,N_757,N_615);
or U935 (N_935,N_790,N_699);
nor U936 (N_936,N_704,N_731);
xor U937 (N_937,N_668,N_717);
xnor U938 (N_938,N_699,N_621);
xnor U939 (N_939,N_607,N_672);
nand U940 (N_940,N_710,N_734);
or U941 (N_941,N_724,N_610);
nor U942 (N_942,N_675,N_603);
nor U943 (N_943,N_669,N_666);
nand U944 (N_944,N_624,N_783);
nor U945 (N_945,N_781,N_614);
nor U946 (N_946,N_613,N_685);
or U947 (N_947,N_725,N_796);
and U948 (N_948,N_664,N_745);
and U949 (N_949,N_714,N_633);
and U950 (N_950,N_728,N_610);
or U951 (N_951,N_792,N_636);
or U952 (N_952,N_693,N_651);
nand U953 (N_953,N_755,N_791);
and U954 (N_954,N_712,N_796);
and U955 (N_955,N_766,N_733);
nand U956 (N_956,N_655,N_719);
and U957 (N_957,N_719,N_653);
xnor U958 (N_958,N_749,N_733);
nand U959 (N_959,N_671,N_657);
and U960 (N_960,N_745,N_704);
and U961 (N_961,N_611,N_622);
nand U962 (N_962,N_615,N_658);
xnor U963 (N_963,N_687,N_773);
or U964 (N_964,N_725,N_768);
or U965 (N_965,N_679,N_612);
xnor U966 (N_966,N_643,N_737);
xor U967 (N_967,N_770,N_701);
and U968 (N_968,N_656,N_642);
nor U969 (N_969,N_629,N_655);
and U970 (N_970,N_685,N_784);
xor U971 (N_971,N_647,N_642);
xor U972 (N_972,N_681,N_799);
nand U973 (N_973,N_783,N_695);
or U974 (N_974,N_746,N_660);
nand U975 (N_975,N_781,N_709);
and U976 (N_976,N_621,N_744);
nand U977 (N_977,N_724,N_736);
nand U978 (N_978,N_604,N_676);
and U979 (N_979,N_672,N_761);
xnor U980 (N_980,N_635,N_689);
and U981 (N_981,N_732,N_659);
nand U982 (N_982,N_770,N_761);
xor U983 (N_983,N_660,N_768);
and U984 (N_984,N_770,N_796);
and U985 (N_985,N_656,N_697);
xor U986 (N_986,N_607,N_673);
nor U987 (N_987,N_702,N_699);
or U988 (N_988,N_787,N_718);
xnor U989 (N_989,N_724,N_731);
nor U990 (N_990,N_742,N_620);
xnor U991 (N_991,N_668,N_605);
nand U992 (N_992,N_677,N_789);
nor U993 (N_993,N_743,N_600);
or U994 (N_994,N_747,N_604);
nor U995 (N_995,N_663,N_719);
nand U996 (N_996,N_729,N_743);
nand U997 (N_997,N_737,N_750);
nand U998 (N_998,N_659,N_684);
nor U999 (N_999,N_741,N_791);
or U1000 (N_1000,N_970,N_886);
nand U1001 (N_1001,N_903,N_871);
or U1002 (N_1002,N_945,N_910);
and U1003 (N_1003,N_900,N_870);
nand U1004 (N_1004,N_956,N_862);
or U1005 (N_1005,N_825,N_931);
xnor U1006 (N_1006,N_979,N_834);
nor U1007 (N_1007,N_845,N_983);
nand U1008 (N_1008,N_892,N_971);
nor U1009 (N_1009,N_876,N_920);
and U1010 (N_1010,N_961,N_957);
or U1011 (N_1011,N_866,N_818);
xor U1012 (N_1012,N_984,N_828);
xor U1013 (N_1013,N_960,N_918);
or U1014 (N_1014,N_952,N_875);
nor U1015 (N_1015,N_829,N_838);
or U1016 (N_1016,N_915,N_954);
or U1017 (N_1017,N_977,N_996);
xor U1018 (N_1018,N_988,N_981);
and U1019 (N_1019,N_946,N_925);
xor U1020 (N_1020,N_923,N_938);
xnor U1021 (N_1021,N_867,N_992);
nand U1022 (N_1022,N_926,N_985);
xnor U1023 (N_1023,N_833,N_901);
xnor U1024 (N_1024,N_819,N_813);
and U1025 (N_1025,N_878,N_831);
xnor U1026 (N_1026,N_824,N_963);
and U1027 (N_1027,N_965,N_858);
nand U1028 (N_1028,N_949,N_815);
and U1029 (N_1029,N_980,N_999);
and U1030 (N_1030,N_941,N_940);
xnor U1031 (N_1031,N_850,N_873);
nor U1032 (N_1032,N_894,N_986);
xor U1033 (N_1033,N_885,N_914);
nor U1034 (N_1034,N_803,N_844);
or U1035 (N_1035,N_859,N_972);
xor U1036 (N_1036,N_806,N_888);
or U1037 (N_1037,N_881,N_820);
xor U1038 (N_1038,N_812,N_978);
and U1039 (N_1039,N_853,N_895);
xnor U1040 (N_1040,N_861,N_913);
nand U1041 (N_1041,N_869,N_809);
nand U1042 (N_1042,N_848,N_933);
xnor U1043 (N_1043,N_880,N_942);
nand U1044 (N_1044,N_922,N_863);
or U1045 (N_1045,N_932,N_976);
nand U1046 (N_1046,N_808,N_994);
nor U1047 (N_1047,N_928,N_800);
xnor U1048 (N_1048,N_997,N_990);
nand U1049 (N_1049,N_917,N_830);
nand U1050 (N_1050,N_935,N_854);
nand U1051 (N_1051,N_899,N_936);
xnor U1052 (N_1052,N_889,N_953);
or U1053 (N_1053,N_840,N_811);
or U1054 (N_1054,N_827,N_930);
xnor U1055 (N_1055,N_912,N_842);
nand U1056 (N_1056,N_849,N_904);
nand U1057 (N_1057,N_958,N_877);
and U1058 (N_1058,N_857,N_929);
nor U1059 (N_1059,N_989,N_968);
xnor U1060 (N_1060,N_874,N_810);
nor U1061 (N_1061,N_967,N_883);
xor U1062 (N_1062,N_982,N_856);
nand U1063 (N_1063,N_839,N_826);
xor U1064 (N_1064,N_804,N_882);
nand U1065 (N_1065,N_890,N_851);
xnor U1066 (N_1066,N_966,N_823);
nand U1067 (N_1067,N_934,N_975);
xnor U1068 (N_1068,N_924,N_887);
xnor U1069 (N_1069,N_962,N_807);
or U1070 (N_1070,N_969,N_821);
or U1071 (N_1071,N_906,N_879);
or U1072 (N_1072,N_896,N_843);
xor U1073 (N_1073,N_816,N_852);
or U1074 (N_1074,N_905,N_891);
or U1075 (N_1075,N_998,N_817);
nand U1076 (N_1076,N_919,N_907);
nor U1077 (N_1077,N_955,N_855);
xnor U1078 (N_1078,N_947,N_836);
nor U1079 (N_1079,N_872,N_835);
nand U1080 (N_1080,N_944,N_908);
nor U1081 (N_1081,N_974,N_847);
nand U1082 (N_1082,N_837,N_865);
and U1083 (N_1083,N_893,N_846);
nand U1084 (N_1084,N_860,N_973);
nor U1085 (N_1085,N_951,N_993);
or U1086 (N_1086,N_964,N_995);
or U1087 (N_1087,N_939,N_802);
nor U1088 (N_1088,N_841,N_991);
or U1089 (N_1089,N_832,N_822);
nor U1090 (N_1090,N_959,N_884);
or U1091 (N_1091,N_916,N_948);
nor U1092 (N_1092,N_943,N_987);
xor U1093 (N_1093,N_921,N_868);
nor U1094 (N_1094,N_864,N_950);
or U1095 (N_1095,N_898,N_897);
and U1096 (N_1096,N_927,N_937);
xnor U1097 (N_1097,N_911,N_805);
nor U1098 (N_1098,N_801,N_902);
and U1099 (N_1099,N_814,N_909);
nand U1100 (N_1100,N_896,N_966);
nand U1101 (N_1101,N_972,N_836);
or U1102 (N_1102,N_885,N_988);
and U1103 (N_1103,N_867,N_859);
nor U1104 (N_1104,N_850,N_830);
nand U1105 (N_1105,N_847,N_894);
and U1106 (N_1106,N_890,N_988);
nor U1107 (N_1107,N_830,N_941);
xnor U1108 (N_1108,N_837,N_818);
nor U1109 (N_1109,N_815,N_909);
and U1110 (N_1110,N_956,N_981);
xor U1111 (N_1111,N_872,N_946);
nor U1112 (N_1112,N_801,N_810);
and U1113 (N_1113,N_846,N_845);
nor U1114 (N_1114,N_931,N_980);
nand U1115 (N_1115,N_869,N_907);
xnor U1116 (N_1116,N_834,N_872);
and U1117 (N_1117,N_816,N_892);
or U1118 (N_1118,N_861,N_859);
nand U1119 (N_1119,N_908,N_986);
and U1120 (N_1120,N_893,N_969);
nor U1121 (N_1121,N_960,N_944);
xnor U1122 (N_1122,N_832,N_811);
nor U1123 (N_1123,N_903,N_932);
or U1124 (N_1124,N_810,N_872);
or U1125 (N_1125,N_827,N_942);
or U1126 (N_1126,N_935,N_898);
nand U1127 (N_1127,N_815,N_825);
or U1128 (N_1128,N_985,N_998);
xnor U1129 (N_1129,N_921,N_867);
or U1130 (N_1130,N_817,N_938);
nand U1131 (N_1131,N_880,N_947);
and U1132 (N_1132,N_991,N_813);
nand U1133 (N_1133,N_868,N_983);
or U1134 (N_1134,N_944,N_942);
xnor U1135 (N_1135,N_839,N_880);
and U1136 (N_1136,N_934,N_996);
or U1137 (N_1137,N_957,N_977);
or U1138 (N_1138,N_800,N_932);
and U1139 (N_1139,N_890,N_814);
and U1140 (N_1140,N_841,N_940);
nor U1141 (N_1141,N_821,N_810);
nand U1142 (N_1142,N_994,N_885);
nor U1143 (N_1143,N_910,N_904);
nor U1144 (N_1144,N_900,N_853);
or U1145 (N_1145,N_946,N_880);
nor U1146 (N_1146,N_870,N_854);
nand U1147 (N_1147,N_991,N_918);
and U1148 (N_1148,N_941,N_927);
or U1149 (N_1149,N_996,N_995);
xnor U1150 (N_1150,N_994,N_852);
and U1151 (N_1151,N_851,N_995);
and U1152 (N_1152,N_829,N_853);
nand U1153 (N_1153,N_864,N_860);
nor U1154 (N_1154,N_865,N_806);
xor U1155 (N_1155,N_923,N_970);
and U1156 (N_1156,N_828,N_885);
or U1157 (N_1157,N_881,N_906);
nor U1158 (N_1158,N_831,N_995);
nand U1159 (N_1159,N_834,N_813);
xnor U1160 (N_1160,N_836,N_863);
or U1161 (N_1161,N_827,N_878);
nand U1162 (N_1162,N_849,N_983);
xnor U1163 (N_1163,N_860,N_909);
xor U1164 (N_1164,N_976,N_950);
xnor U1165 (N_1165,N_927,N_924);
nand U1166 (N_1166,N_884,N_893);
nand U1167 (N_1167,N_941,N_943);
nand U1168 (N_1168,N_889,N_959);
nor U1169 (N_1169,N_809,N_816);
or U1170 (N_1170,N_821,N_940);
nor U1171 (N_1171,N_851,N_976);
and U1172 (N_1172,N_945,N_970);
or U1173 (N_1173,N_875,N_917);
nand U1174 (N_1174,N_929,N_918);
nor U1175 (N_1175,N_997,N_966);
and U1176 (N_1176,N_962,N_918);
or U1177 (N_1177,N_813,N_835);
nand U1178 (N_1178,N_963,N_943);
and U1179 (N_1179,N_872,N_871);
or U1180 (N_1180,N_803,N_867);
nand U1181 (N_1181,N_920,N_912);
or U1182 (N_1182,N_959,N_987);
and U1183 (N_1183,N_960,N_857);
and U1184 (N_1184,N_944,N_990);
nand U1185 (N_1185,N_896,N_815);
nand U1186 (N_1186,N_937,N_891);
and U1187 (N_1187,N_999,N_860);
nand U1188 (N_1188,N_939,N_824);
nand U1189 (N_1189,N_880,N_851);
nand U1190 (N_1190,N_990,N_977);
nor U1191 (N_1191,N_991,N_977);
or U1192 (N_1192,N_982,N_888);
xor U1193 (N_1193,N_968,N_878);
xnor U1194 (N_1194,N_931,N_984);
xor U1195 (N_1195,N_938,N_847);
nor U1196 (N_1196,N_827,N_922);
nor U1197 (N_1197,N_972,N_934);
or U1198 (N_1198,N_846,N_836);
or U1199 (N_1199,N_970,N_878);
nand U1200 (N_1200,N_1006,N_1060);
and U1201 (N_1201,N_1032,N_1184);
or U1202 (N_1202,N_1016,N_1007);
or U1203 (N_1203,N_1104,N_1024);
nor U1204 (N_1204,N_1049,N_1167);
and U1205 (N_1205,N_1005,N_1171);
nand U1206 (N_1206,N_1135,N_1045);
and U1207 (N_1207,N_1132,N_1050);
xor U1208 (N_1208,N_1196,N_1177);
or U1209 (N_1209,N_1084,N_1157);
and U1210 (N_1210,N_1153,N_1080);
nor U1211 (N_1211,N_1047,N_1035);
nor U1212 (N_1212,N_1082,N_1096);
xnor U1213 (N_1213,N_1072,N_1056);
nor U1214 (N_1214,N_1193,N_1166);
nor U1215 (N_1215,N_1009,N_1175);
nand U1216 (N_1216,N_1141,N_1158);
xor U1217 (N_1217,N_1055,N_1123);
nand U1218 (N_1218,N_1041,N_1198);
xnor U1219 (N_1219,N_1105,N_1194);
xnor U1220 (N_1220,N_1090,N_1112);
xnor U1221 (N_1221,N_1183,N_1033);
xnor U1222 (N_1222,N_1074,N_1066);
xor U1223 (N_1223,N_1034,N_1051);
nand U1224 (N_1224,N_1142,N_1162);
nand U1225 (N_1225,N_1190,N_1163);
nor U1226 (N_1226,N_1103,N_1098);
nor U1227 (N_1227,N_1071,N_1111);
xor U1228 (N_1228,N_1092,N_1173);
or U1229 (N_1229,N_1116,N_1180);
and U1230 (N_1230,N_1094,N_1188);
or U1231 (N_1231,N_1021,N_1129);
nand U1232 (N_1232,N_1170,N_1197);
and U1233 (N_1233,N_1078,N_1093);
nor U1234 (N_1234,N_1131,N_1065);
xnor U1235 (N_1235,N_1095,N_1189);
nor U1236 (N_1236,N_1106,N_1037);
nand U1237 (N_1237,N_1185,N_1126);
or U1238 (N_1238,N_1008,N_1086);
nand U1239 (N_1239,N_1079,N_1088);
or U1240 (N_1240,N_1029,N_1022);
or U1241 (N_1241,N_1025,N_1020);
nand U1242 (N_1242,N_1168,N_1182);
nand U1243 (N_1243,N_1097,N_1014);
xnor U1244 (N_1244,N_1109,N_1107);
xor U1245 (N_1245,N_1147,N_1127);
nor U1246 (N_1246,N_1048,N_1039);
xor U1247 (N_1247,N_1091,N_1052);
nor U1248 (N_1248,N_1011,N_1150);
xor U1249 (N_1249,N_1179,N_1159);
or U1250 (N_1250,N_1155,N_1062);
or U1251 (N_1251,N_1192,N_1061);
or U1252 (N_1252,N_1031,N_1070);
and U1253 (N_1253,N_1010,N_1178);
nor U1254 (N_1254,N_1152,N_1114);
nor U1255 (N_1255,N_1156,N_1115);
nor U1256 (N_1256,N_1154,N_1130);
xnor U1257 (N_1257,N_1053,N_1140);
nand U1258 (N_1258,N_1169,N_1017);
nand U1259 (N_1259,N_1172,N_1108);
or U1260 (N_1260,N_1110,N_1139);
nor U1261 (N_1261,N_1145,N_1075);
nor U1262 (N_1262,N_1165,N_1122);
nand U1263 (N_1263,N_1038,N_1143);
or U1264 (N_1264,N_1043,N_1144);
and U1265 (N_1265,N_1125,N_1069);
nor U1266 (N_1266,N_1018,N_1119);
nand U1267 (N_1267,N_1195,N_1004);
and U1268 (N_1268,N_1181,N_1076);
xor U1269 (N_1269,N_1124,N_1089);
and U1270 (N_1270,N_1133,N_1057);
xor U1271 (N_1271,N_1026,N_1067);
and U1272 (N_1272,N_1113,N_1046);
or U1273 (N_1273,N_1015,N_1160);
nand U1274 (N_1274,N_1068,N_1199);
or U1275 (N_1275,N_1013,N_1136);
xor U1276 (N_1276,N_1187,N_1102);
or U1277 (N_1277,N_1118,N_1087);
nor U1278 (N_1278,N_1151,N_1186);
and U1279 (N_1279,N_1027,N_1059);
nor U1280 (N_1280,N_1191,N_1036);
and U1281 (N_1281,N_1019,N_1001);
nor U1282 (N_1282,N_1054,N_1083);
nor U1283 (N_1283,N_1028,N_1012);
or U1284 (N_1284,N_1146,N_1023);
nand U1285 (N_1285,N_1134,N_1044);
xnor U1286 (N_1286,N_1064,N_1085);
nand U1287 (N_1287,N_1137,N_1121);
or U1288 (N_1288,N_1100,N_1058);
nor U1289 (N_1289,N_1128,N_1073);
xnor U1290 (N_1290,N_1120,N_1149);
nand U1291 (N_1291,N_1174,N_1099);
or U1292 (N_1292,N_1040,N_1077);
xor U1293 (N_1293,N_1042,N_1003);
nor U1294 (N_1294,N_1164,N_1101);
xnor U1295 (N_1295,N_1002,N_1081);
xnor U1296 (N_1296,N_1148,N_1176);
xor U1297 (N_1297,N_1063,N_1138);
nand U1298 (N_1298,N_1030,N_1000);
nor U1299 (N_1299,N_1161,N_1117);
nand U1300 (N_1300,N_1111,N_1127);
nor U1301 (N_1301,N_1053,N_1005);
and U1302 (N_1302,N_1132,N_1104);
xnor U1303 (N_1303,N_1120,N_1151);
and U1304 (N_1304,N_1122,N_1011);
and U1305 (N_1305,N_1171,N_1025);
nor U1306 (N_1306,N_1086,N_1117);
xor U1307 (N_1307,N_1195,N_1111);
nor U1308 (N_1308,N_1039,N_1093);
xnor U1309 (N_1309,N_1192,N_1006);
nor U1310 (N_1310,N_1132,N_1171);
or U1311 (N_1311,N_1113,N_1190);
nand U1312 (N_1312,N_1127,N_1176);
nor U1313 (N_1313,N_1131,N_1171);
and U1314 (N_1314,N_1180,N_1159);
or U1315 (N_1315,N_1103,N_1025);
nand U1316 (N_1316,N_1151,N_1117);
nand U1317 (N_1317,N_1087,N_1000);
nor U1318 (N_1318,N_1078,N_1059);
or U1319 (N_1319,N_1130,N_1163);
and U1320 (N_1320,N_1059,N_1170);
nand U1321 (N_1321,N_1057,N_1051);
nor U1322 (N_1322,N_1133,N_1194);
and U1323 (N_1323,N_1006,N_1011);
xnor U1324 (N_1324,N_1022,N_1127);
or U1325 (N_1325,N_1000,N_1180);
nand U1326 (N_1326,N_1157,N_1129);
xnor U1327 (N_1327,N_1110,N_1168);
or U1328 (N_1328,N_1166,N_1160);
and U1329 (N_1329,N_1196,N_1085);
nand U1330 (N_1330,N_1095,N_1083);
xor U1331 (N_1331,N_1062,N_1067);
nor U1332 (N_1332,N_1045,N_1005);
nor U1333 (N_1333,N_1170,N_1191);
xnor U1334 (N_1334,N_1133,N_1073);
nand U1335 (N_1335,N_1021,N_1059);
xnor U1336 (N_1336,N_1052,N_1146);
nand U1337 (N_1337,N_1077,N_1085);
nor U1338 (N_1338,N_1122,N_1089);
xor U1339 (N_1339,N_1166,N_1016);
xnor U1340 (N_1340,N_1190,N_1142);
nand U1341 (N_1341,N_1063,N_1160);
xor U1342 (N_1342,N_1069,N_1164);
nand U1343 (N_1343,N_1155,N_1120);
nand U1344 (N_1344,N_1197,N_1029);
or U1345 (N_1345,N_1186,N_1174);
or U1346 (N_1346,N_1021,N_1155);
nand U1347 (N_1347,N_1131,N_1140);
nor U1348 (N_1348,N_1190,N_1150);
nand U1349 (N_1349,N_1118,N_1101);
or U1350 (N_1350,N_1110,N_1140);
xor U1351 (N_1351,N_1007,N_1086);
and U1352 (N_1352,N_1183,N_1000);
nor U1353 (N_1353,N_1144,N_1057);
or U1354 (N_1354,N_1174,N_1025);
xnor U1355 (N_1355,N_1142,N_1146);
or U1356 (N_1356,N_1000,N_1005);
nor U1357 (N_1357,N_1078,N_1163);
or U1358 (N_1358,N_1037,N_1184);
nor U1359 (N_1359,N_1094,N_1185);
xor U1360 (N_1360,N_1111,N_1070);
nor U1361 (N_1361,N_1144,N_1165);
or U1362 (N_1362,N_1167,N_1101);
nand U1363 (N_1363,N_1094,N_1080);
xor U1364 (N_1364,N_1072,N_1107);
nand U1365 (N_1365,N_1103,N_1044);
and U1366 (N_1366,N_1142,N_1086);
nand U1367 (N_1367,N_1042,N_1073);
xnor U1368 (N_1368,N_1003,N_1024);
or U1369 (N_1369,N_1030,N_1134);
and U1370 (N_1370,N_1125,N_1160);
and U1371 (N_1371,N_1099,N_1070);
xor U1372 (N_1372,N_1129,N_1059);
or U1373 (N_1373,N_1142,N_1193);
nor U1374 (N_1374,N_1184,N_1016);
and U1375 (N_1375,N_1135,N_1079);
nor U1376 (N_1376,N_1149,N_1118);
xor U1377 (N_1377,N_1171,N_1043);
xnor U1378 (N_1378,N_1129,N_1130);
nand U1379 (N_1379,N_1056,N_1167);
nand U1380 (N_1380,N_1053,N_1105);
nor U1381 (N_1381,N_1113,N_1038);
or U1382 (N_1382,N_1109,N_1118);
or U1383 (N_1383,N_1019,N_1087);
nand U1384 (N_1384,N_1130,N_1048);
or U1385 (N_1385,N_1028,N_1143);
xnor U1386 (N_1386,N_1076,N_1104);
nor U1387 (N_1387,N_1173,N_1136);
nor U1388 (N_1388,N_1191,N_1098);
nand U1389 (N_1389,N_1092,N_1141);
xnor U1390 (N_1390,N_1090,N_1047);
nor U1391 (N_1391,N_1052,N_1057);
xor U1392 (N_1392,N_1053,N_1057);
nor U1393 (N_1393,N_1135,N_1056);
or U1394 (N_1394,N_1154,N_1073);
xnor U1395 (N_1395,N_1169,N_1056);
xor U1396 (N_1396,N_1041,N_1137);
and U1397 (N_1397,N_1165,N_1156);
xnor U1398 (N_1398,N_1195,N_1058);
or U1399 (N_1399,N_1079,N_1005);
nand U1400 (N_1400,N_1297,N_1379);
nand U1401 (N_1401,N_1267,N_1207);
nand U1402 (N_1402,N_1331,N_1204);
xor U1403 (N_1403,N_1308,N_1224);
and U1404 (N_1404,N_1388,N_1249);
and U1405 (N_1405,N_1239,N_1387);
nand U1406 (N_1406,N_1385,N_1359);
nand U1407 (N_1407,N_1342,N_1250);
xor U1408 (N_1408,N_1241,N_1231);
xnor U1409 (N_1409,N_1306,N_1268);
and U1410 (N_1410,N_1340,N_1364);
and U1411 (N_1411,N_1339,N_1346);
xor U1412 (N_1412,N_1263,N_1318);
nand U1413 (N_1413,N_1327,N_1301);
and U1414 (N_1414,N_1337,N_1226);
nor U1415 (N_1415,N_1211,N_1215);
nor U1416 (N_1416,N_1252,N_1367);
xnor U1417 (N_1417,N_1278,N_1296);
nand U1418 (N_1418,N_1307,N_1209);
xor U1419 (N_1419,N_1361,N_1245);
nand U1420 (N_1420,N_1377,N_1343);
or U1421 (N_1421,N_1216,N_1279);
or U1422 (N_1422,N_1265,N_1370);
or U1423 (N_1423,N_1376,N_1358);
and U1424 (N_1424,N_1221,N_1356);
nand U1425 (N_1425,N_1257,N_1246);
nor U1426 (N_1426,N_1295,N_1366);
or U1427 (N_1427,N_1371,N_1329);
nand U1428 (N_1428,N_1225,N_1235);
xor U1429 (N_1429,N_1271,N_1372);
nor U1430 (N_1430,N_1321,N_1330);
or U1431 (N_1431,N_1394,N_1270);
nor U1432 (N_1432,N_1254,N_1290);
nand U1433 (N_1433,N_1259,N_1272);
or U1434 (N_1434,N_1368,N_1336);
nand U1435 (N_1435,N_1375,N_1227);
xnor U1436 (N_1436,N_1228,N_1335);
nor U1437 (N_1437,N_1256,N_1242);
or U1438 (N_1438,N_1208,N_1284);
nor U1439 (N_1439,N_1291,N_1381);
and U1440 (N_1440,N_1253,N_1373);
or U1441 (N_1441,N_1386,N_1223);
or U1442 (N_1442,N_1324,N_1300);
nand U1443 (N_1443,N_1354,N_1316);
nand U1444 (N_1444,N_1214,N_1213);
nor U1445 (N_1445,N_1353,N_1383);
and U1446 (N_1446,N_1205,N_1283);
or U1447 (N_1447,N_1389,N_1397);
nand U1448 (N_1448,N_1332,N_1322);
and U1449 (N_1449,N_1251,N_1384);
and U1450 (N_1450,N_1396,N_1392);
nor U1451 (N_1451,N_1304,N_1312);
nand U1452 (N_1452,N_1234,N_1269);
nor U1453 (N_1453,N_1333,N_1277);
xor U1454 (N_1454,N_1286,N_1233);
and U1455 (N_1455,N_1218,N_1317);
or U1456 (N_1456,N_1349,N_1255);
or U1457 (N_1457,N_1276,N_1289);
nor U1458 (N_1458,N_1217,N_1261);
and U1459 (N_1459,N_1369,N_1399);
and U1460 (N_1460,N_1311,N_1391);
nand U1461 (N_1461,N_1288,N_1274);
xnor U1462 (N_1462,N_1260,N_1222);
or U1463 (N_1463,N_1319,N_1344);
xor U1464 (N_1464,N_1320,N_1219);
xor U1465 (N_1465,N_1362,N_1238);
and U1466 (N_1466,N_1293,N_1350);
xor U1467 (N_1467,N_1328,N_1326);
xnor U1468 (N_1468,N_1305,N_1357);
xor U1469 (N_1469,N_1240,N_1285);
xor U1470 (N_1470,N_1315,N_1273);
xor U1471 (N_1471,N_1244,N_1202);
and U1472 (N_1472,N_1264,N_1243);
nor U1473 (N_1473,N_1230,N_1212);
nand U1474 (N_1474,N_1203,N_1236);
and U1475 (N_1475,N_1380,N_1237);
nand U1476 (N_1476,N_1374,N_1341);
or U1477 (N_1477,N_1310,N_1309);
or U1478 (N_1478,N_1355,N_1200);
or U1479 (N_1479,N_1247,N_1314);
and U1480 (N_1480,N_1292,N_1229);
nand U1481 (N_1481,N_1262,N_1348);
and U1482 (N_1482,N_1395,N_1282);
and U1483 (N_1483,N_1302,N_1390);
nand U1484 (N_1484,N_1303,N_1220);
and U1485 (N_1485,N_1325,N_1338);
nand U1486 (N_1486,N_1352,N_1206);
and U1487 (N_1487,N_1398,N_1294);
nor U1488 (N_1488,N_1378,N_1287);
nor U1489 (N_1489,N_1347,N_1248);
xor U1490 (N_1490,N_1201,N_1275);
nand U1491 (N_1491,N_1393,N_1363);
xnor U1492 (N_1492,N_1360,N_1281);
nand U1493 (N_1493,N_1365,N_1382);
and U1494 (N_1494,N_1334,N_1258);
or U1495 (N_1495,N_1351,N_1210);
nand U1496 (N_1496,N_1313,N_1299);
xnor U1497 (N_1497,N_1298,N_1280);
nand U1498 (N_1498,N_1323,N_1232);
nor U1499 (N_1499,N_1266,N_1345);
and U1500 (N_1500,N_1354,N_1251);
or U1501 (N_1501,N_1281,N_1278);
nor U1502 (N_1502,N_1272,N_1364);
and U1503 (N_1503,N_1322,N_1210);
nor U1504 (N_1504,N_1264,N_1325);
xnor U1505 (N_1505,N_1378,N_1264);
or U1506 (N_1506,N_1382,N_1396);
and U1507 (N_1507,N_1339,N_1299);
nand U1508 (N_1508,N_1313,N_1210);
xnor U1509 (N_1509,N_1360,N_1231);
xor U1510 (N_1510,N_1359,N_1323);
nand U1511 (N_1511,N_1304,N_1321);
nor U1512 (N_1512,N_1352,N_1337);
nand U1513 (N_1513,N_1340,N_1380);
and U1514 (N_1514,N_1345,N_1315);
and U1515 (N_1515,N_1277,N_1254);
and U1516 (N_1516,N_1324,N_1326);
or U1517 (N_1517,N_1398,N_1211);
and U1518 (N_1518,N_1205,N_1321);
or U1519 (N_1519,N_1226,N_1344);
nand U1520 (N_1520,N_1391,N_1237);
and U1521 (N_1521,N_1263,N_1205);
and U1522 (N_1522,N_1381,N_1399);
and U1523 (N_1523,N_1253,N_1337);
nor U1524 (N_1524,N_1221,N_1286);
or U1525 (N_1525,N_1261,N_1286);
and U1526 (N_1526,N_1212,N_1386);
xor U1527 (N_1527,N_1360,N_1352);
nand U1528 (N_1528,N_1284,N_1354);
xnor U1529 (N_1529,N_1366,N_1270);
and U1530 (N_1530,N_1253,N_1294);
nor U1531 (N_1531,N_1355,N_1376);
nand U1532 (N_1532,N_1213,N_1395);
xor U1533 (N_1533,N_1311,N_1269);
nor U1534 (N_1534,N_1256,N_1202);
nor U1535 (N_1535,N_1314,N_1287);
and U1536 (N_1536,N_1326,N_1236);
and U1537 (N_1537,N_1326,N_1257);
nand U1538 (N_1538,N_1247,N_1308);
nand U1539 (N_1539,N_1239,N_1229);
and U1540 (N_1540,N_1392,N_1243);
nor U1541 (N_1541,N_1249,N_1218);
nor U1542 (N_1542,N_1266,N_1370);
and U1543 (N_1543,N_1309,N_1362);
and U1544 (N_1544,N_1205,N_1324);
nor U1545 (N_1545,N_1279,N_1215);
nand U1546 (N_1546,N_1319,N_1378);
nor U1547 (N_1547,N_1262,N_1317);
and U1548 (N_1548,N_1257,N_1336);
nand U1549 (N_1549,N_1259,N_1381);
nand U1550 (N_1550,N_1240,N_1385);
or U1551 (N_1551,N_1260,N_1381);
or U1552 (N_1552,N_1216,N_1247);
nor U1553 (N_1553,N_1289,N_1345);
nor U1554 (N_1554,N_1227,N_1326);
and U1555 (N_1555,N_1332,N_1250);
or U1556 (N_1556,N_1252,N_1315);
xnor U1557 (N_1557,N_1382,N_1208);
or U1558 (N_1558,N_1358,N_1205);
and U1559 (N_1559,N_1334,N_1353);
and U1560 (N_1560,N_1276,N_1244);
nor U1561 (N_1561,N_1327,N_1356);
and U1562 (N_1562,N_1384,N_1383);
nor U1563 (N_1563,N_1323,N_1243);
nor U1564 (N_1564,N_1375,N_1300);
nand U1565 (N_1565,N_1210,N_1311);
or U1566 (N_1566,N_1375,N_1382);
nor U1567 (N_1567,N_1330,N_1245);
nand U1568 (N_1568,N_1261,N_1257);
or U1569 (N_1569,N_1250,N_1312);
nor U1570 (N_1570,N_1345,N_1300);
xnor U1571 (N_1571,N_1397,N_1394);
xnor U1572 (N_1572,N_1292,N_1301);
nor U1573 (N_1573,N_1393,N_1376);
or U1574 (N_1574,N_1293,N_1219);
xor U1575 (N_1575,N_1361,N_1321);
nand U1576 (N_1576,N_1362,N_1218);
nor U1577 (N_1577,N_1279,N_1203);
xnor U1578 (N_1578,N_1259,N_1384);
xor U1579 (N_1579,N_1273,N_1349);
and U1580 (N_1580,N_1393,N_1358);
or U1581 (N_1581,N_1354,N_1220);
nand U1582 (N_1582,N_1251,N_1359);
nand U1583 (N_1583,N_1200,N_1331);
xnor U1584 (N_1584,N_1360,N_1285);
nor U1585 (N_1585,N_1317,N_1220);
or U1586 (N_1586,N_1214,N_1208);
nand U1587 (N_1587,N_1252,N_1235);
nor U1588 (N_1588,N_1222,N_1351);
nand U1589 (N_1589,N_1372,N_1383);
and U1590 (N_1590,N_1324,N_1347);
or U1591 (N_1591,N_1216,N_1318);
nand U1592 (N_1592,N_1337,N_1211);
and U1593 (N_1593,N_1375,N_1339);
nand U1594 (N_1594,N_1368,N_1207);
or U1595 (N_1595,N_1256,N_1213);
nor U1596 (N_1596,N_1331,N_1238);
nand U1597 (N_1597,N_1234,N_1384);
nand U1598 (N_1598,N_1308,N_1263);
and U1599 (N_1599,N_1396,N_1366);
and U1600 (N_1600,N_1470,N_1510);
nand U1601 (N_1601,N_1526,N_1557);
nor U1602 (N_1602,N_1535,N_1503);
or U1603 (N_1603,N_1547,N_1409);
nor U1604 (N_1604,N_1499,N_1496);
or U1605 (N_1605,N_1594,N_1536);
nand U1606 (N_1606,N_1491,N_1576);
nor U1607 (N_1607,N_1545,N_1475);
and U1608 (N_1608,N_1456,N_1533);
xnor U1609 (N_1609,N_1513,N_1414);
nand U1610 (N_1610,N_1464,N_1567);
nor U1611 (N_1611,N_1505,N_1445);
nor U1612 (N_1612,N_1479,N_1437);
nor U1613 (N_1613,N_1416,N_1501);
and U1614 (N_1614,N_1467,N_1426);
and U1615 (N_1615,N_1462,N_1570);
xor U1616 (N_1616,N_1530,N_1423);
and U1617 (N_1617,N_1413,N_1419);
or U1618 (N_1618,N_1421,N_1434);
or U1619 (N_1619,N_1585,N_1593);
nor U1620 (N_1620,N_1469,N_1588);
nor U1621 (N_1621,N_1566,N_1439);
nor U1622 (N_1622,N_1506,N_1424);
nand U1623 (N_1623,N_1574,N_1447);
or U1624 (N_1624,N_1402,N_1559);
nor U1625 (N_1625,N_1529,N_1407);
nand U1626 (N_1626,N_1481,N_1569);
or U1627 (N_1627,N_1546,N_1458);
and U1628 (N_1628,N_1441,N_1577);
xnor U1629 (N_1629,N_1583,N_1580);
or U1630 (N_1630,N_1509,N_1524);
nor U1631 (N_1631,N_1400,N_1544);
xnor U1632 (N_1632,N_1488,N_1404);
nor U1633 (N_1633,N_1451,N_1589);
xor U1634 (N_1634,N_1584,N_1568);
nand U1635 (N_1635,N_1512,N_1417);
or U1636 (N_1636,N_1591,N_1579);
xor U1637 (N_1637,N_1477,N_1484);
and U1638 (N_1638,N_1493,N_1438);
xnor U1639 (N_1639,N_1571,N_1540);
nor U1640 (N_1640,N_1595,N_1532);
and U1641 (N_1641,N_1476,N_1539);
xnor U1642 (N_1642,N_1485,N_1587);
or U1643 (N_1643,N_1538,N_1581);
or U1644 (N_1644,N_1582,N_1573);
nand U1645 (N_1645,N_1565,N_1401);
xor U1646 (N_1646,N_1490,N_1541);
or U1647 (N_1647,N_1425,N_1555);
nor U1648 (N_1648,N_1411,N_1598);
nand U1649 (N_1649,N_1422,N_1440);
or U1650 (N_1650,N_1563,N_1410);
xor U1651 (N_1651,N_1516,N_1472);
xnor U1652 (N_1652,N_1432,N_1457);
and U1653 (N_1653,N_1502,N_1537);
nor U1654 (N_1654,N_1596,N_1465);
or U1655 (N_1655,N_1560,N_1406);
xor U1656 (N_1656,N_1519,N_1471);
nand U1657 (N_1657,N_1482,N_1442);
nor U1658 (N_1658,N_1436,N_1507);
or U1659 (N_1659,N_1522,N_1523);
xor U1660 (N_1660,N_1448,N_1599);
nand U1661 (N_1661,N_1578,N_1561);
and U1662 (N_1662,N_1504,N_1500);
or U1663 (N_1663,N_1550,N_1553);
and U1664 (N_1664,N_1558,N_1473);
xnor U1665 (N_1665,N_1549,N_1590);
xor U1666 (N_1666,N_1492,N_1463);
and U1667 (N_1667,N_1444,N_1514);
nand U1668 (N_1668,N_1551,N_1497);
and U1669 (N_1669,N_1433,N_1459);
nor U1670 (N_1670,N_1548,N_1511);
or U1671 (N_1671,N_1486,N_1521);
nand U1672 (N_1672,N_1592,N_1431);
and U1673 (N_1673,N_1468,N_1452);
or U1674 (N_1674,N_1508,N_1427);
xnor U1675 (N_1675,N_1443,N_1498);
or U1676 (N_1676,N_1428,N_1415);
nor U1677 (N_1677,N_1429,N_1487);
and U1678 (N_1678,N_1435,N_1597);
and U1679 (N_1679,N_1575,N_1418);
or U1680 (N_1680,N_1586,N_1495);
nor U1681 (N_1681,N_1543,N_1420);
or U1682 (N_1682,N_1542,N_1518);
nand U1683 (N_1683,N_1527,N_1408);
nor U1684 (N_1684,N_1556,N_1515);
nand U1685 (N_1685,N_1517,N_1572);
nand U1686 (N_1686,N_1534,N_1461);
nand U1687 (N_1687,N_1489,N_1460);
xor U1688 (N_1688,N_1531,N_1455);
xor U1689 (N_1689,N_1474,N_1564);
xnor U1690 (N_1690,N_1446,N_1483);
xor U1691 (N_1691,N_1562,N_1466);
and U1692 (N_1692,N_1454,N_1403);
xnor U1693 (N_1693,N_1525,N_1430);
nor U1694 (N_1694,N_1478,N_1405);
or U1695 (N_1695,N_1450,N_1480);
xor U1696 (N_1696,N_1412,N_1494);
and U1697 (N_1697,N_1552,N_1520);
and U1698 (N_1698,N_1528,N_1449);
xnor U1699 (N_1699,N_1453,N_1554);
xnor U1700 (N_1700,N_1460,N_1471);
nor U1701 (N_1701,N_1475,N_1575);
xnor U1702 (N_1702,N_1594,N_1513);
or U1703 (N_1703,N_1403,N_1591);
xnor U1704 (N_1704,N_1485,N_1410);
and U1705 (N_1705,N_1505,N_1425);
xnor U1706 (N_1706,N_1480,N_1421);
nand U1707 (N_1707,N_1454,N_1546);
nand U1708 (N_1708,N_1545,N_1543);
or U1709 (N_1709,N_1568,N_1459);
nor U1710 (N_1710,N_1545,N_1581);
nor U1711 (N_1711,N_1486,N_1582);
and U1712 (N_1712,N_1550,N_1425);
nor U1713 (N_1713,N_1539,N_1506);
xor U1714 (N_1714,N_1486,N_1493);
nand U1715 (N_1715,N_1442,N_1521);
nand U1716 (N_1716,N_1575,N_1559);
nor U1717 (N_1717,N_1454,N_1561);
nor U1718 (N_1718,N_1409,N_1582);
and U1719 (N_1719,N_1426,N_1401);
xnor U1720 (N_1720,N_1517,N_1511);
nor U1721 (N_1721,N_1570,N_1452);
and U1722 (N_1722,N_1510,N_1591);
or U1723 (N_1723,N_1436,N_1449);
nand U1724 (N_1724,N_1502,N_1487);
nor U1725 (N_1725,N_1525,N_1447);
xnor U1726 (N_1726,N_1562,N_1468);
nand U1727 (N_1727,N_1455,N_1508);
or U1728 (N_1728,N_1593,N_1402);
xnor U1729 (N_1729,N_1448,N_1507);
and U1730 (N_1730,N_1430,N_1528);
nand U1731 (N_1731,N_1420,N_1484);
or U1732 (N_1732,N_1405,N_1567);
and U1733 (N_1733,N_1483,N_1417);
xor U1734 (N_1734,N_1572,N_1456);
xor U1735 (N_1735,N_1427,N_1580);
nor U1736 (N_1736,N_1498,N_1562);
nor U1737 (N_1737,N_1552,N_1464);
or U1738 (N_1738,N_1476,N_1414);
or U1739 (N_1739,N_1475,N_1553);
or U1740 (N_1740,N_1429,N_1566);
and U1741 (N_1741,N_1456,N_1537);
or U1742 (N_1742,N_1536,N_1583);
nor U1743 (N_1743,N_1435,N_1556);
nand U1744 (N_1744,N_1543,N_1519);
xor U1745 (N_1745,N_1545,N_1418);
nand U1746 (N_1746,N_1571,N_1407);
nand U1747 (N_1747,N_1533,N_1526);
nand U1748 (N_1748,N_1506,N_1597);
nor U1749 (N_1749,N_1497,N_1402);
xor U1750 (N_1750,N_1559,N_1482);
nor U1751 (N_1751,N_1441,N_1532);
nand U1752 (N_1752,N_1549,N_1559);
and U1753 (N_1753,N_1445,N_1593);
or U1754 (N_1754,N_1444,N_1482);
xor U1755 (N_1755,N_1498,N_1421);
nor U1756 (N_1756,N_1466,N_1402);
nor U1757 (N_1757,N_1571,N_1528);
or U1758 (N_1758,N_1427,N_1496);
xnor U1759 (N_1759,N_1448,N_1473);
and U1760 (N_1760,N_1540,N_1453);
xnor U1761 (N_1761,N_1504,N_1482);
nor U1762 (N_1762,N_1472,N_1415);
and U1763 (N_1763,N_1468,N_1406);
or U1764 (N_1764,N_1491,N_1549);
and U1765 (N_1765,N_1419,N_1464);
and U1766 (N_1766,N_1565,N_1568);
or U1767 (N_1767,N_1441,N_1479);
xor U1768 (N_1768,N_1449,N_1491);
and U1769 (N_1769,N_1440,N_1543);
and U1770 (N_1770,N_1536,N_1487);
nor U1771 (N_1771,N_1434,N_1568);
nor U1772 (N_1772,N_1596,N_1427);
and U1773 (N_1773,N_1460,N_1588);
and U1774 (N_1774,N_1485,N_1402);
nor U1775 (N_1775,N_1540,N_1593);
or U1776 (N_1776,N_1402,N_1492);
xor U1777 (N_1777,N_1436,N_1495);
or U1778 (N_1778,N_1511,N_1593);
xnor U1779 (N_1779,N_1455,N_1437);
nor U1780 (N_1780,N_1557,N_1509);
nand U1781 (N_1781,N_1436,N_1412);
or U1782 (N_1782,N_1516,N_1502);
nor U1783 (N_1783,N_1536,N_1577);
nand U1784 (N_1784,N_1563,N_1454);
nand U1785 (N_1785,N_1494,N_1418);
nor U1786 (N_1786,N_1560,N_1526);
xor U1787 (N_1787,N_1482,N_1421);
xnor U1788 (N_1788,N_1595,N_1521);
and U1789 (N_1789,N_1567,N_1536);
and U1790 (N_1790,N_1405,N_1470);
nor U1791 (N_1791,N_1577,N_1516);
and U1792 (N_1792,N_1429,N_1579);
nor U1793 (N_1793,N_1448,N_1419);
or U1794 (N_1794,N_1508,N_1509);
nor U1795 (N_1795,N_1511,N_1555);
xnor U1796 (N_1796,N_1426,N_1528);
and U1797 (N_1797,N_1439,N_1537);
or U1798 (N_1798,N_1450,N_1550);
or U1799 (N_1799,N_1558,N_1525);
and U1800 (N_1800,N_1616,N_1701);
nand U1801 (N_1801,N_1796,N_1674);
or U1802 (N_1802,N_1648,N_1798);
nor U1803 (N_1803,N_1668,N_1710);
or U1804 (N_1804,N_1744,N_1765);
and U1805 (N_1805,N_1678,N_1647);
and U1806 (N_1806,N_1649,N_1700);
xor U1807 (N_1807,N_1780,N_1670);
xor U1808 (N_1808,N_1725,N_1611);
or U1809 (N_1809,N_1677,N_1758);
nand U1810 (N_1810,N_1742,N_1608);
nand U1811 (N_1811,N_1759,N_1704);
or U1812 (N_1812,N_1653,N_1644);
and U1813 (N_1813,N_1665,N_1640);
nand U1814 (N_1814,N_1695,N_1694);
and U1815 (N_1815,N_1718,N_1717);
xor U1816 (N_1816,N_1632,N_1779);
nor U1817 (N_1817,N_1620,N_1621);
xnor U1818 (N_1818,N_1757,N_1726);
or U1819 (N_1819,N_1720,N_1722);
nand U1820 (N_1820,N_1797,N_1634);
and U1821 (N_1821,N_1787,N_1724);
and U1822 (N_1822,N_1698,N_1664);
and U1823 (N_1823,N_1773,N_1706);
and U1824 (N_1824,N_1691,N_1771);
and U1825 (N_1825,N_1751,N_1641);
or U1826 (N_1826,N_1754,N_1660);
and U1827 (N_1827,N_1769,N_1713);
nand U1828 (N_1828,N_1659,N_1740);
nand U1829 (N_1829,N_1624,N_1799);
nand U1830 (N_1830,N_1729,N_1623);
or U1831 (N_1831,N_1635,N_1715);
nand U1832 (N_1832,N_1682,N_1708);
or U1833 (N_1833,N_1738,N_1629);
nor U1834 (N_1834,N_1712,N_1709);
nor U1835 (N_1835,N_1749,N_1679);
or U1836 (N_1836,N_1646,N_1636);
nand U1837 (N_1837,N_1723,N_1650);
nand U1838 (N_1838,N_1705,N_1666);
xor U1839 (N_1839,N_1732,N_1685);
nor U1840 (N_1840,N_1673,N_1645);
and U1841 (N_1841,N_1663,N_1711);
xnor U1842 (N_1842,N_1767,N_1760);
xor U1843 (N_1843,N_1631,N_1680);
and U1844 (N_1844,N_1633,N_1794);
xor U1845 (N_1845,N_1747,N_1777);
xnor U1846 (N_1846,N_1768,N_1762);
nand U1847 (N_1847,N_1764,N_1735);
or U1848 (N_1848,N_1693,N_1657);
xor U1849 (N_1849,N_1656,N_1628);
nor U1850 (N_1850,N_1774,N_1783);
xnor U1851 (N_1851,N_1703,N_1688);
and U1852 (N_1852,N_1776,N_1619);
nor U1853 (N_1853,N_1699,N_1627);
nor U1854 (N_1854,N_1612,N_1618);
nand U1855 (N_1855,N_1622,N_1763);
and U1856 (N_1856,N_1692,N_1658);
xnor U1857 (N_1857,N_1790,N_1753);
nand U1858 (N_1858,N_1655,N_1731);
or U1859 (N_1859,N_1637,N_1789);
xor U1860 (N_1860,N_1614,N_1626);
nor U1861 (N_1861,N_1605,N_1756);
and U1862 (N_1862,N_1736,N_1639);
nor U1863 (N_1863,N_1686,N_1721);
or U1864 (N_1864,N_1761,N_1662);
or U1865 (N_1865,N_1625,N_1643);
or U1866 (N_1866,N_1730,N_1707);
or U1867 (N_1867,N_1782,N_1778);
nor U1868 (N_1868,N_1791,N_1697);
xor U1869 (N_1869,N_1788,N_1607);
and U1870 (N_1870,N_1613,N_1781);
nor U1871 (N_1871,N_1746,N_1652);
and U1872 (N_1872,N_1750,N_1690);
and U1873 (N_1873,N_1752,N_1696);
nor U1874 (N_1874,N_1684,N_1786);
or U1875 (N_1875,N_1689,N_1676);
and U1876 (N_1876,N_1719,N_1755);
xnor U1877 (N_1877,N_1667,N_1675);
xnor U1878 (N_1878,N_1714,N_1638);
nand U1879 (N_1879,N_1609,N_1661);
xnor U1880 (N_1880,N_1672,N_1784);
and U1881 (N_1881,N_1785,N_1604);
and U1882 (N_1882,N_1716,N_1792);
or U1883 (N_1883,N_1606,N_1651);
xnor U1884 (N_1884,N_1681,N_1745);
and U1885 (N_1885,N_1770,N_1739);
or U1886 (N_1886,N_1630,N_1728);
and U1887 (N_1887,N_1766,N_1775);
nand U1888 (N_1888,N_1734,N_1748);
or U1889 (N_1889,N_1602,N_1793);
and U1890 (N_1890,N_1601,N_1617);
xnor U1891 (N_1891,N_1702,N_1772);
or U1892 (N_1892,N_1610,N_1727);
xnor U1893 (N_1893,N_1642,N_1733);
xor U1894 (N_1894,N_1741,N_1615);
or U1895 (N_1895,N_1671,N_1600);
or U1896 (N_1896,N_1795,N_1737);
or U1897 (N_1897,N_1603,N_1687);
xnor U1898 (N_1898,N_1683,N_1654);
nor U1899 (N_1899,N_1669,N_1743);
nor U1900 (N_1900,N_1685,N_1726);
xnor U1901 (N_1901,N_1704,N_1771);
or U1902 (N_1902,N_1782,N_1672);
nor U1903 (N_1903,N_1635,N_1694);
or U1904 (N_1904,N_1651,N_1630);
nor U1905 (N_1905,N_1617,N_1671);
nor U1906 (N_1906,N_1659,N_1765);
nor U1907 (N_1907,N_1678,N_1799);
and U1908 (N_1908,N_1685,N_1703);
xnor U1909 (N_1909,N_1782,N_1789);
nor U1910 (N_1910,N_1617,N_1738);
and U1911 (N_1911,N_1607,N_1668);
or U1912 (N_1912,N_1649,N_1660);
nand U1913 (N_1913,N_1761,N_1709);
nand U1914 (N_1914,N_1606,N_1605);
and U1915 (N_1915,N_1792,N_1697);
or U1916 (N_1916,N_1643,N_1613);
or U1917 (N_1917,N_1624,N_1723);
nor U1918 (N_1918,N_1658,N_1728);
nor U1919 (N_1919,N_1644,N_1724);
nor U1920 (N_1920,N_1772,N_1774);
xnor U1921 (N_1921,N_1731,N_1616);
nor U1922 (N_1922,N_1662,N_1673);
nand U1923 (N_1923,N_1747,N_1663);
or U1924 (N_1924,N_1720,N_1699);
xor U1925 (N_1925,N_1798,N_1681);
or U1926 (N_1926,N_1771,N_1785);
nor U1927 (N_1927,N_1662,N_1634);
xnor U1928 (N_1928,N_1770,N_1720);
and U1929 (N_1929,N_1747,N_1762);
nand U1930 (N_1930,N_1744,N_1760);
nand U1931 (N_1931,N_1794,N_1668);
and U1932 (N_1932,N_1791,N_1685);
nor U1933 (N_1933,N_1690,N_1640);
xnor U1934 (N_1934,N_1724,N_1768);
nand U1935 (N_1935,N_1704,N_1670);
or U1936 (N_1936,N_1608,N_1734);
and U1937 (N_1937,N_1744,N_1764);
xnor U1938 (N_1938,N_1668,N_1632);
or U1939 (N_1939,N_1771,N_1769);
and U1940 (N_1940,N_1754,N_1632);
nand U1941 (N_1941,N_1738,N_1693);
xnor U1942 (N_1942,N_1619,N_1798);
and U1943 (N_1943,N_1714,N_1610);
nor U1944 (N_1944,N_1674,N_1612);
nand U1945 (N_1945,N_1678,N_1754);
nor U1946 (N_1946,N_1761,N_1623);
nand U1947 (N_1947,N_1613,N_1688);
and U1948 (N_1948,N_1641,N_1662);
or U1949 (N_1949,N_1689,N_1747);
nand U1950 (N_1950,N_1716,N_1665);
nor U1951 (N_1951,N_1649,N_1735);
nor U1952 (N_1952,N_1709,N_1702);
or U1953 (N_1953,N_1775,N_1669);
nand U1954 (N_1954,N_1614,N_1799);
or U1955 (N_1955,N_1748,N_1704);
nand U1956 (N_1956,N_1659,N_1792);
nor U1957 (N_1957,N_1606,N_1773);
and U1958 (N_1958,N_1681,N_1707);
or U1959 (N_1959,N_1684,N_1626);
and U1960 (N_1960,N_1626,N_1756);
nand U1961 (N_1961,N_1768,N_1657);
and U1962 (N_1962,N_1767,N_1789);
and U1963 (N_1963,N_1774,N_1749);
and U1964 (N_1964,N_1650,N_1684);
xnor U1965 (N_1965,N_1735,N_1626);
and U1966 (N_1966,N_1675,N_1741);
nand U1967 (N_1967,N_1709,N_1767);
and U1968 (N_1968,N_1683,N_1721);
nand U1969 (N_1969,N_1639,N_1649);
xor U1970 (N_1970,N_1727,N_1627);
xor U1971 (N_1971,N_1748,N_1632);
or U1972 (N_1972,N_1658,N_1788);
and U1973 (N_1973,N_1682,N_1666);
nand U1974 (N_1974,N_1751,N_1688);
and U1975 (N_1975,N_1771,N_1753);
and U1976 (N_1976,N_1634,N_1668);
nor U1977 (N_1977,N_1643,N_1671);
and U1978 (N_1978,N_1720,N_1760);
and U1979 (N_1979,N_1686,N_1745);
nand U1980 (N_1980,N_1739,N_1681);
and U1981 (N_1981,N_1699,N_1650);
nand U1982 (N_1982,N_1798,N_1633);
or U1983 (N_1983,N_1604,N_1707);
nand U1984 (N_1984,N_1750,N_1792);
and U1985 (N_1985,N_1686,N_1789);
or U1986 (N_1986,N_1663,N_1652);
nand U1987 (N_1987,N_1677,N_1721);
nor U1988 (N_1988,N_1610,N_1690);
nor U1989 (N_1989,N_1678,N_1640);
nor U1990 (N_1990,N_1669,N_1690);
xnor U1991 (N_1991,N_1768,N_1708);
nand U1992 (N_1992,N_1709,N_1748);
xor U1993 (N_1993,N_1778,N_1629);
xor U1994 (N_1994,N_1702,N_1727);
or U1995 (N_1995,N_1707,N_1688);
or U1996 (N_1996,N_1703,N_1715);
and U1997 (N_1997,N_1695,N_1795);
or U1998 (N_1998,N_1675,N_1799);
and U1999 (N_1999,N_1736,N_1618);
and U2000 (N_2000,N_1938,N_1921);
nand U2001 (N_2001,N_1956,N_1983);
nor U2002 (N_2002,N_1989,N_1904);
or U2003 (N_2003,N_1898,N_1871);
nor U2004 (N_2004,N_1819,N_1912);
nand U2005 (N_2005,N_1852,N_1952);
xnor U2006 (N_2006,N_1829,N_1995);
nand U2007 (N_2007,N_1922,N_1843);
nor U2008 (N_2008,N_1969,N_1932);
nor U2009 (N_2009,N_1907,N_1845);
or U2010 (N_2010,N_1981,N_1985);
nor U2011 (N_2011,N_1901,N_1998);
and U2012 (N_2012,N_1885,N_1838);
xor U2013 (N_2013,N_1880,N_1810);
and U2014 (N_2014,N_1928,N_1870);
nand U2015 (N_2015,N_1973,N_1872);
nor U2016 (N_2016,N_1817,N_1957);
or U2017 (N_2017,N_1818,N_1833);
or U2018 (N_2018,N_1860,N_1888);
or U2019 (N_2019,N_1862,N_1849);
xnor U2020 (N_2020,N_1946,N_1944);
nor U2021 (N_2021,N_1881,N_1966);
nor U2022 (N_2022,N_1903,N_1876);
nand U2023 (N_2023,N_1850,N_1902);
and U2024 (N_2024,N_1964,N_1972);
nand U2025 (N_2025,N_1979,N_1939);
xor U2026 (N_2026,N_1865,N_1851);
and U2027 (N_2027,N_1925,N_1929);
or U2028 (N_2028,N_1858,N_1855);
xnor U2029 (N_2029,N_1967,N_1968);
nand U2030 (N_2030,N_1815,N_1836);
nor U2031 (N_2031,N_1937,N_1971);
or U2032 (N_2032,N_1897,N_1941);
nand U2033 (N_2033,N_1835,N_1878);
nand U2034 (N_2034,N_1824,N_1958);
or U2035 (N_2035,N_1831,N_1820);
nand U2036 (N_2036,N_1804,N_1954);
xor U2037 (N_2037,N_1884,N_1890);
nand U2038 (N_2038,N_1891,N_1924);
nand U2039 (N_2039,N_1866,N_1991);
nor U2040 (N_2040,N_1943,N_1935);
nor U2041 (N_2041,N_1899,N_1803);
xnor U2042 (N_2042,N_1893,N_1854);
nand U2043 (N_2043,N_1977,N_1993);
nor U2044 (N_2044,N_1868,N_1988);
nor U2045 (N_2045,N_1877,N_1900);
nand U2046 (N_2046,N_1840,N_1814);
nand U2047 (N_2047,N_1959,N_1914);
nor U2048 (N_2048,N_1828,N_1913);
nand U2049 (N_2049,N_1951,N_1896);
and U2050 (N_2050,N_1895,N_1978);
nand U2051 (N_2051,N_1984,N_1825);
nor U2052 (N_2052,N_1839,N_1867);
or U2053 (N_2053,N_1832,N_1970);
nor U2054 (N_2054,N_1837,N_1961);
xor U2055 (N_2055,N_1926,N_1962);
xnor U2056 (N_2056,N_1936,N_1864);
nor U2057 (N_2057,N_1945,N_1997);
or U2058 (N_2058,N_1887,N_1942);
xor U2059 (N_2059,N_1992,N_1923);
or U2060 (N_2060,N_1933,N_1996);
and U2061 (N_2061,N_1982,N_1947);
or U2062 (N_2062,N_1809,N_1950);
xnor U2063 (N_2063,N_1861,N_1813);
or U2064 (N_2064,N_1812,N_1910);
xor U2065 (N_2065,N_1986,N_1976);
and U2066 (N_2066,N_1990,N_1919);
or U2067 (N_2067,N_1800,N_1894);
or U2068 (N_2068,N_1807,N_1863);
and U2069 (N_2069,N_1955,N_1987);
or U2070 (N_2070,N_1806,N_1816);
nor U2071 (N_2071,N_1875,N_1874);
nor U2072 (N_2072,N_1930,N_1916);
xnor U2073 (N_2073,N_1869,N_1911);
xor U2074 (N_2074,N_1980,N_1802);
xnor U2075 (N_2075,N_1975,N_1827);
and U2076 (N_2076,N_1920,N_1886);
or U2077 (N_2077,N_1889,N_1953);
nand U2078 (N_2078,N_1841,N_1965);
or U2079 (N_2079,N_1892,N_1844);
and U2080 (N_2080,N_1801,N_1915);
nor U2081 (N_2081,N_1808,N_1856);
xor U2082 (N_2082,N_1908,N_1882);
nand U2083 (N_2083,N_1927,N_1948);
xor U2084 (N_2084,N_1859,N_1918);
xnor U2085 (N_2085,N_1905,N_1842);
nand U2086 (N_2086,N_1879,N_1909);
xor U2087 (N_2087,N_1805,N_1846);
nand U2088 (N_2088,N_1940,N_1906);
or U2089 (N_2089,N_1974,N_1917);
xnor U2090 (N_2090,N_1960,N_1873);
nand U2091 (N_2091,N_1949,N_1883);
and U2092 (N_2092,N_1963,N_1994);
nand U2093 (N_2093,N_1822,N_1853);
xor U2094 (N_2094,N_1821,N_1857);
nor U2095 (N_2095,N_1848,N_1934);
nand U2096 (N_2096,N_1826,N_1811);
and U2097 (N_2097,N_1999,N_1834);
or U2098 (N_2098,N_1823,N_1830);
nand U2099 (N_2099,N_1931,N_1847);
nand U2100 (N_2100,N_1856,N_1965);
and U2101 (N_2101,N_1897,N_1823);
and U2102 (N_2102,N_1970,N_1980);
and U2103 (N_2103,N_1899,N_1954);
nand U2104 (N_2104,N_1826,N_1878);
nor U2105 (N_2105,N_1931,N_1930);
xor U2106 (N_2106,N_1901,N_1836);
xnor U2107 (N_2107,N_1986,N_1844);
and U2108 (N_2108,N_1856,N_1855);
or U2109 (N_2109,N_1923,N_1852);
or U2110 (N_2110,N_1804,N_1842);
xor U2111 (N_2111,N_1825,N_1806);
and U2112 (N_2112,N_1829,N_1863);
and U2113 (N_2113,N_1908,N_1973);
and U2114 (N_2114,N_1812,N_1911);
and U2115 (N_2115,N_1960,N_1949);
or U2116 (N_2116,N_1839,N_1921);
xor U2117 (N_2117,N_1862,N_1879);
nor U2118 (N_2118,N_1873,N_1953);
nand U2119 (N_2119,N_1966,N_1873);
xnor U2120 (N_2120,N_1904,N_1889);
nand U2121 (N_2121,N_1866,N_1989);
or U2122 (N_2122,N_1909,N_1947);
xor U2123 (N_2123,N_1995,N_1917);
nand U2124 (N_2124,N_1945,N_1958);
and U2125 (N_2125,N_1894,N_1879);
nand U2126 (N_2126,N_1911,N_1848);
and U2127 (N_2127,N_1938,N_1831);
or U2128 (N_2128,N_1881,N_1834);
or U2129 (N_2129,N_1929,N_1830);
and U2130 (N_2130,N_1846,N_1912);
nor U2131 (N_2131,N_1937,N_1891);
nor U2132 (N_2132,N_1948,N_1806);
xnor U2133 (N_2133,N_1973,N_1982);
and U2134 (N_2134,N_1962,N_1979);
or U2135 (N_2135,N_1921,N_1900);
nand U2136 (N_2136,N_1898,N_1896);
xor U2137 (N_2137,N_1944,N_1954);
nand U2138 (N_2138,N_1802,N_1981);
xnor U2139 (N_2139,N_1912,N_1870);
nor U2140 (N_2140,N_1852,N_1994);
or U2141 (N_2141,N_1937,N_1962);
or U2142 (N_2142,N_1942,N_1862);
or U2143 (N_2143,N_1872,N_1890);
nor U2144 (N_2144,N_1813,N_1881);
xor U2145 (N_2145,N_1827,N_1836);
xnor U2146 (N_2146,N_1805,N_1921);
xor U2147 (N_2147,N_1810,N_1922);
nand U2148 (N_2148,N_1941,N_1810);
xnor U2149 (N_2149,N_1837,N_1883);
nor U2150 (N_2150,N_1954,N_1828);
nor U2151 (N_2151,N_1969,N_1808);
xnor U2152 (N_2152,N_1890,N_1887);
or U2153 (N_2153,N_1933,N_1859);
xor U2154 (N_2154,N_1864,N_1918);
nor U2155 (N_2155,N_1984,N_1804);
xnor U2156 (N_2156,N_1829,N_1908);
xnor U2157 (N_2157,N_1918,N_1915);
or U2158 (N_2158,N_1976,N_1967);
nor U2159 (N_2159,N_1946,N_1965);
or U2160 (N_2160,N_1811,N_1926);
xnor U2161 (N_2161,N_1891,N_1863);
nand U2162 (N_2162,N_1989,N_1945);
xnor U2163 (N_2163,N_1959,N_1965);
nand U2164 (N_2164,N_1967,N_1830);
and U2165 (N_2165,N_1994,N_1910);
and U2166 (N_2166,N_1842,N_1952);
nand U2167 (N_2167,N_1865,N_1962);
xnor U2168 (N_2168,N_1874,N_1984);
nand U2169 (N_2169,N_1946,N_1995);
xor U2170 (N_2170,N_1856,N_1990);
nor U2171 (N_2171,N_1942,N_1840);
nand U2172 (N_2172,N_1947,N_1923);
xor U2173 (N_2173,N_1889,N_1940);
nor U2174 (N_2174,N_1909,N_1829);
nand U2175 (N_2175,N_1989,N_1997);
nand U2176 (N_2176,N_1937,N_1857);
nor U2177 (N_2177,N_1906,N_1953);
xnor U2178 (N_2178,N_1928,N_1882);
and U2179 (N_2179,N_1855,N_1828);
or U2180 (N_2180,N_1888,N_1810);
xnor U2181 (N_2181,N_1810,N_1860);
nand U2182 (N_2182,N_1911,N_1975);
nand U2183 (N_2183,N_1867,N_1924);
nand U2184 (N_2184,N_1882,N_1910);
nand U2185 (N_2185,N_1867,N_1909);
or U2186 (N_2186,N_1924,N_1996);
or U2187 (N_2187,N_1937,N_1920);
nor U2188 (N_2188,N_1808,N_1924);
or U2189 (N_2189,N_1868,N_1961);
nor U2190 (N_2190,N_1893,N_1981);
nand U2191 (N_2191,N_1872,N_1908);
nor U2192 (N_2192,N_1930,N_1836);
and U2193 (N_2193,N_1967,N_1913);
nand U2194 (N_2194,N_1956,N_1870);
nand U2195 (N_2195,N_1884,N_1851);
and U2196 (N_2196,N_1924,N_1944);
or U2197 (N_2197,N_1995,N_1955);
nand U2198 (N_2198,N_1893,N_1882);
nand U2199 (N_2199,N_1921,N_1888);
and U2200 (N_2200,N_2105,N_2061);
or U2201 (N_2201,N_2124,N_2006);
xnor U2202 (N_2202,N_2140,N_2062);
nand U2203 (N_2203,N_2111,N_2154);
and U2204 (N_2204,N_2018,N_2136);
nand U2205 (N_2205,N_2187,N_2005);
or U2206 (N_2206,N_2102,N_2121);
or U2207 (N_2207,N_2037,N_2001);
xor U2208 (N_2208,N_2125,N_2057);
nor U2209 (N_2209,N_2151,N_2063);
xor U2210 (N_2210,N_2137,N_2119);
or U2211 (N_2211,N_2100,N_2010);
and U2212 (N_2212,N_2107,N_2184);
xnor U2213 (N_2213,N_2157,N_2149);
nor U2214 (N_2214,N_2017,N_2066);
or U2215 (N_2215,N_2168,N_2008);
or U2216 (N_2216,N_2013,N_2040);
and U2217 (N_2217,N_2174,N_2038);
or U2218 (N_2218,N_2036,N_2128);
or U2219 (N_2219,N_2020,N_2082);
nand U2220 (N_2220,N_2050,N_2192);
or U2221 (N_2221,N_2004,N_2025);
and U2222 (N_2222,N_2009,N_2182);
or U2223 (N_2223,N_2019,N_2074);
xor U2224 (N_2224,N_2029,N_2052);
and U2225 (N_2225,N_2164,N_2094);
or U2226 (N_2226,N_2188,N_2172);
or U2227 (N_2227,N_2103,N_2030);
or U2228 (N_2228,N_2167,N_2197);
and U2229 (N_2229,N_2166,N_2110);
and U2230 (N_2230,N_2117,N_2126);
xnor U2231 (N_2231,N_2022,N_2012);
and U2232 (N_2232,N_2088,N_2002);
nand U2233 (N_2233,N_2053,N_2073);
or U2234 (N_2234,N_2090,N_2056);
nand U2235 (N_2235,N_2033,N_2047);
nor U2236 (N_2236,N_2113,N_2060);
nand U2237 (N_2237,N_2087,N_2135);
and U2238 (N_2238,N_2162,N_2122);
or U2239 (N_2239,N_2044,N_2078);
nor U2240 (N_2240,N_2127,N_2046);
xor U2241 (N_2241,N_2141,N_2014);
nand U2242 (N_2242,N_2075,N_2180);
and U2243 (N_2243,N_2028,N_2130);
xor U2244 (N_2244,N_2059,N_2065);
nor U2245 (N_2245,N_2106,N_2067);
and U2246 (N_2246,N_2003,N_2072);
nand U2247 (N_2247,N_2143,N_2134);
and U2248 (N_2248,N_2027,N_2173);
nand U2249 (N_2249,N_2041,N_2161);
nor U2250 (N_2250,N_2007,N_2069);
or U2251 (N_2251,N_2181,N_2015);
and U2252 (N_2252,N_2043,N_2186);
or U2253 (N_2253,N_2064,N_2079);
or U2254 (N_2254,N_2077,N_2175);
or U2255 (N_2255,N_2190,N_2123);
or U2256 (N_2256,N_2032,N_2096);
nand U2257 (N_2257,N_2058,N_2092);
nand U2258 (N_2258,N_2031,N_2158);
nor U2259 (N_2259,N_2035,N_2120);
nand U2260 (N_2260,N_2114,N_2146);
and U2261 (N_2261,N_2112,N_2144);
or U2262 (N_2262,N_2076,N_2039);
nor U2263 (N_2263,N_2115,N_2138);
nand U2264 (N_2264,N_2133,N_2084);
or U2265 (N_2265,N_2150,N_2196);
xor U2266 (N_2266,N_2101,N_2045);
and U2267 (N_2267,N_2142,N_2199);
nor U2268 (N_2268,N_2054,N_2116);
or U2269 (N_2269,N_2023,N_2071);
xnor U2270 (N_2270,N_2086,N_2178);
xor U2271 (N_2271,N_2093,N_2129);
nand U2272 (N_2272,N_2083,N_2159);
xor U2273 (N_2273,N_2155,N_2185);
nand U2274 (N_2274,N_2169,N_2000);
and U2275 (N_2275,N_2021,N_2177);
and U2276 (N_2276,N_2160,N_2026);
or U2277 (N_2277,N_2194,N_2183);
nor U2278 (N_2278,N_2132,N_2156);
nand U2279 (N_2279,N_2070,N_2034);
or U2280 (N_2280,N_2195,N_2108);
and U2281 (N_2281,N_2176,N_2109);
nor U2282 (N_2282,N_2189,N_2049);
nor U2283 (N_2283,N_2171,N_2095);
xor U2284 (N_2284,N_2068,N_2011);
or U2285 (N_2285,N_2147,N_2016);
nor U2286 (N_2286,N_2193,N_2145);
or U2287 (N_2287,N_2048,N_2080);
or U2288 (N_2288,N_2153,N_2165);
and U2289 (N_2289,N_2152,N_2085);
or U2290 (N_2290,N_2148,N_2091);
xor U2291 (N_2291,N_2179,N_2131);
and U2292 (N_2292,N_2097,N_2139);
nand U2293 (N_2293,N_2163,N_2099);
nand U2294 (N_2294,N_2198,N_2170);
nand U2295 (N_2295,N_2081,N_2051);
nand U2296 (N_2296,N_2042,N_2098);
and U2297 (N_2297,N_2024,N_2055);
xor U2298 (N_2298,N_2191,N_2118);
and U2299 (N_2299,N_2089,N_2104);
or U2300 (N_2300,N_2077,N_2051);
nand U2301 (N_2301,N_2119,N_2103);
and U2302 (N_2302,N_2185,N_2011);
nand U2303 (N_2303,N_2114,N_2162);
xor U2304 (N_2304,N_2083,N_2165);
xor U2305 (N_2305,N_2094,N_2149);
nand U2306 (N_2306,N_2192,N_2162);
nand U2307 (N_2307,N_2106,N_2085);
nand U2308 (N_2308,N_2080,N_2065);
and U2309 (N_2309,N_2073,N_2138);
and U2310 (N_2310,N_2132,N_2168);
and U2311 (N_2311,N_2002,N_2199);
xnor U2312 (N_2312,N_2157,N_2002);
and U2313 (N_2313,N_2043,N_2113);
nand U2314 (N_2314,N_2066,N_2044);
or U2315 (N_2315,N_2020,N_2155);
nand U2316 (N_2316,N_2009,N_2117);
nand U2317 (N_2317,N_2075,N_2020);
or U2318 (N_2318,N_2171,N_2062);
or U2319 (N_2319,N_2013,N_2050);
or U2320 (N_2320,N_2051,N_2069);
or U2321 (N_2321,N_2016,N_2104);
xnor U2322 (N_2322,N_2060,N_2126);
and U2323 (N_2323,N_2135,N_2066);
or U2324 (N_2324,N_2148,N_2161);
or U2325 (N_2325,N_2195,N_2157);
or U2326 (N_2326,N_2118,N_2070);
nor U2327 (N_2327,N_2088,N_2124);
nand U2328 (N_2328,N_2058,N_2129);
nor U2329 (N_2329,N_2074,N_2123);
or U2330 (N_2330,N_2168,N_2119);
and U2331 (N_2331,N_2123,N_2050);
nor U2332 (N_2332,N_2031,N_2100);
or U2333 (N_2333,N_2004,N_2098);
nor U2334 (N_2334,N_2157,N_2186);
nor U2335 (N_2335,N_2049,N_2007);
xnor U2336 (N_2336,N_2196,N_2038);
nor U2337 (N_2337,N_2181,N_2143);
nor U2338 (N_2338,N_2188,N_2005);
xor U2339 (N_2339,N_2122,N_2075);
nand U2340 (N_2340,N_2160,N_2141);
xor U2341 (N_2341,N_2048,N_2006);
xor U2342 (N_2342,N_2135,N_2093);
or U2343 (N_2343,N_2035,N_2178);
nand U2344 (N_2344,N_2190,N_2079);
nor U2345 (N_2345,N_2186,N_2093);
nor U2346 (N_2346,N_2175,N_2107);
nor U2347 (N_2347,N_2042,N_2172);
nand U2348 (N_2348,N_2107,N_2173);
xnor U2349 (N_2349,N_2091,N_2177);
or U2350 (N_2350,N_2080,N_2068);
nor U2351 (N_2351,N_2145,N_2050);
nand U2352 (N_2352,N_2199,N_2026);
nand U2353 (N_2353,N_2012,N_2119);
or U2354 (N_2354,N_2133,N_2132);
or U2355 (N_2355,N_2197,N_2073);
xnor U2356 (N_2356,N_2087,N_2122);
xor U2357 (N_2357,N_2173,N_2183);
xnor U2358 (N_2358,N_2170,N_2141);
nand U2359 (N_2359,N_2045,N_2025);
or U2360 (N_2360,N_2174,N_2025);
or U2361 (N_2361,N_2143,N_2123);
nor U2362 (N_2362,N_2152,N_2194);
and U2363 (N_2363,N_2143,N_2161);
and U2364 (N_2364,N_2053,N_2036);
and U2365 (N_2365,N_2170,N_2059);
or U2366 (N_2366,N_2080,N_2165);
or U2367 (N_2367,N_2094,N_2089);
nand U2368 (N_2368,N_2158,N_2049);
xor U2369 (N_2369,N_2196,N_2189);
or U2370 (N_2370,N_2177,N_2034);
or U2371 (N_2371,N_2113,N_2064);
xnor U2372 (N_2372,N_2164,N_2061);
and U2373 (N_2373,N_2055,N_2064);
nand U2374 (N_2374,N_2060,N_2027);
and U2375 (N_2375,N_2022,N_2006);
nand U2376 (N_2376,N_2114,N_2177);
nand U2377 (N_2377,N_2151,N_2030);
or U2378 (N_2378,N_2144,N_2013);
and U2379 (N_2379,N_2049,N_2043);
nor U2380 (N_2380,N_2033,N_2133);
and U2381 (N_2381,N_2148,N_2037);
or U2382 (N_2382,N_2070,N_2042);
or U2383 (N_2383,N_2180,N_2002);
nand U2384 (N_2384,N_2180,N_2136);
xor U2385 (N_2385,N_2166,N_2007);
xnor U2386 (N_2386,N_2130,N_2067);
or U2387 (N_2387,N_2057,N_2028);
or U2388 (N_2388,N_2009,N_2151);
and U2389 (N_2389,N_2027,N_2158);
xnor U2390 (N_2390,N_2103,N_2004);
and U2391 (N_2391,N_2086,N_2198);
nor U2392 (N_2392,N_2000,N_2002);
or U2393 (N_2393,N_2073,N_2021);
and U2394 (N_2394,N_2178,N_2090);
nand U2395 (N_2395,N_2071,N_2146);
nand U2396 (N_2396,N_2093,N_2078);
nand U2397 (N_2397,N_2106,N_2081);
nor U2398 (N_2398,N_2123,N_2002);
xnor U2399 (N_2399,N_2087,N_2093);
xnor U2400 (N_2400,N_2292,N_2249);
xnor U2401 (N_2401,N_2269,N_2299);
nand U2402 (N_2402,N_2386,N_2314);
nor U2403 (N_2403,N_2381,N_2380);
and U2404 (N_2404,N_2224,N_2354);
and U2405 (N_2405,N_2235,N_2345);
nor U2406 (N_2406,N_2279,N_2245);
nand U2407 (N_2407,N_2286,N_2347);
and U2408 (N_2408,N_2255,N_2216);
or U2409 (N_2409,N_2395,N_2204);
or U2410 (N_2410,N_2304,N_2302);
or U2411 (N_2411,N_2202,N_2376);
nand U2412 (N_2412,N_2260,N_2282);
nand U2413 (N_2413,N_2221,N_2271);
or U2414 (N_2414,N_2336,N_2341);
and U2415 (N_2415,N_2277,N_2384);
and U2416 (N_2416,N_2243,N_2268);
nor U2417 (N_2417,N_2360,N_2306);
and U2418 (N_2418,N_2212,N_2311);
or U2419 (N_2419,N_2333,N_2315);
xor U2420 (N_2420,N_2291,N_2200);
xor U2421 (N_2421,N_2280,N_2208);
and U2422 (N_2422,N_2273,N_2262);
xnor U2423 (N_2423,N_2377,N_2364);
nor U2424 (N_2424,N_2305,N_2389);
and U2425 (N_2425,N_2206,N_2267);
nand U2426 (N_2426,N_2371,N_2394);
nand U2427 (N_2427,N_2331,N_2391);
and U2428 (N_2428,N_2214,N_2293);
and U2429 (N_2429,N_2372,N_2387);
or U2430 (N_2430,N_2213,N_2242);
and U2431 (N_2431,N_2309,N_2328);
xnor U2432 (N_2432,N_2295,N_2256);
nor U2433 (N_2433,N_2397,N_2298);
and U2434 (N_2434,N_2303,N_2365);
nand U2435 (N_2435,N_2248,N_2219);
xnor U2436 (N_2436,N_2337,N_2378);
or U2437 (N_2437,N_2375,N_2253);
nor U2438 (N_2438,N_2247,N_2393);
and U2439 (N_2439,N_2319,N_2390);
nand U2440 (N_2440,N_2398,N_2399);
xnor U2441 (N_2441,N_2234,N_2223);
or U2442 (N_2442,N_2258,N_2366);
and U2443 (N_2443,N_2294,N_2263);
nand U2444 (N_2444,N_2322,N_2355);
nor U2445 (N_2445,N_2266,N_2307);
or U2446 (N_2446,N_2257,N_2382);
xor U2447 (N_2447,N_2203,N_2343);
and U2448 (N_2448,N_2209,N_2236);
nor U2449 (N_2449,N_2250,N_2350);
or U2450 (N_2450,N_2321,N_2351);
xnor U2451 (N_2451,N_2251,N_2392);
nand U2452 (N_2452,N_2228,N_2312);
nor U2453 (N_2453,N_2275,N_2231);
nand U2454 (N_2454,N_2361,N_2278);
nand U2455 (N_2455,N_2334,N_2323);
nand U2456 (N_2456,N_2348,N_2296);
xnor U2457 (N_2457,N_2356,N_2207);
nand U2458 (N_2458,N_2383,N_2264);
nand U2459 (N_2459,N_2211,N_2210);
nand U2460 (N_2460,N_2324,N_2344);
and U2461 (N_2461,N_2338,N_2274);
or U2462 (N_2462,N_2201,N_2325);
xor U2463 (N_2463,N_2339,N_2396);
nor U2464 (N_2464,N_2342,N_2352);
and U2465 (N_2465,N_2230,N_2297);
or U2466 (N_2466,N_2374,N_2363);
xnor U2467 (N_2467,N_2388,N_2222);
or U2468 (N_2468,N_2288,N_2335);
or U2469 (N_2469,N_2300,N_2310);
xnor U2470 (N_2470,N_2327,N_2357);
or U2471 (N_2471,N_2346,N_2238);
or U2472 (N_2472,N_2358,N_2227);
nand U2473 (N_2473,N_2270,N_2320);
nor U2474 (N_2474,N_2215,N_2233);
or U2475 (N_2475,N_2349,N_2259);
nor U2476 (N_2476,N_2285,N_2362);
xnor U2477 (N_2477,N_2217,N_2340);
nor U2478 (N_2478,N_2287,N_2284);
xnor U2479 (N_2479,N_2289,N_2373);
xor U2480 (N_2480,N_2254,N_2316);
nand U2481 (N_2481,N_2281,N_2244);
nand U2482 (N_2482,N_2226,N_2276);
nand U2483 (N_2483,N_2218,N_2290);
and U2484 (N_2484,N_2308,N_2265);
xnor U2485 (N_2485,N_2369,N_2370);
nor U2486 (N_2486,N_2329,N_2229);
or U2487 (N_2487,N_2317,N_2367);
and U2488 (N_2488,N_2205,N_2232);
nor U2489 (N_2489,N_2246,N_2313);
xnor U2490 (N_2490,N_2359,N_2237);
xor U2491 (N_2491,N_2220,N_2239);
or U2492 (N_2492,N_2368,N_2252);
or U2493 (N_2493,N_2225,N_2261);
nand U2494 (N_2494,N_2385,N_2301);
and U2495 (N_2495,N_2353,N_2326);
nand U2496 (N_2496,N_2330,N_2379);
nand U2497 (N_2497,N_2332,N_2318);
nand U2498 (N_2498,N_2240,N_2283);
xnor U2499 (N_2499,N_2272,N_2241);
xnor U2500 (N_2500,N_2211,N_2292);
or U2501 (N_2501,N_2385,N_2237);
and U2502 (N_2502,N_2390,N_2291);
nor U2503 (N_2503,N_2327,N_2263);
nand U2504 (N_2504,N_2239,N_2277);
or U2505 (N_2505,N_2279,N_2302);
and U2506 (N_2506,N_2373,N_2302);
nand U2507 (N_2507,N_2210,N_2284);
and U2508 (N_2508,N_2396,N_2290);
xor U2509 (N_2509,N_2280,N_2291);
nand U2510 (N_2510,N_2314,N_2263);
or U2511 (N_2511,N_2225,N_2296);
xnor U2512 (N_2512,N_2381,N_2229);
nand U2513 (N_2513,N_2339,N_2241);
xor U2514 (N_2514,N_2293,N_2281);
and U2515 (N_2515,N_2301,N_2302);
xor U2516 (N_2516,N_2215,N_2256);
or U2517 (N_2517,N_2367,N_2336);
nand U2518 (N_2518,N_2257,N_2330);
or U2519 (N_2519,N_2275,N_2274);
nor U2520 (N_2520,N_2290,N_2255);
nand U2521 (N_2521,N_2398,N_2308);
or U2522 (N_2522,N_2386,N_2383);
nor U2523 (N_2523,N_2335,N_2327);
xor U2524 (N_2524,N_2215,N_2318);
xor U2525 (N_2525,N_2205,N_2242);
or U2526 (N_2526,N_2375,N_2252);
or U2527 (N_2527,N_2365,N_2289);
or U2528 (N_2528,N_2272,N_2215);
xnor U2529 (N_2529,N_2279,N_2291);
nor U2530 (N_2530,N_2224,N_2275);
xor U2531 (N_2531,N_2348,N_2228);
nand U2532 (N_2532,N_2227,N_2205);
xor U2533 (N_2533,N_2240,N_2224);
nand U2534 (N_2534,N_2346,N_2294);
nor U2535 (N_2535,N_2348,N_2329);
xor U2536 (N_2536,N_2204,N_2229);
xor U2537 (N_2537,N_2210,N_2360);
nor U2538 (N_2538,N_2304,N_2266);
or U2539 (N_2539,N_2207,N_2249);
nand U2540 (N_2540,N_2363,N_2335);
nor U2541 (N_2541,N_2269,N_2200);
or U2542 (N_2542,N_2378,N_2374);
or U2543 (N_2543,N_2358,N_2280);
or U2544 (N_2544,N_2306,N_2243);
xor U2545 (N_2545,N_2388,N_2313);
xor U2546 (N_2546,N_2242,N_2327);
nor U2547 (N_2547,N_2358,N_2261);
xnor U2548 (N_2548,N_2309,N_2381);
nand U2549 (N_2549,N_2237,N_2396);
xnor U2550 (N_2550,N_2322,N_2358);
nor U2551 (N_2551,N_2351,N_2265);
or U2552 (N_2552,N_2209,N_2366);
nor U2553 (N_2553,N_2327,N_2366);
nand U2554 (N_2554,N_2297,N_2321);
and U2555 (N_2555,N_2244,N_2374);
or U2556 (N_2556,N_2241,N_2360);
nand U2557 (N_2557,N_2286,N_2241);
and U2558 (N_2558,N_2366,N_2359);
nor U2559 (N_2559,N_2375,N_2347);
xnor U2560 (N_2560,N_2344,N_2293);
xor U2561 (N_2561,N_2324,N_2338);
nand U2562 (N_2562,N_2218,N_2388);
or U2563 (N_2563,N_2289,N_2360);
and U2564 (N_2564,N_2316,N_2326);
and U2565 (N_2565,N_2291,N_2357);
or U2566 (N_2566,N_2206,N_2349);
and U2567 (N_2567,N_2283,N_2290);
xnor U2568 (N_2568,N_2327,N_2362);
nand U2569 (N_2569,N_2298,N_2256);
xor U2570 (N_2570,N_2363,N_2302);
and U2571 (N_2571,N_2237,N_2296);
nor U2572 (N_2572,N_2246,N_2324);
nor U2573 (N_2573,N_2343,N_2380);
or U2574 (N_2574,N_2263,N_2366);
xor U2575 (N_2575,N_2368,N_2339);
nand U2576 (N_2576,N_2223,N_2210);
or U2577 (N_2577,N_2221,N_2373);
nor U2578 (N_2578,N_2388,N_2204);
nand U2579 (N_2579,N_2318,N_2274);
nor U2580 (N_2580,N_2379,N_2369);
or U2581 (N_2581,N_2387,N_2257);
xnor U2582 (N_2582,N_2369,N_2328);
nor U2583 (N_2583,N_2219,N_2202);
xor U2584 (N_2584,N_2351,N_2245);
nand U2585 (N_2585,N_2397,N_2294);
or U2586 (N_2586,N_2253,N_2249);
xor U2587 (N_2587,N_2308,N_2279);
nor U2588 (N_2588,N_2240,N_2249);
xor U2589 (N_2589,N_2238,N_2244);
xnor U2590 (N_2590,N_2305,N_2393);
nor U2591 (N_2591,N_2391,N_2263);
xor U2592 (N_2592,N_2342,N_2276);
and U2593 (N_2593,N_2340,N_2387);
xor U2594 (N_2594,N_2370,N_2215);
or U2595 (N_2595,N_2256,N_2293);
or U2596 (N_2596,N_2256,N_2317);
or U2597 (N_2597,N_2295,N_2211);
nor U2598 (N_2598,N_2372,N_2377);
and U2599 (N_2599,N_2377,N_2232);
and U2600 (N_2600,N_2586,N_2526);
nor U2601 (N_2601,N_2450,N_2441);
or U2602 (N_2602,N_2410,N_2407);
nand U2603 (N_2603,N_2571,N_2413);
and U2604 (N_2604,N_2476,N_2471);
nor U2605 (N_2605,N_2565,N_2408);
nand U2606 (N_2606,N_2593,N_2531);
or U2607 (N_2607,N_2480,N_2467);
and U2608 (N_2608,N_2550,N_2472);
and U2609 (N_2609,N_2463,N_2449);
nand U2610 (N_2610,N_2504,N_2428);
and U2611 (N_2611,N_2533,N_2591);
and U2612 (N_2612,N_2438,N_2460);
and U2613 (N_2613,N_2590,N_2443);
nor U2614 (N_2614,N_2420,N_2566);
xnor U2615 (N_2615,N_2522,N_2430);
nand U2616 (N_2616,N_2418,N_2493);
nand U2617 (N_2617,N_2481,N_2422);
nor U2618 (N_2618,N_2521,N_2411);
or U2619 (N_2619,N_2499,N_2575);
and U2620 (N_2620,N_2542,N_2577);
nand U2621 (N_2621,N_2517,N_2595);
xor U2622 (N_2622,N_2579,N_2425);
nor U2623 (N_2623,N_2576,N_2477);
or U2624 (N_2624,N_2584,N_2540);
nor U2625 (N_2625,N_2541,N_2532);
nand U2626 (N_2626,N_2543,N_2506);
or U2627 (N_2627,N_2554,N_2570);
nor U2628 (N_2628,N_2492,N_2552);
nand U2629 (N_2629,N_2442,N_2465);
or U2630 (N_2630,N_2503,N_2538);
nor U2631 (N_2631,N_2509,N_2487);
nor U2632 (N_2632,N_2578,N_2406);
nand U2633 (N_2633,N_2569,N_2527);
nand U2634 (N_2634,N_2416,N_2434);
nor U2635 (N_2635,N_2551,N_2536);
nor U2636 (N_2636,N_2489,N_2466);
and U2637 (N_2637,N_2417,N_2520);
nand U2638 (N_2638,N_2451,N_2474);
xor U2639 (N_2639,N_2421,N_2558);
xnor U2640 (N_2640,N_2501,N_2412);
nand U2641 (N_2641,N_2462,N_2468);
and U2642 (N_2642,N_2524,N_2515);
xnor U2643 (N_2643,N_2518,N_2404);
and U2644 (N_2644,N_2588,N_2469);
or U2645 (N_2645,N_2401,N_2557);
xor U2646 (N_2646,N_2447,N_2431);
or U2647 (N_2647,N_2419,N_2486);
nor U2648 (N_2648,N_2546,N_2458);
or U2649 (N_2649,N_2562,N_2429);
or U2650 (N_2650,N_2537,N_2400);
nor U2651 (N_2651,N_2519,N_2567);
nor U2652 (N_2652,N_2507,N_2568);
and U2653 (N_2653,N_2402,N_2491);
or U2654 (N_2654,N_2414,N_2525);
nor U2655 (N_2655,N_2454,N_2482);
and U2656 (N_2656,N_2435,N_2455);
xnor U2657 (N_2657,N_2585,N_2502);
nor U2658 (N_2658,N_2510,N_2439);
xor U2659 (N_2659,N_2459,N_2583);
xnor U2660 (N_2660,N_2497,N_2512);
nand U2661 (N_2661,N_2403,N_2508);
or U2662 (N_2662,N_2405,N_2496);
nand U2663 (N_2663,N_2461,N_2559);
xor U2664 (N_2664,N_2573,N_2445);
and U2665 (N_2665,N_2582,N_2423);
nor U2666 (N_2666,N_2514,N_2516);
nor U2667 (N_2667,N_2424,N_2528);
nand U2668 (N_2668,N_2563,N_2484);
nand U2669 (N_2669,N_2490,N_2534);
nor U2670 (N_2670,N_2580,N_2535);
or U2671 (N_2671,N_2594,N_2452);
xor U2672 (N_2672,N_2589,N_2457);
nand U2673 (N_2673,N_2415,N_2427);
and U2674 (N_2674,N_2598,N_2498);
and U2675 (N_2675,N_2495,N_2556);
nor U2676 (N_2676,N_2488,N_2440);
nor U2677 (N_2677,N_2596,N_2529);
or U2678 (N_2678,N_2555,N_2436);
nand U2679 (N_2679,N_2511,N_2560);
nor U2680 (N_2680,N_2494,N_2478);
nand U2681 (N_2681,N_2544,N_2473);
nor U2682 (N_2682,N_2530,N_2581);
nand U2683 (N_2683,N_2453,N_2505);
and U2684 (N_2684,N_2599,N_2597);
nand U2685 (N_2685,N_2539,N_2433);
nor U2686 (N_2686,N_2564,N_2464);
or U2687 (N_2687,N_2545,N_2448);
xnor U2688 (N_2688,N_2483,N_2513);
nor U2689 (N_2689,N_2446,N_2479);
and U2690 (N_2690,N_2444,N_2426);
xnor U2691 (N_2691,N_2574,N_2523);
nor U2692 (N_2692,N_2500,N_2547);
or U2693 (N_2693,N_2587,N_2456);
and U2694 (N_2694,N_2561,N_2409);
or U2695 (N_2695,N_2470,N_2485);
nor U2696 (N_2696,N_2548,N_2432);
and U2697 (N_2697,N_2549,N_2572);
xnor U2698 (N_2698,N_2437,N_2475);
xor U2699 (N_2699,N_2592,N_2553);
nand U2700 (N_2700,N_2589,N_2502);
nand U2701 (N_2701,N_2416,N_2554);
nor U2702 (N_2702,N_2499,N_2436);
nor U2703 (N_2703,N_2418,N_2425);
nor U2704 (N_2704,N_2514,N_2459);
xor U2705 (N_2705,N_2581,N_2542);
nor U2706 (N_2706,N_2553,N_2434);
xor U2707 (N_2707,N_2566,N_2556);
nand U2708 (N_2708,N_2580,N_2579);
or U2709 (N_2709,N_2404,N_2562);
nand U2710 (N_2710,N_2561,N_2593);
and U2711 (N_2711,N_2575,N_2537);
and U2712 (N_2712,N_2445,N_2589);
xor U2713 (N_2713,N_2436,N_2459);
xnor U2714 (N_2714,N_2517,N_2529);
nand U2715 (N_2715,N_2517,N_2475);
or U2716 (N_2716,N_2556,N_2501);
and U2717 (N_2717,N_2401,N_2445);
nor U2718 (N_2718,N_2545,N_2459);
nor U2719 (N_2719,N_2460,N_2546);
xor U2720 (N_2720,N_2577,N_2426);
and U2721 (N_2721,N_2492,N_2583);
nor U2722 (N_2722,N_2550,N_2539);
nand U2723 (N_2723,N_2423,N_2405);
nand U2724 (N_2724,N_2427,N_2445);
or U2725 (N_2725,N_2555,N_2569);
xor U2726 (N_2726,N_2597,N_2542);
and U2727 (N_2727,N_2562,N_2439);
or U2728 (N_2728,N_2543,N_2480);
or U2729 (N_2729,N_2450,N_2414);
or U2730 (N_2730,N_2488,N_2469);
nand U2731 (N_2731,N_2558,N_2479);
xnor U2732 (N_2732,N_2452,N_2575);
nand U2733 (N_2733,N_2540,N_2549);
nand U2734 (N_2734,N_2546,N_2481);
nor U2735 (N_2735,N_2482,N_2484);
and U2736 (N_2736,N_2470,N_2436);
or U2737 (N_2737,N_2422,N_2583);
or U2738 (N_2738,N_2585,N_2562);
nand U2739 (N_2739,N_2560,N_2531);
nand U2740 (N_2740,N_2443,N_2447);
xor U2741 (N_2741,N_2499,N_2412);
nor U2742 (N_2742,N_2424,N_2537);
and U2743 (N_2743,N_2552,N_2599);
or U2744 (N_2744,N_2482,N_2555);
or U2745 (N_2745,N_2537,N_2445);
or U2746 (N_2746,N_2423,N_2471);
nor U2747 (N_2747,N_2598,N_2499);
nand U2748 (N_2748,N_2544,N_2422);
nor U2749 (N_2749,N_2466,N_2499);
nand U2750 (N_2750,N_2510,N_2550);
nand U2751 (N_2751,N_2498,N_2559);
or U2752 (N_2752,N_2464,N_2550);
and U2753 (N_2753,N_2431,N_2427);
or U2754 (N_2754,N_2462,N_2482);
and U2755 (N_2755,N_2505,N_2403);
nor U2756 (N_2756,N_2536,N_2505);
nor U2757 (N_2757,N_2461,N_2574);
xnor U2758 (N_2758,N_2431,N_2475);
nand U2759 (N_2759,N_2561,N_2570);
xor U2760 (N_2760,N_2500,N_2467);
or U2761 (N_2761,N_2488,N_2580);
or U2762 (N_2762,N_2529,N_2442);
or U2763 (N_2763,N_2561,N_2566);
nand U2764 (N_2764,N_2511,N_2507);
nand U2765 (N_2765,N_2415,N_2403);
nand U2766 (N_2766,N_2461,N_2512);
nor U2767 (N_2767,N_2502,N_2449);
or U2768 (N_2768,N_2479,N_2530);
and U2769 (N_2769,N_2566,N_2507);
and U2770 (N_2770,N_2423,N_2502);
and U2771 (N_2771,N_2486,N_2412);
or U2772 (N_2772,N_2499,N_2442);
nor U2773 (N_2773,N_2570,N_2403);
nor U2774 (N_2774,N_2421,N_2531);
xnor U2775 (N_2775,N_2470,N_2466);
and U2776 (N_2776,N_2577,N_2502);
and U2777 (N_2777,N_2528,N_2442);
or U2778 (N_2778,N_2479,N_2501);
xnor U2779 (N_2779,N_2562,N_2589);
xor U2780 (N_2780,N_2496,N_2559);
and U2781 (N_2781,N_2557,N_2412);
or U2782 (N_2782,N_2491,N_2578);
nor U2783 (N_2783,N_2489,N_2452);
nand U2784 (N_2784,N_2425,N_2513);
or U2785 (N_2785,N_2442,N_2481);
nand U2786 (N_2786,N_2543,N_2422);
or U2787 (N_2787,N_2475,N_2496);
or U2788 (N_2788,N_2552,N_2495);
nor U2789 (N_2789,N_2413,N_2534);
nor U2790 (N_2790,N_2454,N_2432);
or U2791 (N_2791,N_2421,N_2550);
and U2792 (N_2792,N_2594,N_2518);
and U2793 (N_2793,N_2474,N_2454);
nor U2794 (N_2794,N_2403,N_2592);
nor U2795 (N_2795,N_2559,N_2480);
or U2796 (N_2796,N_2510,N_2487);
and U2797 (N_2797,N_2441,N_2401);
xnor U2798 (N_2798,N_2457,N_2587);
nand U2799 (N_2799,N_2447,N_2561);
and U2800 (N_2800,N_2728,N_2751);
nor U2801 (N_2801,N_2607,N_2688);
nor U2802 (N_2802,N_2712,N_2740);
xnor U2803 (N_2803,N_2649,N_2746);
or U2804 (N_2804,N_2759,N_2653);
or U2805 (N_2805,N_2778,N_2753);
or U2806 (N_2806,N_2665,N_2672);
and U2807 (N_2807,N_2723,N_2643);
and U2808 (N_2808,N_2652,N_2601);
xnor U2809 (N_2809,N_2678,N_2609);
and U2810 (N_2810,N_2790,N_2730);
xnor U2811 (N_2811,N_2700,N_2625);
nand U2812 (N_2812,N_2704,N_2705);
or U2813 (N_2813,N_2784,N_2788);
nor U2814 (N_2814,N_2693,N_2673);
and U2815 (N_2815,N_2731,N_2634);
nor U2816 (N_2816,N_2747,N_2638);
or U2817 (N_2817,N_2741,N_2613);
and U2818 (N_2818,N_2755,N_2717);
or U2819 (N_2819,N_2776,N_2659);
nand U2820 (N_2820,N_2795,N_2631);
nand U2821 (N_2821,N_2630,N_2658);
and U2822 (N_2822,N_2670,N_2641);
and U2823 (N_2823,N_2635,N_2618);
and U2824 (N_2824,N_2722,N_2789);
nor U2825 (N_2825,N_2629,N_2781);
or U2826 (N_2826,N_2779,N_2765);
or U2827 (N_2827,N_2655,N_2767);
xor U2828 (N_2828,N_2661,N_2745);
or U2829 (N_2829,N_2614,N_2742);
and U2830 (N_2830,N_2640,N_2674);
and U2831 (N_2831,N_2683,N_2726);
nand U2832 (N_2832,N_2725,N_2716);
xor U2833 (N_2833,N_2689,N_2623);
or U2834 (N_2834,N_2737,N_2762);
and U2835 (N_2835,N_2799,N_2603);
nand U2836 (N_2836,N_2713,N_2718);
nand U2837 (N_2837,N_2729,N_2766);
and U2838 (N_2838,N_2710,N_2696);
and U2839 (N_2839,N_2720,N_2791);
xor U2840 (N_2840,N_2651,N_2738);
xor U2841 (N_2841,N_2701,N_2616);
and U2842 (N_2842,N_2605,N_2758);
and U2843 (N_2843,N_2699,N_2604);
xor U2844 (N_2844,N_2782,N_2780);
or U2845 (N_2845,N_2744,N_2787);
nor U2846 (N_2846,N_2692,N_2632);
xnor U2847 (N_2847,N_2733,N_2736);
or U2848 (N_2848,N_2675,N_2702);
or U2849 (N_2849,N_2752,N_2754);
nor U2850 (N_2850,N_2627,N_2687);
nor U2851 (N_2851,N_2783,N_2724);
and U2852 (N_2852,N_2662,N_2721);
and U2853 (N_2853,N_2719,N_2706);
xnor U2854 (N_2854,N_2608,N_2756);
and U2855 (N_2855,N_2685,N_2624);
and U2856 (N_2856,N_2777,N_2743);
nand U2857 (N_2857,N_2642,N_2771);
and U2858 (N_2858,N_2798,N_2694);
xnor U2859 (N_2859,N_2769,N_2647);
xnor U2860 (N_2860,N_2732,N_2727);
nand U2861 (N_2861,N_2711,N_2748);
or U2862 (N_2862,N_2606,N_2708);
nor U2863 (N_2863,N_2600,N_2628);
nor U2864 (N_2864,N_2602,N_2691);
nand U2865 (N_2865,N_2644,N_2610);
xnor U2866 (N_2866,N_2785,N_2792);
nand U2867 (N_2867,N_2757,N_2794);
nor U2868 (N_2868,N_2682,N_2650);
nor U2869 (N_2869,N_2750,N_2622);
xor U2870 (N_2870,N_2663,N_2735);
nor U2871 (N_2871,N_2612,N_2656);
and U2872 (N_2872,N_2646,N_2773);
or U2873 (N_2873,N_2768,N_2637);
xnor U2874 (N_2874,N_2664,N_2793);
nand U2875 (N_2875,N_2657,N_2667);
nor U2876 (N_2876,N_2715,N_2764);
xor U2877 (N_2877,N_2648,N_2734);
or U2878 (N_2878,N_2760,N_2772);
nand U2879 (N_2879,N_2686,N_2669);
nand U2880 (N_2880,N_2645,N_2684);
or U2881 (N_2881,N_2676,N_2763);
nand U2882 (N_2882,N_2619,N_2739);
and U2883 (N_2883,N_2621,N_2654);
nand U2884 (N_2884,N_2714,N_2668);
or U2885 (N_2885,N_2617,N_2797);
nor U2886 (N_2886,N_2770,N_2680);
xor U2887 (N_2887,N_2709,N_2660);
nand U2888 (N_2888,N_2698,N_2620);
nand U2889 (N_2889,N_2615,N_2749);
nor U2890 (N_2890,N_2633,N_2707);
xnor U2891 (N_2891,N_2681,N_2679);
or U2892 (N_2892,N_2666,N_2703);
nand U2893 (N_2893,N_2639,N_2796);
xor U2894 (N_2894,N_2677,N_2695);
nand U2895 (N_2895,N_2786,N_2636);
nor U2896 (N_2896,N_2690,N_2761);
xnor U2897 (N_2897,N_2697,N_2611);
nand U2898 (N_2898,N_2775,N_2626);
nor U2899 (N_2899,N_2774,N_2671);
and U2900 (N_2900,N_2680,N_2747);
xnor U2901 (N_2901,N_2674,N_2746);
and U2902 (N_2902,N_2626,N_2767);
or U2903 (N_2903,N_2639,N_2666);
nand U2904 (N_2904,N_2741,N_2698);
nor U2905 (N_2905,N_2670,N_2665);
and U2906 (N_2906,N_2776,N_2711);
nor U2907 (N_2907,N_2776,N_2767);
nand U2908 (N_2908,N_2752,N_2652);
and U2909 (N_2909,N_2755,N_2665);
nor U2910 (N_2910,N_2798,N_2697);
and U2911 (N_2911,N_2659,N_2678);
xor U2912 (N_2912,N_2689,N_2760);
or U2913 (N_2913,N_2639,N_2624);
nand U2914 (N_2914,N_2657,N_2777);
nand U2915 (N_2915,N_2654,N_2759);
nand U2916 (N_2916,N_2767,N_2609);
xor U2917 (N_2917,N_2697,N_2793);
nor U2918 (N_2918,N_2649,N_2774);
xnor U2919 (N_2919,N_2605,N_2666);
xor U2920 (N_2920,N_2789,N_2752);
xnor U2921 (N_2921,N_2615,N_2660);
or U2922 (N_2922,N_2743,N_2759);
or U2923 (N_2923,N_2794,N_2609);
and U2924 (N_2924,N_2738,N_2751);
or U2925 (N_2925,N_2708,N_2635);
and U2926 (N_2926,N_2781,N_2690);
and U2927 (N_2927,N_2657,N_2637);
or U2928 (N_2928,N_2699,N_2769);
nor U2929 (N_2929,N_2611,N_2626);
and U2930 (N_2930,N_2715,N_2721);
xor U2931 (N_2931,N_2661,N_2712);
xnor U2932 (N_2932,N_2668,N_2755);
and U2933 (N_2933,N_2795,N_2608);
or U2934 (N_2934,N_2795,N_2643);
nor U2935 (N_2935,N_2647,N_2626);
and U2936 (N_2936,N_2799,N_2779);
and U2937 (N_2937,N_2731,N_2695);
or U2938 (N_2938,N_2789,N_2714);
and U2939 (N_2939,N_2649,N_2628);
nand U2940 (N_2940,N_2696,N_2628);
nand U2941 (N_2941,N_2797,N_2682);
xor U2942 (N_2942,N_2735,N_2798);
nor U2943 (N_2943,N_2796,N_2794);
xor U2944 (N_2944,N_2626,N_2792);
nand U2945 (N_2945,N_2782,N_2633);
nor U2946 (N_2946,N_2739,N_2609);
or U2947 (N_2947,N_2766,N_2777);
and U2948 (N_2948,N_2602,N_2739);
nand U2949 (N_2949,N_2742,N_2778);
nor U2950 (N_2950,N_2727,N_2625);
nand U2951 (N_2951,N_2625,N_2663);
and U2952 (N_2952,N_2668,N_2687);
nor U2953 (N_2953,N_2704,N_2671);
or U2954 (N_2954,N_2798,N_2717);
or U2955 (N_2955,N_2755,N_2799);
and U2956 (N_2956,N_2667,N_2628);
or U2957 (N_2957,N_2672,N_2661);
nor U2958 (N_2958,N_2661,N_2632);
nand U2959 (N_2959,N_2645,N_2660);
xor U2960 (N_2960,N_2679,N_2689);
or U2961 (N_2961,N_2705,N_2734);
nand U2962 (N_2962,N_2691,N_2770);
nor U2963 (N_2963,N_2707,N_2664);
xor U2964 (N_2964,N_2781,N_2763);
nand U2965 (N_2965,N_2724,N_2721);
nand U2966 (N_2966,N_2682,N_2645);
nand U2967 (N_2967,N_2649,N_2790);
and U2968 (N_2968,N_2754,N_2786);
or U2969 (N_2969,N_2752,N_2662);
and U2970 (N_2970,N_2654,N_2600);
and U2971 (N_2971,N_2623,N_2676);
nor U2972 (N_2972,N_2677,N_2619);
or U2973 (N_2973,N_2710,N_2724);
nor U2974 (N_2974,N_2755,N_2683);
and U2975 (N_2975,N_2759,N_2685);
and U2976 (N_2976,N_2727,N_2647);
nand U2977 (N_2977,N_2730,N_2674);
xor U2978 (N_2978,N_2703,N_2724);
xnor U2979 (N_2979,N_2608,N_2727);
xor U2980 (N_2980,N_2664,N_2700);
xnor U2981 (N_2981,N_2767,N_2644);
nand U2982 (N_2982,N_2792,N_2764);
xnor U2983 (N_2983,N_2655,N_2707);
xnor U2984 (N_2984,N_2670,N_2624);
nand U2985 (N_2985,N_2639,N_2694);
nor U2986 (N_2986,N_2753,N_2666);
nor U2987 (N_2987,N_2749,N_2758);
nor U2988 (N_2988,N_2730,N_2646);
xor U2989 (N_2989,N_2765,N_2681);
or U2990 (N_2990,N_2680,N_2713);
xor U2991 (N_2991,N_2700,N_2791);
or U2992 (N_2992,N_2649,N_2600);
nor U2993 (N_2993,N_2798,N_2789);
or U2994 (N_2994,N_2632,N_2721);
or U2995 (N_2995,N_2722,N_2642);
nor U2996 (N_2996,N_2660,N_2628);
or U2997 (N_2997,N_2799,N_2673);
and U2998 (N_2998,N_2602,N_2628);
xnor U2999 (N_2999,N_2771,N_2625);
and UO_0 (O_0,N_2911,N_2860);
nor UO_1 (O_1,N_2849,N_2857);
and UO_2 (O_2,N_2929,N_2876);
or UO_3 (O_3,N_2897,N_2984);
and UO_4 (O_4,N_2954,N_2807);
and UO_5 (O_5,N_2996,N_2943);
xnor UO_6 (O_6,N_2856,N_2917);
nand UO_7 (O_7,N_2949,N_2871);
or UO_8 (O_8,N_2942,N_2999);
xor UO_9 (O_9,N_2889,N_2906);
nand UO_10 (O_10,N_2858,N_2835);
or UO_11 (O_11,N_2991,N_2958);
xnor UO_12 (O_12,N_2814,N_2827);
or UO_13 (O_13,N_2888,N_2966);
nor UO_14 (O_14,N_2840,N_2825);
or UO_15 (O_15,N_2819,N_2956);
xor UO_16 (O_16,N_2811,N_2986);
nor UO_17 (O_17,N_2902,N_2859);
or UO_18 (O_18,N_2981,N_2901);
xnor UO_19 (O_19,N_2924,N_2962);
or UO_20 (O_20,N_2868,N_2852);
nand UO_21 (O_21,N_2878,N_2992);
xnor UO_22 (O_22,N_2913,N_2934);
and UO_23 (O_23,N_2826,N_2872);
and UO_24 (O_24,N_2972,N_2945);
nor UO_25 (O_25,N_2862,N_2842);
or UO_26 (O_26,N_2940,N_2967);
nor UO_27 (O_27,N_2973,N_2908);
and UO_28 (O_28,N_2985,N_2989);
or UO_29 (O_29,N_2895,N_2930);
xnor UO_30 (O_30,N_2905,N_2847);
nor UO_31 (O_31,N_2928,N_2993);
nor UO_32 (O_32,N_2939,N_2968);
nand UO_33 (O_33,N_2927,N_2800);
or UO_34 (O_34,N_2964,N_2932);
or UO_35 (O_35,N_2957,N_2994);
or UO_36 (O_36,N_2823,N_2896);
or UO_37 (O_37,N_2880,N_2831);
nand UO_38 (O_38,N_2832,N_2982);
or UO_39 (O_39,N_2863,N_2970);
and UO_40 (O_40,N_2886,N_2834);
nor UO_41 (O_41,N_2894,N_2841);
xor UO_42 (O_42,N_2893,N_2974);
and UO_43 (O_43,N_2898,N_2976);
nor UO_44 (O_44,N_2815,N_2873);
nor UO_45 (O_45,N_2891,N_2998);
or UO_46 (O_46,N_2830,N_2836);
and UO_47 (O_47,N_2965,N_2806);
nor UO_48 (O_48,N_2801,N_2839);
or UO_49 (O_49,N_2944,N_2803);
nand UO_50 (O_50,N_2955,N_2979);
or UO_51 (O_51,N_2892,N_2805);
xnor UO_52 (O_52,N_2874,N_2990);
xor UO_53 (O_53,N_2978,N_2861);
nand UO_54 (O_54,N_2931,N_2953);
or UO_55 (O_55,N_2920,N_2810);
xor UO_56 (O_56,N_2916,N_2884);
nor UO_57 (O_57,N_2977,N_2837);
and UO_58 (O_58,N_2820,N_2919);
nand UO_59 (O_59,N_2882,N_2809);
and UO_60 (O_60,N_2808,N_2870);
nand UO_61 (O_61,N_2845,N_2997);
nor UO_62 (O_62,N_2960,N_2864);
nand UO_63 (O_63,N_2904,N_2875);
nor UO_64 (O_64,N_2855,N_2804);
xnor UO_65 (O_65,N_2914,N_2813);
nor UO_66 (O_66,N_2833,N_2865);
xor UO_67 (O_67,N_2947,N_2925);
and UO_68 (O_68,N_2903,N_2843);
xnor UO_69 (O_69,N_2822,N_2887);
or UO_70 (O_70,N_2933,N_2952);
or UO_71 (O_71,N_2941,N_2938);
and UO_72 (O_72,N_2853,N_2881);
or UO_73 (O_73,N_2969,N_2817);
and UO_74 (O_74,N_2821,N_2912);
nor UO_75 (O_75,N_2877,N_2936);
or UO_76 (O_76,N_2885,N_2848);
nand UO_77 (O_77,N_2851,N_2818);
nor UO_78 (O_78,N_2866,N_2846);
and UO_79 (O_79,N_2910,N_2951);
xnor UO_80 (O_80,N_2918,N_2995);
nand UO_81 (O_81,N_2937,N_2909);
nor UO_82 (O_82,N_2980,N_2900);
xor UO_83 (O_83,N_2879,N_2850);
nand UO_84 (O_84,N_2921,N_2971);
nor UO_85 (O_85,N_2946,N_2828);
and UO_86 (O_86,N_2948,N_2983);
nor UO_87 (O_87,N_2907,N_2935);
nand UO_88 (O_88,N_2963,N_2829);
or UO_89 (O_89,N_2816,N_2854);
and UO_90 (O_90,N_2922,N_2975);
or UO_91 (O_91,N_2926,N_2959);
or UO_92 (O_92,N_2838,N_2812);
nor UO_93 (O_93,N_2869,N_2867);
nand UO_94 (O_94,N_2890,N_2802);
xor UO_95 (O_95,N_2987,N_2844);
nand UO_96 (O_96,N_2950,N_2915);
and UO_97 (O_97,N_2988,N_2824);
nand UO_98 (O_98,N_2883,N_2961);
or UO_99 (O_99,N_2899,N_2923);
nand UO_100 (O_100,N_2928,N_2927);
and UO_101 (O_101,N_2984,N_2803);
xnor UO_102 (O_102,N_2800,N_2840);
xnor UO_103 (O_103,N_2973,N_2816);
or UO_104 (O_104,N_2833,N_2942);
nor UO_105 (O_105,N_2929,N_2961);
xnor UO_106 (O_106,N_2936,N_2908);
or UO_107 (O_107,N_2954,N_2879);
nor UO_108 (O_108,N_2967,N_2880);
nor UO_109 (O_109,N_2851,N_2891);
nor UO_110 (O_110,N_2959,N_2968);
or UO_111 (O_111,N_2904,N_2983);
nand UO_112 (O_112,N_2816,N_2862);
xnor UO_113 (O_113,N_2951,N_2801);
nor UO_114 (O_114,N_2984,N_2908);
and UO_115 (O_115,N_2923,N_2953);
nand UO_116 (O_116,N_2970,N_2845);
nor UO_117 (O_117,N_2892,N_2835);
or UO_118 (O_118,N_2998,N_2948);
xnor UO_119 (O_119,N_2821,N_2852);
and UO_120 (O_120,N_2954,N_2991);
and UO_121 (O_121,N_2801,N_2939);
and UO_122 (O_122,N_2800,N_2906);
xor UO_123 (O_123,N_2939,N_2830);
and UO_124 (O_124,N_2894,N_2811);
and UO_125 (O_125,N_2968,N_2951);
or UO_126 (O_126,N_2964,N_2976);
xnor UO_127 (O_127,N_2946,N_2915);
xor UO_128 (O_128,N_2819,N_2971);
nor UO_129 (O_129,N_2848,N_2802);
nor UO_130 (O_130,N_2898,N_2916);
and UO_131 (O_131,N_2899,N_2987);
nor UO_132 (O_132,N_2961,N_2878);
or UO_133 (O_133,N_2810,N_2850);
nor UO_134 (O_134,N_2879,N_2928);
xor UO_135 (O_135,N_2953,N_2846);
xnor UO_136 (O_136,N_2981,N_2915);
nand UO_137 (O_137,N_2841,N_2874);
nand UO_138 (O_138,N_2875,N_2934);
xnor UO_139 (O_139,N_2863,N_2955);
xnor UO_140 (O_140,N_2859,N_2952);
or UO_141 (O_141,N_2845,N_2874);
xor UO_142 (O_142,N_2965,N_2879);
nor UO_143 (O_143,N_2850,N_2984);
and UO_144 (O_144,N_2884,N_2810);
and UO_145 (O_145,N_2866,N_2848);
and UO_146 (O_146,N_2977,N_2988);
nand UO_147 (O_147,N_2974,N_2857);
and UO_148 (O_148,N_2977,N_2972);
and UO_149 (O_149,N_2949,N_2842);
nor UO_150 (O_150,N_2842,N_2814);
nor UO_151 (O_151,N_2989,N_2901);
or UO_152 (O_152,N_2936,N_2847);
or UO_153 (O_153,N_2959,N_2840);
xor UO_154 (O_154,N_2990,N_2876);
and UO_155 (O_155,N_2918,N_2872);
or UO_156 (O_156,N_2986,N_2822);
nand UO_157 (O_157,N_2811,N_2935);
xnor UO_158 (O_158,N_2985,N_2893);
nand UO_159 (O_159,N_2933,N_2814);
or UO_160 (O_160,N_2884,N_2941);
nand UO_161 (O_161,N_2928,N_2923);
and UO_162 (O_162,N_2854,N_2801);
xnor UO_163 (O_163,N_2862,N_2894);
nand UO_164 (O_164,N_2819,N_2870);
and UO_165 (O_165,N_2942,N_2996);
nand UO_166 (O_166,N_2910,N_2957);
and UO_167 (O_167,N_2820,N_2908);
nor UO_168 (O_168,N_2935,N_2897);
nand UO_169 (O_169,N_2867,N_2992);
xor UO_170 (O_170,N_2822,N_2977);
xor UO_171 (O_171,N_2906,N_2997);
nor UO_172 (O_172,N_2905,N_2873);
nor UO_173 (O_173,N_2852,N_2810);
or UO_174 (O_174,N_2941,N_2987);
or UO_175 (O_175,N_2940,N_2840);
or UO_176 (O_176,N_2868,N_2853);
nand UO_177 (O_177,N_2830,N_2825);
nor UO_178 (O_178,N_2817,N_2885);
nor UO_179 (O_179,N_2926,N_2867);
or UO_180 (O_180,N_2921,N_2947);
nand UO_181 (O_181,N_2924,N_2875);
nand UO_182 (O_182,N_2883,N_2941);
nor UO_183 (O_183,N_2857,N_2822);
or UO_184 (O_184,N_2820,N_2813);
or UO_185 (O_185,N_2987,N_2947);
or UO_186 (O_186,N_2870,N_2932);
or UO_187 (O_187,N_2905,N_2876);
or UO_188 (O_188,N_2885,N_2937);
or UO_189 (O_189,N_2873,N_2858);
xor UO_190 (O_190,N_2829,N_2807);
nor UO_191 (O_191,N_2969,N_2904);
nand UO_192 (O_192,N_2987,N_2858);
and UO_193 (O_193,N_2926,N_2927);
or UO_194 (O_194,N_2847,N_2978);
or UO_195 (O_195,N_2918,N_2868);
xor UO_196 (O_196,N_2934,N_2971);
nand UO_197 (O_197,N_2875,N_2851);
and UO_198 (O_198,N_2917,N_2882);
nand UO_199 (O_199,N_2855,N_2957);
and UO_200 (O_200,N_2873,N_2865);
nand UO_201 (O_201,N_2844,N_2984);
nor UO_202 (O_202,N_2833,N_2841);
and UO_203 (O_203,N_2835,N_2991);
and UO_204 (O_204,N_2970,N_2838);
and UO_205 (O_205,N_2981,N_2808);
nor UO_206 (O_206,N_2843,N_2983);
nand UO_207 (O_207,N_2880,N_2954);
xnor UO_208 (O_208,N_2930,N_2912);
and UO_209 (O_209,N_2868,N_2876);
or UO_210 (O_210,N_2957,N_2831);
nor UO_211 (O_211,N_2936,N_2963);
and UO_212 (O_212,N_2911,N_2901);
xnor UO_213 (O_213,N_2838,N_2892);
and UO_214 (O_214,N_2997,N_2859);
xnor UO_215 (O_215,N_2957,N_2980);
and UO_216 (O_216,N_2983,N_2839);
and UO_217 (O_217,N_2866,N_2942);
and UO_218 (O_218,N_2999,N_2961);
xnor UO_219 (O_219,N_2841,N_2945);
and UO_220 (O_220,N_2976,N_2841);
xnor UO_221 (O_221,N_2884,N_2886);
and UO_222 (O_222,N_2801,N_2876);
and UO_223 (O_223,N_2959,N_2874);
nand UO_224 (O_224,N_2909,N_2893);
xor UO_225 (O_225,N_2949,N_2933);
nand UO_226 (O_226,N_2829,N_2893);
xnor UO_227 (O_227,N_2891,N_2996);
nor UO_228 (O_228,N_2852,N_2838);
nor UO_229 (O_229,N_2842,N_2968);
or UO_230 (O_230,N_2903,N_2934);
nand UO_231 (O_231,N_2881,N_2942);
and UO_232 (O_232,N_2946,N_2813);
or UO_233 (O_233,N_2998,N_2803);
nor UO_234 (O_234,N_2923,N_2996);
nor UO_235 (O_235,N_2820,N_2969);
or UO_236 (O_236,N_2937,N_2873);
xor UO_237 (O_237,N_2937,N_2900);
or UO_238 (O_238,N_2994,N_2841);
and UO_239 (O_239,N_2955,N_2832);
xnor UO_240 (O_240,N_2877,N_2944);
nor UO_241 (O_241,N_2885,N_2978);
xor UO_242 (O_242,N_2830,N_2828);
or UO_243 (O_243,N_2943,N_2832);
xnor UO_244 (O_244,N_2959,N_2822);
nand UO_245 (O_245,N_2868,N_2980);
nor UO_246 (O_246,N_2939,N_2945);
xnor UO_247 (O_247,N_2830,N_2874);
nor UO_248 (O_248,N_2822,N_2886);
nand UO_249 (O_249,N_2830,N_2838);
nand UO_250 (O_250,N_2836,N_2865);
xor UO_251 (O_251,N_2956,N_2858);
nand UO_252 (O_252,N_2983,N_2961);
nand UO_253 (O_253,N_2851,N_2867);
xnor UO_254 (O_254,N_2872,N_2962);
xnor UO_255 (O_255,N_2920,N_2868);
or UO_256 (O_256,N_2954,N_2834);
nor UO_257 (O_257,N_2832,N_2902);
xnor UO_258 (O_258,N_2879,N_2830);
and UO_259 (O_259,N_2834,N_2910);
nor UO_260 (O_260,N_2897,N_2889);
nand UO_261 (O_261,N_2827,N_2937);
or UO_262 (O_262,N_2911,N_2974);
xnor UO_263 (O_263,N_2938,N_2819);
nor UO_264 (O_264,N_2836,N_2955);
nand UO_265 (O_265,N_2908,N_2863);
or UO_266 (O_266,N_2858,N_2910);
nor UO_267 (O_267,N_2889,N_2916);
nor UO_268 (O_268,N_2811,N_2860);
nor UO_269 (O_269,N_2963,N_2859);
nand UO_270 (O_270,N_2976,N_2892);
and UO_271 (O_271,N_2913,N_2867);
or UO_272 (O_272,N_2890,N_2977);
or UO_273 (O_273,N_2932,N_2898);
nor UO_274 (O_274,N_2849,N_2830);
nor UO_275 (O_275,N_2986,N_2876);
xnor UO_276 (O_276,N_2961,N_2852);
nand UO_277 (O_277,N_2898,N_2823);
nand UO_278 (O_278,N_2940,N_2831);
nor UO_279 (O_279,N_2936,N_2929);
nor UO_280 (O_280,N_2887,N_2850);
or UO_281 (O_281,N_2956,N_2894);
xor UO_282 (O_282,N_2928,N_2976);
nor UO_283 (O_283,N_2995,N_2825);
nand UO_284 (O_284,N_2921,N_2910);
nor UO_285 (O_285,N_2952,N_2997);
or UO_286 (O_286,N_2864,N_2895);
and UO_287 (O_287,N_2946,N_2999);
nor UO_288 (O_288,N_2878,N_2970);
nor UO_289 (O_289,N_2873,N_2984);
nand UO_290 (O_290,N_2853,N_2955);
and UO_291 (O_291,N_2931,N_2908);
or UO_292 (O_292,N_2894,N_2887);
and UO_293 (O_293,N_2960,N_2811);
or UO_294 (O_294,N_2889,N_2813);
or UO_295 (O_295,N_2899,N_2938);
or UO_296 (O_296,N_2969,N_2876);
xnor UO_297 (O_297,N_2940,N_2894);
or UO_298 (O_298,N_2840,N_2949);
nand UO_299 (O_299,N_2941,N_2963);
xnor UO_300 (O_300,N_2936,N_2955);
and UO_301 (O_301,N_2883,N_2895);
xnor UO_302 (O_302,N_2877,N_2979);
and UO_303 (O_303,N_2842,N_2866);
nor UO_304 (O_304,N_2804,N_2941);
nor UO_305 (O_305,N_2974,N_2902);
or UO_306 (O_306,N_2896,N_2950);
nand UO_307 (O_307,N_2939,N_2888);
and UO_308 (O_308,N_2913,N_2829);
or UO_309 (O_309,N_2971,N_2821);
nor UO_310 (O_310,N_2956,N_2946);
nand UO_311 (O_311,N_2896,N_2833);
and UO_312 (O_312,N_2806,N_2884);
nand UO_313 (O_313,N_2980,N_2803);
or UO_314 (O_314,N_2840,N_2968);
nand UO_315 (O_315,N_2847,N_2945);
and UO_316 (O_316,N_2989,N_2956);
nand UO_317 (O_317,N_2814,N_2938);
xor UO_318 (O_318,N_2952,N_2897);
or UO_319 (O_319,N_2933,N_2968);
nand UO_320 (O_320,N_2975,N_2885);
and UO_321 (O_321,N_2824,N_2820);
nand UO_322 (O_322,N_2885,N_2831);
nor UO_323 (O_323,N_2977,N_2860);
nor UO_324 (O_324,N_2852,N_2971);
or UO_325 (O_325,N_2859,N_2933);
nor UO_326 (O_326,N_2896,N_2953);
xor UO_327 (O_327,N_2850,N_2838);
nor UO_328 (O_328,N_2987,N_2953);
nor UO_329 (O_329,N_2947,N_2975);
xnor UO_330 (O_330,N_2861,N_2887);
or UO_331 (O_331,N_2941,N_2970);
xnor UO_332 (O_332,N_2853,N_2985);
nand UO_333 (O_333,N_2849,N_2898);
nor UO_334 (O_334,N_2829,N_2954);
xnor UO_335 (O_335,N_2876,N_2982);
and UO_336 (O_336,N_2869,N_2894);
and UO_337 (O_337,N_2908,N_2980);
and UO_338 (O_338,N_2984,N_2829);
nand UO_339 (O_339,N_2808,N_2820);
nor UO_340 (O_340,N_2934,N_2939);
xnor UO_341 (O_341,N_2852,N_2965);
and UO_342 (O_342,N_2854,N_2869);
or UO_343 (O_343,N_2911,N_2800);
nor UO_344 (O_344,N_2847,N_2830);
nor UO_345 (O_345,N_2909,N_2981);
and UO_346 (O_346,N_2911,N_2902);
or UO_347 (O_347,N_2855,N_2987);
or UO_348 (O_348,N_2941,N_2978);
xnor UO_349 (O_349,N_2856,N_2834);
nand UO_350 (O_350,N_2909,N_2873);
and UO_351 (O_351,N_2899,N_2808);
xor UO_352 (O_352,N_2980,N_2825);
nand UO_353 (O_353,N_2880,N_2976);
xnor UO_354 (O_354,N_2801,N_2833);
nand UO_355 (O_355,N_2856,N_2946);
nor UO_356 (O_356,N_2983,N_2973);
and UO_357 (O_357,N_2945,N_2940);
nor UO_358 (O_358,N_2916,N_2883);
or UO_359 (O_359,N_2963,N_2975);
or UO_360 (O_360,N_2867,N_2998);
nor UO_361 (O_361,N_2991,N_2943);
nor UO_362 (O_362,N_2890,N_2909);
or UO_363 (O_363,N_2804,N_2986);
or UO_364 (O_364,N_2934,N_2826);
and UO_365 (O_365,N_2887,N_2952);
or UO_366 (O_366,N_2920,N_2918);
nand UO_367 (O_367,N_2801,N_2950);
xnor UO_368 (O_368,N_2880,N_2855);
nand UO_369 (O_369,N_2981,N_2995);
nor UO_370 (O_370,N_2969,N_2814);
nor UO_371 (O_371,N_2835,N_2872);
or UO_372 (O_372,N_2877,N_2885);
and UO_373 (O_373,N_2974,N_2822);
or UO_374 (O_374,N_2836,N_2832);
nor UO_375 (O_375,N_2976,N_2895);
nand UO_376 (O_376,N_2919,N_2871);
xor UO_377 (O_377,N_2946,N_2953);
or UO_378 (O_378,N_2900,N_2803);
xor UO_379 (O_379,N_2895,N_2820);
nand UO_380 (O_380,N_2984,N_2991);
or UO_381 (O_381,N_2972,N_2924);
and UO_382 (O_382,N_2886,N_2816);
nand UO_383 (O_383,N_2815,N_2943);
or UO_384 (O_384,N_2838,N_2941);
xnor UO_385 (O_385,N_2835,N_2837);
or UO_386 (O_386,N_2974,N_2851);
and UO_387 (O_387,N_2805,N_2989);
and UO_388 (O_388,N_2922,N_2915);
and UO_389 (O_389,N_2802,N_2849);
nand UO_390 (O_390,N_2895,N_2833);
xnor UO_391 (O_391,N_2958,N_2835);
and UO_392 (O_392,N_2870,N_2863);
nor UO_393 (O_393,N_2883,N_2971);
nand UO_394 (O_394,N_2963,N_2913);
or UO_395 (O_395,N_2913,N_2957);
and UO_396 (O_396,N_2881,N_2897);
nor UO_397 (O_397,N_2869,N_2951);
nor UO_398 (O_398,N_2900,N_2901);
xor UO_399 (O_399,N_2940,N_2859);
nor UO_400 (O_400,N_2885,N_2985);
nand UO_401 (O_401,N_2841,N_2904);
xnor UO_402 (O_402,N_2906,N_2818);
or UO_403 (O_403,N_2894,N_2807);
or UO_404 (O_404,N_2992,N_2805);
nor UO_405 (O_405,N_2872,N_2822);
nand UO_406 (O_406,N_2982,N_2823);
and UO_407 (O_407,N_2868,N_2880);
xor UO_408 (O_408,N_2931,N_2973);
or UO_409 (O_409,N_2927,N_2823);
nand UO_410 (O_410,N_2853,N_2959);
nand UO_411 (O_411,N_2926,N_2912);
xnor UO_412 (O_412,N_2845,N_2907);
nor UO_413 (O_413,N_2987,N_2932);
or UO_414 (O_414,N_2958,N_2977);
nand UO_415 (O_415,N_2876,N_2855);
or UO_416 (O_416,N_2801,N_2884);
xnor UO_417 (O_417,N_2843,N_2877);
nand UO_418 (O_418,N_2981,N_2921);
or UO_419 (O_419,N_2999,N_2859);
and UO_420 (O_420,N_2905,N_2913);
or UO_421 (O_421,N_2961,N_2832);
nand UO_422 (O_422,N_2969,N_2869);
nor UO_423 (O_423,N_2966,N_2860);
or UO_424 (O_424,N_2866,N_2957);
and UO_425 (O_425,N_2854,N_2995);
nor UO_426 (O_426,N_2944,N_2902);
and UO_427 (O_427,N_2957,N_2931);
and UO_428 (O_428,N_2988,N_2911);
nand UO_429 (O_429,N_2836,N_2810);
nor UO_430 (O_430,N_2862,N_2922);
or UO_431 (O_431,N_2950,N_2828);
and UO_432 (O_432,N_2831,N_2937);
nand UO_433 (O_433,N_2941,N_2823);
nand UO_434 (O_434,N_2960,N_2927);
and UO_435 (O_435,N_2924,N_2826);
or UO_436 (O_436,N_2802,N_2816);
xnor UO_437 (O_437,N_2861,N_2987);
and UO_438 (O_438,N_2803,N_2847);
xnor UO_439 (O_439,N_2906,N_2817);
xnor UO_440 (O_440,N_2825,N_2872);
xor UO_441 (O_441,N_2838,N_2862);
or UO_442 (O_442,N_2846,N_2919);
and UO_443 (O_443,N_2847,N_2906);
nor UO_444 (O_444,N_2968,N_2852);
or UO_445 (O_445,N_2989,N_2836);
or UO_446 (O_446,N_2894,N_2991);
and UO_447 (O_447,N_2962,N_2838);
xnor UO_448 (O_448,N_2897,N_2834);
nor UO_449 (O_449,N_2820,N_2811);
nand UO_450 (O_450,N_2818,N_2915);
nor UO_451 (O_451,N_2890,N_2874);
nand UO_452 (O_452,N_2903,N_2904);
or UO_453 (O_453,N_2820,N_2891);
or UO_454 (O_454,N_2884,N_2985);
nand UO_455 (O_455,N_2912,N_2870);
nand UO_456 (O_456,N_2923,N_2954);
nand UO_457 (O_457,N_2967,N_2902);
or UO_458 (O_458,N_2991,N_2889);
and UO_459 (O_459,N_2991,N_2967);
xnor UO_460 (O_460,N_2922,N_2842);
nor UO_461 (O_461,N_2850,N_2827);
and UO_462 (O_462,N_2975,N_2854);
nand UO_463 (O_463,N_2834,N_2862);
nand UO_464 (O_464,N_2952,N_2802);
nor UO_465 (O_465,N_2919,N_2852);
xnor UO_466 (O_466,N_2856,N_2923);
or UO_467 (O_467,N_2844,N_2921);
xor UO_468 (O_468,N_2877,N_2951);
nor UO_469 (O_469,N_2933,N_2897);
or UO_470 (O_470,N_2827,N_2946);
xnor UO_471 (O_471,N_2833,N_2846);
nand UO_472 (O_472,N_2925,N_2884);
nor UO_473 (O_473,N_2933,N_2954);
nand UO_474 (O_474,N_2861,N_2838);
or UO_475 (O_475,N_2976,N_2941);
or UO_476 (O_476,N_2802,N_2870);
xor UO_477 (O_477,N_2976,N_2956);
xnor UO_478 (O_478,N_2946,N_2988);
xor UO_479 (O_479,N_2902,N_2874);
xor UO_480 (O_480,N_2880,N_2828);
or UO_481 (O_481,N_2996,N_2881);
nand UO_482 (O_482,N_2876,N_2979);
or UO_483 (O_483,N_2826,N_2947);
xnor UO_484 (O_484,N_2930,N_2848);
nand UO_485 (O_485,N_2869,N_2920);
nand UO_486 (O_486,N_2873,N_2976);
nand UO_487 (O_487,N_2825,N_2865);
xor UO_488 (O_488,N_2807,N_2840);
and UO_489 (O_489,N_2900,N_2805);
nand UO_490 (O_490,N_2897,N_2928);
nand UO_491 (O_491,N_2954,N_2918);
nor UO_492 (O_492,N_2983,N_2981);
xnor UO_493 (O_493,N_2817,N_2943);
nor UO_494 (O_494,N_2844,N_2967);
or UO_495 (O_495,N_2817,N_2919);
nor UO_496 (O_496,N_2990,N_2922);
and UO_497 (O_497,N_2974,N_2845);
and UO_498 (O_498,N_2989,N_2907);
nor UO_499 (O_499,N_2978,N_2838);
endmodule