module basic_2000_20000_2500_80_levels_10xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
xnor U0 (N_0,In_1414,In_422);
nand U1 (N_1,In_1354,In_1517);
or U2 (N_2,In_547,In_1009);
nor U3 (N_3,In_803,In_1756);
or U4 (N_4,In_1987,In_1960);
and U5 (N_5,In_1672,In_1531);
xnor U6 (N_6,In_1236,In_1565);
nor U7 (N_7,In_523,In_1187);
nor U8 (N_8,In_1640,In_702);
nor U9 (N_9,In_790,In_1720);
nand U10 (N_10,In_892,In_622);
or U11 (N_11,In_283,In_797);
nor U12 (N_12,In_1398,In_594);
and U13 (N_13,In_1358,In_1875);
nand U14 (N_14,In_579,In_1740);
nor U15 (N_15,In_15,In_878);
nor U16 (N_16,In_1990,In_459);
nand U17 (N_17,In_1240,In_409);
and U18 (N_18,In_1221,In_1911);
nor U19 (N_19,In_812,In_323);
nand U20 (N_20,In_1915,In_1820);
nand U21 (N_21,In_777,In_209);
or U22 (N_22,In_43,In_50);
xor U23 (N_23,In_1069,In_1397);
xnor U24 (N_24,In_736,In_641);
nand U25 (N_25,In_1577,In_559);
and U26 (N_26,In_183,In_981);
nor U27 (N_27,In_750,In_1762);
nor U28 (N_28,In_1454,In_679);
or U29 (N_29,In_1077,In_1423);
xnor U30 (N_30,In_286,In_584);
nor U31 (N_31,In_476,In_1555);
or U32 (N_32,In_1040,In_566);
and U33 (N_33,In_1348,In_1973);
xnor U34 (N_34,In_1248,In_185);
xor U35 (N_35,In_1859,In_935);
xnor U36 (N_36,In_152,In_222);
or U37 (N_37,In_488,In_1681);
xor U38 (N_38,In_340,In_1266);
xor U39 (N_39,In_1332,In_1614);
or U40 (N_40,In_1778,In_256);
xor U41 (N_41,In_1342,In_901);
and U42 (N_42,In_247,In_1557);
or U43 (N_43,In_1020,In_592);
and U44 (N_44,In_395,In_1387);
and U45 (N_45,In_1508,In_163);
xor U46 (N_46,In_1054,In_174);
xor U47 (N_47,In_426,In_1933);
xor U48 (N_48,In_1195,In_213);
and U49 (N_49,In_1246,In_258);
nor U50 (N_50,In_714,In_1802);
nand U51 (N_51,In_1873,In_1714);
and U52 (N_52,In_985,In_478);
or U53 (N_53,In_79,In_1623);
nor U54 (N_54,In_568,In_1274);
xor U55 (N_55,In_70,In_681);
or U56 (N_56,In_1015,In_632);
or U57 (N_57,In_1719,In_348);
nand U58 (N_58,In_779,In_1463);
or U59 (N_59,In_1854,In_1496);
and U60 (N_60,In_192,In_1901);
or U61 (N_61,In_914,In_1510);
nand U62 (N_62,In_958,In_98);
and U63 (N_63,In_862,In_1660);
xor U64 (N_64,In_1340,In_569);
or U65 (N_65,In_1251,In_1745);
nor U66 (N_66,In_1665,In_438);
nand U67 (N_67,In_1763,In_386);
xnor U68 (N_68,In_166,In_1170);
nor U69 (N_69,In_1619,In_613);
xor U70 (N_70,In_1698,In_895);
or U71 (N_71,In_443,In_1498);
xor U72 (N_72,In_706,In_1796);
xnor U73 (N_73,In_969,In_907);
nand U74 (N_74,In_1606,In_1403);
nor U75 (N_75,In_781,In_1633);
or U76 (N_76,In_87,In_1917);
nand U77 (N_77,In_102,In_886);
xnor U78 (N_78,In_634,In_837);
or U79 (N_79,In_1569,In_505);
nor U80 (N_80,In_1620,In_123);
nor U81 (N_81,In_1514,In_1062);
nor U82 (N_82,In_13,In_446);
xor U83 (N_83,In_1992,In_1029);
or U84 (N_84,In_1417,In_156);
nand U85 (N_85,In_321,In_408);
or U86 (N_86,In_119,In_1902);
nor U87 (N_87,In_1835,In_650);
nand U88 (N_88,In_358,In_1058);
xnor U89 (N_89,In_415,In_503);
xor U90 (N_90,In_684,In_1632);
or U91 (N_91,In_333,In_1439);
xnor U92 (N_92,In_74,In_1458);
xor U93 (N_93,In_1112,In_961);
or U94 (N_94,In_214,In_1663);
xnor U95 (N_95,In_1554,In_1412);
nand U96 (N_96,In_767,In_117);
and U97 (N_97,In_1519,In_1002);
nand U98 (N_98,In_390,In_1539);
nand U99 (N_99,In_1027,In_1704);
xor U100 (N_100,In_1643,In_419);
or U101 (N_101,In_1923,In_179);
or U102 (N_102,In_1083,In_1352);
xnor U103 (N_103,In_282,In_1413);
or U104 (N_104,In_1891,In_73);
nor U105 (N_105,In_1906,In_234);
nor U106 (N_106,In_1401,In_545);
or U107 (N_107,In_1185,In_805);
nor U108 (N_108,In_1922,In_1657);
nor U109 (N_109,In_1427,In_1530);
or U110 (N_110,In_463,In_1064);
or U111 (N_111,In_1026,In_1264);
nor U112 (N_112,In_458,In_265);
xor U113 (N_113,In_1611,In_1886);
or U114 (N_114,In_114,In_1877);
or U115 (N_115,In_487,In_668);
xnor U116 (N_116,In_1318,In_881);
and U117 (N_117,In_1985,In_1154);
nor U118 (N_118,In_1725,In_153);
or U119 (N_119,In_1177,In_1929);
or U120 (N_120,In_91,In_1716);
xor U121 (N_121,In_1741,In_1038);
xor U122 (N_122,In_1882,In_683);
nor U123 (N_123,In_585,In_1344);
and U124 (N_124,In_1007,In_1879);
and U125 (N_125,In_406,In_277);
or U126 (N_126,In_497,In_988);
nor U127 (N_127,In_1225,In_32);
nand U128 (N_128,In_495,In_1356);
and U129 (N_129,In_270,In_77);
or U130 (N_130,In_1031,In_1307);
nand U131 (N_131,In_301,In_93);
and U132 (N_132,In_1809,In_111);
and U133 (N_133,In_1874,In_39);
or U134 (N_134,In_1223,In_1012);
nand U135 (N_135,In_19,In_1085);
or U136 (N_136,In_811,In_1483);
and U137 (N_137,In_1986,In_1919);
and U138 (N_138,In_786,In_1507);
nor U139 (N_139,In_1374,In_751);
or U140 (N_140,In_842,In_852);
nand U141 (N_141,In_1848,In_733);
nand U142 (N_142,In_1495,In_1553);
nand U143 (N_143,In_1789,In_1988);
xnor U144 (N_144,In_610,In_1547);
or U145 (N_145,In_1263,In_972);
nor U146 (N_146,In_1163,In_264);
xnor U147 (N_147,In_479,In_551);
nor U148 (N_148,In_299,In_30);
or U149 (N_149,In_378,In_1831);
and U150 (N_150,In_928,In_1093);
nor U151 (N_151,In_692,In_1474);
nand U152 (N_152,In_1435,In_834);
xor U153 (N_153,In_1057,In_249);
and U154 (N_154,In_1880,In_729);
nand U155 (N_155,In_1978,In_962);
nor U156 (N_156,In_1422,In_1499);
or U157 (N_157,In_8,In_691);
or U158 (N_158,In_1044,In_1883);
nor U159 (N_159,In_1792,In_335);
nor U160 (N_160,In_553,In_1104);
nor U161 (N_161,In_1226,In_1477);
nand U162 (N_162,In_728,In_695);
nand U163 (N_163,In_1864,In_1090);
nand U164 (N_164,In_802,In_565);
nor U165 (N_165,In_1490,In_589);
or U166 (N_166,In_124,In_1543);
nor U167 (N_167,In_1301,In_9);
xor U168 (N_168,In_1816,In_1192);
and U169 (N_169,In_1063,In_489);
xor U170 (N_170,In_1370,In_616);
nor U171 (N_171,In_387,In_61);
or U172 (N_172,In_1126,In_86);
nand U173 (N_173,In_965,In_267);
and U174 (N_174,In_607,In_1636);
or U175 (N_175,In_1216,In_753);
or U176 (N_176,In_850,In_1273);
xor U177 (N_177,In_555,In_59);
or U178 (N_178,In_1829,In_1833);
xor U179 (N_179,In_158,In_311);
nor U180 (N_180,In_693,In_1947);
or U181 (N_181,In_389,In_1100);
xor U182 (N_182,In_998,In_974);
nor U183 (N_183,In_85,In_1535);
nand U184 (N_184,In_383,In_194);
and U185 (N_185,In_745,In_1359);
nor U186 (N_186,In_987,In_732);
or U187 (N_187,In_120,In_1466);
or U188 (N_188,In_1382,In_305);
xor U189 (N_189,In_500,In_891);
xor U190 (N_190,In_288,In_747);
and U191 (N_191,In_1642,In_761);
or U192 (N_192,In_1686,In_1080);
or U193 (N_193,In_1647,In_1727);
nor U194 (N_194,In_314,In_808);
or U195 (N_195,In_1532,In_823);
xor U196 (N_196,In_1047,In_170);
or U197 (N_197,In_1210,In_1825);
or U198 (N_198,In_26,In_1871);
and U199 (N_199,In_1881,In_1337);
nand U200 (N_200,In_1312,In_511);
or U201 (N_201,In_1509,In_947);
nand U202 (N_202,In_1379,In_1147);
or U203 (N_203,In_1323,In_1235);
or U204 (N_204,In_1972,In_587);
or U205 (N_205,In_672,In_544);
and U206 (N_206,In_435,In_1368);
nand U207 (N_207,In_354,In_1229);
and U208 (N_208,In_997,In_1284);
xor U209 (N_209,In_1552,In_1257);
nand U210 (N_210,In_1797,In_1117);
or U211 (N_211,In_135,In_289);
or U212 (N_212,In_626,In_454);
nand U213 (N_213,In_101,In_273);
nor U214 (N_214,In_1476,In_976);
xor U215 (N_215,In_1494,In_1575);
xor U216 (N_216,In_770,In_370);
xor U217 (N_217,In_851,In_597);
nor U218 (N_218,In_82,In_1892);
or U219 (N_219,In_345,In_448);
or U220 (N_220,In_184,In_884);
nand U221 (N_221,In_1380,In_44);
and U222 (N_222,In_903,In_1089);
and U223 (N_223,In_88,In_591);
nand U224 (N_224,In_1980,In_1750);
nand U225 (N_225,In_1869,In_2);
or U226 (N_226,In_1910,In_1781);
nor U227 (N_227,In_1303,In_959);
xor U228 (N_228,In_524,In_1376);
nor U229 (N_229,In_540,In_926);
nor U230 (N_230,In_697,In_104);
and U231 (N_231,In_1479,In_995);
nand U232 (N_232,In_1637,In_1732);
and U233 (N_233,In_1677,In_388);
nand U234 (N_234,In_758,In_1429);
or U235 (N_235,In_466,In_921);
nor U236 (N_236,In_840,In_1308);
nand U237 (N_237,In_1393,In_437);
nand U238 (N_238,In_1161,In_1119);
and U239 (N_239,In_1931,In_240);
and U240 (N_240,In_1484,In_670);
or U241 (N_241,In_1203,In_1655);
nor U242 (N_242,In_1897,In_1433);
or U243 (N_243,In_312,In_1473);
nand U244 (N_244,In_609,In_493);
nand U245 (N_245,In_490,In_1916);
and U246 (N_246,In_468,In_867);
and U247 (N_247,In_731,In_1710);
nand U248 (N_248,In_1219,In_975);
xnor U249 (N_249,In_1288,In_701);
or U250 (N_250,In_1924,In_1037);
and U251 (N_251,In_542,In_1363);
xor U252 (N_252,N_127,In_190);
xnor U253 (N_253,In_703,In_1868);
or U254 (N_254,In_1259,In_1679);
nor U255 (N_255,In_515,In_742);
or U256 (N_256,In_1828,In_212);
xnor U257 (N_257,In_897,In_430);
xor U258 (N_258,In_1735,In_285);
xor U259 (N_259,In_920,N_44);
nand U260 (N_260,N_215,In_1932);
nand U261 (N_261,In_1391,In_902);
or U262 (N_262,In_494,In_7);
and U263 (N_263,N_88,In_1261);
or U264 (N_264,In_665,N_161);
or U265 (N_265,In_1728,In_1239);
nor U266 (N_266,In_943,In_1849);
nor U267 (N_267,In_28,N_176);
nor U268 (N_268,In_1280,In_1141);
and U269 (N_269,N_110,In_1963);
nor U270 (N_270,In_1107,In_1646);
xnor U271 (N_271,In_1810,In_164);
or U272 (N_272,In_825,In_1421);
or U273 (N_273,N_195,In_1262);
nand U274 (N_274,In_217,N_124);
and U275 (N_275,In_1858,In_84);
nor U276 (N_276,In_1768,In_865);
xor U277 (N_277,N_217,In_816);
or U278 (N_278,In_1172,In_1779);
and U279 (N_279,N_99,In_230);
or U280 (N_280,N_202,In_664);
xor U281 (N_281,In_1813,N_30);
nand U282 (N_282,In_1298,In_831);
or U283 (N_283,In_906,In_938);
nor U284 (N_284,In_1110,In_633);
xor U285 (N_285,N_228,In_1587);
xor U286 (N_286,In_483,In_121);
or U287 (N_287,In_640,In_1232);
nand U288 (N_288,In_1049,In_450);
nand U289 (N_289,In_1281,In_939);
and U290 (N_290,N_206,In_983);
and U291 (N_291,In_362,In_244);
nand U292 (N_292,In_611,In_1856);
xnor U293 (N_293,In_1625,In_394);
nand U294 (N_294,In_1299,In_1708);
and U295 (N_295,In_1367,In_198);
or U296 (N_296,In_306,In_659);
xnor U297 (N_297,In_338,In_912);
or U298 (N_298,In_1966,In_5);
nor U299 (N_299,In_241,In_696);
nand U300 (N_300,In_1122,In_1682);
xnor U301 (N_301,In_473,In_480);
or U302 (N_302,In_762,N_138);
xor U303 (N_303,In_374,In_1132);
nand U304 (N_304,In_229,In_1205);
nand U305 (N_305,In_1314,In_182);
nor U306 (N_306,In_1139,N_204);
and U307 (N_307,In_573,In_328);
or U308 (N_308,In_1523,In_24);
nand U309 (N_309,In_1343,In_877);
and U310 (N_310,In_1218,In_882);
and U311 (N_311,In_1157,In_1717);
or U312 (N_312,In_1418,In_1295);
or U313 (N_313,In_1445,In_945);
nor U314 (N_314,In_815,In_1325);
nand U315 (N_315,In_67,In_1692);
xnor U316 (N_316,In_1124,In_482);
nor U317 (N_317,In_1631,In_1194);
nand U318 (N_318,In_1250,In_744);
or U319 (N_319,In_1041,In_1755);
xnor U320 (N_320,In_1608,In_1447);
xor U321 (N_321,In_1390,In_1941);
nor U322 (N_322,In_1217,In_800);
and U323 (N_323,In_982,N_74);
nor U324 (N_324,In_845,In_860);
nand U325 (N_325,In_1939,In_1151);
nand U326 (N_326,In_1355,N_224);
or U327 (N_327,N_49,In_1475);
and U328 (N_328,In_1607,In_1389);
and U329 (N_329,In_643,In_916);
nor U330 (N_330,In_1866,In_1442);
or U331 (N_331,In_1938,In_1827);
xor U332 (N_332,In_1105,In_324);
nor U333 (N_333,N_162,In_826);
or U334 (N_334,In_1073,In_1837);
xor U335 (N_335,In_136,In_588);
nor U336 (N_336,In_1346,In_978);
xor U337 (N_337,In_531,In_1803);
or U338 (N_338,In_1169,In_868);
nand U339 (N_339,In_1648,In_449);
xnor U340 (N_340,In_1513,In_1805);
nand U341 (N_341,In_1184,In_1615);
and U342 (N_342,In_1153,In_1998);
nor U343 (N_343,In_373,In_1405);
and U344 (N_344,In_595,In_129);
xor U345 (N_345,In_1302,In_1574);
xor U346 (N_346,In_228,In_1683);
and U347 (N_347,In_1455,In_1739);
nand U348 (N_348,In_829,In_1247);
or U349 (N_349,In_1198,In_1160);
nand U350 (N_350,In_727,In_735);
or U351 (N_351,In_467,In_989);
nand U352 (N_352,N_225,In_708);
xnor U353 (N_353,In_722,N_31);
or U354 (N_354,In_445,In_1505);
xnor U355 (N_355,In_376,In_1759);
nor U356 (N_356,In_1222,In_1788);
or U357 (N_357,In_1364,In_1357);
or U358 (N_358,In_1841,In_1179);
or U359 (N_359,In_1306,In_1487);
xor U360 (N_360,In_960,N_46);
nand U361 (N_361,In_1061,In_1905);
or U362 (N_362,In_105,In_310);
nor U363 (N_363,In_1667,In_873);
or U364 (N_364,In_1300,In_225);
or U365 (N_365,In_1878,In_269);
nor U366 (N_366,In_1521,In_1214);
and U367 (N_367,N_101,In_1627);
nand U368 (N_368,In_71,In_45);
xnor U369 (N_369,In_1116,In_890);
and U370 (N_370,In_952,In_138);
and U371 (N_371,In_1451,N_182);
and U372 (N_372,In_843,N_91);
xor U373 (N_373,In_331,In_1738);
xor U374 (N_374,In_502,In_1075);
nand U375 (N_375,In_874,In_100);
xor U376 (N_376,In_1688,In_1134);
nor U377 (N_377,In_10,In_262);
xor U378 (N_378,In_280,In_1512);
or U379 (N_379,In_99,In_717);
xnor U380 (N_380,In_973,In_25);
or U381 (N_381,In_516,In_535);
or U382 (N_382,In_20,In_504);
or U383 (N_383,N_175,In_397);
nor U384 (N_384,In_833,In_615);
and U385 (N_385,In_1597,In_1485);
or U386 (N_386,In_1207,In_178);
and U387 (N_387,In_506,In_252);
and U388 (N_388,In_1690,In_1436);
xor U389 (N_389,In_391,In_364);
or U390 (N_390,In_294,In_1043);
nand U391 (N_391,In_1842,In_980);
and U392 (N_392,In_1826,In_858);
xnor U393 (N_393,In_635,In_904);
and U394 (N_394,In_1086,N_207);
nor U395 (N_395,In_1067,In_316);
xor U396 (N_396,N_84,In_861);
xor U397 (N_397,In_940,N_235);
nand U398 (N_398,N_134,In_836);
and U399 (N_399,In_206,In_344);
nand U400 (N_400,N_231,In_1324);
nand U401 (N_401,In_1937,N_118);
xor U402 (N_402,In_1249,In_1680);
nor U403 (N_403,In_1457,N_216);
and U404 (N_404,In_1101,In_196);
or U405 (N_405,In_54,In_1201);
xor U406 (N_406,In_404,In_266);
xor U407 (N_407,In_3,In_1601);
or U408 (N_408,N_98,In_1133);
nor U409 (N_409,In_1995,In_65);
nor U410 (N_410,In_1560,In_1556);
or U411 (N_411,In_620,In_1857);
nor U412 (N_412,In_789,In_402);
nand U413 (N_413,In_618,In_1662);
xor U414 (N_414,N_14,In_1900);
nor U415 (N_415,N_117,In_700);
nor U416 (N_416,In_1258,In_924);
or U417 (N_417,In_413,In_1546);
or U418 (N_418,In_1511,In_1034);
nor U419 (N_419,In_602,In_1087);
and U420 (N_420,In_799,In_963);
nor U421 (N_421,N_222,In_1098);
nor U422 (N_422,N_236,In_1965);
or U423 (N_423,In_1056,In_1138);
nor U424 (N_424,In_22,In_1536);
and U425 (N_425,In_1290,N_6);
xnor U426 (N_426,N_50,In_1730);
nor U427 (N_427,In_534,In_1171);
or U428 (N_428,In_704,In_315);
nand U429 (N_429,In_582,In_1622);
xor U430 (N_430,In_1000,In_716);
or U431 (N_431,In_1005,N_87);
or U432 (N_432,In_1899,In_457);
or U433 (N_433,In_908,In_721);
xnor U434 (N_434,In_1036,In_1890);
nor U435 (N_435,In_1943,In_1066);
and U436 (N_436,In_838,N_63);
nand U437 (N_437,N_37,In_1215);
and U438 (N_438,In_243,In_675);
nor U439 (N_439,In_1658,In_110);
nor U440 (N_440,In_853,In_1074);
and U441 (N_441,N_40,N_62);
or U442 (N_442,In_549,In_1957);
nand U443 (N_443,In_1204,In_517);
nand U444 (N_444,In_1626,In_1599);
or U445 (N_445,In_147,In_1956);
nor U446 (N_446,In_1592,In_1654);
nor U447 (N_447,In_1021,N_66);
and U448 (N_448,In_1538,In_1595);
xor U449 (N_449,In_260,In_403);
and U450 (N_450,In_898,N_187);
xor U451 (N_451,In_232,In_599);
nand U452 (N_452,N_22,In_1936);
nor U453 (N_453,N_78,In_1144);
xnor U454 (N_454,In_423,In_1737);
xor U455 (N_455,In_820,In_550);
or U456 (N_456,In_49,N_238);
nand U457 (N_457,N_148,In_245);
xnor U458 (N_458,In_1310,N_122);
nor U459 (N_459,N_90,In_1754);
or U460 (N_460,In_1920,In_864);
and U461 (N_461,In_349,In_1887);
nor U462 (N_462,In_127,In_1651);
nor U463 (N_463,In_581,In_297);
and U464 (N_464,In_1431,In_876);
and U465 (N_465,In_96,In_1961);
and U466 (N_466,In_526,In_623);
and U467 (N_467,In_1092,In_1470);
nor U468 (N_468,In_63,In_1287);
or U469 (N_469,In_1621,In_1561);
xor U470 (N_470,In_1861,In_760);
nand U471 (N_471,In_1497,In_600);
nor U472 (N_472,In_1594,In_1948);
nand U473 (N_473,In_1807,In_1865);
nor U474 (N_474,In_528,In_1600);
and U475 (N_475,N_155,In_1840);
nor U476 (N_476,In_1734,N_226);
xor U477 (N_477,In_627,N_230);
xnor U478 (N_478,N_60,In_1088);
nand U479 (N_479,In_1743,In_525);
or U480 (N_480,In_278,In_146);
nor U481 (N_481,In_1590,In_856);
nand U482 (N_482,In_271,In_220);
and U483 (N_483,In_4,In_1415);
or U484 (N_484,In_967,In_509);
and U485 (N_485,In_946,In_97);
xnor U486 (N_486,N_17,In_334);
and U487 (N_487,In_496,In_519);
nand U488 (N_488,In_1804,N_144);
nand U489 (N_489,In_456,In_1641);
xnor U490 (N_490,N_152,In_1286);
nand U491 (N_491,In_414,N_214);
nand U492 (N_492,N_70,In_1996);
nor U493 (N_493,In_669,In_1366);
and U494 (N_494,In_532,In_329);
and U495 (N_495,In_472,N_237);
nand U496 (N_496,N_4,N_142);
nand U497 (N_497,In_593,In_444);
nor U498 (N_498,In_1130,N_178);
nor U499 (N_499,In_677,N_168);
xor U500 (N_500,In_977,In_1438);
nand U501 (N_501,In_849,In_1814);
or U502 (N_502,In_23,In_1113);
or U503 (N_503,In_1793,In_636);
and U504 (N_504,N_129,N_71);
and U505 (N_505,In_195,In_188);
and U506 (N_506,N_194,In_1109);
nor U507 (N_507,In_1950,N_496);
and U508 (N_508,In_1908,N_151);
nand U509 (N_509,N_199,In_1824);
and U510 (N_510,N_174,In_1541);
nor U511 (N_511,In_1628,N_45);
nor U512 (N_512,N_240,In_560);
nand U513 (N_513,In_1634,N_58);
or U514 (N_514,In_979,N_402);
xor U515 (N_515,In_224,In_1545);
nand U516 (N_516,In_385,N_2);
xor U517 (N_517,N_334,In_1079);
nand U518 (N_518,In_1976,N_273);
and U519 (N_519,In_211,In_994);
xor U520 (N_520,In_501,N_410);
or U521 (N_521,N_220,In_1492);
nand U522 (N_522,In_221,N_434);
nor U523 (N_523,In_1850,In_1572);
nand U524 (N_524,N_52,In_863);
xor U525 (N_525,In_527,In_1516);
xnor U526 (N_526,In_713,N_462);
xor U527 (N_527,In_1146,In_905);
nand U528 (N_528,In_1396,In_711);
and U529 (N_529,In_1952,In_785);
nand U530 (N_530,In_412,N_437);
xnor U531 (N_531,In_1659,In_796);
and U532 (N_532,N_371,In_1294);
xor U533 (N_533,N_280,In_1563);
or U534 (N_534,In_719,In_1664);
nand U535 (N_535,In_1242,In_1700);
or U536 (N_536,In_1014,In_513);
xor U537 (N_537,N_1,In_485);
or U538 (N_538,N_172,In_888);
and U539 (N_539,In_181,N_329);
or U540 (N_540,In_598,In_580);
xnor U541 (N_541,In_1766,N_476);
and U542 (N_542,N_9,N_141);
xnor U543 (N_543,In_1791,N_257);
nand U544 (N_544,N_53,N_86);
or U545 (N_545,N_314,In_1174);
nand U546 (N_546,In_1771,In_1851);
xnor U547 (N_547,N_456,In_1671);
and U548 (N_548,N_188,In_1155);
or U549 (N_549,N_324,N_139);
and U550 (N_550,N_450,N_365);
nand U551 (N_551,N_317,In_429);
and U552 (N_552,In_720,In_1321);
nand U553 (N_553,In_1610,In_934);
nand U554 (N_554,In_499,In_941);
nand U555 (N_555,In_1722,In_1602);
xor U556 (N_556,In_548,In_1156);
nor U557 (N_557,N_103,In_543);
xnor U558 (N_558,N_452,In_191);
nand U559 (N_559,N_160,N_143);
or U560 (N_560,In_319,In_226);
or U561 (N_561,N_95,In_416);
nand U562 (N_562,In_1870,In_377);
and U563 (N_563,N_287,N_331);
and U564 (N_564,In_1050,N_259);
and U565 (N_565,N_113,In_1570);
nand U566 (N_566,In_1638,N_270);
nor U567 (N_567,N_362,N_183);
xor U568 (N_568,In_1336,In_1320);
or U569 (N_569,N_375,In_1581);
xnor U570 (N_570,In_498,N_391);
nor U571 (N_571,In_647,N_128);
nand U572 (N_572,In_1761,In_1526);
and U573 (N_573,In_1383,N_481);
nand U574 (N_574,In_347,In_1685);
and U575 (N_575,N_311,In_398);
nand U576 (N_576,N_305,N_342);
xor U577 (N_577,In_126,In_410);
or U578 (N_578,N_429,N_42);
or U579 (N_579,In_366,In_686);
and U580 (N_580,In_1395,N_405);
nand U581 (N_581,In_1465,In_1048);
xnor U582 (N_582,In_773,In_1317);
nor U583 (N_583,In_1392,In_1428);
nor U584 (N_584,In_578,N_366);
or U585 (N_585,In_1488,In_562);
or U586 (N_586,In_1189,In_791);
nor U587 (N_587,In_1846,N_140);
nor U588 (N_588,N_380,In_1167);
nand U589 (N_589,In_1598,In_1381);
or U590 (N_590,In_653,N_385);
nand U591 (N_591,In_652,In_360);
and U592 (N_592,In_1618,In_1017);
xor U593 (N_593,In_130,In_37);
xor U594 (N_594,In_1588,In_1253);
or U595 (N_595,In_1528,N_260);
nand U596 (N_596,N_154,N_286);
nor U597 (N_597,In_1549,In_356);
and U598 (N_598,In_1065,N_210);
or U599 (N_599,In_352,N_468);
xor U600 (N_600,N_105,In_1894);
nand U601 (N_601,In_1386,N_67);
nor U602 (N_602,In_1042,In_1168);
or U603 (N_603,In_392,N_353);
and U604 (N_604,In_596,In_361);
nand U605 (N_605,In_1613,In_1702);
nand U606 (N_606,N_83,In_320);
nor U607 (N_607,In_326,N_247);
nand U608 (N_608,In_782,In_514);
or U609 (N_609,N_406,In_202);
nand U610 (N_610,N_373,In_957);
nand U611 (N_611,N_408,In_236);
or U612 (N_612,In_993,In_827);
nand U613 (N_613,In_1503,N_100);
xor U614 (N_614,In_1989,N_328);
nor U615 (N_615,N_399,In_461);
and U616 (N_616,In_630,In_518);
nor U617 (N_617,N_368,In_1668);
xnor U618 (N_618,In_342,In_1921);
or U619 (N_619,N_38,In_554);
and U620 (N_620,In_1925,In_730);
and U621 (N_621,N_319,N_163);
or U622 (N_622,N_120,N_340);
nor U623 (N_623,N_422,N_414);
and U624 (N_624,N_295,In_813);
and U625 (N_625,In_210,N_497);
and U626 (N_626,In_418,In_1265);
nor U627 (N_627,In_1913,In_1289);
xor U628 (N_628,In_639,In_740);
xnor U629 (N_629,In_1930,N_472);
nor U630 (N_630,N_409,In_1033);
xnor U631 (N_631,In_1669,In_538);
and U632 (N_632,In_1958,In_673);
and U633 (N_633,In_199,In_255);
xor U634 (N_634,In_1534,In_756);
nor U635 (N_635,N_77,N_292);
nor U636 (N_636,In_1839,In_899);
and U637 (N_637,In_1845,N_417);
and U638 (N_638,In_583,N_474);
or U639 (N_639,In_1350,In_654);
and U640 (N_640,In_764,N_464);
or U641 (N_641,In_1464,In_1018);
and U642 (N_642,In_667,In_674);
or U643 (N_643,In_1322,N_321);
and U644 (N_644,In_1934,In_971);
nand U645 (N_645,In_869,N_299);
and U646 (N_646,In_216,In_1830);
nand U647 (N_647,In_918,In_208);
or U648 (N_648,In_949,N_131);
xor U649 (N_649,In_1649,In_1777);
nor U650 (N_650,In_1522,N_132);
xnor U651 (N_651,In_1409,In_330);
and U652 (N_652,N_285,N_498);
xor U653 (N_653,In_1885,In_365);
xor U654 (N_654,In_109,In_75);
nor U655 (N_655,In_180,In_451);
nand U656 (N_656,In_748,In_1148);
or U657 (N_657,N_256,In_1991);
and U658 (N_658,In_1853,N_69);
nand U659 (N_659,N_418,In_1121);
xnor U660 (N_660,In_1585,In_1568);
or U661 (N_661,N_477,In_177);
and U662 (N_662,In_1404,In_614);
or U663 (N_663,N_420,In_1770);
xnor U664 (N_664,In_642,In_1125);
or U665 (N_665,In_557,In_1233);
or U666 (N_666,In_655,N_73);
nor U667 (N_667,N_169,In_66);
nand U668 (N_668,In_1441,N_423);
xnor U669 (N_669,In_1907,In_1313);
and U670 (N_670,In_1772,In_625);
nor U671 (N_671,In_1975,In_937);
xnor U672 (N_672,In_1806,In_1001);
nand U673 (N_673,In_1784,In_141);
nand U674 (N_674,In_1202,In_427);
or U675 (N_675,N_341,In_1305);
and U676 (N_676,In_896,N_20);
or U677 (N_677,In_1955,N_315);
and U678 (N_678,N_82,In_162);
xnor U679 (N_679,N_359,N_489);
and U680 (N_680,N_193,In_1378);
and U681 (N_681,N_369,In_1515);
xnor U682 (N_682,In_919,In_1715);
or U683 (N_683,In_556,In_680);
or U684 (N_684,N_108,In_1186);
nor U685 (N_685,N_146,In_712);
or U686 (N_686,N_258,In_1673);
nor U687 (N_687,In_1410,In_1399);
or U688 (N_688,N_381,In_1695);
nand U689 (N_689,In_765,N_370);
nor U690 (N_690,In_132,In_1764);
and U691 (N_691,In_671,In_828);
and U692 (N_692,In_1460,In_715);
nor U693 (N_693,N_411,In_1749);
or U694 (N_694,N_123,In_401);
or U695 (N_695,In_870,In_1006);
or U696 (N_696,In_841,In_133);
nor U697 (N_697,In_1701,In_1402);
or U698 (N_698,In_1801,N_471);
and U699 (N_699,In_1142,In_1744);
nor U700 (N_700,In_46,In_31);
nor U701 (N_701,In_1003,In_522);
or U702 (N_702,N_387,In_619);
nor U703 (N_703,In_368,In_970);
xor U704 (N_704,In_1993,N_268);
or U705 (N_705,In_1970,N_153);
nand U706 (N_706,N_59,In_900);
and U707 (N_707,In_629,In_1566);
nand U708 (N_708,In_1462,N_346);
xnor U709 (N_709,In_336,In_48);
and U710 (N_710,In_433,In_925);
or U711 (N_711,In_570,N_458);
or U712 (N_712,In_250,N_436);
xnor U713 (N_713,In_1983,In_948);
nor U714 (N_714,In_1645,In_795);
nor U715 (N_715,In_1211,In_1334);
nor U716 (N_716,N_289,N_262);
nand U717 (N_717,N_241,In_1624);
nand U718 (N_718,In_11,N_484);
or U719 (N_719,In_1670,N_364);
xnor U720 (N_720,In_1035,In_168);
nand U721 (N_721,In_1843,In_1537);
and U722 (N_722,N_13,In_1296);
and U723 (N_723,In_1967,In_474);
nor U724 (N_724,In_238,N_34);
and U725 (N_725,In_203,In_1889);
nor U726 (N_726,In_215,N_177);
xor U727 (N_727,In_1852,In_1571);
nand U728 (N_728,N_449,N_250);
and U729 (N_729,In_1361,In_1267);
nand U730 (N_730,In_1190,In_460);
nor U731 (N_731,N_3,In_1212);
and U732 (N_732,In_1372,In_875);
or U733 (N_733,In_968,N_5);
nand U734 (N_734,In_1576,In_776);
or U735 (N_735,N_293,In_572);
nand U736 (N_736,In_38,In_1019);
and U737 (N_737,In_1558,In_1518);
nand U738 (N_738,In_40,N_248);
and U739 (N_739,In_1544,In_724);
and U740 (N_740,In_259,In_56);
nor U741 (N_741,N_167,In_1137);
and U742 (N_742,N_276,N_213);
xor U743 (N_743,N_93,In_1103);
nor U744 (N_744,N_397,N_56);
or U745 (N_745,In_689,In_1821);
nand U746 (N_746,In_292,In_1731);
nand U747 (N_747,N_428,In_953);
or U748 (N_748,In_855,N_386);
nand U749 (N_749,In_143,N_48);
and U750 (N_750,In_1165,In_439);
or U751 (N_751,In_1675,In_510);
xor U752 (N_752,In_1694,N_243);
and U753 (N_753,N_500,N_739);
and U754 (N_754,N_737,N_485);
and U755 (N_755,In_991,N_519);
nand U756 (N_756,In_1482,In_246);
or U757 (N_757,In_1834,N_310);
and U758 (N_758,N_274,In_1400);
or U759 (N_759,N_503,N_173);
nor U760 (N_760,In_481,In_1815);
xnor U761 (N_761,N_383,N_16);
or U762 (N_762,In_541,N_0);
and U763 (N_763,In_219,N_447);
xnor U764 (N_764,In_1461,In_1456);
or U765 (N_765,In_1081,N_119);
nand U766 (N_766,N_245,N_244);
nor U767 (N_767,In_1697,N_502);
nor U768 (N_768,In_780,In_1812);
nor U769 (N_769,In_1832,N_656);
xnor U770 (N_770,N_80,In_1818);
nand U771 (N_771,In_1548,In_1529);
and U772 (N_772,N_323,In_436);
or U773 (N_773,In_1297,N_657);
nor U774 (N_774,In_685,In_160);
xnor U775 (N_775,In_879,N_730);
xnor U776 (N_776,N_438,N_590);
and U777 (N_777,In_1178,N_170);
nand U778 (N_778,In_379,In_1078);
or U779 (N_779,N_125,N_707);
nor U780 (N_780,In_428,N_427);
nand U781 (N_781,N_627,In_1183);
nor U782 (N_782,In_1245,In_41);
and U783 (N_783,In_817,In_343);
and U784 (N_784,In_644,In_227);
xor U785 (N_785,N_318,N_595);
and U786 (N_786,N_494,N_446);
nor U787 (N_787,In_1844,In_80);
or U788 (N_788,In_1256,In_367);
or U789 (N_789,N_480,N_539);
and U790 (N_790,N_579,In_1729);
and U791 (N_791,N_165,In_318);
nand U792 (N_792,N_563,In_893);
or U793 (N_793,N_185,In_1120);
nand U794 (N_794,In_806,In_1025);
and U795 (N_795,In_1656,In_718);
or U796 (N_796,N_622,In_1798);
or U797 (N_797,In_281,In_399);
and U798 (N_798,In_769,In_17);
nand U799 (N_799,In_1437,N_130);
nand U800 (N_800,In_821,In_1326);
and U801 (N_801,N_582,N_548);
xnor U802 (N_802,N_734,In_656);
and U803 (N_803,N_478,N_526);
nand U804 (N_804,N_719,In_814);
and U805 (N_805,N_640,N_413);
nor U806 (N_806,N_608,N_249);
xor U807 (N_807,N_486,In_440);
nand U808 (N_808,In_628,N_221);
nand U809 (N_809,N_425,In_1311);
xnor U810 (N_810,In_200,In_1927);
and U811 (N_811,In_300,N_407);
or U812 (N_812,In_1252,In_1096);
nor U813 (N_813,In_83,N_543);
or U814 (N_814,N_252,N_617);
and U815 (N_815,N_439,In_1285);
or U816 (N_816,In_743,In_1115);
nor U817 (N_817,In_1384,In_564);
nor U818 (N_818,In_1942,In_1974);
nand U819 (N_819,In_150,In_1159);
nor U820 (N_820,In_52,In_1748);
and U821 (N_821,In_1783,In_1709);
or U822 (N_822,N_253,In_909);
xor U823 (N_823,N_504,N_112);
nor U824 (N_824,In_149,In_1373);
xnor U825 (N_825,N_677,In_880);
nand U826 (N_826,In_115,N_164);
xnor U827 (N_827,N_388,In_1860);
xnor U828 (N_828,N_121,In_142);
nand U829 (N_829,In_295,In_1525);
xor U830 (N_830,In_1220,N_619);
or U831 (N_831,In_1540,N_506);
and U832 (N_832,In_155,In_866);
or U833 (N_833,In_193,N_89);
nor U834 (N_834,N_363,N_688);
nor U835 (N_835,In_910,N_610);
and U836 (N_836,In_1388,N_511);
or U837 (N_837,In_231,N_27);
nand U838 (N_838,In_151,In_1335);
nand U839 (N_839,In_746,N_106);
xnor U840 (N_840,In_887,In_1951);
nor U841 (N_841,In_1713,N_736);
xor U842 (N_842,N_133,N_85);
nor U843 (N_843,N_465,In_33);
xnor U844 (N_844,In_848,In_605);
and U845 (N_845,In_854,In_1328);
xor U846 (N_846,In_1272,In_1562);
xnor U847 (N_847,In_1365,In_165);
or U848 (N_848,N_682,In_1780);
nand U849 (N_849,N_659,N_554);
nand U850 (N_850,In_844,N_551);
nand U851 (N_851,N_94,In_1746);
or U852 (N_852,N_517,In_1946);
and U853 (N_853,In_1696,N_724);
nor U854 (N_854,In_1684,In_645);
and U855 (N_855,N_569,In_317);
nand U856 (N_856,N_681,In_533);
nand U857 (N_857,N_632,In_112);
xnor U858 (N_858,In_1241,In_172);
or U859 (N_859,In_1440,N_332);
nand U860 (N_860,N_264,In_341);
nand U861 (N_861,N_335,N_355);
nand U862 (N_862,N_239,N_361);
and U863 (N_863,In_1123,In_425);
nand U864 (N_864,N_384,In_1823);
xnor U865 (N_865,N_589,N_583);
or U866 (N_866,N_479,In_363);
xnor U867 (N_867,N_534,In_930);
nor U868 (N_868,In_1108,In_290);
xor U869 (N_869,In_205,N_618);
nand U870 (N_870,N_483,N_689);
xor U871 (N_871,In_1316,In_662);
xor U872 (N_872,N_638,In_1434);
nand U873 (N_873,In_690,In_1617);
or U874 (N_874,In_561,In_577);
or U875 (N_875,In_954,In_1275);
or U876 (N_876,N_404,In_325);
xnor U877 (N_877,N_706,N_609);
xor U878 (N_878,In_1071,In_1230);
and U879 (N_879,N_522,In_393);
and U880 (N_880,N_700,In_1209);
or U881 (N_881,N_24,In_1705);
and U882 (N_882,N_277,N_392);
nor U883 (N_883,In_1954,In_1822);
nor U884 (N_884,In_537,N_745);
and U885 (N_885,In_107,In_894);
nor U886 (N_886,N_23,In_1903);
or U887 (N_887,N_352,In_1753);
and U888 (N_888,In_1045,N_126);
xor U889 (N_889,N_440,N_591);
or U890 (N_890,In_1260,N_278);
nor U891 (N_891,In_263,In_709);
nor U892 (N_892,In_1786,In_471);
xor U893 (N_893,N_611,N_663);
and U894 (N_894,In_734,In_1962);
and U895 (N_895,In_1118,N_717);
xor U896 (N_896,In_1758,N_660);
nor U897 (N_897,In_1520,In_1228);
nor U898 (N_898,In_1039,In_268);
nor U899 (N_899,N_254,In_1278);
and U900 (N_900,N_545,In_1502);
xor U901 (N_901,N_513,N_541);
and U902 (N_902,N_435,N_109);
or U903 (N_903,In_421,In_189);
nor U904 (N_904,In_339,N_670);
nor U905 (N_905,N_189,N_445);
xor U906 (N_906,In_304,In_885);
or U907 (N_907,In_1152,N_653);
nand U908 (N_908,In_1799,In_1411);
nor U909 (N_909,N_744,In_34);
nand U910 (N_910,N_272,In_36);
or U911 (N_911,In_990,In_778);
and U912 (N_912,In_355,In_237);
and U913 (N_913,In_1884,In_1099);
xor U914 (N_914,In_1162,N_114);
and U915 (N_915,N_135,N_431);
or U916 (N_916,In_1271,N_596);
nor U917 (N_917,In_16,N_11);
nor U918 (N_918,In_353,N_448);
and U919 (N_919,In_1994,In_604);
and U920 (N_920,N_686,N_261);
xor U921 (N_921,In_872,N_709);
nand U922 (N_922,In_530,In_261);
nand U923 (N_923,In_173,In_272);
or U924 (N_924,In_536,In_1319);
nand U925 (N_925,In_0,In_1524);
xor U926 (N_926,N_304,In_1652);
and U927 (N_927,In_1629,In_1808);
nor U928 (N_928,In_1787,In_1481);
nor U929 (N_929,In_1500,N_729);
xor U930 (N_930,N_36,N_711);
nand U931 (N_931,In_94,N_654);
xnor U932 (N_932,In_1193,N_219);
xor U933 (N_933,In_60,In_254);
nand U934 (N_934,N_467,N_288);
xor U935 (N_935,N_255,In_1102);
xor U936 (N_936,N_740,N_357);
nor U937 (N_937,In_1330,In_575);
nor U938 (N_938,N_550,In_1888);
nand U939 (N_939,In_1426,In_58);
nor U940 (N_940,In_207,N_624);
nor U941 (N_941,In_55,N_726);
or U942 (N_942,N_742,In_1953);
nor U943 (N_943,N_29,N_416);
nand U944 (N_944,In_1094,In_103);
nor U945 (N_945,In_396,N_282);
xor U946 (N_946,In_586,N_372);
nor U947 (N_947,In_239,In_507);
nand U948 (N_948,In_1896,In_1472);
and U949 (N_949,N_271,In_118);
nor U950 (N_950,In_1208,In_723);
or U951 (N_951,In_932,N_156);
xor U952 (N_952,In_287,N_518);
nor U953 (N_953,In_1408,N_41);
nor U954 (N_954,N_512,In_1416);
and U955 (N_955,In_966,N_316);
xnor U956 (N_956,In_774,In_346);
and U957 (N_957,N_499,N_300);
and U958 (N_958,In_830,N_544);
nand U959 (N_959,In_1480,N_55);
nand U960 (N_960,N_424,In_1459);
and U961 (N_961,In_411,N_308);
nand U962 (N_962,In_1699,N_68);
nand U963 (N_963,N_61,In_741);
or U964 (N_964,In_470,In_822);
xor U965 (N_965,In_725,In_1238);
or U966 (N_966,In_106,In_931);
xor U967 (N_967,In_434,In_68);
nand U968 (N_968,N_412,In_631);
nand U969 (N_969,N_644,In_251);
xor U970 (N_970,In_1206,In_464);
nor U971 (N_971,N_576,In_1718);
nand U972 (N_972,N_695,In_442);
nor U973 (N_973,N_473,N_501);
nor U974 (N_974,In_72,N_540);
xnor U975 (N_975,N_116,N_705);
nor U976 (N_976,N_505,N_602);
nor U977 (N_977,N_32,In_351);
nand U978 (N_978,In_889,N_205);
nor U979 (N_979,N_564,N_196);
or U980 (N_980,In_824,In_1774);
nand U981 (N_981,In_1926,In_1893);
nand U982 (N_982,In_1341,In_950);
or U983 (N_983,In_1243,In_1872);
xor U984 (N_984,N_378,In_1979);
nor U985 (N_985,In_78,In_1687);
xor U986 (N_986,N_421,In_477);
xnor U987 (N_987,In_1898,In_1912);
xnor U988 (N_988,In_694,N_92);
or U989 (N_989,In_1689,In_1909);
nor U990 (N_990,N_104,In_144);
and U991 (N_991,N_444,In_1338);
xor U992 (N_992,N_568,In_807);
nor U993 (N_993,N_374,In_956);
and U994 (N_994,N_697,In_1268);
nor U995 (N_995,In_1283,N_558);
or U996 (N_996,In_1584,N_664);
nand U997 (N_997,In_469,In_1327);
nand U998 (N_998,In_698,N_712);
and U999 (N_999,In_1504,In_1769);
and U1000 (N_1000,N_733,In_1013);
and U1001 (N_1001,N_852,In_1867);
and U1002 (N_1002,In_279,N_96);
or U1003 (N_1003,N_869,In_1450);
nand U1004 (N_1004,In_307,N_893);
or U1005 (N_1005,In_682,In_1114);
xnor U1006 (N_1006,N_266,In_1227);
nor U1007 (N_1007,In_1707,N_983);
xor U1008 (N_1008,In_1564,In_69);
xor U1009 (N_1009,In_139,N_748);
xnor U1010 (N_1010,N_600,N_136);
nand U1011 (N_1011,In_242,N_803);
nand U1012 (N_1012,In_486,In_1551);
xnor U1013 (N_1013,In_663,In_508);
nor U1014 (N_1014,N_715,In_291);
xor U1015 (N_1015,In_1420,In_1028);
xor U1016 (N_1016,In_1589,N_330);
and U1017 (N_1017,In_1191,In_705);
nor U1018 (N_1018,In_1424,N_553);
nand U1019 (N_1019,N_145,N_51);
nand U1020 (N_1020,In_1836,In_274);
or U1021 (N_1021,N_685,In_775);
and U1022 (N_1022,N_884,N_959);
nor U1023 (N_1023,N_827,In_309);
nand U1024 (N_1024,N_851,N_454);
or U1025 (N_1025,In_1362,N_430);
nand U1026 (N_1026,N_181,N_723);
xor U1027 (N_1027,N_25,N_950);
and U1028 (N_1028,N_783,N_459);
nor U1029 (N_1029,N_521,In_1432);
nor U1030 (N_1030,In_1775,N_180);
nor U1031 (N_1031,In_432,N_971);
or U1032 (N_1032,N_888,N_765);
or U1033 (N_1033,In_933,In_1838);
nand U1034 (N_1034,N_646,In_1051);
nand U1035 (N_1035,N_580,In_1430);
xnor U1036 (N_1036,In_1385,N_728);
or U1037 (N_1037,N_900,N_668);
or U1038 (N_1038,N_396,N_832);
and U1039 (N_1039,N_35,N_529);
and U1040 (N_1040,N_957,N_358);
or U1041 (N_1041,In_512,N_792);
nor U1042 (N_1042,N_775,N_794);
nor U1043 (N_1043,In_81,In_1059);
xor U1044 (N_1044,N_981,In_275);
nor U1045 (N_1045,N_634,N_798);
xnor U1046 (N_1046,In_955,N_842);
or U1047 (N_1047,N_8,N_874);
xnor U1048 (N_1048,N_749,In_201);
or U1049 (N_1049,In_1591,N_767);
nand U1050 (N_1050,In_638,In_1292);
nor U1051 (N_1051,N_898,N_830);
nor U1052 (N_1052,N_676,N_933);
and U1053 (N_1053,In_405,N_575);
nand U1054 (N_1054,N_72,In_1469);
xnor U1055 (N_1055,In_1339,N_912);
or U1056 (N_1056,N_649,In_204);
or U1057 (N_1057,N_469,In_175);
and U1058 (N_1058,In_1213,In_1712);
and U1059 (N_1059,In_1982,N_190);
xnor U1060 (N_1060,In_1876,In_53);
or U1061 (N_1061,N_191,In_913);
nor U1062 (N_1062,N_515,N_401);
xor U1063 (N_1063,N_639,In_1070);
nor U1064 (N_1064,In_108,In_1140);
nor U1065 (N_1065,N_75,In_1244);
nand U1066 (N_1066,N_878,N_621);
xnor U1067 (N_1067,N_821,N_891);
nand U1068 (N_1068,N_652,In_676);
and U1069 (N_1069,N_419,N_510);
nor U1070 (N_1070,N_687,N_994);
or U1071 (N_1071,N_566,N_947);
nand U1072 (N_1072,N_790,N_968);
nor U1073 (N_1073,N_781,In_1180);
nor U1074 (N_1074,N_967,N_915);
xor U1075 (N_1075,N_294,N_956);
nor U1076 (N_1076,In_313,In_465);
nand U1077 (N_1077,N_902,N_39);
nand U1078 (N_1078,N_831,N_64);
nand U1079 (N_1079,N_816,In_382);
xnor U1080 (N_1080,N_990,In_159);
and U1081 (N_1081,In_1635,N_298);
and U1082 (N_1082,N_927,In_131);
or U1083 (N_1083,In_357,N_275);
and U1084 (N_1084,N_507,In_420);
xnor U1085 (N_1085,In_1959,In_113);
and U1086 (N_1086,In_1406,In_1471);
and U1087 (N_1087,In_1234,N_301);
nand U1088 (N_1088,N_828,N_606);
and U1089 (N_1089,N_673,N_845);
xor U1090 (N_1090,N_492,N_211);
nand U1091 (N_1091,N_322,In_936);
and U1092 (N_1092,In_1724,N_813);
and U1093 (N_1093,In_752,N_849);
or U1094 (N_1094,N_690,N_797);
xnor U1095 (N_1095,N_963,In_1196);
and U1096 (N_1096,N_658,In_1394);
nand U1097 (N_1097,In_1593,In_651);
or U1098 (N_1098,N_917,N_201);
nand U1099 (N_1099,In_1072,In_1630);
xor U1100 (N_1100,N_389,In_42);
nor U1101 (N_1101,N_556,In_1478);
nand U1102 (N_1102,N_984,In_154);
or U1103 (N_1103,N_43,N_631);
nor U1104 (N_1104,N_333,N_817);
and U1105 (N_1105,N_987,N_242);
xnor U1106 (N_1106,N_970,N_584);
xnor U1107 (N_1107,N_672,N_820);
nand U1108 (N_1108,N_597,N_693);
xor U1109 (N_1109,In_1918,N_887);
or U1110 (N_1110,In_1360,N_771);
nor U1111 (N_1111,N_825,In_1145);
xor U1112 (N_1112,N_54,In_772);
xnor U1113 (N_1113,In_492,In_223);
or U1114 (N_1114,In_18,N_976);
nor U1115 (N_1115,N_871,N_296);
and U1116 (N_1116,In_1863,N_7);
xor U1117 (N_1117,In_1984,In_1304);
or U1118 (N_1118,N_978,N_637);
nor U1119 (N_1119,N_696,N_721);
nand U1120 (N_1120,In_539,N_487);
nand U1121 (N_1121,N_81,N_940);
nor U1122 (N_1122,In_755,N_703);
or U1123 (N_1123,N_367,In_1255);
nand U1124 (N_1124,N_393,N_629);
xnor U1125 (N_1125,In_384,N_523);
or U1126 (N_1126,N_752,N_111);
and U1127 (N_1127,N_630,In_992);
nor U1128 (N_1128,In_89,N_769);
xor U1129 (N_1129,In_447,N_823);
nor U1130 (N_1130,In_1166,N_107);
nor U1131 (N_1131,N_934,In_1765);
or U1132 (N_1132,N_552,N_880);
or U1133 (N_1133,In_1150,N_291);
nand U1134 (N_1134,N_588,N_850);
or U1135 (N_1135,In_819,In_927);
xnor U1136 (N_1136,N_97,N_115);
nand U1137 (N_1137,In_1419,N_636);
and U1138 (N_1138,N_937,In_1586);
and U1139 (N_1139,N_834,N_906);
xor U1140 (N_1140,In_1782,N_166);
or U1141 (N_1141,In_1969,In_157);
and U1142 (N_1142,In_666,N_911);
xor U1143 (N_1143,N_928,N_325);
nand U1144 (N_1144,N_848,N_528);
and U1145 (N_1145,N_691,N_809);
or U1146 (N_1146,In_1862,N_443);
nand U1147 (N_1147,In_809,N_102);
nor U1148 (N_1148,In_1639,In_608);
and U1149 (N_1149,In_1486,N_525);
or U1150 (N_1150,In_1747,In_171);
nor U1151 (N_1151,N_605,N_65);
nor U1152 (N_1152,N_867,N_908);
nand U1153 (N_1153,N_669,N_47);
and U1154 (N_1154,N_675,In_1751);
nand U1155 (N_1155,N_815,N_808);
nand U1156 (N_1156,In_576,N_433);
or U1157 (N_1157,N_470,In_859);
and U1158 (N_1158,In_1199,In_1008);
or U1159 (N_1159,N_811,In_29);
xor U1160 (N_1160,N_796,N_643);
nand U1161 (N_1161,In_1224,In_302);
nand U1162 (N_1162,N_197,N_899);
or U1163 (N_1163,N_527,N_577);
and U1164 (N_1164,In_1757,N_647);
nand U1165 (N_1165,N_279,N_623);
xnor U1166 (N_1166,N_972,N_349);
or U1167 (N_1167,N_594,N_453);
or U1168 (N_1168,N_910,N_920);
xnor U1169 (N_1169,N_157,N_234);
xnor U1170 (N_1170,In_624,N_599);
and U1171 (N_1171,N_960,N_806);
nor U1172 (N_1172,N_754,In_648);
xor U1173 (N_1173,N_836,In_798);
nor U1174 (N_1174,In_749,In_1819);
xnor U1175 (N_1175,In_64,In_529);
nand U1176 (N_1176,N_992,In_1644);
and U1177 (N_1177,In_257,In_1276);
and U1178 (N_1178,In_771,N_841);
and U1179 (N_1179,In_1158,In_1666);
and U1180 (N_1180,In_197,In_1596);
and U1181 (N_1181,In_1721,In_308);
nor U1182 (N_1182,N_916,In_475);
or U1183 (N_1183,In_754,In_996);
or U1184 (N_1184,N_843,N_312);
or U1185 (N_1185,In_90,N_774);
nor U1186 (N_1186,N_10,N_549);
xor U1187 (N_1187,In_792,In_327);
xnor U1188 (N_1188,In_167,N_678);
xor U1189 (N_1189,N_886,In_739);
and U1190 (N_1190,N_232,In_1453);
nor U1191 (N_1191,In_1811,N_655);
nand U1192 (N_1192,In_381,In_145);
nand U1193 (N_1193,In_1082,N_587);
and U1194 (N_1194,In_1790,N_914);
nand U1195 (N_1195,In_1506,N_770);
nand U1196 (N_1196,N_904,In_1449);
nand U1197 (N_1197,In_917,N_18);
and U1198 (N_1198,N_593,N_710);
or U1199 (N_1199,N_403,N_457);
and U1200 (N_1200,N_826,N_79);
or U1201 (N_1201,N_460,N_683);
xor U1202 (N_1202,N_931,In_794);
nor U1203 (N_1203,In_1032,In_1895);
nand U1204 (N_1204,N_651,N_509);
or U1205 (N_1205,N_614,N_641);
nand U1206 (N_1206,N_951,N_212);
and U1207 (N_1207,N_758,In_1188);
and U1208 (N_1208,N_546,In_1055);
nor U1209 (N_1209,In_784,N_961);
or U1210 (N_1210,In_1111,In_1315);
or U1211 (N_1211,In_1703,In_1023);
and U1212 (N_1212,N_698,N_907);
and U1213 (N_1213,In_453,N_777);
or U1214 (N_1214,In_1291,N_854);
nand U1215 (N_1215,N_716,N_838);
or U1216 (N_1216,In_521,In_1785);
and U1217 (N_1217,In_1612,N_757);
nor U1218 (N_1218,In_57,N_755);
xor U1219 (N_1219,N_57,N_535);
nand U1220 (N_1220,In_176,In_332);
nand U1221 (N_1221,N_442,N_998);
nand U1222 (N_1222,N_868,In_1573);
xnor U1223 (N_1223,N_21,N_881);
nor U1224 (N_1224,N_760,In_1128);
nor U1225 (N_1225,N_799,N_674);
nand U1226 (N_1226,In_757,In_687);
or U1227 (N_1227,N_870,N_877);
xor U1228 (N_1228,In_1197,In_1674);
or U1229 (N_1229,N_351,N_807);
nor U1230 (N_1230,N_945,In_1949);
or U1231 (N_1231,In_1371,N_601);
and U1232 (N_1232,N_901,N_598);
nor U1233 (N_1233,N_612,In_1143);
or U1234 (N_1234,N_890,N_865);
and U1235 (N_1235,N_559,N_768);
and U1236 (N_1236,In_1022,N_954);
xnor U1237 (N_1237,In_1331,N_948);
nor U1238 (N_1238,N_995,In_1742);
xor U1239 (N_1239,In_1004,N_732);
xor U1240 (N_1240,N_692,N_209);
nand U1241 (N_1241,N_263,N_883);
xor U1242 (N_1242,N_819,N_303);
and U1243 (N_1243,N_731,In_1968);
nand U1244 (N_1244,N_149,N_400);
and U1245 (N_1245,N_267,N_840);
nand U1246 (N_1246,N_628,N_451);
xnor U1247 (N_1247,In_574,In_1347);
nor U1248 (N_1248,N_578,N_772);
nand U1249 (N_1249,N_856,N_508);
nand U1250 (N_1250,N_812,N_620);
and U1251 (N_1251,N_1041,N_571);
and U1252 (N_1252,N_635,N_1139);
xnor U1253 (N_1253,In_1282,In_911);
or U1254 (N_1254,N_648,N_1075);
nor U1255 (N_1255,In_95,N_269);
xor U1256 (N_1256,In_1024,In_1760);
nand U1257 (N_1257,N_455,N_1056);
or U1258 (N_1258,In_6,N_1051);
or U1259 (N_1259,In_1149,In_1076);
xnor U1260 (N_1260,In_804,N_354);
xor U1261 (N_1261,In_1270,N_1130);
or U1262 (N_1262,In_763,N_1049);
or U1263 (N_1263,N_1090,N_1226);
and U1264 (N_1264,N_1143,N_192);
nor U1265 (N_1265,In_12,N_862);
and U1266 (N_1266,In_1723,N_1039);
xnor U1267 (N_1267,N_1131,In_1800);
and U1268 (N_1268,N_661,N_1021);
nand U1269 (N_1269,In_726,N_895);
or U1270 (N_1270,In_1444,N_805);
or U1271 (N_1271,N_860,N_538);
and U1272 (N_1272,N_1073,N_642);
nor U1273 (N_1273,N_1026,N_722);
xnor U1274 (N_1274,N_186,N_1042);
xnor U1275 (N_1275,N_1054,N_1066);
nor U1276 (N_1276,In_276,In_699);
and U1277 (N_1277,N_864,N_818);
or U1278 (N_1278,N_784,In_407);
xnor U1279 (N_1279,N_1005,In_186);
nand U1280 (N_1280,N_616,N_547);
and U1281 (N_1281,N_938,N_941);
xor U1282 (N_1282,N_789,N_530);
and U1283 (N_1283,N_1105,In_1678);
xor U1284 (N_1284,N_1158,In_372);
or U1285 (N_1285,In_929,N_701);
xnor U1286 (N_1286,In_431,N_1116);
or U1287 (N_1287,N_283,N_615);
or U1288 (N_1288,N_1142,N_1016);
or U1289 (N_1289,In_1691,N_762);
or U1290 (N_1290,In_455,N_1169);
nand U1291 (N_1291,N_491,In_1711);
nand U1292 (N_1292,N_337,N_320);
xnor U1293 (N_1293,N_1135,N_1071);
nand U1294 (N_1294,N_557,N_993);
xor U1295 (N_1295,In_1407,In_1580);
or U1296 (N_1296,In_1550,N_735);
nor U1297 (N_1297,N_1145,N_982);
and U1298 (N_1298,In_590,N_766);
nand U1299 (N_1299,N_1129,In_1084);
or U1300 (N_1300,In_986,N_1153);
or U1301 (N_1301,N_1156,N_1218);
xnor U1302 (N_1302,In_571,In_161);
nand U1303 (N_1303,N_1036,N_1137);
nand U1304 (N_1304,N_863,N_1033);
and U1305 (N_1305,N_751,In_707);
or U1306 (N_1306,In_1046,In_293);
nand U1307 (N_1307,N_1059,In_810);
and U1308 (N_1308,In_296,In_462);
xor U1309 (N_1309,N_1065,N_251);
xnor U1310 (N_1310,In_1693,In_759);
nand U1311 (N_1311,N_1047,N_720);
nand U1312 (N_1312,In_140,N_1223);
or U1313 (N_1313,In_1127,N_855);
or U1314 (N_1314,N_829,In_710);
nor U1315 (N_1315,N_1242,N_1004);
or U1316 (N_1316,In_128,N_1092);
nor U1317 (N_1317,N_463,N_1126);
xnor U1318 (N_1318,N_1248,N_988);
nand U1319 (N_1319,In_1583,N_1219);
xor U1320 (N_1320,N_1089,In_601);
or U1321 (N_1321,N_1178,N_930);
xnor U1322 (N_1322,N_1022,N_894);
and U1323 (N_1323,In_1377,N_1062);
and U1324 (N_1324,N_1233,In_148);
and U1325 (N_1325,N_1076,In_1904);
xor U1326 (N_1326,N_1063,N_974);
nand U1327 (N_1327,N_1053,N_1144);
nand U1328 (N_1328,N_905,In_1095);
or U1329 (N_1329,In_1945,In_1999);
xor U1330 (N_1330,N_977,N_1070);
nand U1331 (N_1331,N_1229,N_1162);
xor U1332 (N_1332,N_203,N_432);
nand U1333 (N_1333,In_1309,N_1157);
xnor U1334 (N_1334,N_377,N_171);
and U1335 (N_1335,In_606,N_943);
or U1336 (N_1336,In_737,N_327);
nand U1337 (N_1337,In_1016,In_923);
xor U1338 (N_1338,In_612,In_14);
and U1339 (N_1339,In_1237,N_918);
or U1340 (N_1340,N_1154,In_688);
or U1341 (N_1341,In_1604,N_991);
nor U1342 (N_1342,N_926,N_1182);
xor U1343 (N_1343,N_802,N_466);
xor U1344 (N_1344,N_879,N_778);
nand U1345 (N_1345,N_1111,N_921);
or U1346 (N_1346,N_297,N_793);
nand U1347 (N_1347,N_1007,N_924);
xnor U1348 (N_1348,N_885,In_235);
nor U1349 (N_1349,N_814,N_1074);
and U1350 (N_1350,N_824,In_801);
xor U1351 (N_1351,N_1238,N_801);
nand U1352 (N_1352,N_1086,N_889);
nor U1353 (N_1353,In_1254,N_233);
and U1354 (N_1354,N_985,In_92);
nand U1355 (N_1355,N_955,N_1055);
and U1356 (N_1356,N_922,In_1676);
and U1357 (N_1357,In_847,N_944);
nor U1358 (N_1358,N_585,N_1196);
nor U1359 (N_1359,N_309,N_218);
nor U1360 (N_1360,In_883,N_306);
nor U1361 (N_1361,In_1068,N_1184);
nand U1362 (N_1362,N_800,N_1064);
xnor U1363 (N_1363,N_1177,N_1106);
nor U1364 (N_1364,N_604,N_1241);
nand U1365 (N_1365,N_147,In_944);
or U1366 (N_1366,N_562,N_750);
nor U1367 (N_1367,N_200,In_857);
xnor U1368 (N_1368,N_1175,N_882);
and U1369 (N_1369,In_839,N_336);
nor U1370 (N_1370,N_1136,N_1220);
and U1371 (N_1371,N_747,N_1037);
or U1372 (N_1372,N_1079,N_495);
nand U1373 (N_1373,N_665,N_1122);
nor U1374 (N_1374,In_1131,In_1940);
and U1375 (N_1375,In_658,In_1847);
or U1376 (N_1376,N_1206,N_516);
and U1377 (N_1377,In_1030,N_1155);
and U1378 (N_1378,N_33,In_1928);
or U1379 (N_1379,N_753,N_776);
nand U1380 (N_1380,N_833,N_804);
xnor U1381 (N_1381,N_1043,N_313);
nor U1382 (N_1382,N_1085,N_607);
nand U1383 (N_1383,N_713,In_1369);
and U1384 (N_1384,In_1231,In_1467);
or U1385 (N_1385,N_531,N_1020);
and U1386 (N_1386,In_380,In_47);
or U1387 (N_1387,N_837,In_1817);
nand U1388 (N_1388,N_1015,In_1559);
xor U1389 (N_1389,In_1653,In_248);
nand U1390 (N_1390,N_964,In_369);
xnor U1391 (N_1391,N_281,In_350);
nand U1392 (N_1392,In_1527,In_646);
nand U1393 (N_1393,In_738,N_394);
nand U1394 (N_1394,N_791,N_1179);
and U1395 (N_1395,In_1349,N_1045);
nand U1396 (N_1396,N_708,N_714);
or U1397 (N_1397,In_1914,N_1152);
nand U1398 (N_1398,N_626,N_1237);
xor U1399 (N_1399,In_491,N_1030);
xnor U1400 (N_1400,N_307,N_759);
nor U1401 (N_1401,In_322,N_1080);
or U1402 (N_1402,In_1997,N_461);
xor U1403 (N_1403,N_625,In_452);
nor U1404 (N_1404,N_1095,In_35);
xnor U1405 (N_1405,N_265,N_1120);
nor U1406 (N_1406,N_835,N_1232);
or U1407 (N_1407,N_997,N_1060);
and U1408 (N_1408,In_1609,N_343);
nor U1409 (N_1409,N_302,N_567);
xnor U1410 (N_1410,N_873,N_785);
nor U1411 (N_1411,N_1061,N_1217);
or U1412 (N_1412,N_847,N_1201);
and U1413 (N_1413,In_1579,In_1425);
and U1414 (N_1414,In_187,In_1468);
and U1415 (N_1415,N_1191,In_169);
or U1416 (N_1416,N_1038,N_150);
or U1417 (N_1417,In_1091,N_866);
or U1418 (N_1418,N_1104,In_793);
nand U1419 (N_1419,N_795,In_766);
and U1420 (N_1420,N_179,N_1040);
nand U1421 (N_1421,N_1082,N_1151);
or U1422 (N_1422,In_964,N_12);
nand U1423 (N_1423,N_137,In_1935);
nor U1424 (N_1424,N_684,N_532);
xor U1425 (N_1425,In_1489,N_1176);
and U1426 (N_1426,In_1971,In_1129);
nor U1427 (N_1427,N_1173,N_572);
or U1428 (N_1428,N_727,N_756);
nor U1429 (N_1429,N_1215,N_1138);
or U1430 (N_1430,N_536,N_1197);
nor U1431 (N_1431,N_1189,N_574);
nand U1432 (N_1432,N_932,N_1121);
xnor U1433 (N_1433,In_424,In_1279);
and U1434 (N_1434,N_1212,N_694);
nand U1435 (N_1435,In_218,N_1024);
nor U1436 (N_1436,N_1208,N_857);
or U1437 (N_1437,N_1008,N_1210);
and U1438 (N_1438,N_488,N_441);
xor U1439 (N_1439,N_1046,In_1060);
and U1440 (N_1440,N_603,N_1246);
and U1441 (N_1441,N_699,In_484);
or U1442 (N_1442,N_782,N_1203);
nand U1443 (N_1443,N_398,In_76);
or U1444 (N_1444,N_356,N_1235);
and U1445 (N_1445,N_344,N_1165);
nor U1446 (N_1446,N_379,N_1140);
or U1447 (N_1447,N_645,N_573);
xnor U1448 (N_1448,N_953,In_1661);
xor U1449 (N_1449,N_1190,N_1186);
nor U1450 (N_1450,N_1174,In_1164);
xor U1451 (N_1451,In_1542,N_1147);
nand U1452 (N_1452,In_1106,N_1134);
nand U1453 (N_1453,N_969,In_1981);
xor U1454 (N_1454,N_1124,N_338);
and U1455 (N_1455,N_1185,N_1097);
xnor U1456 (N_1456,N_939,N_1107);
nand U1457 (N_1457,N_822,In_984);
and U1458 (N_1458,In_1578,N_542);
or U1459 (N_1459,In_563,In_134);
nor U1460 (N_1460,N_1192,N_246);
nor U1461 (N_1461,N_1231,N_1023);
xor U1462 (N_1462,N_1166,N_909);
or U1463 (N_1463,N_1087,In_617);
nand U1464 (N_1464,N_1222,In_1333);
xor U1465 (N_1465,N_555,N_1011);
and U1466 (N_1466,In_1353,In_1010);
nand U1467 (N_1467,N_1093,In_678);
nor U1468 (N_1468,N_1035,In_1097);
and U1469 (N_1469,N_1193,In_1181);
xnor U1470 (N_1470,N_1249,N_426);
or U1471 (N_1471,N_973,N_1028);
or U1472 (N_1472,N_1044,In_1567);
and U1473 (N_1473,In_1329,N_746);
nand U1474 (N_1474,N_1012,In_1351);
nand U1475 (N_1475,N_26,N_859);
nor U1476 (N_1476,In_546,In_1293);
nand U1477 (N_1477,N_561,N_980);
or U1478 (N_1478,N_965,In_116);
or U1479 (N_1479,N_936,N_1132);
xor U1480 (N_1480,N_1209,N_382);
or U1481 (N_1481,N_764,In_999);
or U1482 (N_1482,In_637,N_198);
nand U1483 (N_1483,N_680,N_861);
nand U1484 (N_1484,N_1050,N_475);
nor U1485 (N_1485,N_996,In_1533);
nor U1486 (N_1486,In_1501,N_773);
nand U1487 (N_1487,N_1234,In_1794);
xnor U1488 (N_1488,N_903,In_1135);
xnor U1489 (N_1489,N_1057,In_400);
nor U1490 (N_1490,N_592,N_779);
nand U1491 (N_1491,N_1183,N_1101);
xor U1492 (N_1492,N_1025,N_1109);
nand U1493 (N_1493,In_649,In_375);
xor U1494 (N_1494,In_1443,N_1110);
nor U1495 (N_1495,In_783,In_1773);
and U1496 (N_1496,N_490,In_27);
or U1497 (N_1497,In_1491,In_137);
xor U1498 (N_1498,In_337,N_290);
or U1499 (N_1499,N_741,N_1228);
or U1500 (N_1500,N_1188,N_1492);
and U1501 (N_1501,In_1733,N_1406);
and U1502 (N_1502,N_1357,N_350);
or U1503 (N_1503,N_1420,N_524);
nor U1504 (N_1504,N_76,N_896);
and U1505 (N_1505,N_1475,N_1264);
or U1506 (N_1506,N_1481,N_1251);
xor U1507 (N_1507,N_1440,In_552);
and U1508 (N_1508,N_1245,N_1423);
nand U1509 (N_1509,N_1432,N_1279);
and U1510 (N_1510,N_1362,N_1255);
and U1511 (N_1511,In_846,In_1582);
nand U1512 (N_1512,N_1393,N_962);
nand U1513 (N_1513,N_1254,N_1069);
or U1514 (N_1514,N_1195,N_1150);
nor U1515 (N_1515,N_1052,N_1358);
and U1516 (N_1516,N_667,N_1290);
and U1517 (N_1517,N_1403,N_1390);
xor U1518 (N_1518,N_1017,N_284);
nor U1519 (N_1519,N_1010,In_558);
nand U1520 (N_1520,N_725,In_1448);
xnor U1521 (N_1521,N_15,N_1431);
xor U1522 (N_1522,N_1384,In_787);
and U1523 (N_1523,In_1706,In_1);
nor U1524 (N_1524,N_1364,N_1276);
and U1525 (N_1525,N_1375,N_339);
nor U1526 (N_1526,N_537,N_1417);
xnor U1527 (N_1527,N_846,N_1100);
and U1528 (N_1528,In_1052,N_633);
and U1529 (N_1529,N_1058,N_650);
nand U1530 (N_1530,N_1259,N_1214);
xor U1531 (N_1531,N_1263,N_158);
or U1532 (N_1532,N_1205,N_1455);
nand U1533 (N_1533,N_1293,N_613);
or U1534 (N_1534,N_1252,N_671);
and U1535 (N_1535,N_1485,In_660);
or U1536 (N_1536,In_621,N_1345);
or U1537 (N_1537,N_1376,N_493);
xnor U1538 (N_1538,N_514,N_1227);
and U1539 (N_1539,N_1172,N_1311);
xor U1540 (N_1540,N_390,In_661);
xnor U1541 (N_1541,N_1014,N_1003);
or U1542 (N_1542,N_1283,N_1336);
nor U1543 (N_1543,N_1412,N_923);
xor U1544 (N_1544,N_1404,N_989);
xor U1545 (N_1545,N_1434,N_1330);
nor U1546 (N_1546,N_1298,In_768);
nand U1547 (N_1547,N_1489,N_1318);
or U1548 (N_1548,N_1310,N_1495);
xnor U1549 (N_1549,N_935,N_1468);
xnor U1550 (N_1550,N_1446,N_679);
and U1551 (N_1551,N_1094,N_1148);
xor U1552 (N_1552,N_1449,N_1299);
and U1553 (N_1553,N_1001,N_1244);
nand U1554 (N_1554,N_1284,N_853);
and U1555 (N_1555,N_1401,N_1103);
xnor U1556 (N_1556,N_1427,N_1352);
nand U1557 (N_1557,N_1114,In_21);
and U1558 (N_1558,N_1353,N_581);
or U1559 (N_1559,N_1378,N_1474);
nand U1560 (N_1560,N_704,N_1447);
nor U1561 (N_1561,N_1398,N_1360);
or U1562 (N_1562,N_1307,N_19);
nor U1563 (N_1563,N_1077,N_1425);
or U1564 (N_1564,N_1277,N_1445);
nor U1565 (N_1565,In_125,N_482);
nand U1566 (N_1566,N_1493,In_1446);
nor U1567 (N_1567,N_1411,N_1170);
xor U1568 (N_1568,N_999,N_345);
nand U1569 (N_1569,N_1084,N_1479);
or U1570 (N_1570,N_786,N_1236);
nand U1571 (N_1571,In_871,N_1338);
nand U1572 (N_1572,In_818,N_925);
xnor U1573 (N_1573,N_1312,N_1102);
xnor U1574 (N_1574,N_1324,N_1316);
or U1575 (N_1575,N_1302,N_1395);
nand U1576 (N_1576,In_233,N_1473);
nand U1577 (N_1577,N_1099,N_1303);
nor U1578 (N_1578,N_986,N_913);
xor U1579 (N_1579,N_1443,N_1400);
and U1580 (N_1580,In_1977,In_122);
nor U1581 (N_1581,N_1436,N_1018);
xor U1582 (N_1582,N_227,In_942);
or U1583 (N_1583,N_1442,N_1415);
nor U1584 (N_1584,N_1341,In_1736);
xnor U1585 (N_1585,N_208,N_1159);
nor U1586 (N_1586,N_1346,N_1450);
nor U1587 (N_1587,In_835,N_1292);
xnor U1588 (N_1588,In_1795,N_1413);
and U1589 (N_1589,N_1439,N_1239);
xor U1590 (N_1590,N_702,N_1300);
nand U1591 (N_1591,N_1262,N_1216);
and U1592 (N_1592,N_1477,N_1315);
and U1593 (N_1593,N_1272,In_1375);
nor U1594 (N_1594,N_586,N_1213);
xnor U1595 (N_1595,N_28,N_1367);
xor U1596 (N_1596,N_1112,N_875);
nor U1597 (N_1597,N_1305,In_1277);
nor U1598 (N_1598,N_1032,N_1340);
and U1599 (N_1599,N_1194,N_1359);
xnor U1600 (N_1600,N_1181,N_1348);
xnor U1601 (N_1601,N_1462,N_1289);
nand U1602 (N_1602,N_1392,N_1287);
xnor U1603 (N_1603,N_1332,N_1207);
and U1604 (N_1604,N_1379,N_1471);
nor U1605 (N_1605,N_1428,In_951);
nand U1606 (N_1606,N_1418,N_1383);
or U1607 (N_1607,N_348,N_1499);
and U1608 (N_1608,N_1117,N_780);
xnor U1609 (N_1609,N_929,N_1119);
or U1610 (N_1610,N_958,N_1133);
xor U1611 (N_1611,N_788,N_1366);
nand U1612 (N_1612,N_1354,N_1266);
or U1613 (N_1613,In_1616,In_567);
and U1614 (N_1614,N_1437,N_1230);
nor U1615 (N_1615,N_1271,N_1270);
nand U1616 (N_1616,N_1247,In_603);
and U1617 (N_1617,N_1281,N_1002);
or U1618 (N_1618,N_919,N_520);
nor U1619 (N_1619,N_1261,N_1325);
and U1620 (N_1620,In_788,N_1088);
and U1621 (N_1621,N_1006,N_1484);
nand U1622 (N_1622,N_1288,N_1329);
xor U1623 (N_1623,N_1396,N_892);
and U1624 (N_1624,N_1200,N_1146);
or U1625 (N_1625,N_560,In_915);
and U1626 (N_1626,N_1337,In_1752);
nor U1627 (N_1627,N_1160,N_975);
and U1628 (N_1628,N_1202,N_1260);
nand U1629 (N_1629,N_1350,N_1451);
or U1630 (N_1630,In_284,N_1452);
nor U1631 (N_1631,N_1373,N_949);
nand U1632 (N_1632,N_1072,N_1257);
or U1633 (N_1633,N_1370,In_1605);
xor U1634 (N_1634,N_718,N_1490);
nand U1635 (N_1635,N_1441,N_1430);
xnor U1636 (N_1636,N_1211,N_1083);
nor U1637 (N_1637,N_1399,In_371);
and U1638 (N_1638,In_922,N_1433);
xor U1639 (N_1639,N_1308,N_1331);
xor U1640 (N_1640,N_1274,N_1342);
and U1641 (N_1641,In_1776,In_1269);
or U1642 (N_1642,N_1389,N_159);
nand U1643 (N_1643,N_1108,N_1465);
nand U1644 (N_1644,N_1171,N_1328);
nand U1645 (N_1645,N_1323,N_761);
xnor U1646 (N_1646,N_1448,N_1027);
nor U1647 (N_1647,N_1361,N_1067);
xnor U1648 (N_1648,N_1301,N_1161);
nand U1649 (N_1649,N_876,N_1013);
nor U1650 (N_1650,In_657,N_415);
nor U1651 (N_1651,In_417,N_347);
nor U1652 (N_1652,N_952,N_897);
nand U1653 (N_1653,N_1459,N_1466);
nor U1654 (N_1654,N_1326,N_1355);
or U1655 (N_1655,N_1296,N_1369);
and U1656 (N_1656,N_376,In_1944);
nor U1657 (N_1657,In_1726,N_738);
nand U1658 (N_1658,N_1344,N_1335);
nand U1659 (N_1659,N_787,N_1460);
or U1660 (N_1660,N_1294,N_1243);
or U1661 (N_1661,N_1167,N_666);
xnor U1662 (N_1662,N_1081,N_1461);
and U1663 (N_1663,N_1282,N_1031);
nand U1664 (N_1664,N_1019,N_1327);
xnor U1665 (N_1665,N_1347,In_298);
xnor U1666 (N_1666,N_1494,N_1444);
xnor U1667 (N_1667,N_1421,N_1320);
xnor U1668 (N_1668,N_1048,N_1168);
or U1669 (N_1669,N_1422,N_1382);
and U1670 (N_1670,N_1374,N_565);
nand U1671 (N_1671,N_1269,N_1187);
nor U1672 (N_1672,N_1454,N_872);
nor U1673 (N_1673,In_1175,N_570);
nor U1674 (N_1674,In_1176,N_1204);
xnor U1675 (N_1675,N_223,N_1125);
nand U1676 (N_1676,N_1469,N_1297);
and U1677 (N_1677,N_1068,N_1405);
and U1678 (N_1678,N_1416,N_1322);
and U1679 (N_1679,N_1334,N_1000);
and U1680 (N_1680,N_1397,N_1394);
xor U1681 (N_1681,N_1113,N_1410);
nor U1682 (N_1682,In_1182,N_1391);
nand U1683 (N_1683,N_1457,In_1650);
xnor U1684 (N_1684,In_1964,N_1317);
nor U1685 (N_1685,N_1256,N_1333);
or U1686 (N_1686,N_1319,N_1096);
nor U1687 (N_1687,N_1240,N_1488);
xor U1688 (N_1688,N_1078,N_1268);
or U1689 (N_1689,N_1225,N_1275);
or U1690 (N_1690,N_1273,N_1424);
xnor U1691 (N_1691,N_966,N_1034);
or U1692 (N_1692,N_839,N_1343);
and U1693 (N_1693,N_1123,N_1483);
nor U1694 (N_1694,N_1456,In_253);
and U1695 (N_1695,N_1009,N_1339);
nand U1696 (N_1696,N_662,N_810);
nand U1697 (N_1697,N_1118,N_229);
nand U1698 (N_1698,N_1115,N_1381);
xor U1699 (N_1699,N_1128,In_1493);
nand U1700 (N_1700,N_1498,N_1372);
nor U1701 (N_1701,N_1470,N_1407);
nor U1702 (N_1702,N_1487,N_1199);
and U1703 (N_1703,N_1091,N_1365);
and U1704 (N_1704,N_1497,In_441);
xnor U1705 (N_1705,N_1409,N_1029);
nand U1706 (N_1706,N_1309,N_1351);
nand U1707 (N_1707,In_1767,N_844);
nand U1708 (N_1708,N_1321,In_1011);
or U1709 (N_1709,N_1349,N_1098);
xor U1710 (N_1710,N_743,N_858);
nor U1711 (N_1711,N_1163,N_1221);
and U1712 (N_1712,N_1387,In_520);
or U1713 (N_1713,In_1603,N_1314);
xnor U1714 (N_1714,N_1291,N_946);
or U1715 (N_1715,N_1295,N_763);
xor U1716 (N_1716,N_979,N_1280);
nand U1717 (N_1717,N_1164,N_1224);
or U1718 (N_1718,N_1313,N_1304);
nand U1719 (N_1719,N_1198,N_1491);
and U1720 (N_1720,N_1253,N_1267);
nand U1721 (N_1721,In_1452,N_1141);
nand U1722 (N_1722,In_62,N_1402);
or U1723 (N_1723,N_1180,N_1467);
and U1724 (N_1724,N_1265,N_1258);
xnor U1725 (N_1725,N_395,N_326);
nand U1726 (N_1726,N_184,N_1463);
xnor U1727 (N_1727,In_303,N_1127);
or U1728 (N_1728,N_1286,N_1453);
xor U1729 (N_1729,In_1200,N_1368);
or U1730 (N_1730,N_1458,N_1486);
nor U1731 (N_1731,N_1408,N_1285);
and U1732 (N_1732,N_1426,N_1429);
nor U1733 (N_1733,N_1472,N_1278);
nand U1734 (N_1734,N_942,N_1476);
and U1735 (N_1735,N_1478,N_1149);
nand U1736 (N_1736,In_51,N_1363);
nand U1737 (N_1737,In_1855,In_1053);
nor U1738 (N_1738,N_1464,N_1419);
nand U1739 (N_1739,N_360,In_1173);
and U1740 (N_1740,In_1345,N_1250);
nor U1741 (N_1741,N_1482,In_359);
and U1742 (N_1742,N_1385,N_1438);
nand U1743 (N_1743,N_1480,N_1388);
and U1744 (N_1744,N_1377,In_832);
nand U1745 (N_1745,N_533,N_1386);
and U1746 (N_1746,N_1306,N_1356);
xor U1747 (N_1747,N_1371,N_1435);
or U1748 (N_1748,N_1380,N_1414);
nor U1749 (N_1749,In_1136,N_1496);
nor U1750 (N_1750,N_1664,N_1697);
nor U1751 (N_1751,N_1619,N_1696);
nand U1752 (N_1752,N_1516,N_1695);
nand U1753 (N_1753,N_1581,N_1690);
or U1754 (N_1754,N_1513,N_1741);
xor U1755 (N_1755,N_1717,N_1634);
or U1756 (N_1756,N_1507,N_1512);
nand U1757 (N_1757,N_1510,N_1539);
nand U1758 (N_1758,N_1593,N_1746);
nand U1759 (N_1759,N_1635,N_1705);
xnor U1760 (N_1760,N_1527,N_1551);
or U1761 (N_1761,N_1569,N_1682);
and U1762 (N_1762,N_1647,N_1631);
xor U1763 (N_1763,N_1601,N_1629);
or U1764 (N_1764,N_1704,N_1736);
and U1765 (N_1765,N_1677,N_1531);
nand U1766 (N_1766,N_1622,N_1744);
or U1767 (N_1767,N_1567,N_1597);
nor U1768 (N_1768,N_1501,N_1694);
or U1769 (N_1769,N_1596,N_1637);
nand U1770 (N_1770,N_1670,N_1612);
xor U1771 (N_1771,N_1602,N_1609);
xor U1772 (N_1772,N_1541,N_1578);
xnor U1773 (N_1773,N_1520,N_1714);
and U1774 (N_1774,N_1617,N_1608);
nor U1775 (N_1775,N_1623,N_1676);
xnor U1776 (N_1776,N_1639,N_1656);
and U1777 (N_1777,N_1600,N_1522);
or U1778 (N_1778,N_1657,N_1652);
or U1779 (N_1779,N_1614,N_1679);
and U1780 (N_1780,N_1640,N_1745);
nor U1781 (N_1781,N_1687,N_1620);
or U1782 (N_1782,N_1627,N_1698);
nand U1783 (N_1783,N_1646,N_1613);
and U1784 (N_1784,N_1568,N_1731);
and U1785 (N_1785,N_1708,N_1540);
or U1786 (N_1786,N_1724,N_1590);
nor U1787 (N_1787,N_1533,N_1673);
or U1788 (N_1788,N_1665,N_1716);
and U1789 (N_1789,N_1583,N_1505);
xnor U1790 (N_1790,N_1621,N_1538);
nand U1791 (N_1791,N_1562,N_1732);
or U1792 (N_1792,N_1529,N_1740);
nand U1793 (N_1793,N_1651,N_1519);
xnor U1794 (N_1794,N_1643,N_1730);
or U1795 (N_1795,N_1618,N_1584);
or U1796 (N_1796,N_1645,N_1561);
nand U1797 (N_1797,N_1571,N_1712);
xor U1798 (N_1798,N_1591,N_1729);
nand U1799 (N_1799,N_1550,N_1721);
xnor U1800 (N_1800,N_1615,N_1672);
or U1801 (N_1801,N_1699,N_1560);
or U1802 (N_1802,N_1580,N_1675);
nand U1803 (N_1803,N_1532,N_1749);
xnor U1804 (N_1804,N_1728,N_1678);
or U1805 (N_1805,N_1558,N_1517);
nand U1806 (N_1806,N_1521,N_1528);
nand U1807 (N_1807,N_1579,N_1549);
nor U1808 (N_1808,N_1523,N_1589);
nand U1809 (N_1809,N_1570,N_1604);
or U1810 (N_1810,N_1642,N_1603);
xnor U1811 (N_1811,N_1701,N_1625);
or U1812 (N_1812,N_1530,N_1508);
nand U1813 (N_1813,N_1641,N_1607);
nand U1814 (N_1814,N_1534,N_1654);
and U1815 (N_1815,N_1599,N_1706);
or U1816 (N_1816,N_1648,N_1595);
and U1817 (N_1817,N_1518,N_1655);
or U1818 (N_1818,N_1703,N_1537);
or U1819 (N_1819,N_1734,N_1733);
or U1820 (N_1820,N_1628,N_1693);
nand U1821 (N_1821,N_1559,N_1605);
nor U1822 (N_1822,N_1573,N_1725);
nor U1823 (N_1823,N_1686,N_1633);
and U1824 (N_1824,N_1737,N_1711);
nand U1825 (N_1825,N_1552,N_1536);
nor U1826 (N_1826,N_1577,N_1713);
or U1827 (N_1827,N_1525,N_1684);
nor U1828 (N_1828,N_1660,N_1722);
nand U1829 (N_1829,N_1702,N_1606);
and U1830 (N_1830,N_1626,N_1592);
xnor U1831 (N_1831,N_1526,N_1735);
nand U1832 (N_1832,N_1662,N_1739);
xnor U1833 (N_1833,N_1659,N_1547);
or U1834 (N_1834,N_1554,N_1691);
nor U1835 (N_1835,N_1681,N_1587);
nor U1836 (N_1836,N_1720,N_1683);
nand U1837 (N_1837,N_1565,N_1616);
or U1838 (N_1838,N_1658,N_1715);
xnor U1839 (N_1839,N_1543,N_1630);
nor U1840 (N_1840,N_1611,N_1503);
and U1841 (N_1841,N_1556,N_1514);
nor U1842 (N_1842,N_1742,N_1524);
and U1843 (N_1843,N_1511,N_1588);
or U1844 (N_1844,N_1644,N_1632);
xnor U1845 (N_1845,N_1738,N_1535);
nand U1846 (N_1846,N_1564,N_1669);
and U1847 (N_1847,N_1624,N_1563);
and U1848 (N_1848,N_1723,N_1700);
nand U1849 (N_1849,N_1500,N_1663);
or U1850 (N_1850,N_1553,N_1575);
xnor U1851 (N_1851,N_1598,N_1718);
and U1852 (N_1852,N_1661,N_1707);
or U1853 (N_1853,N_1667,N_1557);
or U1854 (N_1854,N_1638,N_1576);
and U1855 (N_1855,N_1548,N_1689);
or U1856 (N_1856,N_1653,N_1649);
and U1857 (N_1857,N_1502,N_1719);
nor U1858 (N_1858,N_1688,N_1674);
nand U1859 (N_1859,N_1515,N_1727);
nand U1860 (N_1860,N_1594,N_1566);
or U1861 (N_1861,N_1582,N_1680);
or U1862 (N_1862,N_1585,N_1726);
xor U1863 (N_1863,N_1574,N_1586);
nand U1864 (N_1864,N_1572,N_1555);
nor U1865 (N_1865,N_1709,N_1650);
nor U1866 (N_1866,N_1546,N_1504);
or U1867 (N_1867,N_1747,N_1636);
or U1868 (N_1868,N_1666,N_1610);
and U1869 (N_1869,N_1506,N_1685);
xor U1870 (N_1870,N_1545,N_1509);
nor U1871 (N_1871,N_1710,N_1544);
xor U1872 (N_1872,N_1671,N_1748);
nor U1873 (N_1873,N_1542,N_1668);
nor U1874 (N_1874,N_1692,N_1743);
nand U1875 (N_1875,N_1601,N_1573);
nand U1876 (N_1876,N_1706,N_1635);
nor U1877 (N_1877,N_1694,N_1593);
nor U1878 (N_1878,N_1631,N_1655);
xnor U1879 (N_1879,N_1621,N_1562);
and U1880 (N_1880,N_1684,N_1727);
and U1881 (N_1881,N_1682,N_1523);
and U1882 (N_1882,N_1501,N_1749);
xnor U1883 (N_1883,N_1739,N_1633);
nand U1884 (N_1884,N_1511,N_1530);
and U1885 (N_1885,N_1727,N_1557);
and U1886 (N_1886,N_1687,N_1585);
or U1887 (N_1887,N_1734,N_1504);
nor U1888 (N_1888,N_1601,N_1619);
or U1889 (N_1889,N_1600,N_1601);
nor U1890 (N_1890,N_1544,N_1697);
xor U1891 (N_1891,N_1590,N_1580);
nand U1892 (N_1892,N_1669,N_1533);
or U1893 (N_1893,N_1738,N_1602);
nand U1894 (N_1894,N_1636,N_1572);
or U1895 (N_1895,N_1595,N_1591);
xnor U1896 (N_1896,N_1667,N_1551);
and U1897 (N_1897,N_1668,N_1523);
nor U1898 (N_1898,N_1645,N_1680);
and U1899 (N_1899,N_1731,N_1510);
nor U1900 (N_1900,N_1679,N_1582);
xor U1901 (N_1901,N_1722,N_1656);
and U1902 (N_1902,N_1650,N_1671);
or U1903 (N_1903,N_1569,N_1520);
nand U1904 (N_1904,N_1618,N_1662);
and U1905 (N_1905,N_1586,N_1696);
nor U1906 (N_1906,N_1740,N_1609);
nand U1907 (N_1907,N_1525,N_1521);
nand U1908 (N_1908,N_1552,N_1508);
nand U1909 (N_1909,N_1600,N_1705);
or U1910 (N_1910,N_1544,N_1581);
nor U1911 (N_1911,N_1694,N_1689);
xor U1912 (N_1912,N_1725,N_1640);
nor U1913 (N_1913,N_1541,N_1542);
nand U1914 (N_1914,N_1579,N_1643);
nand U1915 (N_1915,N_1743,N_1573);
or U1916 (N_1916,N_1665,N_1565);
nor U1917 (N_1917,N_1511,N_1540);
nand U1918 (N_1918,N_1746,N_1647);
or U1919 (N_1919,N_1697,N_1710);
nor U1920 (N_1920,N_1745,N_1731);
nor U1921 (N_1921,N_1616,N_1651);
and U1922 (N_1922,N_1682,N_1657);
or U1923 (N_1923,N_1624,N_1510);
nand U1924 (N_1924,N_1693,N_1653);
or U1925 (N_1925,N_1710,N_1720);
xnor U1926 (N_1926,N_1712,N_1717);
or U1927 (N_1927,N_1726,N_1533);
and U1928 (N_1928,N_1516,N_1539);
nand U1929 (N_1929,N_1591,N_1505);
nand U1930 (N_1930,N_1581,N_1583);
and U1931 (N_1931,N_1711,N_1621);
nand U1932 (N_1932,N_1587,N_1605);
nor U1933 (N_1933,N_1530,N_1716);
nand U1934 (N_1934,N_1741,N_1527);
nor U1935 (N_1935,N_1551,N_1549);
nor U1936 (N_1936,N_1693,N_1531);
and U1937 (N_1937,N_1512,N_1709);
nand U1938 (N_1938,N_1602,N_1512);
or U1939 (N_1939,N_1598,N_1733);
nor U1940 (N_1940,N_1702,N_1515);
nor U1941 (N_1941,N_1748,N_1717);
and U1942 (N_1942,N_1715,N_1723);
nand U1943 (N_1943,N_1663,N_1554);
and U1944 (N_1944,N_1662,N_1634);
nand U1945 (N_1945,N_1511,N_1670);
nand U1946 (N_1946,N_1536,N_1591);
or U1947 (N_1947,N_1672,N_1745);
xnor U1948 (N_1948,N_1552,N_1732);
xnor U1949 (N_1949,N_1738,N_1684);
or U1950 (N_1950,N_1640,N_1689);
and U1951 (N_1951,N_1699,N_1505);
nand U1952 (N_1952,N_1747,N_1704);
and U1953 (N_1953,N_1621,N_1666);
nor U1954 (N_1954,N_1693,N_1522);
or U1955 (N_1955,N_1560,N_1567);
nand U1956 (N_1956,N_1601,N_1520);
and U1957 (N_1957,N_1645,N_1613);
nand U1958 (N_1958,N_1508,N_1627);
nor U1959 (N_1959,N_1638,N_1508);
xnor U1960 (N_1960,N_1576,N_1525);
nand U1961 (N_1961,N_1569,N_1551);
and U1962 (N_1962,N_1734,N_1747);
nand U1963 (N_1963,N_1612,N_1520);
xor U1964 (N_1964,N_1561,N_1705);
nor U1965 (N_1965,N_1534,N_1748);
and U1966 (N_1966,N_1660,N_1553);
xnor U1967 (N_1967,N_1672,N_1676);
nand U1968 (N_1968,N_1708,N_1717);
nand U1969 (N_1969,N_1735,N_1618);
and U1970 (N_1970,N_1544,N_1631);
nand U1971 (N_1971,N_1549,N_1668);
nor U1972 (N_1972,N_1590,N_1698);
nand U1973 (N_1973,N_1675,N_1608);
nand U1974 (N_1974,N_1643,N_1666);
nand U1975 (N_1975,N_1583,N_1645);
nand U1976 (N_1976,N_1549,N_1591);
and U1977 (N_1977,N_1503,N_1696);
xor U1978 (N_1978,N_1661,N_1552);
xnor U1979 (N_1979,N_1749,N_1643);
and U1980 (N_1980,N_1510,N_1613);
and U1981 (N_1981,N_1507,N_1740);
nor U1982 (N_1982,N_1620,N_1617);
or U1983 (N_1983,N_1706,N_1639);
and U1984 (N_1984,N_1581,N_1520);
xnor U1985 (N_1985,N_1662,N_1502);
and U1986 (N_1986,N_1681,N_1657);
nor U1987 (N_1987,N_1608,N_1749);
and U1988 (N_1988,N_1714,N_1665);
nand U1989 (N_1989,N_1512,N_1544);
or U1990 (N_1990,N_1585,N_1636);
xnor U1991 (N_1991,N_1648,N_1539);
xnor U1992 (N_1992,N_1696,N_1591);
xnor U1993 (N_1993,N_1584,N_1607);
xor U1994 (N_1994,N_1668,N_1670);
xor U1995 (N_1995,N_1654,N_1581);
xnor U1996 (N_1996,N_1667,N_1546);
nand U1997 (N_1997,N_1717,N_1719);
nand U1998 (N_1998,N_1636,N_1732);
nand U1999 (N_1999,N_1617,N_1699);
nor U2000 (N_2000,N_1827,N_1791);
or U2001 (N_2001,N_1913,N_1815);
nor U2002 (N_2002,N_1822,N_1916);
nand U2003 (N_2003,N_1989,N_1774);
or U2004 (N_2004,N_1996,N_1817);
xnor U2005 (N_2005,N_1927,N_1896);
nand U2006 (N_2006,N_1825,N_1810);
nor U2007 (N_2007,N_1767,N_1849);
nor U2008 (N_2008,N_1887,N_1765);
and U2009 (N_2009,N_1976,N_1975);
and U2010 (N_2010,N_1970,N_1836);
xnor U2011 (N_2011,N_1958,N_1813);
and U2012 (N_2012,N_1771,N_1961);
nand U2013 (N_2013,N_1912,N_1966);
nand U2014 (N_2014,N_1934,N_1768);
nand U2015 (N_2015,N_1929,N_1756);
and U2016 (N_2016,N_1925,N_1939);
nor U2017 (N_2017,N_1763,N_1856);
nor U2018 (N_2018,N_1816,N_1840);
and U2019 (N_2019,N_1980,N_1891);
and U2020 (N_2020,N_1898,N_1955);
nor U2021 (N_2021,N_1972,N_1858);
xor U2022 (N_2022,N_1871,N_1773);
nor U2023 (N_2023,N_1909,N_1953);
nand U2024 (N_2024,N_1950,N_1936);
or U2025 (N_2025,N_1819,N_1963);
and U2026 (N_2026,N_1753,N_1841);
or U2027 (N_2027,N_1990,N_1757);
xnor U2028 (N_2028,N_1986,N_1988);
xnor U2029 (N_2029,N_1780,N_1910);
nand U2030 (N_2030,N_1801,N_1894);
and U2031 (N_2031,N_1949,N_1831);
nor U2032 (N_2032,N_1957,N_1799);
xor U2033 (N_2033,N_1755,N_1775);
nand U2034 (N_2034,N_1984,N_1888);
xnor U2035 (N_2035,N_1754,N_1759);
and U2036 (N_2036,N_1863,N_1921);
and U2037 (N_2037,N_1850,N_1964);
or U2038 (N_2038,N_1787,N_1952);
and U2039 (N_2039,N_1944,N_1785);
or U2040 (N_2040,N_1954,N_1778);
and U2041 (N_2041,N_1854,N_1938);
nor U2042 (N_2042,N_1766,N_1917);
nand U2043 (N_2043,N_1832,N_1835);
or U2044 (N_2044,N_1807,N_1999);
xnor U2045 (N_2045,N_1873,N_1793);
nor U2046 (N_2046,N_1907,N_1920);
nor U2047 (N_2047,N_1890,N_1930);
and U2048 (N_2048,N_1770,N_1993);
nor U2049 (N_2049,N_1956,N_1919);
or U2050 (N_2050,N_1977,N_1895);
and U2051 (N_2051,N_1971,N_1779);
nor U2052 (N_2052,N_1940,N_1908);
or U2053 (N_2053,N_1901,N_1973);
or U2054 (N_2054,N_1969,N_1951);
nand U2055 (N_2055,N_1985,N_1877);
nand U2056 (N_2056,N_1783,N_1782);
or U2057 (N_2057,N_1933,N_1842);
xor U2058 (N_2058,N_1884,N_1794);
nor U2059 (N_2059,N_1857,N_1855);
nand U2060 (N_2060,N_1860,N_1862);
nor U2061 (N_2061,N_1983,N_1981);
and U2062 (N_2062,N_1946,N_1828);
or U2063 (N_2063,N_1797,N_1991);
xor U2064 (N_2064,N_1760,N_1848);
nand U2065 (N_2065,N_1897,N_1900);
and U2066 (N_2066,N_1881,N_1859);
nor U2067 (N_2067,N_1750,N_1875);
nand U2068 (N_2068,N_1876,N_1914);
xnor U2069 (N_2069,N_1866,N_1812);
xnor U2070 (N_2070,N_1853,N_1947);
nand U2071 (N_2071,N_1776,N_1792);
nand U2072 (N_2072,N_1962,N_1931);
nor U2073 (N_2073,N_1883,N_1905);
and U2074 (N_2074,N_1761,N_1837);
xor U2075 (N_2075,N_1926,N_1823);
nor U2076 (N_2076,N_1786,N_1790);
xnor U2077 (N_2077,N_1826,N_1903);
or U2078 (N_2078,N_1994,N_1843);
or U2079 (N_2079,N_1751,N_1824);
or U2080 (N_2080,N_1752,N_1924);
xnor U2081 (N_2081,N_1979,N_1874);
xnor U2082 (N_2082,N_1915,N_1800);
and U2083 (N_2083,N_1846,N_1861);
or U2084 (N_2084,N_1889,N_1829);
and U2085 (N_2085,N_1870,N_1784);
nor U2086 (N_2086,N_1802,N_1821);
xnor U2087 (N_2087,N_1762,N_1818);
nor U2088 (N_2088,N_1788,N_1844);
nand U2089 (N_2089,N_1852,N_1808);
nand U2090 (N_2090,N_1880,N_1804);
and U2091 (N_2091,N_1867,N_1959);
nor U2092 (N_2092,N_1928,N_1911);
and U2093 (N_2093,N_1772,N_1878);
xor U2094 (N_2094,N_1918,N_1864);
xnor U2095 (N_2095,N_1798,N_1965);
and U2096 (N_2096,N_1789,N_1838);
nand U2097 (N_2097,N_1968,N_1932);
xor U2098 (N_2098,N_1906,N_1892);
nor U2099 (N_2099,N_1882,N_1997);
nor U2100 (N_2100,N_1904,N_1941);
nor U2101 (N_2101,N_1899,N_1995);
or U2102 (N_2102,N_1839,N_1811);
nor U2103 (N_2103,N_1777,N_1982);
and U2104 (N_2104,N_1945,N_1758);
nand U2105 (N_2105,N_1902,N_1974);
nor U2106 (N_2106,N_1796,N_1764);
and U2107 (N_2107,N_1872,N_1893);
xor U2108 (N_2108,N_1820,N_1869);
nor U2109 (N_2109,N_1942,N_1809);
nor U2110 (N_2110,N_1803,N_1943);
nor U2111 (N_2111,N_1781,N_1885);
xnor U2112 (N_2112,N_1805,N_1967);
xor U2113 (N_2113,N_1845,N_1806);
and U2114 (N_2114,N_1935,N_1960);
or U2115 (N_2115,N_1834,N_1923);
or U2116 (N_2116,N_1922,N_1847);
nand U2117 (N_2117,N_1833,N_1830);
xor U2118 (N_2118,N_1937,N_1992);
and U2119 (N_2119,N_1865,N_1948);
xnor U2120 (N_2120,N_1987,N_1879);
and U2121 (N_2121,N_1769,N_1814);
or U2122 (N_2122,N_1886,N_1978);
nor U2123 (N_2123,N_1868,N_1795);
xnor U2124 (N_2124,N_1851,N_1998);
or U2125 (N_2125,N_1862,N_1813);
and U2126 (N_2126,N_1823,N_1940);
and U2127 (N_2127,N_1991,N_1782);
xnor U2128 (N_2128,N_1767,N_1961);
xnor U2129 (N_2129,N_1871,N_1976);
nor U2130 (N_2130,N_1990,N_1790);
nand U2131 (N_2131,N_1849,N_1922);
xor U2132 (N_2132,N_1980,N_1991);
xor U2133 (N_2133,N_1912,N_1833);
or U2134 (N_2134,N_1879,N_1936);
and U2135 (N_2135,N_1871,N_1958);
or U2136 (N_2136,N_1841,N_1939);
or U2137 (N_2137,N_1849,N_1937);
and U2138 (N_2138,N_1942,N_1930);
and U2139 (N_2139,N_1753,N_1997);
or U2140 (N_2140,N_1811,N_1796);
and U2141 (N_2141,N_1981,N_1878);
xnor U2142 (N_2142,N_1814,N_1964);
xor U2143 (N_2143,N_1763,N_1776);
nor U2144 (N_2144,N_1951,N_1806);
nand U2145 (N_2145,N_1989,N_1937);
nor U2146 (N_2146,N_1797,N_1769);
and U2147 (N_2147,N_1850,N_1767);
nor U2148 (N_2148,N_1982,N_1793);
nand U2149 (N_2149,N_1847,N_1952);
or U2150 (N_2150,N_1792,N_1837);
nor U2151 (N_2151,N_1753,N_1852);
xnor U2152 (N_2152,N_1957,N_1870);
nor U2153 (N_2153,N_1905,N_1940);
nor U2154 (N_2154,N_1781,N_1911);
nor U2155 (N_2155,N_1992,N_1885);
nor U2156 (N_2156,N_1795,N_1843);
and U2157 (N_2157,N_1974,N_1827);
nand U2158 (N_2158,N_1923,N_1936);
nor U2159 (N_2159,N_1892,N_1825);
xor U2160 (N_2160,N_1831,N_1955);
and U2161 (N_2161,N_1805,N_1941);
nor U2162 (N_2162,N_1859,N_1910);
or U2163 (N_2163,N_1921,N_1754);
nor U2164 (N_2164,N_1789,N_1776);
and U2165 (N_2165,N_1976,N_1918);
and U2166 (N_2166,N_1962,N_1780);
and U2167 (N_2167,N_1911,N_1962);
or U2168 (N_2168,N_1815,N_1908);
nand U2169 (N_2169,N_1867,N_1967);
or U2170 (N_2170,N_1883,N_1966);
or U2171 (N_2171,N_1931,N_1880);
nor U2172 (N_2172,N_1834,N_1801);
or U2173 (N_2173,N_1828,N_1914);
nor U2174 (N_2174,N_1980,N_1957);
and U2175 (N_2175,N_1975,N_1763);
xor U2176 (N_2176,N_1960,N_1824);
nand U2177 (N_2177,N_1972,N_1864);
and U2178 (N_2178,N_1868,N_1809);
nand U2179 (N_2179,N_1866,N_1939);
nand U2180 (N_2180,N_1930,N_1800);
or U2181 (N_2181,N_1940,N_1821);
xnor U2182 (N_2182,N_1814,N_1934);
and U2183 (N_2183,N_1890,N_1840);
xnor U2184 (N_2184,N_1998,N_1916);
or U2185 (N_2185,N_1940,N_1827);
nand U2186 (N_2186,N_1925,N_1810);
xor U2187 (N_2187,N_1869,N_1762);
and U2188 (N_2188,N_1751,N_1977);
or U2189 (N_2189,N_1843,N_1881);
and U2190 (N_2190,N_1816,N_1819);
xnor U2191 (N_2191,N_1879,N_1909);
or U2192 (N_2192,N_1835,N_1912);
xnor U2193 (N_2193,N_1934,N_1848);
or U2194 (N_2194,N_1790,N_1785);
nor U2195 (N_2195,N_1873,N_1870);
nand U2196 (N_2196,N_1898,N_1999);
xnor U2197 (N_2197,N_1819,N_1836);
or U2198 (N_2198,N_1921,N_1776);
or U2199 (N_2199,N_1958,N_1812);
or U2200 (N_2200,N_1880,N_1750);
nand U2201 (N_2201,N_1815,N_1817);
xor U2202 (N_2202,N_1787,N_1988);
or U2203 (N_2203,N_1868,N_1857);
xor U2204 (N_2204,N_1974,N_1900);
and U2205 (N_2205,N_1871,N_1829);
and U2206 (N_2206,N_1991,N_1950);
or U2207 (N_2207,N_1983,N_1860);
xor U2208 (N_2208,N_1939,N_1968);
or U2209 (N_2209,N_1819,N_1944);
xnor U2210 (N_2210,N_1907,N_1750);
or U2211 (N_2211,N_1798,N_1865);
and U2212 (N_2212,N_1940,N_1782);
xnor U2213 (N_2213,N_1840,N_1977);
xnor U2214 (N_2214,N_1871,N_1858);
nor U2215 (N_2215,N_1978,N_1806);
nor U2216 (N_2216,N_1973,N_1761);
nand U2217 (N_2217,N_1946,N_1772);
or U2218 (N_2218,N_1811,N_1913);
or U2219 (N_2219,N_1796,N_1965);
and U2220 (N_2220,N_1796,N_1859);
and U2221 (N_2221,N_1907,N_1803);
xnor U2222 (N_2222,N_1809,N_1827);
or U2223 (N_2223,N_1928,N_1962);
xor U2224 (N_2224,N_1908,N_1823);
or U2225 (N_2225,N_1911,N_1775);
nand U2226 (N_2226,N_1882,N_1817);
nand U2227 (N_2227,N_1776,N_1959);
or U2228 (N_2228,N_1864,N_1772);
nor U2229 (N_2229,N_1933,N_1896);
nand U2230 (N_2230,N_1965,N_1869);
nor U2231 (N_2231,N_1854,N_1798);
nand U2232 (N_2232,N_1783,N_1899);
nor U2233 (N_2233,N_1868,N_1752);
or U2234 (N_2234,N_1785,N_1968);
and U2235 (N_2235,N_1791,N_1837);
and U2236 (N_2236,N_1838,N_1957);
or U2237 (N_2237,N_1870,N_1924);
nand U2238 (N_2238,N_1781,N_1832);
or U2239 (N_2239,N_1905,N_1800);
nand U2240 (N_2240,N_1950,N_1967);
or U2241 (N_2241,N_1829,N_1771);
and U2242 (N_2242,N_1764,N_1979);
or U2243 (N_2243,N_1766,N_1774);
and U2244 (N_2244,N_1969,N_1949);
nand U2245 (N_2245,N_1837,N_1957);
nor U2246 (N_2246,N_1869,N_1801);
nor U2247 (N_2247,N_1780,N_1842);
or U2248 (N_2248,N_1791,N_1868);
xor U2249 (N_2249,N_1954,N_1761);
or U2250 (N_2250,N_2213,N_2193);
nand U2251 (N_2251,N_2017,N_2086);
nand U2252 (N_2252,N_2032,N_2013);
xnor U2253 (N_2253,N_2215,N_2173);
or U2254 (N_2254,N_2004,N_2188);
xor U2255 (N_2255,N_2183,N_2127);
nor U2256 (N_2256,N_2245,N_2071);
xor U2257 (N_2257,N_2058,N_2169);
nand U2258 (N_2258,N_2145,N_2014);
xor U2259 (N_2259,N_2234,N_2063);
or U2260 (N_2260,N_2199,N_2196);
xnor U2261 (N_2261,N_2111,N_2008);
nand U2262 (N_2262,N_2003,N_2054);
xnor U2263 (N_2263,N_2040,N_2109);
or U2264 (N_2264,N_2077,N_2221);
or U2265 (N_2265,N_2016,N_2030);
and U2266 (N_2266,N_2052,N_2099);
nand U2267 (N_2267,N_2050,N_2080);
xor U2268 (N_2268,N_2085,N_2118);
xor U2269 (N_2269,N_2102,N_2084);
or U2270 (N_2270,N_2176,N_2222);
nor U2271 (N_2271,N_2185,N_2232);
nor U2272 (N_2272,N_2225,N_2048);
nand U2273 (N_2273,N_2178,N_2010);
or U2274 (N_2274,N_2108,N_2066);
and U2275 (N_2275,N_2165,N_2024);
nand U2276 (N_2276,N_2007,N_2171);
nor U2277 (N_2277,N_2142,N_2131);
or U2278 (N_2278,N_2037,N_2206);
xor U2279 (N_2279,N_2116,N_2212);
nor U2280 (N_2280,N_2235,N_2081);
or U2281 (N_2281,N_2088,N_2233);
nor U2282 (N_2282,N_2208,N_2012);
xnor U2283 (N_2283,N_2097,N_2187);
or U2284 (N_2284,N_2031,N_2190);
nand U2285 (N_2285,N_2049,N_2149);
nor U2286 (N_2286,N_2143,N_2238);
xnor U2287 (N_2287,N_2237,N_2189);
nor U2288 (N_2288,N_2240,N_2159);
xnor U2289 (N_2289,N_2027,N_2115);
and U2290 (N_2290,N_2186,N_2090);
nor U2291 (N_2291,N_2074,N_2140);
xnor U2292 (N_2292,N_2098,N_2020);
or U2293 (N_2293,N_2141,N_2174);
and U2294 (N_2294,N_2104,N_2046);
nor U2295 (N_2295,N_2126,N_2192);
and U2296 (N_2296,N_2194,N_2076);
and U2297 (N_2297,N_2089,N_2248);
nor U2298 (N_2298,N_2091,N_2092);
or U2299 (N_2299,N_2055,N_2095);
or U2300 (N_2300,N_2082,N_2203);
or U2301 (N_2301,N_2035,N_2179);
or U2302 (N_2302,N_2180,N_2167);
or U2303 (N_2303,N_2177,N_2200);
or U2304 (N_2304,N_2152,N_2172);
nor U2305 (N_2305,N_2241,N_2110);
nand U2306 (N_2306,N_2220,N_2019);
nor U2307 (N_2307,N_2057,N_2157);
nand U2308 (N_2308,N_2138,N_2181);
or U2309 (N_2309,N_2029,N_2106);
xor U2310 (N_2310,N_2224,N_2064);
and U2311 (N_2311,N_2103,N_2112);
xnor U2312 (N_2312,N_2202,N_2056);
nor U2313 (N_2313,N_2168,N_2136);
nand U2314 (N_2314,N_2158,N_2053);
nor U2315 (N_2315,N_2228,N_2144);
and U2316 (N_2316,N_2244,N_2025);
nor U2317 (N_2317,N_2107,N_2028);
xnor U2318 (N_2318,N_2207,N_2105);
or U2319 (N_2319,N_2018,N_2022);
nor U2320 (N_2320,N_2044,N_2073);
nor U2321 (N_2321,N_2125,N_2042);
and U2322 (N_2322,N_2039,N_2114);
nor U2323 (N_2323,N_2191,N_2072);
nand U2324 (N_2324,N_2061,N_2083);
nor U2325 (N_2325,N_2006,N_2100);
nand U2326 (N_2326,N_2160,N_2209);
xor U2327 (N_2327,N_2214,N_2021);
nor U2328 (N_2328,N_2227,N_2062);
or U2329 (N_2329,N_2230,N_2069);
nand U2330 (N_2330,N_2005,N_2067);
xnor U2331 (N_2331,N_2117,N_2123);
nand U2332 (N_2332,N_2217,N_2120);
or U2333 (N_2333,N_2231,N_2101);
nand U2334 (N_2334,N_2151,N_2009);
xor U2335 (N_2335,N_2205,N_2043);
nand U2336 (N_2336,N_2243,N_2201);
and U2337 (N_2337,N_2000,N_2175);
or U2338 (N_2338,N_2223,N_2122);
xnor U2339 (N_2339,N_2078,N_2033);
xor U2340 (N_2340,N_2094,N_2164);
and U2341 (N_2341,N_2249,N_2239);
and U2342 (N_2342,N_2060,N_2041);
xnor U2343 (N_2343,N_2129,N_2211);
xnor U2344 (N_2344,N_2045,N_2229);
and U2345 (N_2345,N_2236,N_2075);
nand U2346 (N_2346,N_2148,N_2163);
xnor U2347 (N_2347,N_2197,N_2093);
nand U2348 (N_2348,N_2023,N_2135);
nand U2349 (N_2349,N_2219,N_2134);
xor U2350 (N_2350,N_2153,N_2065);
nand U2351 (N_2351,N_2034,N_2026);
nor U2352 (N_2352,N_2195,N_2146);
nor U2353 (N_2353,N_2170,N_2130);
nand U2354 (N_2354,N_2204,N_2161);
xor U2355 (N_2355,N_2133,N_2139);
xor U2356 (N_2356,N_2121,N_2036);
or U2357 (N_2357,N_2059,N_2155);
xnor U2358 (N_2358,N_2015,N_2068);
nor U2359 (N_2359,N_2070,N_2242);
xor U2360 (N_2360,N_2124,N_2184);
xnor U2361 (N_2361,N_2156,N_2216);
and U2362 (N_2362,N_2011,N_2002);
xnor U2363 (N_2363,N_2132,N_2087);
nand U2364 (N_2364,N_2128,N_2147);
and U2365 (N_2365,N_2038,N_2051);
nor U2366 (N_2366,N_2154,N_2079);
nor U2367 (N_2367,N_2113,N_2166);
or U2368 (N_2368,N_2226,N_2047);
or U2369 (N_2369,N_2198,N_2210);
and U2370 (N_2370,N_2119,N_2137);
nand U2371 (N_2371,N_2218,N_2162);
nor U2372 (N_2372,N_2246,N_2001);
xor U2373 (N_2373,N_2247,N_2096);
nand U2374 (N_2374,N_2182,N_2150);
or U2375 (N_2375,N_2045,N_2007);
or U2376 (N_2376,N_2100,N_2088);
or U2377 (N_2377,N_2230,N_2018);
nand U2378 (N_2378,N_2149,N_2025);
xor U2379 (N_2379,N_2092,N_2243);
xnor U2380 (N_2380,N_2166,N_2025);
nand U2381 (N_2381,N_2203,N_2148);
nand U2382 (N_2382,N_2172,N_2030);
and U2383 (N_2383,N_2113,N_2073);
xor U2384 (N_2384,N_2062,N_2244);
xor U2385 (N_2385,N_2016,N_2090);
xnor U2386 (N_2386,N_2109,N_2146);
nor U2387 (N_2387,N_2034,N_2044);
xor U2388 (N_2388,N_2172,N_2135);
nor U2389 (N_2389,N_2196,N_2166);
nor U2390 (N_2390,N_2085,N_2184);
nor U2391 (N_2391,N_2126,N_2004);
and U2392 (N_2392,N_2194,N_2025);
nor U2393 (N_2393,N_2158,N_2177);
and U2394 (N_2394,N_2030,N_2216);
or U2395 (N_2395,N_2187,N_2164);
nand U2396 (N_2396,N_2055,N_2023);
xnor U2397 (N_2397,N_2081,N_2191);
nor U2398 (N_2398,N_2075,N_2231);
nand U2399 (N_2399,N_2129,N_2141);
nor U2400 (N_2400,N_2189,N_2051);
or U2401 (N_2401,N_2193,N_2167);
nor U2402 (N_2402,N_2026,N_2070);
nor U2403 (N_2403,N_2010,N_2173);
nor U2404 (N_2404,N_2043,N_2052);
xor U2405 (N_2405,N_2159,N_2069);
or U2406 (N_2406,N_2096,N_2215);
xor U2407 (N_2407,N_2011,N_2023);
nand U2408 (N_2408,N_2215,N_2221);
nor U2409 (N_2409,N_2212,N_2030);
xnor U2410 (N_2410,N_2157,N_2231);
nand U2411 (N_2411,N_2079,N_2076);
and U2412 (N_2412,N_2038,N_2108);
or U2413 (N_2413,N_2201,N_2027);
nor U2414 (N_2414,N_2153,N_2005);
nor U2415 (N_2415,N_2082,N_2221);
and U2416 (N_2416,N_2017,N_2192);
or U2417 (N_2417,N_2207,N_2128);
nand U2418 (N_2418,N_2075,N_2191);
or U2419 (N_2419,N_2210,N_2054);
nand U2420 (N_2420,N_2188,N_2097);
or U2421 (N_2421,N_2054,N_2238);
and U2422 (N_2422,N_2144,N_2146);
and U2423 (N_2423,N_2001,N_2027);
nand U2424 (N_2424,N_2110,N_2142);
nand U2425 (N_2425,N_2146,N_2103);
nand U2426 (N_2426,N_2148,N_2041);
or U2427 (N_2427,N_2129,N_2243);
or U2428 (N_2428,N_2229,N_2031);
xor U2429 (N_2429,N_2046,N_2123);
or U2430 (N_2430,N_2180,N_2165);
xnor U2431 (N_2431,N_2188,N_2169);
xor U2432 (N_2432,N_2156,N_2025);
xor U2433 (N_2433,N_2232,N_2039);
xnor U2434 (N_2434,N_2173,N_2177);
nor U2435 (N_2435,N_2120,N_2069);
xor U2436 (N_2436,N_2012,N_2167);
nor U2437 (N_2437,N_2092,N_2134);
nor U2438 (N_2438,N_2112,N_2164);
nand U2439 (N_2439,N_2227,N_2242);
nor U2440 (N_2440,N_2037,N_2066);
and U2441 (N_2441,N_2246,N_2062);
or U2442 (N_2442,N_2117,N_2172);
xnor U2443 (N_2443,N_2084,N_2233);
or U2444 (N_2444,N_2164,N_2024);
or U2445 (N_2445,N_2144,N_2104);
nand U2446 (N_2446,N_2012,N_2019);
or U2447 (N_2447,N_2101,N_2123);
xnor U2448 (N_2448,N_2085,N_2092);
and U2449 (N_2449,N_2154,N_2238);
nand U2450 (N_2450,N_2192,N_2019);
or U2451 (N_2451,N_2032,N_2166);
or U2452 (N_2452,N_2214,N_2058);
nor U2453 (N_2453,N_2017,N_2069);
nand U2454 (N_2454,N_2218,N_2116);
nand U2455 (N_2455,N_2128,N_2227);
nor U2456 (N_2456,N_2244,N_2052);
nand U2457 (N_2457,N_2196,N_2215);
or U2458 (N_2458,N_2204,N_2137);
nand U2459 (N_2459,N_2024,N_2213);
and U2460 (N_2460,N_2052,N_2073);
nand U2461 (N_2461,N_2197,N_2075);
nand U2462 (N_2462,N_2246,N_2078);
or U2463 (N_2463,N_2011,N_2199);
or U2464 (N_2464,N_2129,N_2165);
nand U2465 (N_2465,N_2021,N_2061);
xnor U2466 (N_2466,N_2052,N_2179);
nor U2467 (N_2467,N_2171,N_2191);
xnor U2468 (N_2468,N_2036,N_2188);
nor U2469 (N_2469,N_2239,N_2141);
or U2470 (N_2470,N_2194,N_2004);
nand U2471 (N_2471,N_2117,N_2069);
xnor U2472 (N_2472,N_2083,N_2244);
and U2473 (N_2473,N_2180,N_2128);
nand U2474 (N_2474,N_2171,N_2066);
xnor U2475 (N_2475,N_2183,N_2154);
nand U2476 (N_2476,N_2185,N_2014);
or U2477 (N_2477,N_2080,N_2091);
xnor U2478 (N_2478,N_2018,N_2005);
and U2479 (N_2479,N_2043,N_2102);
or U2480 (N_2480,N_2107,N_2002);
or U2481 (N_2481,N_2217,N_2023);
nor U2482 (N_2482,N_2121,N_2037);
xnor U2483 (N_2483,N_2090,N_2012);
nand U2484 (N_2484,N_2171,N_2220);
and U2485 (N_2485,N_2118,N_2177);
or U2486 (N_2486,N_2038,N_2086);
xor U2487 (N_2487,N_2085,N_2035);
nand U2488 (N_2488,N_2226,N_2098);
and U2489 (N_2489,N_2063,N_2101);
or U2490 (N_2490,N_2134,N_2121);
nor U2491 (N_2491,N_2167,N_2201);
xnor U2492 (N_2492,N_2171,N_2241);
nand U2493 (N_2493,N_2121,N_2141);
nand U2494 (N_2494,N_2186,N_2005);
xor U2495 (N_2495,N_2194,N_2177);
xnor U2496 (N_2496,N_2051,N_2112);
nor U2497 (N_2497,N_2237,N_2108);
and U2498 (N_2498,N_2248,N_2034);
or U2499 (N_2499,N_2155,N_2055);
xor U2500 (N_2500,N_2261,N_2416);
nand U2501 (N_2501,N_2279,N_2420);
xnor U2502 (N_2502,N_2302,N_2490);
nand U2503 (N_2503,N_2267,N_2411);
xnor U2504 (N_2504,N_2404,N_2410);
xnor U2505 (N_2505,N_2364,N_2314);
xor U2506 (N_2506,N_2263,N_2491);
xnor U2507 (N_2507,N_2257,N_2297);
nand U2508 (N_2508,N_2296,N_2481);
and U2509 (N_2509,N_2375,N_2403);
and U2510 (N_2510,N_2483,N_2399);
nand U2511 (N_2511,N_2444,N_2389);
or U2512 (N_2512,N_2370,N_2357);
nand U2513 (N_2513,N_2306,N_2354);
nand U2514 (N_2514,N_2327,N_2480);
xnor U2515 (N_2515,N_2400,N_2280);
nor U2516 (N_2516,N_2360,N_2269);
and U2517 (N_2517,N_2395,N_2468);
or U2518 (N_2518,N_2352,N_2313);
xnor U2519 (N_2519,N_2310,N_2259);
nand U2520 (N_2520,N_2309,N_2287);
or U2521 (N_2521,N_2377,N_2252);
nor U2522 (N_2522,N_2396,N_2356);
and U2523 (N_2523,N_2251,N_2338);
or U2524 (N_2524,N_2429,N_2434);
nand U2525 (N_2525,N_2373,N_2469);
xnor U2526 (N_2526,N_2451,N_2368);
nand U2527 (N_2527,N_2311,N_2367);
nor U2528 (N_2528,N_2378,N_2401);
nand U2529 (N_2529,N_2449,N_2332);
and U2530 (N_2530,N_2328,N_2488);
or U2531 (N_2531,N_2433,N_2336);
nor U2532 (N_2532,N_2255,N_2426);
or U2533 (N_2533,N_2308,N_2331);
nor U2534 (N_2534,N_2325,N_2326);
and U2535 (N_2535,N_2260,N_2254);
or U2536 (N_2536,N_2372,N_2461);
and U2537 (N_2537,N_2348,N_2288);
xor U2538 (N_2538,N_2462,N_2382);
nand U2539 (N_2539,N_2365,N_2475);
xnor U2540 (N_2540,N_2463,N_2290);
and U2541 (N_2541,N_2446,N_2284);
nor U2542 (N_2542,N_2489,N_2472);
or U2543 (N_2543,N_2487,N_2307);
xnor U2544 (N_2544,N_2262,N_2477);
or U2545 (N_2545,N_2391,N_2409);
and U2546 (N_2546,N_2376,N_2436);
or U2547 (N_2547,N_2272,N_2438);
nand U2548 (N_2548,N_2454,N_2393);
and U2549 (N_2549,N_2405,N_2441);
nand U2550 (N_2550,N_2268,N_2492);
or U2551 (N_2551,N_2442,N_2467);
nand U2552 (N_2552,N_2484,N_2270);
xnor U2553 (N_2553,N_2478,N_2371);
nand U2554 (N_2554,N_2406,N_2387);
or U2555 (N_2555,N_2397,N_2407);
or U2556 (N_2556,N_2322,N_2320);
nand U2557 (N_2557,N_2455,N_2292);
nor U2558 (N_2558,N_2448,N_2277);
xnor U2559 (N_2559,N_2447,N_2473);
nand U2560 (N_2560,N_2341,N_2271);
nand U2561 (N_2561,N_2428,N_2415);
and U2562 (N_2562,N_2374,N_2324);
or U2563 (N_2563,N_2298,N_2273);
xnor U2564 (N_2564,N_2497,N_2423);
nor U2565 (N_2565,N_2380,N_2349);
nor U2566 (N_2566,N_2392,N_2351);
and U2567 (N_2567,N_2440,N_2318);
nor U2568 (N_2568,N_2281,N_2353);
nand U2569 (N_2569,N_2276,N_2286);
nor U2570 (N_2570,N_2304,N_2312);
nand U2571 (N_2571,N_2482,N_2432);
nor U2572 (N_2572,N_2294,N_2285);
nand U2573 (N_2573,N_2499,N_2430);
nand U2574 (N_2574,N_2340,N_2435);
xnor U2575 (N_2575,N_2299,N_2274);
nand U2576 (N_2576,N_2474,N_2346);
xnor U2577 (N_2577,N_2443,N_2253);
and U2578 (N_2578,N_2402,N_2398);
xnor U2579 (N_2579,N_2265,N_2300);
nor U2580 (N_2580,N_2342,N_2383);
and U2581 (N_2581,N_2350,N_2323);
or U2582 (N_2582,N_2419,N_2388);
nand U2583 (N_2583,N_2344,N_2355);
and U2584 (N_2584,N_2431,N_2337);
nor U2585 (N_2585,N_2498,N_2394);
nand U2586 (N_2586,N_2439,N_2339);
or U2587 (N_2587,N_2414,N_2418);
or U2588 (N_2588,N_2495,N_2465);
nor U2589 (N_2589,N_2457,N_2330);
nor U2590 (N_2590,N_2494,N_2421);
or U2591 (N_2591,N_2264,N_2450);
nand U2592 (N_2592,N_2424,N_2321);
or U2593 (N_2593,N_2466,N_2379);
or U2594 (N_2594,N_2305,N_2496);
xor U2595 (N_2595,N_2453,N_2427);
nor U2596 (N_2596,N_2460,N_2452);
nand U2597 (N_2597,N_2283,N_2479);
nor U2598 (N_2598,N_2458,N_2413);
nor U2599 (N_2599,N_2295,N_2359);
nand U2600 (N_2600,N_2390,N_2329);
or U2601 (N_2601,N_2381,N_2417);
nor U2602 (N_2602,N_2319,N_2258);
xnor U2603 (N_2603,N_2470,N_2408);
or U2604 (N_2604,N_2486,N_2485);
xnor U2605 (N_2605,N_2291,N_2343);
or U2606 (N_2606,N_2471,N_2422);
and U2607 (N_2607,N_2437,N_2385);
nor U2608 (N_2608,N_2476,N_2366);
nor U2609 (N_2609,N_2456,N_2369);
xnor U2610 (N_2610,N_2256,N_2289);
xnor U2611 (N_2611,N_2250,N_2266);
or U2612 (N_2612,N_2459,N_2384);
and U2613 (N_2613,N_2363,N_2445);
or U2614 (N_2614,N_2301,N_2386);
nand U2615 (N_2615,N_2278,N_2345);
xor U2616 (N_2616,N_2361,N_2333);
nor U2617 (N_2617,N_2275,N_2362);
xor U2618 (N_2618,N_2334,N_2317);
and U2619 (N_2619,N_2282,N_2493);
and U2620 (N_2620,N_2293,N_2347);
nor U2621 (N_2621,N_2425,N_2335);
nor U2622 (N_2622,N_2316,N_2315);
nand U2623 (N_2623,N_2464,N_2303);
and U2624 (N_2624,N_2358,N_2412);
nand U2625 (N_2625,N_2283,N_2366);
nand U2626 (N_2626,N_2457,N_2496);
and U2627 (N_2627,N_2297,N_2362);
and U2628 (N_2628,N_2469,N_2398);
or U2629 (N_2629,N_2258,N_2467);
nor U2630 (N_2630,N_2258,N_2417);
xor U2631 (N_2631,N_2388,N_2315);
and U2632 (N_2632,N_2467,N_2382);
xnor U2633 (N_2633,N_2445,N_2324);
or U2634 (N_2634,N_2259,N_2343);
and U2635 (N_2635,N_2493,N_2477);
xor U2636 (N_2636,N_2382,N_2442);
and U2637 (N_2637,N_2465,N_2402);
xor U2638 (N_2638,N_2393,N_2280);
nand U2639 (N_2639,N_2293,N_2426);
xnor U2640 (N_2640,N_2306,N_2468);
nand U2641 (N_2641,N_2428,N_2281);
nor U2642 (N_2642,N_2451,N_2333);
xnor U2643 (N_2643,N_2254,N_2493);
and U2644 (N_2644,N_2423,N_2483);
nand U2645 (N_2645,N_2288,N_2492);
nor U2646 (N_2646,N_2315,N_2474);
nor U2647 (N_2647,N_2371,N_2489);
nand U2648 (N_2648,N_2474,N_2295);
nor U2649 (N_2649,N_2388,N_2375);
and U2650 (N_2650,N_2264,N_2476);
nand U2651 (N_2651,N_2359,N_2258);
nand U2652 (N_2652,N_2295,N_2338);
xnor U2653 (N_2653,N_2498,N_2438);
xor U2654 (N_2654,N_2266,N_2284);
and U2655 (N_2655,N_2481,N_2365);
xor U2656 (N_2656,N_2487,N_2353);
nor U2657 (N_2657,N_2260,N_2498);
nor U2658 (N_2658,N_2343,N_2325);
nand U2659 (N_2659,N_2386,N_2368);
or U2660 (N_2660,N_2355,N_2263);
or U2661 (N_2661,N_2285,N_2368);
and U2662 (N_2662,N_2392,N_2376);
and U2663 (N_2663,N_2422,N_2315);
or U2664 (N_2664,N_2342,N_2271);
and U2665 (N_2665,N_2499,N_2355);
xnor U2666 (N_2666,N_2416,N_2257);
or U2667 (N_2667,N_2306,N_2261);
or U2668 (N_2668,N_2316,N_2414);
nand U2669 (N_2669,N_2300,N_2461);
and U2670 (N_2670,N_2481,N_2486);
nand U2671 (N_2671,N_2344,N_2459);
nand U2672 (N_2672,N_2423,N_2447);
nand U2673 (N_2673,N_2414,N_2431);
xor U2674 (N_2674,N_2462,N_2362);
nand U2675 (N_2675,N_2485,N_2326);
xor U2676 (N_2676,N_2325,N_2435);
xnor U2677 (N_2677,N_2388,N_2329);
or U2678 (N_2678,N_2387,N_2404);
or U2679 (N_2679,N_2324,N_2291);
nand U2680 (N_2680,N_2298,N_2303);
nand U2681 (N_2681,N_2336,N_2473);
and U2682 (N_2682,N_2258,N_2270);
and U2683 (N_2683,N_2262,N_2353);
xor U2684 (N_2684,N_2264,N_2258);
xnor U2685 (N_2685,N_2319,N_2404);
nor U2686 (N_2686,N_2385,N_2481);
xnor U2687 (N_2687,N_2487,N_2270);
xor U2688 (N_2688,N_2444,N_2378);
nor U2689 (N_2689,N_2413,N_2412);
and U2690 (N_2690,N_2281,N_2412);
nand U2691 (N_2691,N_2305,N_2332);
or U2692 (N_2692,N_2412,N_2431);
nor U2693 (N_2693,N_2425,N_2447);
nand U2694 (N_2694,N_2443,N_2373);
nor U2695 (N_2695,N_2360,N_2476);
nand U2696 (N_2696,N_2347,N_2384);
or U2697 (N_2697,N_2256,N_2487);
xor U2698 (N_2698,N_2254,N_2482);
xnor U2699 (N_2699,N_2291,N_2391);
xor U2700 (N_2700,N_2326,N_2304);
nor U2701 (N_2701,N_2406,N_2443);
xor U2702 (N_2702,N_2409,N_2320);
xnor U2703 (N_2703,N_2415,N_2495);
nor U2704 (N_2704,N_2416,N_2431);
xnor U2705 (N_2705,N_2476,N_2385);
or U2706 (N_2706,N_2364,N_2419);
nand U2707 (N_2707,N_2371,N_2327);
or U2708 (N_2708,N_2357,N_2437);
xnor U2709 (N_2709,N_2407,N_2417);
xnor U2710 (N_2710,N_2392,N_2293);
and U2711 (N_2711,N_2351,N_2436);
nor U2712 (N_2712,N_2271,N_2250);
nand U2713 (N_2713,N_2318,N_2367);
nor U2714 (N_2714,N_2300,N_2448);
nor U2715 (N_2715,N_2365,N_2467);
nand U2716 (N_2716,N_2391,N_2316);
xnor U2717 (N_2717,N_2342,N_2408);
or U2718 (N_2718,N_2295,N_2491);
xor U2719 (N_2719,N_2454,N_2498);
nor U2720 (N_2720,N_2252,N_2465);
and U2721 (N_2721,N_2477,N_2330);
or U2722 (N_2722,N_2341,N_2453);
nand U2723 (N_2723,N_2351,N_2421);
or U2724 (N_2724,N_2278,N_2422);
nor U2725 (N_2725,N_2478,N_2408);
or U2726 (N_2726,N_2365,N_2314);
xor U2727 (N_2727,N_2468,N_2383);
nor U2728 (N_2728,N_2329,N_2470);
and U2729 (N_2729,N_2275,N_2410);
and U2730 (N_2730,N_2495,N_2414);
and U2731 (N_2731,N_2256,N_2339);
and U2732 (N_2732,N_2478,N_2277);
xor U2733 (N_2733,N_2416,N_2355);
nand U2734 (N_2734,N_2343,N_2301);
xnor U2735 (N_2735,N_2272,N_2458);
nand U2736 (N_2736,N_2310,N_2339);
xor U2737 (N_2737,N_2394,N_2384);
and U2738 (N_2738,N_2381,N_2316);
and U2739 (N_2739,N_2309,N_2312);
nor U2740 (N_2740,N_2316,N_2464);
nand U2741 (N_2741,N_2294,N_2404);
nor U2742 (N_2742,N_2253,N_2313);
and U2743 (N_2743,N_2469,N_2461);
xnor U2744 (N_2744,N_2385,N_2465);
xor U2745 (N_2745,N_2465,N_2319);
nand U2746 (N_2746,N_2382,N_2317);
and U2747 (N_2747,N_2333,N_2309);
or U2748 (N_2748,N_2276,N_2323);
nand U2749 (N_2749,N_2485,N_2361);
nor U2750 (N_2750,N_2514,N_2609);
xnor U2751 (N_2751,N_2741,N_2555);
and U2752 (N_2752,N_2686,N_2643);
nand U2753 (N_2753,N_2518,N_2671);
xnor U2754 (N_2754,N_2717,N_2620);
nor U2755 (N_2755,N_2564,N_2687);
and U2756 (N_2756,N_2663,N_2523);
nand U2757 (N_2757,N_2612,N_2611);
nand U2758 (N_2758,N_2530,N_2700);
nor U2759 (N_2759,N_2639,N_2732);
nor U2760 (N_2760,N_2689,N_2571);
and U2761 (N_2761,N_2638,N_2578);
nor U2762 (N_2762,N_2657,N_2685);
nand U2763 (N_2763,N_2624,N_2544);
and U2764 (N_2764,N_2526,N_2708);
or U2765 (N_2765,N_2602,N_2522);
nor U2766 (N_2766,N_2510,N_2617);
nand U2767 (N_2767,N_2625,N_2749);
nor U2768 (N_2768,N_2633,N_2535);
or U2769 (N_2769,N_2576,N_2595);
xnor U2770 (N_2770,N_2582,N_2678);
or U2771 (N_2771,N_2721,N_2604);
nand U2772 (N_2772,N_2742,N_2740);
nand U2773 (N_2773,N_2531,N_2679);
nor U2774 (N_2774,N_2557,N_2527);
or U2775 (N_2775,N_2692,N_2683);
and U2776 (N_2776,N_2501,N_2727);
xor U2777 (N_2777,N_2647,N_2606);
nor U2778 (N_2778,N_2524,N_2723);
nor U2779 (N_2779,N_2634,N_2720);
and U2780 (N_2780,N_2709,N_2521);
xor U2781 (N_2781,N_2610,N_2574);
nand U2782 (N_2782,N_2696,N_2605);
and U2783 (N_2783,N_2559,N_2546);
nand U2784 (N_2784,N_2588,N_2619);
xnor U2785 (N_2785,N_2581,N_2599);
xor U2786 (N_2786,N_2715,N_2684);
or U2787 (N_2787,N_2681,N_2511);
xnor U2788 (N_2788,N_2600,N_2725);
nor U2789 (N_2789,N_2553,N_2738);
nor U2790 (N_2790,N_2666,N_2516);
nand U2791 (N_2791,N_2507,N_2699);
nand U2792 (N_2792,N_2734,N_2566);
nand U2793 (N_2793,N_2662,N_2573);
xnor U2794 (N_2794,N_2735,N_2693);
xor U2795 (N_2795,N_2677,N_2736);
xnor U2796 (N_2796,N_2744,N_2644);
and U2797 (N_2797,N_2691,N_2688);
nor U2798 (N_2798,N_2601,N_2669);
xnor U2799 (N_2799,N_2579,N_2575);
xnor U2800 (N_2800,N_2667,N_2690);
xnor U2801 (N_2801,N_2640,N_2710);
or U2802 (N_2802,N_2593,N_2558);
nand U2803 (N_2803,N_2550,N_2661);
nor U2804 (N_2804,N_2659,N_2655);
or U2805 (N_2805,N_2716,N_2665);
and U2806 (N_2806,N_2594,N_2707);
or U2807 (N_2807,N_2705,N_2551);
nand U2808 (N_2808,N_2728,N_2726);
xor U2809 (N_2809,N_2632,N_2713);
or U2810 (N_2810,N_2642,N_2569);
and U2811 (N_2811,N_2635,N_2508);
xor U2812 (N_2812,N_2517,N_2658);
nand U2813 (N_2813,N_2706,N_2672);
nor U2814 (N_2814,N_2654,N_2562);
or U2815 (N_2815,N_2695,N_2668);
nor U2816 (N_2816,N_2631,N_2556);
nor U2817 (N_2817,N_2701,N_2656);
nor U2818 (N_2818,N_2628,N_2743);
xnor U2819 (N_2819,N_2651,N_2512);
or U2820 (N_2820,N_2580,N_2591);
xnor U2821 (N_2821,N_2627,N_2560);
nand U2822 (N_2822,N_2676,N_2525);
or U2823 (N_2823,N_2731,N_2675);
or U2824 (N_2824,N_2548,N_2549);
or U2825 (N_2825,N_2577,N_2650);
nand U2826 (N_2826,N_2729,N_2583);
nor U2827 (N_2827,N_2653,N_2565);
nand U2828 (N_2828,N_2536,N_2636);
and U2829 (N_2829,N_2540,N_2509);
nor U2830 (N_2830,N_2621,N_2670);
nand U2831 (N_2831,N_2587,N_2589);
xor U2832 (N_2832,N_2704,N_2745);
or U2833 (N_2833,N_2592,N_2739);
xor U2834 (N_2834,N_2598,N_2630);
or U2835 (N_2835,N_2585,N_2534);
or U2836 (N_2836,N_2637,N_2733);
xnor U2837 (N_2837,N_2649,N_2513);
nor U2838 (N_2838,N_2722,N_2529);
nand U2839 (N_2839,N_2660,N_2680);
nor U2840 (N_2840,N_2682,N_2748);
nand U2841 (N_2841,N_2568,N_2623);
nand U2842 (N_2842,N_2505,N_2724);
xnor U2843 (N_2843,N_2652,N_2538);
nor U2844 (N_2844,N_2702,N_2626);
nand U2845 (N_2845,N_2641,N_2506);
nor U2846 (N_2846,N_2561,N_2618);
nand U2847 (N_2847,N_2515,N_2563);
nand U2848 (N_2848,N_2603,N_2572);
nor U2849 (N_2849,N_2570,N_2622);
or U2850 (N_2850,N_2615,N_2567);
nor U2851 (N_2851,N_2519,N_2629);
xnor U2852 (N_2852,N_2608,N_2586);
nand U2853 (N_2853,N_2547,N_2730);
nor U2854 (N_2854,N_2590,N_2614);
nand U2855 (N_2855,N_2545,N_2542);
nand U2856 (N_2856,N_2616,N_2664);
nand U2857 (N_2857,N_2503,N_2719);
nor U2858 (N_2858,N_2584,N_2502);
nor U2859 (N_2859,N_2645,N_2697);
and U2860 (N_2860,N_2543,N_2597);
or U2861 (N_2861,N_2500,N_2541);
xnor U2862 (N_2862,N_2504,N_2711);
and U2863 (N_2863,N_2698,N_2539);
and U2864 (N_2864,N_2646,N_2746);
xnor U2865 (N_2865,N_2607,N_2596);
or U2866 (N_2866,N_2554,N_2673);
and U2867 (N_2867,N_2712,N_2533);
nand U2868 (N_2868,N_2648,N_2737);
nor U2869 (N_2869,N_2694,N_2528);
nor U2870 (N_2870,N_2718,N_2537);
or U2871 (N_2871,N_2532,N_2714);
and U2872 (N_2872,N_2613,N_2703);
nor U2873 (N_2873,N_2552,N_2674);
or U2874 (N_2874,N_2520,N_2747);
nand U2875 (N_2875,N_2749,N_2539);
xnor U2876 (N_2876,N_2703,N_2616);
or U2877 (N_2877,N_2513,N_2719);
nand U2878 (N_2878,N_2689,N_2597);
and U2879 (N_2879,N_2635,N_2713);
nand U2880 (N_2880,N_2625,N_2570);
nor U2881 (N_2881,N_2555,N_2578);
nor U2882 (N_2882,N_2656,N_2668);
or U2883 (N_2883,N_2512,N_2657);
and U2884 (N_2884,N_2732,N_2667);
or U2885 (N_2885,N_2645,N_2512);
and U2886 (N_2886,N_2732,N_2700);
xor U2887 (N_2887,N_2731,N_2541);
and U2888 (N_2888,N_2611,N_2716);
or U2889 (N_2889,N_2599,N_2669);
or U2890 (N_2890,N_2640,N_2587);
nand U2891 (N_2891,N_2541,N_2680);
and U2892 (N_2892,N_2601,N_2699);
nand U2893 (N_2893,N_2585,N_2524);
nor U2894 (N_2894,N_2681,N_2580);
nor U2895 (N_2895,N_2641,N_2541);
and U2896 (N_2896,N_2740,N_2529);
or U2897 (N_2897,N_2517,N_2637);
nor U2898 (N_2898,N_2691,N_2527);
and U2899 (N_2899,N_2514,N_2694);
nand U2900 (N_2900,N_2520,N_2730);
or U2901 (N_2901,N_2552,N_2543);
xor U2902 (N_2902,N_2605,N_2611);
or U2903 (N_2903,N_2585,N_2723);
and U2904 (N_2904,N_2521,N_2529);
and U2905 (N_2905,N_2614,N_2730);
or U2906 (N_2906,N_2736,N_2559);
nor U2907 (N_2907,N_2577,N_2507);
nand U2908 (N_2908,N_2550,N_2626);
or U2909 (N_2909,N_2744,N_2568);
nand U2910 (N_2910,N_2594,N_2597);
or U2911 (N_2911,N_2580,N_2505);
or U2912 (N_2912,N_2654,N_2503);
xnor U2913 (N_2913,N_2625,N_2589);
nor U2914 (N_2914,N_2674,N_2669);
or U2915 (N_2915,N_2634,N_2625);
xnor U2916 (N_2916,N_2560,N_2555);
and U2917 (N_2917,N_2643,N_2507);
nor U2918 (N_2918,N_2740,N_2533);
and U2919 (N_2919,N_2673,N_2749);
nor U2920 (N_2920,N_2673,N_2520);
xnor U2921 (N_2921,N_2607,N_2646);
xnor U2922 (N_2922,N_2671,N_2637);
xor U2923 (N_2923,N_2609,N_2657);
and U2924 (N_2924,N_2676,N_2558);
and U2925 (N_2925,N_2502,N_2553);
or U2926 (N_2926,N_2674,N_2627);
or U2927 (N_2927,N_2724,N_2679);
xor U2928 (N_2928,N_2617,N_2638);
nand U2929 (N_2929,N_2587,N_2644);
or U2930 (N_2930,N_2640,N_2554);
nor U2931 (N_2931,N_2744,N_2707);
nand U2932 (N_2932,N_2533,N_2564);
and U2933 (N_2933,N_2748,N_2645);
and U2934 (N_2934,N_2596,N_2622);
nand U2935 (N_2935,N_2552,N_2548);
nand U2936 (N_2936,N_2502,N_2635);
or U2937 (N_2937,N_2584,N_2737);
nand U2938 (N_2938,N_2602,N_2730);
nor U2939 (N_2939,N_2630,N_2578);
xnor U2940 (N_2940,N_2714,N_2631);
and U2941 (N_2941,N_2664,N_2707);
or U2942 (N_2942,N_2572,N_2517);
xor U2943 (N_2943,N_2611,N_2560);
and U2944 (N_2944,N_2697,N_2702);
and U2945 (N_2945,N_2622,N_2512);
nor U2946 (N_2946,N_2535,N_2664);
nand U2947 (N_2947,N_2623,N_2679);
xnor U2948 (N_2948,N_2561,N_2599);
or U2949 (N_2949,N_2536,N_2523);
nor U2950 (N_2950,N_2533,N_2585);
xnor U2951 (N_2951,N_2686,N_2731);
or U2952 (N_2952,N_2595,N_2653);
nor U2953 (N_2953,N_2534,N_2695);
nand U2954 (N_2954,N_2735,N_2709);
and U2955 (N_2955,N_2698,N_2611);
xor U2956 (N_2956,N_2648,N_2643);
or U2957 (N_2957,N_2517,N_2715);
nor U2958 (N_2958,N_2701,N_2703);
or U2959 (N_2959,N_2706,N_2513);
nor U2960 (N_2960,N_2587,N_2546);
nand U2961 (N_2961,N_2521,N_2624);
xnor U2962 (N_2962,N_2569,N_2660);
or U2963 (N_2963,N_2560,N_2682);
xnor U2964 (N_2964,N_2709,N_2581);
xor U2965 (N_2965,N_2633,N_2576);
or U2966 (N_2966,N_2720,N_2701);
nand U2967 (N_2967,N_2603,N_2619);
or U2968 (N_2968,N_2568,N_2587);
and U2969 (N_2969,N_2522,N_2541);
nor U2970 (N_2970,N_2618,N_2705);
xnor U2971 (N_2971,N_2566,N_2647);
or U2972 (N_2972,N_2518,N_2572);
nor U2973 (N_2973,N_2562,N_2648);
xor U2974 (N_2974,N_2554,N_2566);
or U2975 (N_2975,N_2704,N_2747);
xnor U2976 (N_2976,N_2576,N_2548);
and U2977 (N_2977,N_2698,N_2660);
nand U2978 (N_2978,N_2630,N_2729);
nand U2979 (N_2979,N_2587,N_2509);
or U2980 (N_2980,N_2586,N_2549);
nor U2981 (N_2981,N_2720,N_2544);
nand U2982 (N_2982,N_2620,N_2538);
nand U2983 (N_2983,N_2715,N_2553);
xnor U2984 (N_2984,N_2536,N_2646);
and U2985 (N_2985,N_2737,N_2721);
nor U2986 (N_2986,N_2523,N_2747);
and U2987 (N_2987,N_2738,N_2549);
nand U2988 (N_2988,N_2674,N_2712);
nor U2989 (N_2989,N_2543,N_2609);
or U2990 (N_2990,N_2740,N_2582);
nor U2991 (N_2991,N_2584,N_2554);
and U2992 (N_2992,N_2729,N_2711);
or U2993 (N_2993,N_2620,N_2509);
and U2994 (N_2994,N_2675,N_2666);
xnor U2995 (N_2995,N_2582,N_2567);
and U2996 (N_2996,N_2675,N_2586);
or U2997 (N_2997,N_2687,N_2646);
and U2998 (N_2998,N_2573,N_2594);
or U2999 (N_2999,N_2696,N_2590);
nand U3000 (N_3000,N_2872,N_2841);
nand U3001 (N_3001,N_2851,N_2995);
or U3002 (N_3002,N_2843,N_2998);
nor U3003 (N_3003,N_2877,N_2986);
nor U3004 (N_3004,N_2768,N_2988);
xnor U3005 (N_3005,N_2767,N_2867);
xor U3006 (N_3006,N_2825,N_2908);
nand U3007 (N_3007,N_2903,N_2773);
or U3008 (N_3008,N_2982,N_2922);
nand U3009 (N_3009,N_2751,N_2756);
nor U3010 (N_3010,N_2920,N_2847);
nand U3011 (N_3011,N_2848,N_2772);
nand U3012 (N_3012,N_2792,N_2927);
and U3013 (N_3013,N_2891,N_2961);
or U3014 (N_3014,N_2952,N_2974);
and U3015 (N_3015,N_2786,N_2972);
or U3016 (N_3016,N_2973,N_2858);
or U3017 (N_3017,N_2758,N_2888);
xnor U3018 (N_3018,N_2889,N_2942);
xor U3019 (N_3019,N_2919,N_2782);
xnor U3020 (N_3020,N_2793,N_2983);
and U3021 (N_3021,N_2959,N_2779);
xnor U3022 (N_3022,N_2951,N_2869);
xor U3023 (N_3023,N_2762,N_2814);
nand U3024 (N_3024,N_2956,N_2791);
nor U3025 (N_3025,N_2913,N_2999);
xor U3026 (N_3026,N_2945,N_2829);
xor U3027 (N_3027,N_2895,N_2804);
nor U3028 (N_3028,N_2921,N_2776);
or U3029 (N_3029,N_2834,N_2930);
xnor U3030 (N_3030,N_2898,N_2909);
nor U3031 (N_3031,N_2831,N_2975);
or U3032 (N_3032,N_2868,N_2781);
and U3033 (N_3033,N_2822,N_2996);
xnor U3034 (N_3034,N_2783,N_2940);
xor U3035 (N_3035,N_2980,N_2997);
nand U3036 (N_3036,N_2977,N_2764);
or U3037 (N_3037,N_2830,N_2795);
nand U3038 (N_3038,N_2981,N_2857);
nand U3039 (N_3039,N_2862,N_2842);
nand U3040 (N_3040,N_2810,N_2885);
xnor U3041 (N_3041,N_2876,N_2969);
nand U3042 (N_3042,N_2800,N_2901);
xor U3043 (N_3043,N_2991,N_2778);
or U3044 (N_3044,N_2864,N_2811);
or U3045 (N_3045,N_2798,N_2802);
or U3046 (N_3046,N_2759,N_2949);
nand U3047 (N_3047,N_2849,N_2929);
or U3048 (N_3048,N_2761,N_2854);
or U3049 (N_3049,N_2911,N_2883);
nand U3050 (N_3050,N_2866,N_2939);
xnor U3051 (N_3051,N_2806,N_2875);
nor U3052 (N_3052,N_2808,N_2989);
nand U3053 (N_3053,N_2887,N_2787);
xnor U3054 (N_3054,N_2984,N_2860);
xor U3055 (N_3055,N_2985,N_2979);
xor U3056 (N_3056,N_2839,N_2987);
and U3057 (N_3057,N_2846,N_2923);
or U3058 (N_3058,N_2906,N_2904);
or U3059 (N_3059,N_2790,N_2957);
nand U3060 (N_3060,N_2816,N_2993);
and U3061 (N_3061,N_2917,N_2976);
xor U3062 (N_3062,N_2879,N_2836);
and U3063 (N_3063,N_2852,N_2832);
xor U3064 (N_3064,N_2893,N_2912);
or U3065 (N_3065,N_2937,N_2935);
nand U3066 (N_3066,N_2850,N_2838);
or U3067 (N_3067,N_2833,N_2837);
nor U3068 (N_3068,N_2819,N_2915);
xor U3069 (N_3069,N_2924,N_2907);
or U3070 (N_3070,N_2775,N_2824);
and U3071 (N_3071,N_2941,N_2859);
nand U3072 (N_3072,N_2785,N_2865);
nor U3073 (N_3073,N_2962,N_2902);
nor U3074 (N_3074,N_2827,N_2820);
xnor U3075 (N_3075,N_2788,N_2944);
and U3076 (N_3076,N_2763,N_2789);
nor U3077 (N_3077,N_2966,N_2946);
nor U3078 (N_3078,N_2886,N_2807);
nor U3079 (N_3079,N_2803,N_2938);
xnor U3080 (N_3080,N_2784,N_2884);
or U3081 (N_3081,N_2896,N_2840);
and U3082 (N_3082,N_2916,N_2871);
nor U3083 (N_3083,N_2928,N_2823);
xnor U3084 (N_3084,N_2815,N_2809);
xnor U3085 (N_3085,N_2934,N_2948);
or U3086 (N_3086,N_2978,N_2855);
or U3087 (N_3087,N_2965,N_2878);
or U3088 (N_3088,N_2818,N_2958);
and U3089 (N_3089,N_2821,N_2954);
nand U3090 (N_3090,N_2757,N_2794);
xor U3091 (N_3091,N_2967,N_2835);
xnor U3092 (N_3092,N_2796,N_2766);
nor U3093 (N_3093,N_2918,N_2994);
nor U3094 (N_3094,N_2774,N_2953);
and U3095 (N_3095,N_2752,N_2968);
xnor U3096 (N_3096,N_2894,N_2760);
nand U3097 (N_3097,N_2897,N_2755);
or U3098 (N_3098,N_2828,N_2890);
and U3099 (N_3099,N_2955,N_2936);
nand U3100 (N_3100,N_2769,N_2990);
xnor U3101 (N_3101,N_2797,N_2899);
nor U3102 (N_3102,N_2964,N_2771);
and U3103 (N_3103,N_2932,N_2844);
nand U3104 (N_3104,N_2931,N_2856);
and U3105 (N_3105,N_2817,N_2750);
xor U3106 (N_3106,N_2777,N_2765);
xor U3107 (N_3107,N_2770,N_2826);
nor U3108 (N_3108,N_2947,N_2925);
xnor U3109 (N_3109,N_2905,N_2892);
or U3110 (N_3110,N_2910,N_2874);
nor U3111 (N_3111,N_2926,N_2971);
nor U3112 (N_3112,N_2853,N_2950);
and U3113 (N_3113,N_2943,N_2900);
nand U3114 (N_3114,N_2880,N_2933);
xor U3115 (N_3115,N_2882,N_2805);
nand U3116 (N_3116,N_2992,N_2813);
nor U3117 (N_3117,N_2812,N_2970);
xnor U3118 (N_3118,N_2873,N_2914);
xor U3119 (N_3119,N_2780,N_2753);
xnor U3120 (N_3120,N_2845,N_2799);
nor U3121 (N_3121,N_2960,N_2870);
and U3122 (N_3122,N_2881,N_2754);
nand U3123 (N_3123,N_2863,N_2963);
or U3124 (N_3124,N_2861,N_2801);
or U3125 (N_3125,N_2992,N_2863);
or U3126 (N_3126,N_2857,N_2893);
nand U3127 (N_3127,N_2947,N_2930);
nor U3128 (N_3128,N_2828,N_2905);
nand U3129 (N_3129,N_2984,N_2806);
nor U3130 (N_3130,N_2837,N_2790);
xnor U3131 (N_3131,N_2876,N_2964);
nor U3132 (N_3132,N_2753,N_2833);
xor U3133 (N_3133,N_2774,N_2934);
nor U3134 (N_3134,N_2982,N_2986);
nand U3135 (N_3135,N_2845,N_2863);
nor U3136 (N_3136,N_2997,N_2835);
nand U3137 (N_3137,N_2750,N_2852);
nor U3138 (N_3138,N_2951,N_2919);
xnor U3139 (N_3139,N_2794,N_2975);
and U3140 (N_3140,N_2944,N_2993);
or U3141 (N_3141,N_2812,N_2791);
nand U3142 (N_3142,N_2869,N_2775);
or U3143 (N_3143,N_2940,N_2837);
or U3144 (N_3144,N_2908,N_2809);
nand U3145 (N_3145,N_2815,N_2867);
and U3146 (N_3146,N_2868,N_2940);
nand U3147 (N_3147,N_2864,N_2980);
and U3148 (N_3148,N_2941,N_2755);
nand U3149 (N_3149,N_2811,N_2776);
or U3150 (N_3150,N_2941,N_2753);
nand U3151 (N_3151,N_2863,N_2806);
nor U3152 (N_3152,N_2813,N_2815);
nor U3153 (N_3153,N_2806,N_2897);
nand U3154 (N_3154,N_2768,N_2905);
or U3155 (N_3155,N_2911,N_2777);
xnor U3156 (N_3156,N_2963,N_2765);
xnor U3157 (N_3157,N_2831,N_2771);
xor U3158 (N_3158,N_2867,N_2875);
or U3159 (N_3159,N_2914,N_2843);
and U3160 (N_3160,N_2975,N_2774);
or U3161 (N_3161,N_2890,N_2982);
nor U3162 (N_3162,N_2981,N_2921);
nor U3163 (N_3163,N_2915,N_2834);
xnor U3164 (N_3164,N_2944,N_2800);
or U3165 (N_3165,N_2755,N_2808);
nor U3166 (N_3166,N_2906,N_2860);
nor U3167 (N_3167,N_2847,N_2940);
nand U3168 (N_3168,N_2917,N_2951);
and U3169 (N_3169,N_2884,N_2765);
nor U3170 (N_3170,N_2805,N_2775);
or U3171 (N_3171,N_2787,N_2801);
xor U3172 (N_3172,N_2771,N_2808);
nand U3173 (N_3173,N_2953,N_2876);
nand U3174 (N_3174,N_2840,N_2861);
xor U3175 (N_3175,N_2900,N_2778);
nor U3176 (N_3176,N_2831,N_2948);
xor U3177 (N_3177,N_2985,N_2924);
nand U3178 (N_3178,N_2834,N_2872);
nor U3179 (N_3179,N_2760,N_2925);
or U3180 (N_3180,N_2791,N_2881);
xor U3181 (N_3181,N_2796,N_2802);
and U3182 (N_3182,N_2759,N_2914);
nor U3183 (N_3183,N_2927,N_2795);
xor U3184 (N_3184,N_2816,N_2926);
xnor U3185 (N_3185,N_2970,N_2909);
and U3186 (N_3186,N_2955,N_2910);
or U3187 (N_3187,N_2798,N_2826);
nor U3188 (N_3188,N_2827,N_2771);
nor U3189 (N_3189,N_2911,N_2985);
xor U3190 (N_3190,N_2805,N_2840);
nor U3191 (N_3191,N_2767,N_2801);
and U3192 (N_3192,N_2827,N_2955);
xnor U3193 (N_3193,N_2802,N_2857);
xnor U3194 (N_3194,N_2892,N_2817);
nor U3195 (N_3195,N_2891,N_2805);
nor U3196 (N_3196,N_2759,N_2795);
nor U3197 (N_3197,N_2777,N_2918);
nor U3198 (N_3198,N_2796,N_2895);
and U3199 (N_3199,N_2856,N_2771);
and U3200 (N_3200,N_2843,N_2975);
nand U3201 (N_3201,N_2750,N_2870);
and U3202 (N_3202,N_2866,N_2837);
nand U3203 (N_3203,N_2984,N_2894);
and U3204 (N_3204,N_2920,N_2990);
or U3205 (N_3205,N_2865,N_2796);
nand U3206 (N_3206,N_2875,N_2952);
or U3207 (N_3207,N_2794,N_2836);
nor U3208 (N_3208,N_2893,N_2760);
nor U3209 (N_3209,N_2930,N_2931);
and U3210 (N_3210,N_2974,N_2798);
nand U3211 (N_3211,N_2772,N_2963);
and U3212 (N_3212,N_2903,N_2955);
or U3213 (N_3213,N_2783,N_2936);
or U3214 (N_3214,N_2889,N_2963);
or U3215 (N_3215,N_2805,N_2868);
nand U3216 (N_3216,N_2853,N_2872);
and U3217 (N_3217,N_2911,N_2799);
nor U3218 (N_3218,N_2861,N_2796);
xnor U3219 (N_3219,N_2913,N_2812);
or U3220 (N_3220,N_2912,N_2985);
or U3221 (N_3221,N_2794,N_2899);
nand U3222 (N_3222,N_2948,N_2808);
and U3223 (N_3223,N_2941,N_2897);
and U3224 (N_3224,N_2975,N_2894);
or U3225 (N_3225,N_2886,N_2771);
nor U3226 (N_3226,N_2772,N_2880);
or U3227 (N_3227,N_2980,N_2985);
and U3228 (N_3228,N_2868,N_2918);
xnor U3229 (N_3229,N_2981,N_2820);
nor U3230 (N_3230,N_2836,N_2761);
xor U3231 (N_3231,N_2850,N_2825);
xnor U3232 (N_3232,N_2757,N_2804);
xnor U3233 (N_3233,N_2923,N_2909);
nand U3234 (N_3234,N_2911,N_2862);
xor U3235 (N_3235,N_2808,N_2983);
or U3236 (N_3236,N_2933,N_2976);
nor U3237 (N_3237,N_2956,N_2928);
and U3238 (N_3238,N_2910,N_2937);
nor U3239 (N_3239,N_2974,N_2938);
and U3240 (N_3240,N_2871,N_2977);
or U3241 (N_3241,N_2937,N_2785);
and U3242 (N_3242,N_2771,N_2928);
nand U3243 (N_3243,N_2825,N_2978);
and U3244 (N_3244,N_2800,N_2973);
nor U3245 (N_3245,N_2857,N_2982);
or U3246 (N_3246,N_2883,N_2858);
and U3247 (N_3247,N_2941,N_2975);
xor U3248 (N_3248,N_2951,N_2857);
or U3249 (N_3249,N_2903,N_2894);
or U3250 (N_3250,N_3238,N_3134);
xnor U3251 (N_3251,N_3056,N_3024);
nor U3252 (N_3252,N_3090,N_3203);
nand U3253 (N_3253,N_3248,N_3174);
nor U3254 (N_3254,N_3015,N_3006);
xor U3255 (N_3255,N_3013,N_3144);
and U3256 (N_3256,N_3055,N_3150);
nor U3257 (N_3257,N_3119,N_3147);
or U3258 (N_3258,N_3053,N_3139);
nor U3259 (N_3259,N_3127,N_3035);
nand U3260 (N_3260,N_3033,N_3072);
nor U3261 (N_3261,N_3027,N_3133);
xor U3262 (N_3262,N_3003,N_3224);
xor U3263 (N_3263,N_3047,N_3069);
and U3264 (N_3264,N_3014,N_3121);
nor U3265 (N_3265,N_3219,N_3114);
xor U3266 (N_3266,N_3026,N_3247);
nand U3267 (N_3267,N_3142,N_3039);
nor U3268 (N_3268,N_3156,N_3017);
nor U3269 (N_3269,N_3152,N_3223);
nand U3270 (N_3270,N_3159,N_3103);
nor U3271 (N_3271,N_3001,N_3073);
xor U3272 (N_3272,N_3239,N_3111);
and U3273 (N_3273,N_3200,N_3020);
or U3274 (N_3274,N_3089,N_3234);
nor U3275 (N_3275,N_3209,N_3148);
or U3276 (N_3276,N_3197,N_3045);
or U3277 (N_3277,N_3201,N_3226);
nand U3278 (N_3278,N_3083,N_3093);
or U3279 (N_3279,N_3155,N_3048);
xor U3280 (N_3280,N_3168,N_3004);
or U3281 (N_3281,N_3188,N_3067);
xnor U3282 (N_3282,N_3171,N_3176);
and U3283 (N_3283,N_3204,N_3051);
and U3284 (N_3284,N_3080,N_3005);
xnor U3285 (N_3285,N_3194,N_3059);
xor U3286 (N_3286,N_3216,N_3158);
and U3287 (N_3287,N_3215,N_3102);
or U3288 (N_3288,N_3044,N_3143);
nor U3289 (N_3289,N_3118,N_3208);
xor U3290 (N_3290,N_3079,N_3011);
xnor U3291 (N_3291,N_3207,N_3129);
nand U3292 (N_3292,N_3122,N_3125);
xor U3293 (N_3293,N_3228,N_3240);
or U3294 (N_3294,N_3076,N_3242);
nand U3295 (N_3295,N_3175,N_3243);
nor U3296 (N_3296,N_3153,N_3177);
nor U3297 (N_3297,N_3138,N_3008);
xor U3298 (N_3298,N_3101,N_3236);
or U3299 (N_3299,N_3030,N_3164);
nand U3300 (N_3300,N_3227,N_3063);
nand U3301 (N_3301,N_3041,N_3066);
xor U3302 (N_3302,N_3211,N_3043);
nor U3303 (N_3303,N_3120,N_3112);
or U3304 (N_3304,N_3098,N_3022);
xnor U3305 (N_3305,N_3070,N_3222);
nor U3306 (N_3306,N_3113,N_3212);
nand U3307 (N_3307,N_3179,N_3034);
or U3308 (N_3308,N_3091,N_3166);
and U3309 (N_3309,N_3085,N_3007);
nand U3310 (N_3310,N_3092,N_3115);
nand U3311 (N_3311,N_3145,N_3191);
and U3312 (N_3312,N_3124,N_3135);
xnor U3313 (N_3313,N_3202,N_3206);
or U3314 (N_3314,N_3105,N_3185);
or U3315 (N_3315,N_3050,N_3016);
nor U3316 (N_3316,N_3009,N_3104);
or U3317 (N_3317,N_3163,N_3193);
nand U3318 (N_3318,N_3237,N_3196);
xnor U3319 (N_3319,N_3075,N_3021);
xor U3320 (N_3320,N_3169,N_3181);
nor U3321 (N_3321,N_3217,N_3157);
xnor U3322 (N_3322,N_3231,N_3082);
xor U3323 (N_3323,N_3146,N_3213);
nand U3324 (N_3324,N_3040,N_3097);
xor U3325 (N_3325,N_3096,N_3140);
or U3326 (N_3326,N_3019,N_3167);
and U3327 (N_3327,N_3162,N_3086);
or U3328 (N_3328,N_3099,N_3198);
or U3329 (N_3329,N_3221,N_3108);
and U3330 (N_3330,N_3052,N_3100);
nand U3331 (N_3331,N_3184,N_3235);
and U3332 (N_3332,N_3064,N_3106);
xnor U3333 (N_3333,N_3165,N_3232);
or U3334 (N_3334,N_3154,N_3058);
nor U3335 (N_3335,N_3189,N_3084);
and U3336 (N_3336,N_3136,N_3229);
or U3337 (N_3337,N_3186,N_3032);
and U3338 (N_3338,N_3062,N_3061);
nor U3339 (N_3339,N_3131,N_3029);
nand U3340 (N_3340,N_3220,N_3225);
and U3341 (N_3341,N_3128,N_3246);
nor U3342 (N_3342,N_3110,N_3025);
xor U3343 (N_3343,N_3094,N_3160);
nand U3344 (N_3344,N_3054,N_3183);
nand U3345 (N_3345,N_3095,N_3151);
nor U3346 (N_3346,N_3195,N_3010);
nor U3347 (N_3347,N_3130,N_3081);
nor U3348 (N_3348,N_3057,N_3249);
or U3349 (N_3349,N_3199,N_3107);
or U3350 (N_3350,N_3074,N_3187);
nand U3351 (N_3351,N_3028,N_3210);
nand U3352 (N_3352,N_3233,N_3087);
or U3353 (N_3353,N_3065,N_3117);
nand U3354 (N_3354,N_3245,N_3214);
nor U3355 (N_3355,N_3088,N_3192);
or U3356 (N_3356,N_3002,N_3123);
nand U3357 (N_3357,N_3077,N_3023);
xnor U3358 (N_3358,N_3161,N_3126);
and U3359 (N_3359,N_3137,N_3012);
nand U3360 (N_3360,N_3218,N_3018);
nor U3361 (N_3361,N_3170,N_3230);
xnor U3362 (N_3362,N_3037,N_3180);
xor U3363 (N_3363,N_3049,N_3182);
nor U3364 (N_3364,N_3190,N_3078);
xnor U3365 (N_3365,N_3141,N_3042);
nand U3366 (N_3366,N_3149,N_3244);
and U3367 (N_3367,N_3109,N_3060);
or U3368 (N_3368,N_3241,N_3132);
or U3369 (N_3369,N_3068,N_3205);
xnor U3370 (N_3370,N_3173,N_3046);
xor U3371 (N_3371,N_3000,N_3038);
or U3372 (N_3372,N_3116,N_3036);
xnor U3373 (N_3373,N_3031,N_3071);
or U3374 (N_3374,N_3172,N_3178);
nor U3375 (N_3375,N_3046,N_3151);
or U3376 (N_3376,N_3062,N_3212);
nand U3377 (N_3377,N_3225,N_3169);
or U3378 (N_3378,N_3173,N_3095);
nor U3379 (N_3379,N_3236,N_3006);
nand U3380 (N_3380,N_3057,N_3114);
nand U3381 (N_3381,N_3070,N_3043);
or U3382 (N_3382,N_3062,N_3089);
or U3383 (N_3383,N_3015,N_3070);
nand U3384 (N_3384,N_3044,N_3165);
and U3385 (N_3385,N_3158,N_3072);
nand U3386 (N_3386,N_3030,N_3241);
nor U3387 (N_3387,N_3079,N_3068);
nor U3388 (N_3388,N_3072,N_3049);
xor U3389 (N_3389,N_3153,N_3146);
and U3390 (N_3390,N_3152,N_3163);
xnor U3391 (N_3391,N_3012,N_3032);
xor U3392 (N_3392,N_3050,N_3094);
or U3393 (N_3393,N_3185,N_3098);
xnor U3394 (N_3394,N_3094,N_3143);
nor U3395 (N_3395,N_3228,N_3148);
or U3396 (N_3396,N_3037,N_3030);
or U3397 (N_3397,N_3199,N_3179);
and U3398 (N_3398,N_3235,N_3187);
xor U3399 (N_3399,N_3120,N_3157);
xor U3400 (N_3400,N_3102,N_3143);
and U3401 (N_3401,N_3126,N_3030);
or U3402 (N_3402,N_3087,N_3084);
nand U3403 (N_3403,N_3148,N_3020);
or U3404 (N_3404,N_3129,N_3091);
nand U3405 (N_3405,N_3235,N_3196);
nor U3406 (N_3406,N_3015,N_3096);
or U3407 (N_3407,N_3071,N_3168);
nand U3408 (N_3408,N_3177,N_3014);
xnor U3409 (N_3409,N_3067,N_3122);
or U3410 (N_3410,N_3033,N_3182);
and U3411 (N_3411,N_3216,N_3007);
xor U3412 (N_3412,N_3235,N_3150);
nor U3413 (N_3413,N_3105,N_3089);
and U3414 (N_3414,N_3159,N_3233);
xnor U3415 (N_3415,N_3126,N_3008);
nor U3416 (N_3416,N_3157,N_3211);
nor U3417 (N_3417,N_3173,N_3157);
xnor U3418 (N_3418,N_3173,N_3205);
xor U3419 (N_3419,N_3086,N_3096);
nor U3420 (N_3420,N_3008,N_3228);
and U3421 (N_3421,N_3026,N_3088);
and U3422 (N_3422,N_3095,N_3141);
nor U3423 (N_3423,N_3037,N_3049);
nor U3424 (N_3424,N_3240,N_3010);
and U3425 (N_3425,N_3211,N_3199);
nand U3426 (N_3426,N_3068,N_3118);
or U3427 (N_3427,N_3183,N_3212);
or U3428 (N_3428,N_3181,N_3114);
or U3429 (N_3429,N_3034,N_3145);
nor U3430 (N_3430,N_3122,N_3018);
or U3431 (N_3431,N_3209,N_3135);
xnor U3432 (N_3432,N_3111,N_3060);
or U3433 (N_3433,N_3183,N_3102);
and U3434 (N_3434,N_3050,N_3159);
nor U3435 (N_3435,N_3193,N_3082);
nand U3436 (N_3436,N_3199,N_3186);
nor U3437 (N_3437,N_3129,N_3222);
or U3438 (N_3438,N_3040,N_3129);
or U3439 (N_3439,N_3150,N_3231);
or U3440 (N_3440,N_3107,N_3231);
or U3441 (N_3441,N_3150,N_3103);
nor U3442 (N_3442,N_3065,N_3239);
or U3443 (N_3443,N_3089,N_3082);
xnor U3444 (N_3444,N_3151,N_3056);
xnor U3445 (N_3445,N_3201,N_3187);
nand U3446 (N_3446,N_3056,N_3187);
nor U3447 (N_3447,N_3072,N_3089);
nor U3448 (N_3448,N_3241,N_3044);
nand U3449 (N_3449,N_3015,N_3122);
or U3450 (N_3450,N_3175,N_3158);
xor U3451 (N_3451,N_3202,N_3121);
xnor U3452 (N_3452,N_3134,N_3111);
nor U3453 (N_3453,N_3187,N_3138);
or U3454 (N_3454,N_3224,N_3077);
and U3455 (N_3455,N_3077,N_3054);
and U3456 (N_3456,N_3106,N_3128);
and U3457 (N_3457,N_3166,N_3178);
or U3458 (N_3458,N_3170,N_3048);
nor U3459 (N_3459,N_3228,N_3052);
xor U3460 (N_3460,N_3209,N_3115);
nand U3461 (N_3461,N_3113,N_3074);
nand U3462 (N_3462,N_3053,N_3010);
and U3463 (N_3463,N_3224,N_3235);
and U3464 (N_3464,N_3179,N_3200);
or U3465 (N_3465,N_3084,N_3121);
xor U3466 (N_3466,N_3082,N_3214);
and U3467 (N_3467,N_3049,N_3091);
nand U3468 (N_3468,N_3033,N_3071);
nor U3469 (N_3469,N_3169,N_3007);
nor U3470 (N_3470,N_3171,N_3014);
nor U3471 (N_3471,N_3233,N_3202);
and U3472 (N_3472,N_3087,N_3239);
and U3473 (N_3473,N_3099,N_3167);
nor U3474 (N_3474,N_3167,N_3127);
xor U3475 (N_3475,N_3197,N_3053);
nand U3476 (N_3476,N_3204,N_3154);
nor U3477 (N_3477,N_3194,N_3228);
nor U3478 (N_3478,N_3196,N_3145);
nand U3479 (N_3479,N_3067,N_3130);
nand U3480 (N_3480,N_3152,N_3244);
nand U3481 (N_3481,N_3036,N_3223);
nor U3482 (N_3482,N_3061,N_3109);
nand U3483 (N_3483,N_3211,N_3239);
nor U3484 (N_3484,N_3077,N_3194);
and U3485 (N_3485,N_3245,N_3133);
nand U3486 (N_3486,N_3096,N_3109);
xnor U3487 (N_3487,N_3072,N_3199);
or U3488 (N_3488,N_3207,N_3226);
nand U3489 (N_3489,N_3148,N_3245);
nand U3490 (N_3490,N_3229,N_3027);
xnor U3491 (N_3491,N_3142,N_3172);
nand U3492 (N_3492,N_3246,N_3231);
and U3493 (N_3493,N_3196,N_3097);
xor U3494 (N_3494,N_3034,N_3222);
and U3495 (N_3495,N_3214,N_3213);
xnor U3496 (N_3496,N_3226,N_3003);
nor U3497 (N_3497,N_3234,N_3174);
xnor U3498 (N_3498,N_3056,N_3180);
or U3499 (N_3499,N_3111,N_3112);
nor U3500 (N_3500,N_3380,N_3469);
and U3501 (N_3501,N_3348,N_3361);
nand U3502 (N_3502,N_3287,N_3288);
or U3503 (N_3503,N_3280,N_3381);
and U3504 (N_3504,N_3303,N_3305);
nor U3505 (N_3505,N_3267,N_3443);
nor U3506 (N_3506,N_3256,N_3499);
xor U3507 (N_3507,N_3418,N_3415);
or U3508 (N_3508,N_3286,N_3299);
nor U3509 (N_3509,N_3320,N_3346);
and U3510 (N_3510,N_3301,N_3457);
xor U3511 (N_3511,N_3273,N_3324);
and U3512 (N_3512,N_3485,N_3399);
nor U3513 (N_3513,N_3360,N_3482);
and U3514 (N_3514,N_3385,N_3284);
or U3515 (N_3515,N_3494,N_3438);
nor U3516 (N_3516,N_3261,N_3474);
or U3517 (N_3517,N_3363,N_3362);
and U3518 (N_3518,N_3294,N_3274);
nand U3519 (N_3519,N_3336,N_3251);
and U3520 (N_3520,N_3424,N_3292);
nor U3521 (N_3521,N_3444,N_3341);
nand U3522 (N_3522,N_3400,N_3442);
and U3523 (N_3523,N_3429,N_3460);
and U3524 (N_3524,N_3340,N_3473);
nand U3525 (N_3525,N_3258,N_3322);
xnor U3526 (N_3526,N_3271,N_3426);
and U3527 (N_3527,N_3488,N_3327);
nor U3528 (N_3528,N_3465,N_3475);
nor U3529 (N_3529,N_3479,N_3419);
xnor U3530 (N_3530,N_3383,N_3382);
nand U3531 (N_3531,N_3358,N_3349);
and U3532 (N_3532,N_3262,N_3253);
nand U3533 (N_3533,N_3338,N_3276);
xnor U3534 (N_3534,N_3372,N_3441);
xor U3535 (N_3535,N_3422,N_3490);
xnor U3536 (N_3536,N_3480,N_3483);
xnor U3537 (N_3537,N_3455,N_3407);
or U3538 (N_3538,N_3263,N_3466);
or U3539 (N_3539,N_3272,N_3334);
or U3540 (N_3540,N_3282,N_3376);
nand U3541 (N_3541,N_3255,N_3312);
xnor U3542 (N_3542,N_3329,N_3411);
nand U3543 (N_3543,N_3302,N_3345);
or U3544 (N_3544,N_3357,N_3342);
nor U3545 (N_3545,N_3291,N_3497);
nor U3546 (N_3546,N_3277,N_3498);
nand U3547 (N_3547,N_3454,N_3391);
nor U3548 (N_3548,N_3353,N_3436);
or U3549 (N_3549,N_3264,N_3359);
nor U3550 (N_3550,N_3319,N_3468);
nand U3551 (N_3551,N_3484,N_3311);
or U3552 (N_3552,N_3471,N_3367);
and U3553 (N_3553,N_3478,N_3417);
nand U3554 (N_3554,N_3459,N_3326);
xor U3555 (N_3555,N_3386,N_3423);
or U3556 (N_3556,N_3456,N_3476);
or U3557 (N_3557,N_3496,N_3265);
or U3558 (N_3558,N_3318,N_3278);
xnor U3559 (N_3559,N_3293,N_3308);
nor U3560 (N_3560,N_3435,N_3392);
or U3561 (N_3561,N_3495,N_3332);
xor U3562 (N_3562,N_3390,N_3355);
and U3563 (N_3563,N_3289,N_3270);
xnor U3564 (N_3564,N_3492,N_3304);
or U3565 (N_3565,N_3446,N_3354);
and U3566 (N_3566,N_3493,N_3281);
or U3567 (N_3567,N_3445,N_3409);
or U3568 (N_3568,N_3421,N_3472);
and U3569 (N_3569,N_3463,N_3268);
or U3570 (N_3570,N_3427,N_3335);
nor U3571 (N_3571,N_3283,N_3323);
and U3572 (N_3572,N_3412,N_3350);
nand U3573 (N_3573,N_3339,N_3404);
nand U3574 (N_3574,N_3464,N_3470);
xnor U3575 (N_3575,N_3295,N_3449);
and U3576 (N_3576,N_3347,N_3378);
nor U3577 (N_3577,N_3290,N_3317);
nor U3578 (N_3578,N_3384,N_3313);
xor U3579 (N_3579,N_3370,N_3425);
and U3580 (N_3580,N_3447,N_3451);
nor U3581 (N_3581,N_3397,N_3437);
or U3582 (N_3582,N_3416,N_3379);
nand U3583 (N_3583,N_3439,N_3428);
xnor U3584 (N_3584,N_3394,N_3333);
and U3585 (N_3585,N_3314,N_3398);
and U3586 (N_3586,N_3374,N_3279);
nand U3587 (N_3587,N_3315,N_3406);
nor U3588 (N_3588,N_3461,N_3371);
nor U3589 (N_3589,N_3486,N_3343);
or U3590 (N_3590,N_3491,N_3402);
nand U3591 (N_3591,N_3310,N_3458);
nor U3592 (N_3592,N_3393,N_3413);
or U3593 (N_3593,N_3389,N_3377);
nand U3594 (N_3594,N_3366,N_3405);
xor U3595 (N_3595,N_3298,N_3250);
nor U3596 (N_3596,N_3352,N_3450);
and U3597 (N_3597,N_3388,N_3260);
or U3598 (N_3598,N_3254,N_3477);
nand U3599 (N_3599,N_3440,N_3433);
nor U3600 (N_3600,N_3331,N_3300);
nand U3601 (N_3601,N_3431,N_3420);
nand U3602 (N_3602,N_3481,N_3369);
and U3603 (N_3603,N_3487,N_3395);
nand U3604 (N_3604,N_3365,N_3448);
nor U3605 (N_3605,N_3373,N_3364);
and U3606 (N_3606,N_3309,N_3430);
and U3607 (N_3607,N_3316,N_3296);
and U3608 (N_3608,N_3410,N_3462);
nand U3609 (N_3609,N_3453,N_3252);
and U3610 (N_3610,N_3356,N_3344);
nand U3611 (N_3611,N_3307,N_3325);
xnor U3612 (N_3612,N_3414,N_3452);
nor U3613 (N_3613,N_3408,N_3321);
nand U3614 (N_3614,N_3401,N_3432);
and U3615 (N_3615,N_3266,N_3387);
nand U3616 (N_3616,N_3467,N_3257);
and U3617 (N_3617,N_3306,N_3368);
and U3618 (N_3618,N_3285,N_3489);
nor U3619 (N_3619,N_3403,N_3396);
xnor U3620 (N_3620,N_3328,N_3434);
and U3621 (N_3621,N_3297,N_3259);
xnor U3622 (N_3622,N_3337,N_3351);
nor U3623 (N_3623,N_3275,N_3375);
and U3624 (N_3624,N_3330,N_3269);
nand U3625 (N_3625,N_3486,N_3410);
nor U3626 (N_3626,N_3277,N_3436);
nand U3627 (N_3627,N_3275,N_3378);
and U3628 (N_3628,N_3313,N_3431);
nor U3629 (N_3629,N_3446,N_3347);
nand U3630 (N_3630,N_3272,N_3469);
nor U3631 (N_3631,N_3474,N_3351);
or U3632 (N_3632,N_3345,N_3305);
nor U3633 (N_3633,N_3308,N_3304);
and U3634 (N_3634,N_3413,N_3302);
or U3635 (N_3635,N_3417,N_3428);
nor U3636 (N_3636,N_3407,N_3317);
or U3637 (N_3637,N_3262,N_3260);
nor U3638 (N_3638,N_3277,N_3305);
or U3639 (N_3639,N_3379,N_3274);
nor U3640 (N_3640,N_3384,N_3482);
or U3641 (N_3641,N_3373,N_3385);
or U3642 (N_3642,N_3350,N_3421);
nand U3643 (N_3643,N_3443,N_3392);
or U3644 (N_3644,N_3479,N_3329);
xnor U3645 (N_3645,N_3387,N_3362);
nand U3646 (N_3646,N_3402,N_3440);
and U3647 (N_3647,N_3312,N_3493);
nand U3648 (N_3648,N_3336,N_3275);
and U3649 (N_3649,N_3352,N_3418);
and U3650 (N_3650,N_3483,N_3388);
or U3651 (N_3651,N_3489,N_3470);
and U3652 (N_3652,N_3445,N_3402);
and U3653 (N_3653,N_3430,N_3252);
nor U3654 (N_3654,N_3259,N_3464);
or U3655 (N_3655,N_3438,N_3366);
nor U3656 (N_3656,N_3443,N_3315);
and U3657 (N_3657,N_3454,N_3310);
nand U3658 (N_3658,N_3306,N_3461);
xor U3659 (N_3659,N_3491,N_3256);
nor U3660 (N_3660,N_3461,N_3430);
and U3661 (N_3661,N_3474,N_3401);
nand U3662 (N_3662,N_3428,N_3320);
nand U3663 (N_3663,N_3449,N_3306);
nor U3664 (N_3664,N_3299,N_3495);
nand U3665 (N_3665,N_3483,N_3279);
and U3666 (N_3666,N_3382,N_3261);
nor U3667 (N_3667,N_3260,N_3335);
or U3668 (N_3668,N_3305,N_3359);
and U3669 (N_3669,N_3415,N_3492);
xnor U3670 (N_3670,N_3295,N_3383);
xor U3671 (N_3671,N_3268,N_3468);
and U3672 (N_3672,N_3459,N_3309);
or U3673 (N_3673,N_3435,N_3472);
xnor U3674 (N_3674,N_3425,N_3311);
nor U3675 (N_3675,N_3324,N_3472);
and U3676 (N_3676,N_3279,N_3390);
or U3677 (N_3677,N_3291,N_3341);
nand U3678 (N_3678,N_3297,N_3470);
or U3679 (N_3679,N_3485,N_3343);
or U3680 (N_3680,N_3378,N_3456);
or U3681 (N_3681,N_3329,N_3291);
nand U3682 (N_3682,N_3264,N_3311);
nor U3683 (N_3683,N_3334,N_3366);
or U3684 (N_3684,N_3396,N_3336);
and U3685 (N_3685,N_3416,N_3452);
xor U3686 (N_3686,N_3353,N_3350);
nand U3687 (N_3687,N_3281,N_3328);
or U3688 (N_3688,N_3315,N_3327);
nor U3689 (N_3689,N_3406,N_3492);
nor U3690 (N_3690,N_3334,N_3466);
nor U3691 (N_3691,N_3327,N_3360);
and U3692 (N_3692,N_3470,N_3394);
xor U3693 (N_3693,N_3332,N_3320);
nand U3694 (N_3694,N_3397,N_3337);
and U3695 (N_3695,N_3403,N_3315);
nor U3696 (N_3696,N_3499,N_3410);
and U3697 (N_3697,N_3295,N_3279);
or U3698 (N_3698,N_3293,N_3291);
nor U3699 (N_3699,N_3494,N_3360);
and U3700 (N_3700,N_3487,N_3276);
or U3701 (N_3701,N_3324,N_3391);
nand U3702 (N_3702,N_3484,N_3468);
xor U3703 (N_3703,N_3456,N_3377);
nand U3704 (N_3704,N_3330,N_3439);
nor U3705 (N_3705,N_3275,N_3497);
nor U3706 (N_3706,N_3319,N_3317);
or U3707 (N_3707,N_3251,N_3294);
nand U3708 (N_3708,N_3395,N_3331);
or U3709 (N_3709,N_3337,N_3383);
nor U3710 (N_3710,N_3405,N_3327);
and U3711 (N_3711,N_3389,N_3294);
nand U3712 (N_3712,N_3373,N_3415);
or U3713 (N_3713,N_3267,N_3376);
or U3714 (N_3714,N_3374,N_3405);
nor U3715 (N_3715,N_3352,N_3471);
nor U3716 (N_3716,N_3437,N_3392);
xor U3717 (N_3717,N_3430,N_3254);
xor U3718 (N_3718,N_3275,N_3433);
xnor U3719 (N_3719,N_3414,N_3392);
or U3720 (N_3720,N_3368,N_3415);
xor U3721 (N_3721,N_3495,N_3441);
nor U3722 (N_3722,N_3307,N_3293);
nor U3723 (N_3723,N_3383,N_3429);
nand U3724 (N_3724,N_3260,N_3281);
xnor U3725 (N_3725,N_3419,N_3372);
nor U3726 (N_3726,N_3474,N_3371);
and U3727 (N_3727,N_3279,N_3260);
nor U3728 (N_3728,N_3261,N_3427);
and U3729 (N_3729,N_3320,N_3250);
nor U3730 (N_3730,N_3477,N_3318);
nand U3731 (N_3731,N_3375,N_3338);
and U3732 (N_3732,N_3385,N_3451);
xor U3733 (N_3733,N_3402,N_3371);
and U3734 (N_3734,N_3278,N_3320);
or U3735 (N_3735,N_3471,N_3378);
and U3736 (N_3736,N_3489,N_3344);
or U3737 (N_3737,N_3368,N_3353);
xnor U3738 (N_3738,N_3422,N_3288);
nand U3739 (N_3739,N_3379,N_3254);
and U3740 (N_3740,N_3305,N_3266);
or U3741 (N_3741,N_3447,N_3365);
xnor U3742 (N_3742,N_3485,N_3428);
xnor U3743 (N_3743,N_3367,N_3481);
and U3744 (N_3744,N_3433,N_3301);
and U3745 (N_3745,N_3325,N_3390);
or U3746 (N_3746,N_3289,N_3304);
xor U3747 (N_3747,N_3438,N_3405);
nand U3748 (N_3748,N_3440,N_3404);
nor U3749 (N_3749,N_3443,N_3395);
or U3750 (N_3750,N_3599,N_3651);
or U3751 (N_3751,N_3719,N_3594);
xor U3752 (N_3752,N_3665,N_3514);
or U3753 (N_3753,N_3642,N_3525);
nor U3754 (N_3754,N_3664,N_3583);
xor U3755 (N_3755,N_3663,N_3632);
nor U3756 (N_3756,N_3713,N_3575);
nor U3757 (N_3757,N_3524,N_3513);
and U3758 (N_3758,N_3537,N_3626);
nor U3759 (N_3759,N_3544,N_3704);
and U3760 (N_3760,N_3732,N_3647);
xnor U3761 (N_3761,N_3686,N_3667);
nand U3762 (N_3762,N_3543,N_3641);
nor U3763 (N_3763,N_3697,N_3679);
xnor U3764 (N_3764,N_3576,N_3579);
nand U3765 (N_3765,N_3563,N_3553);
or U3766 (N_3766,N_3520,N_3573);
nand U3767 (N_3767,N_3593,N_3526);
or U3768 (N_3768,N_3712,N_3620);
xor U3769 (N_3769,N_3581,N_3650);
nand U3770 (N_3770,N_3703,N_3658);
or U3771 (N_3771,N_3506,N_3748);
xor U3772 (N_3772,N_3574,N_3603);
xor U3773 (N_3773,N_3547,N_3677);
nand U3774 (N_3774,N_3639,N_3534);
and U3775 (N_3775,N_3622,N_3716);
xor U3776 (N_3776,N_3671,N_3736);
and U3777 (N_3777,N_3542,N_3555);
nor U3778 (N_3778,N_3529,N_3681);
and U3779 (N_3779,N_3597,N_3619);
or U3780 (N_3780,N_3675,N_3731);
and U3781 (N_3781,N_3569,N_3557);
nor U3782 (N_3782,N_3530,N_3721);
nand U3783 (N_3783,N_3680,N_3505);
xor U3784 (N_3784,N_3741,N_3598);
and U3785 (N_3785,N_3552,N_3540);
nor U3786 (N_3786,N_3685,N_3501);
nor U3787 (N_3787,N_3698,N_3657);
or U3788 (N_3788,N_3687,N_3701);
nor U3789 (N_3789,N_3739,N_3695);
or U3790 (N_3790,N_3536,N_3635);
and U3791 (N_3791,N_3609,N_3572);
nand U3792 (N_3792,N_3668,N_3522);
and U3793 (N_3793,N_3561,N_3566);
and U3794 (N_3794,N_3571,N_3627);
and U3795 (N_3795,N_3517,N_3528);
nand U3796 (N_3796,N_3538,N_3611);
nor U3797 (N_3797,N_3694,N_3692);
nand U3798 (N_3798,N_3634,N_3511);
xor U3799 (N_3799,N_3735,N_3503);
and U3800 (N_3800,N_3586,N_3662);
xnor U3801 (N_3801,N_3666,N_3710);
and U3802 (N_3802,N_3560,N_3744);
or U3803 (N_3803,N_3727,N_3684);
nand U3804 (N_3804,N_3607,N_3726);
xor U3805 (N_3805,N_3605,N_3643);
nand U3806 (N_3806,N_3648,N_3523);
and U3807 (N_3807,N_3518,N_3624);
and U3808 (N_3808,N_3653,N_3612);
nand U3809 (N_3809,N_3585,N_3625);
xnor U3810 (N_3810,N_3516,N_3590);
or U3811 (N_3811,N_3584,N_3688);
xor U3812 (N_3812,N_3740,N_3717);
xnor U3813 (N_3813,N_3746,N_3559);
nor U3814 (N_3814,N_3733,N_3527);
or U3815 (N_3815,N_3628,N_3546);
or U3816 (N_3816,N_3661,N_3682);
xor U3817 (N_3817,N_3580,N_3747);
xnor U3818 (N_3818,N_3720,N_3582);
nand U3819 (N_3819,N_3532,N_3570);
and U3820 (N_3820,N_3678,N_3655);
and U3821 (N_3821,N_3595,N_3631);
xnor U3822 (N_3822,N_3539,N_3551);
and U3823 (N_3823,N_3564,N_3743);
and U3824 (N_3824,N_3649,N_3610);
nor U3825 (N_3825,N_3588,N_3707);
or U3826 (N_3826,N_3672,N_3587);
nor U3827 (N_3827,N_3629,N_3693);
or U3828 (N_3828,N_3640,N_3531);
and U3829 (N_3829,N_3745,N_3509);
nand U3830 (N_3830,N_3615,N_3706);
and U3831 (N_3831,N_3708,N_3601);
nand U3832 (N_3832,N_3645,N_3633);
nand U3833 (N_3833,N_3659,N_3623);
or U3834 (N_3834,N_3734,N_3515);
nor U3835 (N_3835,N_3535,N_3674);
and U3836 (N_3836,N_3567,N_3652);
and U3837 (N_3837,N_3702,N_3714);
nand U3838 (N_3838,N_3504,N_3608);
nand U3839 (N_3839,N_3521,N_3502);
and U3840 (N_3840,N_3636,N_3554);
nand U3841 (N_3841,N_3646,N_3742);
and U3842 (N_3842,N_3644,N_3690);
xnor U3843 (N_3843,N_3617,N_3519);
xor U3844 (N_3844,N_3700,N_3638);
and U3845 (N_3845,N_3656,N_3669);
nor U3846 (N_3846,N_3550,N_3562);
nand U3847 (N_3847,N_3725,N_3556);
or U3848 (N_3848,N_3549,N_3614);
or U3849 (N_3849,N_3616,N_3705);
xor U3850 (N_3850,N_3510,N_3600);
or U3851 (N_3851,N_3738,N_3606);
and U3852 (N_3852,N_3724,N_3711);
nor U3853 (N_3853,N_3660,N_3618);
nand U3854 (N_3854,N_3715,N_3613);
and U3855 (N_3855,N_3548,N_3637);
or U3856 (N_3856,N_3699,N_3749);
nand U3857 (N_3857,N_3589,N_3500);
or U3858 (N_3858,N_3737,N_3689);
and U3859 (N_3859,N_3591,N_3558);
nor U3860 (N_3860,N_3728,N_3691);
nand U3861 (N_3861,N_3729,N_3621);
or U3862 (N_3862,N_3683,N_3604);
or U3863 (N_3863,N_3512,N_3654);
nor U3864 (N_3864,N_3696,N_3533);
nor U3865 (N_3865,N_3507,N_3541);
xor U3866 (N_3866,N_3676,N_3718);
xor U3867 (N_3867,N_3723,N_3592);
or U3868 (N_3868,N_3568,N_3673);
and U3869 (N_3869,N_3596,N_3565);
xor U3870 (N_3870,N_3670,N_3730);
nor U3871 (N_3871,N_3545,N_3722);
xnor U3872 (N_3872,N_3602,N_3508);
or U3873 (N_3873,N_3577,N_3578);
nand U3874 (N_3874,N_3630,N_3709);
nand U3875 (N_3875,N_3705,N_3559);
xnor U3876 (N_3876,N_3506,N_3708);
nor U3877 (N_3877,N_3592,N_3695);
xor U3878 (N_3878,N_3618,N_3558);
xor U3879 (N_3879,N_3526,N_3674);
xnor U3880 (N_3880,N_3612,N_3608);
nor U3881 (N_3881,N_3524,N_3503);
and U3882 (N_3882,N_3628,N_3504);
xnor U3883 (N_3883,N_3638,N_3709);
or U3884 (N_3884,N_3595,N_3612);
nor U3885 (N_3885,N_3572,N_3539);
nor U3886 (N_3886,N_3519,N_3731);
nand U3887 (N_3887,N_3717,N_3570);
and U3888 (N_3888,N_3511,N_3686);
and U3889 (N_3889,N_3585,N_3571);
xor U3890 (N_3890,N_3534,N_3739);
or U3891 (N_3891,N_3505,N_3634);
or U3892 (N_3892,N_3616,N_3541);
nand U3893 (N_3893,N_3677,N_3601);
xor U3894 (N_3894,N_3507,N_3598);
xor U3895 (N_3895,N_3695,N_3691);
or U3896 (N_3896,N_3506,N_3611);
nand U3897 (N_3897,N_3714,N_3537);
nor U3898 (N_3898,N_3634,N_3522);
xor U3899 (N_3899,N_3708,N_3598);
nor U3900 (N_3900,N_3667,N_3557);
nand U3901 (N_3901,N_3672,N_3671);
or U3902 (N_3902,N_3712,N_3540);
or U3903 (N_3903,N_3688,N_3697);
or U3904 (N_3904,N_3734,N_3748);
nand U3905 (N_3905,N_3608,N_3726);
nor U3906 (N_3906,N_3749,N_3671);
xnor U3907 (N_3907,N_3660,N_3743);
nand U3908 (N_3908,N_3561,N_3505);
and U3909 (N_3909,N_3575,N_3730);
or U3910 (N_3910,N_3503,N_3528);
nor U3911 (N_3911,N_3569,N_3552);
xor U3912 (N_3912,N_3631,N_3695);
and U3913 (N_3913,N_3690,N_3692);
nand U3914 (N_3914,N_3579,N_3732);
xnor U3915 (N_3915,N_3578,N_3619);
nor U3916 (N_3916,N_3520,N_3682);
xnor U3917 (N_3917,N_3689,N_3565);
nor U3918 (N_3918,N_3624,N_3629);
nor U3919 (N_3919,N_3601,N_3520);
nand U3920 (N_3920,N_3668,N_3500);
or U3921 (N_3921,N_3514,N_3660);
nand U3922 (N_3922,N_3509,N_3521);
xnor U3923 (N_3923,N_3545,N_3513);
or U3924 (N_3924,N_3655,N_3690);
nor U3925 (N_3925,N_3534,N_3689);
nand U3926 (N_3926,N_3594,N_3569);
nand U3927 (N_3927,N_3691,N_3738);
and U3928 (N_3928,N_3538,N_3726);
nand U3929 (N_3929,N_3539,N_3540);
and U3930 (N_3930,N_3745,N_3713);
and U3931 (N_3931,N_3734,N_3575);
nand U3932 (N_3932,N_3667,N_3666);
and U3933 (N_3933,N_3556,N_3692);
xnor U3934 (N_3934,N_3611,N_3730);
nor U3935 (N_3935,N_3643,N_3744);
nand U3936 (N_3936,N_3747,N_3501);
nor U3937 (N_3937,N_3545,N_3747);
nor U3938 (N_3938,N_3547,N_3659);
and U3939 (N_3939,N_3546,N_3660);
nand U3940 (N_3940,N_3650,N_3634);
nand U3941 (N_3941,N_3511,N_3609);
nand U3942 (N_3942,N_3672,N_3691);
nor U3943 (N_3943,N_3695,N_3669);
or U3944 (N_3944,N_3555,N_3554);
and U3945 (N_3945,N_3617,N_3578);
xnor U3946 (N_3946,N_3700,N_3749);
xor U3947 (N_3947,N_3636,N_3628);
xor U3948 (N_3948,N_3566,N_3670);
or U3949 (N_3949,N_3635,N_3522);
or U3950 (N_3950,N_3721,N_3593);
nor U3951 (N_3951,N_3590,N_3729);
nor U3952 (N_3952,N_3501,N_3690);
nor U3953 (N_3953,N_3616,N_3671);
nand U3954 (N_3954,N_3684,N_3656);
and U3955 (N_3955,N_3527,N_3637);
or U3956 (N_3956,N_3505,N_3641);
and U3957 (N_3957,N_3576,N_3637);
nand U3958 (N_3958,N_3602,N_3516);
nand U3959 (N_3959,N_3577,N_3740);
nand U3960 (N_3960,N_3564,N_3532);
or U3961 (N_3961,N_3528,N_3730);
nor U3962 (N_3962,N_3634,N_3604);
nor U3963 (N_3963,N_3529,N_3652);
nor U3964 (N_3964,N_3703,N_3635);
nand U3965 (N_3965,N_3568,N_3589);
and U3966 (N_3966,N_3709,N_3649);
xnor U3967 (N_3967,N_3573,N_3680);
and U3968 (N_3968,N_3540,N_3710);
nand U3969 (N_3969,N_3579,N_3608);
or U3970 (N_3970,N_3737,N_3566);
or U3971 (N_3971,N_3585,N_3570);
and U3972 (N_3972,N_3635,N_3509);
xnor U3973 (N_3973,N_3664,N_3504);
or U3974 (N_3974,N_3572,N_3620);
xor U3975 (N_3975,N_3705,N_3658);
and U3976 (N_3976,N_3572,N_3509);
nand U3977 (N_3977,N_3631,N_3586);
nor U3978 (N_3978,N_3594,N_3628);
or U3979 (N_3979,N_3535,N_3582);
xor U3980 (N_3980,N_3562,N_3746);
nor U3981 (N_3981,N_3610,N_3624);
nand U3982 (N_3982,N_3532,N_3585);
nor U3983 (N_3983,N_3723,N_3545);
and U3984 (N_3984,N_3522,N_3610);
or U3985 (N_3985,N_3547,N_3678);
and U3986 (N_3986,N_3682,N_3532);
and U3987 (N_3987,N_3724,N_3544);
nor U3988 (N_3988,N_3733,N_3591);
nand U3989 (N_3989,N_3573,N_3635);
nand U3990 (N_3990,N_3673,N_3713);
nor U3991 (N_3991,N_3656,N_3640);
and U3992 (N_3992,N_3620,N_3566);
nand U3993 (N_3993,N_3734,N_3724);
nand U3994 (N_3994,N_3742,N_3565);
and U3995 (N_3995,N_3616,N_3531);
or U3996 (N_3996,N_3707,N_3606);
or U3997 (N_3997,N_3515,N_3657);
nor U3998 (N_3998,N_3736,N_3565);
xor U3999 (N_3999,N_3647,N_3684);
or U4000 (N_4000,N_3889,N_3891);
nand U4001 (N_4001,N_3774,N_3871);
and U4002 (N_4002,N_3910,N_3881);
nand U4003 (N_4003,N_3857,N_3811);
nand U4004 (N_4004,N_3938,N_3753);
nand U4005 (N_4005,N_3901,N_3866);
or U4006 (N_4006,N_3752,N_3778);
xnor U4007 (N_4007,N_3942,N_3907);
nor U4008 (N_4008,N_3994,N_3996);
xor U4009 (N_4009,N_3895,N_3872);
xnor U4010 (N_4010,N_3763,N_3972);
or U4011 (N_4011,N_3928,N_3768);
xor U4012 (N_4012,N_3885,N_3973);
xor U4013 (N_4013,N_3977,N_3944);
and U4014 (N_4014,N_3905,N_3770);
xnor U4015 (N_4015,N_3991,N_3842);
and U4016 (N_4016,N_3818,N_3771);
or U4017 (N_4017,N_3927,N_3933);
or U4018 (N_4018,N_3865,N_3940);
nand U4019 (N_4019,N_3984,N_3869);
or U4020 (N_4020,N_3757,N_3961);
and U4021 (N_4021,N_3837,N_3952);
xor U4022 (N_4022,N_3975,N_3765);
and U4023 (N_4023,N_3815,N_3788);
and U4024 (N_4024,N_3833,N_3810);
or U4025 (N_4025,N_3921,N_3935);
nor U4026 (N_4026,N_3999,N_3997);
nand U4027 (N_4027,N_3876,N_3971);
xor U4028 (N_4028,N_3970,N_3819);
nor U4029 (N_4029,N_3978,N_3784);
nand U4030 (N_4030,N_3820,N_3949);
nor U4031 (N_4031,N_3794,N_3924);
xnor U4032 (N_4032,N_3781,N_3754);
and U4033 (N_4033,N_3838,N_3930);
or U4034 (N_4034,N_3858,N_3822);
xor U4035 (N_4035,N_3848,N_3902);
and U4036 (N_4036,N_3845,N_3878);
and U4037 (N_4037,N_3808,N_3824);
and U4038 (N_4038,N_3817,N_3843);
and U4039 (N_4039,N_3862,N_3900);
xnor U4040 (N_4040,N_3948,N_3873);
nand U4041 (N_4041,N_3884,N_3890);
or U4042 (N_4042,N_3931,N_3879);
xor U4043 (N_4043,N_3989,N_3875);
nor U4044 (N_4044,N_3797,N_3751);
or U4045 (N_4045,N_3886,N_3981);
and U4046 (N_4046,N_3919,N_3982);
nand U4047 (N_4047,N_3898,N_3941);
xor U4048 (N_4048,N_3789,N_3897);
and U4049 (N_4049,N_3914,N_3995);
nand U4050 (N_4050,N_3954,N_3979);
or U4051 (N_4051,N_3888,N_3962);
or U4052 (N_4052,N_3790,N_3780);
or U4053 (N_4053,N_3868,N_3782);
or U4054 (N_4054,N_3936,N_3802);
nor U4055 (N_4055,N_3801,N_3805);
or U4056 (N_4056,N_3947,N_3976);
xor U4057 (N_4057,N_3806,N_3849);
nand U4058 (N_4058,N_3983,N_3773);
xor U4059 (N_4059,N_3816,N_3769);
xor U4060 (N_4060,N_3943,N_3785);
nand U4061 (N_4061,N_3985,N_3883);
xnor U4062 (N_4062,N_3899,N_3882);
xor U4063 (N_4063,N_3854,N_3795);
xnor U4064 (N_4064,N_3762,N_3964);
nor U4065 (N_4065,N_3829,N_3809);
nor U4066 (N_4066,N_3755,N_3831);
or U4067 (N_4067,N_3756,N_3870);
xor U4068 (N_4068,N_3787,N_3830);
nand U4069 (N_4069,N_3836,N_3955);
nand U4070 (N_4070,N_3796,N_3793);
and U4071 (N_4071,N_3950,N_3798);
nor U4072 (N_4072,N_3750,N_3917);
or U4073 (N_4073,N_3929,N_3926);
and U4074 (N_4074,N_3987,N_3764);
nand U4075 (N_4075,N_3791,N_3814);
xnor U4076 (N_4076,N_3968,N_3834);
or U4077 (N_4077,N_3759,N_3963);
xor U4078 (N_4078,N_3918,N_3939);
nand U4079 (N_4079,N_3913,N_3877);
or U4080 (N_4080,N_3908,N_3880);
or U4081 (N_4081,N_3894,N_3760);
nand U4082 (N_4082,N_3916,N_3826);
or U4083 (N_4083,N_3967,N_3958);
nand U4084 (N_4084,N_3915,N_3909);
and U4085 (N_4085,N_3786,N_3853);
nand U4086 (N_4086,N_3758,N_3861);
nand U4087 (N_4087,N_3840,N_3799);
and U4088 (N_4088,N_3772,N_3923);
nor U4089 (N_4089,N_3953,N_3951);
and U4090 (N_4090,N_3912,N_3783);
nor U4091 (N_4091,N_3904,N_3767);
nand U4092 (N_4092,N_3803,N_3850);
and U4093 (N_4093,N_3980,N_3969);
nand U4094 (N_4094,N_3874,N_3864);
xor U4095 (N_4095,N_3993,N_3920);
nor U4096 (N_4096,N_3859,N_3925);
nand U4097 (N_4097,N_3932,N_3855);
nand U4098 (N_4098,N_3807,N_3804);
nand U4099 (N_4099,N_3965,N_3896);
nand U4100 (N_4100,N_3800,N_3906);
or U4101 (N_4101,N_3893,N_3986);
xnor U4102 (N_4102,N_3825,N_3863);
or U4103 (N_4103,N_3922,N_3974);
xor U4104 (N_4104,N_3766,N_3776);
or U4105 (N_4105,N_3988,N_3775);
or U4106 (N_4106,N_3911,N_3846);
nand U4107 (N_4107,N_3957,N_3992);
and U4108 (N_4108,N_3990,N_3827);
nor U4109 (N_4109,N_3856,N_3844);
nor U4110 (N_4110,N_3937,N_3934);
nand U4111 (N_4111,N_3839,N_3852);
and U4112 (N_4112,N_3832,N_3847);
nand U4113 (N_4113,N_3966,N_3821);
nor U4114 (N_4114,N_3813,N_3867);
xor U4115 (N_4115,N_3779,N_3956);
nor U4116 (N_4116,N_3792,N_3892);
and U4117 (N_4117,N_3903,N_3761);
and U4118 (N_4118,N_3887,N_3959);
and U4119 (N_4119,N_3945,N_3823);
nor U4120 (N_4120,N_3960,N_3946);
and U4121 (N_4121,N_3851,N_3777);
nor U4122 (N_4122,N_3998,N_3841);
and U4123 (N_4123,N_3828,N_3835);
xor U4124 (N_4124,N_3812,N_3860);
and U4125 (N_4125,N_3764,N_3925);
xnor U4126 (N_4126,N_3807,N_3866);
and U4127 (N_4127,N_3928,N_3885);
xnor U4128 (N_4128,N_3924,N_3800);
xor U4129 (N_4129,N_3881,N_3888);
and U4130 (N_4130,N_3922,N_3806);
and U4131 (N_4131,N_3927,N_3788);
or U4132 (N_4132,N_3775,N_3768);
nor U4133 (N_4133,N_3825,N_3793);
and U4134 (N_4134,N_3931,N_3994);
and U4135 (N_4135,N_3780,N_3777);
and U4136 (N_4136,N_3931,N_3800);
xnor U4137 (N_4137,N_3769,N_3794);
nand U4138 (N_4138,N_3976,N_3879);
or U4139 (N_4139,N_3991,N_3916);
nand U4140 (N_4140,N_3975,N_3973);
nand U4141 (N_4141,N_3924,N_3927);
and U4142 (N_4142,N_3833,N_3889);
and U4143 (N_4143,N_3962,N_3872);
and U4144 (N_4144,N_3915,N_3867);
xor U4145 (N_4145,N_3894,N_3838);
xor U4146 (N_4146,N_3823,N_3908);
or U4147 (N_4147,N_3761,N_3782);
or U4148 (N_4148,N_3843,N_3826);
xor U4149 (N_4149,N_3971,N_3896);
nand U4150 (N_4150,N_3823,N_3801);
or U4151 (N_4151,N_3844,N_3950);
xor U4152 (N_4152,N_3861,N_3768);
or U4153 (N_4153,N_3853,N_3773);
xor U4154 (N_4154,N_3882,N_3839);
or U4155 (N_4155,N_3764,N_3873);
xnor U4156 (N_4156,N_3945,N_3970);
nand U4157 (N_4157,N_3947,N_3965);
nand U4158 (N_4158,N_3986,N_3926);
and U4159 (N_4159,N_3877,N_3791);
or U4160 (N_4160,N_3769,N_3791);
nand U4161 (N_4161,N_3875,N_3977);
xnor U4162 (N_4162,N_3798,N_3832);
xnor U4163 (N_4163,N_3873,N_3840);
nand U4164 (N_4164,N_3792,N_3761);
xor U4165 (N_4165,N_3868,N_3952);
xor U4166 (N_4166,N_3852,N_3959);
nand U4167 (N_4167,N_3835,N_3956);
and U4168 (N_4168,N_3790,N_3846);
or U4169 (N_4169,N_3955,N_3898);
and U4170 (N_4170,N_3854,N_3955);
xnor U4171 (N_4171,N_3799,N_3864);
nor U4172 (N_4172,N_3932,N_3965);
nand U4173 (N_4173,N_3868,N_3873);
xor U4174 (N_4174,N_3920,N_3757);
and U4175 (N_4175,N_3992,N_3990);
and U4176 (N_4176,N_3998,N_3967);
nor U4177 (N_4177,N_3958,N_3833);
and U4178 (N_4178,N_3833,N_3799);
nor U4179 (N_4179,N_3847,N_3984);
nand U4180 (N_4180,N_3922,N_3824);
nand U4181 (N_4181,N_3989,N_3945);
xnor U4182 (N_4182,N_3773,N_3798);
or U4183 (N_4183,N_3925,N_3906);
and U4184 (N_4184,N_3959,N_3904);
and U4185 (N_4185,N_3994,N_3948);
nor U4186 (N_4186,N_3831,N_3924);
and U4187 (N_4187,N_3778,N_3773);
nor U4188 (N_4188,N_3837,N_3947);
and U4189 (N_4189,N_3943,N_3851);
nor U4190 (N_4190,N_3832,N_3949);
and U4191 (N_4191,N_3810,N_3951);
or U4192 (N_4192,N_3965,N_3956);
xor U4193 (N_4193,N_3982,N_3819);
and U4194 (N_4194,N_3935,N_3837);
nand U4195 (N_4195,N_3899,N_3868);
nor U4196 (N_4196,N_3845,N_3761);
nor U4197 (N_4197,N_3752,N_3779);
nand U4198 (N_4198,N_3946,N_3935);
xnor U4199 (N_4199,N_3875,N_3953);
nor U4200 (N_4200,N_3998,N_3758);
and U4201 (N_4201,N_3856,N_3754);
and U4202 (N_4202,N_3833,N_3985);
or U4203 (N_4203,N_3987,N_3949);
xnor U4204 (N_4204,N_3809,N_3968);
xor U4205 (N_4205,N_3800,N_3876);
and U4206 (N_4206,N_3992,N_3754);
nor U4207 (N_4207,N_3924,N_3863);
xnor U4208 (N_4208,N_3855,N_3974);
nand U4209 (N_4209,N_3976,N_3839);
and U4210 (N_4210,N_3829,N_3962);
nor U4211 (N_4211,N_3858,N_3770);
and U4212 (N_4212,N_3767,N_3801);
and U4213 (N_4213,N_3964,N_3899);
and U4214 (N_4214,N_3957,N_3816);
or U4215 (N_4215,N_3763,N_3886);
or U4216 (N_4216,N_3888,N_3912);
or U4217 (N_4217,N_3789,N_3751);
xnor U4218 (N_4218,N_3811,N_3834);
or U4219 (N_4219,N_3798,N_3973);
xor U4220 (N_4220,N_3959,N_3753);
or U4221 (N_4221,N_3923,N_3959);
nand U4222 (N_4222,N_3955,N_3828);
or U4223 (N_4223,N_3827,N_3879);
xnor U4224 (N_4224,N_3899,N_3953);
nor U4225 (N_4225,N_3794,N_3932);
xnor U4226 (N_4226,N_3956,N_3930);
and U4227 (N_4227,N_3892,N_3843);
or U4228 (N_4228,N_3954,N_3991);
nor U4229 (N_4229,N_3789,N_3952);
and U4230 (N_4230,N_3895,N_3862);
nand U4231 (N_4231,N_3824,N_3970);
xor U4232 (N_4232,N_3785,N_3799);
xnor U4233 (N_4233,N_3833,N_3821);
nand U4234 (N_4234,N_3940,N_3989);
xnor U4235 (N_4235,N_3978,N_3898);
nand U4236 (N_4236,N_3996,N_3789);
xor U4237 (N_4237,N_3827,N_3818);
nor U4238 (N_4238,N_3764,N_3813);
or U4239 (N_4239,N_3836,N_3834);
and U4240 (N_4240,N_3761,N_3878);
or U4241 (N_4241,N_3877,N_3770);
xnor U4242 (N_4242,N_3953,N_3946);
nand U4243 (N_4243,N_3913,N_3818);
and U4244 (N_4244,N_3752,N_3965);
nor U4245 (N_4245,N_3813,N_3868);
xor U4246 (N_4246,N_3893,N_3995);
and U4247 (N_4247,N_3892,N_3751);
nor U4248 (N_4248,N_3864,N_3759);
xor U4249 (N_4249,N_3868,N_3771);
xor U4250 (N_4250,N_4087,N_4012);
and U4251 (N_4251,N_4144,N_4014);
nand U4252 (N_4252,N_4184,N_4004);
nor U4253 (N_4253,N_4108,N_4122);
or U4254 (N_4254,N_4165,N_4216);
or U4255 (N_4255,N_4082,N_4151);
nand U4256 (N_4256,N_4041,N_4158);
xnor U4257 (N_4257,N_4197,N_4136);
and U4258 (N_4258,N_4169,N_4243);
nor U4259 (N_4259,N_4021,N_4095);
nand U4260 (N_4260,N_4075,N_4077);
nand U4261 (N_4261,N_4118,N_4067);
and U4262 (N_4262,N_4036,N_4104);
or U4263 (N_4263,N_4061,N_4137);
nor U4264 (N_4264,N_4016,N_4195);
xor U4265 (N_4265,N_4126,N_4006);
nor U4266 (N_4266,N_4102,N_4248);
and U4267 (N_4267,N_4111,N_4143);
nor U4268 (N_4268,N_4022,N_4226);
or U4269 (N_4269,N_4062,N_4053);
and U4270 (N_4270,N_4218,N_4211);
nand U4271 (N_4271,N_4109,N_4249);
xor U4272 (N_4272,N_4009,N_4064);
xor U4273 (N_4273,N_4020,N_4119);
xor U4274 (N_4274,N_4127,N_4084);
xor U4275 (N_4275,N_4206,N_4121);
nor U4276 (N_4276,N_4069,N_4157);
xor U4277 (N_4277,N_4160,N_4170);
and U4278 (N_4278,N_4039,N_4140);
nor U4279 (N_4279,N_4124,N_4083);
or U4280 (N_4280,N_4046,N_4076);
nand U4281 (N_4281,N_4191,N_4026);
nor U4282 (N_4282,N_4107,N_4229);
or U4283 (N_4283,N_4223,N_4193);
nand U4284 (N_4284,N_4187,N_4204);
nand U4285 (N_4285,N_4128,N_4237);
nor U4286 (N_4286,N_4113,N_4150);
and U4287 (N_4287,N_4090,N_4043);
or U4288 (N_4288,N_4156,N_4220);
and U4289 (N_4289,N_4110,N_4068);
or U4290 (N_4290,N_4135,N_4142);
or U4291 (N_4291,N_4152,N_4228);
and U4292 (N_4292,N_4173,N_4018);
nand U4293 (N_4293,N_4080,N_4139);
nor U4294 (N_4294,N_4183,N_4202);
and U4295 (N_4295,N_4171,N_4079);
nand U4296 (N_4296,N_4063,N_4245);
nor U4297 (N_4297,N_4040,N_4133);
nand U4298 (N_4298,N_4167,N_4098);
nor U4299 (N_4299,N_4055,N_4032);
nand U4300 (N_4300,N_4148,N_4130);
or U4301 (N_4301,N_4225,N_4015);
nor U4302 (N_4302,N_4182,N_4112);
and U4303 (N_4303,N_4185,N_4045);
or U4304 (N_4304,N_4166,N_4089);
xor U4305 (N_4305,N_4134,N_4208);
xor U4306 (N_4306,N_4031,N_4232);
or U4307 (N_4307,N_4132,N_4037);
nand U4308 (N_4308,N_4099,N_4101);
xor U4309 (N_4309,N_4005,N_4123);
and U4310 (N_4310,N_4178,N_4050);
nand U4311 (N_4311,N_4141,N_4072);
nand U4312 (N_4312,N_4115,N_4227);
nor U4313 (N_4313,N_4242,N_4205);
xor U4314 (N_4314,N_4233,N_4239);
or U4315 (N_4315,N_4168,N_4159);
nor U4316 (N_4316,N_4081,N_4088);
nor U4317 (N_4317,N_4116,N_4114);
or U4318 (N_4318,N_4154,N_4172);
nand U4319 (N_4319,N_4125,N_4200);
nand U4320 (N_4320,N_4094,N_4246);
nor U4321 (N_4321,N_4213,N_4074);
and U4322 (N_4322,N_4092,N_4044);
nand U4323 (N_4323,N_4146,N_4049);
and U4324 (N_4324,N_4038,N_4238);
xnor U4325 (N_4325,N_4240,N_4207);
nand U4326 (N_4326,N_4052,N_4106);
or U4327 (N_4327,N_4027,N_4222);
nor U4328 (N_4328,N_4174,N_4058);
xor U4329 (N_4329,N_4096,N_4034);
or U4330 (N_4330,N_4085,N_4198);
nor U4331 (N_4331,N_4181,N_4059);
xnor U4332 (N_4332,N_4100,N_4175);
nor U4333 (N_4333,N_4007,N_4013);
or U4334 (N_4334,N_4186,N_4025);
xor U4335 (N_4335,N_4199,N_4149);
or U4336 (N_4336,N_4011,N_4047);
or U4337 (N_4337,N_4145,N_4057);
nand U4338 (N_4338,N_4093,N_4153);
and U4339 (N_4339,N_4086,N_4147);
and U4340 (N_4340,N_4023,N_4210);
xor U4341 (N_4341,N_4164,N_4241);
nand U4342 (N_4342,N_4078,N_4231);
nand U4343 (N_4343,N_4179,N_4017);
or U4344 (N_4344,N_4247,N_4196);
or U4345 (N_4345,N_4177,N_4201);
xnor U4346 (N_4346,N_4214,N_4176);
xnor U4347 (N_4347,N_4001,N_4235);
nand U4348 (N_4348,N_4070,N_4138);
and U4349 (N_4349,N_4097,N_4236);
nor U4350 (N_4350,N_4065,N_4071);
xor U4351 (N_4351,N_4054,N_4189);
xor U4352 (N_4352,N_4203,N_4073);
xnor U4353 (N_4353,N_4019,N_4209);
xor U4354 (N_4354,N_4131,N_4008);
and U4355 (N_4355,N_4221,N_4155);
nor U4356 (N_4356,N_4103,N_4192);
and U4357 (N_4357,N_4162,N_4180);
nor U4358 (N_4358,N_4215,N_4028);
nand U4359 (N_4359,N_4024,N_4033);
and U4360 (N_4360,N_4091,N_4230);
or U4361 (N_4361,N_4105,N_4003);
xor U4362 (N_4362,N_4035,N_4190);
and U4363 (N_4363,N_4120,N_4219);
and U4364 (N_4364,N_4029,N_4194);
and U4365 (N_4365,N_4129,N_4212);
or U4366 (N_4366,N_4161,N_4002);
and U4367 (N_4367,N_4048,N_4010);
nor U4368 (N_4368,N_4117,N_4188);
xor U4369 (N_4369,N_4163,N_4000);
nand U4370 (N_4370,N_4051,N_4056);
xnor U4371 (N_4371,N_4217,N_4030);
or U4372 (N_4372,N_4066,N_4244);
nor U4373 (N_4373,N_4060,N_4234);
xnor U4374 (N_4374,N_4042,N_4224);
xnor U4375 (N_4375,N_4019,N_4113);
nor U4376 (N_4376,N_4177,N_4226);
nand U4377 (N_4377,N_4089,N_4233);
nand U4378 (N_4378,N_4234,N_4135);
nand U4379 (N_4379,N_4003,N_4219);
nor U4380 (N_4380,N_4045,N_4084);
xnor U4381 (N_4381,N_4153,N_4132);
nand U4382 (N_4382,N_4083,N_4245);
xnor U4383 (N_4383,N_4240,N_4087);
and U4384 (N_4384,N_4058,N_4232);
nand U4385 (N_4385,N_4066,N_4216);
xor U4386 (N_4386,N_4097,N_4186);
or U4387 (N_4387,N_4141,N_4075);
and U4388 (N_4388,N_4173,N_4196);
xor U4389 (N_4389,N_4158,N_4162);
and U4390 (N_4390,N_4179,N_4110);
nand U4391 (N_4391,N_4064,N_4100);
nor U4392 (N_4392,N_4173,N_4123);
xnor U4393 (N_4393,N_4211,N_4008);
nor U4394 (N_4394,N_4222,N_4245);
nand U4395 (N_4395,N_4008,N_4011);
nand U4396 (N_4396,N_4174,N_4136);
and U4397 (N_4397,N_4161,N_4134);
nor U4398 (N_4398,N_4225,N_4012);
nand U4399 (N_4399,N_4039,N_4043);
or U4400 (N_4400,N_4229,N_4027);
and U4401 (N_4401,N_4211,N_4065);
or U4402 (N_4402,N_4153,N_4166);
xor U4403 (N_4403,N_4094,N_4201);
xor U4404 (N_4404,N_4222,N_4094);
or U4405 (N_4405,N_4040,N_4211);
nand U4406 (N_4406,N_4046,N_4090);
or U4407 (N_4407,N_4137,N_4155);
and U4408 (N_4408,N_4077,N_4162);
and U4409 (N_4409,N_4079,N_4133);
xor U4410 (N_4410,N_4002,N_4019);
nand U4411 (N_4411,N_4246,N_4140);
or U4412 (N_4412,N_4007,N_4056);
nand U4413 (N_4413,N_4246,N_4103);
xnor U4414 (N_4414,N_4139,N_4246);
nor U4415 (N_4415,N_4142,N_4015);
nand U4416 (N_4416,N_4010,N_4116);
nand U4417 (N_4417,N_4011,N_4048);
nor U4418 (N_4418,N_4111,N_4142);
nor U4419 (N_4419,N_4073,N_4138);
xnor U4420 (N_4420,N_4033,N_4083);
nand U4421 (N_4421,N_4203,N_4043);
nor U4422 (N_4422,N_4179,N_4139);
and U4423 (N_4423,N_4128,N_4062);
xnor U4424 (N_4424,N_4077,N_4148);
and U4425 (N_4425,N_4149,N_4013);
and U4426 (N_4426,N_4248,N_4207);
xnor U4427 (N_4427,N_4196,N_4027);
nand U4428 (N_4428,N_4040,N_4095);
and U4429 (N_4429,N_4114,N_4130);
and U4430 (N_4430,N_4002,N_4103);
and U4431 (N_4431,N_4116,N_4177);
nor U4432 (N_4432,N_4249,N_4172);
nor U4433 (N_4433,N_4202,N_4136);
or U4434 (N_4434,N_4215,N_4117);
nand U4435 (N_4435,N_4233,N_4148);
nand U4436 (N_4436,N_4068,N_4217);
xnor U4437 (N_4437,N_4246,N_4222);
or U4438 (N_4438,N_4225,N_4230);
xor U4439 (N_4439,N_4080,N_4036);
nand U4440 (N_4440,N_4229,N_4039);
nor U4441 (N_4441,N_4120,N_4106);
or U4442 (N_4442,N_4179,N_4038);
and U4443 (N_4443,N_4208,N_4137);
nand U4444 (N_4444,N_4060,N_4133);
nand U4445 (N_4445,N_4070,N_4166);
xnor U4446 (N_4446,N_4144,N_4194);
xnor U4447 (N_4447,N_4210,N_4059);
nor U4448 (N_4448,N_4138,N_4235);
xnor U4449 (N_4449,N_4105,N_4010);
nand U4450 (N_4450,N_4246,N_4064);
xor U4451 (N_4451,N_4008,N_4117);
xor U4452 (N_4452,N_4070,N_4111);
nand U4453 (N_4453,N_4004,N_4128);
or U4454 (N_4454,N_4205,N_4198);
or U4455 (N_4455,N_4183,N_4020);
and U4456 (N_4456,N_4121,N_4228);
nor U4457 (N_4457,N_4115,N_4017);
or U4458 (N_4458,N_4001,N_4174);
or U4459 (N_4459,N_4111,N_4098);
and U4460 (N_4460,N_4006,N_4151);
or U4461 (N_4461,N_4037,N_4004);
and U4462 (N_4462,N_4128,N_4243);
nor U4463 (N_4463,N_4109,N_4030);
or U4464 (N_4464,N_4105,N_4088);
xor U4465 (N_4465,N_4015,N_4184);
or U4466 (N_4466,N_4168,N_4114);
and U4467 (N_4467,N_4222,N_4126);
or U4468 (N_4468,N_4118,N_4138);
nor U4469 (N_4469,N_4223,N_4040);
xnor U4470 (N_4470,N_4064,N_4060);
or U4471 (N_4471,N_4198,N_4068);
nor U4472 (N_4472,N_4034,N_4092);
xnor U4473 (N_4473,N_4091,N_4161);
nand U4474 (N_4474,N_4073,N_4200);
xnor U4475 (N_4475,N_4149,N_4067);
or U4476 (N_4476,N_4052,N_4013);
or U4477 (N_4477,N_4085,N_4038);
nand U4478 (N_4478,N_4121,N_4098);
xor U4479 (N_4479,N_4152,N_4022);
nand U4480 (N_4480,N_4093,N_4180);
and U4481 (N_4481,N_4197,N_4095);
nand U4482 (N_4482,N_4222,N_4169);
and U4483 (N_4483,N_4175,N_4233);
or U4484 (N_4484,N_4073,N_4190);
nor U4485 (N_4485,N_4147,N_4018);
xor U4486 (N_4486,N_4133,N_4160);
nor U4487 (N_4487,N_4077,N_4041);
and U4488 (N_4488,N_4103,N_4217);
nand U4489 (N_4489,N_4204,N_4084);
xor U4490 (N_4490,N_4202,N_4029);
nand U4491 (N_4491,N_4044,N_4151);
xor U4492 (N_4492,N_4246,N_4032);
or U4493 (N_4493,N_4157,N_4153);
nor U4494 (N_4494,N_4089,N_4189);
and U4495 (N_4495,N_4023,N_4173);
or U4496 (N_4496,N_4227,N_4052);
nand U4497 (N_4497,N_4231,N_4015);
and U4498 (N_4498,N_4178,N_4119);
or U4499 (N_4499,N_4230,N_4087);
xor U4500 (N_4500,N_4253,N_4432);
nand U4501 (N_4501,N_4265,N_4441);
xnor U4502 (N_4502,N_4361,N_4256);
or U4503 (N_4503,N_4284,N_4403);
nand U4504 (N_4504,N_4400,N_4398);
and U4505 (N_4505,N_4438,N_4360);
and U4506 (N_4506,N_4419,N_4406);
nand U4507 (N_4507,N_4424,N_4324);
nand U4508 (N_4508,N_4478,N_4381);
or U4509 (N_4509,N_4270,N_4373);
and U4510 (N_4510,N_4405,N_4363);
and U4511 (N_4511,N_4312,N_4313);
and U4512 (N_4512,N_4455,N_4408);
or U4513 (N_4513,N_4495,N_4307);
or U4514 (N_4514,N_4470,N_4283);
and U4515 (N_4515,N_4379,N_4376);
and U4516 (N_4516,N_4453,N_4322);
or U4517 (N_4517,N_4479,N_4450);
xor U4518 (N_4518,N_4466,N_4415);
xnor U4519 (N_4519,N_4459,N_4349);
nand U4520 (N_4520,N_4334,N_4336);
nand U4521 (N_4521,N_4273,N_4250);
nor U4522 (N_4522,N_4282,N_4317);
and U4523 (N_4523,N_4449,N_4343);
xnor U4524 (N_4524,N_4416,N_4402);
nor U4525 (N_4525,N_4325,N_4304);
and U4526 (N_4526,N_4310,N_4393);
or U4527 (N_4527,N_4426,N_4315);
and U4528 (N_4528,N_4401,N_4355);
xnor U4529 (N_4529,N_4346,N_4443);
nand U4530 (N_4530,N_4293,N_4383);
nand U4531 (N_4531,N_4254,N_4366);
nand U4532 (N_4532,N_4338,N_4316);
nand U4533 (N_4533,N_4314,N_4371);
or U4534 (N_4534,N_4414,N_4289);
or U4535 (N_4535,N_4481,N_4431);
nor U4536 (N_4536,N_4380,N_4375);
nand U4537 (N_4537,N_4266,N_4413);
or U4538 (N_4538,N_4494,N_4428);
and U4539 (N_4539,N_4427,N_4412);
and U4540 (N_4540,N_4285,N_4255);
or U4541 (N_4541,N_4276,N_4461);
xor U4542 (N_4542,N_4445,N_4439);
or U4543 (N_4543,N_4287,N_4422);
xnor U4544 (N_4544,N_4446,N_4388);
or U4545 (N_4545,N_4301,N_4295);
or U4546 (N_4546,N_4409,N_4493);
or U4547 (N_4547,N_4430,N_4333);
xnor U4548 (N_4548,N_4264,N_4350);
nand U4549 (N_4549,N_4251,N_4327);
nand U4550 (N_4550,N_4257,N_4384);
or U4551 (N_4551,N_4252,N_4328);
nand U4552 (N_4552,N_4268,N_4407);
or U4553 (N_4553,N_4306,N_4442);
nor U4554 (N_4554,N_4302,N_4353);
xnor U4555 (N_4555,N_4435,N_4492);
xnor U4556 (N_4556,N_4485,N_4434);
and U4557 (N_4557,N_4420,N_4359);
nor U4558 (N_4558,N_4480,N_4299);
nor U4559 (N_4559,N_4364,N_4490);
nand U4560 (N_4560,N_4488,N_4354);
nand U4561 (N_4561,N_4323,N_4332);
nand U4562 (N_4562,N_4344,N_4260);
nor U4563 (N_4563,N_4468,N_4385);
nand U4564 (N_4564,N_4423,N_4374);
nand U4565 (N_4565,N_4464,N_4279);
nand U4566 (N_4566,N_4262,N_4308);
nor U4567 (N_4567,N_4347,N_4362);
nor U4568 (N_4568,N_4271,N_4311);
nor U4569 (N_4569,N_4305,N_4309);
or U4570 (N_4570,N_4281,N_4477);
nand U4571 (N_4571,N_4261,N_4418);
and U4572 (N_4572,N_4369,N_4404);
xor U4573 (N_4573,N_4397,N_4421);
or U4574 (N_4574,N_4280,N_4386);
and U4575 (N_4575,N_4462,N_4278);
nor U4576 (N_4576,N_4291,N_4368);
or U4577 (N_4577,N_4463,N_4473);
xor U4578 (N_4578,N_4319,N_4429);
nor U4579 (N_4579,N_4475,N_4296);
or U4580 (N_4580,N_4392,N_4411);
xor U4581 (N_4581,N_4297,N_4496);
and U4582 (N_4582,N_4274,N_4339);
and U4583 (N_4583,N_4356,N_4318);
and U4584 (N_4584,N_4341,N_4370);
and U4585 (N_4585,N_4436,N_4499);
xor U4586 (N_4586,N_4335,N_4396);
nor U4587 (N_4587,N_4457,N_4321);
and U4588 (N_4588,N_4292,N_4497);
and U4589 (N_4589,N_4377,N_4417);
and U4590 (N_4590,N_4331,N_4474);
and U4591 (N_4591,N_4467,N_4452);
or U4592 (N_4592,N_4342,N_4345);
nor U4593 (N_4593,N_4389,N_4486);
nor U4594 (N_4594,N_4437,N_4352);
and U4595 (N_4595,N_4294,N_4269);
nor U4596 (N_4596,N_4440,N_4382);
nand U4597 (N_4597,N_4348,N_4447);
xor U4598 (N_4598,N_4491,N_4365);
nor U4599 (N_4599,N_4275,N_4472);
and U4600 (N_4600,N_4410,N_4498);
and U4601 (N_4601,N_4337,N_4451);
xnor U4602 (N_4602,N_4367,N_4391);
nand U4603 (N_4603,N_4357,N_4272);
and U4604 (N_4604,N_4458,N_4425);
nor U4605 (N_4605,N_4288,N_4303);
and U4606 (N_4606,N_4465,N_4487);
xor U4607 (N_4607,N_4326,N_4399);
and U4608 (N_4608,N_4358,N_4390);
nand U4609 (N_4609,N_4394,N_4298);
nor U4610 (N_4610,N_4290,N_4395);
xor U4611 (N_4611,N_4263,N_4448);
nor U4612 (N_4612,N_4267,N_4469);
xnor U4613 (N_4613,N_4320,N_4444);
nor U4614 (N_4614,N_4277,N_4476);
xor U4615 (N_4615,N_4259,N_4378);
nor U4616 (N_4616,N_4460,N_4286);
nand U4617 (N_4617,N_4300,N_4433);
nand U4618 (N_4618,N_4387,N_4489);
and U4619 (N_4619,N_4483,N_4454);
nor U4620 (N_4620,N_4351,N_4484);
xnor U4621 (N_4621,N_4258,N_4340);
or U4622 (N_4622,N_4482,N_4329);
nor U4623 (N_4623,N_4372,N_4330);
xor U4624 (N_4624,N_4471,N_4456);
nand U4625 (N_4625,N_4395,N_4431);
nand U4626 (N_4626,N_4361,N_4304);
nand U4627 (N_4627,N_4333,N_4319);
nor U4628 (N_4628,N_4390,N_4447);
or U4629 (N_4629,N_4291,N_4320);
nand U4630 (N_4630,N_4345,N_4301);
or U4631 (N_4631,N_4366,N_4331);
or U4632 (N_4632,N_4467,N_4424);
nor U4633 (N_4633,N_4355,N_4348);
xnor U4634 (N_4634,N_4263,N_4402);
or U4635 (N_4635,N_4433,N_4498);
nor U4636 (N_4636,N_4370,N_4272);
nor U4637 (N_4637,N_4265,N_4467);
xor U4638 (N_4638,N_4349,N_4281);
and U4639 (N_4639,N_4272,N_4383);
nor U4640 (N_4640,N_4330,N_4438);
and U4641 (N_4641,N_4258,N_4486);
or U4642 (N_4642,N_4319,N_4266);
and U4643 (N_4643,N_4464,N_4494);
nand U4644 (N_4644,N_4369,N_4424);
xor U4645 (N_4645,N_4405,N_4487);
xnor U4646 (N_4646,N_4367,N_4402);
xor U4647 (N_4647,N_4263,N_4483);
or U4648 (N_4648,N_4445,N_4359);
and U4649 (N_4649,N_4420,N_4484);
nand U4650 (N_4650,N_4417,N_4361);
xnor U4651 (N_4651,N_4261,N_4380);
or U4652 (N_4652,N_4491,N_4347);
nor U4653 (N_4653,N_4423,N_4403);
xor U4654 (N_4654,N_4303,N_4454);
nand U4655 (N_4655,N_4429,N_4420);
xnor U4656 (N_4656,N_4358,N_4328);
or U4657 (N_4657,N_4388,N_4423);
nor U4658 (N_4658,N_4405,N_4360);
nor U4659 (N_4659,N_4418,N_4455);
and U4660 (N_4660,N_4280,N_4482);
nand U4661 (N_4661,N_4388,N_4284);
xnor U4662 (N_4662,N_4386,N_4301);
nor U4663 (N_4663,N_4374,N_4317);
nand U4664 (N_4664,N_4328,N_4364);
xor U4665 (N_4665,N_4406,N_4376);
nor U4666 (N_4666,N_4384,N_4492);
and U4667 (N_4667,N_4385,N_4292);
and U4668 (N_4668,N_4345,N_4404);
nor U4669 (N_4669,N_4464,N_4405);
or U4670 (N_4670,N_4405,N_4269);
xor U4671 (N_4671,N_4333,N_4496);
xor U4672 (N_4672,N_4306,N_4440);
nand U4673 (N_4673,N_4417,N_4368);
and U4674 (N_4674,N_4380,N_4327);
and U4675 (N_4675,N_4265,N_4281);
or U4676 (N_4676,N_4264,N_4270);
nor U4677 (N_4677,N_4398,N_4292);
xnor U4678 (N_4678,N_4368,N_4281);
nor U4679 (N_4679,N_4298,N_4263);
nand U4680 (N_4680,N_4254,N_4434);
nor U4681 (N_4681,N_4260,N_4434);
and U4682 (N_4682,N_4257,N_4364);
or U4683 (N_4683,N_4308,N_4260);
nand U4684 (N_4684,N_4433,N_4273);
nand U4685 (N_4685,N_4290,N_4250);
nor U4686 (N_4686,N_4495,N_4306);
nor U4687 (N_4687,N_4424,N_4361);
or U4688 (N_4688,N_4306,N_4294);
nand U4689 (N_4689,N_4347,N_4355);
xnor U4690 (N_4690,N_4457,N_4445);
xor U4691 (N_4691,N_4264,N_4420);
or U4692 (N_4692,N_4352,N_4375);
or U4693 (N_4693,N_4487,N_4292);
nor U4694 (N_4694,N_4431,N_4330);
xnor U4695 (N_4695,N_4288,N_4446);
nand U4696 (N_4696,N_4469,N_4494);
or U4697 (N_4697,N_4262,N_4348);
and U4698 (N_4698,N_4281,N_4410);
nand U4699 (N_4699,N_4458,N_4452);
and U4700 (N_4700,N_4307,N_4460);
or U4701 (N_4701,N_4388,N_4384);
nor U4702 (N_4702,N_4353,N_4395);
and U4703 (N_4703,N_4438,N_4290);
xnor U4704 (N_4704,N_4355,N_4333);
nand U4705 (N_4705,N_4497,N_4358);
and U4706 (N_4706,N_4371,N_4351);
nor U4707 (N_4707,N_4345,N_4292);
xor U4708 (N_4708,N_4417,N_4460);
xor U4709 (N_4709,N_4359,N_4407);
nor U4710 (N_4710,N_4257,N_4435);
and U4711 (N_4711,N_4331,N_4498);
and U4712 (N_4712,N_4314,N_4478);
nor U4713 (N_4713,N_4472,N_4376);
nor U4714 (N_4714,N_4309,N_4265);
or U4715 (N_4715,N_4376,N_4349);
xnor U4716 (N_4716,N_4376,N_4420);
and U4717 (N_4717,N_4489,N_4287);
or U4718 (N_4718,N_4318,N_4428);
or U4719 (N_4719,N_4344,N_4471);
or U4720 (N_4720,N_4333,N_4339);
nand U4721 (N_4721,N_4279,N_4331);
nand U4722 (N_4722,N_4366,N_4275);
nand U4723 (N_4723,N_4360,N_4314);
and U4724 (N_4724,N_4356,N_4425);
nor U4725 (N_4725,N_4304,N_4479);
and U4726 (N_4726,N_4361,N_4370);
and U4727 (N_4727,N_4402,N_4379);
nand U4728 (N_4728,N_4379,N_4333);
nor U4729 (N_4729,N_4271,N_4260);
xor U4730 (N_4730,N_4380,N_4439);
or U4731 (N_4731,N_4321,N_4400);
nand U4732 (N_4732,N_4493,N_4333);
nand U4733 (N_4733,N_4287,N_4348);
xnor U4734 (N_4734,N_4357,N_4388);
xnor U4735 (N_4735,N_4288,N_4311);
xnor U4736 (N_4736,N_4474,N_4322);
or U4737 (N_4737,N_4470,N_4363);
and U4738 (N_4738,N_4260,N_4425);
nor U4739 (N_4739,N_4393,N_4371);
and U4740 (N_4740,N_4266,N_4373);
nand U4741 (N_4741,N_4488,N_4370);
or U4742 (N_4742,N_4424,N_4396);
or U4743 (N_4743,N_4431,N_4314);
nand U4744 (N_4744,N_4298,N_4282);
xor U4745 (N_4745,N_4401,N_4282);
and U4746 (N_4746,N_4317,N_4312);
nand U4747 (N_4747,N_4467,N_4349);
and U4748 (N_4748,N_4488,N_4320);
xor U4749 (N_4749,N_4301,N_4488);
nand U4750 (N_4750,N_4729,N_4522);
and U4751 (N_4751,N_4523,N_4706);
nor U4752 (N_4752,N_4574,N_4635);
xnor U4753 (N_4753,N_4695,N_4598);
nand U4754 (N_4754,N_4735,N_4730);
and U4755 (N_4755,N_4543,N_4740);
nand U4756 (N_4756,N_4731,N_4525);
or U4757 (N_4757,N_4514,N_4709);
nand U4758 (N_4758,N_4736,N_4576);
or U4759 (N_4759,N_4542,N_4700);
and U4760 (N_4760,N_4556,N_4668);
or U4761 (N_4761,N_4654,N_4696);
and U4762 (N_4762,N_4573,N_4590);
nor U4763 (N_4763,N_4565,N_4728);
nand U4764 (N_4764,N_4610,N_4656);
nand U4765 (N_4765,N_4640,N_4701);
and U4766 (N_4766,N_4648,N_4680);
nand U4767 (N_4767,N_4732,N_4705);
nor U4768 (N_4768,N_4637,N_4725);
or U4769 (N_4769,N_4734,N_4539);
nand U4770 (N_4770,N_4620,N_4595);
xnor U4771 (N_4771,N_4607,N_4743);
or U4772 (N_4772,N_4739,N_4594);
xnor U4773 (N_4773,N_4692,N_4646);
nor U4774 (N_4774,N_4559,N_4727);
nand U4775 (N_4775,N_4592,N_4506);
nor U4776 (N_4776,N_4624,N_4658);
or U4777 (N_4777,N_4575,N_4512);
or U4778 (N_4778,N_4670,N_4631);
or U4779 (N_4779,N_4652,N_4558);
nand U4780 (N_4780,N_4644,N_4550);
xor U4781 (N_4781,N_4643,N_4665);
nand U4782 (N_4782,N_4638,N_4503);
and U4783 (N_4783,N_4521,N_4713);
nor U4784 (N_4784,N_4747,N_4589);
xnor U4785 (N_4785,N_4615,N_4555);
or U4786 (N_4786,N_4641,N_4642);
nand U4787 (N_4787,N_4714,N_4530);
nand U4788 (N_4788,N_4510,N_4614);
nor U4789 (N_4789,N_4672,N_4623);
and U4790 (N_4790,N_4564,N_4683);
xnor U4791 (N_4791,N_4702,N_4509);
or U4792 (N_4792,N_4679,N_4507);
and U4793 (N_4793,N_4687,N_4669);
nand U4794 (N_4794,N_4676,N_4562);
and U4795 (N_4795,N_4673,N_4529);
nor U4796 (N_4796,N_4712,N_4606);
nand U4797 (N_4797,N_4682,N_4703);
or U4798 (N_4798,N_4536,N_4678);
and U4799 (N_4799,N_4697,N_4519);
nor U4800 (N_4800,N_4588,N_4517);
nand U4801 (N_4801,N_4724,N_4694);
nand U4802 (N_4802,N_4616,N_4563);
xnor U4803 (N_4803,N_4544,N_4561);
nand U4804 (N_4804,N_4653,N_4534);
and U4805 (N_4805,N_4568,N_4508);
nor U4806 (N_4806,N_4632,N_4581);
xor U4807 (N_4807,N_4548,N_4571);
and U4808 (N_4808,N_4600,N_4520);
and U4809 (N_4809,N_4686,N_4621);
xor U4810 (N_4810,N_4546,N_4717);
and U4811 (N_4811,N_4533,N_4605);
nand U4812 (N_4812,N_4578,N_4636);
or U4813 (N_4813,N_4718,N_4720);
nor U4814 (N_4814,N_4707,N_4504);
xor U4815 (N_4815,N_4608,N_4580);
or U4816 (N_4816,N_4723,N_4622);
nand U4817 (N_4817,N_4655,N_4675);
nor U4818 (N_4818,N_4748,N_4500);
and U4819 (N_4819,N_4664,N_4742);
nand U4820 (N_4820,N_4557,N_4587);
or U4821 (N_4821,N_4535,N_4540);
nand U4822 (N_4822,N_4502,N_4560);
and U4823 (N_4823,N_4737,N_4552);
or U4824 (N_4824,N_4721,N_4527);
or U4825 (N_4825,N_4591,N_4567);
xor U4826 (N_4826,N_4667,N_4691);
xnor U4827 (N_4827,N_4746,N_4582);
xor U4828 (N_4828,N_4572,N_4505);
or U4829 (N_4829,N_4526,N_4603);
xnor U4830 (N_4830,N_4639,N_4599);
nand U4831 (N_4831,N_4551,N_4666);
xnor U4832 (N_4832,N_4566,N_4681);
or U4833 (N_4833,N_4733,N_4649);
or U4834 (N_4834,N_4651,N_4515);
or U4835 (N_4835,N_4726,N_4513);
xnor U4836 (N_4836,N_4613,N_4708);
nor U4837 (N_4837,N_4671,N_4627);
xor U4838 (N_4838,N_4518,N_4677);
nand U4839 (N_4839,N_4716,N_4531);
xor U4840 (N_4840,N_4626,N_4541);
nand U4841 (N_4841,N_4659,N_4569);
nand U4842 (N_4842,N_4633,N_4545);
and U4843 (N_4843,N_4593,N_4684);
xnor U4844 (N_4844,N_4538,N_4549);
xnor U4845 (N_4845,N_4617,N_4524);
xor U4846 (N_4846,N_4629,N_4601);
and U4847 (N_4847,N_4647,N_4645);
nand U4848 (N_4848,N_4618,N_4609);
or U4849 (N_4849,N_4602,N_4674);
xor U4850 (N_4850,N_4711,N_4685);
nor U4851 (N_4851,N_4744,N_4710);
or U4852 (N_4852,N_4688,N_4741);
and U4853 (N_4853,N_4570,N_4553);
nor U4854 (N_4854,N_4634,N_4597);
nor U4855 (N_4855,N_4577,N_4689);
nor U4856 (N_4856,N_4619,N_4660);
nand U4857 (N_4857,N_4583,N_4661);
nor U4858 (N_4858,N_4630,N_4690);
and U4859 (N_4859,N_4704,N_4604);
xor U4860 (N_4860,N_4749,N_4586);
or U4861 (N_4861,N_4585,N_4745);
nand U4862 (N_4862,N_4532,N_4596);
and U4863 (N_4863,N_4662,N_4722);
and U4864 (N_4864,N_4547,N_4501);
or U4865 (N_4865,N_4579,N_4693);
and U4866 (N_4866,N_4554,N_4628);
or U4867 (N_4867,N_4528,N_4625);
and U4868 (N_4868,N_4657,N_4715);
xnor U4869 (N_4869,N_4537,N_4663);
or U4870 (N_4870,N_4698,N_4650);
nor U4871 (N_4871,N_4511,N_4738);
or U4872 (N_4872,N_4516,N_4719);
and U4873 (N_4873,N_4584,N_4699);
nor U4874 (N_4874,N_4612,N_4611);
nand U4875 (N_4875,N_4710,N_4593);
nor U4876 (N_4876,N_4742,N_4691);
nor U4877 (N_4877,N_4712,N_4689);
or U4878 (N_4878,N_4666,N_4723);
nand U4879 (N_4879,N_4681,N_4601);
or U4880 (N_4880,N_4590,N_4619);
nand U4881 (N_4881,N_4734,N_4615);
xor U4882 (N_4882,N_4587,N_4676);
nor U4883 (N_4883,N_4652,N_4738);
xor U4884 (N_4884,N_4601,N_4640);
or U4885 (N_4885,N_4502,N_4705);
nor U4886 (N_4886,N_4595,N_4568);
and U4887 (N_4887,N_4527,N_4711);
and U4888 (N_4888,N_4542,N_4630);
or U4889 (N_4889,N_4710,N_4642);
and U4890 (N_4890,N_4574,N_4548);
nor U4891 (N_4891,N_4674,N_4501);
and U4892 (N_4892,N_4514,N_4725);
and U4893 (N_4893,N_4684,N_4525);
or U4894 (N_4894,N_4551,N_4707);
nor U4895 (N_4895,N_4566,N_4729);
or U4896 (N_4896,N_4698,N_4608);
nor U4897 (N_4897,N_4730,N_4536);
nor U4898 (N_4898,N_4688,N_4748);
xnor U4899 (N_4899,N_4661,N_4677);
and U4900 (N_4900,N_4620,N_4719);
nor U4901 (N_4901,N_4554,N_4664);
nand U4902 (N_4902,N_4640,N_4680);
or U4903 (N_4903,N_4542,N_4607);
and U4904 (N_4904,N_4680,N_4721);
nor U4905 (N_4905,N_4672,N_4529);
and U4906 (N_4906,N_4664,N_4530);
nand U4907 (N_4907,N_4708,N_4735);
and U4908 (N_4908,N_4537,N_4510);
or U4909 (N_4909,N_4670,N_4606);
nor U4910 (N_4910,N_4617,N_4555);
nor U4911 (N_4911,N_4677,N_4740);
and U4912 (N_4912,N_4645,N_4549);
or U4913 (N_4913,N_4553,N_4581);
and U4914 (N_4914,N_4716,N_4613);
and U4915 (N_4915,N_4718,N_4651);
nand U4916 (N_4916,N_4667,N_4747);
or U4917 (N_4917,N_4737,N_4536);
nor U4918 (N_4918,N_4576,N_4603);
nand U4919 (N_4919,N_4587,N_4718);
nand U4920 (N_4920,N_4734,N_4547);
or U4921 (N_4921,N_4714,N_4543);
or U4922 (N_4922,N_4570,N_4581);
and U4923 (N_4923,N_4567,N_4533);
nor U4924 (N_4924,N_4684,N_4589);
nand U4925 (N_4925,N_4528,N_4567);
or U4926 (N_4926,N_4713,N_4603);
or U4927 (N_4927,N_4543,N_4709);
xnor U4928 (N_4928,N_4590,N_4676);
xnor U4929 (N_4929,N_4612,N_4691);
nand U4930 (N_4930,N_4573,N_4554);
xnor U4931 (N_4931,N_4700,N_4695);
nor U4932 (N_4932,N_4532,N_4584);
nor U4933 (N_4933,N_4723,N_4572);
nand U4934 (N_4934,N_4604,N_4624);
nand U4935 (N_4935,N_4723,N_4736);
xnor U4936 (N_4936,N_4606,N_4534);
nand U4937 (N_4937,N_4691,N_4714);
or U4938 (N_4938,N_4542,N_4609);
nor U4939 (N_4939,N_4532,N_4531);
xor U4940 (N_4940,N_4541,N_4582);
xnor U4941 (N_4941,N_4691,N_4589);
nand U4942 (N_4942,N_4600,N_4723);
and U4943 (N_4943,N_4692,N_4517);
and U4944 (N_4944,N_4552,N_4668);
or U4945 (N_4945,N_4546,N_4679);
nor U4946 (N_4946,N_4590,N_4520);
nor U4947 (N_4947,N_4676,N_4653);
nor U4948 (N_4948,N_4561,N_4689);
xnor U4949 (N_4949,N_4513,N_4736);
and U4950 (N_4950,N_4618,N_4621);
and U4951 (N_4951,N_4637,N_4747);
nor U4952 (N_4952,N_4554,N_4679);
or U4953 (N_4953,N_4689,N_4704);
or U4954 (N_4954,N_4723,N_4548);
nand U4955 (N_4955,N_4661,N_4609);
or U4956 (N_4956,N_4677,N_4704);
or U4957 (N_4957,N_4587,N_4736);
nand U4958 (N_4958,N_4699,N_4557);
nand U4959 (N_4959,N_4649,N_4585);
and U4960 (N_4960,N_4527,N_4503);
nor U4961 (N_4961,N_4533,N_4548);
or U4962 (N_4962,N_4509,N_4505);
and U4963 (N_4963,N_4643,N_4569);
xor U4964 (N_4964,N_4649,N_4607);
nor U4965 (N_4965,N_4515,N_4585);
and U4966 (N_4966,N_4639,N_4721);
xor U4967 (N_4967,N_4660,N_4708);
nor U4968 (N_4968,N_4603,N_4504);
or U4969 (N_4969,N_4615,N_4670);
nand U4970 (N_4970,N_4728,N_4616);
nand U4971 (N_4971,N_4558,N_4570);
xor U4972 (N_4972,N_4576,N_4577);
nand U4973 (N_4973,N_4515,N_4589);
nand U4974 (N_4974,N_4587,N_4677);
nor U4975 (N_4975,N_4629,N_4549);
nor U4976 (N_4976,N_4697,N_4736);
nor U4977 (N_4977,N_4643,N_4644);
and U4978 (N_4978,N_4557,N_4747);
xnor U4979 (N_4979,N_4601,N_4740);
and U4980 (N_4980,N_4625,N_4717);
nor U4981 (N_4981,N_4646,N_4511);
and U4982 (N_4982,N_4592,N_4597);
nor U4983 (N_4983,N_4559,N_4679);
nand U4984 (N_4984,N_4708,N_4670);
or U4985 (N_4985,N_4576,N_4640);
and U4986 (N_4986,N_4560,N_4597);
xor U4987 (N_4987,N_4544,N_4734);
nor U4988 (N_4988,N_4749,N_4725);
nand U4989 (N_4989,N_4617,N_4540);
nor U4990 (N_4990,N_4641,N_4507);
nor U4991 (N_4991,N_4523,N_4572);
and U4992 (N_4992,N_4508,N_4644);
or U4993 (N_4993,N_4562,N_4555);
nor U4994 (N_4994,N_4721,N_4591);
xnor U4995 (N_4995,N_4596,N_4547);
and U4996 (N_4996,N_4576,N_4571);
nor U4997 (N_4997,N_4735,N_4728);
xor U4998 (N_4998,N_4653,N_4560);
nor U4999 (N_4999,N_4672,N_4683);
and U5000 (N_5000,N_4874,N_4825);
nand U5001 (N_5001,N_4761,N_4852);
nand U5002 (N_5002,N_4848,N_4992);
or U5003 (N_5003,N_4860,N_4797);
xor U5004 (N_5004,N_4876,N_4954);
nand U5005 (N_5005,N_4792,N_4804);
and U5006 (N_5006,N_4779,N_4760);
xnor U5007 (N_5007,N_4914,N_4888);
or U5008 (N_5008,N_4961,N_4824);
xnor U5009 (N_5009,N_4834,N_4894);
nor U5010 (N_5010,N_4999,N_4991);
nor U5011 (N_5011,N_4968,N_4780);
xor U5012 (N_5012,N_4941,N_4892);
or U5013 (N_5013,N_4886,N_4767);
nand U5014 (N_5014,N_4960,N_4762);
or U5015 (N_5015,N_4783,N_4776);
xnor U5016 (N_5016,N_4808,N_4880);
xor U5017 (N_5017,N_4995,N_4922);
nor U5018 (N_5018,N_4869,N_4963);
nor U5019 (N_5019,N_4842,N_4890);
or U5020 (N_5020,N_4847,N_4822);
nor U5021 (N_5021,N_4998,N_4775);
or U5022 (N_5022,N_4840,N_4910);
or U5023 (N_5023,N_4996,N_4994);
nand U5024 (N_5024,N_4906,N_4772);
or U5025 (N_5025,N_4789,N_4782);
and U5026 (N_5026,N_4909,N_4920);
and U5027 (N_5027,N_4974,N_4969);
nand U5028 (N_5028,N_4957,N_4939);
nand U5029 (N_5029,N_4976,N_4793);
nand U5030 (N_5030,N_4943,N_4878);
and U5031 (N_5031,N_4917,N_4815);
and U5032 (N_5032,N_4927,N_4955);
or U5033 (N_5033,N_4811,N_4765);
or U5034 (N_5034,N_4831,N_4981);
nor U5035 (N_5035,N_4774,N_4838);
and U5036 (N_5036,N_4796,N_4865);
xor U5037 (N_5037,N_4889,N_4788);
xor U5038 (N_5038,N_4778,N_4757);
and U5039 (N_5039,N_4752,N_4802);
and U5040 (N_5040,N_4987,N_4785);
or U5041 (N_5041,N_4944,N_4828);
and U5042 (N_5042,N_4826,N_4947);
and U5043 (N_5043,N_4977,N_4845);
and U5044 (N_5044,N_4854,N_4863);
nor U5045 (N_5045,N_4951,N_4931);
xnor U5046 (N_5046,N_4953,N_4884);
or U5047 (N_5047,N_4855,N_4897);
nand U5048 (N_5048,N_4754,N_4933);
nand U5049 (N_5049,N_4769,N_4791);
nor U5050 (N_5050,N_4934,N_4895);
or U5051 (N_5051,N_4965,N_4883);
nand U5052 (N_5052,N_4940,N_4921);
nor U5053 (N_5053,N_4866,N_4758);
xnor U5054 (N_5054,N_4836,N_4784);
nor U5055 (N_5055,N_4989,N_4893);
nor U5056 (N_5056,N_4882,N_4820);
nand U5057 (N_5057,N_4786,N_4835);
nor U5058 (N_5058,N_4972,N_4872);
or U5059 (N_5059,N_4839,N_4849);
and U5060 (N_5060,N_4982,N_4918);
nor U5061 (N_5061,N_4861,N_4912);
xnor U5062 (N_5062,N_4948,N_4794);
nand U5063 (N_5063,N_4807,N_4818);
nand U5064 (N_5064,N_4908,N_4871);
and U5065 (N_5065,N_4873,N_4923);
or U5066 (N_5066,N_4902,N_4952);
or U5067 (N_5067,N_4904,N_4875);
xor U5068 (N_5068,N_4980,N_4870);
or U5069 (N_5069,N_4903,N_4830);
or U5070 (N_5070,N_4853,N_4935);
xor U5071 (N_5071,N_4915,N_4959);
nor U5072 (N_5072,N_4877,N_4958);
xor U5073 (N_5073,N_4984,N_4973);
nor U5074 (N_5074,N_4814,N_4925);
or U5075 (N_5075,N_4881,N_4887);
nand U5076 (N_5076,N_4841,N_4810);
nor U5077 (N_5077,N_4942,N_4805);
or U5078 (N_5078,N_4809,N_4885);
and U5079 (N_5079,N_4898,N_4781);
nand U5080 (N_5080,N_4859,N_4829);
nand U5081 (N_5081,N_4764,N_4905);
and U5082 (N_5082,N_4799,N_4901);
nand U5083 (N_5083,N_4827,N_4879);
nand U5084 (N_5084,N_4756,N_4770);
or U5085 (N_5085,N_4913,N_4993);
and U5086 (N_5086,N_4856,N_4787);
xor U5087 (N_5087,N_4988,N_4766);
nor U5088 (N_5088,N_4819,N_4864);
xor U5089 (N_5089,N_4777,N_4813);
and U5090 (N_5090,N_4946,N_4997);
or U5091 (N_5091,N_4773,N_4753);
xnor U5092 (N_5092,N_4966,N_4983);
or U5093 (N_5093,N_4967,N_4771);
xor U5094 (N_5094,N_4862,N_4978);
xor U5095 (N_5095,N_4800,N_4936);
nand U5096 (N_5096,N_4985,N_4911);
or U5097 (N_5097,N_4962,N_4975);
or U5098 (N_5098,N_4755,N_4812);
and U5099 (N_5099,N_4751,N_4857);
or U5100 (N_5100,N_4945,N_4768);
xnor U5101 (N_5101,N_4896,N_4990);
nor U5102 (N_5102,N_4759,N_4823);
nand U5103 (N_5103,N_4803,N_4801);
nand U5104 (N_5104,N_4900,N_4971);
nor U5105 (N_5105,N_4832,N_4790);
nor U5106 (N_5106,N_4891,N_4795);
nand U5107 (N_5107,N_4816,N_4858);
and U5108 (N_5108,N_4907,N_4916);
and U5109 (N_5109,N_4750,N_4970);
nor U5110 (N_5110,N_4846,N_4821);
nand U5111 (N_5111,N_4964,N_4930);
and U5112 (N_5112,N_4850,N_4950);
nor U5113 (N_5113,N_4937,N_4986);
xor U5114 (N_5114,N_4806,N_4979);
and U5115 (N_5115,N_4798,N_4924);
nand U5116 (N_5116,N_4843,N_4949);
and U5117 (N_5117,N_4851,N_4833);
nor U5118 (N_5118,N_4817,N_4926);
nor U5119 (N_5119,N_4956,N_4938);
or U5120 (N_5120,N_4844,N_4929);
or U5121 (N_5121,N_4919,N_4868);
or U5122 (N_5122,N_4899,N_4932);
nand U5123 (N_5123,N_4837,N_4928);
xnor U5124 (N_5124,N_4867,N_4763);
or U5125 (N_5125,N_4966,N_4795);
nand U5126 (N_5126,N_4834,N_4761);
nand U5127 (N_5127,N_4968,N_4881);
nand U5128 (N_5128,N_4923,N_4937);
nand U5129 (N_5129,N_4831,N_4906);
or U5130 (N_5130,N_4916,N_4956);
and U5131 (N_5131,N_4925,N_4841);
or U5132 (N_5132,N_4858,N_4947);
xor U5133 (N_5133,N_4911,N_4881);
xnor U5134 (N_5134,N_4955,N_4853);
and U5135 (N_5135,N_4981,N_4785);
or U5136 (N_5136,N_4827,N_4885);
or U5137 (N_5137,N_4757,N_4853);
nand U5138 (N_5138,N_4757,N_4892);
xor U5139 (N_5139,N_4984,N_4813);
nor U5140 (N_5140,N_4822,N_4872);
xnor U5141 (N_5141,N_4826,N_4890);
xnor U5142 (N_5142,N_4803,N_4817);
xnor U5143 (N_5143,N_4940,N_4831);
xor U5144 (N_5144,N_4924,N_4855);
or U5145 (N_5145,N_4994,N_4882);
xnor U5146 (N_5146,N_4969,N_4998);
xnor U5147 (N_5147,N_4937,N_4841);
xnor U5148 (N_5148,N_4751,N_4863);
nor U5149 (N_5149,N_4903,N_4796);
or U5150 (N_5150,N_4799,N_4969);
or U5151 (N_5151,N_4912,N_4849);
xnor U5152 (N_5152,N_4928,N_4799);
xor U5153 (N_5153,N_4879,N_4795);
nor U5154 (N_5154,N_4815,N_4956);
xnor U5155 (N_5155,N_4813,N_4809);
nor U5156 (N_5156,N_4982,N_4761);
nand U5157 (N_5157,N_4955,N_4863);
nor U5158 (N_5158,N_4967,N_4812);
nor U5159 (N_5159,N_4902,N_4782);
nor U5160 (N_5160,N_4754,N_4916);
or U5161 (N_5161,N_4829,N_4932);
or U5162 (N_5162,N_4995,N_4849);
nor U5163 (N_5163,N_4794,N_4801);
xor U5164 (N_5164,N_4960,N_4954);
nand U5165 (N_5165,N_4812,N_4898);
nand U5166 (N_5166,N_4752,N_4843);
nor U5167 (N_5167,N_4917,N_4915);
or U5168 (N_5168,N_4916,N_4979);
xnor U5169 (N_5169,N_4830,N_4921);
nand U5170 (N_5170,N_4807,N_4945);
xnor U5171 (N_5171,N_4959,N_4998);
and U5172 (N_5172,N_4759,N_4985);
nor U5173 (N_5173,N_4806,N_4937);
or U5174 (N_5174,N_4992,N_4990);
nor U5175 (N_5175,N_4932,N_4909);
nor U5176 (N_5176,N_4779,N_4859);
xnor U5177 (N_5177,N_4826,N_4908);
nor U5178 (N_5178,N_4955,N_4948);
or U5179 (N_5179,N_4920,N_4781);
and U5180 (N_5180,N_4850,N_4878);
xnor U5181 (N_5181,N_4944,N_4998);
nand U5182 (N_5182,N_4831,N_4862);
and U5183 (N_5183,N_4764,N_4931);
nand U5184 (N_5184,N_4755,N_4943);
or U5185 (N_5185,N_4954,N_4764);
nor U5186 (N_5186,N_4977,N_4804);
xnor U5187 (N_5187,N_4845,N_4836);
and U5188 (N_5188,N_4808,N_4915);
nand U5189 (N_5189,N_4808,N_4769);
nor U5190 (N_5190,N_4864,N_4784);
nand U5191 (N_5191,N_4952,N_4913);
or U5192 (N_5192,N_4799,N_4936);
xnor U5193 (N_5193,N_4833,N_4977);
nand U5194 (N_5194,N_4976,N_4904);
xnor U5195 (N_5195,N_4874,N_4847);
or U5196 (N_5196,N_4953,N_4969);
or U5197 (N_5197,N_4864,N_4840);
or U5198 (N_5198,N_4827,N_4860);
or U5199 (N_5199,N_4993,N_4808);
nor U5200 (N_5200,N_4991,N_4983);
nand U5201 (N_5201,N_4840,N_4924);
or U5202 (N_5202,N_4752,N_4909);
or U5203 (N_5203,N_4808,N_4965);
nor U5204 (N_5204,N_4986,N_4765);
and U5205 (N_5205,N_4754,N_4919);
and U5206 (N_5206,N_4889,N_4896);
or U5207 (N_5207,N_4960,N_4764);
xor U5208 (N_5208,N_4966,N_4816);
nor U5209 (N_5209,N_4886,N_4874);
nand U5210 (N_5210,N_4755,N_4851);
nor U5211 (N_5211,N_4918,N_4922);
or U5212 (N_5212,N_4798,N_4759);
or U5213 (N_5213,N_4896,N_4837);
nand U5214 (N_5214,N_4916,N_4955);
or U5215 (N_5215,N_4954,N_4920);
nand U5216 (N_5216,N_4982,N_4894);
xnor U5217 (N_5217,N_4911,N_4821);
and U5218 (N_5218,N_4806,N_4961);
and U5219 (N_5219,N_4998,N_4997);
and U5220 (N_5220,N_4784,N_4952);
nand U5221 (N_5221,N_4823,N_4752);
xnor U5222 (N_5222,N_4896,N_4867);
xor U5223 (N_5223,N_4754,N_4781);
or U5224 (N_5224,N_4972,N_4954);
nand U5225 (N_5225,N_4758,N_4983);
or U5226 (N_5226,N_4874,N_4831);
nor U5227 (N_5227,N_4944,N_4989);
and U5228 (N_5228,N_4909,N_4768);
and U5229 (N_5229,N_4793,N_4925);
xnor U5230 (N_5230,N_4971,N_4944);
nand U5231 (N_5231,N_4891,N_4920);
xor U5232 (N_5232,N_4967,N_4871);
xnor U5233 (N_5233,N_4846,N_4761);
and U5234 (N_5234,N_4790,N_4844);
or U5235 (N_5235,N_4997,N_4873);
nor U5236 (N_5236,N_4788,N_4824);
nor U5237 (N_5237,N_4917,N_4990);
nand U5238 (N_5238,N_4870,N_4792);
and U5239 (N_5239,N_4866,N_4971);
nor U5240 (N_5240,N_4934,N_4870);
nor U5241 (N_5241,N_4872,N_4979);
nand U5242 (N_5242,N_4764,N_4769);
or U5243 (N_5243,N_4886,N_4904);
or U5244 (N_5244,N_4847,N_4751);
or U5245 (N_5245,N_4971,N_4798);
nand U5246 (N_5246,N_4767,N_4855);
nor U5247 (N_5247,N_4994,N_4984);
and U5248 (N_5248,N_4767,N_4753);
nor U5249 (N_5249,N_4972,N_4996);
nor U5250 (N_5250,N_5083,N_5040);
or U5251 (N_5251,N_5039,N_5063);
nand U5252 (N_5252,N_5117,N_5069);
or U5253 (N_5253,N_5044,N_5137);
nor U5254 (N_5254,N_5087,N_5208);
and U5255 (N_5255,N_5207,N_5158);
xor U5256 (N_5256,N_5170,N_5007);
xor U5257 (N_5257,N_5078,N_5176);
nor U5258 (N_5258,N_5197,N_5179);
nor U5259 (N_5259,N_5169,N_5230);
nor U5260 (N_5260,N_5077,N_5100);
nor U5261 (N_5261,N_5203,N_5235);
nand U5262 (N_5262,N_5177,N_5184);
xnor U5263 (N_5263,N_5062,N_5059);
nand U5264 (N_5264,N_5075,N_5135);
and U5265 (N_5265,N_5181,N_5022);
nand U5266 (N_5266,N_5233,N_5138);
or U5267 (N_5267,N_5157,N_5148);
nor U5268 (N_5268,N_5231,N_5155);
xor U5269 (N_5269,N_5103,N_5133);
nand U5270 (N_5270,N_5162,N_5123);
and U5271 (N_5271,N_5206,N_5191);
nand U5272 (N_5272,N_5125,N_5173);
nor U5273 (N_5273,N_5067,N_5196);
xnor U5274 (N_5274,N_5037,N_5072);
or U5275 (N_5275,N_5029,N_5114);
xor U5276 (N_5276,N_5149,N_5028);
nor U5277 (N_5277,N_5030,N_5056);
or U5278 (N_5278,N_5201,N_5051);
and U5279 (N_5279,N_5036,N_5057);
nand U5280 (N_5280,N_5113,N_5108);
and U5281 (N_5281,N_5175,N_5064);
xor U5282 (N_5282,N_5247,N_5147);
and U5283 (N_5283,N_5046,N_5214);
nand U5284 (N_5284,N_5106,N_5186);
or U5285 (N_5285,N_5033,N_5243);
nor U5286 (N_5286,N_5105,N_5112);
nand U5287 (N_5287,N_5248,N_5084);
and U5288 (N_5288,N_5002,N_5190);
or U5289 (N_5289,N_5187,N_5021);
or U5290 (N_5290,N_5086,N_5094);
nand U5291 (N_5291,N_5145,N_5226);
nand U5292 (N_5292,N_5229,N_5224);
xor U5293 (N_5293,N_5095,N_5150);
nor U5294 (N_5294,N_5042,N_5122);
xnor U5295 (N_5295,N_5134,N_5006);
and U5296 (N_5296,N_5241,N_5058);
or U5297 (N_5297,N_5119,N_5120);
or U5298 (N_5298,N_5128,N_5136);
nor U5299 (N_5299,N_5121,N_5204);
xnor U5300 (N_5300,N_5140,N_5219);
nand U5301 (N_5301,N_5070,N_5003);
and U5302 (N_5302,N_5218,N_5242);
nor U5303 (N_5303,N_5244,N_5188);
xnor U5304 (N_5304,N_5000,N_5160);
and U5305 (N_5305,N_5152,N_5223);
or U5306 (N_5306,N_5054,N_5055);
nor U5307 (N_5307,N_5161,N_5245);
nand U5308 (N_5308,N_5154,N_5142);
and U5309 (N_5309,N_5085,N_5008);
xor U5310 (N_5310,N_5130,N_5004);
and U5311 (N_5311,N_5220,N_5068);
xor U5312 (N_5312,N_5027,N_5045);
or U5313 (N_5313,N_5129,N_5144);
and U5314 (N_5314,N_5111,N_5115);
and U5315 (N_5315,N_5109,N_5227);
nand U5316 (N_5316,N_5092,N_5198);
or U5317 (N_5317,N_5211,N_5168);
nor U5318 (N_5318,N_5182,N_5060);
nor U5319 (N_5319,N_5172,N_5139);
xor U5320 (N_5320,N_5192,N_5165);
and U5321 (N_5321,N_5232,N_5061);
nor U5322 (N_5322,N_5126,N_5228);
or U5323 (N_5323,N_5026,N_5052);
nand U5324 (N_5324,N_5193,N_5038);
nand U5325 (N_5325,N_5163,N_5013);
or U5326 (N_5326,N_5011,N_5239);
xnor U5327 (N_5327,N_5159,N_5215);
or U5328 (N_5328,N_5093,N_5050);
and U5329 (N_5329,N_5189,N_5222);
nor U5330 (N_5330,N_5116,N_5071);
nand U5331 (N_5331,N_5110,N_5143);
xor U5332 (N_5332,N_5020,N_5034);
or U5333 (N_5333,N_5210,N_5019);
and U5334 (N_5334,N_5194,N_5081);
or U5335 (N_5335,N_5164,N_5088);
and U5336 (N_5336,N_5171,N_5049);
nor U5337 (N_5337,N_5225,N_5249);
xnor U5338 (N_5338,N_5018,N_5216);
or U5339 (N_5339,N_5041,N_5066);
or U5340 (N_5340,N_5017,N_5118);
nand U5341 (N_5341,N_5131,N_5209);
nand U5342 (N_5342,N_5174,N_5183);
or U5343 (N_5343,N_5031,N_5202);
nand U5344 (N_5344,N_5153,N_5246);
xnor U5345 (N_5345,N_5200,N_5236);
nand U5346 (N_5346,N_5195,N_5016);
and U5347 (N_5347,N_5014,N_5097);
nand U5348 (N_5348,N_5080,N_5217);
xnor U5349 (N_5349,N_5104,N_5141);
or U5350 (N_5350,N_5151,N_5076);
nor U5351 (N_5351,N_5047,N_5221);
nand U5352 (N_5352,N_5096,N_5180);
xor U5353 (N_5353,N_5032,N_5199);
or U5354 (N_5354,N_5012,N_5107);
nor U5355 (N_5355,N_5127,N_5025);
and U5356 (N_5356,N_5082,N_5098);
or U5357 (N_5357,N_5073,N_5102);
nor U5358 (N_5358,N_5035,N_5132);
xnor U5359 (N_5359,N_5024,N_5237);
or U5360 (N_5360,N_5079,N_5238);
nand U5361 (N_5361,N_5005,N_5001);
or U5362 (N_5362,N_5166,N_5090);
nand U5363 (N_5363,N_5015,N_5234);
or U5364 (N_5364,N_5205,N_5009);
nor U5365 (N_5365,N_5091,N_5213);
nand U5366 (N_5366,N_5146,N_5240);
xor U5367 (N_5367,N_5167,N_5101);
xor U5368 (N_5368,N_5099,N_5156);
and U5369 (N_5369,N_5048,N_5065);
xor U5370 (N_5370,N_5043,N_5023);
or U5371 (N_5371,N_5178,N_5074);
nor U5372 (N_5372,N_5124,N_5089);
nand U5373 (N_5373,N_5010,N_5053);
nand U5374 (N_5374,N_5185,N_5212);
nand U5375 (N_5375,N_5007,N_5038);
xnor U5376 (N_5376,N_5194,N_5056);
nand U5377 (N_5377,N_5033,N_5034);
and U5378 (N_5378,N_5139,N_5099);
and U5379 (N_5379,N_5215,N_5093);
nand U5380 (N_5380,N_5223,N_5239);
or U5381 (N_5381,N_5160,N_5234);
nand U5382 (N_5382,N_5055,N_5064);
nor U5383 (N_5383,N_5042,N_5115);
xnor U5384 (N_5384,N_5053,N_5115);
xnor U5385 (N_5385,N_5097,N_5162);
or U5386 (N_5386,N_5210,N_5000);
nor U5387 (N_5387,N_5163,N_5080);
or U5388 (N_5388,N_5186,N_5051);
xor U5389 (N_5389,N_5074,N_5118);
xor U5390 (N_5390,N_5201,N_5049);
nor U5391 (N_5391,N_5158,N_5133);
xor U5392 (N_5392,N_5148,N_5065);
nor U5393 (N_5393,N_5220,N_5044);
xor U5394 (N_5394,N_5041,N_5110);
or U5395 (N_5395,N_5154,N_5189);
or U5396 (N_5396,N_5166,N_5052);
nand U5397 (N_5397,N_5120,N_5111);
xnor U5398 (N_5398,N_5029,N_5112);
nor U5399 (N_5399,N_5080,N_5052);
and U5400 (N_5400,N_5227,N_5094);
nor U5401 (N_5401,N_5109,N_5212);
nor U5402 (N_5402,N_5089,N_5099);
nand U5403 (N_5403,N_5036,N_5148);
and U5404 (N_5404,N_5189,N_5079);
nor U5405 (N_5405,N_5020,N_5106);
xnor U5406 (N_5406,N_5061,N_5111);
nand U5407 (N_5407,N_5225,N_5126);
nor U5408 (N_5408,N_5158,N_5004);
xnor U5409 (N_5409,N_5216,N_5009);
and U5410 (N_5410,N_5116,N_5017);
nand U5411 (N_5411,N_5095,N_5086);
nor U5412 (N_5412,N_5084,N_5240);
or U5413 (N_5413,N_5224,N_5181);
nor U5414 (N_5414,N_5097,N_5083);
nand U5415 (N_5415,N_5147,N_5241);
and U5416 (N_5416,N_5069,N_5235);
and U5417 (N_5417,N_5196,N_5220);
nor U5418 (N_5418,N_5155,N_5131);
nor U5419 (N_5419,N_5000,N_5111);
nor U5420 (N_5420,N_5072,N_5062);
nor U5421 (N_5421,N_5042,N_5220);
nor U5422 (N_5422,N_5236,N_5146);
nor U5423 (N_5423,N_5210,N_5073);
nor U5424 (N_5424,N_5232,N_5096);
and U5425 (N_5425,N_5215,N_5228);
xor U5426 (N_5426,N_5145,N_5155);
or U5427 (N_5427,N_5144,N_5127);
xnor U5428 (N_5428,N_5140,N_5002);
or U5429 (N_5429,N_5017,N_5141);
xor U5430 (N_5430,N_5168,N_5173);
nor U5431 (N_5431,N_5093,N_5102);
nand U5432 (N_5432,N_5129,N_5175);
or U5433 (N_5433,N_5023,N_5186);
or U5434 (N_5434,N_5192,N_5228);
nand U5435 (N_5435,N_5049,N_5162);
xor U5436 (N_5436,N_5221,N_5134);
and U5437 (N_5437,N_5040,N_5231);
xor U5438 (N_5438,N_5070,N_5211);
or U5439 (N_5439,N_5013,N_5205);
and U5440 (N_5440,N_5012,N_5066);
nor U5441 (N_5441,N_5181,N_5206);
nor U5442 (N_5442,N_5152,N_5237);
xor U5443 (N_5443,N_5195,N_5127);
xnor U5444 (N_5444,N_5100,N_5225);
nor U5445 (N_5445,N_5224,N_5045);
nor U5446 (N_5446,N_5152,N_5069);
nor U5447 (N_5447,N_5051,N_5001);
xnor U5448 (N_5448,N_5149,N_5011);
xnor U5449 (N_5449,N_5207,N_5053);
nor U5450 (N_5450,N_5049,N_5060);
or U5451 (N_5451,N_5146,N_5217);
nor U5452 (N_5452,N_5094,N_5153);
nor U5453 (N_5453,N_5231,N_5024);
nand U5454 (N_5454,N_5220,N_5230);
nand U5455 (N_5455,N_5188,N_5077);
nand U5456 (N_5456,N_5102,N_5081);
or U5457 (N_5457,N_5156,N_5201);
xor U5458 (N_5458,N_5181,N_5174);
nor U5459 (N_5459,N_5136,N_5166);
xor U5460 (N_5460,N_5129,N_5046);
nand U5461 (N_5461,N_5010,N_5042);
and U5462 (N_5462,N_5249,N_5114);
xor U5463 (N_5463,N_5052,N_5180);
nand U5464 (N_5464,N_5038,N_5111);
xor U5465 (N_5465,N_5094,N_5063);
nor U5466 (N_5466,N_5114,N_5200);
nor U5467 (N_5467,N_5009,N_5242);
or U5468 (N_5468,N_5232,N_5092);
or U5469 (N_5469,N_5087,N_5111);
and U5470 (N_5470,N_5174,N_5108);
nor U5471 (N_5471,N_5049,N_5099);
nand U5472 (N_5472,N_5246,N_5184);
and U5473 (N_5473,N_5247,N_5231);
or U5474 (N_5474,N_5211,N_5038);
xor U5475 (N_5475,N_5200,N_5164);
and U5476 (N_5476,N_5092,N_5098);
nor U5477 (N_5477,N_5041,N_5007);
nor U5478 (N_5478,N_5124,N_5218);
and U5479 (N_5479,N_5216,N_5236);
and U5480 (N_5480,N_5042,N_5012);
nor U5481 (N_5481,N_5173,N_5134);
nand U5482 (N_5482,N_5060,N_5170);
and U5483 (N_5483,N_5130,N_5194);
xor U5484 (N_5484,N_5156,N_5157);
nor U5485 (N_5485,N_5080,N_5169);
nand U5486 (N_5486,N_5095,N_5148);
nor U5487 (N_5487,N_5011,N_5066);
or U5488 (N_5488,N_5051,N_5214);
nor U5489 (N_5489,N_5208,N_5221);
and U5490 (N_5490,N_5020,N_5122);
nor U5491 (N_5491,N_5175,N_5248);
xnor U5492 (N_5492,N_5078,N_5031);
xnor U5493 (N_5493,N_5153,N_5123);
xnor U5494 (N_5494,N_5220,N_5229);
or U5495 (N_5495,N_5008,N_5152);
and U5496 (N_5496,N_5174,N_5192);
nand U5497 (N_5497,N_5165,N_5231);
nand U5498 (N_5498,N_5046,N_5175);
or U5499 (N_5499,N_5049,N_5197);
or U5500 (N_5500,N_5346,N_5384);
or U5501 (N_5501,N_5315,N_5336);
and U5502 (N_5502,N_5316,N_5335);
or U5503 (N_5503,N_5269,N_5292);
or U5504 (N_5504,N_5308,N_5264);
and U5505 (N_5505,N_5485,N_5405);
nor U5506 (N_5506,N_5360,N_5395);
and U5507 (N_5507,N_5496,N_5388);
and U5508 (N_5508,N_5494,N_5433);
or U5509 (N_5509,N_5428,N_5353);
nor U5510 (N_5510,N_5293,N_5357);
and U5511 (N_5511,N_5465,N_5459);
nand U5512 (N_5512,N_5463,N_5475);
or U5513 (N_5513,N_5327,N_5362);
nand U5514 (N_5514,N_5471,N_5392);
nor U5515 (N_5515,N_5251,N_5447);
or U5516 (N_5516,N_5396,N_5374);
nand U5517 (N_5517,N_5253,N_5302);
and U5518 (N_5518,N_5371,N_5448);
and U5519 (N_5519,N_5477,N_5452);
or U5520 (N_5520,N_5323,N_5325);
and U5521 (N_5521,N_5339,N_5498);
and U5522 (N_5522,N_5282,N_5410);
and U5523 (N_5523,N_5430,N_5473);
xnor U5524 (N_5524,N_5378,N_5312);
nand U5525 (N_5525,N_5383,N_5466);
or U5526 (N_5526,N_5256,N_5286);
or U5527 (N_5527,N_5261,N_5435);
nor U5528 (N_5528,N_5338,N_5265);
xnor U5529 (N_5529,N_5270,N_5444);
and U5530 (N_5530,N_5390,N_5400);
or U5531 (N_5531,N_5429,N_5404);
nand U5532 (N_5532,N_5391,N_5263);
or U5533 (N_5533,N_5314,N_5277);
nand U5534 (N_5534,N_5385,N_5380);
and U5535 (N_5535,N_5469,N_5387);
or U5536 (N_5536,N_5460,N_5322);
nand U5537 (N_5537,N_5250,N_5446);
and U5538 (N_5538,N_5464,N_5260);
or U5539 (N_5539,N_5412,N_5491);
xor U5540 (N_5540,N_5299,N_5358);
nand U5541 (N_5541,N_5298,N_5375);
or U5542 (N_5542,N_5421,N_5406);
and U5543 (N_5543,N_5356,N_5458);
or U5544 (N_5544,N_5252,N_5402);
nor U5545 (N_5545,N_5397,N_5366);
xnor U5546 (N_5546,N_5438,N_5499);
nor U5547 (N_5547,N_5344,N_5326);
xor U5548 (N_5548,N_5275,N_5394);
or U5549 (N_5549,N_5484,N_5280);
nand U5550 (N_5550,N_5324,N_5285);
and U5551 (N_5551,N_5417,N_5329);
or U5552 (N_5552,N_5377,N_5398);
xor U5553 (N_5553,N_5443,N_5440);
or U5554 (N_5554,N_5311,N_5409);
xnor U5555 (N_5555,N_5363,N_5457);
nor U5556 (N_5556,N_5497,N_5381);
xnor U5557 (N_5557,N_5386,N_5268);
xnor U5558 (N_5558,N_5425,N_5328);
nand U5559 (N_5559,N_5482,N_5305);
nor U5560 (N_5560,N_5296,N_5492);
and U5561 (N_5561,N_5432,N_5373);
or U5562 (N_5562,N_5341,N_5257);
nor U5563 (N_5563,N_5369,N_5413);
xnor U5564 (N_5564,N_5309,N_5468);
nand U5565 (N_5565,N_5364,N_5442);
nand U5566 (N_5566,N_5345,N_5478);
and U5567 (N_5567,N_5331,N_5437);
or U5568 (N_5568,N_5283,N_5297);
nand U5569 (N_5569,N_5359,N_5476);
or U5570 (N_5570,N_5281,N_5354);
and U5571 (N_5571,N_5259,N_5407);
and U5572 (N_5572,N_5495,N_5267);
xor U5573 (N_5573,N_5271,N_5411);
xnor U5574 (N_5574,N_5401,N_5481);
nor U5575 (N_5575,N_5456,N_5287);
and U5576 (N_5576,N_5467,N_5372);
and U5577 (N_5577,N_5342,N_5337);
nand U5578 (N_5578,N_5278,N_5461);
or U5579 (N_5579,N_5262,N_5365);
nor U5580 (N_5580,N_5284,N_5431);
xnor U5581 (N_5581,N_5420,N_5451);
nor U5582 (N_5582,N_5436,N_5418);
xnor U5583 (N_5583,N_5303,N_5274);
xor U5584 (N_5584,N_5368,N_5399);
and U5585 (N_5585,N_5307,N_5351);
xor U5586 (N_5586,N_5454,N_5439);
nor U5587 (N_5587,N_5415,N_5474);
nand U5588 (N_5588,N_5319,N_5350);
xnor U5589 (N_5589,N_5288,N_5422);
nand U5590 (N_5590,N_5470,N_5352);
nor U5591 (N_5591,N_5347,N_5487);
or U5592 (N_5592,N_5434,N_5426);
nor U5593 (N_5593,N_5258,N_5306);
and U5594 (N_5594,N_5408,N_5349);
xnor U5595 (N_5595,N_5304,N_5320);
xnor U5596 (N_5596,N_5419,N_5295);
nand U5597 (N_5597,N_5493,N_5300);
and U5598 (N_5598,N_5379,N_5462);
and U5599 (N_5599,N_5318,N_5273);
and U5600 (N_5600,N_5301,N_5340);
nor U5601 (N_5601,N_5255,N_5441);
nor U5602 (N_5602,N_5480,N_5361);
nor U5603 (N_5603,N_5348,N_5272);
xnor U5604 (N_5604,N_5254,N_5290);
and U5605 (N_5605,N_5334,N_5427);
nand U5606 (N_5606,N_5330,N_5266);
and U5607 (N_5607,N_5310,N_5321);
nand U5608 (N_5608,N_5453,N_5424);
xnor U5609 (N_5609,N_5343,N_5355);
nor U5610 (N_5610,N_5455,N_5370);
xnor U5611 (N_5611,N_5333,N_5488);
nor U5612 (N_5612,N_5279,N_5479);
and U5613 (N_5613,N_5313,N_5449);
and U5614 (N_5614,N_5389,N_5289);
nor U5615 (N_5615,N_5291,N_5276);
xor U5616 (N_5616,N_5317,N_5382);
nand U5617 (N_5617,N_5414,N_5486);
xnor U5618 (N_5618,N_5472,N_5450);
or U5619 (N_5619,N_5445,N_5416);
nand U5620 (N_5620,N_5490,N_5423);
and U5621 (N_5621,N_5403,N_5393);
or U5622 (N_5622,N_5483,N_5367);
nand U5623 (N_5623,N_5489,N_5376);
nor U5624 (N_5624,N_5294,N_5332);
xnor U5625 (N_5625,N_5460,N_5323);
nand U5626 (N_5626,N_5256,N_5489);
or U5627 (N_5627,N_5322,N_5342);
and U5628 (N_5628,N_5327,N_5453);
or U5629 (N_5629,N_5358,N_5250);
and U5630 (N_5630,N_5409,N_5472);
xor U5631 (N_5631,N_5378,N_5431);
xor U5632 (N_5632,N_5391,N_5347);
nand U5633 (N_5633,N_5427,N_5408);
xor U5634 (N_5634,N_5339,N_5311);
or U5635 (N_5635,N_5399,N_5469);
or U5636 (N_5636,N_5298,N_5453);
or U5637 (N_5637,N_5347,N_5427);
nand U5638 (N_5638,N_5346,N_5282);
nand U5639 (N_5639,N_5440,N_5263);
nor U5640 (N_5640,N_5267,N_5358);
or U5641 (N_5641,N_5394,N_5296);
or U5642 (N_5642,N_5412,N_5440);
xnor U5643 (N_5643,N_5451,N_5448);
or U5644 (N_5644,N_5361,N_5279);
xor U5645 (N_5645,N_5458,N_5310);
nor U5646 (N_5646,N_5421,N_5378);
xnor U5647 (N_5647,N_5465,N_5379);
or U5648 (N_5648,N_5333,N_5294);
or U5649 (N_5649,N_5386,N_5318);
nor U5650 (N_5650,N_5315,N_5450);
nor U5651 (N_5651,N_5437,N_5424);
and U5652 (N_5652,N_5274,N_5441);
and U5653 (N_5653,N_5399,N_5405);
nor U5654 (N_5654,N_5469,N_5394);
and U5655 (N_5655,N_5442,N_5275);
or U5656 (N_5656,N_5280,N_5296);
nand U5657 (N_5657,N_5396,N_5325);
nand U5658 (N_5658,N_5312,N_5280);
nand U5659 (N_5659,N_5374,N_5295);
and U5660 (N_5660,N_5469,N_5479);
xor U5661 (N_5661,N_5360,N_5433);
nand U5662 (N_5662,N_5273,N_5296);
and U5663 (N_5663,N_5250,N_5289);
nor U5664 (N_5664,N_5376,N_5351);
and U5665 (N_5665,N_5367,N_5486);
nor U5666 (N_5666,N_5273,N_5431);
nand U5667 (N_5667,N_5338,N_5429);
xor U5668 (N_5668,N_5319,N_5345);
and U5669 (N_5669,N_5291,N_5364);
nor U5670 (N_5670,N_5469,N_5253);
nand U5671 (N_5671,N_5420,N_5356);
nor U5672 (N_5672,N_5448,N_5383);
or U5673 (N_5673,N_5395,N_5467);
nor U5674 (N_5674,N_5292,N_5468);
nor U5675 (N_5675,N_5278,N_5260);
or U5676 (N_5676,N_5386,N_5417);
or U5677 (N_5677,N_5471,N_5250);
xor U5678 (N_5678,N_5372,N_5364);
or U5679 (N_5679,N_5478,N_5359);
or U5680 (N_5680,N_5445,N_5272);
or U5681 (N_5681,N_5373,N_5433);
nand U5682 (N_5682,N_5475,N_5368);
xnor U5683 (N_5683,N_5391,N_5468);
nand U5684 (N_5684,N_5458,N_5304);
or U5685 (N_5685,N_5477,N_5280);
nor U5686 (N_5686,N_5372,N_5355);
nor U5687 (N_5687,N_5281,N_5309);
or U5688 (N_5688,N_5468,N_5382);
nand U5689 (N_5689,N_5321,N_5314);
xor U5690 (N_5690,N_5386,N_5270);
or U5691 (N_5691,N_5279,N_5374);
xnor U5692 (N_5692,N_5489,N_5367);
nand U5693 (N_5693,N_5398,N_5335);
or U5694 (N_5694,N_5493,N_5255);
xnor U5695 (N_5695,N_5465,N_5376);
and U5696 (N_5696,N_5331,N_5357);
xor U5697 (N_5697,N_5481,N_5273);
xnor U5698 (N_5698,N_5367,N_5394);
and U5699 (N_5699,N_5459,N_5334);
nand U5700 (N_5700,N_5436,N_5259);
nand U5701 (N_5701,N_5315,N_5348);
xor U5702 (N_5702,N_5351,N_5440);
nand U5703 (N_5703,N_5495,N_5370);
nand U5704 (N_5704,N_5362,N_5304);
xor U5705 (N_5705,N_5459,N_5497);
and U5706 (N_5706,N_5289,N_5308);
xor U5707 (N_5707,N_5421,N_5445);
and U5708 (N_5708,N_5443,N_5410);
nand U5709 (N_5709,N_5301,N_5366);
or U5710 (N_5710,N_5322,N_5296);
nand U5711 (N_5711,N_5472,N_5339);
or U5712 (N_5712,N_5426,N_5304);
xor U5713 (N_5713,N_5434,N_5493);
and U5714 (N_5714,N_5467,N_5266);
nor U5715 (N_5715,N_5468,N_5475);
nand U5716 (N_5716,N_5390,N_5367);
nand U5717 (N_5717,N_5421,N_5291);
xor U5718 (N_5718,N_5371,N_5436);
or U5719 (N_5719,N_5379,N_5259);
and U5720 (N_5720,N_5261,N_5257);
and U5721 (N_5721,N_5329,N_5425);
and U5722 (N_5722,N_5494,N_5261);
or U5723 (N_5723,N_5403,N_5467);
nor U5724 (N_5724,N_5313,N_5496);
or U5725 (N_5725,N_5468,N_5446);
or U5726 (N_5726,N_5339,N_5277);
and U5727 (N_5727,N_5413,N_5464);
and U5728 (N_5728,N_5304,N_5323);
and U5729 (N_5729,N_5315,N_5415);
and U5730 (N_5730,N_5453,N_5380);
nand U5731 (N_5731,N_5256,N_5453);
nand U5732 (N_5732,N_5400,N_5482);
nand U5733 (N_5733,N_5480,N_5331);
nand U5734 (N_5734,N_5378,N_5465);
and U5735 (N_5735,N_5490,N_5485);
nor U5736 (N_5736,N_5305,N_5324);
xor U5737 (N_5737,N_5407,N_5339);
and U5738 (N_5738,N_5368,N_5431);
xor U5739 (N_5739,N_5317,N_5421);
xnor U5740 (N_5740,N_5305,N_5431);
or U5741 (N_5741,N_5384,N_5319);
and U5742 (N_5742,N_5466,N_5274);
or U5743 (N_5743,N_5363,N_5326);
and U5744 (N_5744,N_5316,N_5301);
xnor U5745 (N_5745,N_5407,N_5328);
nor U5746 (N_5746,N_5322,N_5271);
nand U5747 (N_5747,N_5473,N_5333);
or U5748 (N_5748,N_5455,N_5498);
nand U5749 (N_5749,N_5314,N_5459);
xnor U5750 (N_5750,N_5678,N_5561);
and U5751 (N_5751,N_5579,N_5605);
xor U5752 (N_5752,N_5619,N_5748);
and U5753 (N_5753,N_5610,N_5556);
xnor U5754 (N_5754,N_5568,N_5730);
xnor U5755 (N_5755,N_5728,N_5576);
or U5756 (N_5756,N_5659,N_5512);
and U5757 (N_5757,N_5662,N_5712);
or U5758 (N_5758,N_5572,N_5502);
and U5759 (N_5759,N_5628,N_5669);
or U5760 (N_5760,N_5578,N_5672);
and U5761 (N_5761,N_5703,N_5675);
nand U5762 (N_5762,N_5646,N_5705);
and U5763 (N_5763,N_5639,N_5523);
and U5764 (N_5764,N_5559,N_5624);
xor U5765 (N_5765,N_5530,N_5671);
nor U5766 (N_5766,N_5501,N_5697);
nand U5767 (N_5767,N_5604,N_5535);
nand U5768 (N_5768,N_5707,N_5506);
xor U5769 (N_5769,N_5515,N_5749);
xnor U5770 (N_5770,N_5514,N_5590);
nand U5771 (N_5771,N_5700,N_5622);
nor U5772 (N_5772,N_5618,N_5731);
and U5773 (N_5773,N_5563,N_5743);
nand U5774 (N_5774,N_5607,N_5555);
xor U5775 (N_5775,N_5674,N_5653);
or U5776 (N_5776,N_5736,N_5541);
nand U5777 (N_5777,N_5591,N_5714);
or U5778 (N_5778,N_5596,N_5710);
xnor U5779 (N_5779,N_5740,N_5665);
and U5780 (N_5780,N_5742,N_5695);
nand U5781 (N_5781,N_5706,N_5529);
and U5782 (N_5782,N_5648,N_5533);
xnor U5783 (N_5783,N_5643,N_5650);
nor U5784 (N_5784,N_5676,N_5603);
nor U5785 (N_5785,N_5696,N_5597);
and U5786 (N_5786,N_5519,N_5633);
or U5787 (N_5787,N_5715,N_5593);
or U5788 (N_5788,N_5725,N_5525);
nand U5789 (N_5789,N_5554,N_5685);
nor U5790 (N_5790,N_5536,N_5682);
nor U5791 (N_5791,N_5513,N_5739);
nand U5792 (N_5792,N_5599,N_5557);
nand U5793 (N_5793,N_5687,N_5612);
nor U5794 (N_5794,N_5621,N_5652);
or U5795 (N_5795,N_5716,N_5719);
and U5796 (N_5796,N_5544,N_5588);
nand U5797 (N_5797,N_5699,N_5575);
or U5798 (N_5798,N_5562,N_5668);
nand U5799 (N_5799,N_5510,N_5524);
and U5800 (N_5800,N_5644,N_5690);
nor U5801 (N_5801,N_5522,N_5729);
nor U5802 (N_5802,N_5589,N_5573);
xnor U5803 (N_5803,N_5500,N_5616);
nor U5804 (N_5804,N_5738,N_5598);
and U5805 (N_5805,N_5645,N_5664);
and U5806 (N_5806,N_5571,N_5531);
nor U5807 (N_5807,N_5517,N_5611);
xor U5808 (N_5808,N_5595,N_5640);
nand U5809 (N_5809,N_5503,N_5688);
xor U5810 (N_5810,N_5704,N_5647);
and U5811 (N_5811,N_5508,N_5538);
nand U5812 (N_5812,N_5692,N_5606);
nor U5813 (N_5813,N_5733,N_5708);
nand U5814 (N_5814,N_5681,N_5587);
nand U5815 (N_5815,N_5574,N_5509);
xnor U5816 (N_5816,N_5521,N_5663);
xnor U5817 (N_5817,N_5564,N_5625);
and U5818 (N_5818,N_5582,N_5615);
nand U5819 (N_5819,N_5584,N_5693);
or U5820 (N_5820,N_5717,N_5694);
xnor U5821 (N_5821,N_5580,N_5721);
nor U5822 (N_5822,N_5569,N_5570);
and U5823 (N_5823,N_5601,N_5656);
nor U5824 (N_5824,N_5543,N_5632);
or U5825 (N_5825,N_5528,N_5637);
xnor U5826 (N_5826,N_5547,N_5548);
xor U5827 (N_5827,N_5747,N_5583);
or U5828 (N_5828,N_5642,N_5741);
nor U5829 (N_5829,N_5666,N_5702);
and U5830 (N_5830,N_5542,N_5722);
nor U5831 (N_5831,N_5660,N_5532);
nand U5832 (N_5832,N_5683,N_5627);
or U5833 (N_5833,N_5651,N_5586);
and U5834 (N_5834,N_5516,N_5581);
and U5835 (N_5835,N_5711,N_5511);
or U5836 (N_5836,N_5565,N_5585);
nand U5837 (N_5837,N_5677,N_5520);
nand U5838 (N_5838,N_5609,N_5623);
and U5839 (N_5839,N_5537,N_5608);
or U5840 (N_5840,N_5744,N_5701);
nand U5841 (N_5841,N_5558,N_5661);
or U5842 (N_5842,N_5600,N_5567);
nor U5843 (N_5843,N_5746,N_5551);
xor U5844 (N_5844,N_5505,N_5504);
nand U5845 (N_5845,N_5720,N_5620);
nor U5846 (N_5846,N_5641,N_5552);
nor U5847 (N_5847,N_5655,N_5686);
nor U5848 (N_5848,N_5654,N_5631);
and U5849 (N_5849,N_5592,N_5745);
nand U5850 (N_5850,N_5734,N_5539);
or U5851 (N_5851,N_5629,N_5732);
xnor U5852 (N_5852,N_5636,N_5737);
and U5853 (N_5853,N_5689,N_5649);
or U5854 (N_5854,N_5679,N_5614);
or U5855 (N_5855,N_5577,N_5709);
xor U5856 (N_5856,N_5684,N_5626);
nand U5857 (N_5857,N_5546,N_5518);
xnor U5858 (N_5858,N_5613,N_5507);
nor U5859 (N_5859,N_5723,N_5667);
or U5860 (N_5860,N_5534,N_5630);
xnor U5861 (N_5861,N_5594,N_5634);
nor U5862 (N_5862,N_5724,N_5566);
and U5863 (N_5863,N_5638,N_5540);
and U5864 (N_5864,N_5673,N_5553);
or U5865 (N_5865,N_5727,N_5718);
nand U5866 (N_5866,N_5670,N_5726);
nand U5867 (N_5867,N_5550,N_5549);
or U5868 (N_5868,N_5602,N_5680);
nand U5869 (N_5869,N_5635,N_5545);
and U5870 (N_5870,N_5658,N_5560);
and U5871 (N_5871,N_5657,N_5691);
and U5872 (N_5872,N_5527,N_5526);
or U5873 (N_5873,N_5713,N_5698);
or U5874 (N_5874,N_5617,N_5735);
nor U5875 (N_5875,N_5612,N_5663);
and U5876 (N_5876,N_5568,N_5588);
xnor U5877 (N_5877,N_5656,N_5696);
nor U5878 (N_5878,N_5528,N_5616);
nor U5879 (N_5879,N_5517,N_5658);
and U5880 (N_5880,N_5749,N_5747);
or U5881 (N_5881,N_5543,N_5708);
or U5882 (N_5882,N_5592,N_5646);
and U5883 (N_5883,N_5708,N_5598);
nand U5884 (N_5884,N_5586,N_5608);
xnor U5885 (N_5885,N_5595,N_5628);
or U5886 (N_5886,N_5518,N_5551);
nand U5887 (N_5887,N_5607,N_5695);
and U5888 (N_5888,N_5698,N_5602);
and U5889 (N_5889,N_5582,N_5689);
nor U5890 (N_5890,N_5571,N_5669);
nand U5891 (N_5891,N_5689,N_5679);
and U5892 (N_5892,N_5722,N_5530);
or U5893 (N_5893,N_5655,N_5601);
and U5894 (N_5894,N_5513,N_5672);
xor U5895 (N_5895,N_5614,N_5615);
and U5896 (N_5896,N_5588,N_5580);
nand U5897 (N_5897,N_5664,N_5690);
nand U5898 (N_5898,N_5537,N_5510);
nand U5899 (N_5899,N_5507,N_5666);
nor U5900 (N_5900,N_5662,N_5579);
and U5901 (N_5901,N_5590,N_5664);
or U5902 (N_5902,N_5689,N_5531);
nor U5903 (N_5903,N_5510,N_5555);
and U5904 (N_5904,N_5704,N_5651);
or U5905 (N_5905,N_5565,N_5504);
nand U5906 (N_5906,N_5695,N_5525);
nor U5907 (N_5907,N_5570,N_5511);
xnor U5908 (N_5908,N_5651,N_5747);
or U5909 (N_5909,N_5717,N_5566);
or U5910 (N_5910,N_5631,N_5706);
and U5911 (N_5911,N_5635,N_5552);
xnor U5912 (N_5912,N_5525,N_5606);
nor U5913 (N_5913,N_5521,N_5692);
and U5914 (N_5914,N_5584,N_5588);
nor U5915 (N_5915,N_5714,N_5659);
and U5916 (N_5916,N_5536,N_5613);
and U5917 (N_5917,N_5613,N_5582);
nand U5918 (N_5918,N_5717,N_5704);
nor U5919 (N_5919,N_5559,N_5595);
and U5920 (N_5920,N_5536,N_5606);
or U5921 (N_5921,N_5689,N_5719);
xor U5922 (N_5922,N_5737,N_5700);
or U5923 (N_5923,N_5503,N_5603);
xor U5924 (N_5924,N_5516,N_5745);
nor U5925 (N_5925,N_5557,N_5597);
or U5926 (N_5926,N_5537,N_5540);
nor U5927 (N_5927,N_5608,N_5542);
or U5928 (N_5928,N_5520,N_5629);
nand U5929 (N_5929,N_5740,N_5685);
nand U5930 (N_5930,N_5561,N_5638);
xor U5931 (N_5931,N_5692,N_5585);
nor U5932 (N_5932,N_5738,N_5639);
nand U5933 (N_5933,N_5538,N_5507);
nand U5934 (N_5934,N_5743,N_5616);
nand U5935 (N_5935,N_5672,N_5643);
xor U5936 (N_5936,N_5601,N_5583);
xnor U5937 (N_5937,N_5509,N_5683);
or U5938 (N_5938,N_5652,N_5616);
nor U5939 (N_5939,N_5717,N_5636);
nand U5940 (N_5940,N_5714,N_5618);
nand U5941 (N_5941,N_5524,N_5633);
and U5942 (N_5942,N_5744,N_5736);
nand U5943 (N_5943,N_5533,N_5573);
or U5944 (N_5944,N_5638,N_5549);
nand U5945 (N_5945,N_5647,N_5716);
nand U5946 (N_5946,N_5543,N_5551);
xnor U5947 (N_5947,N_5747,N_5582);
or U5948 (N_5948,N_5587,N_5543);
and U5949 (N_5949,N_5629,N_5652);
and U5950 (N_5950,N_5541,N_5654);
or U5951 (N_5951,N_5665,N_5534);
nor U5952 (N_5952,N_5677,N_5694);
xnor U5953 (N_5953,N_5633,N_5530);
nand U5954 (N_5954,N_5598,N_5683);
xnor U5955 (N_5955,N_5517,N_5686);
and U5956 (N_5956,N_5619,N_5733);
nor U5957 (N_5957,N_5639,N_5538);
nand U5958 (N_5958,N_5622,N_5707);
xnor U5959 (N_5959,N_5542,N_5532);
and U5960 (N_5960,N_5744,N_5604);
and U5961 (N_5961,N_5729,N_5722);
nand U5962 (N_5962,N_5665,N_5602);
xnor U5963 (N_5963,N_5633,N_5508);
or U5964 (N_5964,N_5641,N_5626);
xnor U5965 (N_5965,N_5538,N_5612);
nand U5966 (N_5966,N_5715,N_5577);
nor U5967 (N_5967,N_5560,N_5682);
nor U5968 (N_5968,N_5591,N_5635);
xor U5969 (N_5969,N_5721,N_5732);
nor U5970 (N_5970,N_5668,N_5592);
or U5971 (N_5971,N_5748,N_5749);
nor U5972 (N_5972,N_5721,N_5672);
nand U5973 (N_5973,N_5637,N_5538);
nor U5974 (N_5974,N_5687,N_5705);
or U5975 (N_5975,N_5699,N_5616);
xnor U5976 (N_5976,N_5579,N_5738);
nand U5977 (N_5977,N_5623,N_5640);
nand U5978 (N_5978,N_5658,N_5545);
nor U5979 (N_5979,N_5722,N_5598);
nor U5980 (N_5980,N_5696,N_5621);
or U5981 (N_5981,N_5699,N_5527);
and U5982 (N_5982,N_5663,N_5518);
nor U5983 (N_5983,N_5656,N_5527);
and U5984 (N_5984,N_5513,N_5650);
xor U5985 (N_5985,N_5623,N_5612);
nand U5986 (N_5986,N_5501,N_5619);
and U5987 (N_5987,N_5512,N_5549);
and U5988 (N_5988,N_5551,N_5668);
nor U5989 (N_5989,N_5510,N_5538);
xor U5990 (N_5990,N_5694,N_5513);
nor U5991 (N_5991,N_5654,N_5566);
xnor U5992 (N_5992,N_5540,N_5598);
or U5993 (N_5993,N_5699,N_5729);
xor U5994 (N_5994,N_5567,N_5656);
and U5995 (N_5995,N_5578,N_5682);
or U5996 (N_5996,N_5517,N_5564);
and U5997 (N_5997,N_5728,N_5652);
or U5998 (N_5998,N_5550,N_5666);
or U5999 (N_5999,N_5612,N_5521);
xnor U6000 (N_6000,N_5765,N_5782);
nor U6001 (N_6001,N_5931,N_5770);
and U6002 (N_6002,N_5975,N_5824);
nor U6003 (N_6003,N_5994,N_5844);
or U6004 (N_6004,N_5941,N_5860);
nor U6005 (N_6005,N_5968,N_5767);
nand U6006 (N_6006,N_5918,N_5810);
nand U6007 (N_6007,N_5884,N_5897);
nand U6008 (N_6008,N_5959,N_5754);
nand U6009 (N_6009,N_5958,N_5997);
or U6010 (N_6010,N_5816,N_5835);
nand U6011 (N_6011,N_5951,N_5890);
xor U6012 (N_6012,N_5867,N_5819);
nand U6013 (N_6013,N_5757,N_5928);
nand U6014 (N_6014,N_5783,N_5789);
or U6015 (N_6015,N_5984,N_5776);
nor U6016 (N_6016,N_5779,N_5962);
and U6017 (N_6017,N_5995,N_5854);
and U6018 (N_6018,N_5899,N_5905);
or U6019 (N_6019,N_5882,N_5880);
nor U6020 (N_6020,N_5980,N_5925);
and U6021 (N_6021,N_5977,N_5879);
nor U6022 (N_6022,N_5858,N_5887);
or U6023 (N_6023,N_5811,N_5986);
nand U6024 (N_6024,N_5937,N_5848);
nand U6025 (N_6025,N_5862,N_5885);
nand U6026 (N_6026,N_5839,N_5847);
nor U6027 (N_6027,N_5769,N_5881);
nand U6028 (N_6028,N_5909,N_5875);
nor U6029 (N_6029,N_5762,N_5932);
xor U6030 (N_6030,N_5976,N_5922);
nand U6031 (N_6031,N_5785,N_5952);
nand U6032 (N_6032,N_5773,N_5908);
xnor U6033 (N_6033,N_5828,N_5985);
or U6034 (N_6034,N_5948,N_5945);
and U6035 (N_6035,N_5912,N_5866);
xnor U6036 (N_6036,N_5953,N_5964);
or U6037 (N_6037,N_5838,N_5946);
nor U6038 (N_6038,N_5990,N_5938);
nand U6039 (N_6039,N_5916,N_5904);
nand U6040 (N_6040,N_5914,N_5841);
nand U6041 (N_6041,N_5772,N_5820);
and U6042 (N_6042,N_5944,N_5954);
nand U6043 (N_6043,N_5840,N_5771);
nand U6044 (N_6044,N_5949,N_5775);
nor U6045 (N_6045,N_5821,N_5751);
nor U6046 (N_6046,N_5943,N_5900);
nor U6047 (N_6047,N_5957,N_5855);
xor U6048 (N_6048,N_5935,N_5910);
nand U6049 (N_6049,N_5836,N_5996);
nor U6050 (N_6050,N_5788,N_5792);
and U6051 (N_6051,N_5876,N_5799);
or U6052 (N_6052,N_5791,N_5998);
nand U6053 (N_6053,N_5947,N_5973);
and U6054 (N_6054,N_5845,N_5795);
nand U6055 (N_6055,N_5872,N_5756);
xnor U6056 (N_6056,N_5920,N_5863);
and U6057 (N_6057,N_5934,N_5825);
nor U6058 (N_6058,N_5950,N_5780);
xor U6059 (N_6059,N_5803,N_5806);
and U6060 (N_6060,N_5774,N_5923);
and U6061 (N_6061,N_5978,N_5895);
and U6062 (N_6062,N_5817,N_5830);
nor U6063 (N_6063,N_5955,N_5873);
or U6064 (N_6064,N_5929,N_5768);
and U6065 (N_6065,N_5857,N_5896);
or U6066 (N_6066,N_5842,N_5750);
and U6067 (N_6067,N_5924,N_5898);
and U6068 (N_6068,N_5868,N_5906);
or U6069 (N_6069,N_5960,N_5870);
nand U6070 (N_6070,N_5759,N_5797);
nor U6071 (N_6071,N_5927,N_5888);
nor U6072 (N_6072,N_5861,N_5802);
nor U6073 (N_6073,N_5781,N_5970);
or U6074 (N_6074,N_5758,N_5911);
and U6075 (N_6075,N_5919,N_5966);
or U6076 (N_6076,N_5837,N_5972);
xor U6077 (N_6077,N_5917,N_5753);
and U6078 (N_6078,N_5760,N_5892);
nor U6079 (N_6079,N_5971,N_5859);
nor U6080 (N_6080,N_5823,N_5956);
and U6081 (N_6081,N_5999,N_5883);
nor U6082 (N_6082,N_5804,N_5874);
and U6083 (N_6083,N_5865,N_5913);
nor U6084 (N_6084,N_5807,N_5967);
xor U6085 (N_6085,N_5974,N_5798);
or U6086 (N_6086,N_5988,N_5989);
or U6087 (N_6087,N_5831,N_5983);
xnor U6088 (N_6088,N_5933,N_5815);
or U6089 (N_6089,N_5963,N_5778);
xnor U6090 (N_6090,N_5786,N_5982);
nand U6091 (N_6091,N_5961,N_5764);
and U6092 (N_6092,N_5921,N_5805);
nand U6093 (N_6093,N_5826,N_5777);
and U6094 (N_6094,N_5755,N_5833);
nand U6095 (N_6095,N_5987,N_5766);
and U6096 (N_6096,N_5940,N_5915);
or U6097 (N_6097,N_5851,N_5763);
and U6098 (N_6098,N_5832,N_5891);
nand U6099 (N_6099,N_5794,N_5992);
nor U6100 (N_6100,N_5864,N_5889);
xor U6101 (N_6101,N_5878,N_5856);
nor U6102 (N_6102,N_5834,N_5843);
xor U6103 (N_6103,N_5846,N_5849);
nor U6104 (N_6104,N_5813,N_5991);
and U6105 (N_6105,N_5829,N_5822);
xor U6106 (N_6106,N_5809,N_5853);
nor U6107 (N_6107,N_5942,N_5827);
and U6108 (N_6108,N_5893,N_5903);
xnor U6109 (N_6109,N_5808,N_5752);
nor U6110 (N_6110,N_5894,N_5850);
and U6111 (N_6111,N_5796,N_5793);
nor U6112 (N_6112,N_5993,N_5800);
nand U6113 (N_6113,N_5761,N_5981);
and U6114 (N_6114,N_5869,N_5907);
nor U6115 (N_6115,N_5979,N_5818);
nand U6116 (N_6116,N_5871,N_5969);
nand U6117 (N_6117,N_5801,N_5784);
nand U6118 (N_6118,N_5787,N_5939);
or U6119 (N_6119,N_5852,N_5790);
nand U6120 (N_6120,N_5965,N_5877);
and U6121 (N_6121,N_5930,N_5901);
nand U6122 (N_6122,N_5886,N_5814);
xnor U6123 (N_6123,N_5902,N_5926);
and U6124 (N_6124,N_5936,N_5812);
and U6125 (N_6125,N_5974,N_5994);
and U6126 (N_6126,N_5808,N_5905);
nand U6127 (N_6127,N_5852,N_5975);
xnor U6128 (N_6128,N_5764,N_5972);
and U6129 (N_6129,N_5819,N_5989);
or U6130 (N_6130,N_5915,N_5981);
nand U6131 (N_6131,N_5937,N_5946);
or U6132 (N_6132,N_5963,N_5945);
and U6133 (N_6133,N_5804,N_5818);
or U6134 (N_6134,N_5998,N_5782);
xor U6135 (N_6135,N_5843,N_5967);
nand U6136 (N_6136,N_5798,N_5786);
nor U6137 (N_6137,N_5829,N_5754);
nand U6138 (N_6138,N_5760,N_5862);
and U6139 (N_6139,N_5887,N_5865);
xnor U6140 (N_6140,N_5954,N_5753);
xor U6141 (N_6141,N_5806,N_5861);
nand U6142 (N_6142,N_5957,N_5780);
or U6143 (N_6143,N_5997,N_5943);
or U6144 (N_6144,N_5752,N_5984);
xor U6145 (N_6145,N_5804,N_5937);
nand U6146 (N_6146,N_5912,N_5914);
or U6147 (N_6147,N_5897,N_5877);
and U6148 (N_6148,N_5960,N_5832);
nand U6149 (N_6149,N_5863,N_5814);
nor U6150 (N_6150,N_5838,N_5925);
nand U6151 (N_6151,N_5812,N_5827);
nor U6152 (N_6152,N_5868,N_5858);
xnor U6153 (N_6153,N_5918,N_5935);
nor U6154 (N_6154,N_5797,N_5772);
xor U6155 (N_6155,N_5878,N_5896);
nand U6156 (N_6156,N_5967,N_5891);
nand U6157 (N_6157,N_5814,N_5961);
or U6158 (N_6158,N_5892,N_5864);
nand U6159 (N_6159,N_5896,N_5938);
xnor U6160 (N_6160,N_5988,N_5973);
nand U6161 (N_6161,N_5910,N_5827);
nand U6162 (N_6162,N_5872,N_5822);
and U6163 (N_6163,N_5828,N_5927);
or U6164 (N_6164,N_5962,N_5888);
or U6165 (N_6165,N_5863,N_5834);
or U6166 (N_6166,N_5854,N_5981);
and U6167 (N_6167,N_5983,N_5786);
nand U6168 (N_6168,N_5946,N_5886);
nor U6169 (N_6169,N_5825,N_5971);
or U6170 (N_6170,N_5942,N_5752);
or U6171 (N_6171,N_5931,N_5847);
and U6172 (N_6172,N_5800,N_5785);
nor U6173 (N_6173,N_5825,N_5897);
or U6174 (N_6174,N_5982,N_5905);
nand U6175 (N_6175,N_5892,N_5932);
nor U6176 (N_6176,N_5753,N_5980);
nand U6177 (N_6177,N_5955,N_5937);
or U6178 (N_6178,N_5765,N_5810);
or U6179 (N_6179,N_5793,N_5981);
and U6180 (N_6180,N_5892,N_5898);
nand U6181 (N_6181,N_5998,N_5986);
nand U6182 (N_6182,N_5898,N_5775);
and U6183 (N_6183,N_5839,N_5961);
nor U6184 (N_6184,N_5846,N_5997);
xnor U6185 (N_6185,N_5763,N_5988);
or U6186 (N_6186,N_5937,N_5929);
xnor U6187 (N_6187,N_5809,N_5808);
xor U6188 (N_6188,N_5865,N_5880);
nand U6189 (N_6189,N_5891,N_5976);
nor U6190 (N_6190,N_5778,N_5840);
or U6191 (N_6191,N_5879,N_5956);
and U6192 (N_6192,N_5883,N_5965);
and U6193 (N_6193,N_5759,N_5771);
and U6194 (N_6194,N_5959,N_5852);
and U6195 (N_6195,N_5827,N_5954);
nor U6196 (N_6196,N_5931,N_5906);
xnor U6197 (N_6197,N_5821,N_5966);
and U6198 (N_6198,N_5925,N_5853);
nor U6199 (N_6199,N_5869,N_5920);
and U6200 (N_6200,N_5800,N_5810);
or U6201 (N_6201,N_5946,N_5966);
xor U6202 (N_6202,N_5846,N_5882);
xnor U6203 (N_6203,N_5920,N_5924);
or U6204 (N_6204,N_5928,N_5915);
nand U6205 (N_6205,N_5995,N_5932);
xor U6206 (N_6206,N_5897,N_5752);
nand U6207 (N_6207,N_5924,N_5958);
and U6208 (N_6208,N_5809,N_5803);
nor U6209 (N_6209,N_5894,N_5819);
or U6210 (N_6210,N_5814,N_5903);
or U6211 (N_6211,N_5809,N_5835);
xor U6212 (N_6212,N_5865,N_5832);
and U6213 (N_6213,N_5938,N_5793);
nor U6214 (N_6214,N_5857,N_5908);
or U6215 (N_6215,N_5801,N_5864);
and U6216 (N_6216,N_5780,N_5880);
nand U6217 (N_6217,N_5987,N_5762);
nor U6218 (N_6218,N_5751,N_5840);
nor U6219 (N_6219,N_5762,N_5764);
or U6220 (N_6220,N_5806,N_5995);
or U6221 (N_6221,N_5812,N_5841);
nand U6222 (N_6222,N_5896,N_5970);
nand U6223 (N_6223,N_5827,N_5948);
nand U6224 (N_6224,N_5974,N_5857);
nand U6225 (N_6225,N_5974,N_5755);
and U6226 (N_6226,N_5761,N_5942);
nor U6227 (N_6227,N_5816,N_5858);
xor U6228 (N_6228,N_5916,N_5972);
nand U6229 (N_6229,N_5774,N_5878);
xnor U6230 (N_6230,N_5917,N_5895);
or U6231 (N_6231,N_5785,N_5849);
or U6232 (N_6232,N_5801,N_5958);
nand U6233 (N_6233,N_5931,N_5964);
nor U6234 (N_6234,N_5938,N_5897);
or U6235 (N_6235,N_5980,N_5882);
xnor U6236 (N_6236,N_5930,N_5989);
or U6237 (N_6237,N_5974,N_5896);
nor U6238 (N_6238,N_5925,N_5915);
or U6239 (N_6239,N_5991,N_5761);
or U6240 (N_6240,N_5776,N_5999);
xnor U6241 (N_6241,N_5931,N_5853);
xor U6242 (N_6242,N_5968,N_5883);
nand U6243 (N_6243,N_5998,N_5970);
xor U6244 (N_6244,N_5808,N_5794);
nand U6245 (N_6245,N_5833,N_5750);
nand U6246 (N_6246,N_5943,N_5851);
xnor U6247 (N_6247,N_5817,N_5876);
and U6248 (N_6248,N_5872,N_5810);
xor U6249 (N_6249,N_5958,N_5855);
nand U6250 (N_6250,N_6104,N_6123);
and U6251 (N_6251,N_6197,N_6051);
and U6252 (N_6252,N_6015,N_6194);
and U6253 (N_6253,N_6170,N_6085);
xnor U6254 (N_6254,N_6028,N_6007);
nand U6255 (N_6255,N_6176,N_6247);
nor U6256 (N_6256,N_6212,N_6069);
xor U6257 (N_6257,N_6137,N_6135);
nor U6258 (N_6258,N_6006,N_6206);
or U6259 (N_6259,N_6023,N_6149);
nand U6260 (N_6260,N_6025,N_6177);
nor U6261 (N_6261,N_6072,N_6046);
and U6262 (N_6262,N_6143,N_6211);
xor U6263 (N_6263,N_6110,N_6200);
nor U6264 (N_6264,N_6131,N_6218);
and U6265 (N_6265,N_6107,N_6093);
or U6266 (N_6266,N_6052,N_6002);
xnor U6267 (N_6267,N_6217,N_6117);
and U6268 (N_6268,N_6109,N_6153);
and U6269 (N_6269,N_6000,N_6036);
nor U6270 (N_6270,N_6095,N_6075);
nand U6271 (N_6271,N_6238,N_6103);
xnor U6272 (N_6272,N_6130,N_6113);
nor U6273 (N_6273,N_6210,N_6165);
or U6274 (N_6274,N_6189,N_6124);
or U6275 (N_6275,N_6078,N_6020);
nor U6276 (N_6276,N_6249,N_6061);
nand U6277 (N_6277,N_6196,N_6116);
and U6278 (N_6278,N_6019,N_6155);
xnor U6279 (N_6279,N_6048,N_6221);
nor U6280 (N_6280,N_6105,N_6239);
and U6281 (N_6281,N_6226,N_6160);
nand U6282 (N_6282,N_6074,N_6151);
xor U6283 (N_6283,N_6157,N_6219);
xor U6284 (N_6284,N_6142,N_6220);
and U6285 (N_6285,N_6232,N_6133);
or U6286 (N_6286,N_6144,N_6122);
nor U6287 (N_6287,N_6030,N_6039);
and U6288 (N_6288,N_6014,N_6027);
xor U6289 (N_6289,N_6156,N_6229);
or U6290 (N_6290,N_6008,N_6215);
nand U6291 (N_6291,N_6173,N_6204);
nor U6292 (N_6292,N_6018,N_6024);
nor U6293 (N_6293,N_6083,N_6089);
xnor U6294 (N_6294,N_6208,N_6161);
xor U6295 (N_6295,N_6081,N_6201);
and U6296 (N_6296,N_6047,N_6017);
nand U6297 (N_6297,N_6231,N_6240);
and U6298 (N_6298,N_6057,N_6022);
nor U6299 (N_6299,N_6064,N_6049);
nor U6300 (N_6300,N_6154,N_6066);
nor U6301 (N_6301,N_6132,N_6016);
xnor U6302 (N_6302,N_6235,N_6114);
or U6303 (N_6303,N_6106,N_6125);
and U6304 (N_6304,N_6062,N_6084);
nand U6305 (N_6305,N_6119,N_6077);
nand U6306 (N_6306,N_6096,N_6041);
nor U6307 (N_6307,N_6060,N_6207);
nand U6308 (N_6308,N_6168,N_6205);
or U6309 (N_6309,N_6091,N_6068);
nand U6310 (N_6310,N_6199,N_6134);
nand U6311 (N_6311,N_6053,N_6181);
or U6312 (N_6312,N_6045,N_6115);
or U6313 (N_6313,N_6070,N_6225);
xnor U6314 (N_6314,N_6237,N_6213);
or U6315 (N_6315,N_6005,N_6013);
and U6316 (N_6316,N_6166,N_6086);
or U6317 (N_6317,N_6080,N_6244);
and U6318 (N_6318,N_6245,N_6242);
nand U6319 (N_6319,N_6192,N_6152);
xnor U6320 (N_6320,N_6175,N_6073);
and U6321 (N_6321,N_6183,N_6021);
nor U6322 (N_6322,N_6128,N_6065);
or U6323 (N_6323,N_6230,N_6097);
xor U6324 (N_6324,N_6092,N_6146);
nand U6325 (N_6325,N_6040,N_6228);
nand U6326 (N_6326,N_6120,N_6010);
or U6327 (N_6327,N_6224,N_6079);
xnor U6328 (N_6328,N_6054,N_6167);
nand U6329 (N_6329,N_6108,N_6031);
nand U6330 (N_6330,N_6178,N_6184);
nand U6331 (N_6331,N_6004,N_6034);
nand U6332 (N_6332,N_6098,N_6187);
and U6333 (N_6333,N_6033,N_6140);
and U6334 (N_6334,N_6190,N_6129);
xnor U6335 (N_6335,N_6236,N_6101);
and U6336 (N_6336,N_6233,N_6246);
or U6337 (N_6337,N_6145,N_6026);
nor U6338 (N_6338,N_6141,N_6172);
and U6339 (N_6339,N_6100,N_6063);
nor U6340 (N_6340,N_6127,N_6058);
and U6341 (N_6341,N_6121,N_6009);
or U6342 (N_6342,N_6076,N_6223);
nand U6343 (N_6343,N_6186,N_6050);
nand U6344 (N_6344,N_6067,N_6227);
nor U6345 (N_6345,N_6112,N_6209);
xnor U6346 (N_6346,N_6243,N_6148);
or U6347 (N_6347,N_6032,N_6087);
xnor U6348 (N_6348,N_6164,N_6241);
and U6349 (N_6349,N_6003,N_6163);
or U6350 (N_6350,N_6012,N_6138);
nor U6351 (N_6351,N_6059,N_6248);
and U6352 (N_6352,N_6035,N_6195);
or U6353 (N_6353,N_6198,N_6222);
and U6354 (N_6354,N_6202,N_6162);
and U6355 (N_6355,N_6044,N_6011);
and U6356 (N_6356,N_6234,N_6056);
and U6357 (N_6357,N_6090,N_6185);
and U6358 (N_6358,N_6118,N_6203);
or U6359 (N_6359,N_6158,N_6180);
xor U6360 (N_6360,N_6038,N_6159);
xor U6361 (N_6361,N_6182,N_6029);
and U6362 (N_6362,N_6139,N_6169);
nand U6363 (N_6363,N_6071,N_6037);
nor U6364 (N_6364,N_6099,N_6193);
xor U6365 (N_6365,N_6082,N_6042);
xor U6366 (N_6366,N_6216,N_6191);
xor U6367 (N_6367,N_6001,N_6111);
nor U6368 (N_6368,N_6188,N_6214);
nand U6369 (N_6369,N_6147,N_6136);
nor U6370 (N_6370,N_6179,N_6174);
nor U6371 (N_6371,N_6102,N_6126);
and U6372 (N_6372,N_6094,N_6171);
xor U6373 (N_6373,N_6150,N_6043);
or U6374 (N_6374,N_6055,N_6088);
and U6375 (N_6375,N_6171,N_6009);
nand U6376 (N_6376,N_6086,N_6023);
xor U6377 (N_6377,N_6239,N_6110);
nor U6378 (N_6378,N_6192,N_6008);
and U6379 (N_6379,N_6150,N_6131);
and U6380 (N_6380,N_6123,N_6142);
and U6381 (N_6381,N_6083,N_6150);
or U6382 (N_6382,N_6197,N_6165);
and U6383 (N_6383,N_6154,N_6016);
nor U6384 (N_6384,N_6144,N_6057);
xnor U6385 (N_6385,N_6149,N_6123);
or U6386 (N_6386,N_6198,N_6192);
xnor U6387 (N_6387,N_6234,N_6058);
nor U6388 (N_6388,N_6081,N_6169);
nand U6389 (N_6389,N_6123,N_6140);
and U6390 (N_6390,N_6145,N_6092);
or U6391 (N_6391,N_6184,N_6189);
or U6392 (N_6392,N_6074,N_6178);
xnor U6393 (N_6393,N_6160,N_6086);
nand U6394 (N_6394,N_6173,N_6034);
nand U6395 (N_6395,N_6058,N_6160);
nand U6396 (N_6396,N_6070,N_6083);
nand U6397 (N_6397,N_6043,N_6111);
nor U6398 (N_6398,N_6017,N_6112);
nand U6399 (N_6399,N_6108,N_6213);
or U6400 (N_6400,N_6160,N_6076);
and U6401 (N_6401,N_6141,N_6012);
and U6402 (N_6402,N_6069,N_6093);
and U6403 (N_6403,N_6013,N_6014);
nor U6404 (N_6404,N_6124,N_6063);
or U6405 (N_6405,N_6234,N_6111);
or U6406 (N_6406,N_6102,N_6151);
and U6407 (N_6407,N_6142,N_6232);
nor U6408 (N_6408,N_6018,N_6208);
nand U6409 (N_6409,N_6019,N_6228);
xor U6410 (N_6410,N_6077,N_6029);
and U6411 (N_6411,N_6102,N_6113);
or U6412 (N_6412,N_6047,N_6093);
nor U6413 (N_6413,N_6153,N_6098);
or U6414 (N_6414,N_6182,N_6109);
nor U6415 (N_6415,N_6185,N_6087);
and U6416 (N_6416,N_6206,N_6209);
xnor U6417 (N_6417,N_6091,N_6062);
nor U6418 (N_6418,N_6245,N_6044);
and U6419 (N_6419,N_6186,N_6196);
or U6420 (N_6420,N_6182,N_6085);
nand U6421 (N_6421,N_6240,N_6183);
or U6422 (N_6422,N_6068,N_6076);
nor U6423 (N_6423,N_6015,N_6185);
or U6424 (N_6424,N_6050,N_6096);
nor U6425 (N_6425,N_6156,N_6220);
nor U6426 (N_6426,N_6028,N_6138);
and U6427 (N_6427,N_6238,N_6118);
xnor U6428 (N_6428,N_6083,N_6186);
or U6429 (N_6429,N_6239,N_6114);
nor U6430 (N_6430,N_6131,N_6110);
and U6431 (N_6431,N_6246,N_6114);
and U6432 (N_6432,N_6003,N_6046);
xnor U6433 (N_6433,N_6224,N_6057);
nand U6434 (N_6434,N_6135,N_6235);
nand U6435 (N_6435,N_6183,N_6176);
xnor U6436 (N_6436,N_6097,N_6192);
or U6437 (N_6437,N_6108,N_6151);
and U6438 (N_6438,N_6008,N_6006);
and U6439 (N_6439,N_6178,N_6051);
or U6440 (N_6440,N_6121,N_6019);
nand U6441 (N_6441,N_6184,N_6024);
xnor U6442 (N_6442,N_6146,N_6234);
and U6443 (N_6443,N_6094,N_6120);
nand U6444 (N_6444,N_6073,N_6212);
nand U6445 (N_6445,N_6217,N_6131);
or U6446 (N_6446,N_6028,N_6184);
and U6447 (N_6447,N_6156,N_6084);
or U6448 (N_6448,N_6102,N_6129);
xnor U6449 (N_6449,N_6051,N_6212);
nor U6450 (N_6450,N_6013,N_6065);
xor U6451 (N_6451,N_6019,N_6179);
or U6452 (N_6452,N_6006,N_6072);
and U6453 (N_6453,N_6229,N_6042);
and U6454 (N_6454,N_6038,N_6110);
nand U6455 (N_6455,N_6175,N_6180);
and U6456 (N_6456,N_6051,N_6089);
and U6457 (N_6457,N_6152,N_6197);
and U6458 (N_6458,N_6038,N_6027);
or U6459 (N_6459,N_6022,N_6207);
nand U6460 (N_6460,N_6140,N_6119);
or U6461 (N_6461,N_6059,N_6205);
xnor U6462 (N_6462,N_6114,N_6249);
nand U6463 (N_6463,N_6211,N_6188);
or U6464 (N_6464,N_6167,N_6145);
and U6465 (N_6465,N_6066,N_6091);
nand U6466 (N_6466,N_6001,N_6003);
nor U6467 (N_6467,N_6052,N_6202);
or U6468 (N_6468,N_6066,N_6164);
xnor U6469 (N_6469,N_6057,N_6163);
xnor U6470 (N_6470,N_6071,N_6181);
or U6471 (N_6471,N_6080,N_6135);
xnor U6472 (N_6472,N_6009,N_6101);
xnor U6473 (N_6473,N_6087,N_6103);
xnor U6474 (N_6474,N_6145,N_6056);
and U6475 (N_6475,N_6143,N_6008);
and U6476 (N_6476,N_6057,N_6132);
or U6477 (N_6477,N_6079,N_6188);
and U6478 (N_6478,N_6016,N_6010);
or U6479 (N_6479,N_6158,N_6008);
nor U6480 (N_6480,N_6108,N_6046);
and U6481 (N_6481,N_6106,N_6230);
or U6482 (N_6482,N_6205,N_6200);
xnor U6483 (N_6483,N_6145,N_6099);
xnor U6484 (N_6484,N_6003,N_6072);
and U6485 (N_6485,N_6114,N_6071);
nand U6486 (N_6486,N_6171,N_6029);
or U6487 (N_6487,N_6117,N_6226);
nor U6488 (N_6488,N_6114,N_6121);
nor U6489 (N_6489,N_6171,N_6064);
xnor U6490 (N_6490,N_6087,N_6100);
or U6491 (N_6491,N_6078,N_6029);
xor U6492 (N_6492,N_6072,N_6054);
and U6493 (N_6493,N_6204,N_6160);
nand U6494 (N_6494,N_6119,N_6097);
xnor U6495 (N_6495,N_6136,N_6194);
or U6496 (N_6496,N_6180,N_6161);
or U6497 (N_6497,N_6204,N_6163);
xnor U6498 (N_6498,N_6004,N_6037);
nor U6499 (N_6499,N_6224,N_6175);
or U6500 (N_6500,N_6444,N_6364);
nand U6501 (N_6501,N_6483,N_6353);
or U6502 (N_6502,N_6279,N_6386);
and U6503 (N_6503,N_6282,N_6498);
xor U6504 (N_6504,N_6251,N_6307);
and U6505 (N_6505,N_6427,N_6413);
xor U6506 (N_6506,N_6423,N_6267);
nor U6507 (N_6507,N_6417,N_6477);
nand U6508 (N_6508,N_6481,N_6390);
nand U6509 (N_6509,N_6297,N_6250);
xnor U6510 (N_6510,N_6499,N_6460);
nand U6511 (N_6511,N_6378,N_6440);
or U6512 (N_6512,N_6394,N_6470);
xnor U6513 (N_6513,N_6314,N_6327);
and U6514 (N_6514,N_6308,N_6495);
xor U6515 (N_6515,N_6450,N_6317);
nand U6516 (N_6516,N_6292,N_6332);
and U6517 (N_6517,N_6272,N_6309);
and U6518 (N_6518,N_6262,N_6346);
or U6519 (N_6519,N_6425,N_6428);
nor U6520 (N_6520,N_6438,N_6358);
nor U6521 (N_6521,N_6463,N_6263);
and U6522 (N_6522,N_6312,N_6357);
nor U6523 (N_6523,N_6414,N_6348);
nor U6524 (N_6524,N_6411,N_6393);
nor U6525 (N_6525,N_6431,N_6286);
nor U6526 (N_6526,N_6454,N_6328);
nand U6527 (N_6527,N_6435,N_6416);
and U6528 (N_6528,N_6374,N_6298);
xor U6529 (N_6529,N_6457,N_6274);
and U6530 (N_6530,N_6303,N_6410);
and U6531 (N_6531,N_6468,N_6420);
and U6532 (N_6532,N_6268,N_6379);
nand U6533 (N_6533,N_6255,N_6335);
and U6534 (N_6534,N_6306,N_6270);
xor U6535 (N_6535,N_6269,N_6402);
or U6536 (N_6536,N_6313,N_6344);
or U6537 (N_6537,N_6458,N_6372);
nor U6538 (N_6538,N_6322,N_6369);
xor U6539 (N_6539,N_6434,N_6259);
nor U6540 (N_6540,N_6293,N_6382);
nor U6541 (N_6541,N_6302,N_6461);
nor U6542 (N_6542,N_6253,N_6350);
or U6543 (N_6543,N_6287,N_6254);
nor U6544 (N_6544,N_6453,N_6479);
nor U6545 (N_6545,N_6349,N_6485);
xor U6546 (N_6546,N_6320,N_6490);
xnor U6547 (N_6547,N_6405,N_6432);
xor U6548 (N_6548,N_6278,N_6376);
nor U6549 (N_6549,N_6341,N_6387);
nand U6550 (N_6550,N_6447,N_6475);
or U6551 (N_6551,N_6354,N_6294);
and U6552 (N_6552,N_6482,N_6397);
or U6553 (N_6553,N_6265,N_6396);
xnor U6554 (N_6554,N_6283,N_6363);
or U6555 (N_6555,N_6340,N_6489);
xor U6556 (N_6556,N_6323,N_6399);
and U6557 (N_6557,N_6352,N_6424);
nand U6558 (N_6558,N_6439,N_6462);
nor U6559 (N_6559,N_6351,N_6452);
nand U6560 (N_6560,N_6456,N_6491);
nand U6561 (N_6561,N_6256,N_6449);
nor U6562 (N_6562,N_6448,N_6301);
nor U6563 (N_6563,N_6412,N_6472);
or U6564 (N_6564,N_6391,N_6258);
or U6565 (N_6565,N_6342,N_6260);
or U6566 (N_6566,N_6398,N_6331);
nand U6567 (N_6567,N_6471,N_6252);
and U6568 (N_6568,N_6257,N_6430);
nand U6569 (N_6569,N_6494,N_6336);
nand U6570 (N_6570,N_6326,N_6497);
nand U6571 (N_6571,N_6338,N_6362);
nand U6572 (N_6572,N_6486,N_6373);
or U6573 (N_6573,N_6296,N_6337);
nor U6574 (N_6574,N_6291,N_6377);
nor U6575 (N_6575,N_6464,N_6371);
or U6576 (N_6576,N_6421,N_6266);
nor U6577 (N_6577,N_6488,N_6264);
or U6578 (N_6578,N_6426,N_6492);
or U6579 (N_6579,N_6476,N_6310);
or U6580 (N_6580,N_6469,N_6392);
or U6581 (N_6581,N_6300,N_6415);
xnor U6582 (N_6582,N_6284,N_6408);
or U6583 (N_6583,N_6437,N_6370);
nand U6584 (N_6584,N_6318,N_6321);
nand U6585 (N_6585,N_6459,N_6277);
and U6586 (N_6586,N_6436,N_6389);
nand U6587 (N_6587,N_6484,N_6403);
nand U6588 (N_6588,N_6288,N_6289);
nand U6589 (N_6589,N_6455,N_6333);
nor U6590 (N_6590,N_6466,N_6409);
or U6591 (N_6591,N_6406,N_6445);
and U6592 (N_6592,N_6356,N_6330);
xnor U6593 (N_6593,N_6474,N_6271);
nand U6594 (N_6594,N_6365,N_6367);
and U6595 (N_6595,N_6443,N_6273);
nand U6596 (N_6596,N_6305,N_6366);
xnor U6597 (N_6597,N_6280,N_6325);
nand U6598 (N_6598,N_6276,N_6401);
xor U6599 (N_6599,N_6381,N_6343);
nand U6600 (N_6600,N_6429,N_6304);
and U6601 (N_6601,N_6319,N_6496);
nor U6602 (N_6602,N_6359,N_6290);
nor U6603 (N_6603,N_6311,N_6334);
or U6604 (N_6604,N_6329,N_6433);
or U6605 (N_6605,N_6487,N_6281);
nand U6606 (N_6606,N_6441,N_6395);
nand U6607 (N_6607,N_6361,N_6355);
nor U6608 (N_6608,N_6446,N_6275);
nand U6609 (N_6609,N_6375,N_6316);
nor U6610 (N_6610,N_6480,N_6418);
nand U6611 (N_6611,N_6339,N_6383);
xor U6612 (N_6612,N_6388,N_6384);
nor U6613 (N_6613,N_6324,N_6404);
nand U6614 (N_6614,N_6385,N_6261);
nor U6615 (N_6615,N_6473,N_6380);
xnor U6616 (N_6616,N_6360,N_6478);
or U6617 (N_6617,N_6407,N_6347);
xor U6618 (N_6618,N_6493,N_6368);
nor U6619 (N_6619,N_6295,N_6285);
or U6620 (N_6620,N_6345,N_6419);
and U6621 (N_6621,N_6442,N_6315);
xor U6622 (N_6622,N_6467,N_6422);
and U6623 (N_6623,N_6400,N_6299);
xor U6624 (N_6624,N_6451,N_6465);
nor U6625 (N_6625,N_6339,N_6394);
xnor U6626 (N_6626,N_6253,N_6264);
or U6627 (N_6627,N_6306,N_6298);
nor U6628 (N_6628,N_6298,N_6441);
nand U6629 (N_6629,N_6470,N_6351);
or U6630 (N_6630,N_6300,N_6344);
xor U6631 (N_6631,N_6495,N_6490);
xor U6632 (N_6632,N_6376,N_6454);
or U6633 (N_6633,N_6262,N_6426);
xor U6634 (N_6634,N_6313,N_6366);
nor U6635 (N_6635,N_6380,N_6250);
nor U6636 (N_6636,N_6302,N_6259);
or U6637 (N_6637,N_6273,N_6378);
or U6638 (N_6638,N_6252,N_6498);
or U6639 (N_6639,N_6412,N_6330);
nand U6640 (N_6640,N_6285,N_6416);
xnor U6641 (N_6641,N_6323,N_6341);
xnor U6642 (N_6642,N_6446,N_6426);
or U6643 (N_6643,N_6392,N_6458);
nand U6644 (N_6644,N_6435,N_6443);
nand U6645 (N_6645,N_6278,N_6466);
nor U6646 (N_6646,N_6411,N_6366);
xnor U6647 (N_6647,N_6382,N_6343);
or U6648 (N_6648,N_6255,N_6459);
or U6649 (N_6649,N_6323,N_6430);
nor U6650 (N_6650,N_6458,N_6268);
and U6651 (N_6651,N_6437,N_6299);
and U6652 (N_6652,N_6293,N_6278);
and U6653 (N_6653,N_6416,N_6478);
and U6654 (N_6654,N_6413,N_6488);
nand U6655 (N_6655,N_6432,N_6275);
or U6656 (N_6656,N_6497,N_6437);
nor U6657 (N_6657,N_6448,N_6354);
nand U6658 (N_6658,N_6427,N_6266);
nand U6659 (N_6659,N_6446,N_6274);
nor U6660 (N_6660,N_6279,N_6293);
xor U6661 (N_6661,N_6366,N_6464);
nor U6662 (N_6662,N_6420,N_6455);
and U6663 (N_6663,N_6261,N_6254);
or U6664 (N_6664,N_6267,N_6276);
or U6665 (N_6665,N_6252,N_6328);
and U6666 (N_6666,N_6416,N_6305);
xor U6667 (N_6667,N_6355,N_6461);
xor U6668 (N_6668,N_6342,N_6251);
or U6669 (N_6669,N_6275,N_6412);
xor U6670 (N_6670,N_6296,N_6341);
and U6671 (N_6671,N_6331,N_6317);
and U6672 (N_6672,N_6361,N_6484);
nor U6673 (N_6673,N_6256,N_6370);
nand U6674 (N_6674,N_6376,N_6317);
or U6675 (N_6675,N_6392,N_6491);
and U6676 (N_6676,N_6338,N_6430);
xnor U6677 (N_6677,N_6389,N_6280);
nor U6678 (N_6678,N_6331,N_6380);
xnor U6679 (N_6679,N_6460,N_6264);
nor U6680 (N_6680,N_6337,N_6372);
nor U6681 (N_6681,N_6432,N_6430);
nand U6682 (N_6682,N_6358,N_6382);
xnor U6683 (N_6683,N_6295,N_6453);
nor U6684 (N_6684,N_6369,N_6490);
or U6685 (N_6685,N_6469,N_6292);
and U6686 (N_6686,N_6481,N_6286);
nand U6687 (N_6687,N_6491,N_6411);
and U6688 (N_6688,N_6476,N_6338);
or U6689 (N_6689,N_6456,N_6413);
or U6690 (N_6690,N_6318,N_6465);
or U6691 (N_6691,N_6355,N_6283);
and U6692 (N_6692,N_6297,N_6444);
or U6693 (N_6693,N_6416,N_6297);
nand U6694 (N_6694,N_6337,N_6364);
or U6695 (N_6695,N_6498,N_6491);
nor U6696 (N_6696,N_6374,N_6316);
or U6697 (N_6697,N_6306,N_6350);
and U6698 (N_6698,N_6409,N_6274);
or U6699 (N_6699,N_6368,N_6287);
and U6700 (N_6700,N_6447,N_6405);
and U6701 (N_6701,N_6306,N_6264);
or U6702 (N_6702,N_6431,N_6463);
or U6703 (N_6703,N_6275,N_6420);
or U6704 (N_6704,N_6260,N_6281);
xnor U6705 (N_6705,N_6368,N_6333);
nor U6706 (N_6706,N_6485,N_6366);
nand U6707 (N_6707,N_6445,N_6291);
xnor U6708 (N_6708,N_6261,N_6258);
or U6709 (N_6709,N_6487,N_6402);
and U6710 (N_6710,N_6379,N_6404);
xnor U6711 (N_6711,N_6485,N_6396);
xnor U6712 (N_6712,N_6496,N_6289);
and U6713 (N_6713,N_6345,N_6277);
nand U6714 (N_6714,N_6285,N_6292);
nand U6715 (N_6715,N_6439,N_6326);
or U6716 (N_6716,N_6299,N_6259);
and U6717 (N_6717,N_6443,N_6293);
or U6718 (N_6718,N_6414,N_6298);
xor U6719 (N_6719,N_6402,N_6475);
and U6720 (N_6720,N_6307,N_6342);
or U6721 (N_6721,N_6493,N_6331);
or U6722 (N_6722,N_6447,N_6483);
and U6723 (N_6723,N_6334,N_6459);
or U6724 (N_6724,N_6307,N_6291);
xor U6725 (N_6725,N_6343,N_6499);
or U6726 (N_6726,N_6409,N_6483);
and U6727 (N_6727,N_6426,N_6294);
nand U6728 (N_6728,N_6271,N_6450);
nand U6729 (N_6729,N_6286,N_6386);
xor U6730 (N_6730,N_6376,N_6462);
nand U6731 (N_6731,N_6492,N_6311);
xnor U6732 (N_6732,N_6254,N_6470);
nand U6733 (N_6733,N_6293,N_6405);
nor U6734 (N_6734,N_6417,N_6393);
nand U6735 (N_6735,N_6271,N_6334);
nand U6736 (N_6736,N_6463,N_6399);
nor U6737 (N_6737,N_6261,N_6290);
nand U6738 (N_6738,N_6373,N_6398);
or U6739 (N_6739,N_6462,N_6357);
nand U6740 (N_6740,N_6409,N_6311);
xor U6741 (N_6741,N_6396,N_6291);
xnor U6742 (N_6742,N_6340,N_6428);
and U6743 (N_6743,N_6326,N_6399);
and U6744 (N_6744,N_6328,N_6457);
xor U6745 (N_6745,N_6468,N_6373);
nand U6746 (N_6746,N_6488,N_6317);
nand U6747 (N_6747,N_6499,N_6399);
or U6748 (N_6748,N_6487,N_6350);
nor U6749 (N_6749,N_6434,N_6483);
nor U6750 (N_6750,N_6696,N_6663);
and U6751 (N_6751,N_6748,N_6556);
nand U6752 (N_6752,N_6539,N_6693);
nand U6753 (N_6753,N_6522,N_6613);
nand U6754 (N_6754,N_6713,N_6698);
or U6755 (N_6755,N_6580,N_6731);
or U6756 (N_6756,N_6730,N_6528);
nor U6757 (N_6757,N_6557,N_6509);
or U6758 (N_6758,N_6559,N_6634);
nor U6759 (N_6759,N_6532,N_6664);
and U6760 (N_6760,N_6550,N_6629);
nor U6761 (N_6761,N_6563,N_6720);
and U6762 (N_6762,N_6655,N_6644);
xor U6763 (N_6763,N_6641,N_6501);
or U6764 (N_6764,N_6635,N_6598);
or U6765 (N_6765,N_6533,N_6735);
and U6766 (N_6766,N_6661,N_6685);
or U6767 (N_6767,N_6679,N_6706);
nor U6768 (N_6768,N_6619,N_6584);
and U6769 (N_6769,N_6723,N_6545);
nand U6770 (N_6770,N_6739,N_6627);
and U6771 (N_6771,N_6503,N_6636);
nand U6772 (N_6772,N_6659,N_6595);
xor U6773 (N_6773,N_6649,N_6587);
xor U6774 (N_6774,N_6538,N_6677);
nor U6775 (N_6775,N_6606,N_6570);
xnor U6776 (N_6776,N_6643,N_6589);
xnor U6777 (N_6777,N_6590,N_6702);
nand U6778 (N_6778,N_6530,N_6592);
or U6779 (N_6779,N_6583,N_6704);
nand U6780 (N_6780,N_6588,N_6535);
xnor U6781 (N_6781,N_6682,N_6692);
nor U6782 (N_6782,N_6608,N_6700);
nor U6783 (N_6783,N_6645,N_6746);
xor U6784 (N_6784,N_6604,N_6681);
or U6785 (N_6785,N_6551,N_6579);
xor U6786 (N_6786,N_6591,N_6732);
nand U6787 (N_6787,N_6654,N_6594);
nand U6788 (N_6788,N_6660,N_6582);
xnor U6789 (N_6789,N_6573,N_6615);
or U6790 (N_6790,N_6568,N_6712);
nor U6791 (N_6791,N_6741,N_6718);
xor U6792 (N_6792,N_6737,N_6564);
nand U6793 (N_6793,N_6736,N_6552);
nor U6794 (N_6794,N_6719,N_6734);
xnor U6795 (N_6795,N_6624,N_6724);
nor U6796 (N_6796,N_6558,N_6674);
or U6797 (N_6797,N_6716,N_6524);
and U6798 (N_6798,N_6531,N_6640);
nand U6799 (N_6799,N_6554,N_6586);
or U6800 (N_6800,N_6657,N_6646);
nor U6801 (N_6801,N_6676,N_6507);
xor U6802 (N_6802,N_6622,N_6516);
or U6803 (N_6803,N_6651,N_6658);
nor U6804 (N_6804,N_6717,N_6729);
or U6805 (N_6805,N_6733,N_6697);
xnor U6806 (N_6806,N_6614,N_6705);
or U6807 (N_6807,N_6596,N_6699);
nand U6808 (N_6808,N_6569,N_6662);
and U6809 (N_6809,N_6680,N_6725);
or U6810 (N_6810,N_6514,N_6576);
xor U6811 (N_6811,N_6581,N_6715);
or U6812 (N_6812,N_6525,N_6653);
or U6813 (N_6813,N_6638,N_6668);
and U6814 (N_6814,N_6609,N_6745);
xor U6815 (N_6815,N_6714,N_6572);
nand U6816 (N_6816,N_6728,N_6690);
nor U6817 (N_6817,N_6537,N_6630);
nand U6818 (N_6818,N_6722,N_6626);
nor U6819 (N_6819,N_6519,N_6749);
and U6820 (N_6820,N_6647,N_6505);
xnor U6821 (N_6821,N_6669,N_6665);
nand U6822 (N_6822,N_6546,N_6517);
and U6823 (N_6823,N_6541,N_6744);
and U6824 (N_6824,N_6628,N_6547);
and U6825 (N_6825,N_6510,N_6562);
or U6826 (N_6826,N_6597,N_6603);
xnor U6827 (N_6827,N_6708,N_6549);
nor U6828 (N_6828,N_6512,N_6555);
nor U6829 (N_6829,N_6540,N_6652);
and U6830 (N_6830,N_6574,N_6686);
nand U6831 (N_6831,N_6593,N_6632);
or U6832 (N_6832,N_6513,N_6600);
or U6833 (N_6833,N_6727,N_6648);
or U6834 (N_6834,N_6691,N_6740);
nand U6835 (N_6835,N_6553,N_6672);
xnor U6836 (N_6836,N_6601,N_6534);
and U6837 (N_6837,N_6667,N_6694);
nor U6838 (N_6838,N_6695,N_6504);
nor U6839 (N_6839,N_6738,N_6625);
and U6840 (N_6840,N_6709,N_6612);
or U6841 (N_6841,N_6683,N_6637);
or U6842 (N_6842,N_6571,N_6575);
nand U6843 (N_6843,N_6610,N_6605);
and U6844 (N_6844,N_6602,N_6618);
and U6845 (N_6845,N_6599,N_6567);
and U6846 (N_6846,N_6621,N_6560);
nand U6847 (N_6847,N_6526,N_6721);
nor U6848 (N_6848,N_6536,N_6616);
or U6849 (N_6849,N_6743,N_6515);
xor U6850 (N_6850,N_6561,N_6607);
and U6851 (N_6851,N_6543,N_6650);
xnor U6852 (N_6852,N_6675,N_6703);
nand U6853 (N_6853,N_6633,N_6502);
nor U6854 (N_6854,N_6711,N_6684);
xor U6855 (N_6855,N_6631,N_6639);
nand U6856 (N_6856,N_6707,N_6585);
xnor U6857 (N_6857,N_6620,N_6710);
nand U6858 (N_6858,N_6670,N_6542);
nor U6859 (N_6859,N_6566,N_6687);
and U6860 (N_6860,N_6617,N_6523);
nor U6861 (N_6861,N_6577,N_6521);
xor U6862 (N_6862,N_6506,N_6529);
and U6863 (N_6863,N_6527,N_6688);
and U6864 (N_6864,N_6656,N_6689);
nor U6865 (N_6865,N_6623,N_6611);
nand U6866 (N_6866,N_6671,N_6578);
or U6867 (N_6867,N_6518,N_6511);
xor U6868 (N_6868,N_6701,N_6520);
nand U6869 (N_6869,N_6565,N_6747);
or U6870 (N_6870,N_6508,N_6548);
nand U6871 (N_6871,N_6642,N_6666);
nor U6872 (N_6872,N_6742,N_6500);
nand U6873 (N_6873,N_6726,N_6673);
nor U6874 (N_6874,N_6544,N_6678);
xnor U6875 (N_6875,N_6729,N_6562);
or U6876 (N_6876,N_6546,N_6554);
xnor U6877 (N_6877,N_6553,N_6688);
or U6878 (N_6878,N_6637,N_6749);
or U6879 (N_6879,N_6540,N_6736);
nand U6880 (N_6880,N_6713,N_6586);
nor U6881 (N_6881,N_6536,N_6645);
and U6882 (N_6882,N_6502,N_6593);
and U6883 (N_6883,N_6703,N_6617);
and U6884 (N_6884,N_6519,N_6594);
and U6885 (N_6885,N_6602,N_6582);
nand U6886 (N_6886,N_6684,N_6525);
nand U6887 (N_6887,N_6735,N_6712);
nor U6888 (N_6888,N_6715,N_6652);
xor U6889 (N_6889,N_6708,N_6535);
xor U6890 (N_6890,N_6585,N_6638);
xnor U6891 (N_6891,N_6611,N_6747);
xnor U6892 (N_6892,N_6503,N_6652);
and U6893 (N_6893,N_6551,N_6528);
xor U6894 (N_6894,N_6577,N_6538);
xor U6895 (N_6895,N_6562,N_6509);
nor U6896 (N_6896,N_6569,N_6503);
nand U6897 (N_6897,N_6529,N_6572);
nor U6898 (N_6898,N_6696,N_6715);
or U6899 (N_6899,N_6726,N_6514);
nor U6900 (N_6900,N_6682,N_6627);
and U6901 (N_6901,N_6658,N_6590);
or U6902 (N_6902,N_6546,N_6503);
xor U6903 (N_6903,N_6711,N_6576);
nor U6904 (N_6904,N_6619,N_6727);
nand U6905 (N_6905,N_6550,N_6593);
nand U6906 (N_6906,N_6593,N_6635);
and U6907 (N_6907,N_6648,N_6589);
nor U6908 (N_6908,N_6549,N_6700);
xnor U6909 (N_6909,N_6706,N_6575);
nand U6910 (N_6910,N_6703,N_6700);
and U6911 (N_6911,N_6662,N_6680);
nand U6912 (N_6912,N_6613,N_6591);
nand U6913 (N_6913,N_6601,N_6624);
nor U6914 (N_6914,N_6603,N_6740);
xnor U6915 (N_6915,N_6549,N_6525);
or U6916 (N_6916,N_6681,N_6508);
or U6917 (N_6917,N_6541,N_6646);
nor U6918 (N_6918,N_6652,N_6592);
or U6919 (N_6919,N_6643,N_6504);
xnor U6920 (N_6920,N_6682,N_6622);
and U6921 (N_6921,N_6534,N_6714);
nand U6922 (N_6922,N_6559,N_6732);
or U6923 (N_6923,N_6514,N_6733);
or U6924 (N_6924,N_6688,N_6650);
or U6925 (N_6925,N_6561,N_6666);
and U6926 (N_6926,N_6604,N_6593);
and U6927 (N_6927,N_6522,N_6746);
nor U6928 (N_6928,N_6722,N_6521);
and U6929 (N_6929,N_6588,N_6681);
nand U6930 (N_6930,N_6515,N_6742);
or U6931 (N_6931,N_6664,N_6511);
and U6932 (N_6932,N_6517,N_6696);
and U6933 (N_6933,N_6690,N_6706);
xnor U6934 (N_6934,N_6602,N_6588);
or U6935 (N_6935,N_6653,N_6700);
and U6936 (N_6936,N_6633,N_6501);
or U6937 (N_6937,N_6573,N_6595);
or U6938 (N_6938,N_6682,N_6617);
nand U6939 (N_6939,N_6620,N_6575);
and U6940 (N_6940,N_6733,N_6661);
xor U6941 (N_6941,N_6555,N_6544);
xnor U6942 (N_6942,N_6616,N_6512);
nor U6943 (N_6943,N_6548,N_6670);
nand U6944 (N_6944,N_6636,N_6524);
and U6945 (N_6945,N_6685,N_6560);
or U6946 (N_6946,N_6653,N_6516);
and U6947 (N_6947,N_6543,N_6678);
and U6948 (N_6948,N_6524,N_6593);
nand U6949 (N_6949,N_6684,N_6526);
and U6950 (N_6950,N_6729,N_6722);
nand U6951 (N_6951,N_6736,N_6602);
or U6952 (N_6952,N_6505,N_6648);
or U6953 (N_6953,N_6592,N_6529);
and U6954 (N_6954,N_6735,N_6733);
and U6955 (N_6955,N_6688,N_6614);
nor U6956 (N_6956,N_6502,N_6671);
nand U6957 (N_6957,N_6693,N_6714);
nand U6958 (N_6958,N_6663,N_6662);
and U6959 (N_6959,N_6682,N_6542);
and U6960 (N_6960,N_6745,N_6728);
nand U6961 (N_6961,N_6674,N_6584);
and U6962 (N_6962,N_6680,N_6675);
or U6963 (N_6963,N_6516,N_6600);
or U6964 (N_6964,N_6597,N_6658);
nor U6965 (N_6965,N_6576,N_6528);
nor U6966 (N_6966,N_6733,N_6500);
nand U6967 (N_6967,N_6541,N_6505);
xnor U6968 (N_6968,N_6521,N_6736);
xor U6969 (N_6969,N_6720,N_6516);
nor U6970 (N_6970,N_6582,N_6588);
xnor U6971 (N_6971,N_6729,N_6714);
xor U6972 (N_6972,N_6537,N_6516);
nand U6973 (N_6973,N_6699,N_6591);
and U6974 (N_6974,N_6556,N_6524);
or U6975 (N_6975,N_6727,N_6716);
and U6976 (N_6976,N_6721,N_6588);
or U6977 (N_6977,N_6559,N_6676);
or U6978 (N_6978,N_6662,N_6737);
nor U6979 (N_6979,N_6580,N_6718);
xnor U6980 (N_6980,N_6504,N_6696);
and U6981 (N_6981,N_6542,N_6646);
and U6982 (N_6982,N_6713,N_6723);
nand U6983 (N_6983,N_6711,N_6669);
nand U6984 (N_6984,N_6625,N_6528);
nor U6985 (N_6985,N_6610,N_6634);
xor U6986 (N_6986,N_6686,N_6710);
and U6987 (N_6987,N_6695,N_6696);
nand U6988 (N_6988,N_6682,N_6693);
xnor U6989 (N_6989,N_6732,N_6544);
or U6990 (N_6990,N_6734,N_6627);
or U6991 (N_6991,N_6696,N_6713);
or U6992 (N_6992,N_6585,N_6594);
nor U6993 (N_6993,N_6695,N_6583);
nor U6994 (N_6994,N_6623,N_6539);
xnor U6995 (N_6995,N_6554,N_6704);
and U6996 (N_6996,N_6670,N_6523);
and U6997 (N_6997,N_6666,N_6558);
nor U6998 (N_6998,N_6512,N_6701);
or U6999 (N_6999,N_6516,N_6524);
or U7000 (N_7000,N_6983,N_6816);
nand U7001 (N_7001,N_6930,N_6825);
nor U7002 (N_7002,N_6975,N_6922);
or U7003 (N_7003,N_6818,N_6821);
or U7004 (N_7004,N_6974,N_6913);
nand U7005 (N_7005,N_6814,N_6887);
or U7006 (N_7006,N_6807,N_6938);
nand U7007 (N_7007,N_6968,N_6956);
and U7008 (N_7008,N_6836,N_6905);
or U7009 (N_7009,N_6986,N_6982);
nor U7010 (N_7010,N_6927,N_6962);
nor U7011 (N_7011,N_6969,N_6940);
or U7012 (N_7012,N_6912,N_6906);
and U7013 (N_7013,N_6880,N_6872);
xnor U7014 (N_7014,N_6848,N_6844);
and U7015 (N_7015,N_6754,N_6796);
nand U7016 (N_7016,N_6902,N_6841);
nand U7017 (N_7017,N_6901,N_6998);
xnor U7018 (N_7018,N_6935,N_6764);
xor U7019 (N_7019,N_6869,N_6950);
or U7020 (N_7020,N_6861,N_6772);
and U7021 (N_7021,N_6967,N_6862);
and U7022 (N_7022,N_6804,N_6839);
or U7023 (N_7023,N_6827,N_6881);
xor U7024 (N_7024,N_6971,N_6792);
and U7025 (N_7025,N_6769,N_6959);
nand U7026 (N_7026,N_6970,N_6801);
xor U7027 (N_7027,N_6882,N_6859);
nor U7028 (N_7028,N_6899,N_6832);
or U7029 (N_7029,N_6817,N_6911);
nand U7030 (N_7030,N_6794,N_6851);
nand U7031 (N_7031,N_6919,N_6991);
xnor U7032 (N_7032,N_6757,N_6802);
nand U7033 (N_7033,N_6842,N_6947);
xnor U7034 (N_7034,N_6763,N_6988);
nor U7035 (N_7035,N_6984,N_6907);
nor U7036 (N_7036,N_6820,N_6834);
or U7037 (N_7037,N_6830,N_6756);
nor U7038 (N_7038,N_6944,N_6918);
xnor U7039 (N_7039,N_6767,N_6948);
nor U7040 (N_7040,N_6897,N_6941);
or U7041 (N_7041,N_6992,N_6963);
or U7042 (N_7042,N_6780,N_6961);
xnor U7043 (N_7043,N_6789,N_6972);
nor U7044 (N_7044,N_6876,N_6783);
nor U7045 (N_7045,N_6752,N_6824);
nor U7046 (N_7046,N_6779,N_6893);
nor U7047 (N_7047,N_6954,N_6758);
nor U7048 (N_7048,N_6994,N_6822);
and U7049 (N_7049,N_6985,N_6823);
and U7050 (N_7050,N_6791,N_6955);
or U7051 (N_7051,N_6875,N_6939);
xnor U7052 (N_7052,N_6903,N_6815);
and U7053 (N_7053,N_6781,N_6840);
nor U7054 (N_7054,N_6966,N_6856);
xor U7055 (N_7055,N_6797,N_6803);
nand U7056 (N_7056,N_6999,N_6952);
nor U7057 (N_7057,N_6936,N_6790);
and U7058 (N_7058,N_6852,N_6760);
nor U7059 (N_7059,N_6981,N_6964);
nor U7060 (N_7060,N_6934,N_6879);
or U7061 (N_7061,N_6819,N_6900);
and U7062 (N_7062,N_6896,N_6965);
nand U7063 (N_7063,N_6920,N_6835);
nor U7064 (N_7064,N_6928,N_6909);
or U7065 (N_7065,N_6976,N_6854);
nand U7066 (N_7066,N_6843,N_6812);
xnor U7067 (N_7067,N_6751,N_6777);
nor U7068 (N_7068,N_6782,N_6793);
or U7069 (N_7069,N_6795,N_6951);
nand U7070 (N_7070,N_6785,N_6773);
and U7071 (N_7071,N_6877,N_6858);
or U7072 (N_7072,N_6786,N_6878);
xnor U7073 (N_7073,N_6933,N_6979);
and U7074 (N_7074,N_6813,N_6884);
nand U7075 (N_7075,N_6892,N_6995);
and U7076 (N_7076,N_6808,N_6904);
nor U7077 (N_7077,N_6778,N_6867);
xor U7078 (N_7078,N_6766,N_6921);
nor U7079 (N_7079,N_6868,N_6787);
xnor U7080 (N_7080,N_6949,N_6924);
or U7081 (N_7081,N_6768,N_6847);
or U7082 (N_7082,N_6925,N_6811);
xnor U7083 (N_7083,N_6857,N_6958);
xor U7084 (N_7084,N_6883,N_6957);
xor U7085 (N_7085,N_6891,N_6829);
nor U7086 (N_7086,N_6805,N_6863);
or U7087 (N_7087,N_6929,N_6826);
nor U7088 (N_7088,N_6810,N_6831);
and U7089 (N_7089,N_6889,N_6806);
nor U7090 (N_7090,N_6759,N_6917);
xor U7091 (N_7091,N_6864,N_6770);
xor U7092 (N_7092,N_6978,N_6946);
and U7093 (N_7093,N_6800,N_6845);
and U7094 (N_7094,N_6885,N_6865);
and U7095 (N_7095,N_6850,N_6890);
nand U7096 (N_7096,N_6870,N_6973);
nand U7097 (N_7097,N_6886,N_6788);
nand U7098 (N_7098,N_6915,N_6894);
nand U7099 (N_7099,N_6898,N_6943);
or U7100 (N_7100,N_6855,N_6838);
nand U7101 (N_7101,N_6833,N_6888);
or U7102 (N_7102,N_6873,N_6798);
and U7103 (N_7103,N_6799,N_6846);
or U7104 (N_7104,N_6942,N_6923);
and U7105 (N_7105,N_6753,N_6996);
nor U7106 (N_7106,N_6987,N_6916);
xor U7107 (N_7107,N_6910,N_6953);
xor U7108 (N_7108,N_6776,N_6932);
nor U7109 (N_7109,N_6871,N_6960);
nor U7110 (N_7110,N_6931,N_6849);
nand U7111 (N_7111,N_6945,N_6755);
or U7112 (N_7112,N_6914,N_6775);
and U7113 (N_7113,N_6874,N_6860);
and U7114 (N_7114,N_6853,N_6774);
or U7115 (N_7115,N_6784,N_6771);
or U7116 (N_7116,N_6990,N_6809);
and U7117 (N_7117,N_6993,N_6750);
xor U7118 (N_7118,N_6989,N_6866);
xor U7119 (N_7119,N_6977,N_6980);
xnor U7120 (N_7120,N_6762,N_6828);
and U7121 (N_7121,N_6908,N_6837);
and U7122 (N_7122,N_6761,N_6997);
nand U7123 (N_7123,N_6937,N_6926);
xor U7124 (N_7124,N_6895,N_6765);
nor U7125 (N_7125,N_6802,N_6928);
or U7126 (N_7126,N_6795,N_6952);
or U7127 (N_7127,N_6776,N_6753);
xor U7128 (N_7128,N_6865,N_6967);
nor U7129 (N_7129,N_6754,N_6827);
nand U7130 (N_7130,N_6918,N_6774);
or U7131 (N_7131,N_6895,N_6927);
nand U7132 (N_7132,N_6986,N_6896);
xnor U7133 (N_7133,N_6967,N_6837);
and U7134 (N_7134,N_6838,N_6975);
nor U7135 (N_7135,N_6763,N_6926);
nor U7136 (N_7136,N_6812,N_6835);
nand U7137 (N_7137,N_6906,N_6943);
xnor U7138 (N_7138,N_6887,N_6792);
nand U7139 (N_7139,N_6799,N_6937);
nand U7140 (N_7140,N_6808,N_6882);
nand U7141 (N_7141,N_6905,N_6927);
xnor U7142 (N_7142,N_6862,N_6764);
or U7143 (N_7143,N_6757,N_6949);
and U7144 (N_7144,N_6788,N_6894);
nand U7145 (N_7145,N_6901,N_6947);
and U7146 (N_7146,N_6963,N_6777);
xor U7147 (N_7147,N_6878,N_6971);
or U7148 (N_7148,N_6933,N_6946);
nand U7149 (N_7149,N_6884,N_6847);
nand U7150 (N_7150,N_6846,N_6969);
or U7151 (N_7151,N_6759,N_6900);
nor U7152 (N_7152,N_6942,N_6770);
xnor U7153 (N_7153,N_6985,N_6827);
and U7154 (N_7154,N_6920,N_6930);
xor U7155 (N_7155,N_6958,N_6833);
xor U7156 (N_7156,N_6993,N_6798);
xnor U7157 (N_7157,N_6943,N_6921);
nand U7158 (N_7158,N_6897,N_6958);
nor U7159 (N_7159,N_6945,N_6886);
nand U7160 (N_7160,N_6939,N_6849);
and U7161 (N_7161,N_6873,N_6913);
nor U7162 (N_7162,N_6987,N_6820);
or U7163 (N_7163,N_6790,N_6795);
xor U7164 (N_7164,N_6870,N_6763);
nor U7165 (N_7165,N_6903,N_6930);
or U7166 (N_7166,N_6798,N_6810);
nor U7167 (N_7167,N_6775,N_6843);
nor U7168 (N_7168,N_6805,N_6986);
and U7169 (N_7169,N_6969,N_6803);
xor U7170 (N_7170,N_6927,N_6909);
nand U7171 (N_7171,N_6882,N_6971);
nor U7172 (N_7172,N_6957,N_6960);
nand U7173 (N_7173,N_6988,N_6936);
xnor U7174 (N_7174,N_6965,N_6992);
nand U7175 (N_7175,N_6982,N_6772);
nand U7176 (N_7176,N_6876,N_6858);
nor U7177 (N_7177,N_6802,N_6821);
and U7178 (N_7178,N_6917,N_6945);
and U7179 (N_7179,N_6907,N_6860);
nor U7180 (N_7180,N_6974,N_6955);
nor U7181 (N_7181,N_6769,N_6932);
nor U7182 (N_7182,N_6905,N_6962);
nand U7183 (N_7183,N_6919,N_6987);
nor U7184 (N_7184,N_6876,N_6968);
xnor U7185 (N_7185,N_6790,N_6984);
or U7186 (N_7186,N_6817,N_6898);
and U7187 (N_7187,N_6800,N_6902);
xor U7188 (N_7188,N_6769,N_6775);
and U7189 (N_7189,N_6881,N_6784);
or U7190 (N_7190,N_6921,N_6901);
nor U7191 (N_7191,N_6795,N_6824);
nor U7192 (N_7192,N_6920,N_6902);
xnor U7193 (N_7193,N_6954,N_6830);
nand U7194 (N_7194,N_6777,N_6790);
and U7195 (N_7195,N_6903,N_6752);
nor U7196 (N_7196,N_6898,N_6864);
xor U7197 (N_7197,N_6819,N_6771);
xnor U7198 (N_7198,N_6828,N_6993);
xor U7199 (N_7199,N_6944,N_6992);
or U7200 (N_7200,N_6980,N_6966);
xor U7201 (N_7201,N_6814,N_6774);
nand U7202 (N_7202,N_6875,N_6924);
and U7203 (N_7203,N_6849,N_6801);
nand U7204 (N_7204,N_6942,N_6756);
and U7205 (N_7205,N_6961,N_6771);
nor U7206 (N_7206,N_6929,N_6847);
nor U7207 (N_7207,N_6985,N_6789);
nor U7208 (N_7208,N_6920,N_6839);
nor U7209 (N_7209,N_6832,N_6959);
and U7210 (N_7210,N_6992,N_6923);
or U7211 (N_7211,N_6970,N_6831);
and U7212 (N_7212,N_6836,N_6882);
or U7213 (N_7213,N_6970,N_6799);
nor U7214 (N_7214,N_6783,N_6871);
xor U7215 (N_7215,N_6971,N_6772);
or U7216 (N_7216,N_6971,N_6980);
and U7217 (N_7217,N_6771,N_6869);
and U7218 (N_7218,N_6936,N_6754);
nand U7219 (N_7219,N_6854,N_6827);
or U7220 (N_7220,N_6791,N_6810);
nand U7221 (N_7221,N_6969,N_6920);
xor U7222 (N_7222,N_6768,N_6937);
nor U7223 (N_7223,N_6769,N_6874);
nand U7224 (N_7224,N_6834,N_6784);
nand U7225 (N_7225,N_6751,N_6759);
or U7226 (N_7226,N_6777,N_6847);
nor U7227 (N_7227,N_6846,N_6889);
xor U7228 (N_7228,N_6923,N_6910);
xnor U7229 (N_7229,N_6853,N_6890);
and U7230 (N_7230,N_6984,N_6832);
xnor U7231 (N_7231,N_6844,N_6867);
xnor U7232 (N_7232,N_6761,N_6866);
or U7233 (N_7233,N_6809,N_6903);
nor U7234 (N_7234,N_6859,N_6759);
nor U7235 (N_7235,N_6979,N_6913);
xor U7236 (N_7236,N_6803,N_6891);
nand U7237 (N_7237,N_6794,N_6992);
nand U7238 (N_7238,N_6849,N_6817);
and U7239 (N_7239,N_6823,N_6794);
or U7240 (N_7240,N_6833,N_6752);
and U7241 (N_7241,N_6835,N_6768);
nand U7242 (N_7242,N_6816,N_6852);
xnor U7243 (N_7243,N_6977,N_6774);
and U7244 (N_7244,N_6775,N_6796);
and U7245 (N_7245,N_6992,N_6799);
xnor U7246 (N_7246,N_6792,N_6809);
and U7247 (N_7247,N_6932,N_6860);
nand U7248 (N_7248,N_6945,N_6994);
xor U7249 (N_7249,N_6867,N_6908);
or U7250 (N_7250,N_7143,N_7200);
or U7251 (N_7251,N_7189,N_7214);
nor U7252 (N_7252,N_7158,N_7083);
or U7253 (N_7253,N_7087,N_7166);
nand U7254 (N_7254,N_7058,N_7050);
and U7255 (N_7255,N_7119,N_7227);
and U7256 (N_7256,N_7246,N_7081);
or U7257 (N_7257,N_7192,N_7047);
xnor U7258 (N_7258,N_7066,N_7069);
xor U7259 (N_7259,N_7155,N_7024);
or U7260 (N_7260,N_7028,N_7009);
and U7261 (N_7261,N_7210,N_7106);
xnor U7262 (N_7262,N_7226,N_7188);
nand U7263 (N_7263,N_7000,N_7108);
nor U7264 (N_7264,N_7101,N_7062);
nor U7265 (N_7265,N_7146,N_7113);
nor U7266 (N_7266,N_7038,N_7104);
nand U7267 (N_7267,N_7126,N_7036);
or U7268 (N_7268,N_7079,N_7071);
nand U7269 (N_7269,N_7234,N_7048);
xor U7270 (N_7270,N_7130,N_7098);
or U7271 (N_7271,N_7173,N_7135);
or U7272 (N_7272,N_7212,N_7154);
xnor U7273 (N_7273,N_7010,N_7195);
nand U7274 (N_7274,N_7008,N_7114);
nand U7275 (N_7275,N_7110,N_7190);
xnor U7276 (N_7276,N_7027,N_7142);
xor U7277 (N_7277,N_7165,N_7172);
nor U7278 (N_7278,N_7181,N_7039);
xor U7279 (N_7279,N_7128,N_7199);
and U7280 (N_7280,N_7141,N_7070);
xor U7281 (N_7281,N_7046,N_7120);
nor U7282 (N_7282,N_7231,N_7076);
and U7283 (N_7283,N_7103,N_7015);
or U7284 (N_7284,N_7249,N_7012);
or U7285 (N_7285,N_7137,N_7073);
and U7286 (N_7286,N_7037,N_7213);
nand U7287 (N_7287,N_7068,N_7170);
or U7288 (N_7288,N_7162,N_7171);
or U7289 (N_7289,N_7156,N_7018);
nand U7290 (N_7290,N_7053,N_7030);
or U7291 (N_7291,N_7096,N_7121);
nor U7292 (N_7292,N_7093,N_7014);
nor U7293 (N_7293,N_7125,N_7177);
nor U7294 (N_7294,N_7031,N_7085);
xnor U7295 (N_7295,N_7095,N_7224);
xor U7296 (N_7296,N_7075,N_7034);
nor U7297 (N_7297,N_7094,N_7232);
nand U7298 (N_7298,N_7149,N_7218);
nor U7299 (N_7299,N_7033,N_7049);
nor U7300 (N_7300,N_7145,N_7205);
and U7301 (N_7301,N_7057,N_7140);
xor U7302 (N_7302,N_7164,N_7060);
nor U7303 (N_7303,N_7107,N_7240);
or U7304 (N_7304,N_7115,N_7211);
and U7305 (N_7305,N_7241,N_7132);
nand U7306 (N_7306,N_7157,N_7002);
nor U7307 (N_7307,N_7202,N_7196);
or U7308 (N_7308,N_7163,N_7019);
and U7309 (N_7309,N_7061,N_7133);
or U7310 (N_7310,N_7221,N_7151);
nand U7311 (N_7311,N_7029,N_7016);
nand U7312 (N_7312,N_7204,N_7021);
nor U7313 (N_7313,N_7099,N_7007);
or U7314 (N_7314,N_7032,N_7111);
nor U7315 (N_7315,N_7243,N_7208);
xnor U7316 (N_7316,N_7160,N_7187);
nor U7317 (N_7317,N_7091,N_7242);
or U7318 (N_7318,N_7131,N_7116);
and U7319 (N_7319,N_7040,N_7178);
or U7320 (N_7320,N_7084,N_7223);
or U7321 (N_7321,N_7063,N_7138);
nand U7322 (N_7322,N_7123,N_7059);
and U7323 (N_7323,N_7092,N_7219);
nor U7324 (N_7324,N_7136,N_7052);
and U7325 (N_7325,N_7127,N_7097);
nand U7326 (N_7326,N_7100,N_7051);
xor U7327 (N_7327,N_7023,N_7167);
nand U7328 (N_7328,N_7198,N_7239);
nand U7329 (N_7329,N_7230,N_7174);
nor U7330 (N_7330,N_7089,N_7194);
and U7331 (N_7331,N_7011,N_7112);
nor U7332 (N_7332,N_7054,N_7080);
and U7333 (N_7333,N_7055,N_7176);
nand U7334 (N_7334,N_7229,N_7105);
or U7335 (N_7335,N_7025,N_7102);
nand U7336 (N_7336,N_7004,N_7139);
xor U7337 (N_7337,N_7245,N_7026);
nand U7338 (N_7338,N_7074,N_7185);
nand U7339 (N_7339,N_7045,N_7238);
nand U7340 (N_7340,N_7086,N_7179);
nor U7341 (N_7341,N_7216,N_7041);
or U7342 (N_7342,N_7042,N_7072);
and U7343 (N_7343,N_7077,N_7244);
nor U7344 (N_7344,N_7022,N_7090);
nand U7345 (N_7345,N_7109,N_7043);
nor U7346 (N_7346,N_7152,N_7215);
and U7347 (N_7347,N_7056,N_7191);
or U7348 (N_7348,N_7206,N_7193);
nand U7349 (N_7349,N_7235,N_7169);
nor U7350 (N_7350,N_7129,N_7201);
nor U7351 (N_7351,N_7236,N_7067);
and U7352 (N_7352,N_7197,N_7186);
nand U7353 (N_7353,N_7209,N_7150);
nor U7354 (N_7354,N_7225,N_7147);
xor U7355 (N_7355,N_7044,N_7159);
and U7356 (N_7356,N_7220,N_7001);
nor U7357 (N_7357,N_7153,N_7088);
or U7358 (N_7358,N_7124,N_7134);
xnor U7359 (N_7359,N_7005,N_7168);
and U7360 (N_7360,N_7222,N_7065);
nand U7361 (N_7361,N_7233,N_7182);
xnor U7362 (N_7362,N_7161,N_7082);
or U7363 (N_7363,N_7247,N_7248);
xor U7364 (N_7364,N_7122,N_7013);
and U7365 (N_7365,N_7144,N_7203);
nor U7366 (N_7366,N_7117,N_7020);
nand U7367 (N_7367,N_7237,N_7184);
or U7368 (N_7368,N_7183,N_7175);
and U7369 (N_7369,N_7217,N_7017);
nor U7370 (N_7370,N_7003,N_7228);
or U7371 (N_7371,N_7148,N_7118);
nor U7372 (N_7372,N_7035,N_7078);
nor U7373 (N_7373,N_7006,N_7064);
or U7374 (N_7374,N_7207,N_7180);
nand U7375 (N_7375,N_7209,N_7027);
or U7376 (N_7376,N_7211,N_7077);
xnor U7377 (N_7377,N_7001,N_7248);
and U7378 (N_7378,N_7054,N_7095);
nor U7379 (N_7379,N_7098,N_7025);
nor U7380 (N_7380,N_7039,N_7121);
xnor U7381 (N_7381,N_7024,N_7013);
and U7382 (N_7382,N_7107,N_7249);
nand U7383 (N_7383,N_7173,N_7046);
or U7384 (N_7384,N_7092,N_7075);
and U7385 (N_7385,N_7151,N_7131);
and U7386 (N_7386,N_7152,N_7168);
or U7387 (N_7387,N_7004,N_7113);
or U7388 (N_7388,N_7134,N_7073);
xor U7389 (N_7389,N_7172,N_7168);
xor U7390 (N_7390,N_7013,N_7035);
and U7391 (N_7391,N_7171,N_7224);
nand U7392 (N_7392,N_7023,N_7104);
or U7393 (N_7393,N_7124,N_7207);
xor U7394 (N_7394,N_7151,N_7227);
and U7395 (N_7395,N_7105,N_7015);
or U7396 (N_7396,N_7073,N_7064);
and U7397 (N_7397,N_7133,N_7062);
nand U7398 (N_7398,N_7226,N_7037);
nor U7399 (N_7399,N_7100,N_7080);
nor U7400 (N_7400,N_7121,N_7046);
nand U7401 (N_7401,N_7045,N_7027);
nand U7402 (N_7402,N_7173,N_7219);
nand U7403 (N_7403,N_7140,N_7064);
or U7404 (N_7404,N_7188,N_7185);
xor U7405 (N_7405,N_7243,N_7151);
nand U7406 (N_7406,N_7239,N_7117);
nor U7407 (N_7407,N_7070,N_7246);
and U7408 (N_7408,N_7221,N_7229);
or U7409 (N_7409,N_7192,N_7202);
and U7410 (N_7410,N_7067,N_7035);
and U7411 (N_7411,N_7069,N_7004);
or U7412 (N_7412,N_7101,N_7233);
or U7413 (N_7413,N_7043,N_7147);
and U7414 (N_7414,N_7139,N_7191);
nand U7415 (N_7415,N_7122,N_7111);
and U7416 (N_7416,N_7190,N_7117);
nand U7417 (N_7417,N_7023,N_7066);
nor U7418 (N_7418,N_7215,N_7062);
and U7419 (N_7419,N_7215,N_7202);
xnor U7420 (N_7420,N_7205,N_7017);
xor U7421 (N_7421,N_7020,N_7177);
nand U7422 (N_7422,N_7070,N_7056);
and U7423 (N_7423,N_7235,N_7074);
and U7424 (N_7424,N_7152,N_7123);
or U7425 (N_7425,N_7040,N_7028);
or U7426 (N_7426,N_7052,N_7049);
xor U7427 (N_7427,N_7222,N_7005);
and U7428 (N_7428,N_7049,N_7146);
nand U7429 (N_7429,N_7088,N_7104);
nand U7430 (N_7430,N_7002,N_7134);
nor U7431 (N_7431,N_7087,N_7067);
xnor U7432 (N_7432,N_7165,N_7018);
or U7433 (N_7433,N_7089,N_7116);
nand U7434 (N_7434,N_7206,N_7059);
nor U7435 (N_7435,N_7050,N_7247);
nor U7436 (N_7436,N_7232,N_7218);
or U7437 (N_7437,N_7160,N_7175);
nor U7438 (N_7438,N_7065,N_7245);
nand U7439 (N_7439,N_7152,N_7228);
nand U7440 (N_7440,N_7058,N_7214);
xor U7441 (N_7441,N_7013,N_7061);
and U7442 (N_7442,N_7206,N_7242);
or U7443 (N_7443,N_7211,N_7188);
nor U7444 (N_7444,N_7124,N_7144);
or U7445 (N_7445,N_7129,N_7127);
xnor U7446 (N_7446,N_7085,N_7197);
and U7447 (N_7447,N_7204,N_7066);
nand U7448 (N_7448,N_7072,N_7045);
nand U7449 (N_7449,N_7041,N_7112);
nand U7450 (N_7450,N_7111,N_7126);
nand U7451 (N_7451,N_7080,N_7229);
or U7452 (N_7452,N_7127,N_7002);
and U7453 (N_7453,N_7142,N_7108);
or U7454 (N_7454,N_7020,N_7228);
or U7455 (N_7455,N_7116,N_7041);
nor U7456 (N_7456,N_7033,N_7085);
nor U7457 (N_7457,N_7110,N_7127);
and U7458 (N_7458,N_7113,N_7074);
nor U7459 (N_7459,N_7227,N_7123);
nand U7460 (N_7460,N_7185,N_7248);
and U7461 (N_7461,N_7008,N_7077);
xnor U7462 (N_7462,N_7132,N_7066);
xor U7463 (N_7463,N_7171,N_7090);
or U7464 (N_7464,N_7067,N_7001);
xor U7465 (N_7465,N_7002,N_7125);
or U7466 (N_7466,N_7179,N_7171);
xor U7467 (N_7467,N_7172,N_7241);
xnor U7468 (N_7468,N_7000,N_7225);
nand U7469 (N_7469,N_7114,N_7097);
and U7470 (N_7470,N_7037,N_7215);
nand U7471 (N_7471,N_7169,N_7145);
and U7472 (N_7472,N_7008,N_7229);
and U7473 (N_7473,N_7200,N_7191);
nand U7474 (N_7474,N_7216,N_7219);
xor U7475 (N_7475,N_7018,N_7002);
and U7476 (N_7476,N_7023,N_7078);
nand U7477 (N_7477,N_7175,N_7218);
nand U7478 (N_7478,N_7143,N_7163);
nor U7479 (N_7479,N_7244,N_7049);
nor U7480 (N_7480,N_7140,N_7213);
and U7481 (N_7481,N_7023,N_7192);
and U7482 (N_7482,N_7155,N_7223);
and U7483 (N_7483,N_7217,N_7076);
nand U7484 (N_7484,N_7146,N_7153);
nor U7485 (N_7485,N_7044,N_7047);
nand U7486 (N_7486,N_7077,N_7084);
xnor U7487 (N_7487,N_7192,N_7141);
nand U7488 (N_7488,N_7004,N_7016);
or U7489 (N_7489,N_7105,N_7052);
and U7490 (N_7490,N_7153,N_7205);
nor U7491 (N_7491,N_7106,N_7003);
nand U7492 (N_7492,N_7002,N_7061);
xnor U7493 (N_7493,N_7037,N_7219);
or U7494 (N_7494,N_7170,N_7084);
nor U7495 (N_7495,N_7092,N_7214);
nor U7496 (N_7496,N_7208,N_7197);
nand U7497 (N_7497,N_7161,N_7174);
xnor U7498 (N_7498,N_7181,N_7234);
or U7499 (N_7499,N_7013,N_7145);
xnor U7500 (N_7500,N_7428,N_7361);
and U7501 (N_7501,N_7282,N_7319);
nor U7502 (N_7502,N_7301,N_7337);
xor U7503 (N_7503,N_7492,N_7265);
xnor U7504 (N_7504,N_7408,N_7332);
nor U7505 (N_7505,N_7486,N_7497);
xnor U7506 (N_7506,N_7298,N_7485);
and U7507 (N_7507,N_7254,N_7297);
and U7508 (N_7508,N_7334,N_7461);
or U7509 (N_7509,N_7272,N_7382);
or U7510 (N_7510,N_7451,N_7316);
xnor U7511 (N_7511,N_7406,N_7324);
or U7512 (N_7512,N_7362,N_7420);
nor U7513 (N_7513,N_7251,N_7394);
nor U7514 (N_7514,N_7453,N_7466);
nor U7515 (N_7515,N_7289,N_7437);
and U7516 (N_7516,N_7402,N_7360);
xor U7517 (N_7517,N_7442,N_7400);
or U7518 (N_7518,N_7284,N_7373);
and U7519 (N_7519,N_7342,N_7339);
and U7520 (N_7520,N_7388,N_7318);
or U7521 (N_7521,N_7354,N_7260);
nor U7522 (N_7522,N_7315,N_7412);
xnor U7523 (N_7523,N_7276,N_7454);
nor U7524 (N_7524,N_7398,N_7407);
and U7525 (N_7525,N_7317,N_7474);
nand U7526 (N_7526,N_7422,N_7498);
xnor U7527 (N_7527,N_7445,N_7396);
xnor U7528 (N_7528,N_7264,N_7329);
or U7529 (N_7529,N_7425,N_7262);
nand U7530 (N_7530,N_7424,N_7462);
xnor U7531 (N_7531,N_7326,N_7415);
or U7532 (N_7532,N_7472,N_7393);
and U7533 (N_7533,N_7447,N_7335);
or U7534 (N_7534,N_7482,N_7391);
nand U7535 (N_7535,N_7411,N_7353);
or U7536 (N_7536,N_7488,N_7293);
nand U7537 (N_7537,N_7433,N_7446);
xor U7538 (N_7538,N_7387,N_7292);
and U7539 (N_7539,N_7345,N_7325);
nand U7540 (N_7540,N_7493,N_7385);
nand U7541 (N_7541,N_7307,N_7371);
or U7542 (N_7542,N_7258,N_7463);
or U7543 (N_7543,N_7304,N_7357);
nand U7544 (N_7544,N_7489,N_7495);
or U7545 (N_7545,N_7351,N_7464);
nor U7546 (N_7546,N_7255,N_7367);
and U7547 (N_7547,N_7392,N_7384);
nand U7548 (N_7548,N_7323,N_7491);
nor U7549 (N_7549,N_7483,N_7275);
and U7550 (N_7550,N_7413,N_7321);
or U7551 (N_7551,N_7333,N_7313);
nand U7552 (N_7552,N_7344,N_7414);
xnor U7553 (N_7553,N_7399,N_7452);
nand U7554 (N_7554,N_7409,N_7285);
nand U7555 (N_7555,N_7308,N_7253);
or U7556 (N_7556,N_7465,N_7395);
or U7557 (N_7557,N_7426,N_7456);
nand U7558 (N_7558,N_7341,N_7350);
nand U7559 (N_7559,N_7376,N_7469);
and U7560 (N_7560,N_7397,N_7455);
or U7561 (N_7561,N_7263,N_7312);
xnor U7562 (N_7562,N_7368,N_7372);
nor U7563 (N_7563,N_7405,N_7314);
nor U7564 (N_7564,N_7381,N_7435);
and U7565 (N_7565,N_7338,N_7403);
or U7566 (N_7566,N_7430,N_7444);
and U7567 (N_7567,N_7363,N_7267);
or U7568 (N_7568,N_7457,N_7306);
or U7569 (N_7569,N_7336,N_7434);
and U7570 (N_7570,N_7294,N_7273);
nand U7571 (N_7571,N_7365,N_7295);
nand U7572 (N_7572,N_7269,N_7377);
nand U7573 (N_7573,N_7256,N_7328);
nand U7574 (N_7574,N_7374,N_7421);
nand U7575 (N_7575,N_7305,N_7270);
xnor U7576 (N_7576,N_7458,N_7346);
xnor U7577 (N_7577,N_7443,N_7283);
nor U7578 (N_7578,N_7268,N_7490);
nor U7579 (N_7579,N_7484,N_7274);
or U7580 (N_7580,N_7348,N_7278);
nor U7581 (N_7581,N_7468,N_7378);
nor U7582 (N_7582,N_7475,N_7370);
nand U7583 (N_7583,N_7432,N_7287);
xor U7584 (N_7584,N_7431,N_7390);
or U7585 (N_7585,N_7366,N_7309);
xnor U7586 (N_7586,N_7494,N_7410);
nor U7587 (N_7587,N_7355,N_7266);
or U7588 (N_7588,N_7438,N_7331);
xor U7589 (N_7589,N_7281,N_7300);
or U7590 (N_7590,N_7417,N_7252);
nand U7591 (N_7591,N_7471,N_7416);
nand U7592 (N_7592,N_7330,N_7440);
nor U7593 (N_7593,N_7259,N_7375);
xor U7594 (N_7594,N_7311,N_7383);
xnor U7595 (N_7595,N_7480,N_7441);
nand U7596 (N_7596,N_7347,N_7450);
nand U7597 (N_7597,N_7419,N_7290);
nand U7598 (N_7598,N_7496,N_7349);
nor U7599 (N_7599,N_7343,N_7439);
or U7600 (N_7600,N_7389,N_7478);
xnor U7601 (N_7601,N_7380,N_7310);
nand U7602 (N_7602,N_7327,N_7379);
and U7603 (N_7603,N_7404,N_7476);
and U7604 (N_7604,N_7481,N_7358);
nor U7605 (N_7605,N_7299,N_7364);
xnor U7606 (N_7606,N_7467,N_7303);
nor U7607 (N_7607,N_7356,N_7302);
and U7608 (N_7608,N_7477,N_7352);
xnor U7609 (N_7609,N_7296,N_7418);
nand U7610 (N_7610,N_7257,N_7487);
and U7611 (N_7611,N_7429,N_7288);
or U7612 (N_7612,N_7427,N_7340);
nor U7613 (N_7613,N_7449,N_7479);
and U7614 (N_7614,N_7460,N_7320);
xor U7615 (N_7615,N_7291,N_7459);
nand U7616 (N_7616,N_7359,N_7473);
xnor U7617 (N_7617,N_7280,N_7401);
and U7618 (N_7618,N_7470,N_7499);
xnor U7619 (N_7619,N_7386,N_7369);
and U7620 (N_7620,N_7271,N_7436);
and U7621 (N_7621,N_7322,N_7286);
and U7622 (N_7622,N_7423,N_7448);
or U7623 (N_7623,N_7250,N_7279);
and U7624 (N_7624,N_7261,N_7277);
nor U7625 (N_7625,N_7356,N_7374);
nor U7626 (N_7626,N_7378,N_7492);
nor U7627 (N_7627,N_7458,N_7298);
xor U7628 (N_7628,N_7484,N_7273);
xor U7629 (N_7629,N_7374,N_7393);
nand U7630 (N_7630,N_7374,N_7414);
nand U7631 (N_7631,N_7356,N_7410);
nor U7632 (N_7632,N_7381,N_7344);
xor U7633 (N_7633,N_7332,N_7459);
or U7634 (N_7634,N_7421,N_7336);
and U7635 (N_7635,N_7262,N_7452);
nand U7636 (N_7636,N_7273,N_7267);
nor U7637 (N_7637,N_7396,N_7403);
nand U7638 (N_7638,N_7404,N_7411);
and U7639 (N_7639,N_7470,N_7299);
or U7640 (N_7640,N_7412,N_7318);
xnor U7641 (N_7641,N_7337,N_7311);
nand U7642 (N_7642,N_7398,N_7395);
or U7643 (N_7643,N_7344,N_7280);
xnor U7644 (N_7644,N_7440,N_7392);
xnor U7645 (N_7645,N_7256,N_7442);
nand U7646 (N_7646,N_7305,N_7486);
nand U7647 (N_7647,N_7442,N_7494);
xor U7648 (N_7648,N_7381,N_7294);
xor U7649 (N_7649,N_7407,N_7305);
or U7650 (N_7650,N_7360,N_7455);
and U7651 (N_7651,N_7373,N_7370);
and U7652 (N_7652,N_7374,N_7295);
and U7653 (N_7653,N_7328,N_7265);
nand U7654 (N_7654,N_7481,N_7395);
or U7655 (N_7655,N_7404,N_7299);
or U7656 (N_7656,N_7250,N_7277);
or U7657 (N_7657,N_7366,N_7477);
nand U7658 (N_7658,N_7418,N_7460);
nand U7659 (N_7659,N_7259,N_7459);
nand U7660 (N_7660,N_7463,N_7291);
and U7661 (N_7661,N_7421,N_7450);
nor U7662 (N_7662,N_7269,N_7354);
or U7663 (N_7663,N_7408,N_7286);
nor U7664 (N_7664,N_7325,N_7435);
and U7665 (N_7665,N_7356,N_7347);
or U7666 (N_7666,N_7266,N_7363);
nor U7667 (N_7667,N_7278,N_7392);
nor U7668 (N_7668,N_7301,N_7302);
xor U7669 (N_7669,N_7473,N_7403);
nor U7670 (N_7670,N_7307,N_7377);
nor U7671 (N_7671,N_7282,N_7307);
or U7672 (N_7672,N_7291,N_7470);
nand U7673 (N_7673,N_7455,N_7429);
nor U7674 (N_7674,N_7277,N_7447);
nor U7675 (N_7675,N_7296,N_7442);
xor U7676 (N_7676,N_7438,N_7491);
nand U7677 (N_7677,N_7485,N_7355);
nor U7678 (N_7678,N_7367,N_7474);
nand U7679 (N_7679,N_7450,N_7482);
nand U7680 (N_7680,N_7345,N_7366);
xnor U7681 (N_7681,N_7323,N_7301);
nand U7682 (N_7682,N_7358,N_7277);
nand U7683 (N_7683,N_7308,N_7459);
or U7684 (N_7684,N_7389,N_7497);
xnor U7685 (N_7685,N_7336,N_7341);
or U7686 (N_7686,N_7406,N_7387);
nor U7687 (N_7687,N_7431,N_7256);
xor U7688 (N_7688,N_7277,N_7488);
nand U7689 (N_7689,N_7277,N_7367);
xor U7690 (N_7690,N_7339,N_7312);
nand U7691 (N_7691,N_7255,N_7369);
nand U7692 (N_7692,N_7365,N_7274);
or U7693 (N_7693,N_7271,N_7380);
nor U7694 (N_7694,N_7291,N_7444);
and U7695 (N_7695,N_7399,N_7383);
or U7696 (N_7696,N_7256,N_7466);
xor U7697 (N_7697,N_7487,N_7335);
nor U7698 (N_7698,N_7470,N_7417);
xnor U7699 (N_7699,N_7381,N_7434);
and U7700 (N_7700,N_7256,N_7432);
xor U7701 (N_7701,N_7478,N_7343);
or U7702 (N_7702,N_7476,N_7295);
nor U7703 (N_7703,N_7399,N_7346);
nor U7704 (N_7704,N_7480,N_7414);
and U7705 (N_7705,N_7276,N_7449);
nand U7706 (N_7706,N_7461,N_7342);
or U7707 (N_7707,N_7481,N_7406);
nor U7708 (N_7708,N_7370,N_7372);
or U7709 (N_7709,N_7487,N_7332);
nand U7710 (N_7710,N_7304,N_7310);
or U7711 (N_7711,N_7457,N_7454);
or U7712 (N_7712,N_7283,N_7282);
xor U7713 (N_7713,N_7418,N_7284);
and U7714 (N_7714,N_7343,N_7470);
and U7715 (N_7715,N_7371,N_7334);
and U7716 (N_7716,N_7316,N_7499);
and U7717 (N_7717,N_7386,N_7301);
xor U7718 (N_7718,N_7260,N_7265);
xor U7719 (N_7719,N_7307,N_7413);
and U7720 (N_7720,N_7465,N_7394);
xnor U7721 (N_7721,N_7322,N_7476);
or U7722 (N_7722,N_7436,N_7371);
nand U7723 (N_7723,N_7322,N_7331);
and U7724 (N_7724,N_7265,N_7419);
nand U7725 (N_7725,N_7401,N_7260);
or U7726 (N_7726,N_7469,N_7320);
and U7727 (N_7727,N_7296,N_7338);
xnor U7728 (N_7728,N_7393,N_7474);
and U7729 (N_7729,N_7429,N_7341);
xor U7730 (N_7730,N_7450,N_7320);
nor U7731 (N_7731,N_7302,N_7394);
and U7732 (N_7732,N_7354,N_7410);
nor U7733 (N_7733,N_7270,N_7438);
nand U7734 (N_7734,N_7310,N_7260);
or U7735 (N_7735,N_7296,N_7339);
nor U7736 (N_7736,N_7426,N_7412);
nor U7737 (N_7737,N_7360,N_7475);
nor U7738 (N_7738,N_7252,N_7279);
or U7739 (N_7739,N_7312,N_7486);
xor U7740 (N_7740,N_7478,N_7277);
nor U7741 (N_7741,N_7457,N_7353);
xnor U7742 (N_7742,N_7379,N_7494);
and U7743 (N_7743,N_7416,N_7452);
xnor U7744 (N_7744,N_7396,N_7455);
or U7745 (N_7745,N_7457,N_7324);
xnor U7746 (N_7746,N_7396,N_7303);
xor U7747 (N_7747,N_7318,N_7389);
and U7748 (N_7748,N_7269,N_7291);
and U7749 (N_7749,N_7388,N_7435);
nand U7750 (N_7750,N_7616,N_7586);
nand U7751 (N_7751,N_7547,N_7684);
xor U7752 (N_7752,N_7565,N_7534);
nor U7753 (N_7753,N_7657,N_7551);
xnor U7754 (N_7754,N_7729,N_7689);
nor U7755 (N_7755,N_7738,N_7579);
xnor U7756 (N_7756,N_7699,N_7695);
nor U7757 (N_7757,N_7652,N_7604);
nand U7758 (N_7758,N_7722,N_7585);
xor U7759 (N_7759,N_7618,N_7666);
and U7760 (N_7760,N_7705,N_7563);
xor U7761 (N_7761,N_7671,N_7549);
xor U7762 (N_7762,N_7615,N_7646);
xor U7763 (N_7763,N_7538,N_7676);
nand U7764 (N_7764,N_7726,N_7522);
or U7765 (N_7765,N_7568,N_7701);
xor U7766 (N_7766,N_7527,N_7629);
and U7767 (N_7767,N_7728,N_7611);
or U7768 (N_7768,N_7574,N_7672);
or U7769 (N_7769,N_7623,N_7501);
nand U7770 (N_7770,N_7668,N_7747);
nand U7771 (N_7771,N_7737,N_7720);
or U7772 (N_7772,N_7533,N_7572);
and U7773 (N_7773,N_7554,N_7731);
nand U7774 (N_7774,N_7584,N_7557);
nor U7775 (N_7775,N_7599,N_7704);
or U7776 (N_7776,N_7511,N_7513);
nor U7777 (N_7777,N_7583,N_7597);
xnor U7778 (N_7778,N_7600,N_7706);
and U7779 (N_7779,N_7590,N_7725);
nor U7780 (N_7780,N_7564,N_7667);
and U7781 (N_7781,N_7658,N_7578);
or U7782 (N_7782,N_7598,N_7561);
and U7783 (N_7783,N_7525,N_7632);
nor U7784 (N_7784,N_7727,N_7503);
nand U7785 (N_7785,N_7541,N_7638);
xor U7786 (N_7786,N_7696,N_7636);
nand U7787 (N_7787,N_7575,N_7540);
nor U7788 (N_7788,N_7520,N_7748);
nor U7789 (N_7789,N_7645,N_7682);
nor U7790 (N_7790,N_7723,N_7506);
and U7791 (N_7791,N_7630,N_7651);
nand U7792 (N_7792,N_7544,N_7692);
xnor U7793 (N_7793,N_7673,N_7596);
or U7794 (N_7794,N_7663,N_7530);
nand U7795 (N_7795,N_7620,N_7580);
or U7796 (N_7796,N_7734,N_7573);
xor U7797 (N_7797,N_7550,N_7553);
and U7798 (N_7798,N_7504,N_7685);
or U7799 (N_7799,N_7532,N_7507);
xnor U7800 (N_7800,N_7649,N_7546);
or U7801 (N_7801,N_7736,N_7608);
or U7802 (N_7802,N_7505,N_7593);
xor U7803 (N_7803,N_7612,N_7650);
nand U7804 (N_7804,N_7512,N_7606);
xnor U7805 (N_7805,N_7543,N_7703);
nor U7806 (N_7806,N_7721,N_7717);
nand U7807 (N_7807,N_7719,N_7669);
nand U7808 (N_7808,N_7502,N_7690);
xor U7809 (N_7809,N_7654,N_7661);
xor U7810 (N_7810,N_7714,N_7688);
nor U7811 (N_7811,N_7677,N_7621);
nor U7812 (N_7812,N_7740,N_7655);
nand U7813 (N_7813,N_7745,N_7660);
nand U7814 (N_7814,N_7603,N_7508);
or U7815 (N_7815,N_7560,N_7633);
nor U7816 (N_7816,N_7555,N_7637);
nor U7817 (N_7817,N_7576,N_7531);
xnor U7818 (N_7818,N_7614,N_7698);
xor U7819 (N_7819,N_7521,N_7622);
nand U7820 (N_7820,N_7592,N_7577);
or U7821 (N_7821,N_7524,N_7713);
and U7822 (N_7822,N_7697,N_7617);
nand U7823 (N_7823,N_7562,N_7643);
nand U7824 (N_7824,N_7686,N_7647);
and U7825 (N_7825,N_7744,N_7640);
nand U7826 (N_7826,N_7581,N_7523);
and U7827 (N_7827,N_7595,N_7567);
nand U7828 (N_7828,N_7642,N_7710);
nor U7829 (N_7829,N_7702,N_7733);
or U7830 (N_7830,N_7517,N_7709);
or U7831 (N_7831,N_7635,N_7625);
nand U7832 (N_7832,N_7634,N_7715);
and U7833 (N_7833,N_7749,N_7607);
nor U7834 (N_7834,N_7558,N_7602);
nor U7835 (N_7835,N_7735,N_7631);
and U7836 (N_7836,N_7571,N_7648);
nand U7837 (N_7837,N_7601,N_7624);
or U7838 (N_7838,N_7746,N_7548);
xor U7839 (N_7839,N_7675,N_7742);
and U7840 (N_7840,N_7569,N_7589);
nor U7841 (N_7841,N_7691,N_7588);
nand U7842 (N_7842,N_7528,N_7542);
xor U7843 (N_7843,N_7619,N_7693);
xor U7844 (N_7844,N_7518,N_7656);
or U7845 (N_7845,N_7680,N_7627);
nor U7846 (N_7846,N_7539,N_7514);
nand U7847 (N_7847,N_7659,N_7628);
nand U7848 (N_7848,N_7670,N_7732);
xnor U7849 (N_7849,N_7674,N_7519);
nor U7850 (N_7850,N_7711,N_7529);
nor U7851 (N_7851,N_7545,N_7626);
nor U7852 (N_7852,N_7741,N_7730);
and U7853 (N_7853,N_7700,N_7536);
xnor U7854 (N_7854,N_7641,N_7587);
nor U7855 (N_7855,N_7678,N_7694);
or U7856 (N_7856,N_7556,N_7724);
xor U7857 (N_7857,N_7515,N_7639);
nor U7858 (N_7858,N_7582,N_7594);
nor U7859 (N_7859,N_7537,N_7681);
xnor U7860 (N_7860,N_7662,N_7552);
nor U7861 (N_7861,N_7665,N_7687);
nor U7862 (N_7862,N_7510,N_7535);
xor U7863 (N_7863,N_7610,N_7609);
nor U7864 (N_7864,N_7739,N_7679);
and U7865 (N_7865,N_7526,N_7605);
xor U7866 (N_7866,N_7570,N_7644);
xor U7867 (N_7867,N_7500,N_7591);
nor U7868 (N_7868,N_7708,N_7743);
nor U7869 (N_7869,N_7712,N_7716);
nand U7870 (N_7870,N_7683,N_7653);
or U7871 (N_7871,N_7664,N_7707);
nor U7872 (N_7872,N_7509,N_7613);
nand U7873 (N_7873,N_7516,N_7559);
nand U7874 (N_7874,N_7718,N_7566);
or U7875 (N_7875,N_7707,N_7683);
xor U7876 (N_7876,N_7585,N_7601);
nor U7877 (N_7877,N_7530,N_7692);
and U7878 (N_7878,N_7741,N_7743);
or U7879 (N_7879,N_7713,N_7640);
and U7880 (N_7880,N_7652,N_7679);
and U7881 (N_7881,N_7601,N_7503);
nor U7882 (N_7882,N_7557,N_7668);
or U7883 (N_7883,N_7703,N_7562);
and U7884 (N_7884,N_7507,N_7662);
and U7885 (N_7885,N_7699,N_7732);
xnor U7886 (N_7886,N_7746,N_7738);
nand U7887 (N_7887,N_7719,N_7550);
and U7888 (N_7888,N_7507,N_7667);
or U7889 (N_7889,N_7707,N_7637);
and U7890 (N_7890,N_7514,N_7608);
or U7891 (N_7891,N_7680,N_7612);
nand U7892 (N_7892,N_7744,N_7593);
nor U7893 (N_7893,N_7730,N_7586);
and U7894 (N_7894,N_7608,N_7634);
nor U7895 (N_7895,N_7597,N_7585);
or U7896 (N_7896,N_7643,N_7576);
and U7897 (N_7897,N_7635,N_7567);
nor U7898 (N_7898,N_7678,N_7543);
and U7899 (N_7899,N_7687,N_7592);
xor U7900 (N_7900,N_7721,N_7519);
nor U7901 (N_7901,N_7513,N_7583);
and U7902 (N_7902,N_7649,N_7567);
nand U7903 (N_7903,N_7689,N_7603);
xnor U7904 (N_7904,N_7527,N_7560);
nand U7905 (N_7905,N_7529,N_7630);
nor U7906 (N_7906,N_7664,N_7583);
nor U7907 (N_7907,N_7720,N_7525);
or U7908 (N_7908,N_7500,N_7581);
nor U7909 (N_7909,N_7586,N_7717);
xor U7910 (N_7910,N_7720,N_7557);
xnor U7911 (N_7911,N_7737,N_7597);
or U7912 (N_7912,N_7603,N_7563);
nand U7913 (N_7913,N_7535,N_7749);
nand U7914 (N_7914,N_7677,N_7716);
nand U7915 (N_7915,N_7504,N_7648);
and U7916 (N_7916,N_7665,N_7586);
nor U7917 (N_7917,N_7558,N_7617);
nor U7918 (N_7918,N_7506,N_7578);
xnor U7919 (N_7919,N_7643,N_7711);
xnor U7920 (N_7920,N_7693,N_7715);
xor U7921 (N_7921,N_7612,N_7663);
nand U7922 (N_7922,N_7592,N_7713);
nand U7923 (N_7923,N_7585,N_7525);
or U7924 (N_7924,N_7542,N_7626);
nor U7925 (N_7925,N_7516,N_7590);
xnor U7926 (N_7926,N_7607,N_7640);
nor U7927 (N_7927,N_7713,N_7616);
xnor U7928 (N_7928,N_7724,N_7625);
xnor U7929 (N_7929,N_7738,N_7653);
nand U7930 (N_7930,N_7718,N_7634);
xnor U7931 (N_7931,N_7610,N_7737);
or U7932 (N_7932,N_7663,N_7656);
nand U7933 (N_7933,N_7735,N_7668);
nor U7934 (N_7934,N_7615,N_7735);
and U7935 (N_7935,N_7719,N_7566);
or U7936 (N_7936,N_7677,N_7614);
and U7937 (N_7937,N_7633,N_7746);
and U7938 (N_7938,N_7547,N_7559);
or U7939 (N_7939,N_7696,N_7571);
nand U7940 (N_7940,N_7652,N_7749);
nand U7941 (N_7941,N_7541,N_7736);
xnor U7942 (N_7942,N_7552,N_7648);
xor U7943 (N_7943,N_7531,N_7537);
and U7944 (N_7944,N_7574,N_7738);
and U7945 (N_7945,N_7705,N_7583);
xnor U7946 (N_7946,N_7517,N_7668);
xnor U7947 (N_7947,N_7532,N_7527);
or U7948 (N_7948,N_7599,N_7634);
xor U7949 (N_7949,N_7661,N_7611);
nor U7950 (N_7950,N_7600,N_7619);
nor U7951 (N_7951,N_7694,N_7601);
or U7952 (N_7952,N_7554,N_7585);
or U7953 (N_7953,N_7721,N_7660);
and U7954 (N_7954,N_7559,N_7745);
xnor U7955 (N_7955,N_7564,N_7682);
and U7956 (N_7956,N_7748,N_7691);
nor U7957 (N_7957,N_7643,N_7716);
nor U7958 (N_7958,N_7647,N_7669);
xnor U7959 (N_7959,N_7687,N_7626);
nand U7960 (N_7960,N_7631,N_7617);
nand U7961 (N_7961,N_7739,N_7655);
nand U7962 (N_7962,N_7742,N_7623);
or U7963 (N_7963,N_7690,N_7585);
or U7964 (N_7964,N_7742,N_7643);
nand U7965 (N_7965,N_7518,N_7563);
nor U7966 (N_7966,N_7652,N_7603);
xor U7967 (N_7967,N_7510,N_7550);
or U7968 (N_7968,N_7551,N_7647);
nor U7969 (N_7969,N_7550,N_7536);
or U7970 (N_7970,N_7680,N_7710);
and U7971 (N_7971,N_7520,N_7662);
nand U7972 (N_7972,N_7542,N_7527);
or U7973 (N_7973,N_7629,N_7687);
nor U7974 (N_7974,N_7693,N_7588);
nor U7975 (N_7975,N_7736,N_7741);
nand U7976 (N_7976,N_7645,N_7547);
and U7977 (N_7977,N_7565,N_7743);
or U7978 (N_7978,N_7567,N_7568);
and U7979 (N_7979,N_7658,N_7749);
xor U7980 (N_7980,N_7670,N_7748);
nor U7981 (N_7981,N_7663,N_7592);
nor U7982 (N_7982,N_7727,N_7698);
xnor U7983 (N_7983,N_7627,N_7614);
nor U7984 (N_7984,N_7599,N_7587);
or U7985 (N_7985,N_7621,N_7600);
and U7986 (N_7986,N_7679,N_7671);
nor U7987 (N_7987,N_7622,N_7564);
nor U7988 (N_7988,N_7712,N_7532);
xnor U7989 (N_7989,N_7741,N_7523);
xnor U7990 (N_7990,N_7736,N_7513);
nand U7991 (N_7991,N_7549,N_7529);
xor U7992 (N_7992,N_7721,N_7696);
xor U7993 (N_7993,N_7650,N_7667);
nor U7994 (N_7994,N_7605,N_7658);
nor U7995 (N_7995,N_7552,N_7588);
xnor U7996 (N_7996,N_7741,N_7675);
nand U7997 (N_7997,N_7606,N_7683);
nor U7998 (N_7998,N_7530,N_7682);
xnor U7999 (N_7999,N_7739,N_7694);
xor U8000 (N_8000,N_7812,N_7928);
nor U8001 (N_8001,N_7792,N_7949);
and U8002 (N_8002,N_7852,N_7964);
nor U8003 (N_8003,N_7809,N_7799);
and U8004 (N_8004,N_7796,N_7752);
and U8005 (N_8005,N_7993,N_7791);
nand U8006 (N_8006,N_7991,N_7974);
xor U8007 (N_8007,N_7768,N_7894);
xor U8008 (N_8008,N_7818,N_7882);
nand U8009 (N_8009,N_7827,N_7814);
and U8010 (N_8010,N_7793,N_7878);
nand U8011 (N_8011,N_7824,N_7838);
xnor U8012 (N_8012,N_7750,N_7988);
xnor U8013 (N_8013,N_7948,N_7965);
and U8014 (N_8014,N_7914,N_7817);
nor U8015 (N_8015,N_7918,N_7955);
and U8016 (N_8016,N_7820,N_7961);
nor U8017 (N_8017,N_7939,N_7953);
and U8018 (N_8018,N_7856,N_7813);
or U8019 (N_8019,N_7760,N_7777);
nor U8020 (N_8020,N_7780,N_7978);
xnor U8021 (N_8021,N_7866,N_7862);
or U8022 (N_8022,N_7915,N_7951);
nand U8023 (N_8023,N_7850,N_7963);
and U8024 (N_8024,N_7819,N_7830);
xor U8025 (N_8025,N_7920,N_7895);
nand U8026 (N_8026,N_7945,N_7873);
xnor U8027 (N_8027,N_7903,N_7874);
nor U8028 (N_8028,N_7858,N_7968);
nand U8029 (N_8029,N_7816,N_7922);
or U8030 (N_8030,N_7908,N_7766);
nor U8031 (N_8031,N_7784,N_7962);
or U8032 (N_8032,N_7800,N_7783);
xnor U8033 (N_8033,N_7969,N_7941);
nand U8034 (N_8034,N_7900,N_7888);
nand U8035 (N_8035,N_7801,N_7810);
xnor U8036 (N_8036,N_7901,N_7979);
xnor U8037 (N_8037,N_7757,N_7940);
xnor U8038 (N_8038,N_7835,N_7937);
nand U8039 (N_8039,N_7861,N_7872);
nor U8040 (N_8040,N_7851,N_7758);
nor U8041 (N_8041,N_7855,N_7846);
or U8042 (N_8042,N_7942,N_7854);
or U8043 (N_8043,N_7831,N_7971);
nor U8044 (N_8044,N_7843,N_7825);
and U8045 (N_8045,N_7849,N_7913);
or U8046 (N_8046,N_7970,N_7980);
or U8047 (N_8047,N_7870,N_7805);
nor U8048 (N_8048,N_7997,N_7876);
nor U8049 (N_8049,N_7877,N_7959);
or U8050 (N_8050,N_7926,N_7823);
or U8051 (N_8051,N_7885,N_7925);
nand U8052 (N_8052,N_7803,N_7919);
or U8053 (N_8053,N_7836,N_7763);
nand U8054 (N_8054,N_7938,N_7931);
or U8055 (N_8055,N_7998,N_7898);
or U8056 (N_8056,N_7880,N_7806);
xor U8057 (N_8057,N_7815,N_7773);
or U8058 (N_8058,N_7857,N_7952);
xor U8059 (N_8059,N_7935,N_7807);
nand U8060 (N_8060,N_7776,N_7767);
nand U8061 (N_8061,N_7759,N_7821);
or U8062 (N_8062,N_7797,N_7987);
nand U8063 (N_8063,N_7977,N_7842);
and U8064 (N_8064,N_7957,N_7751);
or U8065 (N_8065,N_7875,N_7999);
nand U8066 (N_8066,N_7984,N_7907);
and U8067 (N_8067,N_7902,N_7867);
xor U8068 (N_8068,N_7921,N_7986);
nor U8069 (N_8069,N_7924,N_7932);
and U8070 (N_8070,N_7782,N_7972);
xnor U8071 (N_8071,N_7860,N_7912);
nor U8072 (N_8072,N_7943,N_7887);
and U8073 (N_8073,N_7983,N_7802);
and U8074 (N_8074,N_7789,N_7833);
nand U8075 (N_8075,N_7884,N_7906);
and U8076 (N_8076,N_7911,N_7905);
or U8077 (N_8077,N_7765,N_7996);
or U8078 (N_8078,N_7770,N_7864);
nand U8079 (N_8079,N_7859,N_7779);
nand U8080 (N_8080,N_7985,N_7891);
nand U8081 (N_8081,N_7853,N_7992);
or U8082 (N_8082,N_7989,N_7771);
xnor U8083 (N_8083,N_7787,N_7990);
xor U8084 (N_8084,N_7995,N_7944);
and U8085 (N_8085,N_7927,N_7865);
xnor U8086 (N_8086,N_7845,N_7909);
xnor U8087 (N_8087,N_7910,N_7761);
or U8088 (N_8088,N_7960,N_7934);
or U8089 (N_8089,N_7804,N_7848);
xnor U8090 (N_8090,N_7764,N_7762);
nor U8091 (N_8091,N_7847,N_7772);
and U8092 (N_8092,N_7795,N_7774);
or U8093 (N_8093,N_7841,N_7946);
nand U8094 (N_8094,N_7755,N_7798);
and U8095 (N_8095,N_7958,N_7889);
and U8096 (N_8096,N_7899,N_7897);
nor U8097 (N_8097,N_7973,N_7863);
nor U8098 (N_8098,N_7936,N_7954);
xnor U8099 (N_8099,N_7868,N_7886);
nor U8100 (N_8100,N_7923,N_7832);
and U8101 (N_8101,N_7904,N_7756);
nand U8102 (N_8102,N_7826,N_7930);
and U8103 (N_8103,N_7929,N_7917);
or U8104 (N_8104,N_7896,N_7822);
xnor U8105 (N_8105,N_7839,N_7775);
nand U8106 (N_8106,N_7786,N_7881);
and U8107 (N_8107,N_7933,N_7976);
or U8108 (N_8108,N_7981,N_7892);
xnor U8109 (N_8109,N_7778,N_7966);
and U8110 (N_8110,N_7883,N_7811);
nand U8111 (N_8111,N_7834,N_7956);
and U8112 (N_8112,N_7879,N_7871);
xor U8113 (N_8113,N_7844,N_7781);
and U8114 (N_8114,N_7788,N_7994);
and U8115 (N_8115,N_7829,N_7840);
or U8116 (N_8116,N_7828,N_7975);
or U8117 (N_8117,N_7753,N_7794);
xnor U8118 (N_8118,N_7808,N_7837);
nor U8119 (N_8119,N_7790,N_7890);
and U8120 (N_8120,N_7754,N_7869);
nor U8121 (N_8121,N_7769,N_7982);
or U8122 (N_8122,N_7950,N_7893);
xor U8123 (N_8123,N_7785,N_7916);
or U8124 (N_8124,N_7967,N_7947);
and U8125 (N_8125,N_7827,N_7850);
nor U8126 (N_8126,N_7839,N_7927);
and U8127 (N_8127,N_7880,N_7907);
nand U8128 (N_8128,N_7778,N_7960);
xnor U8129 (N_8129,N_7833,N_7858);
nand U8130 (N_8130,N_7750,N_7904);
nand U8131 (N_8131,N_7933,N_7949);
xnor U8132 (N_8132,N_7956,N_7846);
or U8133 (N_8133,N_7890,N_7923);
xor U8134 (N_8134,N_7945,N_7821);
or U8135 (N_8135,N_7876,N_7996);
or U8136 (N_8136,N_7758,N_7882);
nor U8137 (N_8137,N_7847,N_7921);
nand U8138 (N_8138,N_7873,N_7763);
nand U8139 (N_8139,N_7839,N_7824);
nand U8140 (N_8140,N_7913,N_7817);
and U8141 (N_8141,N_7767,N_7899);
nand U8142 (N_8142,N_7855,N_7819);
xor U8143 (N_8143,N_7988,N_7763);
nor U8144 (N_8144,N_7801,N_7807);
or U8145 (N_8145,N_7929,N_7908);
and U8146 (N_8146,N_7968,N_7764);
or U8147 (N_8147,N_7788,N_7798);
and U8148 (N_8148,N_7905,N_7865);
xor U8149 (N_8149,N_7902,N_7855);
or U8150 (N_8150,N_7897,N_7962);
and U8151 (N_8151,N_7974,N_7956);
xnor U8152 (N_8152,N_7785,N_7924);
xnor U8153 (N_8153,N_7781,N_7823);
nand U8154 (N_8154,N_7756,N_7971);
and U8155 (N_8155,N_7817,N_7932);
or U8156 (N_8156,N_7918,N_7900);
nor U8157 (N_8157,N_7973,N_7795);
nor U8158 (N_8158,N_7898,N_7965);
xor U8159 (N_8159,N_7930,N_7903);
xor U8160 (N_8160,N_7986,N_7786);
xor U8161 (N_8161,N_7773,N_7825);
xor U8162 (N_8162,N_7968,N_7859);
nor U8163 (N_8163,N_7953,N_7792);
nand U8164 (N_8164,N_7751,N_7939);
xor U8165 (N_8165,N_7897,N_7974);
and U8166 (N_8166,N_7905,N_7868);
nand U8167 (N_8167,N_7774,N_7870);
or U8168 (N_8168,N_7924,N_7887);
xnor U8169 (N_8169,N_7815,N_7974);
xnor U8170 (N_8170,N_7758,N_7911);
or U8171 (N_8171,N_7895,N_7965);
xnor U8172 (N_8172,N_7805,N_7925);
nand U8173 (N_8173,N_7778,N_7883);
xor U8174 (N_8174,N_7892,N_7780);
nor U8175 (N_8175,N_7952,N_7802);
and U8176 (N_8176,N_7915,N_7882);
xnor U8177 (N_8177,N_7824,N_7981);
xor U8178 (N_8178,N_7874,N_7799);
and U8179 (N_8179,N_7801,N_7750);
and U8180 (N_8180,N_7877,N_7801);
and U8181 (N_8181,N_7988,N_7946);
or U8182 (N_8182,N_7972,N_7884);
and U8183 (N_8183,N_7872,N_7755);
and U8184 (N_8184,N_7760,N_7801);
and U8185 (N_8185,N_7851,N_7791);
and U8186 (N_8186,N_7894,N_7952);
and U8187 (N_8187,N_7960,N_7848);
and U8188 (N_8188,N_7815,N_7794);
and U8189 (N_8189,N_7755,N_7910);
nand U8190 (N_8190,N_7817,N_7776);
nor U8191 (N_8191,N_7924,N_7863);
nor U8192 (N_8192,N_7838,N_7890);
nor U8193 (N_8193,N_7954,N_7971);
or U8194 (N_8194,N_7826,N_7802);
or U8195 (N_8195,N_7826,N_7754);
and U8196 (N_8196,N_7761,N_7821);
and U8197 (N_8197,N_7880,N_7995);
nand U8198 (N_8198,N_7798,N_7909);
nor U8199 (N_8199,N_7982,N_7838);
nand U8200 (N_8200,N_7890,N_7983);
nor U8201 (N_8201,N_7971,N_7821);
and U8202 (N_8202,N_7757,N_7862);
and U8203 (N_8203,N_7996,N_7818);
and U8204 (N_8204,N_7991,N_7883);
xnor U8205 (N_8205,N_7948,N_7840);
xor U8206 (N_8206,N_7831,N_7825);
or U8207 (N_8207,N_7880,N_7919);
nor U8208 (N_8208,N_7995,N_7860);
nand U8209 (N_8209,N_7759,N_7822);
nor U8210 (N_8210,N_7985,N_7978);
nand U8211 (N_8211,N_7818,N_7893);
nand U8212 (N_8212,N_7992,N_7946);
xnor U8213 (N_8213,N_7894,N_7803);
nand U8214 (N_8214,N_7979,N_7841);
nor U8215 (N_8215,N_7866,N_7915);
nand U8216 (N_8216,N_7986,N_7845);
xnor U8217 (N_8217,N_7909,N_7782);
xnor U8218 (N_8218,N_7838,N_7812);
or U8219 (N_8219,N_7985,N_7850);
or U8220 (N_8220,N_7887,N_7961);
or U8221 (N_8221,N_7851,N_7933);
xnor U8222 (N_8222,N_7913,N_7828);
or U8223 (N_8223,N_7945,N_7845);
nand U8224 (N_8224,N_7935,N_7773);
nor U8225 (N_8225,N_7851,N_7787);
and U8226 (N_8226,N_7993,N_7898);
nand U8227 (N_8227,N_7964,N_7845);
nor U8228 (N_8228,N_7803,N_7988);
and U8229 (N_8229,N_7879,N_7936);
nand U8230 (N_8230,N_7970,N_7810);
or U8231 (N_8231,N_7767,N_7853);
or U8232 (N_8232,N_7889,N_7917);
nand U8233 (N_8233,N_7818,N_7782);
and U8234 (N_8234,N_7992,N_7825);
xnor U8235 (N_8235,N_7977,N_7889);
xnor U8236 (N_8236,N_7897,N_7864);
nand U8237 (N_8237,N_7823,N_7958);
nand U8238 (N_8238,N_7977,N_7804);
nor U8239 (N_8239,N_7761,N_7942);
and U8240 (N_8240,N_7962,N_7862);
nand U8241 (N_8241,N_7942,N_7904);
xnor U8242 (N_8242,N_7785,N_7751);
xor U8243 (N_8243,N_7935,N_7842);
nor U8244 (N_8244,N_7892,N_7838);
xor U8245 (N_8245,N_7828,N_7959);
and U8246 (N_8246,N_7993,N_7918);
nand U8247 (N_8247,N_7832,N_7942);
nor U8248 (N_8248,N_7937,N_7755);
nand U8249 (N_8249,N_7875,N_7838);
nand U8250 (N_8250,N_8014,N_8045);
nand U8251 (N_8251,N_8005,N_8000);
xor U8252 (N_8252,N_8093,N_8229);
nand U8253 (N_8253,N_8115,N_8010);
nor U8254 (N_8254,N_8058,N_8172);
nand U8255 (N_8255,N_8088,N_8158);
and U8256 (N_8256,N_8166,N_8080);
nand U8257 (N_8257,N_8248,N_8157);
nor U8258 (N_8258,N_8220,N_8242);
nand U8259 (N_8259,N_8222,N_8150);
nand U8260 (N_8260,N_8208,N_8216);
xor U8261 (N_8261,N_8186,N_8090);
nor U8262 (N_8262,N_8237,N_8135);
xnor U8263 (N_8263,N_8230,N_8199);
nor U8264 (N_8264,N_8040,N_8089);
xor U8265 (N_8265,N_8130,N_8205);
nor U8266 (N_8266,N_8162,N_8092);
nor U8267 (N_8267,N_8029,N_8160);
and U8268 (N_8268,N_8132,N_8108);
and U8269 (N_8269,N_8074,N_8110);
xnor U8270 (N_8270,N_8151,N_8038);
nor U8271 (N_8271,N_8169,N_8210);
nor U8272 (N_8272,N_8137,N_8127);
nor U8273 (N_8273,N_8125,N_8138);
or U8274 (N_8274,N_8111,N_8212);
and U8275 (N_8275,N_8214,N_8145);
xnor U8276 (N_8276,N_8224,N_8048);
nor U8277 (N_8277,N_8004,N_8245);
nor U8278 (N_8278,N_8042,N_8188);
or U8279 (N_8279,N_8066,N_8197);
nand U8280 (N_8280,N_8236,N_8034);
nor U8281 (N_8281,N_8116,N_8049);
or U8282 (N_8282,N_8223,N_8241);
or U8283 (N_8283,N_8052,N_8209);
nor U8284 (N_8284,N_8118,N_8023);
xor U8285 (N_8285,N_8202,N_8095);
or U8286 (N_8286,N_8142,N_8140);
or U8287 (N_8287,N_8123,N_8022);
xor U8288 (N_8288,N_8194,N_8035);
nand U8289 (N_8289,N_8215,N_8124);
and U8290 (N_8290,N_8011,N_8185);
or U8291 (N_8291,N_8053,N_8070);
nor U8292 (N_8292,N_8152,N_8064);
nor U8293 (N_8293,N_8012,N_8161);
nand U8294 (N_8294,N_8069,N_8156);
nand U8295 (N_8295,N_8238,N_8027);
nand U8296 (N_8296,N_8146,N_8143);
and U8297 (N_8297,N_8239,N_8244);
nand U8298 (N_8298,N_8184,N_8031);
nor U8299 (N_8299,N_8227,N_8232);
or U8300 (N_8300,N_8191,N_8200);
xnor U8301 (N_8301,N_8065,N_8013);
nor U8302 (N_8302,N_8176,N_8018);
xnor U8303 (N_8303,N_8047,N_8008);
nor U8304 (N_8304,N_8153,N_8078);
nor U8305 (N_8305,N_8059,N_8067);
nand U8306 (N_8306,N_8207,N_8213);
nand U8307 (N_8307,N_8094,N_8086);
xor U8308 (N_8308,N_8003,N_8032);
or U8309 (N_8309,N_8249,N_8006);
or U8310 (N_8310,N_8233,N_8195);
or U8311 (N_8311,N_8148,N_8063);
nor U8312 (N_8312,N_8226,N_8015);
or U8313 (N_8313,N_8025,N_8033);
nand U8314 (N_8314,N_8037,N_8192);
nand U8315 (N_8315,N_8060,N_8225);
and U8316 (N_8316,N_8073,N_8007);
nor U8317 (N_8317,N_8136,N_8087);
and U8318 (N_8318,N_8198,N_8133);
nor U8319 (N_8319,N_8109,N_8147);
nor U8320 (N_8320,N_8046,N_8247);
and U8321 (N_8321,N_8163,N_8174);
xnor U8322 (N_8322,N_8039,N_8019);
nand U8323 (N_8323,N_8113,N_8056);
nand U8324 (N_8324,N_8167,N_8119);
or U8325 (N_8325,N_8082,N_8055);
nor U8326 (N_8326,N_8203,N_8218);
nand U8327 (N_8327,N_8068,N_8170);
xnor U8328 (N_8328,N_8141,N_8001);
nor U8329 (N_8329,N_8009,N_8181);
nor U8330 (N_8330,N_8175,N_8081);
nand U8331 (N_8331,N_8179,N_8149);
xnor U8332 (N_8332,N_8168,N_8120);
nor U8333 (N_8333,N_8024,N_8107);
or U8334 (N_8334,N_8196,N_8129);
and U8335 (N_8335,N_8234,N_8126);
xor U8336 (N_8336,N_8204,N_8096);
nor U8337 (N_8337,N_8097,N_8085);
nand U8338 (N_8338,N_8190,N_8084);
or U8339 (N_8339,N_8102,N_8100);
or U8340 (N_8340,N_8075,N_8182);
xnor U8341 (N_8341,N_8122,N_8144);
nand U8342 (N_8342,N_8187,N_8180);
and U8343 (N_8343,N_8246,N_8072);
and U8344 (N_8344,N_8164,N_8021);
or U8345 (N_8345,N_8206,N_8057);
and U8346 (N_8346,N_8231,N_8183);
xor U8347 (N_8347,N_8114,N_8101);
and U8348 (N_8348,N_8201,N_8211);
xor U8349 (N_8349,N_8016,N_8134);
and U8350 (N_8350,N_8098,N_8221);
xor U8351 (N_8351,N_8178,N_8228);
and U8352 (N_8352,N_8030,N_8155);
nor U8353 (N_8353,N_8139,N_8112);
nor U8354 (N_8354,N_8050,N_8104);
and U8355 (N_8355,N_8217,N_8002);
xor U8356 (N_8356,N_8054,N_8121);
or U8357 (N_8357,N_8131,N_8154);
nor U8358 (N_8358,N_8117,N_8159);
xnor U8359 (N_8359,N_8235,N_8189);
and U8360 (N_8360,N_8083,N_8079);
nand U8361 (N_8361,N_8243,N_8106);
and U8362 (N_8362,N_8043,N_8193);
nand U8363 (N_8363,N_8041,N_8128);
nand U8364 (N_8364,N_8219,N_8036);
xor U8365 (N_8365,N_8028,N_8076);
and U8366 (N_8366,N_8240,N_8099);
nor U8367 (N_8367,N_8165,N_8077);
and U8368 (N_8368,N_8017,N_8062);
or U8369 (N_8369,N_8091,N_8171);
xnor U8370 (N_8370,N_8105,N_8177);
nand U8371 (N_8371,N_8051,N_8173);
or U8372 (N_8372,N_8071,N_8061);
nand U8373 (N_8373,N_8044,N_8026);
nand U8374 (N_8374,N_8020,N_8103);
nand U8375 (N_8375,N_8161,N_8213);
xnor U8376 (N_8376,N_8216,N_8168);
or U8377 (N_8377,N_8247,N_8068);
nor U8378 (N_8378,N_8206,N_8141);
and U8379 (N_8379,N_8083,N_8122);
and U8380 (N_8380,N_8077,N_8143);
nand U8381 (N_8381,N_8005,N_8053);
xor U8382 (N_8382,N_8235,N_8079);
and U8383 (N_8383,N_8230,N_8048);
xor U8384 (N_8384,N_8234,N_8138);
nand U8385 (N_8385,N_8046,N_8174);
xnor U8386 (N_8386,N_8099,N_8160);
nor U8387 (N_8387,N_8184,N_8110);
nor U8388 (N_8388,N_8102,N_8238);
nand U8389 (N_8389,N_8112,N_8196);
xor U8390 (N_8390,N_8032,N_8069);
or U8391 (N_8391,N_8169,N_8086);
and U8392 (N_8392,N_8093,N_8046);
and U8393 (N_8393,N_8090,N_8067);
and U8394 (N_8394,N_8141,N_8187);
xor U8395 (N_8395,N_8061,N_8212);
and U8396 (N_8396,N_8202,N_8144);
xor U8397 (N_8397,N_8063,N_8069);
nor U8398 (N_8398,N_8017,N_8137);
and U8399 (N_8399,N_8179,N_8155);
or U8400 (N_8400,N_8134,N_8160);
xnor U8401 (N_8401,N_8102,N_8034);
or U8402 (N_8402,N_8131,N_8098);
xnor U8403 (N_8403,N_8063,N_8032);
nand U8404 (N_8404,N_8077,N_8160);
or U8405 (N_8405,N_8036,N_8009);
and U8406 (N_8406,N_8198,N_8235);
nor U8407 (N_8407,N_8147,N_8012);
nor U8408 (N_8408,N_8127,N_8015);
nand U8409 (N_8409,N_8160,N_8047);
nand U8410 (N_8410,N_8168,N_8136);
nor U8411 (N_8411,N_8099,N_8111);
xor U8412 (N_8412,N_8215,N_8073);
nand U8413 (N_8413,N_8065,N_8161);
xor U8414 (N_8414,N_8008,N_8186);
nor U8415 (N_8415,N_8004,N_8049);
xor U8416 (N_8416,N_8098,N_8204);
or U8417 (N_8417,N_8201,N_8123);
or U8418 (N_8418,N_8036,N_8141);
or U8419 (N_8419,N_8075,N_8239);
and U8420 (N_8420,N_8108,N_8185);
or U8421 (N_8421,N_8097,N_8042);
or U8422 (N_8422,N_8202,N_8098);
nor U8423 (N_8423,N_8028,N_8194);
xor U8424 (N_8424,N_8050,N_8121);
nand U8425 (N_8425,N_8208,N_8102);
nand U8426 (N_8426,N_8209,N_8119);
xor U8427 (N_8427,N_8142,N_8049);
nor U8428 (N_8428,N_8146,N_8029);
nor U8429 (N_8429,N_8081,N_8151);
or U8430 (N_8430,N_8093,N_8133);
nor U8431 (N_8431,N_8095,N_8246);
xnor U8432 (N_8432,N_8076,N_8070);
nor U8433 (N_8433,N_8198,N_8148);
nand U8434 (N_8434,N_8233,N_8033);
and U8435 (N_8435,N_8099,N_8043);
nand U8436 (N_8436,N_8134,N_8031);
nor U8437 (N_8437,N_8185,N_8083);
nor U8438 (N_8438,N_8125,N_8180);
nand U8439 (N_8439,N_8164,N_8074);
xor U8440 (N_8440,N_8173,N_8162);
xnor U8441 (N_8441,N_8027,N_8048);
nand U8442 (N_8442,N_8020,N_8128);
nor U8443 (N_8443,N_8167,N_8007);
or U8444 (N_8444,N_8170,N_8248);
xor U8445 (N_8445,N_8055,N_8119);
and U8446 (N_8446,N_8044,N_8227);
nand U8447 (N_8447,N_8012,N_8108);
and U8448 (N_8448,N_8136,N_8009);
and U8449 (N_8449,N_8114,N_8039);
or U8450 (N_8450,N_8230,N_8143);
and U8451 (N_8451,N_8018,N_8248);
and U8452 (N_8452,N_8108,N_8102);
xor U8453 (N_8453,N_8002,N_8105);
xnor U8454 (N_8454,N_8093,N_8106);
xor U8455 (N_8455,N_8053,N_8234);
or U8456 (N_8456,N_8051,N_8079);
and U8457 (N_8457,N_8193,N_8099);
nand U8458 (N_8458,N_8090,N_8218);
or U8459 (N_8459,N_8070,N_8213);
nand U8460 (N_8460,N_8075,N_8240);
nor U8461 (N_8461,N_8220,N_8172);
and U8462 (N_8462,N_8121,N_8130);
nand U8463 (N_8463,N_8168,N_8018);
nor U8464 (N_8464,N_8052,N_8236);
nand U8465 (N_8465,N_8121,N_8038);
nor U8466 (N_8466,N_8192,N_8082);
or U8467 (N_8467,N_8047,N_8126);
or U8468 (N_8468,N_8044,N_8171);
nor U8469 (N_8469,N_8246,N_8096);
xnor U8470 (N_8470,N_8249,N_8224);
xnor U8471 (N_8471,N_8033,N_8230);
and U8472 (N_8472,N_8208,N_8144);
or U8473 (N_8473,N_8043,N_8006);
or U8474 (N_8474,N_8099,N_8205);
and U8475 (N_8475,N_8098,N_8176);
nor U8476 (N_8476,N_8167,N_8105);
xor U8477 (N_8477,N_8131,N_8232);
xnor U8478 (N_8478,N_8189,N_8156);
nand U8479 (N_8479,N_8199,N_8046);
or U8480 (N_8480,N_8065,N_8090);
and U8481 (N_8481,N_8059,N_8098);
and U8482 (N_8482,N_8062,N_8244);
nor U8483 (N_8483,N_8014,N_8006);
nor U8484 (N_8484,N_8125,N_8074);
or U8485 (N_8485,N_8194,N_8026);
nor U8486 (N_8486,N_8247,N_8105);
or U8487 (N_8487,N_8113,N_8082);
xnor U8488 (N_8488,N_8202,N_8077);
and U8489 (N_8489,N_8196,N_8166);
nor U8490 (N_8490,N_8110,N_8198);
xor U8491 (N_8491,N_8174,N_8065);
nor U8492 (N_8492,N_8003,N_8011);
nor U8493 (N_8493,N_8077,N_8217);
nand U8494 (N_8494,N_8059,N_8123);
or U8495 (N_8495,N_8093,N_8047);
nand U8496 (N_8496,N_8010,N_8111);
nand U8497 (N_8497,N_8145,N_8207);
or U8498 (N_8498,N_8215,N_8242);
or U8499 (N_8499,N_8174,N_8218);
nand U8500 (N_8500,N_8497,N_8322);
xnor U8501 (N_8501,N_8345,N_8395);
or U8502 (N_8502,N_8296,N_8477);
nand U8503 (N_8503,N_8435,N_8338);
or U8504 (N_8504,N_8342,N_8368);
or U8505 (N_8505,N_8330,N_8311);
nor U8506 (N_8506,N_8366,N_8297);
or U8507 (N_8507,N_8286,N_8272);
nor U8508 (N_8508,N_8351,N_8472);
or U8509 (N_8509,N_8312,N_8495);
nand U8510 (N_8510,N_8421,N_8441);
nor U8511 (N_8511,N_8363,N_8352);
xor U8512 (N_8512,N_8498,N_8316);
xnor U8513 (N_8513,N_8479,N_8277);
xor U8514 (N_8514,N_8261,N_8336);
nor U8515 (N_8515,N_8431,N_8271);
nand U8516 (N_8516,N_8418,N_8433);
xor U8517 (N_8517,N_8458,N_8449);
nand U8518 (N_8518,N_8255,N_8374);
nand U8519 (N_8519,N_8460,N_8411);
nand U8520 (N_8520,N_8402,N_8343);
and U8521 (N_8521,N_8341,N_8378);
nand U8522 (N_8522,N_8388,N_8476);
and U8523 (N_8523,N_8422,N_8386);
or U8524 (N_8524,N_8492,N_8379);
and U8525 (N_8525,N_8425,N_8454);
xor U8526 (N_8526,N_8349,N_8359);
nor U8527 (N_8527,N_8387,N_8300);
or U8528 (N_8528,N_8485,N_8487);
nand U8529 (N_8529,N_8393,N_8302);
xnor U8530 (N_8530,N_8426,N_8265);
xnor U8531 (N_8531,N_8410,N_8438);
and U8532 (N_8532,N_8484,N_8467);
and U8533 (N_8533,N_8290,N_8461);
and U8534 (N_8534,N_8427,N_8450);
and U8535 (N_8535,N_8457,N_8278);
nand U8536 (N_8536,N_8397,N_8493);
nand U8537 (N_8537,N_8453,N_8321);
and U8538 (N_8538,N_8329,N_8443);
xnor U8539 (N_8539,N_8463,N_8376);
nor U8540 (N_8540,N_8417,N_8344);
nor U8541 (N_8541,N_8250,N_8496);
nand U8542 (N_8542,N_8263,N_8491);
nand U8543 (N_8543,N_8273,N_8464);
nand U8544 (N_8544,N_8478,N_8287);
nor U8545 (N_8545,N_8399,N_8456);
xor U8546 (N_8546,N_8306,N_8293);
or U8547 (N_8547,N_8358,N_8281);
or U8548 (N_8548,N_8253,N_8459);
or U8549 (N_8549,N_8434,N_8490);
or U8550 (N_8550,N_8309,N_8367);
or U8551 (N_8551,N_8414,N_8303);
xor U8552 (N_8552,N_8392,N_8371);
or U8553 (N_8553,N_8429,N_8373);
or U8554 (N_8554,N_8447,N_8408);
nor U8555 (N_8555,N_8331,N_8266);
xnor U8556 (N_8556,N_8276,N_8308);
xor U8557 (N_8557,N_8274,N_8357);
or U8558 (N_8558,N_8430,N_8282);
or U8559 (N_8559,N_8468,N_8326);
and U8560 (N_8560,N_8256,N_8314);
and U8561 (N_8561,N_8317,N_8365);
and U8562 (N_8562,N_8494,N_8470);
or U8563 (N_8563,N_8291,N_8318);
xnor U8564 (N_8564,N_8356,N_8424);
nand U8565 (N_8565,N_8489,N_8398);
nor U8566 (N_8566,N_8400,N_8334);
nand U8567 (N_8567,N_8324,N_8251);
nand U8568 (N_8568,N_8348,N_8471);
nor U8569 (N_8569,N_8375,N_8482);
nor U8570 (N_8570,N_8455,N_8279);
nand U8571 (N_8571,N_8262,N_8328);
nand U8572 (N_8572,N_8298,N_8372);
xor U8573 (N_8573,N_8369,N_8313);
nand U8574 (N_8574,N_8407,N_8275);
nand U8575 (N_8575,N_8416,N_8361);
xor U8576 (N_8576,N_8270,N_8269);
nand U8577 (N_8577,N_8258,N_8299);
nand U8578 (N_8578,N_8448,N_8315);
xor U8579 (N_8579,N_8267,N_8444);
xnor U8580 (N_8580,N_8486,N_8377);
nand U8581 (N_8581,N_8360,N_8499);
and U8582 (N_8582,N_8320,N_8442);
xor U8583 (N_8583,N_8339,N_8362);
xor U8584 (N_8584,N_8446,N_8335);
nor U8585 (N_8585,N_8288,N_8264);
nor U8586 (N_8586,N_8289,N_8346);
or U8587 (N_8587,N_8384,N_8404);
nand U8588 (N_8588,N_8268,N_8370);
and U8589 (N_8589,N_8340,N_8292);
nand U8590 (N_8590,N_8304,N_8383);
nor U8591 (N_8591,N_8380,N_8475);
or U8592 (N_8592,N_8428,N_8364);
or U8593 (N_8593,N_8480,N_8432);
xnor U8594 (N_8594,N_8252,N_8310);
and U8595 (N_8595,N_8403,N_8394);
nand U8596 (N_8596,N_8409,N_8469);
xor U8597 (N_8597,N_8285,N_8259);
nor U8598 (N_8598,N_8436,N_8415);
and U8599 (N_8599,N_8488,N_8355);
nor U8600 (N_8600,N_8257,N_8437);
xor U8601 (N_8601,N_8381,N_8473);
or U8602 (N_8602,N_8332,N_8353);
nand U8603 (N_8603,N_8445,N_8419);
nand U8604 (N_8604,N_8301,N_8307);
xnor U8605 (N_8605,N_8327,N_8350);
and U8606 (N_8606,N_8294,N_8405);
xnor U8607 (N_8607,N_8413,N_8333);
nand U8608 (N_8608,N_8465,N_8483);
or U8609 (N_8609,N_8323,N_8466);
xor U8610 (N_8610,N_8406,N_8325);
and U8611 (N_8611,N_8385,N_8390);
nand U8612 (N_8612,N_8481,N_8391);
and U8613 (N_8613,N_8283,N_8474);
nor U8614 (N_8614,N_8319,N_8462);
or U8615 (N_8615,N_8423,N_8347);
nor U8616 (N_8616,N_8439,N_8280);
nor U8617 (N_8617,N_8260,N_8337);
xor U8618 (N_8618,N_8440,N_8401);
nand U8619 (N_8619,N_8451,N_8452);
nand U8620 (N_8620,N_8284,N_8389);
xnor U8621 (N_8621,N_8412,N_8396);
nor U8622 (N_8622,N_8354,N_8382);
xor U8623 (N_8623,N_8295,N_8420);
and U8624 (N_8624,N_8254,N_8305);
nand U8625 (N_8625,N_8489,N_8480);
and U8626 (N_8626,N_8416,N_8309);
nand U8627 (N_8627,N_8350,N_8464);
xnor U8628 (N_8628,N_8374,N_8359);
xnor U8629 (N_8629,N_8385,N_8266);
or U8630 (N_8630,N_8358,N_8431);
or U8631 (N_8631,N_8334,N_8441);
or U8632 (N_8632,N_8365,N_8384);
or U8633 (N_8633,N_8366,N_8422);
xnor U8634 (N_8634,N_8323,N_8434);
nor U8635 (N_8635,N_8350,N_8283);
and U8636 (N_8636,N_8419,N_8411);
nand U8637 (N_8637,N_8490,N_8421);
and U8638 (N_8638,N_8338,N_8292);
and U8639 (N_8639,N_8304,N_8293);
nand U8640 (N_8640,N_8455,N_8399);
xor U8641 (N_8641,N_8469,N_8476);
xnor U8642 (N_8642,N_8282,N_8411);
xnor U8643 (N_8643,N_8329,N_8372);
nor U8644 (N_8644,N_8492,N_8288);
and U8645 (N_8645,N_8358,N_8332);
xnor U8646 (N_8646,N_8342,N_8350);
or U8647 (N_8647,N_8310,N_8340);
xor U8648 (N_8648,N_8469,N_8293);
and U8649 (N_8649,N_8313,N_8406);
or U8650 (N_8650,N_8491,N_8414);
nand U8651 (N_8651,N_8392,N_8468);
and U8652 (N_8652,N_8490,N_8269);
and U8653 (N_8653,N_8350,N_8365);
xor U8654 (N_8654,N_8343,N_8264);
xor U8655 (N_8655,N_8306,N_8395);
nand U8656 (N_8656,N_8451,N_8474);
xor U8657 (N_8657,N_8333,N_8389);
and U8658 (N_8658,N_8304,N_8385);
nor U8659 (N_8659,N_8282,N_8408);
nor U8660 (N_8660,N_8311,N_8399);
xor U8661 (N_8661,N_8420,N_8399);
nand U8662 (N_8662,N_8489,N_8435);
and U8663 (N_8663,N_8297,N_8343);
and U8664 (N_8664,N_8440,N_8313);
and U8665 (N_8665,N_8295,N_8293);
or U8666 (N_8666,N_8368,N_8339);
and U8667 (N_8667,N_8476,N_8405);
xnor U8668 (N_8668,N_8416,N_8301);
and U8669 (N_8669,N_8357,N_8406);
nand U8670 (N_8670,N_8327,N_8482);
nor U8671 (N_8671,N_8345,N_8436);
or U8672 (N_8672,N_8269,N_8432);
or U8673 (N_8673,N_8435,N_8458);
nand U8674 (N_8674,N_8407,N_8346);
nor U8675 (N_8675,N_8321,N_8480);
nor U8676 (N_8676,N_8360,N_8416);
nand U8677 (N_8677,N_8378,N_8377);
or U8678 (N_8678,N_8349,N_8480);
or U8679 (N_8679,N_8467,N_8258);
and U8680 (N_8680,N_8296,N_8393);
or U8681 (N_8681,N_8424,N_8410);
or U8682 (N_8682,N_8309,N_8319);
xor U8683 (N_8683,N_8378,N_8388);
xor U8684 (N_8684,N_8474,N_8473);
nand U8685 (N_8685,N_8332,N_8348);
xnor U8686 (N_8686,N_8270,N_8378);
and U8687 (N_8687,N_8447,N_8271);
nor U8688 (N_8688,N_8315,N_8365);
and U8689 (N_8689,N_8477,N_8366);
xnor U8690 (N_8690,N_8379,N_8330);
nor U8691 (N_8691,N_8442,N_8257);
nand U8692 (N_8692,N_8298,N_8414);
and U8693 (N_8693,N_8275,N_8463);
nor U8694 (N_8694,N_8367,N_8277);
nand U8695 (N_8695,N_8306,N_8493);
and U8696 (N_8696,N_8450,N_8277);
or U8697 (N_8697,N_8486,N_8348);
xor U8698 (N_8698,N_8290,N_8266);
xnor U8699 (N_8699,N_8396,N_8274);
nor U8700 (N_8700,N_8483,N_8469);
nand U8701 (N_8701,N_8463,N_8374);
nor U8702 (N_8702,N_8384,N_8443);
and U8703 (N_8703,N_8349,N_8371);
nor U8704 (N_8704,N_8329,N_8363);
xnor U8705 (N_8705,N_8267,N_8326);
nand U8706 (N_8706,N_8321,N_8486);
nor U8707 (N_8707,N_8419,N_8342);
nand U8708 (N_8708,N_8378,N_8409);
nand U8709 (N_8709,N_8483,N_8467);
xor U8710 (N_8710,N_8348,N_8334);
nand U8711 (N_8711,N_8377,N_8365);
nor U8712 (N_8712,N_8462,N_8395);
nor U8713 (N_8713,N_8470,N_8411);
nand U8714 (N_8714,N_8468,N_8365);
xor U8715 (N_8715,N_8396,N_8400);
nand U8716 (N_8716,N_8352,N_8334);
nor U8717 (N_8717,N_8434,N_8388);
nand U8718 (N_8718,N_8404,N_8291);
and U8719 (N_8719,N_8308,N_8293);
nor U8720 (N_8720,N_8299,N_8313);
or U8721 (N_8721,N_8252,N_8386);
or U8722 (N_8722,N_8323,N_8305);
or U8723 (N_8723,N_8306,N_8353);
xnor U8724 (N_8724,N_8482,N_8394);
nand U8725 (N_8725,N_8496,N_8255);
nand U8726 (N_8726,N_8382,N_8331);
nor U8727 (N_8727,N_8491,N_8319);
or U8728 (N_8728,N_8478,N_8472);
nand U8729 (N_8729,N_8327,N_8330);
or U8730 (N_8730,N_8398,N_8467);
xnor U8731 (N_8731,N_8498,N_8351);
xor U8732 (N_8732,N_8435,N_8305);
or U8733 (N_8733,N_8447,N_8482);
nor U8734 (N_8734,N_8464,N_8267);
and U8735 (N_8735,N_8300,N_8459);
and U8736 (N_8736,N_8267,N_8339);
and U8737 (N_8737,N_8388,N_8252);
xor U8738 (N_8738,N_8410,N_8279);
or U8739 (N_8739,N_8254,N_8338);
xnor U8740 (N_8740,N_8253,N_8361);
and U8741 (N_8741,N_8262,N_8274);
nand U8742 (N_8742,N_8490,N_8305);
nand U8743 (N_8743,N_8337,N_8316);
nand U8744 (N_8744,N_8389,N_8264);
and U8745 (N_8745,N_8359,N_8341);
xor U8746 (N_8746,N_8270,N_8395);
nand U8747 (N_8747,N_8434,N_8498);
nor U8748 (N_8748,N_8369,N_8271);
xnor U8749 (N_8749,N_8373,N_8404);
nor U8750 (N_8750,N_8743,N_8527);
and U8751 (N_8751,N_8723,N_8565);
or U8752 (N_8752,N_8688,N_8728);
and U8753 (N_8753,N_8732,N_8513);
or U8754 (N_8754,N_8611,N_8654);
nand U8755 (N_8755,N_8550,N_8626);
xor U8756 (N_8756,N_8543,N_8710);
nand U8757 (N_8757,N_8713,N_8556);
or U8758 (N_8758,N_8555,N_8532);
xnor U8759 (N_8759,N_8623,N_8712);
nor U8760 (N_8760,N_8718,N_8722);
nor U8761 (N_8761,N_8515,N_8686);
xor U8762 (N_8762,N_8531,N_8707);
or U8763 (N_8763,N_8501,N_8733);
nor U8764 (N_8764,N_8639,N_8582);
and U8765 (N_8765,N_8680,N_8508);
or U8766 (N_8766,N_8689,N_8641);
nand U8767 (N_8767,N_8627,N_8669);
or U8768 (N_8768,N_8603,N_8534);
xor U8769 (N_8769,N_8505,N_8564);
nor U8770 (N_8770,N_8706,N_8574);
xor U8771 (N_8771,N_8636,N_8651);
or U8772 (N_8772,N_8648,N_8642);
or U8773 (N_8773,N_8570,N_8700);
xnor U8774 (N_8774,N_8609,N_8561);
or U8775 (N_8775,N_8553,N_8587);
nor U8776 (N_8776,N_8682,N_8640);
or U8777 (N_8777,N_8579,N_8568);
nand U8778 (N_8778,N_8672,N_8657);
nand U8779 (N_8779,N_8719,N_8649);
or U8780 (N_8780,N_8738,N_8591);
nand U8781 (N_8781,N_8677,N_8745);
xor U8782 (N_8782,N_8542,N_8646);
or U8783 (N_8783,N_8716,N_8573);
nor U8784 (N_8784,N_8597,N_8662);
or U8785 (N_8785,N_8504,N_8638);
nor U8786 (N_8786,N_8666,N_8506);
or U8787 (N_8787,N_8607,N_8625);
or U8788 (N_8788,N_8678,N_8746);
xnor U8789 (N_8789,N_8604,N_8530);
nor U8790 (N_8790,N_8708,N_8509);
and U8791 (N_8791,N_8599,N_8727);
xor U8792 (N_8792,N_8747,N_8588);
and U8793 (N_8793,N_8724,N_8748);
nor U8794 (N_8794,N_8720,N_8537);
and U8795 (N_8795,N_8517,N_8554);
and U8796 (N_8796,N_8549,N_8668);
or U8797 (N_8797,N_8528,N_8575);
nor U8798 (N_8798,N_8730,N_8526);
and U8799 (N_8799,N_8551,N_8659);
and U8800 (N_8800,N_8613,N_8622);
nand U8801 (N_8801,N_8578,N_8619);
xnor U8802 (N_8802,N_8698,N_8624);
nor U8803 (N_8803,N_8630,N_8637);
nor U8804 (N_8804,N_8699,N_8692);
nor U8805 (N_8805,N_8594,N_8545);
xnor U8806 (N_8806,N_8548,N_8695);
or U8807 (N_8807,N_8691,N_8671);
and U8808 (N_8808,N_8701,N_8581);
or U8809 (N_8809,N_8563,N_8664);
and U8810 (N_8810,N_8584,N_8737);
or U8811 (N_8811,N_8559,N_8608);
nand U8812 (N_8812,N_8679,N_8705);
or U8813 (N_8813,N_8523,N_8616);
nand U8814 (N_8814,N_8596,N_8725);
and U8815 (N_8815,N_8661,N_8512);
or U8816 (N_8816,N_8557,N_8602);
nor U8817 (N_8817,N_8562,N_8632);
and U8818 (N_8818,N_8676,N_8572);
xnor U8819 (N_8819,N_8538,N_8714);
and U8820 (N_8820,N_8577,N_8580);
nand U8821 (N_8821,N_8711,N_8703);
nor U8822 (N_8822,N_8566,N_8631);
nand U8823 (N_8823,N_8629,N_8734);
and U8824 (N_8824,N_8628,N_8735);
nand U8825 (N_8825,N_8558,N_8620);
xor U8826 (N_8826,N_8571,N_8618);
xnor U8827 (N_8827,N_8600,N_8612);
nand U8828 (N_8828,N_8583,N_8576);
nor U8829 (N_8829,N_8541,N_8511);
nor U8830 (N_8830,N_8552,N_8655);
nand U8831 (N_8831,N_8749,N_8521);
nand U8832 (N_8832,N_8593,N_8643);
nand U8833 (N_8833,N_8653,N_8697);
xnor U8834 (N_8834,N_8633,N_8634);
nor U8835 (N_8835,N_8673,N_8665);
nor U8836 (N_8836,N_8614,N_8739);
nand U8837 (N_8837,N_8721,N_8670);
or U8838 (N_8838,N_8507,N_8717);
nor U8839 (N_8839,N_8621,N_8687);
and U8840 (N_8840,N_8740,N_8742);
nand U8841 (N_8841,N_8533,N_8585);
nor U8842 (N_8842,N_8544,N_8610);
and U8843 (N_8843,N_8715,N_8606);
nand U8844 (N_8844,N_8503,N_8589);
nand U8845 (N_8845,N_8518,N_8536);
nand U8846 (N_8846,N_8617,N_8519);
xor U8847 (N_8847,N_8598,N_8693);
and U8848 (N_8848,N_8726,N_8510);
nor U8849 (N_8849,N_8529,N_8685);
nand U8850 (N_8850,N_8516,N_8595);
nor U8851 (N_8851,N_8667,N_8635);
and U8852 (N_8852,N_8681,N_8709);
nor U8853 (N_8853,N_8500,N_8615);
nand U8854 (N_8854,N_8663,N_8656);
nor U8855 (N_8855,N_8684,N_8702);
nand U8856 (N_8856,N_8652,N_8683);
and U8857 (N_8857,N_8694,N_8569);
nor U8858 (N_8858,N_8675,N_8744);
and U8859 (N_8859,N_8586,N_8524);
and U8860 (N_8860,N_8658,N_8736);
and U8861 (N_8861,N_8567,N_8704);
or U8862 (N_8862,N_8645,N_8592);
xnor U8863 (N_8863,N_8650,N_8546);
or U8864 (N_8864,N_8644,N_8605);
xnor U8865 (N_8865,N_8560,N_8590);
xnor U8866 (N_8866,N_8514,N_8674);
and U8867 (N_8867,N_8696,N_8690);
or U8868 (N_8868,N_8741,N_8647);
nand U8869 (N_8869,N_8660,N_8502);
nand U8870 (N_8870,N_8520,N_8539);
or U8871 (N_8871,N_8535,N_8547);
xor U8872 (N_8872,N_8522,N_8601);
xor U8873 (N_8873,N_8525,N_8731);
nand U8874 (N_8874,N_8729,N_8540);
nand U8875 (N_8875,N_8639,N_8650);
xnor U8876 (N_8876,N_8637,N_8732);
or U8877 (N_8877,N_8586,N_8636);
or U8878 (N_8878,N_8718,N_8563);
nor U8879 (N_8879,N_8729,N_8632);
nand U8880 (N_8880,N_8722,N_8573);
nand U8881 (N_8881,N_8717,N_8542);
or U8882 (N_8882,N_8578,N_8713);
xor U8883 (N_8883,N_8541,N_8588);
and U8884 (N_8884,N_8547,N_8662);
or U8885 (N_8885,N_8730,N_8587);
xnor U8886 (N_8886,N_8660,N_8626);
xor U8887 (N_8887,N_8591,N_8655);
or U8888 (N_8888,N_8526,N_8626);
nand U8889 (N_8889,N_8578,N_8509);
or U8890 (N_8890,N_8528,N_8504);
or U8891 (N_8891,N_8543,N_8741);
and U8892 (N_8892,N_8656,N_8646);
xor U8893 (N_8893,N_8579,N_8673);
nand U8894 (N_8894,N_8610,N_8607);
nand U8895 (N_8895,N_8712,N_8671);
nand U8896 (N_8896,N_8684,N_8627);
or U8897 (N_8897,N_8534,N_8575);
and U8898 (N_8898,N_8674,N_8692);
nand U8899 (N_8899,N_8517,N_8500);
nand U8900 (N_8900,N_8621,N_8544);
nor U8901 (N_8901,N_8536,N_8723);
and U8902 (N_8902,N_8688,N_8738);
or U8903 (N_8903,N_8714,N_8721);
and U8904 (N_8904,N_8655,N_8725);
and U8905 (N_8905,N_8504,N_8748);
and U8906 (N_8906,N_8530,N_8589);
xor U8907 (N_8907,N_8581,N_8724);
and U8908 (N_8908,N_8670,N_8719);
and U8909 (N_8909,N_8653,N_8611);
xor U8910 (N_8910,N_8680,N_8585);
xnor U8911 (N_8911,N_8717,N_8683);
or U8912 (N_8912,N_8710,N_8512);
xnor U8913 (N_8913,N_8609,N_8714);
nand U8914 (N_8914,N_8505,N_8704);
nor U8915 (N_8915,N_8573,N_8547);
and U8916 (N_8916,N_8585,N_8527);
nor U8917 (N_8917,N_8614,N_8627);
or U8918 (N_8918,N_8674,N_8633);
or U8919 (N_8919,N_8651,N_8517);
nor U8920 (N_8920,N_8671,N_8591);
nor U8921 (N_8921,N_8659,N_8612);
nor U8922 (N_8922,N_8530,N_8700);
or U8923 (N_8923,N_8569,N_8547);
nand U8924 (N_8924,N_8644,N_8519);
nor U8925 (N_8925,N_8732,N_8558);
or U8926 (N_8926,N_8501,N_8619);
nand U8927 (N_8927,N_8741,N_8600);
and U8928 (N_8928,N_8552,N_8559);
nor U8929 (N_8929,N_8746,N_8646);
nor U8930 (N_8930,N_8531,N_8534);
xor U8931 (N_8931,N_8526,N_8603);
xnor U8932 (N_8932,N_8574,N_8604);
nor U8933 (N_8933,N_8722,N_8506);
xnor U8934 (N_8934,N_8705,N_8670);
nor U8935 (N_8935,N_8734,N_8695);
xnor U8936 (N_8936,N_8632,N_8731);
or U8937 (N_8937,N_8600,N_8599);
xor U8938 (N_8938,N_8641,N_8540);
nand U8939 (N_8939,N_8599,N_8709);
xnor U8940 (N_8940,N_8528,N_8596);
or U8941 (N_8941,N_8586,N_8679);
nand U8942 (N_8942,N_8619,N_8738);
and U8943 (N_8943,N_8743,N_8719);
xnor U8944 (N_8944,N_8649,N_8651);
nand U8945 (N_8945,N_8699,N_8558);
xnor U8946 (N_8946,N_8649,N_8601);
nand U8947 (N_8947,N_8593,N_8649);
nand U8948 (N_8948,N_8582,N_8528);
and U8949 (N_8949,N_8664,N_8745);
xor U8950 (N_8950,N_8651,N_8660);
or U8951 (N_8951,N_8722,N_8697);
nand U8952 (N_8952,N_8625,N_8577);
nand U8953 (N_8953,N_8576,N_8738);
nor U8954 (N_8954,N_8740,N_8628);
xnor U8955 (N_8955,N_8649,N_8576);
or U8956 (N_8956,N_8713,N_8634);
nor U8957 (N_8957,N_8693,N_8676);
nor U8958 (N_8958,N_8704,N_8529);
or U8959 (N_8959,N_8525,N_8622);
nor U8960 (N_8960,N_8545,N_8659);
nand U8961 (N_8961,N_8657,N_8707);
or U8962 (N_8962,N_8629,N_8745);
and U8963 (N_8963,N_8576,N_8715);
nand U8964 (N_8964,N_8517,N_8693);
xnor U8965 (N_8965,N_8510,N_8644);
xnor U8966 (N_8966,N_8541,N_8529);
nand U8967 (N_8967,N_8717,N_8731);
and U8968 (N_8968,N_8593,N_8658);
nor U8969 (N_8969,N_8519,N_8591);
nand U8970 (N_8970,N_8621,N_8525);
nand U8971 (N_8971,N_8661,N_8559);
xor U8972 (N_8972,N_8646,N_8633);
xor U8973 (N_8973,N_8548,N_8540);
or U8974 (N_8974,N_8725,N_8621);
nor U8975 (N_8975,N_8740,N_8510);
xnor U8976 (N_8976,N_8651,N_8543);
or U8977 (N_8977,N_8615,N_8613);
nand U8978 (N_8978,N_8642,N_8568);
and U8979 (N_8979,N_8584,N_8650);
xor U8980 (N_8980,N_8747,N_8643);
xor U8981 (N_8981,N_8531,N_8511);
nand U8982 (N_8982,N_8745,N_8549);
and U8983 (N_8983,N_8652,N_8542);
nor U8984 (N_8984,N_8666,N_8565);
nor U8985 (N_8985,N_8685,N_8515);
xor U8986 (N_8986,N_8672,N_8650);
nand U8987 (N_8987,N_8629,N_8527);
xnor U8988 (N_8988,N_8649,N_8588);
nand U8989 (N_8989,N_8504,N_8622);
nand U8990 (N_8990,N_8701,N_8572);
nor U8991 (N_8991,N_8580,N_8687);
xnor U8992 (N_8992,N_8501,N_8627);
or U8993 (N_8993,N_8740,N_8616);
xor U8994 (N_8994,N_8574,N_8739);
and U8995 (N_8995,N_8692,N_8715);
xnor U8996 (N_8996,N_8706,N_8516);
nand U8997 (N_8997,N_8649,N_8688);
nand U8998 (N_8998,N_8527,N_8552);
or U8999 (N_8999,N_8588,N_8571);
and U9000 (N_9000,N_8845,N_8859);
nand U9001 (N_9001,N_8902,N_8912);
or U9002 (N_9002,N_8883,N_8875);
nor U9003 (N_9003,N_8795,N_8932);
nor U9004 (N_9004,N_8942,N_8980);
xor U9005 (N_9005,N_8950,N_8807);
xnor U9006 (N_9006,N_8931,N_8789);
xor U9007 (N_9007,N_8787,N_8842);
xnor U9008 (N_9008,N_8753,N_8802);
or U9009 (N_9009,N_8885,N_8974);
and U9010 (N_9010,N_8817,N_8997);
xor U9011 (N_9011,N_8949,N_8811);
nand U9012 (N_9012,N_8969,N_8962);
nand U9013 (N_9013,N_8994,N_8840);
xor U9014 (N_9014,N_8781,N_8979);
nor U9015 (N_9015,N_8884,N_8854);
xor U9016 (N_9016,N_8768,N_8846);
nor U9017 (N_9017,N_8847,N_8995);
nand U9018 (N_9018,N_8867,N_8920);
nor U9019 (N_9019,N_8798,N_8864);
or U9020 (N_9020,N_8946,N_8973);
xor U9021 (N_9021,N_8900,N_8861);
and U9022 (N_9022,N_8830,N_8794);
nor U9023 (N_9023,N_8917,N_8869);
or U9024 (N_9024,N_8848,N_8851);
xor U9025 (N_9025,N_8831,N_8919);
xnor U9026 (N_9026,N_8907,N_8956);
and U9027 (N_9027,N_8750,N_8903);
and U9028 (N_9028,N_8982,N_8918);
or U9029 (N_9029,N_8836,N_8799);
and U9030 (N_9030,N_8924,N_8893);
nand U9031 (N_9031,N_8986,N_8769);
or U9032 (N_9032,N_8923,N_8780);
nand U9033 (N_9033,N_8987,N_8877);
and U9034 (N_9034,N_8977,N_8911);
nor U9035 (N_9035,N_8910,N_8758);
xnor U9036 (N_9036,N_8975,N_8819);
and U9037 (N_9037,N_8870,N_8872);
or U9038 (N_9038,N_8958,N_8981);
or U9039 (N_9039,N_8887,N_8940);
or U9040 (N_9040,N_8897,N_8952);
nor U9041 (N_9041,N_8808,N_8921);
nor U9042 (N_9042,N_8909,N_8783);
nand U9043 (N_9043,N_8810,N_8823);
or U9044 (N_9044,N_8880,N_8757);
or U9045 (N_9045,N_8820,N_8844);
and U9046 (N_9046,N_8879,N_8760);
or U9047 (N_9047,N_8908,N_8983);
xnor U9048 (N_9048,N_8825,N_8906);
xnor U9049 (N_9049,N_8899,N_8855);
and U9050 (N_9050,N_8863,N_8796);
or U9051 (N_9051,N_8874,N_8775);
xor U9052 (N_9052,N_8927,N_8866);
xor U9053 (N_9053,N_8770,N_8901);
nor U9054 (N_9054,N_8764,N_8925);
xnor U9055 (N_9055,N_8793,N_8826);
nor U9056 (N_9056,N_8878,N_8941);
xor U9057 (N_9057,N_8970,N_8773);
or U9058 (N_9058,N_8961,N_8858);
nor U9059 (N_9059,N_8754,N_8957);
nand U9060 (N_9060,N_8837,N_8882);
or U9061 (N_9061,N_8841,N_8803);
nand U9062 (N_9062,N_8776,N_8865);
nand U9063 (N_9063,N_8971,N_8938);
nor U9064 (N_9064,N_8944,N_8800);
and U9065 (N_9065,N_8822,N_8976);
xnor U9066 (N_9066,N_8945,N_8955);
nand U9067 (N_9067,N_8838,N_8934);
or U9068 (N_9068,N_8774,N_8862);
or U9069 (N_9069,N_8896,N_8886);
nor U9070 (N_9070,N_8812,N_8892);
nand U9071 (N_9071,N_8937,N_8929);
or U9072 (N_9072,N_8939,N_8778);
xor U9073 (N_9073,N_8876,N_8806);
and U9074 (N_9074,N_8914,N_8960);
or U9075 (N_9075,N_8992,N_8972);
nor U9076 (N_9076,N_8821,N_8894);
or U9077 (N_9077,N_8813,N_8756);
nand U9078 (N_9078,N_8978,N_8948);
nor U9079 (N_9079,N_8833,N_8857);
and U9080 (N_9080,N_8791,N_8834);
and U9081 (N_9081,N_8759,N_8943);
nor U9082 (N_9082,N_8809,N_8933);
or U9083 (N_9083,N_8904,N_8930);
or U9084 (N_9084,N_8829,N_8751);
xnor U9085 (N_9085,N_8965,N_8990);
nor U9086 (N_9086,N_8832,N_8963);
or U9087 (N_9087,N_8755,N_8853);
nand U9088 (N_9088,N_8849,N_8788);
and U9089 (N_9089,N_8889,N_8989);
nor U9090 (N_9090,N_8905,N_8947);
and U9091 (N_9091,N_8797,N_8922);
nand U9092 (N_9092,N_8763,N_8890);
or U9093 (N_9093,N_8785,N_8777);
xor U9094 (N_9094,N_8765,N_8815);
nor U9095 (N_9095,N_8839,N_8964);
nor U9096 (N_9096,N_8850,N_8993);
nor U9097 (N_9097,N_8860,N_8998);
xor U9098 (N_9098,N_8843,N_8784);
xnor U9099 (N_9099,N_8873,N_8868);
or U9100 (N_9100,N_8951,N_8772);
xnor U9101 (N_9101,N_8782,N_8752);
and U9102 (N_9102,N_8953,N_8814);
and U9103 (N_9103,N_8888,N_8928);
nor U9104 (N_9104,N_8805,N_8895);
or U9105 (N_9105,N_8816,N_8792);
and U9106 (N_9106,N_8881,N_8835);
nor U9107 (N_9107,N_8779,N_8801);
nand U9108 (N_9108,N_8828,N_8968);
and U9109 (N_9109,N_8824,N_8891);
xor U9110 (N_9110,N_8988,N_8954);
or U9111 (N_9111,N_8871,N_8898);
xor U9112 (N_9112,N_8915,N_8818);
nand U9113 (N_9113,N_8856,N_8936);
xnor U9114 (N_9114,N_8984,N_8852);
xor U9115 (N_9115,N_8766,N_8991);
or U9116 (N_9116,N_8926,N_8804);
xnor U9117 (N_9117,N_8913,N_8767);
or U9118 (N_9118,N_8966,N_8771);
or U9119 (N_9119,N_8935,N_8827);
nand U9120 (N_9120,N_8786,N_8916);
or U9121 (N_9121,N_8790,N_8996);
nand U9122 (N_9122,N_8761,N_8967);
and U9123 (N_9123,N_8959,N_8985);
nor U9124 (N_9124,N_8762,N_8999);
nor U9125 (N_9125,N_8779,N_8915);
nor U9126 (N_9126,N_8831,N_8763);
nor U9127 (N_9127,N_8837,N_8766);
nor U9128 (N_9128,N_8869,N_8914);
nand U9129 (N_9129,N_8788,N_8873);
or U9130 (N_9130,N_8909,N_8860);
and U9131 (N_9131,N_8976,N_8791);
xor U9132 (N_9132,N_8896,N_8898);
and U9133 (N_9133,N_8933,N_8843);
or U9134 (N_9134,N_8780,N_8959);
or U9135 (N_9135,N_8950,N_8765);
nand U9136 (N_9136,N_8860,N_8894);
nand U9137 (N_9137,N_8801,N_8797);
nand U9138 (N_9138,N_8934,N_8908);
and U9139 (N_9139,N_8997,N_8899);
xor U9140 (N_9140,N_8986,N_8938);
nand U9141 (N_9141,N_8935,N_8978);
and U9142 (N_9142,N_8857,N_8877);
nor U9143 (N_9143,N_8783,N_8890);
nand U9144 (N_9144,N_8957,N_8861);
nand U9145 (N_9145,N_8929,N_8847);
nand U9146 (N_9146,N_8767,N_8938);
or U9147 (N_9147,N_8905,N_8858);
nor U9148 (N_9148,N_8839,N_8756);
nand U9149 (N_9149,N_8804,N_8886);
xnor U9150 (N_9150,N_8904,N_8781);
xor U9151 (N_9151,N_8861,N_8822);
xnor U9152 (N_9152,N_8782,N_8879);
and U9153 (N_9153,N_8957,N_8997);
nand U9154 (N_9154,N_8994,N_8986);
xnor U9155 (N_9155,N_8750,N_8782);
xor U9156 (N_9156,N_8913,N_8857);
or U9157 (N_9157,N_8988,N_8909);
xor U9158 (N_9158,N_8847,N_8834);
xnor U9159 (N_9159,N_8814,N_8975);
nor U9160 (N_9160,N_8825,N_8772);
or U9161 (N_9161,N_8964,N_8961);
xor U9162 (N_9162,N_8907,N_8981);
nand U9163 (N_9163,N_8982,N_8799);
and U9164 (N_9164,N_8855,N_8915);
and U9165 (N_9165,N_8831,N_8861);
or U9166 (N_9166,N_8873,N_8850);
and U9167 (N_9167,N_8817,N_8937);
nand U9168 (N_9168,N_8942,N_8936);
or U9169 (N_9169,N_8960,N_8861);
or U9170 (N_9170,N_8765,N_8813);
and U9171 (N_9171,N_8852,N_8949);
nand U9172 (N_9172,N_8772,N_8945);
nand U9173 (N_9173,N_8858,N_8754);
xnor U9174 (N_9174,N_8991,N_8804);
or U9175 (N_9175,N_8961,N_8870);
or U9176 (N_9176,N_8937,N_8920);
nand U9177 (N_9177,N_8865,N_8883);
or U9178 (N_9178,N_8931,N_8908);
or U9179 (N_9179,N_8903,N_8826);
and U9180 (N_9180,N_8860,N_8851);
and U9181 (N_9181,N_8921,N_8786);
xnor U9182 (N_9182,N_8778,N_8815);
nand U9183 (N_9183,N_8796,N_8780);
nor U9184 (N_9184,N_8803,N_8844);
xor U9185 (N_9185,N_8984,N_8772);
xor U9186 (N_9186,N_8863,N_8806);
xnor U9187 (N_9187,N_8852,N_8773);
or U9188 (N_9188,N_8814,N_8848);
or U9189 (N_9189,N_8962,N_8857);
or U9190 (N_9190,N_8831,N_8820);
xnor U9191 (N_9191,N_8925,N_8795);
nand U9192 (N_9192,N_8990,N_8930);
or U9193 (N_9193,N_8954,N_8991);
and U9194 (N_9194,N_8879,N_8815);
or U9195 (N_9195,N_8953,N_8887);
nand U9196 (N_9196,N_8931,N_8952);
nor U9197 (N_9197,N_8861,N_8806);
nand U9198 (N_9198,N_8921,N_8980);
and U9199 (N_9199,N_8918,N_8965);
nor U9200 (N_9200,N_8874,N_8783);
nor U9201 (N_9201,N_8915,N_8825);
and U9202 (N_9202,N_8752,N_8882);
nor U9203 (N_9203,N_8817,N_8924);
or U9204 (N_9204,N_8998,N_8863);
or U9205 (N_9205,N_8970,N_8796);
nor U9206 (N_9206,N_8800,N_8967);
nand U9207 (N_9207,N_8933,N_8815);
and U9208 (N_9208,N_8996,N_8783);
xor U9209 (N_9209,N_8873,N_8915);
and U9210 (N_9210,N_8942,N_8911);
or U9211 (N_9211,N_8849,N_8903);
nor U9212 (N_9212,N_8971,N_8945);
nand U9213 (N_9213,N_8988,N_8754);
or U9214 (N_9214,N_8918,N_8753);
nand U9215 (N_9215,N_8995,N_8764);
xnor U9216 (N_9216,N_8812,N_8848);
xnor U9217 (N_9217,N_8797,N_8826);
nor U9218 (N_9218,N_8810,N_8796);
or U9219 (N_9219,N_8805,N_8913);
nand U9220 (N_9220,N_8843,N_8967);
nand U9221 (N_9221,N_8832,N_8856);
and U9222 (N_9222,N_8828,N_8860);
or U9223 (N_9223,N_8891,N_8902);
and U9224 (N_9224,N_8948,N_8812);
nand U9225 (N_9225,N_8951,N_8775);
nand U9226 (N_9226,N_8820,N_8986);
and U9227 (N_9227,N_8924,N_8796);
nand U9228 (N_9228,N_8928,N_8918);
nor U9229 (N_9229,N_8917,N_8973);
nor U9230 (N_9230,N_8793,N_8984);
or U9231 (N_9231,N_8995,N_8776);
nand U9232 (N_9232,N_8955,N_8844);
and U9233 (N_9233,N_8833,N_8868);
xnor U9234 (N_9234,N_8979,N_8954);
and U9235 (N_9235,N_8803,N_8819);
nor U9236 (N_9236,N_8840,N_8751);
nand U9237 (N_9237,N_8957,N_8945);
xnor U9238 (N_9238,N_8880,N_8899);
xor U9239 (N_9239,N_8972,N_8952);
nor U9240 (N_9240,N_8982,N_8939);
nand U9241 (N_9241,N_8949,N_8869);
and U9242 (N_9242,N_8847,N_8820);
or U9243 (N_9243,N_8930,N_8931);
or U9244 (N_9244,N_8853,N_8943);
xor U9245 (N_9245,N_8940,N_8756);
xor U9246 (N_9246,N_8939,N_8923);
or U9247 (N_9247,N_8894,N_8923);
nor U9248 (N_9248,N_8937,N_8829);
nor U9249 (N_9249,N_8798,N_8757);
or U9250 (N_9250,N_9099,N_9025);
xor U9251 (N_9251,N_9147,N_9164);
or U9252 (N_9252,N_9110,N_9015);
xnor U9253 (N_9253,N_9105,N_9121);
xnor U9254 (N_9254,N_9136,N_9095);
nor U9255 (N_9255,N_9034,N_9031);
nand U9256 (N_9256,N_9010,N_9063);
nor U9257 (N_9257,N_9238,N_9093);
nand U9258 (N_9258,N_9175,N_9038);
or U9259 (N_9259,N_9155,N_9132);
and U9260 (N_9260,N_9204,N_9165);
nand U9261 (N_9261,N_9094,N_9070);
or U9262 (N_9262,N_9080,N_9153);
nor U9263 (N_9263,N_9124,N_9211);
nor U9264 (N_9264,N_9189,N_9233);
nor U9265 (N_9265,N_9019,N_9041);
and U9266 (N_9266,N_9247,N_9225);
xor U9267 (N_9267,N_9018,N_9188);
nand U9268 (N_9268,N_9023,N_9008);
nor U9269 (N_9269,N_9020,N_9213);
and U9270 (N_9270,N_9221,N_9079);
or U9271 (N_9271,N_9214,N_9119);
xnor U9272 (N_9272,N_9172,N_9064);
nand U9273 (N_9273,N_9006,N_9026);
or U9274 (N_9274,N_9126,N_9111);
nand U9275 (N_9275,N_9205,N_9192);
xnor U9276 (N_9276,N_9045,N_9013);
nor U9277 (N_9277,N_9215,N_9073);
xor U9278 (N_9278,N_9199,N_9120);
xnor U9279 (N_9279,N_9075,N_9146);
and U9280 (N_9280,N_9187,N_9246);
xnor U9281 (N_9281,N_9201,N_9134);
nand U9282 (N_9282,N_9158,N_9237);
or U9283 (N_9283,N_9004,N_9179);
nand U9284 (N_9284,N_9171,N_9176);
nand U9285 (N_9285,N_9059,N_9113);
or U9286 (N_9286,N_9162,N_9066);
and U9287 (N_9287,N_9048,N_9043);
nand U9288 (N_9288,N_9245,N_9032);
nand U9289 (N_9289,N_9050,N_9216);
nand U9290 (N_9290,N_9055,N_9249);
xnor U9291 (N_9291,N_9218,N_9226);
or U9292 (N_9292,N_9223,N_9125);
nor U9293 (N_9293,N_9077,N_9083);
or U9294 (N_9294,N_9003,N_9014);
nand U9295 (N_9295,N_9044,N_9235);
and U9296 (N_9296,N_9116,N_9035);
nor U9297 (N_9297,N_9000,N_9011);
xor U9298 (N_9298,N_9033,N_9229);
xor U9299 (N_9299,N_9129,N_9166);
and U9300 (N_9300,N_9060,N_9057);
or U9301 (N_9301,N_9047,N_9085);
nor U9302 (N_9302,N_9090,N_9163);
or U9303 (N_9303,N_9024,N_9149);
or U9304 (N_9304,N_9012,N_9236);
or U9305 (N_9305,N_9069,N_9206);
nor U9306 (N_9306,N_9182,N_9139);
or U9307 (N_9307,N_9061,N_9122);
and U9308 (N_9308,N_9217,N_9207);
and U9309 (N_9309,N_9194,N_9091);
and U9310 (N_9310,N_9037,N_9184);
or U9311 (N_9311,N_9185,N_9150);
or U9312 (N_9312,N_9128,N_9102);
nand U9313 (N_9313,N_9046,N_9030);
nand U9314 (N_9314,N_9097,N_9228);
or U9315 (N_9315,N_9240,N_9183);
or U9316 (N_9316,N_9203,N_9100);
xnor U9317 (N_9317,N_9036,N_9178);
or U9318 (N_9318,N_9161,N_9168);
xor U9319 (N_9319,N_9210,N_9088);
xnor U9320 (N_9320,N_9123,N_9200);
or U9321 (N_9321,N_9145,N_9159);
nand U9322 (N_9322,N_9092,N_9148);
or U9323 (N_9323,N_9174,N_9191);
and U9324 (N_9324,N_9029,N_9114);
xnor U9325 (N_9325,N_9181,N_9127);
xor U9326 (N_9326,N_9005,N_9137);
xor U9327 (N_9327,N_9170,N_9156);
nor U9328 (N_9328,N_9202,N_9115);
or U9329 (N_9329,N_9016,N_9062);
xor U9330 (N_9330,N_9112,N_9051);
or U9331 (N_9331,N_9106,N_9058);
or U9332 (N_9332,N_9130,N_9118);
and U9333 (N_9333,N_9186,N_9109);
xnor U9334 (N_9334,N_9234,N_9195);
or U9335 (N_9335,N_9103,N_9067);
or U9336 (N_9336,N_9071,N_9028);
xor U9337 (N_9337,N_9089,N_9086);
xor U9338 (N_9338,N_9027,N_9098);
nand U9339 (N_9339,N_9173,N_9151);
and U9340 (N_9340,N_9241,N_9104);
or U9341 (N_9341,N_9222,N_9141);
or U9342 (N_9342,N_9002,N_9230);
nor U9343 (N_9343,N_9239,N_9209);
or U9344 (N_9344,N_9052,N_9096);
and U9345 (N_9345,N_9157,N_9177);
and U9346 (N_9346,N_9056,N_9042);
or U9347 (N_9347,N_9087,N_9143);
nor U9348 (N_9348,N_9196,N_9107);
nand U9349 (N_9349,N_9068,N_9212);
xor U9350 (N_9350,N_9076,N_9065);
or U9351 (N_9351,N_9039,N_9227);
nor U9352 (N_9352,N_9220,N_9133);
and U9353 (N_9353,N_9082,N_9072);
nand U9354 (N_9354,N_9101,N_9242);
and U9355 (N_9355,N_9138,N_9208);
xor U9356 (N_9356,N_9232,N_9169);
and U9357 (N_9357,N_9017,N_9131);
nand U9358 (N_9358,N_9140,N_9021);
nand U9359 (N_9359,N_9007,N_9180);
and U9360 (N_9360,N_9054,N_9198);
nand U9361 (N_9361,N_9117,N_9074);
nor U9362 (N_9362,N_9135,N_9144);
xnor U9363 (N_9363,N_9244,N_9219);
nor U9364 (N_9364,N_9243,N_9108);
nor U9365 (N_9365,N_9053,N_9142);
or U9366 (N_9366,N_9001,N_9231);
and U9367 (N_9367,N_9084,N_9248);
nor U9368 (N_9368,N_9022,N_9152);
nand U9369 (N_9369,N_9197,N_9009);
or U9370 (N_9370,N_9193,N_9224);
nor U9371 (N_9371,N_9167,N_9160);
nand U9372 (N_9372,N_9078,N_9081);
xor U9373 (N_9373,N_9040,N_9049);
or U9374 (N_9374,N_9154,N_9190);
nand U9375 (N_9375,N_9238,N_9169);
and U9376 (N_9376,N_9117,N_9060);
nor U9377 (N_9377,N_9190,N_9096);
nor U9378 (N_9378,N_9027,N_9109);
nand U9379 (N_9379,N_9036,N_9058);
xnor U9380 (N_9380,N_9017,N_9105);
xnor U9381 (N_9381,N_9117,N_9189);
or U9382 (N_9382,N_9118,N_9233);
and U9383 (N_9383,N_9184,N_9136);
nand U9384 (N_9384,N_9220,N_9014);
nor U9385 (N_9385,N_9083,N_9185);
and U9386 (N_9386,N_9113,N_9022);
and U9387 (N_9387,N_9223,N_9023);
and U9388 (N_9388,N_9004,N_9111);
or U9389 (N_9389,N_9051,N_9005);
and U9390 (N_9390,N_9181,N_9165);
xnor U9391 (N_9391,N_9149,N_9060);
and U9392 (N_9392,N_9238,N_9214);
and U9393 (N_9393,N_9031,N_9093);
and U9394 (N_9394,N_9126,N_9206);
nand U9395 (N_9395,N_9114,N_9221);
nor U9396 (N_9396,N_9117,N_9124);
nor U9397 (N_9397,N_9035,N_9102);
and U9398 (N_9398,N_9146,N_9098);
xnor U9399 (N_9399,N_9199,N_9031);
nor U9400 (N_9400,N_9053,N_9044);
and U9401 (N_9401,N_9012,N_9107);
xnor U9402 (N_9402,N_9141,N_9031);
xnor U9403 (N_9403,N_9087,N_9148);
nor U9404 (N_9404,N_9100,N_9058);
xnor U9405 (N_9405,N_9025,N_9208);
nand U9406 (N_9406,N_9215,N_9138);
or U9407 (N_9407,N_9175,N_9229);
or U9408 (N_9408,N_9231,N_9089);
nand U9409 (N_9409,N_9114,N_9064);
nand U9410 (N_9410,N_9194,N_9064);
and U9411 (N_9411,N_9086,N_9128);
nor U9412 (N_9412,N_9169,N_9130);
and U9413 (N_9413,N_9246,N_9079);
nand U9414 (N_9414,N_9227,N_9208);
or U9415 (N_9415,N_9012,N_9116);
or U9416 (N_9416,N_9158,N_9200);
nand U9417 (N_9417,N_9033,N_9234);
xnor U9418 (N_9418,N_9142,N_9159);
nand U9419 (N_9419,N_9158,N_9037);
nand U9420 (N_9420,N_9019,N_9107);
nor U9421 (N_9421,N_9193,N_9019);
nor U9422 (N_9422,N_9163,N_9141);
nor U9423 (N_9423,N_9101,N_9096);
nand U9424 (N_9424,N_9163,N_9240);
and U9425 (N_9425,N_9198,N_9104);
nand U9426 (N_9426,N_9247,N_9148);
or U9427 (N_9427,N_9004,N_9236);
xor U9428 (N_9428,N_9220,N_9020);
and U9429 (N_9429,N_9132,N_9112);
or U9430 (N_9430,N_9202,N_9054);
nor U9431 (N_9431,N_9020,N_9215);
xnor U9432 (N_9432,N_9009,N_9123);
nor U9433 (N_9433,N_9099,N_9171);
or U9434 (N_9434,N_9035,N_9111);
nor U9435 (N_9435,N_9195,N_9085);
and U9436 (N_9436,N_9001,N_9188);
xnor U9437 (N_9437,N_9236,N_9100);
nor U9438 (N_9438,N_9041,N_9074);
nand U9439 (N_9439,N_9068,N_9214);
nor U9440 (N_9440,N_9241,N_9050);
and U9441 (N_9441,N_9160,N_9125);
nor U9442 (N_9442,N_9158,N_9018);
and U9443 (N_9443,N_9091,N_9241);
nand U9444 (N_9444,N_9053,N_9234);
or U9445 (N_9445,N_9184,N_9096);
or U9446 (N_9446,N_9235,N_9241);
nand U9447 (N_9447,N_9164,N_9228);
and U9448 (N_9448,N_9218,N_9081);
nand U9449 (N_9449,N_9137,N_9105);
or U9450 (N_9450,N_9093,N_9155);
nor U9451 (N_9451,N_9248,N_9108);
or U9452 (N_9452,N_9202,N_9111);
or U9453 (N_9453,N_9145,N_9059);
nand U9454 (N_9454,N_9207,N_9209);
nand U9455 (N_9455,N_9078,N_9189);
nand U9456 (N_9456,N_9219,N_9120);
and U9457 (N_9457,N_9107,N_9061);
or U9458 (N_9458,N_9116,N_9222);
xor U9459 (N_9459,N_9170,N_9168);
nor U9460 (N_9460,N_9116,N_9061);
nor U9461 (N_9461,N_9235,N_9110);
nand U9462 (N_9462,N_9104,N_9153);
or U9463 (N_9463,N_9137,N_9169);
xnor U9464 (N_9464,N_9076,N_9120);
and U9465 (N_9465,N_9122,N_9115);
nor U9466 (N_9466,N_9031,N_9046);
and U9467 (N_9467,N_9192,N_9035);
nand U9468 (N_9468,N_9051,N_9135);
or U9469 (N_9469,N_9233,N_9031);
and U9470 (N_9470,N_9126,N_9051);
xnor U9471 (N_9471,N_9228,N_9172);
nor U9472 (N_9472,N_9216,N_9113);
nor U9473 (N_9473,N_9221,N_9204);
nand U9474 (N_9474,N_9241,N_9229);
and U9475 (N_9475,N_9016,N_9054);
xnor U9476 (N_9476,N_9072,N_9021);
or U9477 (N_9477,N_9149,N_9240);
xnor U9478 (N_9478,N_9215,N_9063);
nand U9479 (N_9479,N_9049,N_9157);
and U9480 (N_9480,N_9196,N_9235);
or U9481 (N_9481,N_9022,N_9079);
nor U9482 (N_9482,N_9155,N_9235);
and U9483 (N_9483,N_9125,N_9070);
xor U9484 (N_9484,N_9060,N_9183);
xnor U9485 (N_9485,N_9015,N_9194);
and U9486 (N_9486,N_9032,N_9063);
nor U9487 (N_9487,N_9134,N_9130);
or U9488 (N_9488,N_9189,N_9041);
or U9489 (N_9489,N_9075,N_9190);
and U9490 (N_9490,N_9236,N_9018);
nand U9491 (N_9491,N_9173,N_9165);
or U9492 (N_9492,N_9242,N_9000);
nor U9493 (N_9493,N_9186,N_9054);
and U9494 (N_9494,N_9194,N_9144);
or U9495 (N_9495,N_9065,N_9224);
nand U9496 (N_9496,N_9034,N_9006);
xnor U9497 (N_9497,N_9212,N_9046);
or U9498 (N_9498,N_9206,N_9211);
and U9499 (N_9499,N_9172,N_9049);
nand U9500 (N_9500,N_9300,N_9366);
nand U9501 (N_9501,N_9363,N_9308);
nand U9502 (N_9502,N_9496,N_9413);
xnor U9503 (N_9503,N_9442,N_9254);
nand U9504 (N_9504,N_9423,N_9417);
nor U9505 (N_9505,N_9447,N_9252);
and U9506 (N_9506,N_9327,N_9260);
xnor U9507 (N_9507,N_9481,N_9486);
xor U9508 (N_9508,N_9351,N_9272);
and U9509 (N_9509,N_9398,N_9455);
xnor U9510 (N_9510,N_9492,N_9409);
nand U9511 (N_9511,N_9378,N_9335);
and U9512 (N_9512,N_9290,N_9281);
nor U9513 (N_9513,N_9433,N_9493);
or U9514 (N_9514,N_9499,N_9436);
xor U9515 (N_9515,N_9410,N_9372);
and U9516 (N_9516,N_9253,N_9497);
xnor U9517 (N_9517,N_9469,N_9344);
nand U9518 (N_9518,N_9263,N_9371);
and U9519 (N_9519,N_9353,N_9307);
and U9520 (N_9520,N_9444,N_9289);
or U9521 (N_9521,N_9419,N_9412);
or U9522 (N_9522,N_9386,N_9389);
and U9523 (N_9523,N_9293,N_9275);
nand U9524 (N_9524,N_9399,N_9451);
and U9525 (N_9525,N_9375,N_9473);
nor U9526 (N_9526,N_9323,N_9251);
nand U9527 (N_9527,N_9302,N_9402);
or U9528 (N_9528,N_9355,N_9431);
or U9529 (N_9529,N_9397,N_9296);
or U9530 (N_9530,N_9277,N_9405);
or U9531 (N_9531,N_9332,N_9333);
xnor U9532 (N_9532,N_9458,N_9374);
nor U9533 (N_9533,N_9257,N_9314);
nand U9534 (N_9534,N_9471,N_9325);
nand U9535 (N_9535,N_9264,N_9286);
nor U9536 (N_9536,N_9396,N_9424);
xor U9537 (N_9537,N_9420,N_9352);
or U9538 (N_9538,N_9370,N_9348);
or U9539 (N_9539,N_9256,N_9491);
nor U9540 (N_9540,N_9324,N_9316);
or U9541 (N_9541,N_9421,N_9448);
nor U9542 (N_9542,N_9360,N_9288);
and U9543 (N_9543,N_9416,N_9401);
or U9544 (N_9544,N_9285,N_9346);
nor U9545 (N_9545,N_9490,N_9443);
or U9546 (N_9546,N_9259,N_9428);
or U9547 (N_9547,N_9376,N_9310);
nor U9548 (N_9548,N_9270,N_9488);
xor U9549 (N_9549,N_9474,N_9303);
nand U9550 (N_9550,N_9341,N_9321);
and U9551 (N_9551,N_9317,N_9391);
or U9552 (N_9552,N_9468,N_9425);
or U9553 (N_9553,N_9439,N_9337);
xnor U9554 (N_9554,N_9465,N_9380);
xor U9555 (N_9555,N_9438,N_9477);
nand U9556 (N_9556,N_9326,N_9279);
and U9557 (N_9557,N_9268,N_9261);
and U9558 (N_9558,N_9364,N_9322);
or U9559 (N_9559,N_9462,N_9475);
or U9560 (N_9560,N_9358,N_9388);
nor U9561 (N_9561,N_9385,N_9450);
nand U9562 (N_9562,N_9422,N_9482);
xnor U9563 (N_9563,N_9362,N_9258);
or U9564 (N_9564,N_9373,N_9298);
or U9565 (N_9565,N_9449,N_9336);
nand U9566 (N_9566,N_9356,N_9459);
and U9567 (N_9567,N_9415,N_9487);
or U9568 (N_9568,N_9379,N_9434);
or U9569 (N_9569,N_9483,N_9287);
or U9570 (N_9570,N_9390,N_9480);
or U9571 (N_9571,N_9394,N_9343);
or U9572 (N_9572,N_9342,N_9274);
and U9573 (N_9573,N_9411,N_9456);
and U9574 (N_9574,N_9466,N_9400);
nor U9575 (N_9575,N_9276,N_9311);
nor U9576 (N_9576,N_9478,N_9291);
nand U9577 (N_9577,N_9345,N_9349);
xnor U9578 (N_9578,N_9320,N_9347);
and U9579 (N_9579,N_9467,N_9359);
xor U9580 (N_9580,N_9318,N_9452);
xnor U9581 (N_9581,N_9494,N_9304);
and U9582 (N_9582,N_9445,N_9418);
and U9583 (N_9583,N_9334,N_9384);
xnor U9584 (N_9584,N_9407,N_9269);
nand U9585 (N_9585,N_9457,N_9387);
nand U9586 (N_9586,N_9377,N_9495);
or U9587 (N_9587,N_9454,N_9406);
nand U9588 (N_9588,N_9295,N_9265);
nand U9589 (N_9589,N_9313,N_9381);
and U9590 (N_9590,N_9441,N_9404);
and U9591 (N_9591,N_9292,N_9393);
nor U9592 (N_9592,N_9382,N_9403);
and U9593 (N_9593,N_9392,N_9299);
xor U9594 (N_9594,N_9470,N_9453);
nor U9595 (N_9595,N_9461,N_9479);
nor U9596 (N_9596,N_9432,N_9330);
nand U9597 (N_9597,N_9312,N_9340);
xnor U9598 (N_9598,N_9369,N_9331);
nand U9599 (N_9599,N_9301,N_9485);
and U9600 (N_9600,N_9368,N_9294);
xnor U9601 (N_9601,N_9354,N_9271);
xor U9602 (N_9602,N_9267,N_9437);
xnor U9603 (N_9603,N_9361,N_9339);
and U9604 (N_9604,N_9319,N_9273);
nand U9605 (N_9605,N_9315,N_9357);
or U9606 (N_9606,N_9305,N_9463);
or U9607 (N_9607,N_9435,N_9338);
xnor U9608 (N_9608,N_9309,N_9498);
nor U9609 (N_9609,N_9440,N_9255);
nor U9610 (N_9610,N_9262,N_9328);
nand U9611 (N_9611,N_9365,N_9278);
or U9612 (N_9612,N_9284,N_9427);
nand U9613 (N_9613,N_9429,N_9489);
xnor U9614 (N_9614,N_9250,N_9476);
and U9615 (N_9615,N_9266,N_9297);
xnor U9616 (N_9616,N_9350,N_9408);
nand U9617 (N_9617,N_9464,N_9460);
xnor U9618 (N_9618,N_9283,N_9414);
xnor U9619 (N_9619,N_9472,N_9426);
or U9620 (N_9620,N_9484,N_9280);
xnor U9621 (N_9621,N_9367,N_9395);
or U9622 (N_9622,N_9329,N_9383);
and U9623 (N_9623,N_9282,N_9430);
nor U9624 (N_9624,N_9306,N_9446);
xor U9625 (N_9625,N_9303,N_9390);
nand U9626 (N_9626,N_9397,N_9436);
nand U9627 (N_9627,N_9284,N_9250);
and U9628 (N_9628,N_9334,N_9443);
or U9629 (N_9629,N_9290,N_9474);
nor U9630 (N_9630,N_9467,N_9392);
nand U9631 (N_9631,N_9454,N_9363);
or U9632 (N_9632,N_9381,N_9296);
and U9633 (N_9633,N_9387,N_9393);
xor U9634 (N_9634,N_9262,N_9380);
xnor U9635 (N_9635,N_9461,N_9430);
nor U9636 (N_9636,N_9333,N_9365);
or U9637 (N_9637,N_9466,N_9388);
and U9638 (N_9638,N_9403,N_9295);
and U9639 (N_9639,N_9480,N_9397);
and U9640 (N_9640,N_9491,N_9328);
xnor U9641 (N_9641,N_9434,N_9479);
or U9642 (N_9642,N_9257,N_9311);
or U9643 (N_9643,N_9276,N_9454);
nor U9644 (N_9644,N_9264,N_9381);
xor U9645 (N_9645,N_9291,N_9429);
and U9646 (N_9646,N_9446,N_9385);
and U9647 (N_9647,N_9443,N_9398);
or U9648 (N_9648,N_9283,N_9318);
nor U9649 (N_9649,N_9383,N_9259);
nor U9650 (N_9650,N_9336,N_9315);
nor U9651 (N_9651,N_9385,N_9331);
and U9652 (N_9652,N_9305,N_9293);
and U9653 (N_9653,N_9326,N_9358);
and U9654 (N_9654,N_9355,N_9489);
and U9655 (N_9655,N_9432,N_9435);
and U9656 (N_9656,N_9411,N_9301);
or U9657 (N_9657,N_9335,N_9384);
nor U9658 (N_9658,N_9337,N_9252);
nor U9659 (N_9659,N_9349,N_9457);
or U9660 (N_9660,N_9262,N_9263);
nand U9661 (N_9661,N_9460,N_9429);
nor U9662 (N_9662,N_9281,N_9363);
and U9663 (N_9663,N_9389,N_9489);
nor U9664 (N_9664,N_9381,N_9462);
and U9665 (N_9665,N_9442,N_9466);
nor U9666 (N_9666,N_9484,N_9264);
or U9667 (N_9667,N_9483,N_9351);
xnor U9668 (N_9668,N_9285,N_9428);
nor U9669 (N_9669,N_9264,N_9363);
nor U9670 (N_9670,N_9359,N_9423);
and U9671 (N_9671,N_9280,N_9409);
xnor U9672 (N_9672,N_9364,N_9332);
xor U9673 (N_9673,N_9274,N_9400);
xor U9674 (N_9674,N_9321,N_9389);
xnor U9675 (N_9675,N_9388,N_9438);
or U9676 (N_9676,N_9413,N_9268);
nand U9677 (N_9677,N_9420,N_9438);
xor U9678 (N_9678,N_9375,N_9451);
nor U9679 (N_9679,N_9342,N_9415);
xnor U9680 (N_9680,N_9392,N_9321);
or U9681 (N_9681,N_9259,N_9374);
nor U9682 (N_9682,N_9256,N_9359);
xnor U9683 (N_9683,N_9471,N_9351);
nand U9684 (N_9684,N_9316,N_9347);
nor U9685 (N_9685,N_9364,N_9321);
or U9686 (N_9686,N_9334,N_9476);
xor U9687 (N_9687,N_9426,N_9389);
xor U9688 (N_9688,N_9408,N_9351);
nand U9689 (N_9689,N_9447,N_9317);
nor U9690 (N_9690,N_9273,N_9316);
nand U9691 (N_9691,N_9359,N_9300);
xnor U9692 (N_9692,N_9424,N_9287);
and U9693 (N_9693,N_9461,N_9473);
nand U9694 (N_9694,N_9323,N_9475);
xnor U9695 (N_9695,N_9447,N_9313);
nor U9696 (N_9696,N_9438,N_9269);
and U9697 (N_9697,N_9250,N_9307);
and U9698 (N_9698,N_9322,N_9313);
nor U9699 (N_9699,N_9434,N_9375);
and U9700 (N_9700,N_9271,N_9435);
nand U9701 (N_9701,N_9476,N_9446);
nand U9702 (N_9702,N_9412,N_9444);
nor U9703 (N_9703,N_9406,N_9346);
nor U9704 (N_9704,N_9278,N_9416);
nand U9705 (N_9705,N_9311,N_9499);
and U9706 (N_9706,N_9383,N_9478);
nor U9707 (N_9707,N_9389,N_9259);
nand U9708 (N_9708,N_9294,N_9466);
or U9709 (N_9709,N_9269,N_9393);
and U9710 (N_9710,N_9263,N_9493);
or U9711 (N_9711,N_9354,N_9478);
or U9712 (N_9712,N_9333,N_9347);
nor U9713 (N_9713,N_9401,N_9290);
or U9714 (N_9714,N_9410,N_9440);
xor U9715 (N_9715,N_9413,N_9380);
nor U9716 (N_9716,N_9404,N_9250);
nand U9717 (N_9717,N_9314,N_9482);
nand U9718 (N_9718,N_9439,N_9412);
xor U9719 (N_9719,N_9417,N_9478);
xnor U9720 (N_9720,N_9370,N_9432);
nor U9721 (N_9721,N_9433,N_9494);
xnor U9722 (N_9722,N_9393,N_9284);
nor U9723 (N_9723,N_9450,N_9400);
or U9724 (N_9724,N_9282,N_9478);
and U9725 (N_9725,N_9354,N_9339);
and U9726 (N_9726,N_9385,N_9427);
xor U9727 (N_9727,N_9350,N_9422);
and U9728 (N_9728,N_9369,N_9480);
or U9729 (N_9729,N_9338,N_9411);
xor U9730 (N_9730,N_9494,N_9372);
xnor U9731 (N_9731,N_9270,N_9321);
and U9732 (N_9732,N_9355,N_9357);
nand U9733 (N_9733,N_9334,N_9296);
and U9734 (N_9734,N_9495,N_9438);
nor U9735 (N_9735,N_9391,N_9284);
nand U9736 (N_9736,N_9314,N_9372);
nand U9737 (N_9737,N_9316,N_9496);
nor U9738 (N_9738,N_9262,N_9294);
nand U9739 (N_9739,N_9383,N_9378);
nor U9740 (N_9740,N_9433,N_9294);
xor U9741 (N_9741,N_9263,N_9480);
nor U9742 (N_9742,N_9489,N_9312);
nand U9743 (N_9743,N_9419,N_9379);
and U9744 (N_9744,N_9440,N_9267);
or U9745 (N_9745,N_9489,N_9448);
nor U9746 (N_9746,N_9409,N_9294);
or U9747 (N_9747,N_9420,N_9493);
xor U9748 (N_9748,N_9300,N_9420);
nand U9749 (N_9749,N_9322,N_9395);
and U9750 (N_9750,N_9601,N_9544);
nand U9751 (N_9751,N_9632,N_9541);
or U9752 (N_9752,N_9697,N_9642);
xnor U9753 (N_9753,N_9617,N_9560);
and U9754 (N_9754,N_9629,N_9516);
and U9755 (N_9755,N_9711,N_9509);
xnor U9756 (N_9756,N_9550,N_9539);
xor U9757 (N_9757,N_9698,N_9596);
and U9758 (N_9758,N_9715,N_9625);
nand U9759 (N_9759,N_9546,N_9590);
nor U9760 (N_9760,N_9524,N_9639);
nor U9761 (N_9761,N_9643,N_9635);
or U9762 (N_9762,N_9520,N_9681);
and U9763 (N_9763,N_9615,N_9621);
nor U9764 (N_9764,N_9679,N_9511);
or U9765 (N_9765,N_9559,N_9626);
and U9766 (N_9766,N_9510,N_9659);
or U9767 (N_9767,N_9543,N_9609);
and U9768 (N_9768,N_9567,N_9529);
nor U9769 (N_9769,N_9630,N_9731);
and U9770 (N_9770,N_9628,N_9655);
nand U9771 (N_9771,N_9651,N_9605);
and U9772 (N_9772,N_9582,N_9707);
nand U9773 (N_9773,N_9547,N_9537);
and U9774 (N_9774,N_9568,N_9523);
or U9775 (N_9775,N_9746,N_9744);
nand U9776 (N_9776,N_9552,N_9737);
nand U9777 (N_9777,N_9576,N_9636);
nand U9778 (N_9778,N_9500,N_9563);
or U9779 (N_9779,N_9591,N_9647);
and U9780 (N_9780,N_9745,N_9555);
xor U9781 (N_9781,N_9666,N_9665);
nor U9782 (N_9782,N_9506,N_9536);
or U9783 (N_9783,N_9699,N_9686);
nor U9784 (N_9784,N_9689,N_9557);
xor U9785 (N_9785,N_9504,N_9574);
and U9786 (N_9786,N_9706,N_9503);
or U9787 (N_9787,N_9719,N_9712);
and U9788 (N_9788,N_9589,N_9627);
or U9789 (N_9789,N_9723,N_9733);
nand U9790 (N_9790,N_9739,N_9556);
nor U9791 (N_9791,N_9508,N_9736);
xor U9792 (N_9792,N_9695,N_9728);
nor U9793 (N_9793,N_9549,N_9595);
xnor U9794 (N_9794,N_9606,N_9604);
nor U9795 (N_9795,N_9741,N_9518);
xor U9796 (N_9796,N_9545,N_9717);
nand U9797 (N_9797,N_9684,N_9577);
and U9798 (N_9798,N_9661,N_9743);
nor U9799 (N_9799,N_9502,N_9522);
nand U9800 (N_9800,N_9533,N_9517);
nor U9801 (N_9801,N_9685,N_9648);
xor U9802 (N_9802,N_9564,N_9730);
and U9803 (N_9803,N_9571,N_9521);
or U9804 (N_9804,N_9603,N_9548);
and U9805 (N_9805,N_9578,N_9593);
and U9806 (N_9806,N_9586,N_9507);
nor U9807 (N_9807,N_9670,N_9663);
xor U9808 (N_9808,N_9569,N_9703);
nor U9809 (N_9809,N_9718,N_9727);
and U9810 (N_9810,N_9734,N_9722);
or U9811 (N_9811,N_9662,N_9608);
xnor U9812 (N_9812,N_9677,N_9542);
xnor U9813 (N_9813,N_9638,N_9554);
xnor U9814 (N_9814,N_9641,N_9614);
and U9815 (N_9815,N_9724,N_9602);
xnor U9816 (N_9816,N_9505,N_9624);
and U9817 (N_9817,N_9740,N_9579);
nor U9818 (N_9818,N_9599,N_9742);
nand U9819 (N_9819,N_9683,N_9652);
nor U9820 (N_9820,N_9696,N_9725);
or U9821 (N_9821,N_9610,N_9738);
nor U9822 (N_9822,N_9688,N_9553);
nand U9823 (N_9823,N_9583,N_9588);
nor U9824 (N_9824,N_9747,N_9716);
and U9825 (N_9825,N_9534,N_9540);
xor U9826 (N_9826,N_9708,N_9721);
and U9827 (N_9827,N_9748,N_9620);
nand U9828 (N_9828,N_9607,N_9519);
or U9829 (N_9829,N_9700,N_9565);
nand U9830 (N_9830,N_9640,N_9678);
nand U9831 (N_9831,N_9575,N_9616);
nor U9832 (N_9832,N_9501,N_9594);
nand U9833 (N_9833,N_9581,N_9649);
xnor U9834 (N_9834,N_9633,N_9551);
and U9835 (N_9835,N_9644,N_9668);
nand U9836 (N_9836,N_9514,N_9680);
and U9837 (N_9837,N_9654,N_9623);
nand U9838 (N_9838,N_9713,N_9729);
xor U9839 (N_9839,N_9515,N_9611);
nor U9840 (N_9840,N_9597,N_9527);
and U9841 (N_9841,N_9704,N_9584);
or U9842 (N_9842,N_9732,N_9587);
nor U9843 (N_9843,N_9573,N_9671);
or U9844 (N_9844,N_9709,N_9580);
or U9845 (N_9845,N_9714,N_9622);
or U9846 (N_9846,N_9674,N_9562);
or U9847 (N_9847,N_9600,N_9528);
or U9848 (N_9848,N_9676,N_9613);
or U9849 (N_9849,N_9705,N_9702);
xor U9850 (N_9850,N_9653,N_9512);
or U9851 (N_9851,N_9561,N_9720);
nor U9852 (N_9852,N_9592,N_9657);
or U9853 (N_9853,N_9735,N_9646);
and U9854 (N_9854,N_9694,N_9691);
and U9855 (N_9855,N_9585,N_9532);
and U9856 (N_9856,N_9667,N_9669);
and U9857 (N_9857,N_9538,N_9634);
xor U9858 (N_9858,N_9618,N_9650);
nand U9859 (N_9859,N_9558,N_9726);
nor U9860 (N_9860,N_9749,N_9526);
nor U9861 (N_9861,N_9692,N_9598);
or U9862 (N_9862,N_9572,N_9612);
xnor U9863 (N_9863,N_9690,N_9660);
and U9864 (N_9864,N_9535,N_9710);
nand U9865 (N_9865,N_9525,N_9656);
and U9866 (N_9866,N_9513,N_9664);
or U9867 (N_9867,N_9619,N_9693);
and U9868 (N_9868,N_9531,N_9530);
or U9869 (N_9869,N_9637,N_9701);
nor U9870 (N_9870,N_9645,N_9570);
xor U9871 (N_9871,N_9682,N_9672);
and U9872 (N_9872,N_9675,N_9658);
nand U9873 (N_9873,N_9631,N_9566);
or U9874 (N_9874,N_9673,N_9687);
and U9875 (N_9875,N_9605,N_9719);
nor U9876 (N_9876,N_9596,N_9530);
nor U9877 (N_9877,N_9577,N_9606);
or U9878 (N_9878,N_9536,N_9552);
nand U9879 (N_9879,N_9680,N_9709);
xnor U9880 (N_9880,N_9681,N_9567);
or U9881 (N_9881,N_9694,N_9581);
or U9882 (N_9882,N_9515,N_9667);
xnor U9883 (N_9883,N_9652,N_9669);
and U9884 (N_9884,N_9604,N_9631);
xnor U9885 (N_9885,N_9598,N_9550);
xor U9886 (N_9886,N_9639,N_9718);
or U9887 (N_9887,N_9707,N_9535);
nand U9888 (N_9888,N_9737,N_9668);
xor U9889 (N_9889,N_9580,N_9740);
xor U9890 (N_9890,N_9650,N_9676);
and U9891 (N_9891,N_9561,N_9731);
or U9892 (N_9892,N_9539,N_9730);
xor U9893 (N_9893,N_9577,N_9647);
nand U9894 (N_9894,N_9646,N_9529);
and U9895 (N_9895,N_9549,N_9639);
nor U9896 (N_9896,N_9610,N_9524);
xnor U9897 (N_9897,N_9609,N_9501);
or U9898 (N_9898,N_9522,N_9566);
or U9899 (N_9899,N_9602,N_9720);
nand U9900 (N_9900,N_9708,N_9571);
and U9901 (N_9901,N_9593,N_9596);
xor U9902 (N_9902,N_9675,N_9690);
nor U9903 (N_9903,N_9562,N_9654);
nand U9904 (N_9904,N_9663,N_9557);
nor U9905 (N_9905,N_9586,N_9644);
nor U9906 (N_9906,N_9616,N_9647);
or U9907 (N_9907,N_9734,N_9549);
nand U9908 (N_9908,N_9739,N_9684);
or U9909 (N_9909,N_9655,N_9684);
xor U9910 (N_9910,N_9570,N_9678);
nand U9911 (N_9911,N_9697,N_9539);
and U9912 (N_9912,N_9608,N_9530);
nand U9913 (N_9913,N_9516,N_9709);
or U9914 (N_9914,N_9743,N_9540);
xnor U9915 (N_9915,N_9704,N_9598);
and U9916 (N_9916,N_9542,N_9693);
xnor U9917 (N_9917,N_9514,N_9740);
and U9918 (N_9918,N_9531,N_9535);
nand U9919 (N_9919,N_9530,N_9545);
xnor U9920 (N_9920,N_9662,N_9637);
nor U9921 (N_9921,N_9667,N_9549);
nor U9922 (N_9922,N_9514,N_9722);
and U9923 (N_9923,N_9729,N_9543);
nor U9924 (N_9924,N_9581,N_9562);
nand U9925 (N_9925,N_9664,N_9503);
or U9926 (N_9926,N_9503,N_9538);
xor U9927 (N_9927,N_9577,N_9505);
xor U9928 (N_9928,N_9507,N_9749);
nor U9929 (N_9929,N_9729,N_9657);
nor U9930 (N_9930,N_9669,N_9512);
or U9931 (N_9931,N_9746,N_9570);
nor U9932 (N_9932,N_9679,N_9594);
and U9933 (N_9933,N_9548,N_9567);
or U9934 (N_9934,N_9645,N_9739);
xnor U9935 (N_9935,N_9747,N_9656);
xnor U9936 (N_9936,N_9741,N_9662);
xnor U9937 (N_9937,N_9634,N_9622);
or U9938 (N_9938,N_9649,N_9742);
nand U9939 (N_9939,N_9718,N_9690);
xor U9940 (N_9940,N_9533,N_9519);
or U9941 (N_9941,N_9534,N_9694);
nor U9942 (N_9942,N_9541,N_9621);
and U9943 (N_9943,N_9597,N_9708);
xor U9944 (N_9944,N_9647,N_9501);
xnor U9945 (N_9945,N_9609,N_9716);
xnor U9946 (N_9946,N_9610,N_9586);
and U9947 (N_9947,N_9733,N_9594);
nor U9948 (N_9948,N_9732,N_9593);
and U9949 (N_9949,N_9567,N_9596);
xor U9950 (N_9950,N_9517,N_9644);
and U9951 (N_9951,N_9555,N_9535);
or U9952 (N_9952,N_9503,N_9671);
xnor U9953 (N_9953,N_9705,N_9725);
and U9954 (N_9954,N_9551,N_9593);
nand U9955 (N_9955,N_9600,N_9568);
and U9956 (N_9956,N_9671,N_9579);
nor U9957 (N_9957,N_9592,N_9501);
xor U9958 (N_9958,N_9511,N_9593);
or U9959 (N_9959,N_9569,N_9613);
xor U9960 (N_9960,N_9695,N_9552);
or U9961 (N_9961,N_9567,N_9726);
and U9962 (N_9962,N_9634,N_9568);
and U9963 (N_9963,N_9607,N_9643);
and U9964 (N_9964,N_9746,N_9612);
or U9965 (N_9965,N_9547,N_9536);
nand U9966 (N_9966,N_9557,N_9573);
xnor U9967 (N_9967,N_9606,N_9529);
nand U9968 (N_9968,N_9697,N_9637);
nand U9969 (N_9969,N_9593,N_9641);
and U9970 (N_9970,N_9744,N_9745);
nand U9971 (N_9971,N_9744,N_9542);
nor U9972 (N_9972,N_9538,N_9730);
or U9973 (N_9973,N_9634,N_9723);
or U9974 (N_9974,N_9636,N_9710);
and U9975 (N_9975,N_9615,N_9515);
xor U9976 (N_9976,N_9698,N_9690);
or U9977 (N_9977,N_9720,N_9663);
and U9978 (N_9978,N_9602,N_9570);
nor U9979 (N_9979,N_9620,N_9547);
xnor U9980 (N_9980,N_9523,N_9505);
xor U9981 (N_9981,N_9622,N_9673);
xor U9982 (N_9982,N_9516,N_9607);
or U9983 (N_9983,N_9617,N_9562);
xnor U9984 (N_9984,N_9597,N_9749);
nor U9985 (N_9985,N_9681,N_9713);
nand U9986 (N_9986,N_9569,N_9713);
nor U9987 (N_9987,N_9729,N_9578);
or U9988 (N_9988,N_9510,N_9503);
nand U9989 (N_9989,N_9515,N_9725);
nand U9990 (N_9990,N_9730,N_9685);
xor U9991 (N_9991,N_9633,N_9500);
xor U9992 (N_9992,N_9560,N_9588);
or U9993 (N_9993,N_9713,N_9603);
xnor U9994 (N_9994,N_9717,N_9571);
nand U9995 (N_9995,N_9601,N_9564);
nand U9996 (N_9996,N_9536,N_9523);
xnor U9997 (N_9997,N_9506,N_9745);
and U9998 (N_9998,N_9724,N_9733);
nor U9999 (N_9999,N_9660,N_9607);
or U10000 (N_10000,N_9864,N_9983);
and U10001 (N_10001,N_9754,N_9777);
xnor U10002 (N_10002,N_9898,N_9902);
or U10003 (N_10003,N_9882,N_9766);
or U10004 (N_10004,N_9886,N_9827);
or U10005 (N_10005,N_9877,N_9867);
or U10006 (N_10006,N_9883,N_9838);
nor U10007 (N_10007,N_9800,N_9993);
nand U10008 (N_10008,N_9881,N_9973);
or U10009 (N_10009,N_9907,N_9940);
or U10010 (N_10010,N_9924,N_9795);
nor U10011 (N_10011,N_9843,N_9820);
nand U10012 (N_10012,N_9975,N_9752);
or U10013 (N_10013,N_9824,N_9835);
and U10014 (N_10014,N_9999,N_9914);
and U10015 (N_10015,N_9775,N_9758);
and U10016 (N_10016,N_9773,N_9751);
nor U10017 (N_10017,N_9842,N_9812);
nor U10018 (N_10018,N_9779,N_9788);
or U10019 (N_10019,N_9992,N_9929);
nand U10020 (N_10020,N_9998,N_9792);
nor U10021 (N_10021,N_9833,N_9997);
nand U10022 (N_10022,N_9769,N_9778);
nor U10023 (N_10023,N_9958,N_9826);
or U10024 (N_10024,N_9763,N_9834);
or U10025 (N_10025,N_9938,N_9948);
nor U10026 (N_10026,N_9819,N_9985);
nor U10027 (N_10027,N_9863,N_9967);
or U10028 (N_10028,N_9846,N_9950);
xor U10029 (N_10029,N_9815,N_9793);
nand U10030 (N_10030,N_9963,N_9784);
and U10031 (N_10031,N_9830,N_9771);
xor U10032 (N_10032,N_9971,N_9980);
nand U10033 (N_10033,N_9908,N_9951);
or U10034 (N_10034,N_9874,N_9939);
nand U10035 (N_10035,N_9935,N_9959);
nand U10036 (N_10036,N_9803,N_9957);
or U10037 (N_10037,N_9813,N_9972);
nand U10038 (N_10038,N_9979,N_9945);
xnor U10039 (N_10039,N_9790,N_9926);
nor U10040 (N_10040,N_9756,N_9851);
nor U10041 (N_10041,N_9844,N_9901);
and U10042 (N_10042,N_9772,N_9974);
or U10043 (N_10043,N_9767,N_9782);
or U10044 (N_10044,N_9814,N_9955);
nor U10045 (N_10045,N_9761,N_9854);
or U10046 (N_10046,N_9903,N_9866);
and U10047 (N_10047,N_9991,N_9897);
nor U10048 (N_10048,N_9910,N_9783);
and U10049 (N_10049,N_9934,N_9978);
and U10050 (N_10050,N_9868,N_9941);
and U10051 (N_10051,N_9984,N_9911);
nor U10052 (N_10052,N_9956,N_9770);
and U10053 (N_10053,N_9832,N_9762);
and U10054 (N_10054,N_9841,N_9930);
nand U10055 (N_10055,N_9927,N_9857);
xor U10056 (N_10056,N_9915,N_9932);
nand U10057 (N_10057,N_9764,N_9920);
nor U10058 (N_10058,N_9807,N_9797);
or U10059 (N_10059,N_9885,N_9946);
nand U10060 (N_10060,N_9949,N_9786);
nand U10061 (N_10061,N_9964,N_9858);
nor U10062 (N_10062,N_9892,N_9872);
xor U10063 (N_10063,N_9928,N_9899);
nor U10064 (N_10064,N_9982,N_9850);
xor U10065 (N_10065,N_9760,N_9925);
nor U10066 (N_10066,N_9869,N_9776);
xor U10067 (N_10067,N_9861,N_9822);
xnor U10068 (N_10068,N_9953,N_9961);
xnor U10069 (N_10069,N_9952,N_9848);
xnor U10070 (N_10070,N_9917,N_9798);
or U10071 (N_10071,N_9968,N_9805);
and U10072 (N_10072,N_9787,N_9870);
and U10073 (N_10073,N_9794,N_9876);
nor U10074 (N_10074,N_9774,N_9919);
xnor U10075 (N_10075,N_9871,N_9753);
or U10076 (N_10076,N_9806,N_9816);
xnor U10077 (N_10077,N_9913,N_9969);
nand U10078 (N_10078,N_9921,N_9799);
and U10079 (N_10079,N_9933,N_9765);
and U10080 (N_10080,N_9789,N_9845);
or U10081 (N_10081,N_9862,N_9994);
and U10082 (N_10082,N_9804,N_9852);
or U10083 (N_10083,N_9780,N_9900);
and U10084 (N_10084,N_9990,N_9808);
nor U10085 (N_10085,N_9890,N_9879);
and U10086 (N_10086,N_9801,N_9889);
xnor U10087 (N_10087,N_9759,N_9865);
or U10088 (N_10088,N_9965,N_9894);
nor U10089 (N_10089,N_9896,N_9937);
xor U10090 (N_10090,N_9856,N_9880);
and U10091 (N_10091,N_9796,N_9904);
nor U10092 (N_10092,N_9860,N_9916);
nor U10093 (N_10093,N_9887,N_9931);
or U10094 (N_10094,N_9970,N_9823);
and U10095 (N_10095,N_9986,N_9757);
xor U10096 (N_10096,N_9875,N_9909);
or U10097 (N_10097,N_9847,N_9987);
xor U10098 (N_10098,N_9923,N_9895);
or U10099 (N_10099,N_9849,N_9831);
xnor U10100 (N_10100,N_9791,N_9817);
nand U10101 (N_10101,N_9981,N_9878);
nand U10102 (N_10102,N_9977,N_9855);
or U10103 (N_10103,N_9809,N_9960);
xor U10104 (N_10104,N_9829,N_9966);
nand U10105 (N_10105,N_9922,N_9947);
nand U10106 (N_10106,N_9884,N_9810);
or U10107 (N_10107,N_9839,N_9785);
xor U10108 (N_10108,N_9821,N_9781);
xor U10109 (N_10109,N_9825,N_9853);
nor U10110 (N_10110,N_9840,N_9918);
and U10111 (N_10111,N_9768,N_9905);
and U10112 (N_10112,N_9818,N_9906);
and U10113 (N_10113,N_9888,N_9962);
nor U10114 (N_10114,N_9837,N_9954);
nor U10115 (N_10115,N_9755,N_9988);
or U10116 (N_10116,N_9859,N_9943);
xnor U10117 (N_10117,N_9828,N_9836);
nand U10118 (N_10118,N_9944,N_9893);
and U10119 (N_10119,N_9802,N_9873);
nor U10120 (N_10120,N_9989,N_9912);
nand U10121 (N_10121,N_9976,N_9995);
and U10122 (N_10122,N_9936,N_9811);
and U10123 (N_10123,N_9942,N_9750);
nor U10124 (N_10124,N_9996,N_9891);
or U10125 (N_10125,N_9863,N_9873);
and U10126 (N_10126,N_9842,N_9795);
or U10127 (N_10127,N_9995,N_9885);
xor U10128 (N_10128,N_9867,N_9787);
and U10129 (N_10129,N_9865,N_9811);
and U10130 (N_10130,N_9947,N_9907);
and U10131 (N_10131,N_9970,N_9888);
and U10132 (N_10132,N_9959,N_9957);
and U10133 (N_10133,N_9772,N_9759);
nor U10134 (N_10134,N_9904,N_9798);
nor U10135 (N_10135,N_9873,N_9940);
and U10136 (N_10136,N_9929,N_9790);
nand U10137 (N_10137,N_9882,N_9834);
xnor U10138 (N_10138,N_9897,N_9988);
nor U10139 (N_10139,N_9850,N_9774);
and U10140 (N_10140,N_9823,N_9948);
xnor U10141 (N_10141,N_9881,N_9798);
xor U10142 (N_10142,N_9776,N_9800);
and U10143 (N_10143,N_9875,N_9873);
xor U10144 (N_10144,N_9894,N_9957);
or U10145 (N_10145,N_9925,N_9757);
nor U10146 (N_10146,N_9794,N_9958);
nor U10147 (N_10147,N_9995,N_9809);
or U10148 (N_10148,N_9797,N_9946);
or U10149 (N_10149,N_9933,N_9756);
or U10150 (N_10150,N_9936,N_9868);
xor U10151 (N_10151,N_9931,N_9820);
nand U10152 (N_10152,N_9857,N_9982);
nor U10153 (N_10153,N_9944,N_9806);
nand U10154 (N_10154,N_9921,N_9775);
nor U10155 (N_10155,N_9811,N_9750);
or U10156 (N_10156,N_9932,N_9953);
and U10157 (N_10157,N_9835,N_9831);
and U10158 (N_10158,N_9942,N_9863);
xnor U10159 (N_10159,N_9752,N_9781);
or U10160 (N_10160,N_9908,N_9929);
nor U10161 (N_10161,N_9763,N_9779);
nor U10162 (N_10162,N_9989,N_9890);
and U10163 (N_10163,N_9889,N_9819);
nor U10164 (N_10164,N_9862,N_9999);
nand U10165 (N_10165,N_9954,N_9851);
xor U10166 (N_10166,N_9840,N_9980);
and U10167 (N_10167,N_9751,N_9910);
xor U10168 (N_10168,N_9805,N_9907);
nand U10169 (N_10169,N_9832,N_9952);
and U10170 (N_10170,N_9816,N_9926);
xor U10171 (N_10171,N_9885,N_9840);
xnor U10172 (N_10172,N_9941,N_9812);
nor U10173 (N_10173,N_9988,N_9809);
nor U10174 (N_10174,N_9812,N_9939);
and U10175 (N_10175,N_9923,N_9959);
nand U10176 (N_10176,N_9939,N_9752);
xnor U10177 (N_10177,N_9872,N_9930);
or U10178 (N_10178,N_9997,N_9809);
nand U10179 (N_10179,N_9915,N_9975);
and U10180 (N_10180,N_9870,N_9977);
nand U10181 (N_10181,N_9932,N_9772);
xor U10182 (N_10182,N_9844,N_9764);
or U10183 (N_10183,N_9775,N_9976);
or U10184 (N_10184,N_9795,N_9952);
and U10185 (N_10185,N_9925,N_9872);
xor U10186 (N_10186,N_9899,N_9924);
xor U10187 (N_10187,N_9888,N_9765);
nor U10188 (N_10188,N_9861,N_9817);
xnor U10189 (N_10189,N_9984,N_9959);
xnor U10190 (N_10190,N_9887,N_9925);
nor U10191 (N_10191,N_9998,N_9788);
nand U10192 (N_10192,N_9799,N_9855);
xor U10193 (N_10193,N_9957,N_9850);
nor U10194 (N_10194,N_9816,N_9918);
nand U10195 (N_10195,N_9843,N_9953);
xor U10196 (N_10196,N_9938,N_9898);
or U10197 (N_10197,N_9798,N_9901);
and U10198 (N_10198,N_9823,N_9946);
or U10199 (N_10199,N_9771,N_9941);
nor U10200 (N_10200,N_9908,N_9980);
nor U10201 (N_10201,N_9802,N_9939);
nand U10202 (N_10202,N_9890,N_9911);
or U10203 (N_10203,N_9809,N_9864);
nand U10204 (N_10204,N_9923,N_9854);
or U10205 (N_10205,N_9974,N_9944);
and U10206 (N_10206,N_9979,N_9922);
nand U10207 (N_10207,N_9844,N_9756);
xnor U10208 (N_10208,N_9779,N_9967);
or U10209 (N_10209,N_9781,N_9909);
xnor U10210 (N_10210,N_9802,N_9821);
nand U10211 (N_10211,N_9959,N_9876);
xnor U10212 (N_10212,N_9775,N_9785);
nand U10213 (N_10213,N_9900,N_9918);
and U10214 (N_10214,N_9959,N_9854);
nand U10215 (N_10215,N_9796,N_9882);
nand U10216 (N_10216,N_9929,N_9753);
and U10217 (N_10217,N_9934,N_9999);
and U10218 (N_10218,N_9876,N_9995);
nor U10219 (N_10219,N_9750,N_9792);
xnor U10220 (N_10220,N_9856,N_9841);
or U10221 (N_10221,N_9988,N_9780);
or U10222 (N_10222,N_9945,N_9914);
nand U10223 (N_10223,N_9797,N_9973);
xnor U10224 (N_10224,N_9983,N_9970);
and U10225 (N_10225,N_9778,N_9877);
or U10226 (N_10226,N_9962,N_9797);
nand U10227 (N_10227,N_9768,N_9931);
xnor U10228 (N_10228,N_9878,N_9776);
and U10229 (N_10229,N_9818,N_9988);
and U10230 (N_10230,N_9954,N_9771);
or U10231 (N_10231,N_9933,N_9895);
nand U10232 (N_10232,N_9907,N_9753);
or U10233 (N_10233,N_9800,N_9891);
and U10234 (N_10234,N_9997,N_9807);
nand U10235 (N_10235,N_9943,N_9852);
nand U10236 (N_10236,N_9907,N_9950);
xnor U10237 (N_10237,N_9905,N_9885);
nand U10238 (N_10238,N_9977,N_9958);
nor U10239 (N_10239,N_9795,N_9910);
or U10240 (N_10240,N_9757,N_9980);
nand U10241 (N_10241,N_9808,N_9904);
and U10242 (N_10242,N_9756,N_9987);
and U10243 (N_10243,N_9923,N_9873);
and U10244 (N_10244,N_9933,N_9793);
and U10245 (N_10245,N_9819,N_9958);
nand U10246 (N_10246,N_9780,N_9913);
and U10247 (N_10247,N_9856,N_9991);
nand U10248 (N_10248,N_9868,N_9886);
xor U10249 (N_10249,N_9964,N_9989);
nand U10250 (N_10250,N_10105,N_10236);
nand U10251 (N_10251,N_10219,N_10147);
xnor U10252 (N_10252,N_10052,N_10034);
or U10253 (N_10253,N_10031,N_10049);
and U10254 (N_10254,N_10177,N_10004);
nor U10255 (N_10255,N_10104,N_10142);
xor U10256 (N_10256,N_10221,N_10126);
nand U10257 (N_10257,N_10077,N_10240);
nand U10258 (N_10258,N_10124,N_10214);
and U10259 (N_10259,N_10098,N_10204);
nand U10260 (N_10260,N_10080,N_10216);
xnor U10261 (N_10261,N_10001,N_10086);
xor U10262 (N_10262,N_10011,N_10066);
and U10263 (N_10263,N_10097,N_10170);
or U10264 (N_10264,N_10195,N_10133);
nand U10265 (N_10265,N_10184,N_10227);
nand U10266 (N_10266,N_10128,N_10106);
or U10267 (N_10267,N_10220,N_10159);
nor U10268 (N_10268,N_10182,N_10012);
or U10269 (N_10269,N_10215,N_10107);
or U10270 (N_10270,N_10055,N_10043);
or U10271 (N_10271,N_10030,N_10063);
nand U10272 (N_10272,N_10051,N_10189);
nand U10273 (N_10273,N_10226,N_10158);
and U10274 (N_10274,N_10244,N_10185);
or U10275 (N_10275,N_10025,N_10103);
or U10276 (N_10276,N_10153,N_10115);
nand U10277 (N_10277,N_10246,N_10074);
nand U10278 (N_10278,N_10238,N_10163);
nor U10279 (N_10279,N_10019,N_10209);
and U10280 (N_10280,N_10053,N_10151);
or U10281 (N_10281,N_10213,N_10002);
nand U10282 (N_10282,N_10165,N_10175);
and U10283 (N_10283,N_10041,N_10248);
xor U10284 (N_10284,N_10181,N_10218);
and U10285 (N_10285,N_10167,N_10241);
nand U10286 (N_10286,N_10135,N_10129);
xnor U10287 (N_10287,N_10130,N_10060);
xnor U10288 (N_10288,N_10040,N_10143);
xor U10289 (N_10289,N_10186,N_10026);
and U10290 (N_10290,N_10206,N_10141);
nand U10291 (N_10291,N_10071,N_10148);
nand U10292 (N_10292,N_10044,N_10162);
nand U10293 (N_10293,N_10078,N_10145);
or U10294 (N_10294,N_10171,N_10229);
nand U10295 (N_10295,N_10082,N_10146);
xnor U10296 (N_10296,N_10038,N_10224);
nor U10297 (N_10297,N_10211,N_10247);
and U10298 (N_10298,N_10111,N_10007);
nand U10299 (N_10299,N_10168,N_10010);
nor U10300 (N_10300,N_10203,N_10091);
nand U10301 (N_10301,N_10072,N_10099);
or U10302 (N_10302,N_10188,N_10137);
or U10303 (N_10303,N_10174,N_10056);
nor U10304 (N_10304,N_10036,N_10197);
xnor U10305 (N_10305,N_10102,N_10067);
and U10306 (N_10306,N_10008,N_10176);
and U10307 (N_10307,N_10085,N_10234);
nand U10308 (N_10308,N_10222,N_10233);
nand U10309 (N_10309,N_10155,N_10088);
nand U10310 (N_10310,N_10015,N_10118);
nand U10311 (N_10311,N_10054,N_10033);
nor U10312 (N_10312,N_10223,N_10164);
xor U10313 (N_10313,N_10122,N_10050);
and U10314 (N_10314,N_10200,N_10110);
or U10315 (N_10315,N_10138,N_10140);
xor U10316 (N_10316,N_10125,N_10112);
and U10317 (N_10317,N_10190,N_10009);
or U10318 (N_10318,N_10210,N_10076);
and U10319 (N_10319,N_10139,N_10116);
xnor U10320 (N_10320,N_10114,N_10178);
nand U10321 (N_10321,N_10230,N_10196);
xnor U10322 (N_10322,N_10021,N_10217);
xor U10323 (N_10323,N_10149,N_10160);
or U10324 (N_10324,N_10023,N_10006);
xnor U10325 (N_10325,N_10249,N_10132);
and U10326 (N_10326,N_10027,N_10192);
nor U10327 (N_10327,N_10093,N_10113);
or U10328 (N_10328,N_10003,N_10117);
xor U10329 (N_10329,N_10096,N_10144);
nand U10330 (N_10330,N_10119,N_10242);
or U10331 (N_10331,N_10013,N_10205);
or U10332 (N_10332,N_10069,N_10062);
xnor U10333 (N_10333,N_10235,N_10231);
nand U10334 (N_10334,N_10068,N_10032);
and U10335 (N_10335,N_10123,N_10014);
nand U10336 (N_10336,N_10207,N_10092);
nor U10337 (N_10337,N_10059,N_10057);
nor U10338 (N_10338,N_10191,N_10081);
nand U10339 (N_10339,N_10198,N_10073);
or U10340 (N_10340,N_10161,N_10193);
xnor U10341 (N_10341,N_10212,N_10187);
and U10342 (N_10342,N_10134,N_10087);
xnor U10343 (N_10343,N_10228,N_10039);
xor U10344 (N_10344,N_10243,N_10048);
or U10345 (N_10345,N_10127,N_10237);
or U10346 (N_10346,N_10180,N_10100);
xnor U10347 (N_10347,N_10016,N_10037);
nand U10348 (N_10348,N_10108,N_10109);
xor U10349 (N_10349,N_10183,N_10199);
or U10350 (N_10350,N_10046,N_10131);
and U10351 (N_10351,N_10232,N_10121);
nor U10352 (N_10352,N_10194,N_10064);
nand U10353 (N_10353,N_10154,N_10061);
xnor U10354 (N_10354,N_10156,N_10101);
xnor U10355 (N_10355,N_10208,N_10172);
or U10356 (N_10356,N_10045,N_10173);
xor U10357 (N_10357,N_10042,N_10090);
or U10358 (N_10358,N_10245,N_10065);
xor U10359 (N_10359,N_10169,N_10239);
and U10360 (N_10360,N_10084,N_10157);
xnor U10361 (N_10361,N_10058,N_10202);
nor U10362 (N_10362,N_10029,N_10152);
and U10363 (N_10363,N_10094,N_10075);
or U10364 (N_10364,N_10047,N_10028);
xor U10365 (N_10365,N_10089,N_10166);
nand U10366 (N_10366,N_10018,N_10005);
xor U10367 (N_10367,N_10120,N_10136);
nand U10368 (N_10368,N_10017,N_10035);
or U10369 (N_10369,N_10024,N_10225);
or U10370 (N_10370,N_10020,N_10000);
or U10371 (N_10371,N_10083,N_10095);
and U10372 (N_10372,N_10070,N_10179);
or U10373 (N_10373,N_10079,N_10201);
nand U10374 (N_10374,N_10022,N_10150);
or U10375 (N_10375,N_10032,N_10241);
and U10376 (N_10376,N_10069,N_10197);
nand U10377 (N_10377,N_10221,N_10212);
and U10378 (N_10378,N_10218,N_10214);
nand U10379 (N_10379,N_10024,N_10069);
or U10380 (N_10380,N_10113,N_10248);
xor U10381 (N_10381,N_10096,N_10207);
and U10382 (N_10382,N_10071,N_10235);
xnor U10383 (N_10383,N_10235,N_10060);
xor U10384 (N_10384,N_10237,N_10081);
nand U10385 (N_10385,N_10180,N_10078);
nor U10386 (N_10386,N_10183,N_10162);
nor U10387 (N_10387,N_10093,N_10227);
or U10388 (N_10388,N_10149,N_10055);
xnor U10389 (N_10389,N_10078,N_10021);
xor U10390 (N_10390,N_10021,N_10188);
xor U10391 (N_10391,N_10246,N_10052);
nand U10392 (N_10392,N_10165,N_10226);
nor U10393 (N_10393,N_10215,N_10051);
nand U10394 (N_10394,N_10218,N_10201);
or U10395 (N_10395,N_10086,N_10128);
and U10396 (N_10396,N_10033,N_10240);
xnor U10397 (N_10397,N_10131,N_10154);
nor U10398 (N_10398,N_10165,N_10114);
and U10399 (N_10399,N_10209,N_10005);
and U10400 (N_10400,N_10132,N_10115);
or U10401 (N_10401,N_10163,N_10157);
nor U10402 (N_10402,N_10044,N_10056);
and U10403 (N_10403,N_10125,N_10003);
nor U10404 (N_10404,N_10211,N_10106);
nor U10405 (N_10405,N_10123,N_10233);
and U10406 (N_10406,N_10024,N_10103);
xnor U10407 (N_10407,N_10128,N_10244);
nor U10408 (N_10408,N_10179,N_10005);
xnor U10409 (N_10409,N_10225,N_10013);
nor U10410 (N_10410,N_10075,N_10074);
nor U10411 (N_10411,N_10110,N_10231);
and U10412 (N_10412,N_10128,N_10076);
and U10413 (N_10413,N_10175,N_10062);
xnor U10414 (N_10414,N_10032,N_10236);
nand U10415 (N_10415,N_10132,N_10045);
xor U10416 (N_10416,N_10223,N_10056);
nor U10417 (N_10417,N_10227,N_10049);
nand U10418 (N_10418,N_10136,N_10206);
and U10419 (N_10419,N_10203,N_10187);
nand U10420 (N_10420,N_10076,N_10192);
and U10421 (N_10421,N_10238,N_10079);
nor U10422 (N_10422,N_10096,N_10012);
nand U10423 (N_10423,N_10170,N_10079);
nor U10424 (N_10424,N_10185,N_10201);
nor U10425 (N_10425,N_10118,N_10192);
and U10426 (N_10426,N_10234,N_10163);
and U10427 (N_10427,N_10207,N_10183);
or U10428 (N_10428,N_10137,N_10072);
nand U10429 (N_10429,N_10121,N_10144);
nor U10430 (N_10430,N_10246,N_10195);
nor U10431 (N_10431,N_10047,N_10140);
or U10432 (N_10432,N_10089,N_10203);
or U10433 (N_10433,N_10143,N_10062);
xnor U10434 (N_10434,N_10193,N_10042);
and U10435 (N_10435,N_10053,N_10244);
nand U10436 (N_10436,N_10087,N_10183);
xor U10437 (N_10437,N_10102,N_10168);
or U10438 (N_10438,N_10064,N_10117);
nand U10439 (N_10439,N_10243,N_10239);
xor U10440 (N_10440,N_10123,N_10101);
nor U10441 (N_10441,N_10214,N_10217);
or U10442 (N_10442,N_10130,N_10044);
nor U10443 (N_10443,N_10104,N_10033);
nand U10444 (N_10444,N_10050,N_10086);
and U10445 (N_10445,N_10198,N_10096);
xor U10446 (N_10446,N_10229,N_10133);
nor U10447 (N_10447,N_10061,N_10191);
and U10448 (N_10448,N_10176,N_10032);
and U10449 (N_10449,N_10199,N_10053);
nand U10450 (N_10450,N_10222,N_10244);
xnor U10451 (N_10451,N_10024,N_10166);
or U10452 (N_10452,N_10206,N_10150);
xor U10453 (N_10453,N_10241,N_10080);
nand U10454 (N_10454,N_10005,N_10165);
and U10455 (N_10455,N_10137,N_10228);
or U10456 (N_10456,N_10192,N_10046);
nor U10457 (N_10457,N_10169,N_10240);
and U10458 (N_10458,N_10013,N_10248);
nand U10459 (N_10459,N_10068,N_10130);
and U10460 (N_10460,N_10169,N_10067);
and U10461 (N_10461,N_10199,N_10127);
and U10462 (N_10462,N_10180,N_10175);
nand U10463 (N_10463,N_10176,N_10036);
nor U10464 (N_10464,N_10021,N_10060);
and U10465 (N_10465,N_10236,N_10184);
xnor U10466 (N_10466,N_10025,N_10193);
xor U10467 (N_10467,N_10076,N_10119);
nor U10468 (N_10468,N_10191,N_10028);
xor U10469 (N_10469,N_10248,N_10217);
and U10470 (N_10470,N_10106,N_10031);
and U10471 (N_10471,N_10245,N_10093);
nand U10472 (N_10472,N_10212,N_10004);
xnor U10473 (N_10473,N_10147,N_10169);
and U10474 (N_10474,N_10214,N_10170);
nand U10475 (N_10475,N_10033,N_10207);
and U10476 (N_10476,N_10222,N_10067);
nor U10477 (N_10477,N_10070,N_10048);
and U10478 (N_10478,N_10044,N_10224);
nor U10479 (N_10479,N_10109,N_10224);
nor U10480 (N_10480,N_10133,N_10138);
or U10481 (N_10481,N_10163,N_10155);
nor U10482 (N_10482,N_10089,N_10038);
or U10483 (N_10483,N_10151,N_10007);
or U10484 (N_10484,N_10036,N_10231);
nand U10485 (N_10485,N_10084,N_10099);
xor U10486 (N_10486,N_10102,N_10012);
or U10487 (N_10487,N_10098,N_10009);
nand U10488 (N_10488,N_10243,N_10148);
or U10489 (N_10489,N_10225,N_10057);
nor U10490 (N_10490,N_10185,N_10128);
or U10491 (N_10491,N_10171,N_10203);
and U10492 (N_10492,N_10114,N_10069);
nor U10493 (N_10493,N_10116,N_10164);
xnor U10494 (N_10494,N_10142,N_10191);
nand U10495 (N_10495,N_10234,N_10079);
and U10496 (N_10496,N_10007,N_10231);
and U10497 (N_10497,N_10075,N_10178);
nand U10498 (N_10498,N_10004,N_10102);
or U10499 (N_10499,N_10243,N_10039);
and U10500 (N_10500,N_10423,N_10404);
or U10501 (N_10501,N_10360,N_10431);
nor U10502 (N_10502,N_10275,N_10399);
nand U10503 (N_10503,N_10499,N_10298);
or U10504 (N_10504,N_10428,N_10293);
and U10505 (N_10505,N_10424,N_10339);
nor U10506 (N_10506,N_10322,N_10351);
nor U10507 (N_10507,N_10392,N_10391);
nor U10508 (N_10508,N_10343,N_10363);
xnor U10509 (N_10509,N_10472,N_10478);
or U10510 (N_10510,N_10488,N_10303);
or U10511 (N_10511,N_10356,N_10301);
or U10512 (N_10512,N_10324,N_10496);
nand U10513 (N_10513,N_10443,N_10290);
nor U10514 (N_10514,N_10385,N_10331);
nor U10515 (N_10515,N_10476,N_10349);
xnor U10516 (N_10516,N_10289,N_10381);
xnor U10517 (N_10517,N_10276,N_10283);
nand U10518 (N_10518,N_10386,N_10317);
or U10519 (N_10519,N_10461,N_10483);
or U10520 (N_10520,N_10313,N_10361);
or U10521 (N_10521,N_10414,N_10316);
nand U10522 (N_10522,N_10440,N_10256);
nand U10523 (N_10523,N_10375,N_10444);
nor U10524 (N_10524,N_10305,N_10364);
nand U10525 (N_10525,N_10449,N_10353);
nand U10526 (N_10526,N_10441,N_10292);
or U10527 (N_10527,N_10480,N_10378);
nor U10528 (N_10528,N_10346,N_10421);
or U10529 (N_10529,N_10307,N_10314);
nor U10530 (N_10530,N_10420,N_10335);
or U10531 (N_10531,N_10451,N_10485);
nor U10532 (N_10532,N_10255,N_10296);
and U10533 (N_10533,N_10416,N_10342);
nand U10534 (N_10534,N_10358,N_10474);
xor U10535 (N_10535,N_10332,N_10365);
or U10536 (N_10536,N_10486,N_10250);
nor U10537 (N_10537,N_10412,N_10409);
and U10538 (N_10538,N_10294,N_10334);
and U10539 (N_10539,N_10415,N_10453);
and U10540 (N_10540,N_10446,N_10475);
xnor U10541 (N_10541,N_10284,N_10460);
or U10542 (N_10542,N_10271,N_10394);
nand U10543 (N_10543,N_10434,N_10437);
or U10544 (N_10544,N_10436,N_10253);
nor U10545 (N_10545,N_10383,N_10388);
and U10546 (N_10546,N_10273,N_10297);
nor U10547 (N_10547,N_10291,N_10479);
or U10548 (N_10548,N_10402,N_10477);
or U10549 (N_10549,N_10310,N_10309);
nand U10550 (N_10550,N_10393,N_10493);
nor U10551 (N_10551,N_10374,N_10265);
nand U10552 (N_10552,N_10400,N_10266);
or U10553 (N_10553,N_10379,N_10376);
or U10554 (N_10554,N_10464,N_10347);
xor U10555 (N_10555,N_10492,N_10359);
and U10556 (N_10556,N_10278,N_10405);
or U10557 (N_10557,N_10457,N_10319);
nand U10558 (N_10558,N_10491,N_10348);
or U10559 (N_10559,N_10323,N_10268);
xnor U10560 (N_10560,N_10261,N_10368);
or U10561 (N_10561,N_10272,N_10285);
nor U10562 (N_10562,N_10338,N_10411);
and U10563 (N_10563,N_10419,N_10299);
xnor U10564 (N_10564,N_10279,N_10321);
or U10565 (N_10565,N_10287,N_10442);
and U10566 (N_10566,N_10466,N_10468);
and U10567 (N_10567,N_10328,N_10270);
and U10568 (N_10568,N_10395,N_10311);
xor U10569 (N_10569,N_10445,N_10280);
or U10570 (N_10570,N_10295,N_10315);
nand U10571 (N_10571,N_10462,N_10403);
or U10572 (N_10572,N_10465,N_10390);
nor U10573 (N_10573,N_10470,N_10267);
and U10574 (N_10574,N_10452,N_10432);
nor U10575 (N_10575,N_10454,N_10329);
and U10576 (N_10576,N_10447,N_10357);
nand U10577 (N_10577,N_10340,N_10387);
or U10578 (N_10578,N_10308,N_10281);
and U10579 (N_10579,N_10397,N_10463);
or U10580 (N_10580,N_10302,N_10481);
and U10581 (N_10581,N_10337,N_10254);
or U10582 (N_10582,N_10330,N_10352);
nor U10583 (N_10583,N_10336,N_10427);
nand U10584 (N_10584,N_10407,N_10258);
xor U10585 (N_10585,N_10277,N_10413);
or U10586 (N_10586,N_10372,N_10312);
xnor U10587 (N_10587,N_10433,N_10429);
or U10588 (N_10588,N_10450,N_10344);
and U10589 (N_10589,N_10487,N_10435);
nor U10590 (N_10590,N_10467,N_10439);
nor U10591 (N_10591,N_10426,N_10469);
xnor U10592 (N_10592,N_10326,N_10497);
or U10593 (N_10593,N_10263,N_10389);
nor U10594 (N_10594,N_10373,N_10382);
or U10595 (N_10595,N_10396,N_10471);
and U10596 (N_10596,N_10425,N_10341);
nor U10597 (N_10597,N_10345,N_10448);
or U10598 (N_10598,N_10438,N_10430);
or U10599 (N_10599,N_10362,N_10484);
or U10600 (N_10600,N_10300,N_10350);
nor U10601 (N_10601,N_10417,N_10251);
and U10602 (N_10602,N_10274,N_10327);
xnor U10603 (N_10603,N_10366,N_10418);
xor U10604 (N_10604,N_10354,N_10288);
nand U10605 (N_10605,N_10286,N_10380);
and U10606 (N_10606,N_10406,N_10259);
nand U10607 (N_10607,N_10422,N_10495);
or U10608 (N_10608,N_10490,N_10252);
nand U10609 (N_10609,N_10456,N_10369);
nor U10610 (N_10610,N_10257,N_10384);
nand U10611 (N_10611,N_10498,N_10458);
nand U10612 (N_10612,N_10408,N_10282);
nand U10613 (N_10613,N_10370,N_10264);
and U10614 (N_10614,N_10455,N_10489);
nor U10615 (N_10615,N_10410,N_10401);
and U10616 (N_10616,N_10333,N_10260);
nor U10617 (N_10617,N_10318,N_10398);
nor U10618 (N_10618,N_10325,N_10269);
xnor U10619 (N_10619,N_10320,N_10494);
xnor U10620 (N_10620,N_10473,N_10304);
nand U10621 (N_10621,N_10482,N_10367);
and U10622 (N_10622,N_10355,N_10459);
or U10623 (N_10623,N_10306,N_10377);
nor U10624 (N_10624,N_10371,N_10262);
nor U10625 (N_10625,N_10405,N_10376);
nor U10626 (N_10626,N_10458,N_10300);
nor U10627 (N_10627,N_10369,N_10286);
nand U10628 (N_10628,N_10416,N_10494);
nor U10629 (N_10629,N_10470,N_10429);
or U10630 (N_10630,N_10428,N_10475);
nor U10631 (N_10631,N_10456,N_10402);
nor U10632 (N_10632,N_10342,N_10465);
nor U10633 (N_10633,N_10424,N_10479);
nand U10634 (N_10634,N_10477,N_10443);
xor U10635 (N_10635,N_10456,N_10395);
nor U10636 (N_10636,N_10469,N_10265);
or U10637 (N_10637,N_10330,N_10441);
and U10638 (N_10638,N_10410,N_10468);
xnor U10639 (N_10639,N_10376,N_10274);
or U10640 (N_10640,N_10268,N_10365);
xnor U10641 (N_10641,N_10330,N_10361);
and U10642 (N_10642,N_10488,N_10292);
xnor U10643 (N_10643,N_10344,N_10267);
and U10644 (N_10644,N_10366,N_10335);
or U10645 (N_10645,N_10364,N_10286);
xnor U10646 (N_10646,N_10322,N_10477);
or U10647 (N_10647,N_10348,N_10342);
xor U10648 (N_10648,N_10385,N_10409);
nor U10649 (N_10649,N_10495,N_10406);
nand U10650 (N_10650,N_10282,N_10275);
nor U10651 (N_10651,N_10441,N_10346);
or U10652 (N_10652,N_10260,N_10327);
nor U10653 (N_10653,N_10401,N_10408);
nand U10654 (N_10654,N_10485,N_10362);
nor U10655 (N_10655,N_10466,N_10445);
nand U10656 (N_10656,N_10436,N_10373);
nand U10657 (N_10657,N_10365,N_10435);
nor U10658 (N_10658,N_10482,N_10475);
xor U10659 (N_10659,N_10465,N_10433);
nor U10660 (N_10660,N_10431,N_10347);
nor U10661 (N_10661,N_10431,N_10358);
and U10662 (N_10662,N_10309,N_10436);
or U10663 (N_10663,N_10364,N_10371);
nand U10664 (N_10664,N_10272,N_10290);
nor U10665 (N_10665,N_10475,N_10341);
xor U10666 (N_10666,N_10464,N_10293);
nand U10667 (N_10667,N_10376,N_10371);
and U10668 (N_10668,N_10442,N_10497);
or U10669 (N_10669,N_10431,N_10463);
xnor U10670 (N_10670,N_10448,N_10254);
and U10671 (N_10671,N_10299,N_10468);
xnor U10672 (N_10672,N_10270,N_10337);
xnor U10673 (N_10673,N_10364,N_10398);
nand U10674 (N_10674,N_10415,N_10425);
nand U10675 (N_10675,N_10494,N_10289);
and U10676 (N_10676,N_10340,N_10477);
or U10677 (N_10677,N_10263,N_10258);
nand U10678 (N_10678,N_10471,N_10441);
nand U10679 (N_10679,N_10365,N_10429);
or U10680 (N_10680,N_10390,N_10426);
or U10681 (N_10681,N_10460,N_10339);
and U10682 (N_10682,N_10429,N_10258);
or U10683 (N_10683,N_10492,N_10402);
nor U10684 (N_10684,N_10272,N_10388);
nand U10685 (N_10685,N_10415,N_10407);
and U10686 (N_10686,N_10345,N_10456);
or U10687 (N_10687,N_10330,N_10281);
nor U10688 (N_10688,N_10370,N_10365);
nand U10689 (N_10689,N_10269,N_10439);
or U10690 (N_10690,N_10265,N_10311);
or U10691 (N_10691,N_10405,N_10328);
nand U10692 (N_10692,N_10326,N_10335);
xor U10693 (N_10693,N_10332,N_10436);
nor U10694 (N_10694,N_10298,N_10272);
nor U10695 (N_10695,N_10445,N_10480);
and U10696 (N_10696,N_10312,N_10350);
nand U10697 (N_10697,N_10427,N_10309);
nand U10698 (N_10698,N_10258,N_10340);
and U10699 (N_10699,N_10322,N_10406);
nor U10700 (N_10700,N_10361,N_10323);
or U10701 (N_10701,N_10286,N_10387);
nor U10702 (N_10702,N_10337,N_10442);
and U10703 (N_10703,N_10385,N_10422);
or U10704 (N_10704,N_10423,N_10460);
or U10705 (N_10705,N_10440,N_10449);
or U10706 (N_10706,N_10469,N_10276);
xnor U10707 (N_10707,N_10460,N_10436);
xnor U10708 (N_10708,N_10347,N_10326);
and U10709 (N_10709,N_10446,N_10388);
and U10710 (N_10710,N_10436,N_10375);
or U10711 (N_10711,N_10456,N_10265);
nand U10712 (N_10712,N_10299,N_10405);
and U10713 (N_10713,N_10293,N_10364);
xor U10714 (N_10714,N_10272,N_10394);
nand U10715 (N_10715,N_10311,N_10357);
and U10716 (N_10716,N_10424,N_10318);
or U10717 (N_10717,N_10470,N_10433);
nand U10718 (N_10718,N_10446,N_10339);
and U10719 (N_10719,N_10446,N_10334);
nand U10720 (N_10720,N_10311,N_10490);
or U10721 (N_10721,N_10282,N_10318);
nand U10722 (N_10722,N_10275,N_10453);
nand U10723 (N_10723,N_10466,N_10488);
xor U10724 (N_10724,N_10426,N_10498);
nand U10725 (N_10725,N_10432,N_10488);
nor U10726 (N_10726,N_10424,N_10387);
nand U10727 (N_10727,N_10318,N_10309);
nand U10728 (N_10728,N_10353,N_10345);
or U10729 (N_10729,N_10328,N_10436);
and U10730 (N_10730,N_10337,N_10252);
nor U10731 (N_10731,N_10468,N_10424);
xor U10732 (N_10732,N_10466,N_10253);
or U10733 (N_10733,N_10363,N_10255);
xnor U10734 (N_10734,N_10465,N_10327);
or U10735 (N_10735,N_10334,N_10435);
nand U10736 (N_10736,N_10334,N_10479);
nand U10737 (N_10737,N_10372,N_10274);
and U10738 (N_10738,N_10357,N_10364);
xnor U10739 (N_10739,N_10445,N_10339);
nor U10740 (N_10740,N_10438,N_10400);
or U10741 (N_10741,N_10414,N_10299);
or U10742 (N_10742,N_10329,N_10410);
nor U10743 (N_10743,N_10382,N_10288);
nor U10744 (N_10744,N_10251,N_10295);
xnor U10745 (N_10745,N_10468,N_10328);
or U10746 (N_10746,N_10412,N_10350);
nor U10747 (N_10747,N_10447,N_10375);
xnor U10748 (N_10748,N_10286,N_10390);
or U10749 (N_10749,N_10448,N_10310);
and U10750 (N_10750,N_10591,N_10614);
or U10751 (N_10751,N_10556,N_10653);
or U10752 (N_10752,N_10646,N_10601);
and U10753 (N_10753,N_10713,N_10658);
xor U10754 (N_10754,N_10534,N_10520);
nand U10755 (N_10755,N_10710,N_10530);
and U10756 (N_10756,N_10631,N_10542);
xnor U10757 (N_10757,N_10674,N_10627);
nand U10758 (N_10758,N_10505,N_10625);
nor U10759 (N_10759,N_10667,N_10599);
or U10760 (N_10760,N_10579,N_10689);
or U10761 (N_10761,N_10551,N_10654);
xor U10762 (N_10762,N_10616,N_10660);
xor U10763 (N_10763,N_10637,N_10528);
nand U10764 (N_10764,N_10736,N_10571);
and U10765 (N_10765,N_10547,N_10749);
or U10766 (N_10766,N_10583,N_10729);
nor U10767 (N_10767,N_10665,N_10582);
nor U10768 (N_10768,N_10629,N_10544);
and U10769 (N_10769,N_10586,N_10731);
nand U10770 (N_10770,N_10573,N_10561);
nand U10771 (N_10771,N_10694,N_10587);
and U10772 (N_10772,N_10640,N_10515);
or U10773 (N_10773,N_10503,N_10555);
nand U10774 (N_10774,N_10645,N_10568);
or U10775 (N_10775,N_10504,N_10572);
xor U10776 (N_10776,N_10514,N_10527);
and U10777 (N_10777,N_10558,N_10549);
and U10778 (N_10778,N_10683,N_10565);
or U10779 (N_10779,N_10663,N_10563);
and U10780 (N_10780,N_10622,N_10672);
and U10781 (N_10781,N_10747,N_10541);
and U10782 (N_10782,N_10634,N_10506);
nand U10783 (N_10783,N_10721,N_10662);
nand U10784 (N_10784,N_10709,N_10737);
and U10785 (N_10785,N_10724,N_10650);
or U10786 (N_10786,N_10589,N_10513);
nor U10787 (N_10787,N_10691,N_10636);
and U10788 (N_10788,N_10661,N_10603);
and U10789 (N_10789,N_10546,N_10562);
xor U10790 (N_10790,N_10719,N_10666);
xor U10791 (N_10791,N_10620,N_10693);
nand U10792 (N_10792,N_10669,N_10714);
nand U10793 (N_10793,N_10698,N_10643);
nand U10794 (N_10794,N_10604,N_10580);
and U10795 (N_10795,N_10681,N_10621);
nand U10796 (N_10796,N_10602,N_10739);
xnor U10797 (N_10797,N_10685,N_10688);
or U10798 (N_10798,N_10626,N_10679);
or U10799 (N_10799,N_10690,N_10639);
nor U10800 (N_10800,N_10595,N_10684);
nor U10801 (N_10801,N_10612,N_10619);
or U10802 (N_10802,N_10687,N_10536);
or U10803 (N_10803,N_10677,N_10664);
nor U10804 (N_10804,N_10744,N_10581);
or U10805 (N_10805,N_10577,N_10697);
and U10806 (N_10806,N_10720,N_10680);
xnor U10807 (N_10807,N_10559,N_10523);
nor U10808 (N_10808,N_10651,N_10567);
and U10809 (N_10809,N_10743,N_10531);
nand U10810 (N_10810,N_10524,N_10708);
and U10811 (N_10811,N_10598,N_10647);
and U10812 (N_10812,N_10615,N_10532);
or U10813 (N_10813,N_10593,N_10566);
xnor U10814 (N_10814,N_10733,N_10618);
xor U10815 (N_10815,N_10607,N_10500);
nand U10816 (N_10816,N_10734,N_10742);
xor U10817 (N_10817,N_10671,N_10537);
or U10818 (N_10818,N_10656,N_10746);
or U10819 (N_10819,N_10611,N_10699);
nand U10820 (N_10820,N_10552,N_10609);
nand U10821 (N_10821,N_10545,N_10550);
and U10822 (N_10822,N_10659,N_10707);
nand U10823 (N_10823,N_10727,N_10594);
xnor U10824 (N_10824,N_10512,N_10543);
nand U10825 (N_10825,N_10519,N_10738);
xnor U10826 (N_10826,N_10518,N_10717);
xnor U10827 (N_10827,N_10732,N_10696);
nor U10828 (N_10828,N_10722,N_10554);
nor U10829 (N_10829,N_10522,N_10592);
or U10830 (N_10830,N_10557,N_10569);
nand U10831 (N_10831,N_10501,N_10705);
nand U10832 (N_10832,N_10700,N_10649);
nand U10833 (N_10833,N_10570,N_10723);
nand U10834 (N_10834,N_10735,N_10711);
xor U10835 (N_10835,N_10686,N_10675);
nand U10836 (N_10836,N_10633,N_10624);
nand U10837 (N_10837,N_10652,N_10718);
or U10838 (N_10838,N_10578,N_10597);
or U10839 (N_10839,N_10668,N_10678);
or U10840 (N_10840,N_10682,N_10540);
and U10841 (N_10841,N_10517,N_10642);
xor U10842 (N_10842,N_10725,N_10605);
nor U10843 (N_10843,N_10606,N_10715);
and U10844 (N_10844,N_10521,N_10628);
and U10845 (N_10845,N_10730,N_10695);
nor U10846 (N_10846,N_10745,N_10638);
or U10847 (N_10847,N_10608,N_10748);
or U10848 (N_10848,N_10641,N_10526);
xor U10849 (N_10849,N_10701,N_10655);
xor U10850 (N_10850,N_10740,N_10692);
or U10851 (N_10851,N_10509,N_10535);
nand U10852 (N_10852,N_10673,N_10553);
xnor U10853 (N_10853,N_10574,N_10657);
and U10854 (N_10854,N_10644,N_10632);
or U10855 (N_10855,N_10617,N_10623);
and U10856 (N_10856,N_10511,N_10635);
or U10857 (N_10857,N_10548,N_10728);
or U10858 (N_10858,N_10610,N_10741);
nor U10859 (N_10859,N_10704,N_10510);
nand U10860 (N_10860,N_10670,N_10584);
nand U10861 (N_10861,N_10590,N_10596);
and U10862 (N_10862,N_10613,N_10676);
or U10863 (N_10863,N_10533,N_10716);
xor U10864 (N_10864,N_10600,N_10560);
nand U10865 (N_10865,N_10525,N_10508);
nor U10866 (N_10866,N_10702,N_10502);
or U10867 (N_10867,N_10507,N_10706);
and U10868 (N_10868,N_10564,N_10516);
nand U10869 (N_10869,N_10575,N_10588);
nand U10870 (N_10870,N_10726,N_10576);
xor U10871 (N_10871,N_10585,N_10539);
and U10872 (N_10872,N_10529,N_10648);
nand U10873 (N_10873,N_10538,N_10630);
nand U10874 (N_10874,N_10703,N_10712);
or U10875 (N_10875,N_10736,N_10664);
and U10876 (N_10876,N_10516,N_10693);
nand U10877 (N_10877,N_10542,N_10720);
nor U10878 (N_10878,N_10566,N_10602);
nand U10879 (N_10879,N_10514,N_10592);
nand U10880 (N_10880,N_10593,N_10743);
xnor U10881 (N_10881,N_10654,N_10711);
xor U10882 (N_10882,N_10749,N_10640);
nor U10883 (N_10883,N_10722,N_10505);
nand U10884 (N_10884,N_10554,N_10573);
and U10885 (N_10885,N_10586,N_10548);
xnor U10886 (N_10886,N_10555,N_10720);
nand U10887 (N_10887,N_10573,N_10569);
xor U10888 (N_10888,N_10712,N_10663);
nor U10889 (N_10889,N_10574,N_10529);
or U10890 (N_10890,N_10595,N_10589);
and U10891 (N_10891,N_10558,N_10502);
or U10892 (N_10892,N_10537,N_10684);
nor U10893 (N_10893,N_10708,N_10598);
or U10894 (N_10894,N_10728,N_10662);
or U10895 (N_10895,N_10577,N_10736);
nand U10896 (N_10896,N_10689,N_10644);
nand U10897 (N_10897,N_10607,N_10734);
and U10898 (N_10898,N_10566,N_10654);
nor U10899 (N_10899,N_10556,N_10737);
nand U10900 (N_10900,N_10549,N_10692);
or U10901 (N_10901,N_10675,N_10548);
xnor U10902 (N_10902,N_10690,N_10518);
or U10903 (N_10903,N_10675,N_10632);
nor U10904 (N_10904,N_10679,N_10605);
or U10905 (N_10905,N_10504,N_10628);
or U10906 (N_10906,N_10502,N_10726);
and U10907 (N_10907,N_10652,N_10557);
nor U10908 (N_10908,N_10725,N_10695);
and U10909 (N_10909,N_10602,N_10729);
or U10910 (N_10910,N_10621,N_10540);
and U10911 (N_10911,N_10701,N_10733);
and U10912 (N_10912,N_10518,N_10650);
and U10913 (N_10913,N_10536,N_10553);
xnor U10914 (N_10914,N_10592,N_10656);
nor U10915 (N_10915,N_10711,N_10586);
nor U10916 (N_10916,N_10635,N_10706);
nor U10917 (N_10917,N_10728,N_10516);
or U10918 (N_10918,N_10668,N_10685);
and U10919 (N_10919,N_10647,N_10612);
nand U10920 (N_10920,N_10537,N_10717);
nor U10921 (N_10921,N_10565,N_10512);
xnor U10922 (N_10922,N_10740,N_10507);
xnor U10923 (N_10923,N_10519,N_10692);
or U10924 (N_10924,N_10651,N_10598);
xor U10925 (N_10925,N_10727,N_10549);
and U10926 (N_10926,N_10695,N_10723);
nor U10927 (N_10927,N_10580,N_10546);
nand U10928 (N_10928,N_10525,N_10708);
or U10929 (N_10929,N_10608,N_10536);
nand U10930 (N_10930,N_10538,N_10670);
xor U10931 (N_10931,N_10538,N_10687);
nor U10932 (N_10932,N_10584,N_10659);
xor U10933 (N_10933,N_10539,N_10542);
nor U10934 (N_10934,N_10600,N_10559);
or U10935 (N_10935,N_10611,N_10551);
xor U10936 (N_10936,N_10743,N_10546);
or U10937 (N_10937,N_10569,N_10628);
and U10938 (N_10938,N_10672,N_10520);
nor U10939 (N_10939,N_10713,N_10670);
or U10940 (N_10940,N_10651,N_10641);
xnor U10941 (N_10941,N_10538,N_10552);
or U10942 (N_10942,N_10730,N_10689);
or U10943 (N_10943,N_10614,N_10598);
xnor U10944 (N_10944,N_10583,N_10567);
or U10945 (N_10945,N_10641,N_10659);
nand U10946 (N_10946,N_10542,N_10705);
and U10947 (N_10947,N_10715,N_10683);
or U10948 (N_10948,N_10695,N_10656);
or U10949 (N_10949,N_10646,N_10686);
or U10950 (N_10950,N_10733,N_10524);
or U10951 (N_10951,N_10643,N_10681);
nand U10952 (N_10952,N_10602,N_10626);
or U10953 (N_10953,N_10513,N_10705);
nor U10954 (N_10954,N_10587,N_10616);
xnor U10955 (N_10955,N_10511,N_10700);
nor U10956 (N_10956,N_10535,N_10717);
or U10957 (N_10957,N_10709,N_10662);
nor U10958 (N_10958,N_10514,N_10661);
xnor U10959 (N_10959,N_10605,N_10517);
and U10960 (N_10960,N_10530,N_10550);
and U10961 (N_10961,N_10677,N_10682);
nor U10962 (N_10962,N_10663,N_10678);
and U10963 (N_10963,N_10545,N_10576);
or U10964 (N_10964,N_10559,N_10571);
and U10965 (N_10965,N_10596,N_10667);
or U10966 (N_10966,N_10523,N_10688);
or U10967 (N_10967,N_10738,N_10740);
nor U10968 (N_10968,N_10527,N_10627);
and U10969 (N_10969,N_10688,N_10501);
nor U10970 (N_10970,N_10594,N_10509);
and U10971 (N_10971,N_10582,N_10544);
nor U10972 (N_10972,N_10728,N_10518);
or U10973 (N_10973,N_10516,N_10521);
or U10974 (N_10974,N_10616,N_10554);
and U10975 (N_10975,N_10591,N_10628);
nor U10976 (N_10976,N_10559,N_10529);
and U10977 (N_10977,N_10681,N_10716);
nand U10978 (N_10978,N_10721,N_10641);
or U10979 (N_10979,N_10671,N_10686);
xor U10980 (N_10980,N_10622,N_10530);
nand U10981 (N_10981,N_10598,N_10673);
nand U10982 (N_10982,N_10659,N_10506);
and U10983 (N_10983,N_10553,N_10521);
xor U10984 (N_10984,N_10595,N_10737);
nand U10985 (N_10985,N_10590,N_10712);
nand U10986 (N_10986,N_10540,N_10661);
nand U10987 (N_10987,N_10719,N_10581);
nand U10988 (N_10988,N_10529,N_10676);
nor U10989 (N_10989,N_10558,N_10552);
and U10990 (N_10990,N_10568,N_10648);
xnor U10991 (N_10991,N_10636,N_10505);
or U10992 (N_10992,N_10727,N_10501);
and U10993 (N_10993,N_10603,N_10537);
xor U10994 (N_10994,N_10565,N_10598);
and U10995 (N_10995,N_10606,N_10628);
nor U10996 (N_10996,N_10641,N_10551);
xor U10997 (N_10997,N_10727,N_10732);
and U10998 (N_10998,N_10697,N_10519);
and U10999 (N_10999,N_10674,N_10625);
nor U11000 (N_11000,N_10973,N_10986);
and U11001 (N_11001,N_10879,N_10815);
and U11002 (N_11002,N_10849,N_10866);
xor U11003 (N_11003,N_10772,N_10756);
and U11004 (N_11004,N_10942,N_10854);
xor U11005 (N_11005,N_10867,N_10775);
or U11006 (N_11006,N_10933,N_10840);
nand U11007 (N_11007,N_10856,N_10813);
nor U11008 (N_11008,N_10770,N_10972);
nand U11009 (N_11009,N_10932,N_10871);
xnor U11010 (N_11010,N_10801,N_10807);
or U11011 (N_11011,N_10994,N_10918);
nor U11012 (N_11012,N_10948,N_10841);
nand U11013 (N_11013,N_10914,N_10851);
nor U11014 (N_11014,N_10889,N_10799);
nand U11015 (N_11015,N_10999,N_10901);
nor U11016 (N_11016,N_10830,N_10824);
or U11017 (N_11017,N_10868,N_10876);
nand U11018 (N_11018,N_10892,N_10922);
or U11019 (N_11019,N_10752,N_10896);
or U11020 (N_11020,N_10795,N_10891);
and U11021 (N_11021,N_10898,N_10760);
nand U11022 (N_11022,N_10822,N_10971);
xor U11023 (N_11023,N_10959,N_10771);
nand U11024 (N_11024,N_10991,N_10833);
nand U11025 (N_11025,N_10863,N_10951);
or U11026 (N_11026,N_10827,N_10938);
nand U11027 (N_11027,N_10970,N_10888);
nor U11028 (N_11028,N_10817,N_10913);
xnor U11029 (N_11029,N_10819,N_10870);
and U11030 (N_11030,N_10777,N_10809);
and U11031 (N_11031,N_10875,N_10964);
or U11032 (N_11032,N_10821,N_10916);
xor U11033 (N_11033,N_10763,N_10757);
nand U11034 (N_11034,N_10769,N_10784);
nand U11035 (N_11035,N_10865,N_10845);
and U11036 (N_11036,N_10900,N_10953);
xor U11037 (N_11037,N_10930,N_10869);
nor U11038 (N_11038,N_10931,N_10982);
and U11039 (N_11039,N_10993,N_10855);
xor U11040 (N_11040,N_10890,N_10820);
or U11041 (N_11041,N_10759,N_10909);
xnor U11042 (N_11042,N_10980,N_10995);
or U11043 (N_11043,N_10793,N_10786);
xor U11044 (N_11044,N_10794,N_10887);
nor U11045 (N_11045,N_10996,N_10903);
nand U11046 (N_11046,N_10975,N_10850);
xnor U11047 (N_11047,N_10810,N_10842);
and U11048 (N_11048,N_10804,N_10874);
xnor U11049 (N_11049,N_10968,N_10751);
or U11050 (N_11050,N_10788,N_10773);
nor U11051 (N_11051,N_10829,N_10967);
nor U11052 (N_11052,N_10792,N_10977);
or U11053 (N_11053,N_10803,N_10861);
or U11054 (N_11054,N_10997,N_10877);
nand U11055 (N_11055,N_10782,N_10956);
or U11056 (N_11056,N_10910,N_10945);
xnor U11057 (N_11057,N_10939,N_10998);
xor U11058 (N_11058,N_10755,N_10765);
and U11059 (N_11059,N_10785,N_10783);
nand U11060 (N_11060,N_10912,N_10862);
xnor U11061 (N_11061,N_10844,N_10988);
and U11062 (N_11062,N_10966,N_10990);
nand U11063 (N_11063,N_10992,N_10848);
and U11064 (N_11064,N_10886,N_10872);
nor U11065 (N_11065,N_10979,N_10976);
and U11066 (N_11066,N_10895,N_10963);
and U11067 (N_11067,N_10762,N_10904);
nor U11068 (N_11068,N_10826,N_10983);
and U11069 (N_11069,N_10860,N_10835);
or U11070 (N_11070,N_10882,N_10905);
and U11071 (N_11071,N_10857,N_10936);
nor U11072 (N_11072,N_10960,N_10885);
or U11073 (N_11073,N_10802,N_10899);
or U11074 (N_11074,N_10776,N_10881);
nor U11075 (N_11075,N_10944,N_10915);
and U11076 (N_11076,N_10873,N_10926);
xor U11077 (N_11077,N_10780,N_10781);
nand U11078 (N_11078,N_10923,N_10750);
or U11079 (N_11079,N_10949,N_10934);
or U11080 (N_11080,N_10843,N_10758);
xor U11081 (N_11081,N_10906,N_10836);
nand U11082 (N_11082,N_10768,N_10778);
nor U11083 (N_11083,N_10921,N_10927);
or U11084 (N_11084,N_10911,N_10853);
or U11085 (N_11085,N_10754,N_10985);
nand U11086 (N_11086,N_10950,N_10946);
or U11087 (N_11087,N_10825,N_10834);
xnor U11088 (N_11088,N_10958,N_10796);
xor U11089 (N_11089,N_10954,N_10928);
nand U11090 (N_11090,N_10957,N_10791);
and U11091 (N_11091,N_10761,N_10818);
nand U11092 (N_11092,N_10965,N_10955);
and U11093 (N_11093,N_10907,N_10940);
or U11094 (N_11094,N_10952,N_10947);
and U11095 (N_11095,N_10989,N_10846);
nand U11096 (N_11096,N_10859,N_10779);
or U11097 (N_11097,N_10937,N_10917);
xnor U11098 (N_11098,N_10978,N_10878);
and U11099 (N_11099,N_10766,N_10894);
nand U11100 (N_11100,N_10893,N_10935);
or U11101 (N_11101,N_10831,N_10832);
xor U11102 (N_11102,N_10823,N_10924);
and U11103 (N_11103,N_10838,N_10798);
or U11104 (N_11104,N_10812,N_10897);
nor U11105 (N_11105,N_10961,N_10902);
and U11106 (N_11106,N_10774,N_10974);
nand U11107 (N_11107,N_10987,N_10943);
nor U11108 (N_11108,N_10919,N_10880);
nor U11109 (N_11109,N_10962,N_10789);
nand U11110 (N_11110,N_10814,N_10920);
and U11111 (N_11111,N_10908,N_10929);
or U11112 (N_11112,N_10941,N_10753);
or U11113 (N_11113,N_10800,N_10837);
xnor U11114 (N_11114,N_10816,N_10969);
xnor U11115 (N_11115,N_10828,N_10811);
nand U11116 (N_11116,N_10764,N_10852);
or U11117 (N_11117,N_10858,N_10839);
nand U11118 (N_11118,N_10767,N_10787);
nor U11119 (N_11119,N_10805,N_10884);
or U11120 (N_11120,N_10806,N_10790);
xor U11121 (N_11121,N_10981,N_10984);
xnor U11122 (N_11122,N_10847,N_10797);
or U11123 (N_11123,N_10808,N_10883);
xor U11124 (N_11124,N_10925,N_10864);
or U11125 (N_11125,N_10964,N_10916);
nor U11126 (N_11126,N_10883,N_10974);
nor U11127 (N_11127,N_10972,N_10832);
nor U11128 (N_11128,N_10896,N_10900);
and U11129 (N_11129,N_10830,N_10946);
nor U11130 (N_11130,N_10821,N_10777);
and U11131 (N_11131,N_10898,N_10865);
and U11132 (N_11132,N_10784,N_10983);
xor U11133 (N_11133,N_10939,N_10822);
nand U11134 (N_11134,N_10762,N_10989);
nand U11135 (N_11135,N_10830,N_10948);
or U11136 (N_11136,N_10792,N_10807);
and U11137 (N_11137,N_10943,N_10863);
xor U11138 (N_11138,N_10937,N_10831);
nand U11139 (N_11139,N_10959,N_10923);
and U11140 (N_11140,N_10950,N_10894);
and U11141 (N_11141,N_10876,N_10797);
xor U11142 (N_11142,N_10798,N_10910);
or U11143 (N_11143,N_10810,N_10980);
nor U11144 (N_11144,N_10838,N_10868);
nor U11145 (N_11145,N_10896,N_10919);
nor U11146 (N_11146,N_10962,N_10922);
or U11147 (N_11147,N_10893,N_10766);
xor U11148 (N_11148,N_10861,N_10820);
nor U11149 (N_11149,N_10857,N_10884);
xor U11150 (N_11150,N_10939,N_10930);
and U11151 (N_11151,N_10754,N_10934);
nor U11152 (N_11152,N_10799,N_10753);
or U11153 (N_11153,N_10782,N_10803);
xnor U11154 (N_11154,N_10799,N_10823);
or U11155 (N_11155,N_10843,N_10819);
or U11156 (N_11156,N_10842,N_10933);
nand U11157 (N_11157,N_10764,N_10797);
or U11158 (N_11158,N_10788,N_10847);
and U11159 (N_11159,N_10933,N_10899);
and U11160 (N_11160,N_10754,N_10794);
and U11161 (N_11161,N_10892,N_10951);
nand U11162 (N_11162,N_10870,N_10784);
or U11163 (N_11163,N_10956,N_10905);
and U11164 (N_11164,N_10935,N_10988);
or U11165 (N_11165,N_10946,N_10899);
nand U11166 (N_11166,N_10933,N_10871);
nand U11167 (N_11167,N_10929,N_10981);
and U11168 (N_11168,N_10754,N_10964);
nor U11169 (N_11169,N_10751,N_10831);
nor U11170 (N_11170,N_10847,N_10953);
nand U11171 (N_11171,N_10811,N_10773);
xnor U11172 (N_11172,N_10886,N_10756);
nand U11173 (N_11173,N_10822,N_10922);
and U11174 (N_11174,N_10935,N_10778);
or U11175 (N_11175,N_10962,N_10875);
xnor U11176 (N_11176,N_10945,N_10887);
nand U11177 (N_11177,N_10926,N_10950);
xnor U11178 (N_11178,N_10971,N_10817);
nand U11179 (N_11179,N_10855,N_10807);
xor U11180 (N_11180,N_10989,N_10893);
xor U11181 (N_11181,N_10780,N_10912);
nand U11182 (N_11182,N_10799,N_10858);
xnor U11183 (N_11183,N_10871,N_10987);
nor U11184 (N_11184,N_10780,N_10799);
and U11185 (N_11185,N_10885,N_10855);
nand U11186 (N_11186,N_10787,N_10906);
nand U11187 (N_11187,N_10761,N_10785);
xnor U11188 (N_11188,N_10958,N_10908);
nor U11189 (N_11189,N_10780,N_10963);
or U11190 (N_11190,N_10752,N_10823);
nor U11191 (N_11191,N_10776,N_10782);
and U11192 (N_11192,N_10803,N_10773);
nand U11193 (N_11193,N_10874,N_10887);
or U11194 (N_11194,N_10977,N_10986);
and U11195 (N_11195,N_10860,N_10833);
nand U11196 (N_11196,N_10945,N_10964);
nor U11197 (N_11197,N_10845,N_10778);
or U11198 (N_11198,N_10937,N_10851);
or U11199 (N_11199,N_10763,N_10750);
or U11200 (N_11200,N_10856,N_10976);
nand U11201 (N_11201,N_10816,N_10859);
and U11202 (N_11202,N_10799,N_10804);
and U11203 (N_11203,N_10992,N_10882);
and U11204 (N_11204,N_10895,N_10940);
or U11205 (N_11205,N_10752,N_10824);
nor U11206 (N_11206,N_10946,N_10816);
nor U11207 (N_11207,N_10874,N_10851);
xor U11208 (N_11208,N_10773,N_10750);
nor U11209 (N_11209,N_10897,N_10793);
and U11210 (N_11210,N_10840,N_10978);
xor U11211 (N_11211,N_10837,N_10927);
and U11212 (N_11212,N_10946,N_10953);
nand U11213 (N_11213,N_10913,N_10930);
nor U11214 (N_11214,N_10885,N_10919);
and U11215 (N_11215,N_10982,N_10808);
xnor U11216 (N_11216,N_10852,N_10989);
nor U11217 (N_11217,N_10936,N_10921);
xnor U11218 (N_11218,N_10950,N_10776);
or U11219 (N_11219,N_10898,N_10847);
xor U11220 (N_11220,N_10907,N_10976);
nand U11221 (N_11221,N_10886,N_10956);
nor U11222 (N_11222,N_10825,N_10935);
nor U11223 (N_11223,N_10888,N_10931);
or U11224 (N_11224,N_10817,N_10868);
and U11225 (N_11225,N_10782,N_10888);
nand U11226 (N_11226,N_10823,N_10769);
nand U11227 (N_11227,N_10880,N_10979);
or U11228 (N_11228,N_10761,N_10893);
or U11229 (N_11229,N_10832,N_10788);
and U11230 (N_11230,N_10763,N_10812);
nor U11231 (N_11231,N_10768,N_10942);
nand U11232 (N_11232,N_10981,N_10818);
and U11233 (N_11233,N_10861,N_10907);
nor U11234 (N_11234,N_10996,N_10780);
nand U11235 (N_11235,N_10796,N_10931);
or U11236 (N_11236,N_10763,N_10878);
xnor U11237 (N_11237,N_10875,N_10928);
or U11238 (N_11238,N_10927,N_10843);
nand U11239 (N_11239,N_10754,N_10759);
and U11240 (N_11240,N_10984,N_10975);
nor U11241 (N_11241,N_10787,N_10922);
nand U11242 (N_11242,N_10766,N_10768);
and U11243 (N_11243,N_10960,N_10917);
nand U11244 (N_11244,N_10940,N_10839);
nand U11245 (N_11245,N_10889,N_10883);
nand U11246 (N_11246,N_10877,N_10930);
or U11247 (N_11247,N_10865,N_10986);
nor U11248 (N_11248,N_10810,N_10903);
and U11249 (N_11249,N_10965,N_10807);
nand U11250 (N_11250,N_11062,N_11127);
or U11251 (N_11251,N_11143,N_11113);
xnor U11252 (N_11252,N_11164,N_11119);
or U11253 (N_11253,N_11128,N_11003);
or U11254 (N_11254,N_11080,N_11189);
xnor U11255 (N_11255,N_11101,N_11055);
nand U11256 (N_11256,N_11138,N_11031);
nand U11257 (N_11257,N_11249,N_11060);
and U11258 (N_11258,N_11122,N_11118);
xor U11259 (N_11259,N_11232,N_11084);
nor U11260 (N_11260,N_11206,N_11099);
xor U11261 (N_11261,N_11009,N_11241);
nor U11262 (N_11262,N_11216,N_11220);
or U11263 (N_11263,N_11109,N_11131);
nand U11264 (N_11264,N_11058,N_11212);
or U11265 (N_11265,N_11204,N_11098);
nand U11266 (N_11266,N_11090,N_11202);
nand U11267 (N_11267,N_11108,N_11100);
nor U11268 (N_11268,N_11208,N_11116);
xnor U11269 (N_11269,N_11183,N_11225);
nor U11270 (N_11270,N_11175,N_11048);
and U11271 (N_11271,N_11078,N_11089);
nor U11272 (N_11272,N_11016,N_11196);
or U11273 (N_11273,N_11137,N_11247);
nor U11274 (N_11274,N_11026,N_11178);
nor U11275 (N_11275,N_11068,N_11197);
nand U11276 (N_11276,N_11152,N_11168);
nor U11277 (N_11277,N_11029,N_11157);
and U11278 (N_11278,N_11171,N_11222);
or U11279 (N_11279,N_11240,N_11075);
nand U11280 (N_11280,N_11043,N_11007);
or U11281 (N_11281,N_11107,N_11000);
xor U11282 (N_11282,N_11161,N_11184);
or U11283 (N_11283,N_11018,N_11226);
and U11284 (N_11284,N_11010,N_11181);
nand U11285 (N_11285,N_11150,N_11190);
or U11286 (N_11286,N_11085,N_11053);
xnor U11287 (N_11287,N_11012,N_11063);
and U11288 (N_11288,N_11038,N_11231);
nand U11289 (N_11289,N_11230,N_11141);
nand U11290 (N_11290,N_11054,N_11027);
xor U11291 (N_11291,N_11059,N_11154);
or U11292 (N_11292,N_11242,N_11174);
nor U11293 (N_11293,N_11142,N_11153);
or U11294 (N_11294,N_11163,N_11248);
and U11295 (N_11295,N_11229,N_11151);
nor U11296 (N_11296,N_11082,N_11166);
or U11297 (N_11297,N_11004,N_11037);
xnor U11298 (N_11298,N_11134,N_11083);
nand U11299 (N_11299,N_11147,N_11030);
nand U11300 (N_11300,N_11073,N_11176);
and U11301 (N_11301,N_11050,N_11072);
nand U11302 (N_11302,N_11041,N_11077);
nand U11303 (N_11303,N_11104,N_11001);
nor U11304 (N_11304,N_11102,N_11211);
nand U11305 (N_11305,N_11180,N_11092);
nand U11306 (N_11306,N_11071,N_11214);
nand U11307 (N_11307,N_11021,N_11065);
and U11308 (N_11308,N_11091,N_11020);
nand U11309 (N_11309,N_11132,N_11115);
or U11310 (N_11310,N_11195,N_11097);
or U11311 (N_11311,N_11246,N_11056);
and U11312 (N_11312,N_11042,N_11193);
and U11313 (N_11313,N_11133,N_11033);
nor U11314 (N_11314,N_11219,N_11201);
or U11315 (N_11315,N_11014,N_11044);
and U11316 (N_11316,N_11106,N_11187);
nor U11317 (N_11317,N_11112,N_11243);
nand U11318 (N_11318,N_11117,N_11129);
nor U11319 (N_11319,N_11136,N_11076);
nand U11320 (N_11320,N_11093,N_11172);
and U11321 (N_11321,N_11067,N_11040);
xor U11322 (N_11322,N_11169,N_11130);
or U11323 (N_11323,N_11158,N_11160);
nor U11324 (N_11324,N_11177,N_11124);
nor U11325 (N_11325,N_11203,N_11199);
nor U11326 (N_11326,N_11025,N_11019);
or U11327 (N_11327,N_11022,N_11188);
and U11328 (N_11328,N_11061,N_11051);
nand U11329 (N_11329,N_11224,N_11221);
or U11330 (N_11330,N_11244,N_11148);
or U11331 (N_11331,N_11049,N_11064);
xor U11332 (N_11332,N_11167,N_11145);
nand U11333 (N_11333,N_11209,N_11005);
and U11334 (N_11334,N_11032,N_11095);
nor U11335 (N_11335,N_11235,N_11213);
nand U11336 (N_11336,N_11165,N_11023);
nand U11337 (N_11337,N_11173,N_11227);
or U11338 (N_11338,N_11123,N_11046);
and U11339 (N_11339,N_11002,N_11149);
nor U11340 (N_11340,N_11139,N_11179);
nand U11341 (N_11341,N_11207,N_11081);
nor U11342 (N_11342,N_11006,N_11146);
or U11343 (N_11343,N_11015,N_11036);
and U11344 (N_11344,N_11215,N_11237);
and U11345 (N_11345,N_11086,N_11170);
and U11346 (N_11346,N_11191,N_11200);
nand U11347 (N_11347,N_11135,N_11047);
and U11348 (N_11348,N_11114,N_11234);
and U11349 (N_11349,N_11217,N_11070);
nor U11350 (N_11350,N_11186,N_11011);
or U11351 (N_11351,N_11144,N_11198);
and U11352 (N_11352,N_11024,N_11126);
xor U11353 (N_11353,N_11228,N_11121);
and U11354 (N_11354,N_11120,N_11087);
or U11355 (N_11355,N_11039,N_11192);
or U11356 (N_11356,N_11103,N_11105);
nor U11357 (N_11357,N_11218,N_11094);
nor U11358 (N_11358,N_11156,N_11140);
or U11359 (N_11359,N_11223,N_11088);
nor U11360 (N_11360,N_11013,N_11110);
and U11361 (N_11361,N_11236,N_11245);
or U11362 (N_11362,N_11162,N_11017);
xnor U11363 (N_11363,N_11205,N_11034);
nor U11364 (N_11364,N_11066,N_11079);
xnor U11365 (N_11365,N_11074,N_11008);
and U11366 (N_11366,N_11035,N_11238);
and U11367 (N_11367,N_11028,N_11233);
or U11368 (N_11368,N_11194,N_11239);
nand U11369 (N_11369,N_11045,N_11182);
and U11370 (N_11370,N_11125,N_11069);
xnor U11371 (N_11371,N_11052,N_11210);
xnor U11372 (N_11372,N_11096,N_11155);
xnor U11373 (N_11373,N_11159,N_11057);
nand U11374 (N_11374,N_11185,N_11111);
nor U11375 (N_11375,N_11121,N_11199);
nand U11376 (N_11376,N_11094,N_11005);
or U11377 (N_11377,N_11047,N_11166);
nand U11378 (N_11378,N_11050,N_11030);
nor U11379 (N_11379,N_11140,N_11243);
xnor U11380 (N_11380,N_11040,N_11034);
xnor U11381 (N_11381,N_11192,N_11196);
xnor U11382 (N_11382,N_11099,N_11081);
and U11383 (N_11383,N_11164,N_11045);
and U11384 (N_11384,N_11084,N_11019);
xor U11385 (N_11385,N_11057,N_11109);
nand U11386 (N_11386,N_11089,N_11038);
xnor U11387 (N_11387,N_11138,N_11191);
or U11388 (N_11388,N_11161,N_11063);
or U11389 (N_11389,N_11152,N_11140);
and U11390 (N_11390,N_11131,N_11197);
and U11391 (N_11391,N_11154,N_11212);
xor U11392 (N_11392,N_11058,N_11119);
or U11393 (N_11393,N_11112,N_11230);
nand U11394 (N_11394,N_11151,N_11027);
and U11395 (N_11395,N_11000,N_11167);
nand U11396 (N_11396,N_11171,N_11132);
and U11397 (N_11397,N_11229,N_11211);
nand U11398 (N_11398,N_11020,N_11139);
or U11399 (N_11399,N_11136,N_11204);
or U11400 (N_11400,N_11203,N_11195);
nand U11401 (N_11401,N_11222,N_11185);
and U11402 (N_11402,N_11137,N_11131);
xnor U11403 (N_11403,N_11170,N_11128);
or U11404 (N_11404,N_11131,N_11208);
nor U11405 (N_11405,N_11183,N_11238);
xnor U11406 (N_11406,N_11126,N_11099);
or U11407 (N_11407,N_11065,N_11196);
nand U11408 (N_11408,N_11139,N_11226);
xor U11409 (N_11409,N_11049,N_11192);
xor U11410 (N_11410,N_11088,N_11069);
or U11411 (N_11411,N_11185,N_11003);
nand U11412 (N_11412,N_11131,N_11082);
nor U11413 (N_11413,N_11038,N_11130);
xor U11414 (N_11414,N_11217,N_11139);
nor U11415 (N_11415,N_11103,N_11038);
or U11416 (N_11416,N_11192,N_11040);
xor U11417 (N_11417,N_11028,N_11137);
and U11418 (N_11418,N_11177,N_11226);
nand U11419 (N_11419,N_11188,N_11087);
nand U11420 (N_11420,N_11149,N_11239);
nand U11421 (N_11421,N_11108,N_11220);
nand U11422 (N_11422,N_11005,N_11129);
nand U11423 (N_11423,N_11165,N_11249);
nand U11424 (N_11424,N_11151,N_11163);
xor U11425 (N_11425,N_11215,N_11168);
nand U11426 (N_11426,N_11134,N_11201);
or U11427 (N_11427,N_11085,N_11123);
and U11428 (N_11428,N_11164,N_11160);
nor U11429 (N_11429,N_11242,N_11169);
xnor U11430 (N_11430,N_11144,N_11063);
nor U11431 (N_11431,N_11150,N_11092);
and U11432 (N_11432,N_11030,N_11003);
xnor U11433 (N_11433,N_11152,N_11225);
and U11434 (N_11434,N_11165,N_11114);
nand U11435 (N_11435,N_11023,N_11232);
nand U11436 (N_11436,N_11227,N_11168);
nand U11437 (N_11437,N_11123,N_11020);
and U11438 (N_11438,N_11116,N_11022);
xnor U11439 (N_11439,N_11004,N_11182);
xnor U11440 (N_11440,N_11130,N_11006);
and U11441 (N_11441,N_11049,N_11044);
nand U11442 (N_11442,N_11233,N_11142);
nand U11443 (N_11443,N_11203,N_11070);
and U11444 (N_11444,N_11215,N_11177);
or U11445 (N_11445,N_11018,N_11032);
xor U11446 (N_11446,N_11165,N_11094);
or U11447 (N_11447,N_11234,N_11021);
and U11448 (N_11448,N_11032,N_11078);
nor U11449 (N_11449,N_11106,N_11239);
nor U11450 (N_11450,N_11241,N_11226);
or U11451 (N_11451,N_11045,N_11040);
or U11452 (N_11452,N_11152,N_11105);
or U11453 (N_11453,N_11045,N_11025);
nor U11454 (N_11454,N_11049,N_11006);
nor U11455 (N_11455,N_11158,N_11203);
or U11456 (N_11456,N_11223,N_11040);
and U11457 (N_11457,N_11153,N_11193);
nor U11458 (N_11458,N_11197,N_11233);
and U11459 (N_11459,N_11160,N_11203);
and U11460 (N_11460,N_11115,N_11123);
or U11461 (N_11461,N_11169,N_11097);
nand U11462 (N_11462,N_11136,N_11027);
nand U11463 (N_11463,N_11141,N_11024);
nor U11464 (N_11464,N_11007,N_11179);
nor U11465 (N_11465,N_11071,N_11141);
nor U11466 (N_11466,N_11100,N_11014);
and U11467 (N_11467,N_11096,N_11078);
nand U11468 (N_11468,N_11173,N_11167);
nand U11469 (N_11469,N_11177,N_11135);
or U11470 (N_11470,N_11014,N_11138);
nand U11471 (N_11471,N_11194,N_11151);
nor U11472 (N_11472,N_11179,N_11108);
or U11473 (N_11473,N_11177,N_11028);
nand U11474 (N_11474,N_11001,N_11137);
nor U11475 (N_11475,N_11142,N_11027);
nand U11476 (N_11476,N_11009,N_11197);
xor U11477 (N_11477,N_11191,N_11127);
or U11478 (N_11478,N_11040,N_11216);
and U11479 (N_11479,N_11053,N_11038);
nor U11480 (N_11480,N_11126,N_11113);
xor U11481 (N_11481,N_11067,N_11151);
or U11482 (N_11482,N_11201,N_11156);
xor U11483 (N_11483,N_11069,N_11215);
nor U11484 (N_11484,N_11080,N_11078);
nor U11485 (N_11485,N_11133,N_11142);
nor U11486 (N_11486,N_11021,N_11038);
xnor U11487 (N_11487,N_11217,N_11117);
or U11488 (N_11488,N_11189,N_11245);
nand U11489 (N_11489,N_11105,N_11230);
nand U11490 (N_11490,N_11126,N_11175);
nor U11491 (N_11491,N_11098,N_11035);
nor U11492 (N_11492,N_11075,N_11155);
and U11493 (N_11493,N_11101,N_11004);
nor U11494 (N_11494,N_11180,N_11059);
xnor U11495 (N_11495,N_11238,N_11071);
or U11496 (N_11496,N_11002,N_11198);
nand U11497 (N_11497,N_11003,N_11231);
and U11498 (N_11498,N_11170,N_11027);
or U11499 (N_11499,N_11218,N_11040);
nand U11500 (N_11500,N_11471,N_11392);
or U11501 (N_11501,N_11368,N_11383);
nand U11502 (N_11502,N_11488,N_11266);
nor U11503 (N_11503,N_11341,N_11258);
xor U11504 (N_11504,N_11410,N_11444);
nor U11505 (N_11505,N_11291,N_11298);
and U11506 (N_11506,N_11374,N_11295);
or U11507 (N_11507,N_11492,N_11478);
nor U11508 (N_11508,N_11311,N_11423);
xor U11509 (N_11509,N_11303,N_11393);
nor U11510 (N_11510,N_11281,N_11468);
nor U11511 (N_11511,N_11402,N_11387);
nand U11512 (N_11512,N_11270,N_11405);
or U11513 (N_11513,N_11339,N_11260);
nor U11514 (N_11514,N_11411,N_11255);
or U11515 (N_11515,N_11359,N_11494);
nor U11516 (N_11516,N_11330,N_11479);
or U11517 (N_11517,N_11332,N_11475);
nand U11518 (N_11518,N_11490,N_11307);
xnor U11519 (N_11519,N_11347,N_11484);
and U11520 (N_11520,N_11304,N_11456);
nand U11521 (N_11521,N_11319,N_11296);
xnor U11522 (N_11522,N_11459,N_11434);
nor U11523 (N_11523,N_11465,N_11324);
nor U11524 (N_11524,N_11289,N_11406);
xor U11525 (N_11525,N_11353,N_11476);
or U11526 (N_11526,N_11428,N_11425);
nor U11527 (N_11527,N_11299,N_11499);
or U11528 (N_11528,N_11466,N_11433);
nor U11529 (N_11529,N_11297,N_11305);
and U11530 (N_11530,N_11306,N_11278);
xor U11531 (N_11531,N_11349,N_11293);
nor U11532 (N_11532,N_11446,N_11421);
nand U11533 (N_11533,N_11390,N_11438);
xnor U11534 (N_11534,N_11254,N_11321);
xnor U11535 (N_11535,N_11315,N_11395);
nand U11536 (N_11536,N_11461,N_11382);
and U11537 (N_11537,N_11400,N_11338);
xnor U11538 (N_11538,N_11313,N_11399);
nor U11539 (N_11539,N_11489,N_11337);
and U11540 (N_11540,N_11285,N_11407);
or U11541 (N_11541,N_11263,N_11449);
or U11542 (N_11542,N_11371,N_11389);
nor U11543 (N_11543,N_11327,N_11415);
nor U11544 (N_11544,N_11323,N_11498);
nand U11545 (N_11545,N_11472,N_11427);
xor U11546 (N_11546,N_11437,N_11442);
or U11547 (N_11547,N_11398,N_11381);
or U11548 (N_11548,N_11300,N_11355);
or U11549 (N_11549,N_11350,N_11362);
nand U11550 (N_11550,N_11346,N_11443);
or U11551 (N_11551,N_11403,N_11343);
or U11552 (N_11552,N_11336,N_11414);
xnor U11553 (N_11553,N_11474,N_11329);
nor U11554 (N_11554,N_11409,N_11301);
and U11555 (N_11555,N_11317,N_11252);
xor U11556 (N_11556,N_11372,N_11376);
nand U11557 (N_11557,N_11309,N_11441);
and U11558 (N_11558,N_11396,N_11432);
and U11559 (N_11559,N_11451,N_11377);
nand U11560 (N_11560,N_11369,N_11375);
nor U11561 (N_11561,N_11480,N_11334);
xor U11562 (N_11562,N_11276,N_11360);
and U11563 (N_11563,N_11325,N_11250);
nand U11564 (N_11564,N_11470,N_11271);
and U11565 (N_11565,N_11496,N_11275);
nor U11566 (N_11566,N_11386,N_11431);
nor U11567 (N_11567,N_11458,N_11257);
or U11568 (N_11568,N_11380,N_11314);
nand U11569 (N_11569,N_11436,N_11284);
and U11570 (N_11570,N_11331,N_11420);
and U11571 (N_11571,N_11342,N_11286);
xor U11572 (N_11572,N_11455,N_11473);
or U11573 (N_11573,N_11495,N_11356);
xor U11574 (N_11574,N_11357,N_11429);
xnor U11575 (N_11575,N_11435,N_11460);
and U11576 (N_11576,N_11316,N_11401);
nor U11577 (N_11577,N_11354,N_11477);
or U11578 (N_11578,N_11417,N_11290);
and U11579 (N_11579,N_11312,N_11345);
xor U11580 (N_11580,N_11486,N_11283);
and U11581 (N_11581,N_11485,N_11450);
or U11582 (N_11582,N_11373,N_11365);
nor U11583 (N_11583,N_11256,N_11262);
nand U11584 (N_11584,N_11378,N_11408);
nor U11585 (N_11585,N_11367,N_11388);
nor U11586 (N_11586,N_11364,N_11320);
and U11587 (N_11587,N_11482,N_11413);
nand U11588 (N_11588,N_11481,N_11292);
xnor U11589 (N_11589,N_11335,N_11322);
and U11590 (N_11590,N_11440,N_11430);
or U11591 (N_11591,N_11261,N_11394);
and U11592 (N_11592,N_11497,N_11267);
or U11593 (N_11593,N_11363,N_11272);
nand U11594 (N_11594,N_11351,N_11328);
nand U11595 (N_11595,N_11391,N_11462);
nor U11596 (N_11596,N_11467,N_11302);
xor U11597 (N_11597,N_11253,N_11422);
nand U11598 (N_11598,N_11348,N_11352);
or U11599 (N_11599,N_11274,N_11344);
xnor U11600 (N_11600,N_11279,N_11318);
xnor U11601 (N_11601,N_11419,N_11277);
or U11602 (N_11602,N_11404,N_11308);
or U11603 (N_11603,N_11447,N_11259);
nand U11604 (N_11604,N_11483,N_11264);
nor U11605 (N_11605,N_11361,N_11491);
xnor U11606 (N_11606,N_11418,N_11333);
nand U11607 (N_11607,N_11469,N_11454);
nor U11608 (N_11608,N_11453,N_11439);
xor U11609 (N_11609,N_11269,N_11370);
and U11610 (N_11610,N_11397,N_11412);
and U11611 (N_11611,N_11379,N_11457);
nand U11612 (N_11612,N_11448,N_11384);
and U11613 (N_11613,N_11385,N_11251);
nand U11614 (N_11614,N_11445,N_11282);
or U11615 (N_11615,N_11416,N_11452);
nor U11616 (N_11616,N_11426,N_11463);
or U11617 (N_11617,N_11493,N_11358);
nor U11618 (N_11618,N_11464,N_11366);
nor U11619 (N_11619,N_11273,N_11280);
nor U11620 (N_11620,N_11340,N_11310);
nand U11621 (N_11621,N_11294,N_11268);
nand U11622 (N_11622,N_11265,N_11487);
and U11623 (N_11623,N_11424,N_11288);
nor U11624 (N_11624,N_11326,N_11287);
nand U11625 (N_11625,N_11365,N_11417);
and U11626 (N_11626,N_11391,N_11449);
and U11627 (N_11627,N_11471,N_11433);
xor U11628 (N_11628,N_11313,N_11489);
nor U11629 (N_11629,N_11342,N_11282);
xor U11630 (N_11630,N_11437,N_11272);
and U11631 (N_11631,N_11409,N_11481);
nand U11632 (N_11632,N_11394,N_11302);
xnor U11633 (N_11633,N_11406,N_11365);
nand U11634 (N_11634,N_11308,N_11414);
and U11635 (N_11635,N_11370,N_11407);
or U11636 (N_11636,N_11334,N_11375);
xor U11637 (N_11637,N_11315,N_11328);
xnor U11638 (N_11638,N_11355,N_11365);
nor U11639 (N_11639,N_11484,N_11325);
nand U11640 (N_11640,N_11424,N_11412);
nand U11641 (N_11641,N_11256,N_11270);
xnor U11642 (N_11642,N_11335,N_11491);
or U11643 (N_11643,N_11281,N_11385);
nor U11644 (N_11644,N_11317,N_11432);
or U11645 (N_11645,N_11273,N_11477);
nand U11646 (N_11646,N_11440,N_11309);
xor U11647 (N_11647,N_11365,N_11449);
and U11648 (N_11648,N_11370,N_11343);
and U11649 (N_11649,N_11299,N_11283);
and U11650 (N_11650,N_11390,N_11310);
xnor U11651 (N_11651,N_11256,N_11365);
or U11652 (N_11652,N_11388,N_11260);
xor U11653 (N_11653,N_11344,N_11484);
nand U11654 (N_11654,N_11324,N_11398);
nor U11655 (N_11655,N_11367,N_11306);
or U11656 (N_11656,N_11255,N_11272);
nor U11657 (N_11657,N_11348,N_11252);
xor U11658 (N_11658,N_11254,N_11455);
nand U11659 (N_11659,N_11399,N_11479);
and U11660 (N_11660,N_11363,N_11256);
nand U11661 (N_11661,N_11377,N_11417);
nor U11662 (N_11662,N_11480,N_11443);
xor U11663 (N_11663,N_11302,N_11419);
nor U11664 (N_11664,N_11433,N_11283);
xnor U11665 (N_11665,N_11419,N_11259);
nor U11666 (N_11666,N_11289,N_11327);
nor U11667 (N_11667,N_11468,N_11414);
xnor U11668 (N_11668,N_11410,N_11474);
and U11669 (N_11669,N_11386,N_11424);
nor U11670 (N_11670,N_11444,N_11446);
and U11671 (N_11671,N_11294,N_11281);
nand U11672 (N_11672,N_11463,N_11440);
xnor U11673 (N_11673,N_11372,N_11380);
nor U11674 (N_11674,N_11359,N_11484);
and U11675 (N_11675,N_11451,N_11257);
and U11676 (N_11676,N_11413,N_11320);
xor U11677 (N_11677,N_11335,N_11332);
nand U11678 (N_11678,N_11379,N_11464);
and U11679 (N_11679,N_11360,N_11395);
nand U11680 (N_11680,N_11338,N_11415);
xor U11681 (N_11681,N_11444,N_11356);
xor U11682 (N_11682,N_11298,N_11302);
nand U11683 (N_11683,N_11398,N_11315);
xor U11684 (N_11684,N_11404,N_11273);
nand U11685 (N_11685,N_11319,N_11359);
nand U11686 (N_11686,N_11487,N_11365);
or U11687 (N_11687,N_11489,N_11475);
and U11688 (N_11688,N_11473,N_11470);
and U11689 (N_11689,N_11463,N_11280);
nor U11690 (N_11690,N_11309,N_11394);
xnor U11691 (N_11691,N_11471,N_11418);
nand U11692 (N_11692,N_11440,N_11377);
and U11693 (N_11693,N_11484,N_11413);
nand U11694 (N_11694,N_11444,N_11311);
and U11695 (N_11695,N_11343,N_11351);
and U11696 (N_11696,N_11368,N_11381);
nand U11697 (N_11697,N_11329,N_11468);
nor U11698 (N_11698,N_11424,N_11398);
nor U11699 (N_11699,N_11494,N_11349);
and U11700 (N_11700,N_11370,N_11285);
and U11701 (N_11701,N_11475,N_11409);
or U11702 (N_11702,N_11278,N_11417);
or U11703 (N_11703,N_11469,N_11359);
and U11704 (N_11704,N_11261,N_11250);
or U11705 (N_11705,N_11446,N_11479);
nand U11706 (N_11706,N_11266,N_11470);
nand U11707 (N_11707,N_11452,N_11393);
or U11708 (N_11708,N_11379,N_11371);
xnor U11709 (N_11709,N_11308,N_11498);
nand U11710 (N_11710,N_11487,N_11319);
or U11711 (N_11711,N_11331,N_11266);
and U11712 (N_11712,N_11357,N_11330);
xnor U11713 (N_11713,N_11444,N_11272);
nor U11714 (N_11714,N_11261,N_11428);
nor U11715 (N_11715,N_11474,N_11337);
nor U11716 (N_11716,N_11345,N_11265);
xor U11717 (N_11717,N_11363,N_11361);
and U11718 (N_11718,N_11281,N_11337);
xnor U11719 (N_11719,N_11360,N_11469);
nor U11720 (N_11720,N_11392,N_11307);
or U11721 (N_11721,N_11420,N_11270);
xor U11722 (N_11722,N_11414,N_11470);
nand U11723 (N_11723,N_11412,N_11468);
nor U11724 (N_11724,N_11453,N_11390);
nand U11725 (N_11725,N_11399,N_11429);
nand U11726 (N_11726,N_11410,N_11252);
or U11727 (N_11727,N_11319,N_11304);
or U11728 (N_11728,N_11258,N_11464);
and U11729 (N_11729,N_11432,N_11290);
xor U11730 (N_11730,N_11330,N_11470);
nor U11731 (N_11731,N_11391,N_11289);
nand U11732 (N_11732,N_11436,N_11398);
nor U11733 (N_11733,N_11270,N_11393);
nor U11734 (N_11734,N_11386,N_11250);
nor U11735 (N_11735,N_11455,N_11272);
nor U11736 (N_11736,N_11292,N_11328);
nor U11737 (N_11737,N_11342,N_11252);
and U11738 (N_11738,N_11402,N_11385);
nand U11739 (N_11739,N_11409,N_11369);
or U11740 (N_11740,N_11465,N_11489);
nor U11741 (N_11741,N_11327,N_11296);
and U11742 (N_11742,N_11314,N_11253);
nor U11743 (N_11743,N_11305,N_11322);
xor U11744 (N_11744,N_11383,N_11330);
and U11745 (N_11745,N_11255,N_11458);
nand U11746 (N_11746,N_11348,N_11455);
nand U11747 (N_11747,N_11274,N_11357);
or U11748 (N_11748,N_11263,N_11442);
nor U11749 (N_11749,N_11320,N_11417);
xnor U11750 (N_11750,N_11548,N_11722);
or U11751 (N_11751,N_11745,N_11523);
nor U11752 (N_11752,N_11688,N_11730);
or U11753 (N_11753,N_11710,N_11698);
nand U11754 (N_11754,N_11708,N_11669);
xor U11755 (N_11755,N_11566,N_11540);
nor U11756 (N_11756,N_11551,N_11646);
or U11757 (N_11757,N_11629,N_11623);
xor U11758 (N_11758,N_11524,N_11601);
or U11759 (N_11759,N_11676,N_11563);
xor U11760 (N_11760,N_11565,N_11530);
nand U11761 (N_11761,N_11561,N_11593);
nand U11762 (N_11762,N_11699,N_11596);
nor U11763 (N_11763,N_11554,N_11539);
and U11764 (N_11764,N_11543,N_11624);
nor U11765 (N_11765,N_11740,N_11610);
and U11766 (N_11766,N_11590,N_11679);
nand U11767 (N_11767,N_11545,N_11580);
nor U11768 (N_11768,N_11536,N_11707);
xnor U11769 (N_11769,N_11528,N_11559);
nand U11770 (N_11770,N_11547,N_11725);
and U11771 (N_11771,N_11518,N_11643);
or U11772 (N_11772,N_11746,N_11668);
nand U11773 (N_11773,N_11644,N_11597);
nor U11774 (N_11774,N_11682,N_11656);
or U11775 (N_11775,N_11739,N_11504);
xnor U11776 (N_11776,N_11572,N_11742);
xnor U11777 (N_11777,N_11599,N_11744);
nor U11778 (N_11778,N_11655,N_11639);
or U11779 (N_11779,N_11712,N_11615);
nand U11780 (N_11780,N_11532,N_11684);
nor U11781 (N_11781,N_11625,N_11607);
nand U11782 (N_11782,N_11716,N_11697);
nand U11783 (N_11783,N_11603,N_11595);
xor U11784 (N_11784,N_11531,N_11560);
and U11785 (N_11785,N_11631,N_11529);
nor U11786 (N_11786,N_11736,N_11741);
xnor U11787 (N_11787,N_11588,N_11609);
or U11788 (N_11788,N_11534,N_11672);
nand U11789 (N_11789,N_11585,N_11748);
or U11790 (N_11790,N_11706,N_11608);
xor U11791 (N_11791,N_11632,N_11680);
nand U11792 (N_11792,N_11501,N_11509);
xor U11793 (N_11793,N_11577,N_11503);
xor U11794 (N_11794,N_11723,N_11506);
xor U11795 (N_11795,N_11541,N_11605);
nand U11796 (N_11796,N_11692,N_11579);
and U11797 (N_11797,N_11521,N_11726);
xor U11798 (N_11798,N_11512,N_11515);
or U11799 (N_11799,N_11641,N_11729);
nor U11800 (N_11800,N_11696,N_11606);
xor U11801 (N_11801,N_11634,N_11568);
xnor U11802 (N_11802,N_11627,N_11620);
nand U11803 (N_11803,N_11738,N_11701);
nand U11804 (N_11804,N_11535,N_11616);
or U11805 (N_11805,N_11619,N_11573);
nor U11806 (N_11806,N_11686,N_11645);
nand U11807 (N_11807,N_11558,N_11553);
and U11808 (N_11808,N_11584,N_11678);
xor U11809 (N_11809,N_11648,N_11600);
nor U11810 (N_11810,N_11613,N_11693);
or U11811 (N_11811,N_11576,N_11526);
xor U11812 (N_11812,N_11651,N_11510);
and U11813 (N_11813,N_11626,N_11652);
nor U11814 (N_11814,N_11511,N_11578);
nand U11815 (N_11815,N_11592,N_11611);
and U11816 (N_11816,N_11647,N_11552);
xnor U11817 (N_11817,N_11617,N_11614);
nand U11818 (N_11818,N_11516,N_11546);
xnor U11819 (N_11819,N_11747,N_11618);
nor U11820 (N_11820,N_11500,N_11653);
xor U11821 (N_11821,N_11520,N_11636);
or U11822 (N_11822,N_11743,N_11542);
nand U11823 (N_11823,N_11658,N_11640);
xnor U11824 (N_11824,N_11550,N_11670);
or U11825 (N_11825,N_11695,N_11721);
and U11826 (N_11826,N_11628,N_11677);
nor U11827 (N_11827,N_11522,N_11727);
nor U11828 (N_11828,N_11527,N_11513);
xor U11829 (N_11829,N_11519,N_11734);
nor U11830 (N_11830,N_11717,N_11557);
and U11831 (N_11831,N_11703,N_11583);
xnor U11832 (N_11832,N_11538,N_11673);
nor U11833 (N_11833,N_11714,N_11728);
xnor U11834 (N_11834,N_11570,N_11638);
nand U11835 (N_11835,N_11683,N_11662);
and U11836 (N_11836,N_11675,N_11689);
nand U11837 (N_11837,N_11574,N_11581);
nor U11838 (N_11838,N_11718,N_11749);
or U11839 (N_11839,N_11544,N_11681);
or U11840 (N_11840,N_11690,N_11582);
or U11841 (N_11841,N_11713,N_11671);
nor U11842 (N_11842,N_11642,N_11587);
nor U11843 (N_11843,N_11514,N_11517);
nand U11844 (N_11844,N_11724,N_11664);
xor U11845 (N_11845,N_11569,N_11564);
and U11846 (N_11846,N_11715,N_11586);
nand U11847 (N_11847,N_11635,N_11562);
xnor U11848 (N_11848,N_11589,N_11659);
xnor U11849 (N_11849,N_11525,N_11649);
nor U11850 (N_11850,N_11700,N_11502);
nor U11851 (N_11851,N_11691,N_11556);
or U11852 (N_11852,N_11654,N_11719);
and U11853 (N_11853,N_11731,N_11567);
nand U11854 (N_11854,N_11737,N_11694);
and U11855 (N_11855,N_11602,N_11667);
and U11856 (N_11856,N_11555,N_11735);
or U11857 (N_11857,N_11533,N_11711);
or U11858 (N_11858,N_11630,N_11702);
nor U11859 (N_11859,N_11621,N_11604);
nand U11860 (N_11860,N_11537,N_11622);
nor U11861 (N_11861,N_11598,N_11591);
nor U11862 (N_11862,N_11575,N_11666);
xnor U11863 (N_11863,N_11685,N_11687);
nor U11864 (N_11864,N_11704,N_11733);
nand U11865 (N_11865,N_11660,N_11507);
and U11866 (N_11866,N_11637,N_11612);
nand U11867 (N_11867,N_11508,N_11594);
nor U11868 (N_11868,N_11732,N_11505);
nand U11869 (N_11869,N_11663,N_11549);
nand U11870 (N_11870,N_11650,N_11705);
nand U11871 (N_11871,N_11633,N_11720);
and U11872 (N_11872,N_11657,N_11709);
or U11873 (N_11873,N_11661,N_11674);
or U11874 (N_11874,N_11571,N_11665);
xnor U11875 (N_11875,N_11594,N_11572);
nor U11876 (N_11876,N_11653,N_11619);
nor U11877 (N_11877,N_11623,N_11745);
or U11878 (N_11878,N_11639,N_11726);
xnor U11879 (N_11879,N_11526,N_11705);
or U11880 (N_11880,N_11601,N_11639);
or U11881 (N_11881,N_11622,N_11687);
xor U11882 (N_11882,N_11676,N_11646);
and U11883 (N_11883,N_11587,N_11653);
or U11884 (N_11884,N_11516,N_11571);
or U11885 (N_11885,N_11669,N_11699);
and U11886 (N_11886,N_11518,N_11736);
or U11887 (N_11887,N_11513,N_11575);
nand U11888 (N_11888,N_11531,N_11743);
or U11889 (N_11889,N_11526,N_11724);
or U11890 (N_11890,N_11719,N_11741);
xor U11891 (N_11891,N_11644,N_11680);
and U11892 (N_11892,N_11515,N_11589);
or U11893 (N_11893,N_11527,N_11730);
and U11894 (N_11894,N_11640,N_11607);
or U11895 (N_11895,N_11629,N_11699);
and U11896 (N_11896,N_11667,N_11579);
xnor U11897 (N_11897,N_11654,N_11632);
nor U11898 (N_11898,N_11505,N_11518);
nor U11899 (N_11899,N_11740,N_11715);
xor U11900 (N_11900,N_11569,N_11735);
nor U11901 (N_11901,N_11512,N_11699);
and U11902 (N_11902,N_11709,N_11615);
nand U11903 (N_11903,N_11588,N_11718);
nand U11904 (N_11904,N_11532,N_11715);
xnor U11905 (N_11905,N_11592,N_11619);
xor U11906 (N_11906,N_11639,N_11645);
or U11907 (N_11907,N_11659,N_11696);
nor U11908 (N_11908,N_11741,N_11720);
and U11909 (N_11909,N_11717,N_11583);
xnor U11910 (N_11910,N_11642,N_11513);
nand U11911 (N_11911,N_11712,N_11727);
or U11912 (N_11912,N_11716,N_11620);
nor U11913 (N_11913,N_11739,N_11715);
or U11914 (N_11914,N_11515,N_11684);
nor U11915 (N_11915,N_11689,N_11510);
nand U11916 (N_11916,N_11533,N_11504);
or U11917 (N_11917,N_11702,N_11624);
nand U11918 (N_11918,N_11703,N_11642);
xor U11919 (N_11919,N_11593,N_11548);
or U11920 (N_11920,N_11508,N_11728);
nand U11921 (N_11921,N_11663,N_11614);
or U11922 (N_11922,N_11675,N_11739);
nor U11923 (N_11923,N_11515,N_11552);
or U11924 (N_11924,N_11630,N_11698);
or U11925 (N_11925,N_11513,N_11707);
and U11926 (N_11926,N_11704,N_11727);
or U11927 (N_11927,N_11696,N_11743);
and U11928 (N_11928,N_11530,N_11670);
and U11929 (N_11929,N_11534,N_11709);
nor U11930 (N_11930,N_11522,N_11705);
or U11931 (N_11931,N_11553,N_11675);
and U11932 (N_11932,N_11567,N_11659);
and U11933 (N_11933,N_11687,N_11745);
or U11934 (N_11934,N_11559,N_11712);
or U11935 (N_11935,N_11600,N_11598);
and U11936 (N_11936,N_11508,N_11646);
and U11937 (N_11937,N_11596,N_11681);
nor U11938 (N_11938,N_11584,N_11607);
nand U11939 (N_11939,N_11510,N_11601);
nor U11940 (N_11940,N_11643,N_11651);
and U11941 (N_11941,N_11576,N_11564);
nand U11942 (N_11942,N_11548,N_11517);
and U11943 (N_11943,N_11615,N_11652);
or U11944 (N_11944,N_11741,N_11728);
nor U11945 (N_11945,N_11690,N_11524);
and U11946 (N_11946,N_11513,N_11738);
or U11947 (N_11947,N_11675,N_11670);
xor U11948 (N_11948,N_11620,N_11747);
nor U11949 (N_11949,N_11638,N_11555);
or U11950 (N_11950,N_11728,N_11731);
and U11951 (N_11951,N_11714,N_11507);
or U11952 (N_11952,N_11670,N_11660);
or U11953 (N_11953,N_11737,N_11613);
nand U11954 (N_11954,N_11505,N_11689);
nor U11955 (N_11955,N_11539,N_11695);
nand U11956 (N_11956,N_11530,N_11629);
nor U11957 (N_11957,N_11571,N_11533);
nor U11958 (N_11958,N_11524,N_11545);
nor U11959 (N_11959,N_11590,N_11655);
and U11960 (N_11960,N_11518,N_11644);
nor U11961 (N_11961,N_11734,N_11655);
nand U11962 (N_11962,N_11658,N_11685);
nand U11963 (N_11963,N_11553,N_11641);
and U11964 (N_11964,N_11704,N_11523);
or U11965 (N_11965,N_11572,N_11672);
xnor U11966 (N_11966,N_11669,N_11727);
xor U11967 (N_11967,N_11510,N_11660);
nor U11968 (N_11968,N_11711,N_11507);
nor U11969 (N_11969,N_11610,N_11530);
nor U11970 (N_11970,N_11649,N_11518);
nor U11971 (N_11971,N_11602,N_11707);
xnor U11972 (N_11972,N_11649,N_11670);
nor U11973 (N_11973,N_11722,N_11630);
nor U11974 (N_11974,N_11682,N_11531);
and U11975 (N_11975,N_11560,N_11648);
nor U11976 (N_11976,N_11722,N_11673);
xnor U11977 (N_11977,N_11663,N_11556);
and U11978 (N_11978,N_11709,N_11513);
nor U11979 (N_11979,N_11553,N_11678);
and U11980 (N_11980,N_11625,N_11606);
nor U11981 (N_11981,N_11570,N_11666);
and U11982 (N_11982,N_11550,N_11604);
nor U11983 (N_11983,N_11743,N_11547);
xor U11984 (N_11984,N_11579,N_11633);
nand U11985 (N_11985,N_11748,N_11626);
xor U11986 (N_11986,N_11508,N_11528);
and U11987 (N_11987,N_11686,N_11574);
nand U11988 (N_11988,N_11610,N_11745);
xor U11989 (N_11989,N_11620,N_11628);
or U11990 (N_11990,N_11660,N_11636);
nand U11991 (N_11991,N_11520,N_11727);
nor U11992 (N_11992,N_11742,N_11618);
and U11993 (N_11993,N_11553,N_11639);
and U11994 (N_11994,N_11718,N_11584);
or U11995 (N_11995,N_11686,N_11602);
nor U11996 (N_11996,N_11507,N_11504);
nand U11997 (N_11997,N_11694,N_11547);
and U11998 (N_11998,N_11660,N_11694);
nor U11999 (N_11999,N_11578,N_11553);
xor U12000 (N_12000,N_11877,N_11991);
xnor U12001 (N_12001,N_11825,N_11973);
and U12002 (N_12002,N_11983,N_11831);
xor U12003 (N_12003,N_11799,N_11979);
and U12004 (N_12004,N_11987,N_11802);
nor U12005 (N_12005,N_11855,N_11892);
or U12006 (N_12006,N_11833,N_11969);
or U12007 (N_12007,N_11863,N_11811);
nand U12008 (N_12008,N_11797,N_11858);
and U12009 (N_12009,N_11787,N_11912);
and U12010 (N_12010,N_11988,N_11792);
nand U12011 (N_12011,N_11813,N_11924);
xor U12012 (N_12012,N_11975,N_11793);
and U12013 (N_12013,N_11849,N_11812);
and U12014 (N_12014,N_11967,N_11822);
xnor U12015 (N_12015,N_11814,N_11996);
and U12016 (N_12016,N_11868,N_11864);
and U12017 (N_12017,N_11982,N_11838);
nand U12018 (N_12018,N_11885,N_11754);
nor U12019 (N_12019,N_11872,N_11840);
or U12020 (N_12020,N_11945,N_11919);
nor U12021 (N_12021,N_11893,N_11785);
and U12022 (N_12022,N_11980,N_11974);
or U12023 (N_12023,N_11894,N_11837);
nand U12024 (N_12024,N_11835,N_11800);
xor U12025 (N_12025,N_11907,N_11901);
nor U12026 (N_12026,N_11751,N_11803);
nand U12027 (N_12027,N_11777,N_11816);
or U12028 (N_12028,N_11949,N_11761);
and U12029 (N_12029,N_11795,N_11783);
or U12030 (N_12030,N_11961,N_11990);
or U12031 (N_12031,N_11915,N_11847);
xnor U12032 (N_12032,N_11756,N_11852);
nand U12033 (N_12033,N_11778,N_11917);
and U12034 (N_12034,N_11869,N_11794);
nand U12035 (N_12035,N_11750,N_11832);
nor U12036 (N_12036,N_11827,N_11861);
nand U12037 (N_12037,N_11879,N_11776);
or U12038 (N_12038,N_11986,N_11817);
xnor U12039 (N_12039,N_11779,N_11759);
nor U12040 (N_12040,N_11804,N_11888);
xnor U12041 (N_12041,N_11758,N_11989);
or U12042 (N_12042,N_11834,N_11951);
xor U12043 (N_12043,N_11752,N_11952);
and U12044 (N_12044,N_11881,N_11993);
nand U12045 (N_12045,N_11981,N_11931);
nand U12046 (N_12046,N_11788,N_11824);
or U12047 (N_12047,N_11760,N_11866);
nand U12048 (N_12048,N_11998,N_11851);
or U12049 (N_12049,N_11842,N_11845);
nor U12050 (N_12050,N_11929,N_11918);
or U12051 (N_12051,N_11768,N_11906);
and U12052 (N_12052,N_11920,N_11939);
xor U12053 (N_12053,N_11977,N_11870);
nor U12054 (N_12054,N_11798,N_11934);
or U12055 (N_12055,N_11757,N_11927);
nor U12056 (N_12056,N_11908,N_11957);
nand U12057 (N_12057,N_11926,N_11904);
or U12058 (N_12058,N_11942,N_11876);
or U12059 (N_12059,N_11997,N_11883);
nor U12060 (N_12060,N_11950,N_11763);
and U12061 (N_12061,N_11999,N_11959);
or U12062 (N_12062,N_11910,N_11905);
xor U12063 (N_12063,N_11958,N_11772);
or U12064 (N_12064,N_11859,N_11805);
xnor U12065 (N_12065,N_11955,N_11923);
and U12066 (N_12066,N_11829,N_11815);
or U12067 (N_12067,N_11984,N_11790);
nor U12068 (N_12068,N_11765,N_11878);
or U12069 (N_12069,N_11806,N_11947);
nor U12070 (N_12070,N_11911,N_11871);
nor U12071 (N_12071,N_11935,N_11887);
and U12072 (N_12072,N_11930,N_11895);
nor U12073 (N_12073,N_11964,N_11938);
or U12074 (N_12074,N_11862,N_11995);
and U12075 (N_12075,N_11775,N_11966);
nor U12076 (N_12076,N_11928,N_11786);
nor U12077 (N_12077,N_11922,N_11826);
and U12078 (N_12078,N_11965,N_11774);
nand U12079 (N_12079,N_11850,N_11769);
and U12080 (N_12080,N_11963,N_11882);
or U12081 (N_12081,N_11857,N_11909);
xnor U12082 (N_12082,N_11985,N_11978);
nand U12083 (N_12083,N_11860,N_11903);
and U12084 (N_12084,N_11767,N_11773);
nor U12085 (N_12085,N_11994,N_11784);
nand U12086 (N_12086,N_11886,N_11764);
or U12087 (N_12087,N_11921,N_11770);
or U12088 (N_12088,N_11970,N_11753);
or U12089 (N_12089,N_11846,N_11941);
nand U12090 (N_12090,N_11916,N_11960);
nor U12091 (N_12091,N_11899,N_11809);
and U12092 (N_12092,N_11801,N_11914);
xor U12093 (N_12093,N_11925,N_11953);
nor U12094 (N_12094,N_11766,N_11856);
or U12095 (N_12095,N_11796,N_11884);
nor U12096 (N_12096,N_11962,N_11830);
xnor U12097 (N_12097,N_11854,N_11972);
and U12098 (N_12098,N_11940,N_11913);
or U12099 (N_12099,N_11808,N_11755);
xnor U12100 (N_12100,N_11762,N_11976);
nor U12101 (N_12101,N_11874,N_11848);
nor U12102 (N_12102,N_11954,N_11841);
or U12103 (N_12103,N_11898,N_11844);
nor U12104 (N_12104,N_11821,N_11791);
or U12105 (N_12105,N_11880,N_11946);
and U12106 (N_12106,N_11971,N_11828);
and U12107 (N_12107,N_11865,N_11902);
xnor U12108 (N_12108,N_11948,N_11943);
or U12109 (N_12109,N_11823,N_11789);
or U12110 (N_12110,N_11944,N_11819);
or U12111 (N_12111,N_11936,N_11896);
and U12112 (N_12112,N_11781,N_11932);
xnor U12113 (N_12113,N_11807,N_11810);
or U12114 (N_12114,N_11873,N_11771);
nor U12115 (N_12115,N_11968,N_11780);
nor U12116 (N_12116,N_11782,N_11889);
nand U12117 (N_12117,N_11933,N_11890);
and U12118 (N_12118,N_11891,N_11956);
nor U12119 (N_12119,N_11836,N_11867);
xnor U12120 (N_12120,N_11992,N_11897);
nor U12121 (N_12121,N_11820,N_11875);
nand U12122 (N_12122,N_11839,N_11900);
or U12123 (N_12123,N_11843,N_11937);
xor U12124 (N_12124,N_11853,N_11818);
xor U12125 (N_12125,N_11952,N_11842);
nor U12126 (N_12126,N_11819,N_11975);
and U12127 (N_12127,N_11998,N_11794);
nor U12128 (N_12128,N_11821,N_11840);
or U12129 (N_12129,N_11959,N_11857);
nor U12130 (N_12130,N_11953,N_11901);
xnor U12131 (N_12131,N_11797,N_11962);
and U12132 (N_12132,N_11946,N_11837);
and U12133 (N_12133,N_11783,N_11817);
or U12134 (N_12134,N_11785,N_11819);
xor U12135 (N_12135,N_11878,N_11902);
xor U12136 (N_12136,N_11962,N_11890);
nand U12137 (N_12137,N_11877,N_11840);
or U12138 (N_12138,N_11912,N_11783);
or U12139 (N_12139,N_11796,N_11904);
xnor U12140 (N_12140,N_11881,N_11825);
or U12141 (N_12141,N_11810,N_11893);
nand U12142 (N_12142,N_11952,N_11775);
nor U12143 (N_12143,N_11905,N_11784);
or U12144 (N_12144,N_11763,N_11934);
and U12145 (N_12145,N_11992,N_11921);
or U12146 (N_12146,N_11922,N_11993);
and U12147 (N_12147,N_11920,N_11753);
and U12148 (N_12148,N_11916,N_11975);
nand U12149 (N_12149,N_11953,N_11811);
nor U12150 (N_12150,N_11842,N_11859);
or U12151 (N_12151,N_11864,N_11962);
nor U12152 (N_12152,N_11760,N_11983);
xnor U12153 (N_12153,N_11990,N_11757);
or U12154 (N_12154,N_11878,N_11940);
nor U12155 (N_12155,N_11972,N_11825);
xnor U12156 (N_12156,N_11909,N_11866);
and U12157 (N_12157,N_11817,N_11892);
or U12158 (N_12158,N_11856,N_11788);
and U12159 (N_12159,N_11989,N_11811);
xnor U12160 (N_12160,N_11963,N_11943);
nand U12161 (N_12161,N_11887,N_11965);
nand U12162 (N_12162,N_11832,N_11773);
xor U12163 (N_12163,N_11834,N_11975);
nor U12164 (N_12164,N_11981,N_11818);
nand U12165 (N_12165,N_11896,N_11871);
nor U12166 (N_12166,N_11764,N_11771);
nor U12167 (N_12167,N_11912,N_11857);
and U12168 (N_12168,N_11886,N_11776);
nand U12169 (N_12169,N_11906,N_11976);
nand U12170 (N_12170,N_11997,N_11773);
or U12171 (N_12171,N_11911,N_11756);
or U12172 (N_12172,N_11976,N_11911);
nand U12173 (N_12173,N_11904,N_11838);
nor U12174 (N_12174,N_11774,N_11885);
nand U12175 (N_12175,N_11974,N_11915);
nor U12176 (N_12176,N_11854,N_11751);
xor U12177 (N_12177,N_11876,N_11846);
xor U12178 (N_12178,N_11835,N_11754);
and U12179 (N_12179,N_11827,N_11862);
or U12180 (N_12180,N_11783,N_11772);
nand U12181 (N_12181,N_11901,N_11971);
nand U12182 (N_12182,N_11848,N_11901);
or U12183 (N_12183,N_11934,N_11864);
and U12184 (N_12184,N_11755,N_11765);
and U12185 (N_12185,N_11971,N_11976);
and U12186 (N_12186,N_11784,N_11956);
nand U12187 (N_12187,N_11829,N_11882);
or U12188 (N_12188,N_11783,N_11816);
nor U12189 (N_12189,N_11997,N_11841);
nand U12190 (N_12190,N_11849,N_11889);
xor U12191 (N_12191,N_11940,N_11840);
and U12192 (N_12192,N_11761,N_11835);
and U12193 (N_12193,N_11807,N_11799);
and U12194 (N_12194,N_11926,N_11936);
xnor U12195 (N_12195,N_11829,N_11816);
nor U12196 (N_12196,N_11899,N_11824);
xor U12197 (N_12197,N_11924,N_11773);
or U12198 (N_12198,N_11841,N_11862);
nand U12199 (N_12199,N_11859,N_11846);
nand U12200 (N_12200,N_11853,N_11766);
nor U12201 (N_12201,N_11852,N_11837);
or U12202 (N_12202,N_11800,N_11887);
or U12203 (N_12203,N_11989,N_11967);
or U12204 (N_12204,N_11854,N_11883);
and U12205 (N_12205,N_11823,N_11756);
xnor U12206 (N_12206,N_11824,N_11982);
and U12207 (N_12207,N_11775,N_11882);
or U12208 (N_12208,N_11941,N_11821);
xnor U12209 (N_12209,N_11985,N_11827);
nor U12210 (N_12210,N_11877,N_11842);
nand U12211 (N_12211,N_11920,N_11851);
xor U12212 (N_12212,N_11906,N_11960);
xor U12213 (N_12213,N_11873,N_11790);
xor U12214 (N_12214,N_11758,N_11756);
nand U12215 (N_12215,N_11801,N_11989);
or U12216 (N_12216,N_11973,N_11826);
xor U12217 (N_12217,N_11878,N_11845);
and U12218 (N_12218,N_11869,N_11805);
nand U12219 (N_12219,N_11902,N_11917);
and U12220 (N_12220,N_11839,N_11803);
xnor U12221 (N_12221,N_11962,N_11775);
nor U12222 (N_12222,N_11860,N_11844);
nand U12223 (N_12223,N_11914,N_11818);
xor U12224 (N_12224,N_11856,N_11949);
and U12225 (N_12225,N_11750,N_11939);
nor U12226 (N_12226,N_11902,N_11758);
nor U12227 (N_12227,N_11867,N_11829);
nand U12228 (N_12228,N_11925,N_11783);
nand U12229 (N_12229,N_11835,N_11785);
nor U12230 (N_12230,N_11880,N_11963);
nor U12231 (N_12231,N_11839,N_11977);
nand U12232 (N_12232,N_11822,N_11777);
and U12233 (N_12233,N_11971,N_11938);
and U12234 (N_12234,N_11774,N_11849);
xnor U12235 (N_12235,N_11938,N_11982);
xnor U12236 (N_12236,N_11934,N_11844);
or U12237 (N_12237,N_11977,N_11854);
nand U12238 (N_12238,N_11899,N_11906);
xnor U12239 (N_12239,N_11905,N_11846);
nor U12240 (N_12240,N_11872,N_11856);
and U12241 (N_12241,N_11888,N_11975);
or U12242 (N_12242,N_11939,N_11968);
nor U12243 (N_12243,N_11848,N_11789);
or U12244 (N_12244,N_11811,N_11870);
nor U12245 (N_12245,N_11995,N_11977);
nor U12246 (N_12246,N_11902,N_11951);
or U12247 (N_12247,N_11882,N_11989);
nor U12248 (N_12248,N_11932,N_11910);
or U12249 (N_12249,N_11774,N_11872);
or U12250 (N_12250,N_12228,N_12004);
xnor U12251 (N_12251,N_12000,N_12174);
nand U12252 (N_12252,N_12186,N_12005);
and U12253 (N_12253,N_12203,N_12189);
nand U12254 (N_12254,N_12077,N_12212);
or U12255 (N_12255,N_12145,N_12168);
nand U12256 (N_12256,N_12011,N_12040);
xnor U12257 (N_12257,N_12080,N_12218);
nand U12258 (N_12258,N_12137,N_12060);
xnor U12259 (N_12259,N_12133,N_12209);
and U12260 (N_12260,N_12113,N_12217);
and U12261 (N_12261,N_12206,N_12117);
xnor U12262 (N_12262,N_12086,N_12207);
nor U12263 (N_12263,N_12041,N_12219);
xnor U12264 (N_12264,N_12239,N_12025);
and U12265 (N_12265,N_12061,N_12127);
nand U12266 (N_12266,N_12130,N_12231);
or U12267 (N_12267,N_12033,N_12043);
nor U12268 (N_12268,N_12120,N_12048);
nor U12269 (N_12269,N_12112,N_12224);
or U12270 (N_12270,N_12072,N_12021);
xor U12271 (N_12271,N_12173,N_12109);
or U12272 (N_12272,N_12099,N_12028);
or U12273 (N_12273,N_12039,N_12079);
or U12274 (N_12274,N_12153,N_12074);
nor U12275 (N_12275,N_12053,N_12183);
nand U12276 (N_12276,N_12190,N_12070);
or U12277 (N_12277,N_12069,N_12066);
nor U12278 (N_12278,N_12124,N_12129);
xnor U12279 (N_12279,N_12215,N_12096);
and U12280 (N_12280,N_12233,N_12042);
xor U12281 (N_12281,N_12022,N_12199);
nand U12282 (N_12282,N_12010,N_12227);
nor U12283 (N_12283,N_12152,N_12101);
xor U12284 (N_12284,N_12121,N_12017);
nor U12285 (N_12285,N_12193,N_12135);
xor U12286 (N_12286,N_12095,N_12093);
xor U12287 (N_12287,N_12001,N_12034);
or U12288 (N_12288,N_12157,N_12177);
nor U12289 (N_12289,N_12084,N_12210);
and U12290 (N_12290,N_12092,N_12027);
xor U12291 (N_12291,N_12223,N_12214);
nand U12292 (N_12292,N_12160,N_12136);
or U12293 (N_12293,N_12155,N_12081);
nand U12294 (N_12294,N_12110,N_12014);
and U12295 (N_12295,N_12198,N_12104);
or U12296 (N_12296,N_12038,N_12171);
and U12297 (N_12297,N_12073,N_12058);
and U12298 (N_12298,N_12249,N_12143);
nor U12299 (N_12299,N_12119,N_12003);
and U12300 (N_12300,N_12236,N_12242);
nor U12301 (N_12301,N_12024,N_12147);
nand U12302 (N_12302,N_12063,N_12082);
nand U12303 (N_12303,N_12123,N_12019);
xor U12304 (N_12304,N_12184,N_12241);
and U12305 (N_12305,N_12037,N_12220);
xor U12306 (N_12306,N_12205,N_12179);
or U12307 (N_12307,N_12211,N_12094);
nand U12308 (N_12308,N_12248,N_12194);
nor U12309 (N_12309,N_12122,N_12100);
and U12310 (N_12310,N_12140,N_12162);
nor U12311 (N_12311,N_12055,N_12247);
xnor U12312 (N_12312,N_12149,N_12196);
nor U12313 (N_12313,N_12240,N_12114);
nand U12314 (N_12314,N_12046,N_12204);
or U12315 (N_12315,N_12076,N_12195);
and U12316 (N_12316,N_12208,N_12134);
nor U12317 (N_12317,N_12016,N_12246);
nor U12318 (N_12318,N_12181,N_12222);
or U12319 (N_12319,N_12185,N_12059);
nand U12320 (N_12320,N_12178,N_12243);
nor U12321 (N_12321,N_12029,N_12083);
nand U12322 (N_12322,N_12244,N_12148);
nand U12323 (N_12323,N_12051,N_12180);
and U12324 (N_12324,N_12187,N_12151);
and U12325 (N_12325,N_12049,N_12031);
nor U12326 (N_12326,N_12126,N_12216);
nor U12327 (N_12327,N_12163,N_12197);
nor U12328 (N_12328,N_12125,N_12237);
nor U12329 (N_12329,N_12230,N_12030);
nor U12330 (N_12330,N_12026,N_12090);
nand U12331 (N_12331,N_12008,N_12146);
nor U12332 (N_12332,N_12118,N_12050);
nor U12333 (N_12333,N_12002,N_12062);
or U12334 (N_12334,N_12235,N_12045);
nand U12335 (N_12335,N_12226,N_12103);
xnor U12336 (N_12336,N_12091,N_12154);
xnor U12337 (N_12337,N_12161,N_12064);
xor U12338 (N_12338,N_12023,N_12191);
or U12339 (N_12339,N_12105,N_12229);
xnor U12340 (N_12340,N_12044,N_12035);
and U12341 (N_12341,N_12175,N_12057);
nor U12342 (N_12342,N_12166,N_12144);
nand U12343 (N_12343,N_12232,N_12102);
xor U12344 (N_12344,N_12188,N_12159);
xnor U12345 (N_12345,N_12116,N_12018);
or U12346 (N_12346,N_12158,N_12007);
nor U12347 (N_12347,N_12139,N_12097);
and U12348 (N_12348,N_12098,N_12172);
or U12349 (N_12349,N_12170,N_12167);
nand U12350 (N_12350,N_12164,N_12213);
and U12351 (N_12351,N_12150,N_12115);
or U12352 (N_12352,N_12065,N_12054);
and U12353 (N_12353,N_12141,N_12245);
nor U12354 (N_12354,N_12032,N_12089);
and U12355 (N_12355,N_12132,N_12087);
and U12356 (N_12356,N_12013,N_12107);
xor U12357 (N_12357,N_12085,N_12075);
xor U12358 (N_12358,N_12128,N_12200);
xor U12359 (N_12359,N_12111,N_12182);
nand U12360 (N_12360,N_12012,N_12052);
nand U12361 (N_12361,N_12221,N_12015);
nor U12362 (N_12362,N_12156,N_12020);
nor U12363 (N_12363,N_12088,N_12108);
nand U12364 (N_12364,N_12176,N_12071);
and U12365 (N_12365,N_12106,N_12078);
and U12366 (N_12366,N_12009,N_12165);
nand U12367 (N_12367,N_12192,N_12138);
nor U12368 (N_12368,N_12006,N_12238);
or U12369 (N_12369,N_12234,N_12131);
nand U12370 (N_12370,N_12202,N_12142);
xor U12371 (N_12371,N_12036,N_12225);
or U12372 (N_12372,N_12169,N_12067);
nand U12373 (N_12373,N_12056,N_12068);
and U12374 (N_12374,N_12047,N_12201);
nand U12375 (N_12375,N_12090,N_12205);
and U12376 (N_12376,N_12113,N_12071);
or U12377 (N_12377,N_12090,N_12011);
nand U12378 (N_12378,N_12193,N_12132);
xor U12379 (N_12379,N_12245,N_12083);
nor U12380 (N_12380,N_12030,N_12084);
nand U12381 (N_12381,N_12117,N_12193);
or U12382 (N_12382,N_12011,N_12002);
or U12383 (N_12383,N_12222,N_12233);
xor U12384 (N_12384,N_12138,N_12015);
xnor U12385 (N_12385,N_12056,N_12194);
and U12386 (N_12386,N_12239,N_12012);
and U12387 (N_12387,N_12202,N_12119);
nor U12388 (N_12388,N_12166,N_12225);
and U12389 (N_12389,N_12086,N_12081);
nor U12390 (N_12390,N_12247,N_12132);
nor U12391 (N_12391,N_12088,N_12035);
nand U12392 (N_12392,N_12112,N_12248);
nor U12393 (N_12393,N_12226,N_12113);
nor U12394 (N_12394,N_12013,N_12182);
nand U12395 (N_12395,N_12057,N_12183);
and U12396 (N_12396,N_12232,N_12240);
nand U12397 (N_12397,N_12243,N_12200);
and U12398 (N_12398,N_12208,N_12204);
nand U12399 (N_12399,N_12028,N_12151);
or U12400 (N_12400,N_12002,N_12061);
and U12401 (N_12401,N_12117,N_12246);
xnor U12402 (N_12402,N_12175,N_12002);
or U12403 (N_12403,N_12046,N_12229);
nor U12404 (N_12404,N_12247,N_12123);
xor U12405 (N_12405,N_12010,N_12162);
and U12406 (N_12406,N_12207,N_12231);
or U12407 (N_12407,N_12001,N_12133);
nand U12408 (N_12408,N_12193,N_12003);
xnor U12409 (N_12409,N_12161,N_12169);
or U12410 (N_12410,N_12032,N_12186);
or U12411 (N_12411,N_12034,N_12188);
xor U12412 (N_12412,N_12023,N_12075);
nor U12413 (N_12413,N_12202,N_12071);
and U12414 (N_12414,N_12010,N_12190);
or U12415 (N_12415,N_12046,N_12132);
nor U12416 (N_12416,N_12008,N_12048);
nand U12417 (N_12417,N_12238,N_12164);
or U12418 (N_12418,N_12044,N_12007);
nor U12419 (N_12419,N_12014,N_12033);
nor U12420 (N_12420,N_12231,N_12094);
and U12421 (N_12421,N_12035,N_12010);
and U12422 (N_12422,N_12202,N_12168);
xnor U12423 (N_12423,N_12197,N_12017);
xnor U12424 (N_12424,N_12171,N_12070);
nand U12425 (N_12425,N_12226,N_12152);
or U12426 (N_12426,N_12127,N_12099);
and U12427 (N_12427,N_12105,N_12124);
xor U12428 (N_12428,N_12169,N_12152);
nor U12429 (N_12429,N_12019,N_12174);
and U12430 (N_12430,N_12221,N_12233);
and U12431 (N_12431,N_12171,N_12084);
nand U12432 (N_12432,N_12100,N_12205);
xnor U12433 (N_12433,N_12076,N_12169);
xnor U12434 (N_12434,N_12058,N_12071);
or U12435 (N_12435,N_12236,N_12192);
or U12436 (N_12436,N_12095,N_12136);
or U12437 (N_12437,N_12148,N_12242);
xor U12438 (N_12438,N_12092,N_12171);
and U12439 (N_12439,N_12204,N_12115);
or U12440 (N_12440,N_12112,N_12231);
nor U12441 (N_12441,N_12225,N_12202);
nand U12442 (N_12442,N_12073,N_12051);
and U12443 (N_12443,N_12100,N_12022);
nand U12444 (N_12444,N_12241,N_12217);
and U12445 (N_12445,N_12083,N_12072);
nand U12446 (N_12446,N_12012,N_12083);
or U12447 (N_12447,N_12157,N_12060);
or U12448 (N_12448,N_12039,N_12101);
nand U12449 (N_12449,N_12180,N_12162);
and U12450 (N_12450,N_12131,N_12096);
or U12451 (N_12451,N_12024,N_12240);
nor U12452 (N_12452,N_12148,N_12220);
xor U12453 (N_12453,N_12173,N_12200);
or U12454 (N_12454,N_12055,N_12007);
or U12455 (N_12455,N_12200,N_12150);
nand U12456 (N_12456,N_12129,N_12064);
or U12457 (N_12457,N_12099,N_12136);
nor U12458 (N_12458,N_12098,N_12187);
nand U12459 (N_12459,N_12053,N_12086);
or U12460 (N_12460,N_12100,N_12026);
nand U12461 (N_12461,N_12002,N_12145);
nor U12462 (N_12462,N_12150,N_12235);
or U12463 (N_12463,N_12175,N_12097);
nand U12464 (N_12464,N_12226,N_12181);
xnor U12465 (N_12465,N_12077,N_12083);
xnor U12466 (N_12466,N_12141,N_12103);
nor U12467 (N_12467,N_12000,N_12163);
xor U12468 (N_12468,N_12207,N_12210);
nand U12469 (N_12469,N_12008,N_12087);
or U12470 (N_12470,N_12144,N_12238);
nand U12471 (N_12471,N_12136,N_12153);
and U12472 (N_12472,N_12145,N_12021);
or U12473 (N_12473,N_12229,N_12241);
xnor U12474 (N_12474,N_12058,N_12070);
nand U12475 (N_12475,N_12247,N_12174);
or U12476 (N_12476,N_12034,N_12128);
xor U12477 (N_12477,N_12185,N_12011);
xor U12478 (N_12478,N_12125,N_12094);
xor U12479 (N_12479,N_12043,N_12170);
or U12480 (N_12480,N_12221,N_12163);
or U12481 (N_12481,N_12035,N_12213);
xnor U12482 (N_12482,N_12152,N_12086);
xor U12483 (N_12483,N_12040,N_12192);
or U12484 (N_12484,N_12144,N_12030);
nand U12485 (N_12485,N_12190,N_12085);
nor U12486 (N_12486,N_12087,N_12239);
or U12487 (N_12487,N_12081,N_12160);
xnor U12488 (N_12488,N_12224,N_12107);
nand U12489 (N_12489,N_12064,N_12202);
or U12490 (N_12490,N_12015,N_12201);
nand U12491 (N_12491,N_12090,N_12004);
xnor U12492 (N_12492,N_12055,N_12196);
xor U12493 (N_12493,N_12090,N_12100);
nand U12494 (N_12494,N_12069,N_12181);
nor U12495 (N_12495,N_12057,N_12042);
xnor U12496 (N_12496,N_12026,N_12132);
xnor U12497 (N_12497,N_12066,N_12221);
nor U12498 (N_12498,N_12174,N_12015);
nand U12499 (N_12499,N_12152,N_12002);
xnor U12500 (N_12500,N_12275,N_12296);
nor U12501 (N_12501,N_12320,N_12298);
or U12502 (N_12502,N_12454,N_12352);
nor U12503 (N_12503,N_12277,N_12403);
nand U12504 (N_12504,N_12332,N_12377);
and U12505 (N_12505,N_12467,N_12395);
or U12506 (N_12506,N_12444,N_12300);
nand U12507 (N_12507,N_12365,N_12495);
and U12508 (N_12508,N_12258,N_12453);
and U12509 (N_12509,N_12416,N_12415);
nor U12510 (N_12510,N_12351,N_12482);
nor U12511 (N_12511,N_12497,N_12355);
nand U12512 (N_12512,N_12478,N_12435);
nand U12513 (N_12513,N_12265,N_12317);
or U12514 (N_12514,N_12329,N_12369);
nor U12515 (N_12515,N_12385,N_12259);
xor U12516 (N_12516,N_12262,N_12330);
nor U12517 (N_12517,N_12489,N_12486);
nand U12518 (N_12518,N_12480,N_12382);
or U12519 (N_12519,N_12418,N_12407);
and U12520 (N_12520,N_12255,N_12284);
and U12521 (N_12521,N_12368,N_12384);
nor U12522 (N_12522,N_12370,N_12421);
or U12523 (N_12523,N_12286,N_12272);
and U12524 (N_12524,N_12305,N_12357);
nand U12525 (N_12525,N_12432,N_12391);
xor U12526 (N_12526,N_12303,N_12412);
or U12527 (N_12527,N_12427,N_12322);
and U12528 (N_12528,N_12267,N_12372);
and U12529 (N_12529,N_12440,N_12419);
nor U12530 (N_12530,N_12269,N_12359);
or U12531 (N_12531,N_12316,N_12289);
nor U12532 (N_12532,N_12402,N_12491);
nand U12533 (N_12533,N_12420,N_12270);
nand U12534 (N_12534,N_12460,N_12333);
nor U12535 (N_12535,N_12297,N_12381);
or U12536 (N_12536,N_12302,N_12490);
nor U12537 (N_12537,N_12325,N_12276);
nand U12538 (N_12538,N_12310,N_12362);
xnor U12539 (N_12539,N_12346,N_12283);
and U12540 (N_12540,N_12442,N_12438);
xnor U12541 (N_12541,N_12373,N_12383);
xnor U12542 (N_12542,N_12363,N_12339);
nor U12543 (N_12543,N_12471,N_12446);
nand U12544 (N_12544,N_12304,N_12464);
nor U12545 (N_12545,N_12301,N_12293);
xor U12546 (N_12546,N_12413,N_12430);
and U12547 (N_12547,N_12319,N_12281);
and U12548 (N_12548,N_12290,N_12498);
or U12549 (N_12549,N_12343,N_12345);
nand U12550 (N_12550,N_12306,N_12285);
and U12551 (N_12551,N_12447,N_12307);
or U12552 (N_12552,N_12251,N_12387);
or U12553 (N_12553,N_12424,N_12459);
nor U12554 (N_12554,N_12308,N_12493);
nand U12555 (N_12555,N_12392,N_12436);
nor U12556 (N_12556,N_12401,N_12326);
xor U12557 (N_12557,N_12474,N_12449);
xnor U12558 (N_12558,N_12280,N_12475);
nor U12559 (N_12559,N_12263,N_12254);
nand U12560 (N_12560,N_12428,N_12426);
and U12561 (N_12561,N_12452,N_12279);
xnor U12562 (N_12562,N_12439,N_12389);
and U12563 (N_12563,N_12484,N_12434);
and U12564 (N_12564,N_12311,N_12398);
nand U12565 (N_12565,N_12410,N_12394);
nor U12566 (N_12566,N_12312,N_12250);
or U12567 (N_12567,N_12399,N_12390);
nand U12568 (N_12568,N_12455,N_12376);
nand U12569 (N_12569,N_12378,N_12462);
and U12570 (N_12570,N_12406,N_12314);
nor U12571 (N_12571,N_12379,N_12386);
nor U12572 (N_12572,N_12487,N_12409);
xor U12573 (N_12573,N_12485,N_12349);
and U12574 (N_12574,N_12331,N_12338);
xnor U12575 (N_12575,N_12469,N_12336);
and U12576 (N_12576,N_12496,N_12252);
xnor U12577 (N_12577,N_12356,N_12294);
nor U12578 (N_12578,N_12422,N_12282);
and U12579 (N_12579,N_12445,N_12268);
or U12580 (N_12580,N_12309,N_12353);
nand U12581 (N_12581,N_12324,N_12463);
xor U12582 (N_12582,N_12492,N_12273);
nand U12583 (N_12583,N_12354,N_12417);
nand U12584 (N_12584,N_12397,N_12340);
and U12585 (N_12585,N_12472,N_12451);
and U12586 (N_12586,N_12466,N_12374);
or U12587 (N_12587,N_12465,N_12347);
nand U12588 (N_12588,N_12358,N_12488);
xnor U12589 (N_12589,N_12425,N_12494);
and U12590 (N_12590,N_12321,N_12456);
xnor U12591 (N_12591,N_12256,N_12360);
or U12592 (N_12592,N_12388,N_12393);
xnor U12593 (N_12593,N_12271,N_12334);
or U12594 (N_12594,N_12364,N_12299);
nor U12595 (N_12595,N_12350,N_12450);
nand U12596 (N_12596,N_12429,N_12375);
xnor U12597 (N_12597,N_12266,N_12405);
and U12598 (N_12598,N_12366,N_12318);
or U12599 (N_12599,N_12291,N_12287);
and U12600 (N_12600,N_12443,N_12433);
and U12601 (N_12601,N_12313,N_12437);
nor U12602 (N_12602,N_12461,N_12361);
and U12603 (N_12603,N_12457,N_12260);
nor U12604 (N_12604,N_12288,N_12264);
and U12605 (N_12605,N_12257,N_12477);
nor U12606 (N_12606,N_12470,N_12274);
nand U12607 (N_12607,N_12448,N_12414);
or U12608 (N_12608,N_12481,N_12328);
nand U12609 (N_12609,N_12335,N_12423);
nand U12610 (N_12610,N_12468,N_12396);
or U12611 (N_12611,N_12344,N_12476);
or U12612 (N_12612,N_12327,N_12431);
nor U12613 (N_12613,N_12278,N_12342);
and U12614 (N_12614,N_12323,N_12483);
and U12615 (N_12615,N_12441,N_12458);
xor U12616 (N_12616,N_12341,N_12404);
nand U12617 (N_12617,N_12292,N_12499);
or U12618 (N_12618,N_12261,N_12253);
or U12619 (N_12619,N_12348,N_12371);
or U12620 (N_12620,N_12408,N_12473);
nand U12621 (N_12621,N_12315,N_12295);
nor U12622 (N_12622,N_12367,N_12337);
nor U12623 (N_12623,N_12411,N_12479);
xnor U12624 (N_12624,N_12380,N_12400);
xor U12625 (N_12625,N_12313,N_12342);
and U12626 (N_12626,N_12434,N_12276);
or U12627 (N_12627,N_12417,N_12256);
or U12628 (N_12628,N_12390,N_12364);
nor U12629 (N_12629,N_12347,N_12257);
xnor U12630 (N_12630,N_12303,N_12456);
and U12631 (N_12631,N_12389,N_12487);
nand U12632 (N_12632,N_12301,N_12391);
and U12633 (N_12633,N_12250,N_12260);
xor U12634 (N_12634,N_12464,N_12429);
nand U12635 (N_12635,N_12320,N_12287);
nand U12636 (N_12636,N_12342,N_12431);
xnor U12637 (N_12637,N_12439,N_12399);
nor U12638 (N_12638,N_12490,N_12470);
xor U12639 (N_12639,N_12451,N_12449);
xnor U12640 (N_12640,N_12319,N_12470);
xor U12641 (N_12641,N_12414,N_12323);
nor U12642 (N_12642,N_12290,N_12305);
and U12643 (N_12643,N_12381,N_12375);
and U12644 (N_12644,N_12300,N_12473);
xor U12645 (N_12645,N_12446,N_12449);
xnor U12646 (N_12646,N_12456,N_12481);
xor U12647 (N_12647,N_12417,N_12360);
nand U12648 (N_12648,N_12290,N_12327);
or U12649 (N_12649,N_12329,N_12389);
xnor U12650 (N_12650,N_12263,N_12413);
nand U12651 (N_12651,N_12342,N_12471);
and U12652 (N_12652,N_12498,N_12336);
xnor U12653 (N_12653,N_12415,N_12319);
xor U12654 (N_12654,N_12314,N_12447);
and U12655 (N_12655,N_12394,N_12359);
nor U12656 (N_12656,N_12479,N_12390);
xnor U12657 (N_12657,N_12363,N_12404);
and U12658 (N_12658,N_12290,N_12337);
nor U12659 (N_12659,N_12282,N_12480);
or U12660 (N_12660,N_12385,N_12396);
xnor U12661 (N_12661,N_12327,N_12442);
xnor U12662 (N_12662,N_12296,N_12416);
and U12663 (N_12663,N_12379,N_12477);
and U12664 (N_12664,N_12454,N_12411);
and U12665 (N_12665,N_12474,N_12366);
and U12666 (N_12666,N_12436,N_12296);
nand U12667 (N_12667,N_12320,N_12374);
nor U12668 (N_12668,N_12491,N_12450);
and U12669 (N_12669,N_12398,N_12418);
nor U12670 (N_12670,N_12360,N_12312);
nor U12671 (N_12671,N_12461,N_12360);
nor U12672 (N_12672,N_12304,N_12307);
xnor U12673 (N_12673,N_12388,N_12349);
xnor U12674 (N_12674,N_12266,N_12306);
xnor U12675 (N_12675,N_12351,N_12316);
xnor U12676 (N_12676,N_12393,N_12419);
xor U12677 (N_12677,N_12487,N_12460);
nor U12678 (N_12678,N_12263,N_12372);
nand U12679 (N_12679,N_12461,N_12472);
nor U12680 (N_12680,N_12262,N_12474);
and U12681 (N_12681,N_12389,N_12275);
or U12682 (N_12682,N_12440,N_12389);
or U12683 (N_12683,N_12276,N_12344);
xor U12684 (N_12684,N_12394,N_12339);
nand U12685 (N_12685,N_12289,N_12439);
and U12686 (N_12686,N_12332,N_12395);
xnor U12687 (N_12687,N_12290,N_12471);
and U12688 (N_12688,N_12443,N_12465);
nor U12689 (N_12689,N_12314,N_12382);
nand U12690 (N_12690,N_12436,N_12394);
and U12691 (N_12691,N_12375,N_12377);
nand U12692 (N_12692,N_12369,N_12345);
xnor U12693 (N_12693,N_12365,N_12450);
nand U12694 (N_12694,N_12268,N_12276);
or U12695 (N_12695,N_12328,N_12386);
and U12696 (N_12696,N_12341,N_12439);
nor U12697 (N_12697,N_12392,N_12266);
nor U12698 (N_12698,N_12391,N_12469);
and U12699 (N_12699,N_12462,N_12390);
xnor U12700 (N_12700,N_12456,N_12459);
nor U12701 (N_12701,N_12410,N_12379);
nor U12702 (N_12702,N_12482,N_12451);
and U12703 (N_12703,N_12250,N_12290);
nand U12704 (N_12704,N_12462,N_12389);
nor U12705 (N_12705,N_12397,N_12478);
nand U12706 (N_12706,N_12384,N_12346);
or U12707 (N_12707,N_12266,N_12358);
nand U12708 (N_12708,N_12359,N_12432);
or U12709 (N_12709,N_12329,N_12443);
nor U12710 (N_12710,N_12369,N_12310);
and U12711 (N_12711,N_12315,N_12374);
or U12712 (N_12712,N_12346,N_12350);
nor U12713 (N_12713,N_12413,N_12437);
nand U12714 (N_12714,N_12287,N_12348);
xnor U12715 (N_12715,N_12472,N_12288);
and U12716 (N_12716,N_12389,N_12281);
nor U12717 (N_12717,N_12452,N_12263);
nor U12718 (N_12718,N_12431,N_12305);
or U12719 (N_12719,N_12375,N_12353);
nand U12720 (N_12720,N_12466,N_12271);
nor U12721 (N_12721,N_12256,N_12311);
xor U12722 (N_12722,N_12460,N_12454);
nor U12723 (N_12723,N_12492,N_12290);
or U12724 (N_12724,N_12252,N_12280);
nand U12725 (N_12725,N_12464,N_12446);
and U12726 (N_12726,N_12386,N_12393);
and U12727 (N_12727,N_12378,N_12433);
nor U12728 (N_12728,N_12340,N_12296);
or U12729 (N_12729,N_12407,N_12294);
and U12730 (N_12730,N_12463,N_12384);
xor U12731 (N_12731,N_12271,N_12340);
nand U12732 (N_12732,N_12410,N_12355);
nor U12733 (N_12733,N_12427,N_12420);
nand U12734 (N_12734,N_12380,N_12489);
or U12735 (N_12735,N_12316,N_12359);
and U12736 (N_12736,N_12421,N_12360);
and U12737 (N_12737,N_12286,N_12325);
and U12738 (N_12738,N_12358,N_12263);
or U12739 (N_12739,N_12380,N_12311);
xor U12740 (N_12740,N_12342,N_12425);
or U12741 (N_12741,N_12490,N_12320);
xor U12742 (N_12742,N_12302,N_12359);
and U12743 (N_12743,N_12460,N_12408);
or U12744 (N_12744,N_12301,N_12498);
nor U12745 (N_12745,N_12291,N_12444);
and U12746 (N_12746,N_12354,N_12338);
nand U12747 (N_12747,N_12441,N_12293);
nor U12748 (N_12748,N_12297,N_12466);
nand U12749 (N_12749,N_12485,N_12359);
xnor U12750 (N_12750,N_12535,N_12615);
nand U12751 (N_12751,N_12627,N_12578);
or U12752 (N_12752,N_12719,N_12565);
nor U12753 (N_12753,N_12669,N_12692);
xnor U12754 (N_12754,N_12539,N_12525);
nand U12755 (N_12755,N_12595,N_12637);
xnor U12756 (N_12756,N_12629,N_12665);
nand U12757 (N_12757,N_12700,N_12567);
or U12758 (N_12758,N_12653,N_12675);
and U12759 (N_12759,N_12544,N_12717);
and U12760 (N_12760,N_12620,N_12704);
or U12761 (N_12761,N_12518,N_12531);
and U12762 (N_12762,N_12687,N_12603);
nor U12763 (N_12763,N_12695,N_12621);
and U12764 (N_12764,N_12540,N_12672);
or U12765 (N_12765,N_12721,N_12688);
nor U12766 (N_12766,N_12584,N_12645);
nand U12767 (N_12767,N_12677,N_12650);
xor U12768 (N_12768,N_12566,N_12701);
xnor U12769 (N_12769,N_12682,N_12707);
nand U12770 (N_12770,N_12668,N_12735);
nor U12771 (N_12771,N_12661,N_12689);
nor U12772 (N_12772,N_12607,N_12663);
or U12773 (N_12773,N_12670,N_12749);
nor U12774 (N_12774,N_12593,N_12683);
xnor U12775 (N_12775,N_12555,N_12557);
nand U12776 (N_12776,N_12723,N_12667);
nand U12777 (N_12777,N_12722,N_12718);
nand U12778 (N_12778,N_12710,N_12716);
nand U12779 (N_12779,N_12537,N_12529);
xnor U12780 (N_12780,N_12680,N_12638);
xor U12781 (N_12781,N_12631,N_12737);
nor U12782 (N_12782,N_12583,N_12734);
or U12783 (N_12783,N_12625,N_12523);
and U12784 (N_12784,N_12504,N_12698);
xor U12785 (N_12785,N_12501,N_12724);
nor U12786 (N_12786,N_12727,N_12634);
xnor U12787 (N_12787,N_12635,N_12568);
nand U12788 (N_12788,N_12508,N_12577);
or U12789 (N_12789,N_12736,N_12705);
nand U12790 (N_12790,N_12608,N_12709);
or U12791 (N_12791,N_12641,N_12617);
nand U12792 (N_12792,N_12513,N_12678);
nand U12793 (N_12793,N_12611,N_12626);
nand U12794 (N_12794,N_12706,N_12549);
and U12795 (N_12795,N_12609,N_12624);
or U12796 (N_12796,N_12671,N_12686);
or U12797 (N_12797,N_12576,N_12512);
or U12798 (N_12798,N_12574,N_12536);
or U12799 (N_12799,N_12684,N_12636);
and U12800 (N_12800,N_12703,N_12679);
and U12801 (N_12801,N_12545,N_12569);
nor U12802 (N_12802,N_12581,N_12541);
or U12803 (N_12803,N_12519,N_12509);
xnor U12804 (N_12804,N_12664,N_12674);
nor U12805 (N_12805,N_12511,N_12681);
xnor U12806 (N_12806,N_12748,N_12708);
xnor U12807 (N_12807,N_12628,N_12599);
and U12808 (N_12808,N_12573,N_12690);
nand U12809 (N_12809,N_12622,N_12510);
and U12810 (N_12810,N_12592,N_12676);
xnor U12811 (N_12811,N_12715,N_12600);
or U12812 (N_12812,N_12514,N_12623);
xnor U12813 (N_12813,N_12742,N_12729);
and U12814 (N_12814,N_12740,N_12658);
nor U12815 (N_12815,N_12711,N_12651);
or U12816 (N_12816,N_12613,N_12522);
xnor U12817 (N_12817,N_12575,N_12550);
nor U12818 (N_12818,N_12712,N_12553);
xnor U12819 (N_12819,N_12561,N_12551);
nand U12820 (N_12820,N_12558,N_12570);
nor U12821 (N_12821,N_12702,N_12733);
or U12822 (N_12822,N_12632,N_12604);
and U12823 (N_12823,N_12725,N_12591);
and U12824 (N_12824,N_12521,N_12588);
and U12825 (N_12825,N_12543,N_12647);
nor U12826 (N_12826,N_12554,N_12589);
xnor U12827 (N_12827,N_12560,N_12559);
or U12828 (N_12828,N_12699,N_12696);
or U12829 (N_12829,N_12597,N_12552);
nand U12830 (N_12830,N_12655,N_12659);
nand U12831 (N_12831,N_12547,N_12546);
nor U12832 (N_12832,N_12503,N_12612);
or U12833 (N_12833,N_12614,N_12630);
or U12834 (N_12834,N_12602,N_12713);
nor U12835 (N_12835,N_12657,N_12685);
nand U12836 (N_12836,N_12662,N_12594);
or U12837 (N_12837,N_12744,N_12587);
xnor U12838 (N_12838,N_12601,N_12741);
or U12839 (N_12839,N_12517,N_12526);
or U12840 (N_12840,N_12694,N_12652);
nand U12841 (N_12841,N_12747,N_12738);
or U12842 (N_12842,N_12714,N_12728);
nand U12843 (N_12843,N_12743,N_12580);
xnor U12844 (N_12844,N_12564,N_12562);
and U12845 (N_12845,N_12730,N_12532);
xor U12846 (N_12846,N_12563,N_12582);
nand U12847 (N_12847,N_12691,N_12507);
xnor U12848 (N_12848,N_12640,N_12644);
xnor U12849 (N_12849,N_12520,N_12619);
or U12850 (N_12850,N_12585,N_12596);
and U12851 (N_12851,N_12610,N_12642);
nor U12852 (N_12852,N_12666,N_12660);
nand U12853 (N_12853,N_12746,N_12654);
and U12854 (N_12854,N_12745,N_12524);
xnor U12855 (N_12855,N_12605,N_12542);
nand U12856 (N_12856,N_12506,N_12505);
or U12857 (N_12857,N_12538,N_12673);
nor U12858 (N_12858,N_12739,N_12572);
and U12859 (N_12859,N_12643,N_12516);
nand U12860 (N_12860,N_12548,N_12590);
xor U12861 (N_12861,N_12649,N_12515);
nand U12862 (N_12862,N_12639,N_12646);
and U12863 (N_12863,N_12720,N_12500);
or U12864 (N_12864,N_12618,N_12726);
nor U12865 (N_12865,N_12586,N_12731);
and U12866 (N_12866,N_12571,N_12502);
or U12867 (N_12867,N_12556,N_12656);
nor U12868 (N_12868,N_12530,N_12527);
and U12869 (N_12869,N_12598,N_12693);
or U12870 (N_12870,N_12616,N_12606);
nand U12871 (N_12871,N_12528,N_12633);
nor U12872 (N_12872,N_12697,N_12533);
or U12873 (N_12873,N_12534,N_12732);
nor U12874 (N_12874,N_12579,N_12648);
xnor U12875 (N_12875,N_12714,N_12619);
xnor U12876 (N_12876,N_12607,N_12645);
nand U12877 (N_12877,N_12715,N_12522);
or U12878 (N_12878,N_12659,N_12687);
nor U12879 (N_12879,N_12711,N_12745);
nor U12880 (N_12880,N_12648,N_12612);
or U12881 (N_12881,N_12643,N_12588);
xor U12882 (N_12882,N_12613,N_12646);
xor U12883 (N_12883,N_12583,N_12571);
or U12884 (N_12884,N_12647,N_12558);
or U12885 (N_12885,N_12667,N_12587);
and U12886 (N_12886,N_12605,N_12600);
xor U12887 (N_12887,N_12711,N_12623);
xor U12888 (N_12888,N_12560,N_12558);
or U12889 (N_12889,N_12541,N_12626);
and U12890 (N_12890,N_12669,N_12624);
and U12891 (N_12891,N_12695,N_12532);
nand U12892 (N_12892,N_12684,N_12730);
nor U12893 (N_12893,N_12710,N_12621);
xnor U12894 (N_12894,N_12557,N_12554);
and U12895 (N_12895,N_12648,N_12733);
and U12896 (N_12896,N_12682,N_12609);
xor U12897 (N_12897,N_12507,N_12534);
xnor U12898 (N_12898,N_12616,N_12642);
and U12899 (N_12899,N_12679,N_12685);
xnor U12900 (N_12900,N_12694,N_12517);
and U12901 (N_12901,N_12620,N_12712);
or U12902 (N_12902,N_12717,N_12694);
or U12903 (N_12903,N_12668,N_12636);
nand U12904 (N_12904,N_12628,N_12531);
or U12905 (N_12905,N_12715,N_12564);
and U12906 (N_12906,N_12596,N_12661);
or U12907 (N_12907,N_12577,N_12679);
or U12908 (N_12908,N_12616,N_12706);
nand U12909 (N_12909,N_12625,N_12560);
nand U12910 (N_12910,N_12551,N_12651);
or U12911 (N_12911,N_12721,N_12746);
and U12912 (N_12912,N_12501,N_12538);
nor U12913 (N_12913,N_12724,N_12530);
nor U12914 (N_12914,N_12535,N_12540);
xnor U12915 (N_12915,N_12683,N_12654);
nor U12916 (N_12916,N_12711,N_12703);
or U12917 (N_12917,N_12685,N_12744);
nand U12918 (N_12918,N_12606,N_12534);
nand U12919 (N_12919,N_12727,N_12743);
nand U12920 (N_12920,N_12529,N_12595);
and U12921 (N_12921,N_12539,N_12513);
nand U12922 (N_12922,N_12677,N_12636);
nor U12923 (N_12923,N_12693,N_12560);
nand U12924 (N_12924,N_12561,N_12613);
xnor U12925 (N_12925,N_12682,N_12659);
nor U12926 (N_12926,N_12650,N_12741);
nor U12927 (N_12927,N_12533,N_12557);
or U12928 (N_12928,N_12505,N_12681);
xnor U12929 (N_12929,N_12744,N_12573);
or U12930 (N_12930,N_12714,N_12572);
nand U12931 (N_12931,N_12534,N_12668);
nand U12932 (N_12932,N_12662,N_12744);
or U12933 (N_12933,N_12720,N_12584);
or U12934 (N_12934,N_12689,N_12692);
nor U12935 (N_12935,N_12740,N_12565);
or U12936 (N_12936,N_12613,N_12543);
or U12937 (N_12937,N_12735,N_12610);
xor U12938 (N_12938,N_12518,N_12730);
or U12939 (N_12939,N_12743,N_12518);
nand U12940 (N_12940,N_12709,N_12522);
or U12941 (N_12941,N_12545,N_12542);
or U12942 (N_12942,N_12512,N_12519);
xor U12943 (N_12943,N_12503,N_12668);
or U12944 (N_12944,N_12575,N_12627);
xnor U12945 (N_12945,N_12674,N_12651);
xor U12946 (N_12946,N_12533,N_12674);
or U12947 (N_12947,N_12563,N_12738);
and U12948 (N_12948,N_12651,N_12649);
nand U12949 (N_12949,N_12634,N_12740);
nand U12950 (N_12950,N_12568,N_12698);
nor U12951 (N_12951,N_12596,N_12600);
nand U12952 (N_12952,N_12520,N_12539);
xor U12953 (N_12953,N_12569,N_12662);
nor U12954 (N_12954,N_12713,N_12618);
xnor U12955 (N_12955,N_12661,N_12578);
nor U12956 (N_12956,N_12560,N_12716);
and U12957 (N_12957,N_12512,N_12555);
xnor U12958 (N_12958,N_12595,N_12624);
nand U12959 (N_12959,N_12727,N_12534);
xnor U12960 (N_12960,N_12533,N_12605);
or U12961 (N_12961,N_12583,N_12505);
nor U12962 (N_12962,N_12636,N_12584);
and U12963 (N_12963,N_12540,N_12685);
and U12964 (N_12964,N_12694,N_12576);
or U12965 (N_12965,N_12720,N_12601);
nand U12966 (N_12966,N_12734,N_12710);
and U12967 (N_12967,N_12508,N_12733);
or U12968 (N_12968,N_12574,N_12555);
nand U12969 (N_12969,N_12538,N_12607);
nand U12970 (N_12970,N_12741,N_12514);
and U12971 (N_12971,N_12550,N_12584);
nor U12972 (N_12972,N_12614,N_12693);
xor U12973 (N_12973,N_12543,N_12703);
nor U12974 (N_12974,N_12650,N_12658);
nor U12975 (N_12975,N_12526,N_12536);
xor U12976 (N_12976,N_12553,N_12612);
nor U12977 (N_12977,N_12666,N_12580);
xor U12978 (N_12978,N_12507,N_12675);
xnor U12979 (N_12979,N_12540,N_12659);
and U12980 (N_12980,N_12737,N_12703);
xnor U12981 (N_12981,N_12522,N_12654);
and U12982 (N_12982,N_12536,N_12641);
nand U12983 (N_12983,N_12536,N_12582);
xor U12984 (N_12984,N_12526,N_12578);
and U12985 (N_12985,N_12636,N_12620);
xnor U12986 (N_12986,N_12718,N_12589);
and U12987 (N_12987,N_12576,N_12610);
xnor U12988 (N_12988,N_12502,N_12629);
nand U12989 (N_12989,N_12513,N_12592);
xor U12990 (N_12990,N_12514,N_12639);
nor U12991 (N_12991,N_12537,N_12706);
and U12992 (N_12992,N_12718,N_12671);
and U12993 (N_12993,N_12708,N_12696);
and U12994 (N_12994,N_12563,N_12621);
and U12995 (N_12995,N_12746,N_12606);
nand U12996 (N_12996,N_12668,N_12728);
xnor U12997 (N_12997,N_12648,N_12635);
xor U12998 (N_12998,N_12733,N_12684);
nor U12999 (N_12999,N_12730,N_12680);
nor U13000 (N_13000,N_12792,N_12870);
nand U13001 (N_13001,N_12967,N_12986);
and U13002 (N_13002,N_12771,N_12826);
nand U13003 (N_13003,N_12985,N_12820);
nand U13004 (N_13004,N_12893,N_12908);
nand U13005 (N_13005,N_12960,N_12800);
or U13006 (N_13006,N_12807,N_12890);
and U13007 (N_13007,N_12880,N_12858);
and U13008 (N_13008,N_12815,N_12806);
nand U13009 (N_13009,N_12910,N_12899);
xnor U13010 (N_13010,N_12949,N_12816);
or U13011 (N_13011,N_12852,N_12991);
and U13012 (N_13012,N_12918,N_12947);
and U13013 (N_13013,N_12941,N_12838);
xnor U13014 (N_13014,N_12917,N_12886);
nand U13015 (N_13015,N_12773,N_12840);
and U13016 (N_13016,N_12762,N_12769);
nand U13017 (N_13017,N_12878,N_12849);
nor U13018 (N_13018,N_12854,N_12931);
nor U13019 (N_13019,N_12857,N_12760);
nor U13020 (N_13020,N_12959,N_12934);
xnor U13021 (N_13021,N_12909,N_12980);
nand U13022 (N_13022,N_12928,N_12763);
and U13023 (N_13023,N_12919,N_12864);
xor U13024 (N_13024,N_12896,N_12836);
or U13025 (N_13025,N_12932,N_12984);
nor U13026 (N_13026,N_12901,N_12859);
and U13027 (N_13027,N_12784,N_12979);
or U13028 (N_13028,N_12787,N_12781);
and U13029 (N_13029,N_12866,N_12817);
nand U13030 (N_13030,N_12767,N_12798);
nor U13031 (N_13031,N_12923,N_12829);
or U13032 (N_13032,N_12965,N_12810);
and U13033 (N_13033,N_12915,N_12830);
xnor U13034 (N_13034,N_12823,N_12912);
xor U13035 (N_13035,N_12832,N_12873);
and U13036 (N_13036,N_12988,N_12945);
and U13037 (N_13037,N_12944,N_12775);
nor U13038 (N_13038,N_12754,N_12846);
and U13039 (N_13039,N_12990,N_12755);
xor U13040 (N_13040,N_12921,N_12814);
or U13041 (N_13041,N_12853,N_12956);
nand U13042 (N_13042,N_12963,N_12977);
xnor U13043 (N_13043,N_12833,N_12872);
xor U13044 (N_13044,N_12897,N_12793);
nand U13045 (N_13045,N_12939,N_12969);
nand U13046 (N_13046,N_12861,N_12971);
nor U13047 (N_13047,N_12957,N_12879);
or U13048 (N_13048,N_12804,N_12774);
nand U13049 (N_13049,N_12953,N_12785);
and U13050 (N_13050,N_12819,N_12831);
nand U13051 (N_13051,N_12848,N_12906);
and U13052 (N_13052,N_12948,N_12863);
nor U13053 (N_13053,N_12962,N_12885);
nand U13054 (N_13054,N_12779,N_12843);
xor U13055 (N_13055,N_12847,N_12881);
nor U13056 (N_13056,N_12968,N_12751);
nand U13057 (N_13057,N_12976,N_12996);
nand U13058 (N_13058,N_12809,N_12808);
and U13059 (N_13059,N_12877,N_12860);
nand U13060 (N_13060,N_12777,N_12927);
or U13061 (N_13061,N_12835,N_12776);
nor U13062 (N_13062,N_12750,N_12803);
nand U13063 (N_13063,N_12753,N_12812);
xor U13064 (N_13064,N_12994,N_12821);
xnor U13065 (N_13065,N_12813,N_12850);
nand U13066 (N_13066,N_12770,N_12898);
or U13067 (N_13067,N_12936,N_12958);
xnor U13068 (N_13068,N_12995,N_12938);
nand U13069 (N_13069,N_12757,N_12894);
nor U13070 (N_13070,N_12913,N_12801);
nand U13071 (N_13071,N_12768,N_12791);
or U13072 (N_13072,N_12998,N_12972);
and U13073 (N_13073,N_12778,N_12954);
xnor U13074 (N_13074,N_12758,N_12788);
xor U13075 (N_13075,N_12902,N_12765);
nor U13076 (N_13076,N_12865,N_12871);
or U13077 (N_13077,N_12834,N_12891);
nand U13078 (N_13078,N_12887,N_12822);
and U13079 (N_13079,N_12974,N_12895);
nor U13080 (N_13080,N_12935,N_12920);
xor U13081 (N_13081,N_12818,N_12955);
nor U13082 (N_13082,N_12914,N_12855);
or U13083 (N_13083,N_12828,N_12759);
or U13084 (N_13084,N_12876,N_12929);
or U13085 (N_13085,N_12795,N_12827);
or U13086 (N_13086,N_12916,N_12883);
or U13087 (N_13087,N_12761,N_12796);
or U13088 (N_13088,N_12997,N_12797);
nand U13089 (N_13089,N_12951,N_12922);
nor U13090 (N_13090,N_12942,N_12987);
nor U13091 (N_13091,N_12856,N_12904);
xnor U13092 (N_13092,N_12862,N_12766);
or U13093 (N_13093,N_12841,N_12874);
nor U13094 (N_13094,N_12802,N_12952);
nor U13095 (N_13095,N_12845,N_12937);
nor U13096 (N_13096,N_12756,N_12790);
xnor U13097 (N_13097,N_12973,N_12786);
xnor U13098 (N_13098,N_12978,N_12930);
xnor U13099 (N_13099,N_12940,N_12837);
nand U13100 (N_13100,N_12868,N_12842);
or U13101 (N_13101,N_12783,N_12933);
or U13102 (N_13102,N_12946,N_12903);
nor U13103 (N_13103,N_12884,N_12844);
or U13104 (N_13104,N_12888,N_12811);
xnor U13105 (N_13105,N_12825,N_12805);
nor U13106 (N_13106,N_12981,N_12970);
or U13107 (N_13107,N_12875,N_12989);
xnor U13108 (N_13108,N_12889,N_12772);
nand U13109 (N_13109,N_12950,N_12993);
xnor U13110 (N_13110,N_12999,N_12905);
or U13111 (N_13111,N_12982,N_12925);
nand U13112 (N_13112,N_12961,N_12975);
nor U13113 (N_13113,N_12926,N_12764);
xnor U13114 (N_13114,N_12782,N_12839);
and U13115 (N_13115,N_12789,N_12799);
xor U13116 (N_13116,N_12900,N_12869);
nand U13117 (N_13117,N_12882,N_12943);
and U13118 (N_13118,N_12851,N_12964);
xor U13119 (N_13119,N_12780,N_12924);
or U13120 (N_13120,N_12867,N_12824);
nand U13121 (N_13121,N_12907,N_12752);
nand U13122 (N_13122,N_12983,N_12992);
xnor U13123 (N_13123,N_12911,N_12892);
or U13124 (N_13124,N_12794,N_12966);
xor U13125 (N_13125,N_12754,N_12799);
nand U13126 (N_13126,N_12918,N_12764);
nor U13127 (N_13127,N_12777,N_12862);
xor U13128 (N_13128,N_12761,N_12897);
and U13129 (N_13129,N_12962,N_12852);
or U13130 (N_13130,N_12884,N_12813);
and U13131 (N_13131,N_12854,N_12965);
or U13132 (N_13132,N_12919,N_12818);
xor U13133 (N_13133,N_12917,N_12833);
nor U13134 (N_13134,N_12810,N_12916);
xnor U13135 (N_13135,N_12886,N_12853);
and U13136 (N_13136,N_12898,N_12921);
or U13137 (N_13137,N_12813,N_12921);
nor U13138 (N_13138,N_12841,N_12768);
nor U13139 (N_13139,N_12852,N_12824);
or U13140 (N_13140,N_12896,N_12853);
xor U13141 (N_13141,N_12973,N_12975);
and U13142 (N_13142,N_12824,N_12896);
nand U13143 (N_13143,N_12801,N_12902);
xnor U13144 (N_13144,N_12751,N_12952);
nor U13145 (N_13145,N_12928,N_12885);
nor U13146 (N_13146,N_12918,N_12881);
xnor U13147 (N_13147,N_12810,N_12914);
xnor U13148 (N_13148,N_12822,N_12776);
or U13149 (N_13149,N_12933,N_12830);
or U13150 (N_13150,N_12889,N_12943);
nand U13151 (N_13151,N_12774,N_12961);
nand U13152 (N_13152,N_12842,N_12954);
nor U13153 (N_13153,N_12939,N_12964);
xor U13154 (N_13154,N_12984,N_12820);
and U13155 (N_13155,N_12814,N_12982);
and U13156 (N_13156,N_12950,N_12863);
nor U13157 (N_13157,N_12901,N_12811);
and U13158 (N_13158,N_12756,N_12782);
or U13159 (N_13159,N_12803,N_12868);
and U13160 (N_13160,N_12910,N_12757);
nor U13161 (N_13161,N_12998,N_12777);
nand U13162 (N_13162,N_12983,N_12870);
nand U13163 (N_13163,N_12982,N_12804);
nand U13164 (N_13164,N_12790,N_12922);
nor U13165 (N_13165,N_12769,N_12995);
xnor U13166 (N_13166,N_12960,N_12817);
or U13167 (N_13167,N_12813,N_12808);
xor U13168 (N_13168,N_12971,N_12794);
nand U13169 (N_13169,N_12784,N_12792);
xor U13170 (N_13170,N_12960,N_12920);
nor U13171 (N_13171,N_12855,N_12957);
nor U13172 (N_13172,N_12987,N_12800);
nand U13173 (N_13173,N_12811,N_12866);
nor U13174 (N_13174,N_12931,N_12862);
or U13175 (N_13175,N_12794,N_12892);
xnor U13176 (N_13176,N_12850,N_12821);
xor U13177 (N_13177,N_12854,N_12902);
and U13178 (N_13178,N_12971,N_12898);
and U13179 (N_13179,N_12944,N_12878);
xnor U13180 (N_13180,N_12796,N_12876);
nor U13181 (N_13181,N_12786,N_12975);
nand U13182 (N_13182,N_12981,N_12984);
xnor U13183 (N_13183,N_12929,N_12843);
and U13184 (N_13184,N_12927,N_12780);
and U13185 (N_13185,N_12994,N_12853);
xor U13186 (N_13186,N_12767,N_12803);
nand U13187 (N_13187,N_12883,N_12780);
nand U13188 (N_13188,N_12999,N_12909);
and U13189 (N_13189,N_12881,N_12820);
nor U13190 (N_13190,N_12797,N_12999);
nand U13191 (N_13191,N_12836,N_12812);
xor U13192 (N_13192,N_12876,N_12896);
or U13193 (N_13193,N_12984,N_12802);
xor U13194 (N_13194,N_12966,N_12854);
xnor U13195 (N_13195,N_12911,N_12752);
nor U13196 (N_13196,N_12752,N_12926);
nor U13197 (N_13197,N_12856,N_12917);
or U13198 (N_13198,N_12793,N_12827);
nor U13199 (N_13199,N_12986,N_12899);
xor U13200 (N_13200,N_12849,N_12900);
xor U13201 (N_13201,N_12814,N_12915);
and U13202 (N_13202,N_12759,N_12916);
nor U13203 (N_13203,N_12960,N_12772);
xnor U13204 (N_13204,N_12939,N_12792);
or U13205 (N_13205,N_12915,N_12754);
nand U13206 (N_13206,N_12976,N_12774);
or U13207 (N_13207,N_12793,N_12848);
or U13208 (N_13208,N_12811,N_12937);
and U13209 (N_13209,N_12845,N_12835);
and U13210 (N_13210,N_12869,N_12831);
nor U13211 (N_13211,N_12935,N_12799);
xor U13212 (N_13212,N_12796,N_12922);
and U13213 (N_13213,N_12902,N_12787);
and U13214 (N_13214,N_12827,N_12808);
and U13215 (N_13215,N_12781,N_12854);
nor U13216 (N_13216,N_12940,N_12987);
xnor U13217 (N_13217,N_12895,N_12881);
nand U13218 (N_13218,N_12814,N_12960);
xor U13219 (N_13219,N_12901,N_12819);
nor U13220 (N_13220,N_12820,N_12965);
or U13221 (N_13221,N_12879,N_12914);
nand U13222 (N_13222,N_12795,N_12816);
nor U13223 (N_13223,N_12975,N_12847);
and U13224 (N_13224,N_12778,N_12799);
xnor U13225 (N_13225,N_12964,N_12969);
nor U13226 (N_13226,N_12750,N_12782);
xor U13227 (N_13227,N_12847,N_12923);
nor U13228 (N_13228,N_12784,N_12864);
xor U13229 (N_13229,N_12811,N_12767);
or U13230 (N_13230,N_12766,N_12864);
or U13231 (N_13231,N_12830,N_12965);
or U13232 (N_13232,N_12932,N_12886);
nand U13233 (N_13233,N_12887,N_12795);
xnor U13234 (N_13234,N_12974,N_12788);
or U13235 (N_13235,N_12830,N_12866);
and U13236 (N_13236,N_12915,N_12766);
and U13237 (N_13237,N_12837,N_12960);
nor U13238 (N_13238,N_12839,N_12977);
nor U13239 (N_13239,N_12862,N_12761);
xnor U13240 (N_13240,N_12774,N_12765);
and U13241 (N_13241,N_12924,N_12901);
and U13242 (N_13242,N_12952,N_12817);
or U13243 (N_13243,N_12888,N_12857);
nor U13244 (N_13244,N_12836,N_12981);
and U13245 (N_13245,N_12983,N_12751);
and U13246 (N_13246,N_12942,N_12903);
or U13247 (N_13247,N_12961,N_12786);
nand U13248 (N_13248,N_12911,N_12804);
xnor U13249 (N_13249,N_12765,N_12843);
or U13250 (N_13250,N_13087,N_13146);
xnor U13251 (N_13251,N_13098,N_13217);
and U13252 (N_13252,N_13001,N_13214);
or U13253 (N_13253,N_13111,N_13216);
nand U13254 (N_13254,N_13014,N_13188);
nand U13255 (N_13255,N_13169,N_13059);
xor U13256 (N_13256,N_13152,N_13164);
and U13257 (N_13257,N_13238,N_13208);
nor U13258 (N_13258,N_13226,N_13107);
nor U13259 (N_13259,N_13078,N_13176);
xnor U13260 (N_13260,N_13029,N_13149);
nand U13261 (N_13261,N_13131,N_13187);
nand U13262 (N_13262,N_13018,N_13097);
nand U13263 (N_13263,N_13086,N_13112);
and U13264 (N_13264,N_13142,N_13245);
or U13265 (N_13265,N_13104,N_13051);
and U13266 (N_13266,N_13065,N_13076);
nand U13267 (N_13267,N_13190,N_13241);
nand U13268 (N_13268,N_13175,N_13088);
or U13269 (N_13269,N_13074,N_13004);
and U13270 (N_13270,N_13060,N_13235);
nor U13271 (N_13271,N_13181,N_13171);
nor U13272 (N_13272,N_13047,N_13194);
and U13273 (N_13273,N_13201,N_13093);
xnor U13274 (N_13274,N_13222,N_13031);
xor U13275 (N_13275,N_13027,N_13167);
and U13276 (N_13276,N_13206,N_13158);
xnor U13277 (N_13277,N_13230,N_13148);
nor U13278 (N_13278,N_13044,N_13134);
xor U13279 (N_13279,N_13139,N_13096);
and U13280 (N_13280,N_13079,N_13191);
and U13281 (N_13281,N_13034,N_13198);
xor U13282 (N_13282,N_13002,N_13140);
and U13283 (N_13283,N_13114,N_13117);
xor U13284 (N_13284,N_13227,N_13077);
and U13285 (N_13285,N_13035,N_13143);
nand U13286 (N_13286,N_13013,N_13160);
or U13287 (N_13287,N_13124,N_13066);
and U13288 (N_13288,N_13000,N_13009);
or U13289 (N_13289,N_13224,N_13023);
nand U13290 (N_13290,N_13089,N_13068);
nand U13291 (N_13291,N_13126,N_13057);
and U13292 (N_13292,N_13172,N_13105);
and U13293 (N_13293,N_13150,N_13177);
nand U13294 (N_13294,N_13130,N_13162);
nand U13295 (N_13295,N_13248,N_13006);
nor U13296 (N_13296,N_13147,N_13189);
nor U13297 (N_13297,N_13128,N_13115);
nand U13298 (N_13298,N_13005,N_13081);
or U13299 (N_13299,N_13030,N_13062);
or U13300 (N_13300,N_13050,N_13157);
nand U13301 (N_13301,N_13012,N_13022);
and U13302 (N_13302,N_13102,N_13218);
xor U13303 (N_13303,N_13003,N_13053);
nand U13304 (N_13304,N_13244,N_13151);
xor U13305 (N_13305,N_13174,N_13213);
and U13306 (N_13306,N_13072,N_13084);
or U13307 (N_13307,N_13196,N_13136);
nand U13308 (N_13308,N_13163,N_13122);
nor U13309 (N_13309,N_13073,N_13120);
xor U13310 (N_13310,N_13094,N_13090);
nor U13311 (N_13311,N_13186,N_13135);
or U13312 (N_13312,N_13103,N_13118);
xnor U13313 (N_13313,N_13211,N_13116);
xor U13314 (N_13314,N_13108,N_13199);
or U13315 (N_13315,N_13125,N_13138);
or U13316 (N_13316,N_13168,N_13010);
nor U13317 (N_13317,N_13246,N_13166);
xor U13318 (N_13318,N_13011,N_13080);
nor U13319 (N_13319,N_13215,N_13210);
nor U13320 (N_13320,N_13247,N_13082);
xor U13321 (N_13321,N_13231,N_13165);
xor U13322 (N_13322,N_13159,N_13219);
or U13323 (N_13323,N_13036,N_13161);
xor U13324 (N_13324,N_13209,N_13178);
nand U13325 (N_13325,N_13155,N_13121);
nand U13326 (N_13326,N_13234,N_13048);
nor U13327 (N_13327,N_13067,N_13026);
nand U13328 (N_13328,N_13055,N_13095);
nor U13329 (N_13329,N_13046,N_13032);
xnor U13330 (N_13330,N_13239,N_13020);
nor U13331 (N_13331,N_13229,N_13041);
xnor U13332 (N_13332,N_13156,N_13207);
or U13333 (N_13333,N_13233,N_13184);
xor U13334 (N_13334,N_13069,N_13123);
xor U13335 (N_13335,N_13039,N_13110);
xor U13336 (N_13336,N_13145,N_13049);
nand U13337 (N_13337,N_13232,N_13202);
or U13338 (N_13338,N_13043,N_13173);
and U13339 (N_13339,N_13058,N_13085);
and U13340 (N_13340,N_13025,N_13242);
nor U13341 (N_13341,N_13154,N_13064);
nand U13342 (N_13342,N_13223,N_13197);
nor U13343 (N_13343,N_13007,N_13192);
xor U13344 (N_13344,N_13204,N_13017);
nand U13345 (N_13345,N_13237,N_13170);
xnor U13346 (N_13346,N_13249,N_13052);
or U13347 (N_13347,N_13042,N_13091);
nand U13348 (N_13348,N_13033,N_13040);
nor U13349 (N_13349,N_13100,N_13071);
nand U13350 (N_13350,N_13180,N_13119);
and U13351 (N_13351,N_13129,N_13061);
nand U13352 (N_13352,N_13153,N_13028);
nor U13353 (N_13353,N_13016,N_13133);
or U13354 (N_13354,N_13070,N_13021);
or U13355 (N_13355,N_13024,N_13008);
or U13356 (N_13356,N_13179,N_13240);
or U13357 (N_13357,N_13185,N_13109);
or U13358 (N_13358,N_13054,N_13193);
nor U13359 (N_13359,N_13144,N_13225);
nand U13360 (N_13360,N_13243,N_13220);
nand U13361 (N_13361,N_13056,N_13101);
or U13362 (N_13362,N_13045,N_13099);
or U13363 (N_13363,N_13182,N_13075);
nor U13364 (N_13364,N_13183,N_13127);
and U13365 (N_13365,N_13083,N_13113);
nor U13366 (N_13366,N_13137,N_13195);
and U13367 (N_13367,N_13236,N_13038);
xnor U13368 (N_13368,N_13132,N_13141);
xor U13369 (N_13369,N_13037,N_13212);
or U13370 (N_13370,N_13015,N_13200);
xnor U13371 (N_13371,N_13221,N_13203);
nor U13372 (N_13372,N_13106,N_13205);
nand U13373 (N_13373,N_13019,N_13063);
xnor U13374 (N_13374,N_13228,N_13092);
or U13375 (N_13375,N_13168,N_13052);
nand U13376 (N_13376,N_13013,N_13087);
xnor U13377 (N_13377,N_13107,N_13056);
xor U13378 (N_13378,N_13028,N_13082);
and U13379 (N_13379,N_13075,N_13044);
and U13380 (N_13380,N_13003,N_13135);
or U13381 (N_13381,N_13195,N_13238);
xnor U13382 (N_13382,N_13089,N_13000);
nor U13383 (N_13383,N_13206,N_13088);
and U13384 (N_13384,N_13085,N_13239);
and U13385 (N_13385,N_13144,N_13188);
xnor U13386 (N_13386,N_13010,N_13164);
xnor U13387 (N_13387,N_13142,N_13170);
nand U13388 (N_13388,N_13213,N_13154);
nand U13389 (N_13389,N_13164,N_13016);
or U13390 (N_13390,N_13088,N_13239);
xnor U13391 (N_13391,N_13134,N_13045);
or U13392 (N_13392,N_13196,N_13203);
nor U13393 (N_13393,N_13050,N_13059);
or U13394 (N_13394,N_13247,N_13108);
or U13395 (N_13395,N_13066,N_13141);
or U13396 (N_13396,N_13189,N_13243);
or U13397 (N_13397,N_13026,N_13236);
or U13398 (N_13398,N_13143,N_13019);
nor U13399 (N_13399,N_13002,N_13096);
nand U13400 (N_13400,N_13117,N_13100);
nor U13401 (N_13401,N_13230,N_13144);
nand U13402 (N_13402,N_13142,N_13123);
or U13403 (N_13403,N_13161,N_13123);
or U13404 (N_13404,N_13146,N_13191);
nor U13405 (N_13405,N_13214,N_13117);
nand U13406 (N_13406,N_13197,N_13005);
or U13407 (N_13407,N_13012,N_13203);
nand U13408 (N_13408,N_13122,N_13157);
xor U13409 (N_13409,N_13209,N_13196);
or U13410 (N_13410,N_13035,N_13024);
nand U13411 (N_13411,N_13090,N_13144);
nor U13412 (N_13412,N_13100,N_13234);
or U13413 (N_13413,N_13034,N_13204);
nand U13414 (N_13414,N_13235,N_13154);
xor U13415 (N_13415,N_13100,N_13075);
nand U13416 (N_13416,N_13053,N_13041);
or U13417 (N_13417,N_13104,N_13154);
xnor U13418 (N_13418,N_13191,N_13001);
nand U13419 (N_13419,N_13229,N_13085);
nand U13420 (N_13420,N_13041,N_13192);
and U13421 (N_13421,N_13060,N_13140);
and U13422 (N_13422,N_13113,N_13151);
nor U13423 (N_13423,N_13126,N_13176);
nor U13424 (N_13424,N_13082,N_13200);
nor U13425 (N_13425,N_13136,N_13216);
and U13426 (N_13426,N_13171,N_13154);
and U13427 (N_13427,N_13172,N_13115);
nor U13428 (N_13428,N_13009,N_13022);
xor U13429 (N_13429,N_13079,N_13234);
nor U13430 (N_13430,N_13153,N_13184);
or U13431 (N_13431,N_13077,N_13201);
and U13432 (N_13432,N_13013,N_13241);
nor U13433 (N_13433,N_13202,N_13016);
and U13434 (N_13434,N_13061,N_13084);
xor U13435 (N_13435,N_13152,N_13068);
or U13436 (N_13436,N_13051,N_13186);
and U13437 (N_13437,N_13055,N_13166);
or U13438 (N_13438,N_13012,N_13166);
nand U13439 (N_13439,N_13043,N_13225);
nand U13440 (N_13440,N_13214,N_13235);
and U13441 (N_13441,N_13004,N_13042);
or U13442 (N_13442,N_13163,N_13082);
and U13443 (N_13443,N_13046,N_13222);
or U13444 (N_13444,N_13105,N_13212);
and U13445 (N_13445,N_13221,N_13143);
and U13446 (N_13446,N_13099,N_13231);
xor U13447 (N_13447,N_13184,N_13132);
and U13448 (N_13448,N_13018,N_13159);
xnor U13449 (N_13449,N_13074,N_13220);
and U13450 (N_13450,N_13014,N_13095);
or U13451 (N_13451,N_13207,N_13029);
and U13452 (N_13452,N_13030,N_13012);
or U13453 (N_13453,N_13241,N_13221);
and U13454 (N_13454,N_13175,N_13153);
and U13455 (N_13455,N_13196,N_13052);
nand U13456 (N_13456,N_13222,N_13061);
or U13457 (N_13457,N_13016,N_13092);
nand U13458 (N_13458,N_13047,N_13158);
xnor U13459 (N_13459,N_13227,N_13228);
nand U13460 (N_13460,N_13148,N_13012);
nor U13461 (N_13461,N_13114,N_13023);
nor U13462 (N_13462,N_13172,N_13175);
or U13463 (N_13463,N_13150,N_13043);
nand U13464 (N_13464,N_13245,N_13249);
xor U13465 (N_13465,N_13005,N_13131);
nand U13466 (N_13466,N_13074,N_13246);
or U13467 (N_13467,N_13003,N_13066);
or U13468 (N_13468,N_13232,N_13225);
xnor U13469 (N_13469,N_13235,N_13240);
and U13470 (N_13470,N_13239,N_13198);
or U13471 (N_13471,N_13014,N_13036);
or U13472 (N_13472,N_13240,N_13086);
or U13473 (N_13473,N_13126,N_13087);
nand U13474 (N_13474,N_13248,N_13104);
nand U13475 (N_13475,N_13245,N_13102);
and U13476 (N_13476,N_13072,N_13182);
nor U13477 (N_13477,N_13075,N_13228);
nor U13478 (N_13478,N_13241,N_13125);
or U13479 (N_13479,N_13240,N_13183);
nor U13480 (N_13480,N_13147,N_13145);
nor U13481 (N_13481,N_13128,N_13015);
nor U13482 (N_13482,N_13054,N_13187);
nand U13483 (N_13483,N_13203,N_13201);
nand U13484 (N_13484,N_13081,N_13136);
and U13485 (N_13485,N_13184,N_13109);
nor U13486 (N_13486,N_13110,N_13063);
and U13487 (N_13487,N_13082,N_13086);
or U13488 (N_13488,N_13190,N_13103);
xnor U13489 (N_13489,N_13056,N_13133);
and U13490 (N_13490,N_13105,N_13076);
xor U13491 (N_13491,N_13225,N_13068);
or U13492 (N_13492,N_13205,N_13014);
xor U13493 (N_13493,N_13074,N_13169);
and U13494 (N_13494,N_13166,N_13181);
nor U13495 (N_13495,N_13102,N_13052);
and U13496 (N_13496,N_13007,N_13182);
nor U13497 (N_13497,N_13085,N_13176);
xor U13498 (N_13498,N_13168,N_13067);
and U13499 (N_13499,N_13187,N_13188);
and U13500 (N_13500,N_13331,N_13429);
nand U13501 (N_13501,N_13472,N_13345);
and U13502 (N_13502,N_13366,N_13466);
xnor U13503 (N_13503,N_13498,N_13393);
nor U13504 (N_13504,N_13399,N_13297);
nor U13505 (N_13505,N_13317,N_13314);
xnor U13506 (N_13506,N_13383,N_13417);
xor U13507 (N_13507,N_13382,N_13456);
nor U13508 (N_13508,N_13302,N_13435);
and U13509 (N_13509,N_13334,N_13269);
nor U13510 (N_13510,N_13405,N_13279);
and U13511 (N_13511,N_13367,N_13360);
nand U13512 (N_13512,N_13316,N_13319);
nor U13513 (N_13513,N_13357,N_13292);
nor U13514 (N_13514,N_13368,N_13401);
and U13515 (N_13515,N_13352,N_13305);
nand U13516 (N_13516,N_13274,N_13315);
or U13517 (N_13517,N_13348,N_13273);
or U13518 (N_13518,N_13496,N_13422);
or U13519 (N_13519,N_13369,N_13350);
nor U13520 (N_13520,N_13445,N_13493);
xor U13521 (N_13521,N_13388,N_13485);
and U13522 (N_13522,N_13324,N_13270);
nand U13523 (N_13523,N_13252,N_13387);
and U13524 (N_13524,N_13303,N_13403);
nand U13525 (N_13525,N_13420,N_13278);
xor U13526 (N_13526,N_13386,N_13371);
nand U13527 (N_13527,N_13475,N_13397);
and U13528 (N_13528,N_13459,N_13277);
and U13529 (N_13529,N_13436,N_13370);
nor U13530 (N_13530,N_13447,N_13455);
or U13531 (N_13531,N_13355,N_13284);
and U13532 (N_13532,N_13413,N_13379);
xnor U13533 (N_13533,N_13288,N_13294);
and U13534 (N_13534,N_13261,N_13462);
xor U13535 (N_13535,N_13260,N_13442);
nand U13536 (N_13536,N_13257,N_13372);
nor U13537 (N_13537,N_13268,N_13421);
or U13538 (N_13538,N_13451,N_13264);
xor U13539 (N_13539,N_13253,N_13342);
xor U13540 (N_13540,N_13453,N_13416);
nor U13541 (N_13541,N_13365,N_13439);
xor U13542 (N_13542,N_13359,N_13446);
nand U13543 (N_13543,N_13289,N_13255);
and U13544 (N_13544,N_13310,N_13437);
and U13545 (N_13545,N_13259,N_13349);
nor U13546 (N_13546,N_13376,N_13452);
or U13547 (N_13547,N_13250,N_13378);
xnor U13548 (N_13548,N_13384,N_13391);
nor U13549 (N_13549,N_13444,N_13313);
xnor U13550 (N_13550,N_13415,N_13408);
nor U13551 (N_13551,N_13483,N_13341);
or U13552 (N_13552,N_13291,N_13467);
xor U13553 (N_13553,N_13312,N_13428);
xnor U13554 (N_13554,N_13337,N_13364);
xnor U13555 (N_13555,N_13332,N_13263);
xor U13556 (N_13556,N_13308,N_13375);
and U13557 (N_13557,N_13470,N_13419);
or U13558 (N_13558,N_13450,N_13468);
nand U13559 (N_13559,N_13301,N_13344);
xor U13560 (N_13560,N_13356,N_13458);
or U13561 (N_13561,N_13488,N_13374);
xnor U13562 (N_13562,N_13276,N_13290);
nand U13563 (N_13563,N_13339,N_13394);
nand U13564 (N_13564,N_13327,N_13262);
nor U13565 (N_13565,N_13373,N_13463);
and U13566 (N_13566,N_13410,N_13400);
xnor U13567 (N_13567,N_13398,N_13492);
or U13568 (N_13568,N_13361,N_13266);
nor U13569 (N_13569,N_13418,N_13461);
nand U13570 (N_13570,N_13295,N_13333);
xnor U13571 (N_13571,N_13395,N_13473);
xnor U13572 (N_13572,N_13254,N_13487);
xor U13573 (N_13573,N_13464,N_13280);
or U13574 (N_13574,N_13335,N_13265);
or U13575 (N_13575,N_13286,N_13460);
nor U13576 (N_13576,N_13406,N_13469);
nand U13577 (N_13577,N_13304,N_13427);
nand U13578 (N_13578,N_13449,N_13321);
nor U13579 (N_13579,N_13381,N_13283);
xnor U13580 (N_13580,N_13362,N_13499);
or U13581 (N_13581,N_13271,N_13293);
xor U13582 (N_13582,N_13486,N_13340);
nor U13583 (N_13583,N_13402,N_13409);
nand U13584 (N_13584,N_13434,N_13347);
or U13585 (N_13585,N_13484,N_13328);
xor U13586 (N_13586,N_13258,N_13474);
xnor U13587 (N_13587,N_13296,N_13477);
nor U13588 (N_13588,N_13482,N_13354);
and U13589 (N_13589,N_13457,N_13358);
or U13590 (N_13590,N_13256,N_13431);
nand U13591 (N_13591,N_13404,N_13433);
and U13592 (N_13592,N_13251,N_13389);
or U13593 (N_13593,N_13272,N_13299);
or U13594 (N_13594,N_13281,N_13489);
xnor U13595 (N_13595,N_13282,N_13392);
or U13596 (N_13596,N_13432,N_13443);
nand U13597 (N_13597,N_13380,N_13287);
or U13598 (N_13598,N_13298,N_13275);
or U13599 (N_13599,N_13481,N_13407);
and U13600 (N_13600,N_13479,N_13440);
and U13601 (N_13601,N_13497,N_13448);
nor U13602 (N_13602,N_13430,N_13318);
xnor U13603 (N_13603,N_13414,N_13411);
xor U13604 (N_13604,N_13351,N_13385);
nor U13605 (N_13605,N_13320,N_13325);
or U13606 (N_13606,N_13390,N_13311);
xnor U13607 (N_13607,N_13471,N_13478);
nand U13608 (N_13608,N_13438,N_13338);
nor U13609 (N_13609,N_13329,N_13424);
and U13610 (N_13610,N_13346,N_13300);
or U13611 (N_13611,N_13322,N_13480);
or U13612 (N_13612,N_13377,N_13396);
and U13613 (N_13613,N_13490,N_13330);
nand U13614 (N_13614,N_13309,N_13465);
and U13615 (N_13615,N_13426,N_13494);
nand U13616 (N_13616,N_13491,N_13336);
xnor U13617 (N_13617,N_13307,N_13412);
or U13618 (N_13618,N_13495,N_13353);
and U13619 (N_13619,N_13267,N_13476);
nand U13620 (N_13620,N_13285,N_13323);
and U13621 (N_13621,N_13363,N_13425);
nor U13622 (N_13622,N_13441,N_13423);
nor U13623 (N_13623,N_13306,N_13454);
and U13624 (N_13624,N_13326,N_13343);
nand U13625 (N_13625,N_13299,N_13387);
or U13626 (N_13626,N_13386,N_13307);
nand U13627 (N_13627,N_13466,N_13487);
or U13628 (N_13628,N_13482,N_13420);
nand U13629 (N_13629,N_13362,N_13264);
and U13630 (N_13630,N_13425,N_13365);
and U13631 (N_13631,N_13337,N_13481);
or U13632 (N_13632,N_13498,N_13405);
or U13633 (N_13633,N_13357,N_13400);
xor U13634 (N_13634,N_13472,N_13466);
or U13635 (N_13635,N_13394,N_13459);
xor U13636 (N_13636,N_13273,N_13337);
and U13637 (N_13637,N_13412,N_13464);
xnor U13638 (N_13638,N_13431,N_13364);
nor U13639 (N_13639,N_13426,N_13343);
nor U13640 (N_13640,N_13386,N_13449);
and U13641 (N_13641,N_13305,N_13306);
and U13642 (N_13642,N_13348,N_13383);
or U13643 (N_13643,N_13373,N_13331);
nor U13644 (N_13644,N_13269,N_13422);
xor U13645 (N_13645,N_13288,N_13437);
nand U13646 (N_13646,N_13402,N_13326);
nand U13647 (N_13647,N_13489,N_13363);
nor U13648 (N_13648,N_13448,N_13322);
nor U13649 (N_13649,N_13263,N_13408);
nor U13650 (N_13650,N_13344,N_13340);
nor U13651 (N_13651,N_13297,N_13344);
and U13652 (N_13652,N_13285,N_13491);
and U13653 (N_13653,N_13452,N_13442);
nand U13654 (N_13654,N_13314,N_13374);
nor U13655 (N_13655,N_13331,N_13267);
nand U13656 (N_13656,N_13387,N_13467);
nand U13657 (N_13657,N_13341,N_13286);
nand U13658 (N_13658,N_13436,N_13284);
or U13659 (N_13659,N_13339,N_13438);
nor U13660 (N_13660,N_13455,N_13442);
nor U13661 (N_13661,N_13285,N_13390);
nor U13662 (N_13662,N_13305,N_13390);
nor U13663 (N_13663,N_13466,N_13446);
nand U13664 (N_13664,N_13422,N_13493);
xor U13665 (N_13665,N_13343,N_13389);
and U13666 (N_13666,N_13286,N_13492);
nand U13667 (N_13667,N_13287,N_13447);
xor U13668 (N_13668,N_13439,N_13493);
and U13669 (N_13669,N_13274,N_13319);
and U13670 (N_13670,N_13294,N_13427);
nand U13671 (N_13671,N_13321,N_13371);
or U13672 (N_13672,N_13396,N_13498);
nand U13673 (N_13673,N_13320,N_13318);
and U13674 (N_13674,N_13257,N_13262);
and U13675 (N_13675,N_13481,N_13319);
or U13676 (N_13676,N_13338,N_13331);
and U13677 (N_13677,N_13424,N_13498);
nor U13678 (N_13678,N_13445,N_13273);
nor U13679 (N_13679,N_13361,N_13396);
xor U13680 (N_13680,N_13360,N_13450);
nand U13681 (N_13681,N_13357,N_13265);
and U13682 (N_13682,N_13402,N_13480);
nor U13683 (N_13683,N_13310,N_13312);
nor U13684 (N_13684,N_13282,N_13449);
and U13685 (N_13685,N_13296,N_13265);
or U13686 (N_13686,N_13260,N_13346);
and U13687 (N_13687,N_13271,N_13479);
or U13688 (N_13688,N_13404,N_13330);
and U13689 (N_13689,N_13282,N_13382);
nand U13690 (N_13690,N_13409,N_13263);
or U13691 (N_13691,N_13342,N_13390);
and U13692 (N_13692,N_13492,N_13340);
xnor U13693 (N_13693,N_13471,N_13474);
nand U13694 (N_13694,N_13353,N_13368);
and U13695 (N_13695,N_13381,N_13463);
or U13696 (N_13696,N_13439,N_13424);
and U13697 (N_13697,N_13413,N_13434);
xnor U13698 (N_13698,N_13336,N_13375);
and U13699 (N_13699,N_13269,N_13262);
nand U13700 (N_13700,N_13444,N_13437);
or U13701 (N_13701,N_13344,N_13317);
xnor U13702 (N_13702,N_13376,N_13442);
or U13703 (N_13703,N_13391,N_13448);
xnor U13704 (N_13704,N_13274,N_13326);
or U13705 (N_13705,N_13290,N_13389);
nor U13706 (N_13706,N_13341,N_13345);
or U13707 (N_13707,N_13418,N_13472);
xnor U13708 (N_13708,N_13360,N_13466);
xnor U13709 (N_13709,N_13354,N_13401);
and U13710 (N_13710,N_13282,N_13495);
nor U13711 (N_13711,N_13325,N_13381);
and U13712 (N_13712,N_13432,N_13331);
nand U13713 (N_13713,N_13430,N_13427);
nor U13714 (N_13714,N_13498,N_13420);
xnor U13715 (N_13715,N_13483,N_13409);
xor U13716 (N_13716,N_13272,N_13432);
nor U13717 (N_13717,N_13398,N_13367);
nor U13718 (N_13718,N_13421,N_13491);
or U13719 (N_13719,N_13438,N_13269);
nand U13720 (N_13720,N_13272,N_13346);
nor U13721 (N_13721,N_13471,N_13480);
nand U13722 (N_13722,N_13475,N_13310);
and U13723 (N_13723,N_13459,N_13412);
and U13724 (N_13724,N_13353,N_13418);
nand U13725 (N_13725,N_13402,N_13471);
or U13726 (N_13726,N_13336,N_13325);
or U13727 (N_13727,N_13287,N_13453);
nand U13728 (N_13728,N_13342,N_13285);
nand U13729 (N_13729,N_13251,N_13399);
or U13730 (N_13730,N_13402,N_13346);
and U13731 (N_13731,N_13457,N_13321);
and U13732 (N_13732,N_13458,N_13295);
nand U13733 (N_13733,N_13344,N_13311);
nor U13734 (N_13734,N_13438,N_13446);
or U13735 (N_13735,N_13480,N_13403);
nor U13736 (N_13736,N_13452,N_13340);
nand U13737 (N_13737,N_13448,N_13288);
xnor U13738 (N_13738,N_13429,N_13355);
xor U13739 (N_13739,N_13452,N_13285);
nand U13740 (N_13740,N_13292,N_13428);
or U13741 (N_13741,N_13253,N_13302);
nand U13742 (N_13742,N_13277,N_13404);
and U13743 (N_13743,N_13421,N_13346);
xor U13744 (N_13744,N_13396,N_13348);
nand U13745 (N_13745,N_13438,N_13316);
and U13746 (N_13746,N_13439,N_13360);
xnor U13747 (N_13747,N_13363,N_13462);
or U13748 (N_13748,N_13428,N_13476);
nand U13749 (N_13749,N_13331,N_13273);
nand U13750 (N_13750,N_13741,N_13537);
xor U13751 (N_13751,N_13659,N_13623);
or U13752 (N_13752,N_13727,N_13608);
or U13753 (N_13753,N_13574,N_13640);
and U13754 (N_13754,N_13615,N_13590);
nand U13755 (N_13755,N_13735,N_13561);
nor U13756 (N_13756,N_13602,N_13576);
xor U13757 (N_13757,N_13690,N_13664);
xor U13758 (N_13758,N_13725,N_13538);
and U13759 (N_13759,N_13545,N_13655);
and U13760 (N_13760,N_13672,N_13709);
nand U13761 (N_13761,N_13745,N_13631);
and U13762 (N_13762,N_13604,N_13562);
nand U13763 (N_13763,N_13575,N_13714);
or U13764 (N_13764,N_13612,N_13547);
nor U13765 (N_13765,N_13596,N_13606);
and U13766 (N_13766,N_13662,N_13543);
or U13767 (N_13767,N_13658,N_13603);
nor U13768 (N_13768,N_13651,N_13584);
nand U13769 (N_13769,N_13539,N_13694);
nor U13770 (N_13770,N_13678,N_13583);
nor U13771 (N_13771,N_13571,N_13744);
or U13772 (N_13772,N_13724,N_13653);
nor U13773 (N_13773,N_13614,N_13531);
xor U13774 (N_13774,N_13611,N_13564);
nand U13775 (N_13775,N_13514,N_13645);
or U13776 (N_13776,N_13685,N_13568);
xnor U13777 (N_13777,N_13505,N_13675);
nor U13778 (N_13778,N_13665,N_13519);
nand U13779 (N_13779,N_13617,N_13699);
xor U13780 (N_13780,N_13719,N_13679);
nand U13781 (N_13781,N_13683,N_13706);
xnor U13782 (N_13782,N_13667,N_13629);
nand U13783 (N_13783,N_13549,N_13656);
or U13784 (N_13784,N_13573,N_13532);
and U13785 (N_13785,N_13533,N_13668);
xor U13786 (N_13786,N_13593,N_13703);
xor U13787 (N_13787,N_13715,N_13591);
nor U13788 (N_13788,N_13558,N_13747);
and U13789 (N_13789,N_13648,N_13550);
xor U13790 (N_13790,N_13646,N_13647);
xnor U13791 (N_13791,N_13517,N_13691);
or U13792 (N_13792,N_13508,N_13737);
nor U13793 (N_13793,N_13619,N_13693);
xor U13794 (N_13794,N_13594,N_13644);
nor U13795 (N_13795,N_13536,N_13628);
and U13796 (N_13796,N_13605,N_13743);
nand U13797 (N_13797,N_13613,N_13625);
nor U13798 (N_13798,N_13579,N_13524);
or U13799 (N_13799,N_13700,N_13633);
and U13800 (N_13800,N_13513,N_13638);
nor U13801 (N_13801,N_13728,N_13677);
or U13802 (N_13802,N_13726,N_13600);
or U13803 (N_13803,N_13515,N_13541);
nor U13804 (N_13804,N_13544,N_13572);
nor U13805 (N_13805,N_13522,N_13510);
xnor U13806 (N_13806,N_13710,N_13697);
or U13807 (N_13807,N_13501,N_13509);
nor U13808 (N_13808,N_13518,N_13698);
or U13809 (N_13809,N_13618,N_13681);
and U13810 (N_13810,N_13529,N_13595);
and U13811 (N_13811,N_13684,N_13566);
and U13812 (N_13812,N_13707,N_13502);
nand U13813 (N_13813,N_13692,N_13671);
nor U13814 (N_13814,N_13673,N_13557);
nor U13815 (N_13815,N_13704,N_13731);
xor U13816 (N_13816,N_13587,N_13701);
nand U13817 (N_13817,N_13657,N_13551);
xnor U13818 (N_13818,N_13695,N_13607);
or U13819 (N_13819,N_13663,N_13733);
xor U13820 (N_13820,N_13500,N_13530);
or U13821 (N_13821,N_13601,N_13621);
nand U13822 (N_13822,N_13516,N_13748);
and U13823 (N_13823,N_13643,N_13680);
xor U13824 (N_13824,N_13702,N_13676);
or U13825 (N_13825,N_13616,N_13712);
and U13826 (N_13826,N_13555,N_13687);
nand U13827 (N_13827,N_13708,N_13512);
xnor U13828 (N_13828,N_13717,N_13589);
or U13829 (N_13829,N_13540,N_13620);
nand U13830 (N_13830,N_13598,N_13682);
xnor U13831 (N_13831,N_13636,N_13674);
nand U13832 (N_13832,N_13713,N_13736);
xnor U13833 (N_13833,N_13732,N_13506);
nor U13834 (N_13834,N_13634,N_13542);
nor U13835 (N_13835,N_13520,N_13609);
nor U13836 (N_13836,N_13688,N_13632);
nor U13837 (N_13837,N_13592,N_13581);
and U13838 (N_13838,N_13552,N_13718);
or U13839 (N_13839,N_13742,N_13556);
or U13840 (N_13840,N_13548,N_13641);
nor U13841 (N_13841,N_13730,N_13660);
or U13842 (N_13842,N_13720,N_13661);
nor U13843 (N_13843,N_13670,N_13686);
or U13844 (N_13844,N_13585,N_13569);
nor U13845 (N_13845,N_13563,N_13729);
nand U13846 (N_13846,N_13504,N_13630);
and U13847 (N_13847,N_13722,N_13578);
and U13848 (N_13848,N_13734,N_13521);
xor U13849 (N_13849,N_13559,N_13577);
or U13850 (N_13850,N_13553,N_13666);
nand U13851 (N_13851,N_13696,N_13738);
or U13852 (N_13852,N_13586,N_13652);
xnor U13853 (N_13853,N_13639,N_13637);
nor U13854 (N_13854,N_13565,N_13689);
nor U13855 (N_13855,N_13554,N_13740);
xnor U13856 (N_13856,N_13570,N_13716);
and U13857 (N_13857,N_13503,N_13650);
nor U13858 (N_13858,N_13567,N_13534);
xnor U13859 (N_13859,N_13535,N_13749);
nor U13860 (N_13860,N_13711,N_13746);
xor U13861 (N_13861,N_13610,N_13588);
nand U13862 (N_13862,N_13669,N_13599);
nor U13863 (N_13863,N_13654,N_13582);
nor U13864 (N_13864,N_13511,N_13723);
nand U13865 (N_13865,N_13624,N_13626);
or U13866 (N_13866,N_13635,N_13721);
or U13867 (N_13867,N_13580,N_13627);
or U13868 (N_13868,N_13649,N_13705);
nor U13869 (N_13869,N_13507,N_13622);
nor U13870 (N_13870,N_13526,N_13739);
nor U13871 (N_13871,N_13560,N_13642);
xor U13872 (N_13872,N_13597,N_13528);
xnor U13873 (N_13873,N_13546,N_13527);
xor U13874 (N_13874,N_13523,N_13525);
and U13875 (N_13875,N_13647,N_13724);
xnor U13876 (N_13876,N_13653,N_13607);
and U13877 (N_13877,N_13749,N_13520);
and U13878 (N_13878,N_13568,N_13720);
and U13879 (N_13879,N_13736,N_13517);
and U13880 (N_13880,N_13674,N_13567);
and U13881 (N_13881,N_13747,N_13716);
xnor U13882 (N_13882,N_13532,N_13741);
or U13883 (N_13883,N_13663,N_13521);
nor U13884 (N_13884,N_13717,N_13580);
or U13885 (N_13885,N_13738,N_13568);
and U13886 (N_13886,N_13620,N_13626);
xnor U13887 (N_13887,N_13575,N_13560);
nor U13888 (N_13888,N_13719,N_13690);
xnor U13889 (N_13889,N_13553,N_13648);
nor U13890 (N_13890,N_13573,N_13674);
and U13891 (N_13891,N_13737,N_13528);
and U13892 (N_13892,N_13634,N_13712);
xor U13893 (N_13893,N_13508,N_13667);
nand U13894 (N_13894,N_13714,N_13584);
nor U13895 (N_13895,N_13666,N_13529);
and U13896 (N_13896,N_13545,N_13735);
xnor U13897 (N_13897,N_13729,N_13543);
and U13898 (N_13898,N_13696,N_13659);
nand U13899 (N_13899,N_13666,N_13511);
nor U13900 (N_13900,N_13621,N_13669);
and U13901 (N_13901,N_13523,N_13573);
nand U13902 (N_13902,N_13625,N_13652);
xor U13903 (N_13903,N_13736,N_13747);
nand U13904 (N_13904,N_13663,N_13501);
and U13905 (N_13905,N_13668,N_13633);
nor U13906 (N_13906,N_13529,N_13641);
and U13907 (N_13907,N_13673,N_13543);
or U13908 (N_13908,N_13534,N_13684);
or U13909 (N_13909,N_13693,N_13590);
or U13910 (N_13910,N_13587,N_13630);
and U13911 (N_13911,N_13700,N_13501);
nand U13912 (N_13912,N_13508,N_13505);
or U13913 (N_13913,N_13713,N_13603);
nor U13914 (N_13914,N_13577,N_13599);
and U13915 (N_13915,N_13747,N_13526);
nor U13916 (N_13916,N_13689,N_13700);
nand U13917 (N_13917,N_13563,N_13586);
xor U13918 (N_13918,N_13599,N_13572);
xor U13919 (N_13919,N_13663,N_13537);
and U13920 (N_13920,N_13712,N_13710);
nor U13921 (N_13921,N_13508,N_13705);
xnor U13922 (N_13922,N_13571,N_13504);
and U13923 (N_13923,N_13613,N_13609);
and U13924 (N_13924,N_13707,N_13691);
nand U13925 (N_13925,N_13501,N_13598);
and U13926 (N_13926,N_13605,N_13583);
or U13927 (N_13927,N_13533,N_13585);
nand U13928 (N_13928,N_13653,N_13705);
or U13929 (N_13929,N_13559,N_13679);
and U13930 (N_13930,N_13539,N_13707);
nor U13931 (N_13931,N_13726,N_13550);
or U13932 (N_13932,N_13686,N_13571);
or U13933 (N_13933,N_13668,N_13676);
nand U13934 (N_13934,N_13543,N_13716);
or U13935 (N_13935,N_13738,N_13714);
nor U13936 (N_13936,N_13630,N_13560);
or U13937 (N_13937,N_13530,N_13716);
xnor U13938 (N_13938,N_13734,N_13609);
xor U13939 (N_13939,N_13557,N_13742);
xor U13940 (N_13940,N_13606,N_13715);
nand U13941 (N_13941,N_13661,N_13503);
or U13942 (N_13942,N_13506,N_13630);
and U13943 (N_13943,N_13544,N_13655);
and U13944 (N_13944,N_13570,N_13505);
nand U13945 (N_13945,N_13528,N_13534);
or U13946 (N_13946,N_13508,N_13686);
or U13947 (N_13947,N_13651,N_13687);
or U13948 (N_13948,N_13612,N_13721);
nor U13949 (N_13949,N_13685,N_13744);
nand U13950 (N_13950,N_13651,N_13684);
nand U13951 (N_13951,N_13608,N_13582);
and U13952 (N_13952,N_13680,N_13718);
or U13953 (N_13953,N_13674,N_13620);
xor U13954 (N_13954,N_13524,N_13603);
nor U13955 (N_13955,N_13708,N_13689);
xor U13956 (N_13956,N_13596,N_13710);
xor U13957 (N_13957,N_13559,N_13646);
nor U13958 (N_13958,N_13522,N_13669);
and U13959 (N_13959,N_13744,N_13705);
xor U13960 (N_13960,N_13681,N_13540);
nand U13961 (N_13961,N_13724,N_13587);
nand U13962 (N_13962,N_13667,N_13604);
nand U13963 (N_13963,N_13544,N_13517);
or U13964 (N_13964,N_13641,N_13504);
and U13965 (N_13965,N_13615,N_13693);
or U13966 (N_13966,N_13505,N_13516);
xnor U13967 (N_13967,N_13664,N_13739);
xnor U13968 (N_13968,N_13574,N_13502);
xor U13969 (N_13969,N_13743,N_13649);
nor U13970 (N_13970,N_13740,N_13597);
or U13971 (N_13971,N_13716,N_13685);
xor U13972 (N_13972,N_13652,N_13708);
nor U13973 (N_13973,N_13538,N_13653);
and U13974 (N_13974,N_13632,N_13683);
and U13975 (N_13975,N_13603,N_13587);
nor U13976 (N_13976,N_13513,N_13678);
and U13977 (N_13977,N_13713,N_13652);
nand U13978 (N_13978,N_13660,N_13686);
nand U13979 (N_13979,N_13726,N_13529);
nand U13980 (N_13980,N_13604,N_13716);
and U13981 (N_13981,N_13612,N_13607);
and U13982 (N_13982,N_13578,N_13560);
xor U13983 (N_13983,N_13687,N_13611);
and U13984 (N_13984,N_13507,N_13660);
xnor U13985 (N_13985,N_13586,N_13641);
xnor U13986 (N_13986,N_13641,N_13703);
xor U13987 (N_13987,N_13625,N_13527);
and U13988 (N_13988,N_13510,N_13573);
or U13989 (N_13989,N_13501,N_13517);
xor U13990 (N_13990,N_13630,N_13566);
or U13991 (N_13991,N_13546,N_13569);
nand U13992 (N_13992,N_13628,N_13541);
nand U13993 (N_13993,N_13700,N_13612);
or U13994 (N_13994,N_13512,N_13640);
xor U13995 (N_13995,N_13664,N_13597);
and U13996 (N_13996,N_13500,N_13637);
or U13997 (N_13997,N_13647,N_13501);
and U13998 (N_13998,N_13579,N_13749);
and U13999 (N_13999,N_13633,N_13583);
xnor U14000 (N_14000,N_13973,N_13980);
nor U14001 (N_14001,N_13889,N_13761);
xor U14002 (N_14002,N_13842,N_13881);
nor U14003 (N_14003,N_13957,N_13932);
nor U14004 (N_14004,N_13794,N_13783);
xor U14005 (N_14005,N_13813,N_13995);
and U14006 (N_14006,N_13928,N_13873);
or U14007 (N_14007,N_13766,N_13943);
xnor U14008 (N_14008,N_13874,N_13937);
or U14009 (N_14009,N_13836,N_13790);
or U14010 (N_14010,N_13905,N_13996);
and U14011 (N_14011,N_13885,N_13965);
nand U14012 (N_14012,N_13960,N_13899);
or U14013 (N_14013,N_13827,N_13806);
or U14014 (N_14014,N_13918,N_13848);
or U14015 (N_14015,N_13851,N_13812);
or U14016 (N_14016,N_13936,N_13755);
or U14017 (N_14017,N_13803,N_13849);
or U14018 (N_14018,N_13771,N_13951);
xnor U14019 (N_14019,N_13880,N_13789);
nor U14020 (N_14020,N_13954,N_13979);
and U14021 (N_14021,N_13955,N_13784);
or U14022 (N_14022,N_13984,N_13922);
nand U14023 (N_14023,N_13863,N_13909);
nor U14024 (N_14024,N_13990,N_13860);
or U14025 (N_14025,N_13940,N_13752);
xor U14026 (N_14026,N_13769,N_13770);
and U14027 (N_14027,N_13877,N_13974);
and U14028 (N_14028,N_13958,N_13981);
nor U14029 (N_14029,N_13982,N_13792);
xnor U14030 (N_14030,N_13967,N_13826);
xor U14031 (N_14031,N_13798,N_13775);
or U14032 (N_14032,N_13782,N_13938);
nand U14033 (N_14033,N_13994,N_13805);
nand U14034 (N_14034,N_13855,N_13935);
nand U14035 (N_14035,N_13910,N_13912);
xor U14036 (N_14036,N_13866,N_13971);
nand U14037 (N_14037,N_13925,N_13976);
or U14038 (N_14038,N_13953,N_13883);
and U14039 (N_14039,N_13926,N_13787);
and U14040 (N_14040,N_13751,N_13754);
or U14041 (N_14041,N_13944,N_13924);
nand U14042 (N_14042,N_13875,N_13985);
or U14043 (N_14043,N_13818,N_13908);
nor U14044 (N_14044,N_13862,N_13781);
nor U14045 (N_14045,N_13821,N_13966);
nand U14046 (N_14046,N_13872,N_13952);
and U14047 (N_14047,N_13869,N_13948);
nand U14048 (N_14048,N_13864,N_13956);
and U14049 (N_14049,N_13838,N_13823);
nor U14050 (N_14050,N_13799,N_13768);
nor U14051 (N_14051,N_13945,N_13765);
and U14052 (N_14052,N_13993,N_13773);
xnor U14053 (N_14053,N_13941,N_13764);
and U14054 (N_14054,N_13774,N_13837);
nor U14055 (N_14055,N_13999,N_13978);
nor U14056 (N_14056,N_13913,N_13961);
or U14057 (N_14057,N_13856,N_13898);
and U14058 (N_14058,N_13931,N_13970);
or U14059 (N_14059,N_13815,N_13824);
xor U14060 (N_14060,N_13777,N_13830);
or U14061 (N_14061,N_13989,N_13964);
and U14062 (N_14062,N_13897,N_13933);
and U14063 (N_14063,N_13795,N_13896);
nand U14064 (N_14064,N_13882,N_13939);
and U14065 (N_14065,N_13903,N_13804);
and U14066 (N_14066,N_13968,N_13949);
nand U14067 (N_14067,N_13963,N_13844);
and U14068 (N_14068,N_13921,N_13893);
nand U14069 (N_14069,N_13776,N_13758);
xor U14070 (N_14070,N_13919,N_13942);
xor U14071 (N_14071,N_13870,N_13772);
and U14072 (N_14072,N_13847,N_13760);
nor U14073 (N_14073,N_13811,N_13857);
nand U14074 (N_14074,N_13962,N_13901);
nor U14075 (N_14075,N_13950,N_13802);
or U14076 (N_14076,N_13793,N_13756);
or U14077 (N_14077,N_13762,N_13865);
xor U14078 (N_14078,N_13916,N_13785);
nand U14079 (N_14079,N_13843,N_13977);
nand U14080 (N_14080,N_13876,N_13853);
nor U14081 (N_14081,N_13894,N_13797);
and U14082 (N_14082,N_13809,N_13934);
nor U14083 (N_14083,N_13859,N_13819);
nor U14084 (N_14084,N_13778,N_13927);
nor U14085 (N_14085,N_13923,N_13759);
xnor U14086 (N_14086,N_13902,N_13845);
nor U14087 (N_14087,N_13796,N_13895);
nor U14088 (N_14088,N_13914,N_13763);
xnor U14089 (N_14089,N_13891,N_13904);
or U14090 (N_14090,N_13816,N_13808);
or U14091 (N_14091,N_13900,N_13892);
or U14092 (N_14092,N_13890,N_13801);
nand U14093 (N_14093,N_13992,N_13987);
or U14094 (N_14094,N_13839,N_13991);
xor U14095 (N_14095,N_13959,N_13757);
nand U14096 (N_14096,N_13888,N_13753);
or U14097 (N_14097,N_13814,N_13854);
xnor U14098 (N_14098,N_13868,N_13786);
xor U14099 (N_14099,N_13867,N_13907);
and U14100 (N_14100,N_13998,N_13930);
and U14101 (N_14101,N_13861,N_13988);
and U14102 (N_14102,N_13871,N_13828);
and U14103 (N_14103,N_13887,N_13915);
or U14104 (N_14104,N_13834,N_13767);
nor U14105 (N_14105,N_13800,N_13841);
nor U14106 (N_14106,N_13975,N_13820);
nor U14107 (N_14107,N_13807,N_13997);
nor U14108 (N_14108,N_13831,N_13779);
xnor U14109 (N_14109,N_13850,N_13780);
and U14110 (N_14110,N_13846,N_13879);
and U14111 (N_14111,N_13906,N_13884);
nor U14112 (N_14112,N_13929,N_13986);
nor U14113 (N_14113,N_13829,N_13878);
or U14114 (N_14114,N_13833,N_13972);
or U14115 (N_14115,N_13886,N_13946);
nor U14116 (N_14116,N_13810,N_13911);
nand U14117 (N_14117,N_13917,N_13947);
or U14118 (N_14118,N_13835,N_13791);
xor U14119 (N_14119,N_13858,N_13983);
nand U14120 (N_14120,N_13969,N_13825);
nand U14121 (N_14121,N_13750,N_13920);
nand U14122 (N_14122,N_13832,N_13817);
nand U14123 (N_14123,N_13822,N_13852);
or U14124 (N_14124,N_13840,N_13788);
or U14125 (N_14125,N_13777,N_13900);
or U14126 (N_14126,N_13776,N_13980);
nor U14127 (N_14127,N_13829,N_13914);
nand U14128 (N_14128,N_13781,N_13803);
nor U14129 (N_14129,N_13977,N_13957);
or U14130 (N_14130,N_13849,N_13864);
nor U14131 (N_14131,N_13885,N_13848);
or U14132 (N_14132,N_13762,N_13902);
nand U14133 (N_14133,N_13914,N_13821);
nor U14134 (N_14134,N_13847,N_13869);
nor U14135 (N_14135,N_13987,N_13756);
xor U14136 (N_14136,N_13808,N_13956);
nand U14137 (N_14137,N_13910,N_13946);
and U14138 (N_14138,N_13827,N_13908);
or U14139 (N_14139,N_13940,N_13889);
nand U14140 (N_14140,N_13836,N_13861);
nor U14141 (N_14141,N_13862,N_13754);
nor U14142 (N_14142,N_13758,N_13819);
or U14143 (N_14143,N_13989,N_13893);
nand U14144 (N_14144,N_13835,N_13913);
and U14145 (N_14145,N_13828,N_13754);
xor U14146 (N_14146,N_13952,N_13834);
or U14147 (N_14147,N_13915,N_13897);
xor U14148 (N_14148,N_13991,N_13850);
nor U14149 (N_14149,N_13840,N_13899);
xnor U14150 (N_14150,N_13927,N_13756);
and U14151 (N_14151,N_13917,N_13763);
or U14152 (N_14152,N_13987,N_13795);
nand U14153 (N_14153,N_13942,N_13980);
nor U14154 (N_14154,N_13801,N_13907);
xnor U14155 (N_14155,N_13798,N_13916);
xor U14156 (N_14156,N_13942,N_13962);
or U14157 (N_14157,N_13941,N_13962);
nor U14158 (N_14158,N_13925,N_13853);
and U14159 (N_14159,N_13820,N_13886);
and U14160 (N_14160,N_13789,N_13779);
nand U14161 (N_14161,N_13851,N_13843);
nand U14162 (N_14162,N_13754,N_13903);
nand U14163 (N_14163,N_13924,N_13839);
nand U14164 (N_14164,N_13968,N_13966);
and U14165 (N_14165,N_13913,N_13786);
and U14166 (N_14166,N_13764,N_13979);
and U14167 (N_14167,N_13883,N_13776);
or U14168 (N_14168,N_13821,N_13921);
xor U14169 (N_14169,N_13964,N_13863);
or U14170 (N_14170,N_13920,N_13890);
xnor U14171 (N_14171,N_13923,N_13947);
and U14172 (N_14172,N_13800,N_13888);
nor U14173 (N_14173,N_13937,N_13930);
xor U14174 (N_14174,N_13916,N_13983);
xor U14175 (N_14175,N_13844,N_13917);
nand U14176 (N_14176,N_13806,N_13946);
and U14177 (N_14177,N_13985,N_13980);
nand U14178 (N_14178,N_13768,N_13931);
nand U14179 (N_14179,N_13956,N_13936);
nand U14180 (N_14180,N_13918,N_13887);
and U14181 (N_14181,N_13816,N_13880);
or U14182 (N_14182,N_13949,N_13988);
nor U14183 (N_14183,N_13989,N_13965);
or U14184 (N_14184,N_13794,N_13796);
nor U14185 (N_14185,N_13867,N_13805);
nor U14186 (N_14186,N_13887,N_13999);
or U14187 (N_14187,N_13885,N_13847);
nand U14188 (N_14188,N_13949,N_13975);
and U14189 (N_14189,N_13904,N_13798);
and U14190 (N_14190,N_13996,N_13927);
and U14191 (N_14191,N_13805,N_13963);
nor U14192 (N_14192,N_13948,N_13826);
nand U14193 (N_14193,N_13871,N_13844);
nand U14194 (N_14194,N_13887,N_13763);
or U14195 (N_14195,N_13822,N_13963);
nand U14196 (N_14196,N_13813,N_13769);
nor U14197 (N_14197,N_13804,N_13911);
xnor U14198 (N_14198,N_13783,N_13886);
nand U14199 (N_14199,N_13776,N_13915);
xnor U14200 (N_14200,N_13790,N_13978);
nor U14201 (N_14201,N_13775,N_13781);
nand U14202 (N_14202,N_13964,N_13901);
and U14203 (N_14203,N_13965,N_13867);
and U14204 (N_14204,N_13872,N_13833);
or U14205 (N_14205,N_13873,N_13831);
and U14206 (N_14206,N_13870,N_13797);
nand U14207 (N_14207,N_13974,N_13988);
nand U14208 (N_14208,N_13972,N_13901);
nor U14209 (N_14209,N_13907,N_13789);
or U14210 (N_14210,N_13757,N_13781);
or U14211 (N_14211,N_13861,N_13998);
and U14212 (N_14212,N_13947,N_13952);
nand U14213 (N_14213,N_13809,N_13913);
and U14214 (N_14214,N_13968,N_13843);
nor U14215 (N_14215,N_13927,N_13865);
nand U14216 (N_14216,N_13848,N_13860);
nand U14217 (N_14217,N_13847,N_13820);
or U14218 (N_14218,N_13800,N_13940);
xor U14219 (N_14219,N_13950,N_13905);
nand U14220 (N_14220,N_13826,N_13845);
nand U14221 (N_14221,N_13987,N_13894);
or U14222 (N_14222,N_13995,N_13854);
and U14223 (N_14223,N_13799,N_13810);
nor U14224 (N_14224,N_13929,N_13918);
nand U14225 (N_14225,N_13986,N_13930);
or U14226 (N_14226,N_13941,N_13901);
nand U14227 (N_14227,N_13773,N_13862);
or U14228 (N_14228,N_13925,N_13954);
nand U14229 (N_14229,N_13866,N_13756);
and U14230 (N_14230,N_13909,N_13834);
and U14231 (N_14231,N_13833,N_13996);
xor U14232 (N_14232,N_13772,N_13871);
nand U14233 (N_14233,N_13874,N_13776);
or U14234 (N_14234,N_13959,N_13911);
and U14235 (N_14235,N_13871,N_13976);
or U14236 (N_14236,N_13766,N_13981);
xnor U14237 (N_14237,N_13910,N_13829);
xor U14238 (N_14238,N_13863,N_13914);
nor U14239 (N_14239,N_13847,N_13879);
xnor U14240 (N_14240,N_13937,N_13801);
nand U14241 (N_14241,N_13778,N_13793);
xnor U14242 (N_14242,N_13755,N_13778);
nor U14243 (N_14243,N_13879,N_13789);
xnor U14244 (N_14244,N_13874,N_13993);
nand U14245 (N_14245,N_13967,N_13803);
nand U14246 (N_14246,N_13809,N_13927);
nand U14247 (N_14247,N_13875,N_13855);
nor U14248 (N_14248,N_13789,N_13949);
xor U14249 (N_14249,N_13790,N_13769);
or U14250 (N_14250,N_14140,N_14070);
and U14251 (N_14251,N_14142,N_14155);
nor U14252 (N_14252,N_14024,N_14017);
nor U14253 (N_14253,N_14160,N_14247);
nor U14254 (N_14254,N_14203,N_14188);
xor U14255 (N_14255,N_14166,N_14128);
xnor U14256 (N_14256,N_14179,N_14196);
and U14257 (N_14257,N_14236,N_14000);
nand U14258 (N_14258,N_14156,N_14135);
xnor U14259 (N_14259,N_14147,N_14127);
or U14260 (N_14260,N_14032,N_14162);
nand U14261 (N_14261,N_14242,N_14053);
nor U14262 (N_14262,N_14050,N_14089);
nor U14263 (N_14263,N_14194,N_14060);
nand U14264 (N_14264,N_14123,N_14065);
xnor U14265 (N_14265,N_14074,N_14144);
nor U14266 (N_14266,N_14101,N_14022);
nor U14267 (N_14267,N_14034,N_14224);
nor U14268 (N_14268,N_14072,N_14002);
nand U14269 (N_14269,N_14126,N_14043);
nor U14270 (N_14270,N_14057,N_14173);
nand U14271 (N_14271,N_14161,N_14009);
and U14272 (N_14272,N_14030,N_14239);
and U14273 (N_14273,N_14087,N_14149);
and U14274 (N_14274,N_14099,N_14092);
nand U14275 (N_14275,N_14192,N_14201);
or U14276 (N_14276,N_14185,N_14001);
xnor U14277 (N_14277,N_14199,N_14210);
or U14278 (N_14278,N_14103,N_14088);
and U14279 (N_14279,N_14125,N_14231);
nor U14280 (N_14280,N_14221,N_14133);
or U14281 (N_14281,N_14102,N_14091);
and U14282 (N_14282,N_14229,N_14068);
nor U14283 (N_14283,N_14019,N_14211);
and U14284 (N_14284,N_14051,N_14096);
nand U14285 (N_14285,N_14136,N_14115);
xor U14286 (N_14286,N_14045,N_14163);
and U14287 (N_14287,N_14146,N_14207);
xor U14288 (N_14288,N_14226,N_14181);
and U14289 (N_14289,N_14197,N_14040);
nand U14290 (N_14290,N_14159,N_14167);
xnor U14291 (N_14291,N_14031,N_14107);
and U14292 (N_14292,N_14122,N_14047);
or U14293 (N_14293,N_14183,N_14212);
nor U14294 (N_14294,N_14238,N_14036);
nand U14295 (N_14295,N_14130,N_14071);
xnor U14296 (N_14296,N_14033,N_14180);
and U14297 (N_14297,N_14028,N_14113);
nor U14298 (N_14298,N_14220,N_14190);
xor U14299 (N_14299,N_14164,N_14094);
nand U14300 (N_14300,N_14139,N_14066);
nor U14301 (N_14301,N_14178,N_14129);
nor U14302 (N_14302,N_14058,N_14061);
nor U14303 (N_14303,N_14174,N_14069);
and U14304 (N_14304,N_14137,N_14154);
nand U14305 (N_14305,N_14084,N_14073);
nand U14306 (N_14306,N_14079,N_14222);
or U14307 (N_14307,N_14014,N_14240);
and U14308 (N_14308,N_14241,N_14219);
nand U14309 (N_14309,N_14108,N_14081);
or U14310 (N_14310,N_14186,N_14213);
xor U14311 (N_14311,N_14052,N_14012);
nand U14312 (N_14312,N_14170,N_14193);
xnor U14313 (N_14313,N_14118,N_14175);
or U14314 (N_14314,N_14208,N_14029);
nor U14315 (N_14315,N_14037,N_14225);
or U14316 (N_14316,N_14243,N_14041);
and U14317 (N_14317,N_14223,N_14067);
nor U14318 (N_14318,N_14228,N_14143);
xnor U14319 (N_14319,N_14076,N_14027);
nand U14320 (N_14320,N_14086,N_14075);
nor U14321 (N_14321,N_14004,N_14152);
nor U14322 (N_14322,N_14165,N_14177);
and U14323 (N_14323,N_14011,N_14080);
nor U14324 (N_14324,N_14049,N_14200);
nor U14325 (N_14325,N_14098,N_14018);
and U14326 (N_14326,N_14205,N_14209);
or U14327 (N_14327,N_14189,N_14046);
nand U14328 (N_14328,N_14120,N_14090);
nor U14329 (N_14329,N_14010,N_14006);
xnor U14330 (N_14330,N_14187,N_14106);
and U14331 (N_14331,N_14008,N_14230);
xnor U14332 (N_14332,N_14114,N_14169);
nor U14333 (N_14333,N_14248,N_14117);
nor U14334 (N_14334,N_14100,N_14148);
xnor U14335 (N_14335,N_14153,N_14131);
nor U14336 (N_14336,N_14138,N_14056);
xnor U14337 (N_14337,N_14063,N_14237);
or U14338 (N_14338,N_14015,N_14121);
and U14339 (N_14339,N_14083,N_14116);
xor U14340 (N_14340,N_14195,N_14202);
xor U14341 (N_14341,N_14059,N_14171);
nand U14342 (N_14342,N_14038,N_14227);
nand U14343 (N_14343,N_14168,N_14244);
and U14344 (N_14344,N_14078,N_14214);
nor U14345 (N_14345,N_14218,N_14206);
and U14346 (N_14346,N_14132,N_14124);
and U14347 (N_14347,N_14003,N_14039);
or U14348 (N_14348,N_14182,N_14042);
nor U14349 (N_14349,N_14054,N_14233);
and U14350 (N_14350,N_14246,N_14025);
or U14351 (N_14351,N_14216,N_14023);
or U14352 (N_14352,N_14016,N_14151);
and U14353 (N_14353,N_14215,N_14112);
or U14354 (N_14354,N_14044,N_14134);
xor U14355 (N_14355,N_14184,N_14191);
xnor U14356 (N_14356,N_14062,N_14235);
and U14357 (N_14357,N_14105,N_14082);
nand U14358 (N_14358,N_14217,N_14026);
xnor U14359 (N_14359,N_14150,N_14232);
xor U14360 (N_14360,N_14198,N_14204);
nand U14361 (N_14361,N_14020,N_14093);
xor U14362 (N_14362,N_14055,N_14110);
nor U14363 (N_14363,N_14109,N_14234);
nor U14364 (N_14364,N_14007,N_14104);
and U14365 (N_14365,N_14085,N_14172);
or U14366 (N_14366,N_14249,N_14097);
and U14367 (N_14367,N_14021,N_14013);
xor U14368 (N_14368,N_14141,N_14119);
and U14369 (N_14369,N_14145,N_14245);
nand U14370 (N_14370,N_14095,N_14048);
nand U14371 (N_14371,N_14005,N_14035);
or U14372 (N_14372,N_14176,N_14158);
nor U14373 (N_14373,N_14157,N_14064);
xor U14374 (N_14374,N_14077,N_14111);
nand U14375 (N_14375,N_14150,N_14054);
xnor U14376 (N_14376,N_14232,N_14081);
xnor U14377 (N_14377,N_14162,N_14057);
or U14378 (N_14378,N_14199,N_14209);
nor U14379 (N_14379,N_14025,N_14125);
or U14380 (N_14380,N_14050,N_14086);
and U14381 (N_14381,N_14189,N_14246);
xnor U14382 (N_14382,N_14215,N_14022);
nor U14383 (N_14383,N_14122,N_14056);
or U14384 (N_14384,N_14078,N_14247);
xor U14385 (N_14385,N_14125,N_14082);
xor U14386 (N_14386,N_14218,N_14187);
nor U14387 (N_14387,N_14071,N_14025);
nand U14388 (N_14388,N_14114,N_14117);
and U14389 (N_14389,N_14125,N_14249);
or U14390 (N_14390,N_14175,N_14138);
nand U14391 (N_14391,N_14146,N_14048);
or U14392 (N_14392,N_14199,N_14043);
nand U14393 (N_14393,N_14007,N_14017);
or U14394 (N_14394,N_14200,N_14230);
nor U14395 (N_14395,N_14240,N_14033);
and U14396 (N_14396,N_14202,N_14205);
nand U14397 (N_14397,N_14077,N_14003);
nor U14398 (N_14398,N_14187,N_14057);
or U14399 (N_14399,N_14088,N_14021);
nand U14400 (N_14400,N_14007,N_14119);
nand U14401 (N_14401,N_14128,N_14161);
or U14402 (N_14402,N_14155,N_14070);
or U14403 (N_14403,N_14205,N_14167);
xor U14404 (N_14404,N_14088,N_14229);
or U14405 (N_14405,N_14227,N_14002);
xor U14406 (N_14406,N_14215,N_14002);
nand U14407 (N_14407,N_14056,N_14077);
and U14408 (N_14408,N_14101,N_14245);
nor U14409 (N_14409,N_14158,N_14059);
or U14410 (N_14410,N_14066,N_14024);
or U14411 (N_14411,N_14180,N_14175);
nor U14412 (N_14412,N_14073,N_14062);
nor U14413 (N_14413,N_14097,N_14160);
xnor U14414 (N_14414,N_14178,N_14006);
and U14415 (N_14415,N_14048,N_14204);
nand U14416 (N_14416,N_14095,N_14059);
nand U14417 (N_14417,N_14001,N_14094);
or U14418 (N_14418,N_14008,N_14240);
xor U14419 (N_14419,N_14193,N_14096);
and U14420 (N_14420,N_14158,N_14081);
nor U14421 (N_14421,N_14023,N_14044);
xnor U14422 (N_14422,N_14033,N_14095);
nand U14423 (N_14423,N_14189,N_14223);
nor U14424 (N_14424,N_14047,N_14111);
nor U14425 (N_14425,N_14176,N_14073);
or U14426 (N_14426,N_14230,N_14069);
nand U14427 (N_14427,N_14046,N_14217);
or U14428 (N_14428,N_14233,N_14040);
nor U14429 (N_14429,N_14138,N_14144);
nand U14430 (N_14430,N_14240,N_14020);
xor U14431 (N_14431,N_14021,N_14238);
xnor U14432 (N_14432,N_14245,N_14199);
and U14433 (N_14433,N_14111,N_14185);
and U14434 (N_14434,N_14018,N_14032);
xor U14435 (N_14435,N_14180,N_14235);
nor U14436 (N_14436,N_14197,N_14079);
xor U14437 (N_14437,N_14126,N_14054);
and U14438 (N_14438,N_14073,N_14207);
nor U14439 (N_14439,N_14125,N_14028);
nor U14440 (N_14440,N_14082,N_14022);
xor U14441 (N_14441,N_14222,N_14085);
nor U14442 (N_14442,N_14047,N_14137);
and U14443 (N_14443,N_14048,N_14155);
xor U14444 (N_14444,N_14154,N_14050);
and U14445 (N_14445,N_14237,N_14119);
xnor U14446 (N_14446,N_14221,N_14083);
nand U14447 (N_14447,N_14022,N_14132);
or U14448 (N_14448,N_14054,N_14156);
nand U14449 (N_14449,N_14131,N_14186);
and U14450 (N_14450,N_14053,N_14198);
or U14451 (N_14451,N_14142,N_14079);
nand U14452 (N_14452,N_14211,N_14153);
and U14453 (N_14453,N_14181,N_14135);
xor U14454 (N_14454,N_14098,N_14053);
or U14455 (N_14455,N_14015,N_14142);
or U14456 (N_14456,N_14027,N_14060);
nor U14457 (N_14457,N_14002,N_14046);
xnor U14458 (N_14458,N_14091,N_14157);
xor U14459 (N_14459,N_14036,N_14152);
and U14460 (N_14460,N_14159,N_14243);
and U14461 (N_14461,N_14109,N_14129);
nand U14462 (N_14462,N_14165,N_14226);
nor U14463 (N_14463,N_14056,N_14007);
nor U14464 (N_14464,N_14004,N_14168);
nor U14465 (N_14465,N_14114,N_14152);
or U14466 (N_14466,N_14177,N_14190);
or U14467 (N_14467,N_14226,N_14065);
xnor U14468 (N_14468,N_14210,N_14169);
and U14469 (N_14469,N_14087,N_14015);
nor U14470 (N_14470,N_14188,N_14091);
or U14471 (N_14471,N_14153,N_14101);
nor U14472 (N_14472,N_14161,N_14108);
nor U14473 (N_14473,N_14049,N_14130);
xnor U14474 (N_14474,N_14222,N_14205);
nor U14475 (N_14475,N_14080,N_14135);
nor U14476 (N_14476,N_14157,N_14218);
nand U14477 (N_14477,N_14159,N_14093);
xnor U14478 (N_14478,N_14036,N_14230);
xor U14479 (N_14479,N_14106,N_14026);
and U14480 (N_14480,N_14137,N_14211);
and U14481 (N_14481,N_14143,N_14006);
nor U14482 (N_14482,N_14053,N_14105);
xor U14483 (N_14483,N_14076,N_14227);
nand U14484 (N_14484,N_14115,N_14056);
or U14485 (N_14485,N_14080,N_14085);
nand U14486 (N_14486,N_14054,N_14039);
nor U14487 (N_14487,N_14033,N_14216);
nor U14488 (N_14488,N_14065,N_14105);
or U14489 (N_14489,N_14214,N_14144);
nand U14490 (N_14490,N_14133,N_14029);
nand U14491 (N_14491,N_14082,N_14214);
nand U14492 (N_14492,N_14025,N_14218);
and U14493 (N_14493,N_14127,N_14216);
xnor U14494 (N_14494,N_14125,N_14008);
or U14495 (N_14495,N_14249,N_14178);
xor U14496 (N_14496,N_14032,N_14114);
and U14497 (N_14497,N_14044,N_14209);
xnor U14498 (N_14498,N_14004,N_14043);
xnor U14499 (N_14499,N_14245,N_14127);
nand U14500 (N_14500,N_14465,N_14295);
xnor U14501 (N_14501,N_14336,N_14488);
nor U14502 (N_14502,N_14396,N_14395);
and U14503 (N_14503,N_14475,N_14346);
nor U14504 (N_14504,N_14397,N_14408);
xor U14505 (N_14505,N_14283,N_14264);
nor U14506 (N_14506,N_14381,N_14262);
and U14507 (N_14507,N_14252,N_14380);
nand U14508 (N_14508,N_14481,N_14403);
or U14509 (N_14509,N_14472,N_14293);
nand U14510 (N_14510,N_14494,N_14431);
nor U14511 (N_14511,N_14423,N_14255);
nand U14512 (N_14512,N_14261,N_14329);
and U14513 (N_14513,N_14299,N_14268);
nand U14514 (N_14514,N_14406,N_14464);
and U14515 (N_14515,N_14487,N_14489);
and U14516 (N_14516,N_14250,N_14445);
nand U14517 (N_14517,N_14368,N_14342);
xor U14518 (N_14518,N_14411,N_14367);
nand U14519 (N_14519,N_14451,N_14458);
xor U14520 (N_14520,N_14450,N_14360);
xor U14521 (N_14521,N_14316,N_14428);
and U14522 (N_14522,N_14492,N_14254);
xor U14523 (N_14523,N_14412,N_14290);
nor U14524 (N_14524,N_14333,N_14476);
and U14525 (N_14525,N_14491,N_14379);
nor U14526 (N_14526,N_14383,N_14343);
and U14527 (N_14527,N_14317,N_14328);
nor U14528 (N_14528,N_14312,N_14345);
and U14529 (N_14529,N_14253,N_14313);
xnor U14530 (N_14530,N_14358,N_14277);
or U14531 (N_14531,N_14448,N_14352);
nand U14532 (N_14532,N_14462,N_14334);
xor U14533 (N_14533,N_14393,N_14292);
nor U14534 (N_14534,N_14394,N_14302);
and U14535 (N_14535,N_14390,N_14427);
and U14536 (N_14536,N_14351,N_14327);
and U14537 (N_14537,N_14256,N_14386);
or U14538 (N_14538,N_14330,N_14442);
nand U14539 (N_14539,N_14400,N_14468);
xor U14540 (N_14540,N_14260,N_14444);
nand U14541 (N_14541,N_14361,N_14371);
and U14542 (N_14542,N_14306,N_14471);
xnor U14543 (N_14543,N_14375,N_14482);
xor U14544 (N_14544,N_14272,N_14259);
and U14545 (N_14545,N_14389,N_14473);
nand U14546 (N_14546,N_14296,N_14314);
nor U14547 (N_14547,N_14307,N_14469);
xor U14548 (N_14548,N_14440,N_14282);
and U14549 (N_14549,N_14294,N_14339);
xor U14550 (N_14550,N_14300,N_14486);
and U14551 (N_14551,N_14422,N_14366);
and U14552 (N_14552,N_14466,N_14439);
and U14553 (N_14553,N_14279,N_14435);
xor U14554 (N_14554,N_14478,N_14474);
nand U14555 (N_14555,N_14387,N_14477);
or U14556 (N_14556,N_14303,N_14480);
or U14557 (N_14557,N_14369,N_14278);
xnor U14558 (N_14558,N_14483,N_14453);
and U14559 (N_14559,N_14308,N_14298);
nor U14560 (N_14560,N_14430,N_14415);
or U14561 (N_14561,N_14407,N_14452);
and U14562 (N_14562,N_14322,N_14349);
nand U14563 (N_14563,N_14271,N_14385);
xor U14564 (N_14564,N_14325,N_14355);
xor U14565 (N_14565,N_14417,N_14461);
xnor U14566 (N_14566,N_14286,N_14350);
nand U14567 (N_14567,N_14401,N_14391);
nand U14568 (N_14568,N_14323,N_14324);
and U14569 (N_14569,N_14421,N_14347);
xnor U14570 (N_14570,N_14269,N_14354);
xor U14571 (N_14571,N_14340,N_14344);
nor U14572 (N_14572,N_14359,N_14257);
nand U14573 (N_14573,N_14485,N_14356);
nor U14574 (N_14574,N_14341,N_14392);
or U14575 (N_14575,N_14495,N_14363);
or U14576 (N_14576,N_14319,N_14398);
xnor U14577 (N_14577,N_14413,N_14365);
or U14578 (N_14578,N_14384,N_14362);
and U14579 (N_14579,N_14479,N_14251);
nor U14580 (N_14580,N_14310,N_14456);
nor U14581 (N_14581,N_14370,N_14467);
xnor U14582 (N_14582,N_14455,N_14420);
and U14583 (N_14583,N_14263,N_14457);
or U14584 (N_14584,N_14402,N_14364);
or U14585 (N_14585,N_14490,N_14425);
and U14586 (N_14586,N_14291,N_14372);
and U14587 (N_14587,N_14348,N_14463);
nand U14588 (N_14588,N_14496,N_14493);
nand U14589 (N_14589,N_14459,N_14416);
and U14590 (N_14590,N_14266,N_14304);
or U14591 (N_14591,N_14353,N_14280);
nor U14592 (N_14592,N_14497,N_14443);
or U14593 (N_14593,N_14331,N_14434);
nand U14594 (N_14594,N_14419,N_14318);
nand U14595 (N_14595,N_14357,N_14399);
or U14596 (N_14596,N_14426,N_14409);
xnor U14597 (N_14597,N_14436,N_14446);
nand U14598 (N_14598,N_14499,N_14433);
nand U14599 (N_14599,N_14382,N_14373);
or U14600 (N_14600,N_14309,N_14258);
or U14601 (N_14601,N_14335,N_14404);
xor U14602 (N_14602,N_14270,N_14311);
xor U14603 (N_14603,N_14388,N_14438);
and U14604 (N_14604,N_14305,N_14281);
nand U14605 (N_14605,N_14321,N_14275);
nor U14606 (N_14606,N_14301,N_14410);
nor U14607 (N_14607,N_14470,N_14284);
and U14608 (N_14608,N_14276,N_14418);
or U14609 (N_14609,N_14405,N_14460);
and U14610 (N_14610,N_14338,N_14337);
xnor U14611 (N_14611,N_14287,N_14273);
nor U14612 (N_14612,N_14432,N_14265);
xor U14613 (N_14613,N_14285,N_14267);
nand U14614 (N_14614,N_14326,N_14437);
nor U14615 (N_14615,N_14289,N_14377);
or U14616 (N_14616,N_14441,N_14320);
nor U14617 (N_14617,N_14315,N_14424);
and U14618 (N_14618,N_14378,N_14498);
or U14619 (N_14619,N_14374,N_14429);
xor U14620 (N_14620,N_14449,N_14297);
and U14621 (N_14621,N_14484,N_14447);
and U14622 (N_14622,N_14454,N_14376);
nor U14623 (N_14623,N_14274,N_14332);
and U14624 (N_14624,N_14414,N_14288);
and U14625 (N_14625,N_14390,N_14350);
xor U14626 (N_14626,N_14295,N_14416);
xor U14627 (N_14627,N_14282,N_14469);
xor U14628 (N_14628,N_14341,N_14480);
xnor U14629 (N_14629,N_14349,N_14448);
nand U14630 (N_14630,N_14405,N_14423);
nor U14631 (N_14631,N_14402,N_14410);
and U14632 (N_14632,N_14292,N_14430);
nand U14633 (N_14633,N_14272,N_14426);
nand U14634 (N_14634,N_14329,N_14266);
nand U14635 (N_14635,N_14338,N_14314);
nor U14636 (N_14636,N_14499,N_14286);
nor U14637 (N_14637,N_14343,N_14317);
or U14638 (N_14638,N_14254,N_14295);
xnor U14639 (N_14639,N_14420,N_14294);
nor U14640 (N_14640,N_14433,N_14468);
nand U14641 (N_14641,N_14485,N_14437);
xnor U14642 (N_14642,N_14338,N_14415);
nand U14643 (N_14643,N_14267,N_14307);
or U14644 (N_14644,N_14265,N_14387);
nor U14645 (N_14645,N_14286,N_14295);
xnor U14646 (N_14646,N_14499,N_14476);
or U14647 (N_14647,N_14491,N_14319);
or U14648 (N_14648,N_14398,N_14459);
xor U14649 (N_14649,N_14479,N_14263);
xor U14650 (N_14650,N_14295,N_14459);
or U14651 (N_14651,N_14445,N_14328);
nand U14652 (N_14652,N_14382,N_14496);
xor U14653 (N_14653,N_14494,N_14268);
nand U14654 (N_14654,N_14265,N_14372);
nor U14655 (N_14655,N_14400,N_14475);
or U14656 (N_14656,N_14273,N_14413);
xor U14657 (N_14657,N_14460,N_14375);
xor U14658 (N_14658,N_14313,N_14428);
xor U14659 (N_14659,N_14301,N_14416);
or U14660 (N_14660,N_14386,N_14400);
nand U14661 (N_14661,N_14253,N_14491);
xor U14662 (N_14662,N_14260,N_14253);
and U14663 (N_14663,N_14373,N_14405);
and U14664 (N_14664,N_14452,N_14406);
nand U14665 (N_14665,N_14451,N_14466);
nor U14666 (N_14666,N_14283,N_14400);
nor U14667 (N_14667,N_14322,N_14418);
xnor U14668 (N_14668,N_14436,N_14302);
or U14669 (N_14669,N_14375,N_14326);
nand U14670 (N_14670,N_14273,N_14449);
and U14671 (N_14671,N_14256,N_14432);
xnor U14672 (N_14672,N_14429,N_14261);
xnor U14673 (N_14673,N_14419,N_14337);
xor U14674 (N_14674,N_14474,N_14481);
nor U14675 (N_14675,N_14472,N_14306);
nand U14676 (N_14676,N_14315,N_14310);
nor U14677 (N_14677,N_14352,N_14461);
and U14678 (N_14678,N_14432,N_14352);
nand U14679 (N_14679,N_14431,N_14261);
nand U14680 (N_14680,N_14267,N_14350);
nor U14681 (N_14681,N_14410,N_14478);
and U14682 (N_14682,N_14313,N_14282);
or U14683 (N_14683,N_14449,N_14426);
nand U14684 (N_14684,N_14252,N_14411);
or U14685 (N_14685,N_14332,N_14336);
nand U14686 (N_14686,N_14433,N_14364);
or U14687 (N_14687,N_14299,N_14481);
nand U14688 (N_14688,N_14455,N_14348);
or U14689 (N_14689,N_14334,N_14303);
nor U14690 (N_14690,N_14370,N_14287);
nand U14691 (N_14691,N_14452,N_14278);
nor U14692 (N_14692,N_14383,N_14496);
xor U14693 (N_14693,N_14359,N_14329);
nor U14694 (N_14694,N_14348,N_14432);
xor U14695 (N_14695,N_14270,N_14293);
nor U14696 (N_14696,N_14272,N_14444);
and U14697 (N_14697,N_14422,N_14259);
nand U14698 (N_14698,N_14486,N_14308);
nor U14699 (N_14699,N_14427,N_14280);
nand U14700 (N_14700,N_14350,N_14402);
or U14701 (N_14701,N_14460,N_14271);
nand U14702 (N_14702,N_14365,N_14286);
and U14703 (N_14703,N_14305,N_14291);
nor U14704 (N_14704,N_14343,N_14337);
nor U14705 (N_14705,N_14300,N_14458);
nor U14706 (N_14706,N_14296,N_14425);
nor U14707 (N_14707,N_14279,N_14304);
nand U14708 (N_14708,N_14350,N_14488);
xnor U14709 (N_14709,N_14308,N_14435);
nor U14710 (N_14710,N_14449,N_14320);
and U14711 (N_14711,N_14255,N_14395);
nand U14712 (N_14712,N_14476,N_14360);
or U14713 (N_14713,N_14471,N_14329);
nand U14714 (N_14714,N_14267,N_14473);
nor U14715 (N_14715,N_14303,N_14268);
or U14716 (N_14716,N_14287,N_14308);
nand U14717 (N_14717,N_14251,N_14338);
nand U14718 (N_14718,N_14425,N_14431);
xnor U14719 (N_14719,N_14347,N_14278);
and U14720 (N_14720,N_14445,N_14399);
xnor U14721 (N_14721,N_14337,N_14379);
and U14722 (N_14722,N_14430,N_14408);
nand U14723 (N_14723,N_14456,N_14495);
nand U14724 (N_14724,N_14496,N_14341);
nand U14725 (N_14725,N_14457,N_14423);
or U14726 (N_14726,N_14377,N_14421);
nand U14727 (N_14727,N_14326,N_14254);
and U14728 (N_14728,N_14250,N_14437);
nand U14729 (N_14729,N_14460,N_14265);
or U14730 (N_14730,N_14335,N_14396);
xor U14731 (N_14731,N_14303,N_14292);
and U14732 (N_14732,N_14314,N_14367);
or U14733 (N_14733,N_14479,N_14430);
nor U14734 (N_14734,N_14381,N_14284);
nand U14735 (N_14735,N_14422,N_14351);
and U14736 (N_14736,N_14280,N_14452);
and U14737 (N_14737,N_14407,N_14442);
xor U14738 (N_14738,N_14471,N_14265);
nor U14739 (N_14739,N_14417,N_14333);
and U14740 (N_14740,N_14472,N_14494);
and U14741 (N_14741,N_14388,N_14437);
nor U14742 (N_14742,N_14266,N_14453);
xnor U14743 (N_14743,N_14312,N_14269);
xnor U14744 (N_14744,N_14474,N_14465);
nand U14745 (N_14745,N_14497,N_14308);
or U14746 (N_14746,N_14400,N_14304);
or U14747 (N_14747,N_14469,N_14495);
and U14748 (N_14748,N_14442,N_14472);
or U14749 (N_14749,N_14304,N_14357);
or U14750 (N_14750,N_14596,N_14719);
or U14751 (N_14751,N_14743,N_14675);
nand U14752 (N_14752,N_14672,N_14604);
and U14753 (N_14753,N_14564,N_14576);
and U14754 (N_14754,N_14607,N_14640);
nand U14755 (N_14755,N_14630,N_14571);
or U14756 (N_14756,N_14600,N_14693);
xnor U14757 (N_14757,N_14637,N_14708);
xnor U14758 (N_14758,N_14540,N_14658);
or U14759 (N_14759,N_14507,N_14558);
xnor U14760 (N_14760,N_14639,N_14695);
xor U14761 (N_14761,N_14681,N_14522);
and U14762 (N_14762,N_14618,N_14673);
or U14763 (N_14763,N_14602,N_14668);
xnor U14764 (N_14764,N_14570,N_14539);
nor U14765 (N_14765,N_14704,N_14617);
and U14766 (N_14766,N_14710,N_14711);
nor U14767 (N_14767,N_14562,N_14520);
nand U14768 (N_14768,N_14557,N_14548);
nand U14769 (N_14769,N_14587,N_14651);
xor U14770 (N_14770,N_14531,N_14735);
nand U14771 (N_14771,N_14671,N_14578);
xor U14772 (N_14772,N_14688,N_14715);
or U14773 (N_14773,N_14720,N_14633);
nor U14774 (N_14774,N_14670,N_14638);
nor U14775 (N_14775,N_14556,N_14572);
nor U14776 (N_14776,N_14620,N_14510);
nor U14777 (N_14777,N_14549,N_14685);
nor U14778 (N_14778,N_14701,N_14598);
nor U14779 (N_14779,N_14629,N_14677);
nor U14780 (N_14780,N_14712,N_14736);
nand U14781 (N_14781,N_14729,N_14626);
and U14782 (N_14782,N_14666,N_14517);
nand U14783 (N_14783,N_14724,N_14608);
or U14784 (N_14784,N_14655,N_14749);
and U14785 (N_14785,N_14580,N_14742);
xor U14786 (N_14786,N_14547,N_14583);
nand U14787 (N_14787,N_14631,N_14527);
nand U14788 (N_14788,N_14663,N_14590);
nor U14789 (N_14789,N_14744,N_14678);
and U14790 (N_14790,N_14731,N_14702);
nor U14791 (N_14791,N_14727,N_14627);
or U14792 (N_14792,N_14709,N_14560);
nand U14793 (N_14793,N_14714,N_14676);
xor U14794 (N_14794,N_14559,N_14532);
nor U14795 (N_14795,N_14603,N_14732);
nand U14796 (N_14796,N_14519,N_14746);
and U14797 (N_14797,N_14725,N_14660);
nor U14798 (N_14798,N_14609,N_14504);
nor U14799 (N_14799,N_14533,N_14523);
nand U14800 (N_14800,N_14636,N_14707);
xor U14801 (N_14801,N_14705,N_14740);
and U14802 (N_14802,N_14619,N_14646);
nor U14803 (N_14803,N_14541,N_14722);
and U14804 (N_14804,N_14652,N_14664);
nand U14805 (N_14805,N_14573,N_14534);
and U14806 (N_14806,N_14593,N_14625);
and U14807 (N_14807,N_14544,N_14700);
nor U14808 (N_14808,N_14529,N_14659);
xnor U14809 (N_14809,N_14605,N_14622);
or U14810 (N_14810,N_14584,N_14542);
xnor U14811 (N_14811,N_14594,N_14551);
nor U14812 (N_14812,N_14657,N_14632);
or U14813 (N_14813,N_14643,N_14734);
or U14814 (N_14814,N_14610,N_14521);
or U14815 (N_14815,N_14500,N_14623);
and U14816 (N_14816,N_14661,N_14577);
or U14817 (N_14817,N_14690,N_14509);
nand U14818 (N_14818,N_14513,N_14545);
nand U14819 (N_14819,N_14574,N_14501);
or U14820 (N_14820,N_14595,N_14703);
or U14821 (N_14821,N_14716,N_14567);
nand U14822 (N_14822,N_14730,N_14667);
nor U14823 (N_14823,N_14505,N_14597);
xnor U14824 (N_14824,N_14699,N_14554);
nor U14825 (N_14825,N_14528,N_14514);
nand U14826 (N_14826,N_14615,N_14641);
or U14827 (N_14827,N_14745,N_14747);
or U14828 (N_14828,N_14679,N_14546);
and U14829 (N_14829,N_14726,N_14717);
xnor U14830 (N_14830,N_14535,N_14656);
nor U14831 (N_14831,N_14674,N_14516);
xnor U14832 (N_14832,N_14647,N_14582);
nor U14833 (N_14833,N_14662,N_14665);
nor U14834 (N_14834,N_14682,N_14624);
nor U14835 (N_14835,N_14586,N_14648);
xnor U14836 (N_14836,N_14599,N_14575);
xnor U14837 (N_14837,N_14524,N_14536);
or U14838 (N_14838,N_14686,N_14553);
or U14839 (N_14839,N_14669,N_14649);
and U14840 (N_14840,N_14691,N_14650);
nor U14841 (N_14841,N_14538,N_14739);
nand U14842 (N_14842,N_14621,N_14569);
nor U14843 (N_14843,N_14692,N_14697);
nor U14844 (N_14844,N_14728,N_14654);
xnor U14845 (N_14845,N_14680,N_14634);
xor U14846 (N_14846,N_14550,N_14644);
and U14847 (N_14847,N_14741,N_14684);
and U14848 (N_14848,N_14689,N_14585);
nand U14849 (N_14849,N_14694,N_14687);
and U14850 (N_14850,N_14738,N_14635);
nand U14851 (N_14851,N_14511,N_14698);
nor U14852 (N_14852,N_14506,N_14733);
nand U14853 (N_14853,N_14518,N_14612);
xnor U14854 (N_14854,N_14565,N_14579);
and U14855 (N_14855,N_14591,N_14723);
nand U14856 (N_14856,N_14526,N_14748);
and U14857 (N_14857,N_14616,N_14581);
xnor U14858 (N_14858,N_14601,N_14552);
nor U14859 (N_14859,N_14721,N_14589);
nand U14860 (N_14860,N_14530,N_14642);
xor U14861 (N_14861,N_14588,N_14696);
xor U14862 (N_14862,N_14592,N_14653);
nand U14863 (N_14863,N_14645,N_14628);
and U14864 (N_14864,N_14713,N_14563);
and U14865 (N_14865,N_14525,N_14537);
nand U14866 (N_14866,N_14555,N_14508);
xor U14867 (N_14867,N_14737,N_14614);
and U14868 (N_14868,N_14566,N_14502);
xnor U14869 (N_14869,N_14568,N_14706);
and U14870 (N_14870,N_14683,N_14611);
xnor U14871 (N_14871,N_14606,N_14561);
xor U14872 (N_14872,N_14718,N_14512);
and U14873 (N_14873,N_14503,N_14515);
and U14874 (N_14874,N_14543,N_14613);
nand U14875 (N_14875,N_14650,N_14741);
xor U14876 (N_14876,N_14743,N_14649);
nor U14877 (N_14877,N_14652,N_14506);
and U14878 (N_14878,N_14637,N_14615);
nor U14879 (N_14879,N_14634,N_14616);
and U14880 (N_14880,N_14525,N_14509);
nand U14881 (N_14881,N_14733,N_14581);
nor U14882 (N_14882,N_14587,N_14623);
and U14883 (N_14883,N_14709,N_14685);
nor U14884 (N_14884,N_14642,N_14506);
nand U14885 (N_14885,N_14613,N_14633);
xnor U14886 (N_14886,N_14646,N_14644);
nand U14887 (N_14887,N_14543,N_14682);
xnor U14888 (N_14888,N_14693,N_14591);
xnor U14889 (N_14889,N_14511,N_14516);
nand U14890 (N_14890,N_14529,N_14519);
nor U14891 (N_14891,N_14744,N_14501);
or U14892 (N_14892,N_14720,N_14670);
nor U14893 (N_14893,N_14555,N_14662);
nand U14894 (N_14894,N_14531,N_14580);
or U14895 (N_14895,N_14667,N_14678);
and U14896 (N_14896,N_14571,N_14642);
or U14897 (N_14897,N_14519,N_14634);
or U14898 (N_14898,N_14693,N_14725);
nor U14899 (N_14899,N_14657,N_14685);
nor U14900 (N_14900,N_14698,N_14520);
xor U14901 (N_14901,N_14568,N_14705);
xnor U14902 (N_14902,N_14543,N_14665);
nand U14903 (N_14903,N_14521,N_14665);
and U14904 (N_14904,N_14541,N_14531);
or U14905 (N_14905,N_14601,N_14500);
nand U14906 (N_14906,N_14543,N_14617);
nor U14907 (N_14907,N_14538,N_14733);
xor U14908 (N_14908,N_14540,N_14608);
nor U14909 (N_14909,N_14741,N_14703);
xnor U14910 (N_14910,N_14561,N_14740);
and U14911 (N_14911,N_14634,N_14746);
nor U14912 (N_14912,N_14639,N_14735);
nand U14913 (N_14913,N_14690,N_14502);
xor U14914 (N_14914,N_14644,N_14706);
or U14915 (N_14915,N_14540,N_14700);
nand U14916 (N_14916,N_14699,N_14646);
or U14917 (N_14917,N_14710,N_14598);
nor U14918 (N_14918,N_14707,N_14652);
xnor U14919 (N_14919,N_14657,N_14618);
or U14920 (N_14920,N_14528,N_14597);
and U14921 (N_14921,N_14556,N_14579);
or U14922 (N_14922,N_14560,N_14540);
and U14923 (N_14923,N_14622,N_14695);
nand U14924 (N_14924,N_14689,N_14642);
nand U14925 (N_14925,N_14635,N_14658);
xnor U14926 (N_14926,N_14696,N_14524);
and U14927 (N_14927,N_14730,N_14697);
nor U14928 (N_14928,N_14737,N_14736);
or U14929 (N_14929,N_14530,N_14588);
or U14930 (N_14930,N_14621,N_14736);
nor U14931 (N_14931,N_14574,N_14612);
or U14932 (N_14932,N_14562,N_14620);
nand U14933 (N_14933,N_14581,N_14519);
or U14934 (N_14934,N_14749,N_14513);
nand U14935 (N_14935,N_14658,N_14687);
and U14936 (N_14936,N_14601,N_14675);
and U14937 (N_14937,N_14688,N_14691);
or U14938 (N_14938,N_14642,N_14507);
nand U14939 (N_14939,N_14560,N_14686);
and U14940 (N_14940,N_14584,N_14626);
xnor U14941 (N_14941,N_14688,N_14716);
xnor U14942 (N_14942,N_14631,N_14504);
nand U14943 (N_14943,N_14550,N_14578);
and U14944 (N_14944,N_14655,N_14731);
and U14945 (N_14945,N_14537,N_14704);
and U14946 (N_14946,N_14682,N_14611);
nor U14947 (N_14947,N_14518,N_14600);
nor U14948 (N_14948,N_14513,N_14675);
nand U14949 (N_14949,N_14658,N_14741);
nor U14950 (N_14950,N_14616,N_14670);
xor U14951 (N_14951,N_14643,N_14732);
nor U14952 (N_14952,N_14607,N_14615);
and U14953 (N_14953,N_14719,N_14559);
and U14954 (N_14954,N_14748,N_14638);
nand U14955 (N_14955,N_14615,N_14683);
xor U14956 (N_14956,N_14636,N_14654);
nand U14957 (N_14957,N_14660,N_14502);
or U14958 (N_14958,N_14515,N_14661);
nand U14959 (N_14959,N_14748,N_14714);
or U14960 (N_14960,N_14686,N_14550);
nand U14961 (N_14961,N_14718,N_14539);
nand U14962 (N_14962,N_14720,N_14740);
and U14963 (N_14963,N_14736,N_14544);
and U14964 (N_14964,N_14631,N_14584);
or U14965 (N_14965,N_14657,N_14738);
and U14966 (N_14966,N_14746,N_14693);
nor U14967 (N_14967,N_14701,N_14541);
nor U14968 (N_14968,N_14667,N_14611);
nand U14969 (N_14969,N_14576,N_14726);
and U14970 (N_14970,N_14714,N_14582);
and U14971 (N_14971,N_14666,N_14532);
xnor U14972 (N_14972,N_14536,N_14749);
xnor U14973 (N_14973,N_14530,N_14616);
or U14974 (N_14974,N_14531,N_14542);
nor U14975 (N_14975,N_14579,N_14567);
nand U14976 (N_14976,N_14514,N_14559);
and U14977 (N_14977,N_14603,N_14581);
xor U14978 (N_14978,N_14623,N_14642);
xnor U14979 (N_14979,N_14700,N_14596);
xnor U14980 (N_14980,N_14558,N_14583);
or U14981 (N_14981,N_14667,N_14658);
nor U14982 (N_14982,N_14627,N_14529);
xor U14983 (N_14983,N_14550,N_14597);
nand U14984 (N_14984,N_14669,N_14547);
xor U14985 (N_14985,N_14596,N_14527);
or U14986 (N_14986,N_14514,N_14574);
and U14987 (N_14987,N_14722,N_14585);
nand U14988 (N_14988,N_14598,N_14528);
or U14989 (N_14989,N_14522,N_14546);
xnor U14990 (N_14990,N_14596,N_14546);
or U14991 (N_14991,N_14692,N_14587);
or U14992 (N_14992,N_14698,N_14587);
nor U14993 (N_14993,N_14660,N_14514);
or U14994 (N_14994,N_14616,N_14675);
nand U14995 (N_14995,N_14649,N_14594);
and U14996 (N_14996,N_14729,N_14602);
or U14997 (N_14997,N_14554,N_14681);
and U14998 (N_14998,N_14546,N_14508);
or U14999 (N_14999,N_14523,N_14687);
and U15000 (N_15000,N_14943,N_14920);
nand U15001 (N_15001,N_14839,N_14819);
nor U15002 (N_15002,N_14921,N_14838);
nand U15003 (N_15003,N_14836,N_14853);
xnor U15004 (N_15004,N_14926,N_14831);
xnor U15005 (N_15005,N_14843,N_14857);
nand U15006 (N_15006,N_14890,N_14905);
or U15007 (N_15007,N_14870,N_14881);
nor U15008 (N_15008,N_14766,N_14958);
and U15009 (N_15009,N_14820,N_14859);
nand U15010 (N_15010,N_14871,N_14752);
xnor U15011 (N_15011,N_14930,N_14841);
or U15012 (N_15012,N_14972,N_14848);
and U15013 (N_15013,N_14847,N_14882);
nand U15014 (N_15014,N_14975,N_14998);
or U15015 (N_15015,N_14783,N_14765);
nor U15016 (N_15016,N_14868,N_14751);
nand U15017 (N_15017,N_14812,N_14773);
or U15018 (N_15018,N_14824,N_14912);
nor U15019 (N_15019,N_14851,N_14984);
and U15020 (N_15020,N_14979,N_14767);
xor U15021 (N_15021,N_14821,N_14802);
or U15022 (N_15022,N_14761,N_14891);
nand U15023 (N_15023,N_14937,N_14777);
xnor U15024 (N_15024,N_14939,N_14988);
xnor U15025 (N_15025,N_14828,N_14915);
xor U15026 (N_15026,N_14902,N_14948);
xnor U15027 (N_15027,N_14807,N_14909);
nor U15028 (N_15028,N_14755,N_14946);
nand U15029 (N_15029,N_14840,N_14994);
and U15030 (N_15030,N_14918,N_14950);
nand U15031 (N_15031,N_14806,N_14794);
or U15032 (N_15032,N_14856,N_14827);
nor U15033 (N_15033,N_14753,N_14759);
nand U15034 (N_15034,N_14760,N_14981);
or U15035 (N_15035,N_14850,N_14814);
nor U15036 (N_15036,N_14957,N_14780);
or U15037 (N_15037,N_14858,N_14945);
xor U15038 (N_15038,N_14974,N_14833);
nor U15039 (N_15039,N_14865,N_14869);
or U15040 (N_15040,N_14788,N_14986);
xnor U15041 (N_15041,N_14883,N_14997);
xnor U15042 (N_15042,N_14795,N_14976);
xor U15043 (N_15043,N_14911,N_14875);
or U15044 (N_15044,N_14846,N_14892);
and U15045 (N_15045,N_14964,N_14770);
xor U15046 (N_15046,N_14786,N_14778);
and U15047 (N_15047,N_14886,N_14798);
or U15048 (N_15048,N_14774,N_14936);
nand U15049 (N_15049,N_14951,N_14811);
nand U15050 (N_15050,N_14923,N_14762);
nand U15051 (N_15051,N_14934,N_14860);
nand U15052 (N_15052,N_14989,N_14919);
xnor U15053 (N_15053,N_14913,N_14967);
xnor U15054 (N_15054,N_14944,N_14818);
or U15055 (N_15055,N_14849,N_14880);
xnor U15056 (N_15056,N_14901,N_14887);
nor U15057 (N_15057,N_14803,N_14985);
xor U15058 (N_15058,N_14970,N_14917);
xnor U15059 (N_15059,N_14845,N_14983);
nor U15060 (N_15060,N_14965,N_14900);
xnor U15061 (N_15061,N_14982,N_14942);
or U15062 (N_15062,N_14929,N_14854);
or U15063 (N_15063,N_14793,N_14897);
nand U15064 (N_15064,N_14935,N_14789);
xor U15065 (N_15065,N_14813,N_14792);
xnor U15066 (N_15066,N_14889,N_14888);
or U15067 (N_15067,N_14924,N_14823);
xor U15068 (N_15068,N_14885,N_14872);
xor U15069 (N_15069,N_14817,N_14916);
nor U15070 (N_15070,N_14782,N_14877);
xor U15071 (N_15071,N_14829,N_14835);
xor U15072 (N_15072,N_14757,N_14987);
nand U15073 (N_15073,N_14804,N_14878);
nor U15074 (N_15074,N_14977,N_14771);
nor U15075 (N_15075,N_14776,N_14784);
xnor U15076 (N_15076,N_14769,N_14775);
xor U15077 (N_15077,N_14953,N_14866);
and U15078 (N_15078,N_14933,N_14864);
and U15079 (N_15079,N_14893,N_14910);
and U15080 (N_15080,N_14922,N_14861);
or U15081 (N_15081,N_14973,N_14756);
nand U15082 (N_15082,N_14862,N_14928);
and U15083 (N_15083,N_14844,N_14808);
and U15084 (N_15084,N_14993,N_14990);
xnor U15085 (N_15085,N_14898,N_14907);
or U15086 (N_15086,N_14781,N_14855);
nor U15087 (N_15087,N_14876,N_14895);
nor U15088 (N_15088,N_14966,N_14927);
nand U15089 (N_15089,N_14852,N_14903);
nand U15090 (N_15090,N_14980,N_14894);
nor U15091 (N_15091,N_14932,N_14963);
or U15092 (N_15092,N_14992,N_14816);
xnor U15093 (N_15093,N_14805,N_14815);
or U15094 (N_15094,N_14940,N_14906);
or U15095 (N_15095,N_14768,N_14879);
nor U15096 (N_15096,N_14999,N_14954);
and U15097 (N_15097,N_14938,N_14949);
or U15098 (N_15098,N_14826,N_14863);
and U15099 (N_15099,N_14842,N_14908);
and U15100 (N_15100,N_14925,N_14790);
and U15101 (N_15101,N_14779,N_14764);
or U15102 (N_15102,N_14961,N_14968);
xor U15103 (N_15103,N_14796,N_14960);
or U15104 (N_15104,N_14810,N_14941);
and U15105 (N_15105,N_14754,N_14830);
nand U15106 (N_15106,N_14914,N_14947);
nand U15107 (N_15107,N_14899,N_14799);
or U15108 (N_15108,N_14772,N_14837);
nand U15109 (N_15109,N_14787,N_14969);
nor U15110 (N_15110,N_14959,N_14832);
or U15111 (N_15111,N_14971,N_14822);
or U15112 (N_15112,N_14931,N_14834);
xnor U15113 (N_15113,N_14791,N_14800);
nor U15114 (N_15114,N_14996,N_14955);
nor U15115 (N_15115,N_14873,N_14867);
or U15116 (N_15116,N_14758,N_14809);
nand U15117 (N_15117,N_14785,N_14962);
and U15118 (N_15118,N_14978,N_14995);
and U15119 (N_15119,N_14763,N_14991);
and U15120 (N_15120,N_14884,N_14801);
nand U15121 (N_15121,N_14952,N_14904);
and U15122 (N_15122,N_14956,N_14825);
nor U15123 (N_15123,N_14750,N_14896);
xnor U15124 (N_15124,N_14874,N_14797);
xnor U15125 (N_15125,N_14941,N_14815);
or U15126 (N_15126,N_14882,N_14980);
or U15127 (N_15127,N_14873,N_14929);
xnor U15128 (N_15128,N_14752,N_14829);
xor U15129 (N_15129,N_14873,N_14762);
nor U15130 (N_15130,N_14932,N_14937);
or U15131 (N_15131,N_14785,N_14793);
nand U15132 (N_15132,N_14997,N_14957);
and U15133 (N_15133,N_14769,N_14985);
xnor U15134 (N_15134,N_14962,N_14934);
nor U15135 (N_15135,N_14804,N_14783);
nor U15136 (N_15136,N_14796,N_14907);
nand U15137 (N_15137,N_14841,N_14820);
or U15138 (N_15138,N_14761,N_14967);
nor U15139 (N_15139,N_14783,N_14947);
nand U15140 (N_15140,N_14894,N_14952);
and U15141 (N_15141,N_14825,N_14936);
nor U15142 (N_15142,N_14894,N_14929);
xor U15143 (N_15143,N_14775,N_14888);
nand U15144 (N_15144,N_14876,N_14942);
or U15145 (N_15145,N_14750,N_14906);
and U15146 (N_15146,N_14774,N_14928);
nand U15147 (N_15147,N_14753,N_14905);
nor U15148 (N_15148,N_14767,N_14907);
xnor U15149 (N_15149,N_14981,N_14829);
and U15150 (N_15150,N_14757,N_14944);
and U15151 (N_15151,N_14929,N_14947);
and U15152 (N_15152,N_14894,N_14866);
and U15153 (N_15153,N_14802,N_14761);
and U15154 (N_15154,N_14852,N_14863);
xnor U15155 (N_15155,N_14842,N_14926);
nand U15156 (N_15156,N_14772,N_14828);
xor U15157 (N_15157,N_14954,N_14893);
xnor U15158 (N_15158,N_14825,N_14759);
nand U15159 (N_15159,N_14789,N_14923);
nor U15160 (N_15160,N_14882,N_14856);
or U15161 (N_15161,N_14953,N_14947);
and U15162 (N_15162,N_14796,N_14753);
nor U15163 (N_15163,N_14984,N_14921);
and U15164 (N_15164,N_14865,N_14812);
xnor U15165 (N_15165,N_14837,N_14824);
nor U15166 (N_15166,N_14795,N_14944);
xor U15167 (N_15167,N_14997,N_14814);
nand U15168 (N_15168,N_14785,N_14887);
or U15169 (N_15169,N_14951,N_14813);
nor U15170 (N_15170,N_14784,N_14936);
or U15171 (N_15171,N_14843,N_14914);
nor U15172 (N_15172,N_14967,N_14926);
xnor U15173 (N_15173,N_14934,N_14793);
or U15174 (N_15174,N_14889,N_14930);
or U15175 (N_15175,N_14786,N_14940);
or U15176 (N_15176,N_14927,N_14882);
and U15177 (N_15177,N_14991,N_14777);
nand U15178 (N_15178,N_14863,N_14832);
or U15179 (N_15179,N_14797,N_14804);
nand U15180 (N_15180,N_14948,N_14940);
nand U15181 (N_15181,N_14857,N_14856);
nand U15182 (N_15182,N_14836,N_14825);
nand U15183 (N_15183,N_14778,N_14768);
nand U15184 (N_15184,N_14772,N_14965);
nand U15185 (N_15185,N_14852,N_14810);
xnor U15186 (N_15186,N_14933,N_14983);
nor U15187 (N_15187,N_14982,N_14861);
nand U15188 (N_15188,N_14789,N_14879);
or U15189 (N_15189,N_14909,N_14785);
nor U15190 (N_15190,N_14970,N_14767);
and U15191 (N_15191,N_14866,N_14988);
nand U15192 (N_15192,N_14968,N_14882);
nor U15193 (N_15193,N_14841,N_14838);
nand U15194 (N_15194,N_14995,N_14894);
nor U15195 (N_15195,N_14808,N_14867);
and U15196 (N_15196,N_14857,N_14783);
nand U15197 (N_15197,N_14933,N_14884);
nand U15198 (N_15198,N_14907,N_14801);
nand U15199 (N_15199,N_14751,N_14925);
nand U15200 (N_15200,N_14853,N_14787);
or U15201 (N_15201,N_14997,N_14981);
nand U15202 (N_15202,N_14841,N_14789);
and U15203 (N_15203,N_14990,N_14849);
nor U15204 (N_15204,N_14996,N_14774);
nand U15205 (N_15205,N_14914,N_14877);
or U15206 (N_15206,N_14918,N_14920);
nor U15207 (N_15207,N_14904,N_14818);
or U15208 (N_15208,N_14970,N_14994);
xnor U15209 (N_15209,N_14989,N_14754);
or U15210 (N_15210,N_14856,N_14877);
or U15211 (N_15211,N_14989,N_14985);
or U15212 (N_15212,N_14967,N_14754);
nor U15213 (N_15213,N_14995,N_14945);
or U15214 (N_15214,N_14767,N_14866);
or U15215 (N_15215,N_14853,N_14848);
nand U15216 (N_15216,N_14814,N_14880);
xnor U15217 (N_15217,N_14807,N_14944);
and U15218 (N_15218,N_14952,N_14787);
or U15219 (N_15219,N_14914,N_14769);
nor U15220 (N_15220,N_14881,N_14958);
or U15221 (N_15221,N_14838,N_14850);
or U15222 (N_15222,N_14949,N_14958);
xor U15223 (N_15223,N_14916,N_14818);
nor U15224 (N_15224,N_14943,N_14785);
xor U15225 (N_15225,N_14769,N_14965);
nand U15226 (N_15226,N_14768,N_14900);
and U15227 (N_15227,N_14820,N_14801);
nor U15228 (N_15228,N_14945,N_14992);
and U15229 (N_15229,N_14973,N_14767);
or U15230 (N_15230,N_14983,N_14826);
nand U15231 (N_15231,N_14948,N_14819);
or U15232 (N_15232,N_14788,N_14864);
or U15233 (N_15233,N_14866,N_14781);
nand U15234 (N_15234,N_14809,N_14987);
or U15235 (N_15235,N_14960,N_14883);
nand U15236 (N_15236,N_14801,N_14978);
nor U15237 (N_15237,N_14921,N_14983);
or U15238 (N_15238,N_14810,N_14845);
or U15239 (N_15239,N_14842,N_14888);
and U15240 (N_15240,N_14799,N_14935);
xor U15241 (N_15241,N_14989,N_14758);
and U15242 (N_15242,N_14791,N_14837);
xor U15243 (N_15243,N_14897,N_14855);
and U15244 (N_15244,N_14899,N_14970);
or U15245 (N_15245,N_14917,N_14916);
xor U15246 (N_15246,N_14771,N_14964);
nor U15247 (N_15247,N_14922,N_14776);
nand U15248 (N_15248,N_14957,N_14896);
nand U15249 (N_15249,N_14898,N_14939);
nor U15250 (N_15250,N_15099,N_15193);
nor U15251 (N_15251,N_15164,N_15067);
nor U15252 (N_15252,N_15211,N_15033);
or U15253 (N_15253,N_15116,N_15079);
or U15254 (N_15254,N_15104,N_15108);
or U15255 (N_15255,N_15204,N_15012);
xnor U15256 (N_15256,N_15171,N_15072);
or U15257 (N_15257,N_15014,N_15201);
xor U15258 (N_15258,N_15063,N_15209);
and U15259 (N_15259,N_15162,N_15200);
nor U15260 (N_15260,N_15194,N_15028);
or U15261 (N_15261,N_15089,N_15221);
or U15262 (N_15262,N_15084,N_15032);
nand U15263 (N_15263,N_15149,N_15009);
nor U15264 (N_15264,N_15215,N_15167);
or U15265 (N_15265,N_15095,N_15154);
or U15266 (N_15266,N_15128,N_15127);
nor U15267 (N_15267,N_15216,N_15048);
or U15268 (N_15268,N_15055,N_15142);
and U15269 (N_15269,N_15006,N_15246);
xnor U15270 (N_15270,N_15073,N_15069);
or U15271 (N_15271,N_15096,N_15120);
nor U15272 (N_15272,N_15081,N_15231);
xnor U15273 (N_15273,N_15210,N_15126);
xnor U15274 (N_15274,N_15090,N_15035);
nand U15275 (N_15275,N_15051,N_15161);
nand U15276 (N_15276,N_15004,N_15034);
or U15277 (N_15277,N_15119,N_15043);
and U15278 (N_15278,N_15001,N_15183);
nand U15279 (N_15279,N_15042,N_15057);
xor U15280 (N_15280,N_15002,N_15065);
xor U15281 (N_15281,N_15085,N_15223);
nand U15282 (N_15282,N_15025,N_15172);
xor U15283 (N_15283,N_15036,N_15109);
and U15284 (N_15284,N_15179,N_15117);
nand U15285 (N_15285,N_15061,N_15180);
nand U15286 (N_15286,N_15207,N_15219);
or U15287 (N_15287,N_15236,N_15101);
nor U15288 (N_15288,N_15205,N_15198);
and U15289 (N_15289,N_15074,N_15160);
or U15290 (N_15290,N_15064,N_15019);
and U15291 (N_15291,N_15052,N_15011);
or U15292 (N_15292,N_15247,N_15112);
nand U15293 (N_15293,N_15082,N_15137);
xnor U15294 (N_15294,N_15232,N_15206);
xor U15295 (N_15295,N_15103,N_15233);
and U15296 (N_15296,N_15075,N_15047);
and U15297 (N_15297,N_15169,N_15058);
and U15298 (N_15298,N_15195,N_15097);
nor U15299 (N_15299,N_15187,N_15220);
nor U15300 (N_15300,N_15086,N_15145);
and U15301 (N_15301,N_15030,N_15023);
or U15302 (N_15302,N_15131,N_15111);
nand U15303 (N_15303,N_15044,N_15166);
nor U15304 (N_15304,N_15024,N_15045);
and U15305 (N_15305,N_15100,N_15088);
nand U15306 (N_15306,N_15174,N_15182);
nand U15307 (N_15307,N_15078,N_15240);
nand U15308 (N_15308,N_15152,N_15000);
and U15309 (N_15309,N_15225,N_15054);
xnor U15310 (N_15310,N_15184,N_15018);
nand U15311 (N_15311,N_15015,N_15071);
nor U15312 (N_15312,N_15199,N_15170);
or U15313 (N_15313,N_15141,N_15202);
or U15314 (N_15314,N_15053,N_15062);
xor U15315 (N_15315,N_15155,N_15114);
or U15316 (N_15316,N_15189,N_15157);
and U15317 (N_15317,N_15020,N_15050);
or U15318 (N_15318,N_15230,N_15245);
nand U15319 (N_15319,N_15242,N_15005);
and U15320 (N_15320,N_15178,N_15159);
or U15321 (N_15321,N_15106,N_15177);
nand U15322 (N_15322,N_15234,N_15016);
and U15323 (N_15323,N_15008,N_15091);
or U15324 (N_15324,N_15049,N_15191);
xnor U15325 (N_15325,N_15070,N_15241);
xor U15326 (N_15326,N_15176,N_15129);
nand U15327 (N_15327,N_15229,N_15188);
and U15328 (N_15328,N_15144,N_15046);
nor U15329 (N_15329,N_15094,N_15124);
xnor U15330 (N_15330,N_15003,N_15163);
xnor U15331 (N_15331,N_15228,N_15010);
nor U15332 (N_15332,N_15158,N_15186);
nor U15333 (N_15333,N_15113,N_15203);
nor U15334 (N_15334,N_15227,N_15041);
nor U15335 (N_15335,N_15139,N_15037);
or U15336 (N_15336,N_15118,N_15248);
nor U15337 (N_15337,N_15098,N_15123);
and U15338 (N_15338,N_15066,N_15092);
nand U15339 (N_15339,N_15132,N_15192);
and U15340 (N_15340,N_15105,N_15208);
nand U15341 (N_15341,N_15143,N_15235);
nand U15342 (N_15342,N_15238,N_15196);
xor U15343 (N_15343,N_15068,N_15217);
nor U15344 (N_15344,N_15115,N_15244);
nand U15345 (N_15345,N_15181,N_15022);
or U15346 (N_15346,N_15107,N_15039);
xnor U15347 (N_15347,N_15213,N_15165);
nand U15348 (N_15348,N_15185,N_15239);
nand U15349 (N_15349,N_15168,N_15007);
or U15350 (N_15350,N_15110,N_15121);
nor U15351 (N_15351,N_15130,N_15146);
xor U15352 (N_15352,N_15151,N_15021);
and U15353 (N_15353,N_15083,N_15237);
or U15354 (N_15354,N_15197,N_15138);
nand U15355 (N_15355,N_15102,N_15013);
nand U15356 (N_15356,N_15150,N_15218);
nor U15357 (N_15357,N_15249,N_15134);
nor U15358 (N_15358,N_15147,N_15135);
xor U15359 (N_15359,N_15214,N_15038);
nor U15360 (N_15360,N_15026,N_15060);
or U15361 (N_15361,N_15156,N_15029);
nor U15362 (N_15362,N_15076,N_15173);
xnor U15363 (N_15363,N_15027,N_15226);
xor U15364 (N_15364,N_15077,N_15031);
or U15365 (N_15365,N_15222,N_15212);
nor U15366 (N_15366,N_15133,N_15153);
and U15367 (N_15367,N_15140,N_15080);
and U15368 (N_15368,N_15040,N_15136);
nand U15369 (N_15369,N_15148,N_15224);
nand U15370 (N_15370,N_15093,N_15190);
nor U15371 (N_15371,N_15056,N_15017);
xnor U15372 (N_15372,N_15087,N_15059);
xor U15373 (N_15373,N_15243,N_15125);
nor U15374 (N_15374,N_15175,N_15122);
and U15375 (N_15375,N_15229,N_15165);
and U15376 (N_15376,N_15095,N_15054);
and U15377 (N_15377,N_15153,N_15119);
xnor U15378 (N_15378,N_15189,N_15121);
or U15379 (N_15379,N_15217,N_15211);
or U15380 (N_15380,N_15220,N_15233);
or U15381 (N_15381,N_15245,N_15048);
xnor U15382 (N_15382,N_15213,N_15164);
nor U15383 (N_15383,N_15194,N_15165);
or U15384 (N_15384,N_15209,N_15170);
nor U15385 (N_15385,N_15099,N_15051);
nor U15386 (N_15386,N_15007,N_15054);
nor U15387 (N_15387,N_15057,N_15235);
nand U15388 (N_15388,N_15219,N_15241);
nand U15389 (N_15389,N_15090,N_15022);
or U15390 (N_15390,N_15111,N_15108);
nand U15391 (N_15391,N_15136,N_15007);
or U15392 (N_15392,N_15007,N_15069);
and U15393 (N_15393,N_15118,N_15082);
or U15394 (N_15394,N_15089,N_15108);
and U15395 (N_15395,N_15035,N_15149);
nand U15396 (N_15396,N_15157,N_15053);
nand U15397 (N_15397,N_15006,N_15156);
xor U15398 (N_15398,N_15203,N_15035);
nand U15399 (N_15399,N_15239,N_15091);
nor U15400 (N_15400,N_15146,N_15248);
xor U15401 (N_15401,N_15089,N_15036);
or U15402 (N_15402,N_15225,N_15019);
or U15403 (N_15403,N_15060,N_15209);
nor U15404 (N_15404,N_15239,N_15111);
and U15405 (N_15405,N_15136,N_15132);
xor U15406 (N_15406,N_15201,N_15077);
and U15407 (N_15407,N_15140,N_15192);
and U15408 (N_15408,N_15183,N_15230);
nand U15409 (N_15409,N_15140,N_15166);
xor U15410 (N_15410,N_15173,N_15136);
nor U15411 (N_15411,N_15018,N_15202);
or U15412 (N_15412,N_15218,N_15221);
nor U15413 (N_15413,N_15190,N_15096);
nor U15414 (N_15414,N_15013,N_15115);
xor U15415 (N_15415,N_15079,N_15150);
and U15416 (N_15416,N_15075,N_15054);
and U15417 (N_15417,N_15019,N_15081);
and U15418 (N_15418,N_15185,N_15034);
nor U15419 (N_15419,N_15242,N_15121);
xnor U15420 (N_15420,N_15003,N_15114);
or U15421 (N_15421,N_15033,N_15037);
nand U15422 (N_15422,N_15051,N_15072);
or U15423 (N_15423,N_15203,N_15026);
xor U15424 (N_15424,N_15085,N_15114);
and U15425 (N_15425,N_15046,N_15174);
nand U15426 (N_15426,N_15157,N_15194);
nor U15427 (N_15427,N_15196,N_15246);
nand U15428 (N_15428,N_15000,N_15249);
or U15429 (N_15429,N_15099,N_15149);
xnor U15430 (N_15430,N_15202,N_15231);
xnor U15431 (N_15431,N_15070,N_15034);
xor U15432 (N_15432,N_15184,N_15062);
and U15433 (N_15433,N_15121,N_15205);
nor U15434 (N_15434,N_15070,N_15233);
nor U15435 (N_15435,N_15032,N_15005);
nand U15436 (N_15436,N_15207,N_15222);
and U15437 (N_15437,N_15207,N_15183);
xor U15438 (N_15438,N_15111,N_15119);
and U15439 (N_15439,N_15172,N_15036);
and U15440 (N_15440,N_15002,N_15025);
and U15441 (N_15441,N_15137,N_15180);
nand U15442 (N_15442,N_15143,N_15151);
nand U15443 (N_15443,N_15230,N_15000);
or U15444 (N_15444,N_15162,N_15058);
xnor U15445 (N_15445,N_15076,N_15080);
or U15446 (N_15446,N_15228,N_15214);
and U15447 (N_15447,N_15183,N_15095);
nand U15448 (N_15448,N_15062,N_15205);
nor U15449 (N_15449,N_15119,N_15100);
xor U15450 (N_15450,N_15130,N_15161);
xnor U15451 (N_15451,N_15022,N_15242);
nand U15452 (N_15452,N_15121,N_15160);
nor U15453 (N_15453,N_15231,N_15219);
nor U15454 (N_15454,N_15085,N_15060);
and U15455 (N_15455,N_15180,N_15186);
or U15456 (N_15456,N_15159,N_15067);
nor U15457 (N_15457,N_15128,N_15016);
or U15458 (N_15458,N_15148,N_15183);
and U15459 (N_15459,N_15182,N_15193);
xnor U15460 (N_15460,N_15073,N_15244);
nand U15461 (N_15461,N_15194,N_15024);
xnor U15462 (N_15462,N_15091,N_15138);
or U15463 (N_15463,N_15212,N_15126);
or U15464 (N_15464,N_15096,N_15032);
xor U15465 (N_15465,N_15127,N_15075);
nor U15466 (N_15466,N_15242,N_15054);
or U15467 (N_15467,N_15021,N_15215);
nor U15468 (N_15468,N_15176,N_15108);
or U15469 (N_15469,N_15203,N_15079);
xor U15470 (N_15470,N_15079,N_15051);
nor U15471 (N_15471,N_15057,N_15006);
nand U15472 (N_15472,N_15117,N_15146);
nor U15473 (N_15473,N_15079,N_15194);
nor U15474 (N_15474,N_15233,N_15120);
nor U15475 (N_15475,N_15025,N_15189);
nand U15476 (N_15476,N_15065,N_15102);
nand U15477 (N_15477,N_15231,N_15192);
and U15478 (N_15478,N_15045,N_15003);
xor U15479 (N_15479,N_15035,N_15014);
xor U15480 (N_15480,N_15245,N_15196);
and U15481 (N_15481,N_15032,N_15033);
or U15482 (N_15482,N_15196,N_15019);
and U15483 (N_15483,N_15041,N_15068);
nor U15484 (N_15484,N_15086,N_15021);
or U15485 (N_15485,N_15136,N_15201);
nand U15486 (N_15486,N_15006,N_15083);
xor U15487 (N_15487,N_15212,N_15225);
nor U15488 (N_15488,N_15159,N_15016);
xor U15489 (N_15489,N_15058,N_15051);
nor U15490 (N_15490,N_15004,N_15202);
and U15491 (N_15491,N_15058,N_15153);
nand U15492 (N_15492,N_15232,N_15095);
nor U15493 (N_15493,N_15199,N_15066);
xnor U15494 (N_15494,N_15238,N_15045);
or U15495 (N_15495,N_15105,N_15146);
xor U15496 (N_15496,N_15245,N_15121);
and U15497 (N_15497,N_15103,N_15232);
xor U15498 (N_15498,N_15025,N_15232);
nand U15499 (N_15499,N_15052,N_15128);
and U15500 (N_15500,N_15303,N_15319);
or U15501 (N_15501,N_15496,N_15487);
nand U15502 (N_15502,N_15264,N_15464);
or U15503 (N_15503,N_15331,N_15291);
and U15504 (N_15504,N_15397,N_15390);
and U15505 (N_15505,N_15419,N_15306);
nor U15506 (N_15506,N_15418,N_15386);
and U15507 (N_15507,N_15268,N_15295);
nand U15508 (N_15508,N_15337,N_15346);
or U15509 (N_15509,N_15254,N_15339);
nand U15510 (N_15510,N_15326,N_15356);
nor U15511 (N_15511,N_15357,N_15336);
nand U15512 (N_15512,N_15412,N_15282);
or U15513 (N_15513,N_15494,N_15408);
and U15514 (N_15514,N_15279,N_15313);
and U15515 (N_15515,N_15424,N_15352);
xnor U15516 (N_15516,N_15422,N_15348);
or U15517 (N_15517,N_15455,N_15258);
nand U15518 (N_15518,N_15314,N_15385);
or U15519 (N_15519,N_15406,N_15344);
nor U15520 (N_15520,N_15370,N_15304);
and U15521 (N_15521,N_15469,N_15456);
or U15522 (N_15522,N_15353,N_15471);
nand U15523 (N_15523,N_15444,N_15489);
and U15524 (N_15524,N_15465,N_15498);
nand U15525 (N_15525,N_15350,N_15287);
nor U15526 (N_15526,N_15286,N_15332);
nor U15527 (N_15527,N_15476,N_15269);
and U15528 (N_15528,N_15460,N_15318);
nand U15529 (N_15529,N_15328,N_15363);
and U15530 (N_15530,N_15420,N_15367);
or U15531 (N_15531,N_15392,N_15273);
nand U15532 (N_15532,N_15265,N_15461);
nand U15533 (N_15533,N_15395,N_15492);
nand U15534 (N_15534,N_15333,N_15340);
nand U15535 (N_15535,N_15393,N_15470);
xnor U15536 (N_15536,N_15414,N_15296);
nand U15537 (N_15537,N_15473,N_15480);
or U15538 (N_15538,N_15443,N_15371);
or U15539 (N_15539,N_15377,N_15302);
and U15540 (N_15540,N_15477,N_15285);
xnor U15541 (N_15541,N_15366,N_15283);
nor U15542 (N_15542,N_15447,N_15369);
or U15543 (N_15543,N_15301,N_15361);
and U15544 (N_15544,N_15467,N_15468);
and U15545 (N_15545,N_15310,N_15440);
nor U15546 (N_15546,N_15458,N_15288);
and U15547 (N_15547,N_15450,N_15497);
nand U15548 (N_15548,N_15441,N_15488);
nor U15549 (N_15549,N_15376,N_15409);
xor U15550 (N_15550,N_15427,N_15449);
or U15551 (N_15551,N_15278,N_15275);
nor U15552 (N_15552,N_15391,N_15266);
and U15553 (N_15553,N_15325,N_15297);
nand U15554 (N_15554,N_15415,N_15445);
xnor U15555 (N_15555,N_15410,N_15342);
and U15556 (N_15556,N_15430,N_15413);
or U15557 (N_15557,N_15389,N_15388);
or U15558 (N_15558,N_15439,N_15423);
nand U15559 (N_15559,N_15431,N_15429);
and U15560 (N_15560,N_15250,N_15323);
nand U15561 (N_15561,N_15490,N_15425);
nand U15562 (N_15562,N_15405,N_15387);
nand U15563 (N_15563,N_15478,N_15378);
or U15564 (N_15564,N_15479,N_15454);
and U15565 (N_15565,N_15475,N_15316);
or U15566 (N_15566,N_15417,N_15358);
nor U15567 (N_15567,N_15483,N_15421);
nor U15568 (N_15568,N_15432,N_15491);
and U15569 (N_15569,N_15463,N_15485);
and U15570 (N_15570,N_15267,N_15394);
or U15571 (N_15571,N_15320,N_15398);
nand U15572 (N_15572,N_15403,N_15355);
nor U15573 (N_15573,N_15374,N_15372);
and U15574 (N_15574,N_15277,N_15298);
and U15575 (N_15575,N_15472,N_15349);
and U15576 (N_15576,N_15338,N_15334);
nand U15577 (N_15577,N_15311,N_15402);
nor U15578 (N_15578,N_15255,N_15442);
nor U15579 (N_15579,N_15299,N_15257);
and U15580 (N_15580,N_15309,N_15292);
and U15581 (N_15581,N_15452,N_15459);
or U15582 (N_15582,N_15308,N_15384);
or U15583 (N_15583,N_15271,N_15457);
nor U15584 (N_15584,N_15434,N_15274);
and U15585 (N_15585,N_15321,N_15379);
xnor U15586 (N_15586,N_15411,N_15484);
or U15587 (N_15587,N_15252,N_15347);
and U15588 (N_15588,N_15466,N_15373);
and U15589 (N_15589,N_15307,N_15294);
nand U15590 (N_15590,N_15359,N_15253);
xnor U15591 (N_15591,N_15380,N_15446);
nand U15592 (N_15592,N_15474,N_15451);
nand U15593 (N_15593,N_15284,N_15407);
xor U15594 (N_15594,N_15399,N_15251);
nor U15595 (N_15595,N_15435,N_15453);
nand U15596 (N_15596,N_15341,N_15263);
nand U15597 (N_15597,N_15260,N_15482);
nor U15598 (N_15598,N_15400,N_15322);
nor U15599 (N_15599,N_15280,N_15259);
nor U15600 (N_15600,N_15261,N_15272);
nor U15601 (N_15601,N_15300,N_15416);
nand U15602 (N_15602,N_15428,N_15462);
and U15603 (N_15603,N_15486,N_15312);
xnor U15604 (N_15604,N_15329,N_15493);
nand U15605 (N_15605,N_15436,N_15354);
nor U15606 (N_15606,N_15433,N_15383);
or U15607 (N_15607,N_15290,N_15437);
and U15608 (N_15608,N_15360,N_15293);
and U15609 (N_15609,N_15324,N_15343);
and U15610 (N_15610,N_15481,N_15381);
nor U15611 (N_15611,N_15375,N_15276);
nor U15612 (N_15612,N_15305,N_15396);
nor U15613 (N_15613,N_15330,N_15448);
or U15614 (N_15614,N_15262,N_15317);
nand U15615 (N_15615,N_15362,N_15382);
nand U15616 (N_15616,N_15327,N_15351);
xnor U15617 (N_15617,N_15270,N_15281);
and U15618 (N_15618,N_15315,N_15368);
nor U15619 (N_15619,N_15345,N_15256);
and U15620 (N_15620,N_15426,N_15499);
xor U15621 (N_15621,N_15335,N_15404);
xnor U15622 (N_15622,N_15289,N_15401);
and U15623 (N_15623,N_15495,N_15438);
or U15624 (N_15624,N_15365,N_15364);
nor U15625 (N_15625,N_15488,N_15397);
nand U15626 (N_15626,N_15345,N_15351);
and U15627 (N_15627,N_15436,N_15251);
nand U15628 (N_15628,N_15301,N_15297);
and U15629 (N_15629,N_15359,N_15456);
nor U15630 (N_15630,N_15484,N_15264);
or U15631 (N_15631,N_15499,N_15346);
nor U15632 (N_15632,N_15284,N_15487);
xor U15633 (N_15633,N_15463,N_15375);
xor U15634 (N_15634,N_15483,N_15405);
nand U15635 (N_15635,N_15306,N_15274);
and U15636 (N_15636,N_15376,N_15286);
nand U15637 (N_15637,N_15360,N_15434);
xor U15638 (N_15638,N_15307,N_15458);
xor U15639 (N_15639,N_15416,N_15458);
nor U15640 (N_15640,N_15276,N_15313);
nor U15641 (N_15641,N_15445,N_15325);
nand U15642 (N_15642,N_15418,N_15421);
nand U15643 (N_15643,N_15411,N_15261);
and U15644 (N_15644,N_15407,N_15381);
nand U15645 (N_15645,N_15408,N_15437);
nor U15646 (N_15646,N_15382,N_15263);
nand U15647 (N_15647,N_15498,N_15488);
nor U15648 (N_15648,N_15283,N_15488);
or U15649 (N_15649,N_15257,N_15432);
nor U15650 (N_15650,N_15379,N_15344);
and U15651 (N_15651,N_15419,N_15468);
nand U15652 (N_15652,N_15275,N_15259);
or U15653 (N_15653,N_15419,N_15445);
nor U15654 (N_15654,N_15261,N_15371);
nand U15655 (N_15655,N_15430,N_15434);
xor U15656 (N_15656,N_15376,N_15471);
or U15657 (N_15657,N_15321,N_15353);
nor U15658 (N_15658,N_15417,N_15455);
or U15659 (N_15659,N_15270,N_15271);
nand U15660 (N_15660,N_15391,N_15397);
nor U15661 (N_15661,N_15492,N_15268);
or U15662 (N_15662,N_15417,N_15457);
nand U15663 (N_15663,N_15298,N_15352);
and U15664 (N_15664,N_15319,N_15343);
or U15665 (N_15665,N_15312,N_15308);
nor U15666 (N_15666,N_15450,N_15291);
xor U15667 (N_15667,N_15474,N_15311);
xor U15668 (N_15668,N_15388,N_15292);
nor U15669 (N_15669,N_15330,N_15350);
xnor U15670 (N_15670,N_15470,N_15282);
and U15671 (N_15671,N_15409,N_15466);
or U15672 (N_15672,N_15293,N_15440);
nand U15673 (N_15673,N_15389,N_15298);
and U15674 (N_15674,N_15382,N_15325);
and U15675 (N_15675,N_15308,N_15428);
nand U15676 (N_15676,N_15374,N_15323);
and U15677 (N_15677,N_15490,N_15355);
nand U15678 (N_15678,N_15335,N_15338);
nand U15679 (N_15679,N_15338,N_15395);
xnor U15680 (N_15680,N_15455,N_15437);
or U15681 (N_15681,N_15328,N_15479);
xnor U15682 (N_15682,N_15259,N_15493);
xnor U15683 (N_15683,N_15321,N_15260);
or U15684 (N_15684,N_15370,N_15368);
xor U15685 (N_15685,N_15351,N_15433);
nor U15686 (N_15686,N_15324,N_15435);
xnor U15687 (N_15687,N_15449,N_15417);
nand U15688 (N_15688,N_15314,N_15498);
nor U15689 (N_15689,N_15289,N_15355);
nand U15690 (N_15690,N_15266,N_15300);
nand U15691 (N_15691,N_15397,N_15445);
and U15692 (N_15692,N_15356,N_15423);
and U15693 (N_15693,N_15428,N_15418);
or U15694 (N_15694,N_15386,N_15254);
nand U15695 (N_15695,N_15259,N_15361);
xnor U15696 (N_15696,N_15387,N_15491);
nand U15697 (N_15697,N_15406,N_15416);
nand U15698 (N_15698,N_15458,N_15443);
nor U15699 (N_15699,N_15364,N_15251);
xor U15700 (N_15700,N_15362,N_15292);
xor U15701 (N_15701,N_15416,N_15334);
nand U15702 (N_15702,N_15466,N_15390);
or U15703 (N_15703,N_15298,N_15319);
and U15704 (N_15704,N_15488,N_15334);
nor U15705 (N_15705,N_15474,N_15456);
nand U15706 (N_15706,N_15294,N_15383);
xnor U15707 (N_15707,N_15338,N_15461);
or U15708 (N_15708,N_15459,N_15422);
and U15709 (N_15709,N_15371,N_15480);
or U15710 (N_15710,N_15380,N_15475);
xor U15711 (N_15711,N_15412,N_15380);
or U15712 (N_15712,N_15412,N_15498);
nor U15713 (N_15713,N_15475,N_15279);
nor U15714 (N_15714,N_15369,N_15376);
xor U15715 (N_15715,N_15307,N_15456);
nor U15716 (N_15716,N_15393,N_15305);
nand U15717 (N_15717,N_15428,N_15250);
nand U15718 (N_15718,N_15438,N_15346);
nand U15719 (N_15719,N_15376,N_15343);
or U15720 (N_15720,N_15455,N_15255);
and U15721 (N_15721,N_15358,N_15388);
nor U15722 (N_15722,N_15489,N_15289);
xor U15723 (N_15723,N_15464,N_15287);
nor U15724 (N_15724,N_15272,N_15370);
or U15725 (N_15725,N_15474,N_15418);
xnor U15726 (N_15726,N_15400,N_15353);
and U15727 (N_15727,N_15297,N_15421);
xnor U15728 (N_15728,N_15496,N_15488);
xnor U15729 (N_15729,N_15288,N_15388);
xor U15730 (N_15730,N_15433,N_15361);
xor U15731 (N_15731,N_15421,N_15250);
and U15732 (N_15732,N_15341,N_15343);
and U15733 (N_15733,N_15390,N_15451);
and U15734 (N_15734,N_15475,N_15273);
nand U15735 (N_15735,N_15295,N_15301);
nand U15736 (N_15736,N_15418,N_15494);
nand U15737 (N_15737,N_15324,N_15281);
nand U15738 (N_15738,N_15297,N_15327);
nand U15739 (N_15739,N_15398,N_15258);
nand U15740 (N_15740,N_15270,N_15434);
nor U15741 (N_15741,N_15449,N_15287);
and U15742 (N_15742,N_15367,N_15269);
or U15743 (N_15743,N_15372,N_15352);
nor U15744 (N_15744,N_15422,N_15377);
xnor U15745 (N_15745,N_15461,N_15469);
or U15746 (N_15746,N_15322,N_15333);
or U15747 (N_15747,N_15424,N_15411);
nor U15748 (N_15748,N_15318,N_15262);
and U15749 (N_15749,N_15255,N_15279);
and U15750 (N_15750,N_15534,N_15697);
nand U15751 (N_15751,N_15510,N_15587);
xnor U15752 (N_15752,N_15689,N_15664);
nor U15753 (N_15753,N_15521,N_15725);
or U15754 (N_15754,N_15729,N_15734);
xnor U15755 (N_15755,N_15609,N_15677);
and U15756 (N_15756,N_15512,N_15706);
and U15757 (N_15757,N_15552,N_15633);
nor U15758 (N_15758,N_15730,N_15508);
nand U15759 (N_15759,N_15567,N_15568);
or U15760 (N_15760,N_15631,N_15716);
nor U15761 (N_15761,N_15577,N_15747);
and U15762 (N_15762,N_15583,N_15678);
xnor U15763 (N_15763,N_15647,N_15711);
nor U15764 (N_15764,N_15603,N_15691);
or U15765 (N_15765,N_15586,N_15606);
nand U15766 (N_15766,N_15565,N_15721);
nor U15767 (N_15767,N_15524,N_15511);
nor U15768 (N_15768,N_15671,N_15654);
nor U15769 (N_15769,N_15544,N_15522);
nor U15770 (N_15770,N_15621,N_15741);
xnor U15771 (N_15771,N_15722,N_15723);
or U15772 (N_15772,N_15748,N_15597);
nor U15773 (N_15773,N_15739,N_15728);
or U15774 (N_15774,N_15690,N_15638);
or U15775 (N_15775,N_15529,N_15500);
nand U15776 (N_15776,N_15736,N_15648);
or U15777 (N_15777,N_15708,N_15559);
and U15778 (N_15778,N_15607,N_15662);
nor U15779 (N_15779,N_15669,N_15514);
and U15780 (N_15780,N_15566,N_15573);
xor U15781 (N_15781,N_15602,N_15718);
and U15782 (N_15782,N_15657,N_15539);
and U15783 (N_15783,N_15712,N_15526);
nor U15784 (N_15784,N_15554,N_15640);
and U15785 (N_15785,N_15555,N_15720);
nand U15786 (N_15786,N_15695,N_15639);
nor U15787 (N_15787,N_15692,N_15724);
nand U15788 (N_15788,N_15737,N_15744);
xnor U15789 (N_15789,N_15746,N_15742);
or U15790 (N_15790,N_15507,N_15649);
and U15791 (N_15791,N_15513,N_15593);
and U15792 (N_15792,N_15674,N_15580);
or U15793 (N_15793,N_15656,N_15731);
nor U15794 (N_15794,N_15541,N_15591);
and U15795 (N_15795,N_15642,N_15619);
and U15796 (N_15796,N_15616,N_15509);
nand U15797 (N_15797,N_15704,N_15743);
xor U15798 (N_15798,N_15681,N_15715);
or U15799 (N_15799,N_15628,N_15661);
xnor U15800 (N_15800,N_15658,N_15643);
and U15801 (N_15801,N_15545,N_15667);
and U15802 (N_15802,N_15668,N_15575);
nand U15803 (N_15803,N_15564,N_15523);
nand U15804 (N_15804,N_15733,N_15663);
xor U15805 (N_15805,N_15738,N_15687);
xnor U15806 (N_15806,N_15740,N_15613);
nand U15807 (N_15807,N_15683,N_15634);
and U15808 (N_15808,N_15680,N_15506);
nor U15809 (N_15809,N_15735,N_15536);
xor U15810 (N_15810,N_15703,N_15605);
nand U15811 (N_15811,N_15629,N_15531);
and U15812 (N_15812,N_15726,N_15614);
or U15813 (N_15813,N_15732,N_15682);
xor U15814 (N_15814,N_15625,N_15581);
or U15815 (N_15815,N_15557,N_15652);
nor U15816 (N_15816,N_15561,N_15540);
or U15817 (N_15817,N_15645,N_15572);
or U15818 (N_15818,N_15543,N_15717);
and U15819 (N_15819,N_15562,N_15701);
and U15820 (N_15820,N_15626,N_15713);
xor U15821 (N_15821,N_15705,N_15535);
or U15822 (N_15822,N_15502,N_15556);
nor U15823 (N_15823,N_15653,N_15595);
nor U15824 (N_15824,N_15574,N_15636);
and U15825 (N_15825,N_15599,N_15659);
or U15826 (N_15826,N_15630,N_15578);
or U15827 (N_15827,N_15660,N_15589);
and U15828 (N_15828,N_15655,N_15612);
and U15829 (N_15829,N_15505,N_15688);
and U15830 (N_15830,N_15624,N_15579);
or U15831 (N_15831,N_15617,N_15501);
and U15832 (N_15832,N_15623,N_15611);
nor U15833 (N_15833,N_15503,N_15622);
nor U15834 (N_15834,N_15596,N_15699);
xor U15835 (N_15835,N_15601,N_15582);
or U15836 (N_15836,N_15528,N_15585);
xor U15837 (N_15837,N_15694,N_15650);
nor U15838 (N_15838,N_15515,N_15673);
or U15839 (N_15839,N_15530,N_15641);
xor U15840 (N_15840,N_15698,N_15686);
and U15841 (N_15841,N_15666,N_15672);
and U15842 (N_15842,N_15651,N_15533);
and U15843 (N_15843,N_15676,N_15538);
nor U15844 (N_15844,N_15707,N_15570);
xor U15845 (N_15845,N_15569,N_15714);
and U15846 (N_15846,N_15675,N_15504);
xnor U15847 (N_15847,N_15588,N_15550);
and U15848 (N_15848,N_15558,N_15745);
and U15849 (N_15849,N_15632,N_15685);
nand U15850 (N_15850,N_15679,N_15563);
nor U15851 (N_15851,N_15670,N_15610);
nor U15852 (N_15852,N_15537,N_15527);
nand U15853 (N_15853,N_15542,N_15546);
xor U15854 (N_15854,N_15620,N_15598);
and U15855 (N_15855,N_15684,N_15519);
and U15856 (N_15856,N_15560,N_15576);
or U15857 (N_15857,N_15719,N_15604);
or U15858 (N_15858,N_15749,N_15600);
nor U15859 (N_15859,N_15644,N_15627);
and U15860 (N_15860,N_15517,N_15635);
and U15861 (N_15861,N_15553,N_15608);
xor U15862 (N_15862,N_15693,N_15516);
nand U15863 (N_15863,N_15727,N_15551);
and U15864 (N_15864,N_15710,N_15532);
or U15865 (N_15865,N_15646,N_15571);
xor U15866 (N_15866,N_15665,N_15520);
or U15867 (N_15867,N_15518,N_15709);
xor U15868 (N_15868,N_15584,N_15700);
nand U15869 (N_15869,N_15525,N_15594);
nand U15870 (N_15870,N_15590,N_15702);
nand U15871 (N_15871,N_15592,N_15615);
nor U15872 (N_15872,N_15618,N_15547);
and U15873 (N_15873,N_15548,N_15637);
nor U15874 (N_15874,N_15549,N_15696);
nand U15875 (N_15875,N_15513,N_15612);
and U15876 (N_15876,N_15709,N_15680);
nor U15877 (N_15877,N_15603,N_15685);
and U15878 (N_15878,N_15609,N_15711);
or U15879 (N_15879,N_15737,N_15548);
nor U15880 (N_15880,N_15705,N_15548);
and U15881 (N_15881,N_15677,N_15719);
or U15882 (N_15882,N_15500,N_15563);
nor U15883 (N_15883,N_15602,N_15632);
xnor U15884 (N_15884,N_15702,N_15556);
and U15885 (N_15885,N_15667,N_15662);
or U15886 (N_15886,N_15566,N_15578);
or U15887 (N_15887,N_15702,N_15596);
xor U15888 (N_15888,N_15646,N_15736);
nand U15889 (N_15889,N_15589,N_15545);
and U15890 (N_15890,N_15524,N_15579);
nor U15891 (N_15891,N_15664,N_15549);
or U15892 (N_15892,N_15718,N_15565);
and U15893 (N_15893,N_15654,N_15713);
nor U15894 (N_15894,N_15726,N_15608);
or U15895 (N_15895,N_15709,N_15693);
nand U15896 (N_15896,N_15528,N_15562);
or U15897 (N_15897,N_15564,N_15655);
and U15898 (N_15898,N_15674,N_15745);
and U15899 (N_15899,N_15689,N_15548);
or U15900 (N_15900,N_15649,N_15739);
or U15901 (N_15901,N_15587,N_15680);
nand U15902 (N_15902,N_15568,N_15714);
nor U15903 (N_15903,N_15619,N_15632);
xnor U15904 (N_15904,N_15667,N_15698);
nor U15905 (N_15905,N_15713,N_15625);
nand U15906 (N_15906,N_15672,N_15558);
nor U15907 (N_15907,N_15569,N_15518);
nand U15908 (N_15908,N_15599,N_15683);
nand U15909 (N_15909,N_15593,N_15559);
xnor U15910 (N_15910,N_15584,N_15711);
and U15911 (N_15911,N_15667,N_15577);
nand U15912 (N_15912,N_15650,N_15675);
and U15913 (N_15913,N_15634,N_15670);
and U15914 (N_15914,N_15573,N_15677);
nor U15915 (N_15915,N_15543,N_15514);
xnor U15916 (N_15916,N_15604,N_15726);
nand U15917 (N_15917,N_15580,N_15522);
nor U15918 (N_15918,N_15720,N_15538);
or U15919 (N_15919,N_15590,N_15739);
and U15920 (N_15920,N_15697,N_15673);
nand U15921 (N_15921,N_15577,N_15583);
or U15922 (N_15922,N_15577,N_15644);
xor U15923 (N_15923,N_15702,N_15699);
and U15924 (N_15924,N_15575,N_15615);
nand U15925 (N_15925,N_15530,N_15625);
nand U15926 (N_15926,N_15636,N_15730);
xor U15927 (N_15927,N_15676,N_15599);
or U15928 (N_15928,N_15540,N_15575);
and U15929 (N_15929,N_15613,N_15541);
xor U15930 (N_15930,N_15516,N_15654);
nand U15931 (N_15931,N_15711,N_15529);
and U15932 (N_15932,N_15613,N_15691);
xnor U15933 (N_15933,N_15664,N_15530);
nand U15934 (N_15934,N_15715,N_15738);
or U15935 (N_15935,N_15701,N_15609);
or U15936 (N_15936,N_15593,N_15574);
and U15937 (N_15937,N_15588,N_15551);
or U15938 (N_15938,N_15701,N_15724);
and U15939 (N_15939,N_15568,N_15609);
nand U15940 (N_15940,N_15563,N_15572);
xor U15941 (N_15941,N_15626,N_15501);
nand U15942 (N_15942,N_15534,N_15581);
and U15943 (N_15943,N_15569,N_15651);
and U15944 (N_15944,N_15567,N_15528);
xor U15945 (N_15945,N_15574,N_15520);
nor U15946 (N_15946,N_15669,N_15682);
or U15947 (N_15947,N_15501,N_15570);
xnor U15948 (N_15948,N_15718,N_15702);
xnor U15949 (N_15949,N_15682,N_15534);
nand U15950 (N_15950,N_15573,N_15633);
nand U15951 (N_15951,N_15649,N_15748);
and U15952 (N_15952,N_15613,N_15589);
nor U15953 (N_15953,N_15533,N_15612);
xnor U15954 (N_15954,N_15643,N_15503);
nor U15955 (N_15955,N_15526,N_15641);
nor U15956 (N_15956,N_15642,N_15746);
xor U15957 (N_15957,N_15639,N_15567);
xnor U15958 (N_15958,N_15645,N_15567);
nor U15959 (N_15959,N_15698,N_15547);
nor U15960 (N_15960,N_15663,N_15658);
or U15961 (N_15961,N_15676,N_15716);
or U15962 (N_15962,N_15723,N_15631);
and U15963 (N_15963,N_15577,N_15616);
and U15964 (N_15964,N_15683,N_15612);
nand U15965 (N_15965,N_15723,N_15714);
nor U15966 (N_15966,N_15717,N_15694);
or U15967 (N_15967,N_15565,N_15690);
nand U15968 (N_15968,N_15736,N_15557);
nor U15969 (N_15969,N_15691,N_15545);
nand U15970 (N_15970,N_15523,N_15576);
or U15971 (N_15971,N_15665,N_15648);
xor U15972 (N_15972,N_15612,N_15599);
and U15973 (N_15973,N_15609,N_15631);
and U15974 (N_15974,N_15508,N_15545);
nand U15975 (N_15975,N_15701,N_15630);
xor U15976 (N_15976,N_15747,N_15602);
and U15977 (N_15977,N_15610,N_15510);
nor U15978 (N_15978,N_15594,N_15640);
or U15979 (N_15979,N_15614,N_15507);
xnor U15980 (N_15980,N_15537,N_15589);
xor U15981 (N_15981,N_15746,N_15712);
or U15982 (N_15982,N_15615,N_15611);
nor U15983 (N_15983,N_15536,N_15615);
nand U15984 (N_15984,N_15705,N_15517);
or U15985 (N_15985,N_15663,N_15566);
xor U15986 (N_15986,N_15679,N_15578);
and U15987 (N_15987,N_15578,N_15552);
or U15988 (N_15988,N_15720,N_15713);
xnor U15989 (N_15989,N_15642,N_15644);
and U15990 (N_15990,N_15636,N_15566);
and U15991 (N_15991,N_15603,N_15588);
or U15992 (N_15992,N_15647,N_15713);
xor U15993 (N_15993,N_15745,N_15658);
nor U15994 (N_15994,N_15588,N_15654);
or U15995 (N_15995,N_15731,N_15587);
nand U15996 (N_15996,N_15734,N_15748);
and U15997 (N_15997,N_15679,N_15643);
and U15998 (N_15998,N_15638,N_15716);
nand U15999 (N_15999,N_15565,N_15726);
nor U16000 (N_16000,N_15867,N_15786);
or U16001 (N_16001,N_15908,N_15764);
and U16002 (N_16002,N_15998,N_15788);
nand U16003 (N_16003,N_15811,N_15758);
nand U16004 (N_16004,N_15876,N_15969);
xnor U16005 (N_16005,N_15902,N_15870);
xor U16006 (N_16006,N_15755,N_15946);
xnor U16007 (N_16007,N_15795,N_15851);
or U16008 (N_16008,N_15874,N_15956);
xnor U16009 (N_16009,N_15925,N_15915);
and U16010 (N_16010,N_15873,N_15960);
nand U16011 (N_16011,N_15994,N_15937);
nand U16012 (N_16012,N_15978,N_15975);
xnor U16013 (N_16013,N_15772,N_15865);
xnor U16014 (N_16014,N_15776,N_15914);
xor U16015 (N_16015,N_15927,N_15922);
xor U16016 (N_16016,N_15973,N_15942);
or U16017 (N_16017,N_15910,N_15947);
or U16018 (N_16018,N_15905,N_15808);
nand U16019 (N_16019,N_15948,N_15923);
nor U16020 (N_16020,N_15751,N_15752);
nor U16021 (N_16021,N_15968,N_15831);
or U16022 (N_16022,N_15896,N_15880);
xnor U16023 (N_16023,N_15853,N_15839);
nand U16024 (N_16024,N_15785,N_15816);
nand U16025 (N_16025,N_15797,N_15988);
nor U16026 (N_16026,N_15818,N_15835);
nand U16027 (N_16027,N_15939,N_15763);
and U16028 (N_16028,N_15997,N_15836);
xor U16029 (N_16029,N_15966,N_15829);
or U16030 (N_16030,N_15809,N_15825);
and U16031 (N_16031,N_15753,N_15787);
xor U16032 (N_16032,N_15928,N_15857);
nor U16033 (N_16033,N_15961,N_15990);
and U16034 (N_16034,N_15893,N_15985);
or U16035 (N_16035,N_15805,N_15815);
and U16036 (N_16036,N_15850,N_15982);
nand U16037 (N_16037,N_15898,N_15983);
nor U16038 (N_16038,N_15989,N_15761);
nor U16039 (N_16039,N_15800,N_15897);
xnor U16040 (N_16040,N_15931,N_15771);
and U16041 (N_16041,N_15812,N_15762);
and U16042 (N_16042,N_15862,N_15930);
and U16043 (N_16043,N_15855,N_15885);
and U16044 (N_16044,N_15819,N_15806);
nor U16045 (N_16045,N_15760,N_15912);
xnor U16046 (N_16046,N_15813,N_15833);
xor U16047 (N_16047,N_15777,N_15859);
xor U16048 (N_16048,N_15909,N_15860);
and U16049 (N_16049,N_15953,N_15974);
and U16050 (N_16050,N_15796,N_15767);
or U16051 (N_16051,N_15972,N_15954);
xor U16052 (N_16052,N_15878,N_15828);
nand U16053 (N_16053,N_15826,N_15849);
and U16054 (N_16054,N_15863,N_15790);
nor U16055 (N_16055,N_15801,N_15951);
xor U16056 (N_16056,N_15827,N_15992);
nor U16057 (N_16057,N_15881,N_15793);
or U16058 (N_16058,N_15964,N_15963);
xnor U16059 (N_16059,N_15929,N_15916);
nand U16060 (N_16060,N_15892,N_15765);
or U16061 (N_16061,N_15759,N_15775);
and U16062 (N_16062,N_15841,N_15903);
or U16063 (N_16063,N_15814,N_15875);
or U16064 (N_16064,N_15976,N_15784);
or U16065 (N_16065,N_15770,N_15934);
xnor U16066 (N_16066,N_15944,N_15821);
or U16067 (N_16067,N_15952,N_15757);
xnor U16068 (N_16068,N_15958,N_15803);
nor U16069 (N_16069,N_15766,N_15991);
nand U16070 (N_16070,N_15807,N_15884);
or U16071 (N_16071,N_15769,N_15750);
nor U16072 (N_16072,N_15773,N_15913);
and U16073 (N_16073,N_15887,N_15844);
nand U16074 (N_16074,N_15965,N_15941);
and U16075 (N_16075,N_15779,N_15993);
nand U16076 (N_16076,N_15890,N_15798);
nand U16077 (N_16077,N_15856,N_15879);
or U16078 (N_16078,N_15971,N_15926);
nand U16079 (N_16079,N_15906,N_15888);
nand U16080 (N_16080,N_15987,N_15780);
or U16081 (N_16081,N_15962,N_15783);
or U16082 (N_16082,N_15904,N_15891);
nor U16083 (N_16083,N_15936,N_15768);
xnor U16084 (N_16084,N_15935,N_15921);
nand U16085 (N_16085,N_15918,N_15846);
nor U16086 (N_16086,N_15981,N_15756);
nor U16087 (N_16087,N_15945,N_15864);
or U16088 (N_16088,N_15834,N_15843);
nor U16089 (N_16089,N_15996,N_15858);
nand U16090 (N_16090,N_15920,N_15822);
nor U16091 (N_16091,N_15868,N_15802);
and U16092 (N_16092,N_15817,N_15791);
and U16093 (N_16093,N_15866,N_15877);
or U16094 (N_16094,N_15933,N_15882);
or U16095 (N_16095,N_15792,N_15949);
xor U16096 (N_16096,N_15781,N_15782);
nor U16097 (N_16097,N_15901,N_15900);
nand U16098 (N_16098,N_15979,N_15957);
xnor U16099 (N_16099,N_15799,N_15840);
or U16100 (N_16100,N_15919,N_15977);
or U16101 (N_16101,N_15889,N_15911);
or U16102 (N_16102,N_15861,N_15838);
or U16103 (N_16103,N_15943,N_15830);
nor U16104 (N_16104,N_15847,N_15886);
nor U16105 (N_16105,N_15832,N_15940);
and U16106 (N_16106,N_15824,N_15894);
xor U16107 (N_16107,N_15842,N_15899);
and U16108 (N_16108,N_15895,N_15774);
nor U16109 (N_16109,N_15820,N_15810);
nor U16110 (N_16110,N_15959,N_15883);
or U16111 (N_16111,N_15955,N_15984);
and U16112 (N_16112,N_15872,N_15907);
or U16113 (N_16113,N_15871,N_15938);
xor U16114 (N_16114,N_15778,N_15794);
and U16115 (N_16115,N_15999,N_15932);
nor U16116 (N_16116,N_15837,N_15950);
nor U16117 (N_16117,N_15848,N_15986);
nand U16118 (N_16118,N_15995,N_15917);
or U16119 (N_16119,N_15845,N_15869);
or U16120 (N_16120,N_15980,N_15823);
nor U16121 (N_16121,N_15754,N_15789);
or U16122 (N_16122,N_15854,N_15924);
or U16123 (N_16123,N_15970,N_15852);
and U16124 (N_16124,N_15804,N_15967);
or U16125 (N_16125,N_15871,N_15844);
or U16126 (N_16126,N_15798,N_15813);
xnor U16127 (N_16127,N_15924,N_15810);
nor U16128 (N_16128,N_15752,N_15982);
xor U16129 (N_16129,N_15809,N_15993);
nand U16130 (N_16130,N_15876,N_15976);
nor U16131 (N_16131,N_15930,N_15880);
and U16132 (N_16132,N_15952,N_15985);
xor U16133 (N_16133,N_15952,N_15927);
nor U16134 (N_16134,N_15943,N_15760);
nand U16135 (N_16135,N_15938,N_15972);
nor U16136 (N_16136,N_15801,N_15852);
or U16137 (N_16137,N_15916,N_15825);
nor U16138 (N_16138,N_15954,N_15860);
nor U16139 (N_16139,N_15921,N_15978);
xor U16140 (N_16140,N_15789,N_15854);
and U16141 (N_16141,N_15969,N_15792);
and U16142 (N_16142,N_15950,N_15889);
nor U16143 (N_16143,N_15883,N_15801);
or U16144 (N_16144,N_15806,N_15947);
nor U16145 (N_16145,N_15948,N_15865);
xnor U16146 (N_16146,N_15831,N_15959);
nand U16147 (N_16147,N_15959,N_15834);
nand U16148 (N_16148,N_15755,N_15839);
or U16149 (N_16149,N_15916,N_15812);
and U16150 (N_16150,N_15820,N_15915);
nor U16151 (N_16151,N_15928,N_15803);
and U16152 (N_16152,N_15910,N_15878);
nor U16153 (N_16153,N_15998,N_15913);
xnor U16154 (N_16154,N_15823,N_15988);
and U16155 (N_16155,N_15938,N_15975);
nor U16156 (N_16156,N_15789,N_15892);
nand U16157 (N_16157,N_15764,N_15911);
and U16158 (N_16158,N_15948,N_15830);
and U16159 (N_16159,N_15792,N_15892);
xnor U16160 (N_16160,N_15923,N_15841);
xor U16161 (N_16161,N_15992,N_15794);
nand U16162 (N_16162,N_15764,N_15831);
nand U16163 (N_16163,N_15782,N_15951);
nor U16164 (N_16164,N_15899,N_15890);
and U16165 (N_16165,N_15782,N_15950);
nor U16166 (N_16166,N_15880,N_15910);
nand U16167 (N_16167,N_15851,N_15867);
nand U16168 (N_16168,N_15964,N_15822);
xor U16169 (N_16169,N_15998,N_15824);
xnor U16170 (N_16170,N_15955,N_15938);
xor U16171 (N_16171,N_15999,N_15935);
nor U16172 (N_16172,N_15946,N_15958);
nor U16173 (N_16173,N_15884,N_15976);
nor U16174 (N_16174,N_15794,N_15762);
or U16175 (N_16175,N_15927,N_15827);
nand U16176 (N_16176,N_15894,N_15810);
xor U16177 (N_16177,N_15816,N_15981);
xor U16178 (N_16178,N_15943,N_15884);
nand U16179 (N_16179,N_15776,N_15761);
and U16180 (N_16180,N_15750,N_15927);
xor U16181 (N_16181,N_15809,N_15937);
nor U16182 (N_16182,N_15954,N_15776);
nand U16183 (N_16183,N_15955,N_15754);
nor U16184 (N_16184,N_15788,N_15957);
and U16185 (N_16185,N_15851,N_15818);
and U16186 (N_16186,N_15997,N_15938);
xor U16187 (N_16187,N_15928,N_15900);
and U16188 (N_16188,N_15855,N_15867);
xor U16189 (N_16189,N_15892,N_15884);
or U16190 (N_16190,N_15920,N_15883);
nand U16191 (N_16191,N_15902,N_15768);
and U16192 (N_16192,N_15765,N_15913);
or U16193 (N_16193,N_15856,N_15921);
xor U16194 (N_16194,N_15752,N_15811);
nor U16195 (N_16195,N_15801,N_15832);
xor U16196 (N_16196,N_15986,N_15923);
nor U16197 (N_16197,N_15833,N_15761);
xor U16198 (N_16198,N_15839,N_15837);
xor U16199 (N_16199,N_15906,N_15772);
xnor U16200 (N_16200,N_15936,N_15954);
nor U16201 (N_16201,N_15772,N_15929);
nand U16202 (N_16202,N_15927,N_15888);
or U16203 (N_16203,N_15763,N_15767);
nor U16204 (N_16204,N_15893,N_15972);
xor U16205 (N_16205,N_15842,N_15988);
and U16206 (N_16206,N_15826,N_15824);
nand U16207 (N_16207,N_15864,N_15906);
xor U16208 (N_16208,N_15803,N_15809);
or U16209 (N_16209,N_15764,N_15819);
nor U16210 (N_16210,N_15988,N_15907);
nand U16211 (N_16211,N_15874,N_15959);
nor U16212 (N_16212,N_15941,N_15873);
and U16213 (N_16213,N_15870,N_15844);
and U16214 (N_16214,N_15937,N_15812);
nor U16215 (N_16215,N_15756,N_15886);
and U16216 (N_16216,N_15818,N_15958);
nand U16217 (N_16217,N_15957,N_15915);
and U16218 (N_16218,N_15948,N_15810);
xor U16219 (N_16219,N_15838,N_15943);
xor U16220 (N_16220,N_15869,N_15878);
and U16221 (N_16221,N_15879,N_15898);
or U16222 (N_16222,N_15976,N_15929);
or U16223 (N_16223,N_15947,N_15949);
and U16224 (N_16224,N_15949,N_15764);
and U16225 (N_16225,N_15915,N_15980);
and U16226 (N_16226,N_15791,N_15753);
xnor U16227 (N_16227,N_15983,N_15821);
nor U16228 (N_16228,N_15886,N_15852);
nand U16229 (N_16229,N_15913,N_15965);
xnor U16230 (N_16230,N_15932,N_15822);
nor U16231 (N_16231,N_15978,N_15972);
nor U16232 (N_16232,N_15864,N_15815);
xnor U16233 (N_16233,N_15995,N_15859);
or U16234 (N_16234,N_15882,N_15824);
xor U16235 (N_16235,N_15933,N_15818);
xnor U16236 (N_16236,N_15845,N_15915);
nor U16237 (N_16237,N_15856,N_15905);
and U16238 (N_16238,N_15797,N_15804);
and U16239 (N_16239,N_15990,N_15790);
nor U16240 (N_16240,N_15987,N_15916);
nor U16241 (N_16241,N_15948,N_15771);
xor U16242 (N_16242,N_15905,N_15864);
xor U16243 (N_16243,N_15797,N_15864);
nor U16244 (N_16244,N_15909,N_15917);
xnor U16245 (N_16245,N_15930,N_15914);
and U16246 (N_16246,N_15863,N_15906);
nand U16247 (N_16247,N_15999,N_15800);
nor U16248 (N_16248,N_15781,N_15925);
or U16249 (N_16249,N_15792,N_15831);
nor U16250 (N_16250,N_16085,N_16024);
nand U16251 (N_16251,N_16097,N_16094);
or U16252 (N_16252,N_16234,N_16147);
or U16253 (N_16253,N_16110,N_16125);
or U16254 (N_16254,N_16003,N_16068);
and U16255 (N_16255,N_16166,N_16145);
nor U16256 (N_16256,N_16242,N_16170);
nand U16257 (N_16257,N_16129,N_16067);
xor U16258 (N_16258,N_16058,N_16049);
nor U16259 (N_16259,N_16059,N_16137);
and U16260 (N_16260,N_16022,N_16134);
xnor U16261 (N_16261,N_16161,N_16036);
nand U16262 (N_16262,N_16245,N_16168);
nand U16263 (N_16263,N_16207,N_16159);
or U16264 (N_16264,N_16146,N_16064);
nand U16265 (N_16265,N_16009,N_16186);
xor U16266 (N_16266,N_16238,N_16192);
xor U16267 (N_16267,N_16176,N_16201);
nand U16268 (N_16268,N_16047,N_16039);
and U16269 (N_16269,N_16179,N_16101);
or U16270 (N_16270,N_16174,N_16127);
and U16271 (N_16271,N_16209,N_16220);
nand U16272 (N_16272,N_16196,N_16045);
and U16273 (N_16273,N_16093,N_16126);
or U16274 (N_16274,N_16099,N_16212);
nand U16275 (N_16275,N_16183,N_16041);
and U16276 (N_16276,N_16107,N_16138);
nor U16277 (N_16277,N_16164,N_16066);
nand U16278 (N_16278,N_16032,N_16157);
nand U16279 (N_16279,N_16084,N_16105);
nor U16280 (N_16280,N_16154,N_16246);
nor U16281 (N_16281,N_16232,N_16029);
xor U16282 (N_16282,N_16240,N_16076);
nor U16283 (N_16283,N_16208,N_16187);
nor U16284 (N_16284,N_16016,N_16158);
nor U16285 (N_16285,N_16004,N_16162);
xnor U16286 (N_16286,N_16079,N_16102);
xor U16287 (N_16287,N_16199,N_16062);
xor U16288 (N_16288,N_16113,N_16108);
and U16289 (N_16289,N_16198,N_16033);
nand U16290 (N_16290,N_16046,N_16218);
nor U16291 (N_16291,N_16028,N_16120);
nor U16292 (N_16292,N_16075,N_16103);
nand U16293 (N_16293,N_16098,N_16155);
nor U16294 (N_16294,N_16061,N_16226);
xor U16295 (N_16295,N_16136,N_16019);
and U16296 (N_16296,N_16082,N_16141);
or U16297 (N_16297,N_16030,N_16178);
nor U16298 (N_16298,N_16215,N_16050);
xnor U16299 (N_16299,N_16228,N_16048);
or U16300 (N_16300,N_16160,N_16006);
nand U16301 (N_16301,N_16195,N_16181);
or U16302 (N_16302,N_16005,N_16132);
and U16303 (N_16303,N_16221,N_16071);
or U16304 (N_16304,N_16051,N_16247);
or U16305 (N_16305,N_16153,N_16193);
or U16306 (N_16306,N_16149,N_16189);
or U16307 (N_16307,N_16185,N_16092);
xnor U16308 (N_16308,N_16026,N_16000);
or U16309 (N_16309,N_16167,N_16057);
or U16310 (N_16310,N_16236,N_16008);
or U16311 (N_16311,N_16089,N_16063);
xor U16312 (N_16312,N_16015,N_16197);
nand U16313 (N_16313,N_16217,N_16073);
or U16314 (N_16314,N_16111,N_16190);
nand U16315 (N_16315,N_16114,N_16130);
nor U16316 (N_16316,N_16038,N_16202);
and U16317 (N_16317,N_16031,N_16229);
or U16318 (N_16318,N_16227,N_16011);
xnor U16319 (N_16319,N_16241,N_16204);
nor U16320 (N_16320,N_16018,N_16025);
and U16321 (N_16321,N_16072,N_16117);
nand U16322 (N_16322,N_16078,N_16135);
xnor U16323 (N_16323,N_16007,N_16148);
xor U16324 (N_16324,N_16224,N_16222);
xor U16325 (N_16325,N_16194,N_16177);
or U16326 (N_16326,N_16054,N_16121);
nor U16327 (N_16327,N_16017,N_16090);
nor U16328 (N_16328,N_16010,N_16172);
nand U16329 (N_16329,N_16230,N_16128);
nand U16330 (N_16330,N_16211,N_16052);
nand U16331 (N_16331,N_16069,N_16091);
xor U16332 (N_16332,N_16248,N_16070);
or U16333 (N_16333,N_16225,N_16144);
and U16334 (N_16334,N_16180,N_16165);
or U16335 (N_16335,N_16118,N_16055);
nand U16336 (N_16336,N_16083,N_16001);
xnor U16337 (N_16337,N_16216,N_16231);
nand U16338 (N_16338,N_16034,N_16020);
and U16339 (N_16339,N_16239,N_16140);
xnor U16340 (N_16340,N_16081,N_16219);
nand U16341 (N_16341,N_16205,N_16088);
xnor U16342 (N_16342,N_16214,N_16115);
xnor U16343 (N_16343,N_16012,N_16056);
or U16344 (N_16344,N_16123,N_16095);
nand U16345 (N_16345,N_16171,N_16060);
xnor U16346 (N_16346,N_16233,N_16087);
or U16347 (N_16347,N_16044,N_16013);
nor U16348 (N_16348,N_16151,N_16156);
xor U16349 (N_16349,N_16191,N_16188);
nand U16350 (N_16350,N_16037,N_16109);
nor U16351 (N_16351,N_16139,N_16169);
nor U16352 (N_16352,N_16210,N_16243);
xor U16353 (N_16353,N_16142,N_16106);
nor U16354 (N_16354,N_16235,N_16116);
or U16355 (N_16355,N_16143,N_16131);
or U16356 (N_16356,N_16065,N_16023);
nand U16357 (N_16357,N_16042,N_16112);
and U16358 (N_16358,N_16133,N_16249);
and U16359 (N_16359,N_16021,N_16182);
nand U16360 (N_16360,N_16027,N_16223);
xnor U16361 (N_16361,N_16213,N_16100);
or U16362 (N_16362,N_16206,N_16096);
nand U16363 (N_16363,N_16203,N_16040);
or U16364 (N_16364,N_16150,N_16014);
nor U16365 (N_16365,N_16053,N_16244);
xnor U16366 (N_16366,N_16163,N_16086);
nor U16367 (N_16367,N_16152,N_16035);
or U16368 (N_16368,N_16104,N_16122);
xnor U16369 (N_16369,N_16043,N_16173);
or U16370 (N_16370,N_16119,N_16002);
or U16371 (N_16371,N_16175,N_16237);
xnor U16372 (N_16372,N_16184,N_16074);
or U16373 (N_16373,N_16077,N_16080);
nor U16374 (N_16374,N_16200,N_16124);
or U16375 (N_16375,N_16239,N_16011);
xnor U16376 (N_16376,N_16243,N_16015);
or U16377 (N_16377,N_16019,N_16153);
xor U16378 (N_16378,N_16150,N_16000);
nor U16379 (N_16379,N_16231,N_16090);
or U16380 (N_16380,N_16017,N_16151);
and U16381 (N_16381,N_16146,N_16126);
nor U16382 (N_16382,N_16184,N_16031);
and U16383 (N_16383,N_16056,N_16057);
nand U16384 (N_16384,N_16158,N_16233);
xor U16385 (N_16385,N_16171,N_16045);
nand U16386 (N_16386,N_16201,N_16033);
nor U16387 (N_16387,N_16241,N_16005);
nor U16388 (N_16388,N_16182,N_16128);
nor U16389 (N_16389,N_16226,N_16174);
nor U16390 (N_16390,N_16057,N_16045);
and U16391 (N_16391,N_16121,N_16115);
nor U16392 (N_16392,N_16051,N_16014);
xor U16393 (N_16393,N_16124,N_16216);
nand U16394 (N_16394,N_16187,N_16171);
nor U16395 (N_16395,N_16246,N_16182);
xor U16396 (N_16396,N_16165,N_16245);
nor U16397 (N_16397,N_16219,N_16141);
and U16398 (N_16398,N_16046,N_16181);
xnor U16399 (N_16399,N_16114,N_16208);
nand U16400 (N_16400,N_16112,N_16191);
xnor U16401 (N_16401,N_16101,N_16037);
nand U16402 (N_16402,N_16056,N_16050);
or U16403 (N_16403,N_16198,N_16154);
and U16404 (N_16404,N_16056,N_16156);
xnor U16405 (N_16405,N_16081,N_16106);
nand U16406 (N_16406,N_16001,N_16239);
xnor U16407 (N_16407,N_16101,N_16084);
nand U16408 (N_16408,N_16054,N_16206);
xnor U16409 (N_16409,N_16078,N_16150);
and U16410 (N_16410,N_16232,N_16037);
nor U16411 (N_16411,N_16117,N_16004);
xnor U16412 (N_16412,N_16057,N_16113);
or U16413 (N_16413,N_16094,N_16152);
nor U16414 (N_16414,N_16149,N_16043);
xnor U16415 (N_16415,N_16081,N_16121);
and U16416 (N_16416,N_16218,N_16155);
xnor U16417 (N_16417,N_16133,N_16226);
xnor U16418 (N_16418,N_16197,N_16140);
nand U16419 (N_16419,N_16183,N_16075);
nand U16420 (N_16420,N_16054,N_16136);
and U16421 (N_16421,N_16130,N_16160);
or U16422 (N_16422,N_16159,N_16071);
nand U16423 (N_16423,N_16102,N_16037);
nor U16424 (N_16424,N_16140,N_16055);
and U16425 (N_16425,N_16051,N_16024);
and U16426 (N_16426,N_16057,N_16235);
and U16427 (N_16427,N_16084,N_16125);
xnor U16428 (N_16428,N_16098,N_16047);
and U16429 (N_16429,N_16127,N_16214);
nor U16430 (N_16430,N_16152,N_16044);
and U16431 (N_16431,N_16082,N_16190);
and U16432 (N_16432,N_16069,N_16181);
and U16433 (N_16433,N_16198,N_16105);
nor U16434 (N_16434,N_16224,N_16237);
xor U16435 (N_16435,N_16033,N_16108);
nor U16436 (N_16436,N_16155,N_16126);
nor U16437 (N_16437,N_16201,N_16152);
or U16438 (N_16438,N_16003,N_16130);
and U16439 (N_16439,N_16071,N_16009);
nor U16440 (N_16440,N_16142,N_16025);
nand U16441 (N_16441,N_16122,N_16016);
nand U16442 (N_16442,N_16218,N_16160);
and U16443 (N_16443,N_16128,N_16086);
or U16444 (N_16444,N_16184,N_16102);
nand U16445 (N_16445,N_16180,N_16085);
and U16446 (N_16446,N_16207,N_16033);
nand U16447 (N_16447,N_16165,N_16064);
and U16448 (N_16448,N_16134,N_16011);
or U16449 (N_16449,N_16108,N_16125);
nor U16450 (N_16450,N_16023,N_16117);
and U16451 (N_16451,N_16200,N_16133);
nor U16452 (N_16452,N_16235,N_16219);
nand U16453 (N_16453,N_16173,N_16039);
and U16454 (N_16454,N_16082,N_16203);
nand U16455 (N_16455,N_16048,N_16018);
and U16456 (N_16456,N_16249,N_16015);
nand U16457 (N_16457,N_16200,N_16118);
xor U16458 (N_16458,N_16003,N_16238);
nor U16459 (N_16459,N_16073,N_16004);
and U16460 (N_16460,N_16245,N_16230);
or U16461 (N_16461,N_16241,N_16206);
nand U16462 (N_16462,N_16240,N_16222);
nor U16463 (N_16463,N_16206,N_16168);
nand U16464 (N_16464,N_16151,N_16219);
nand U16465 (N_16465,N_16225,N_16132);
xor U16466 (N_16466,N_16221,N_16040);
nand U16467 (N_16467,N_16170,N_16000);
or U16468 (N_16468,N_16107,N_16050);
or U16469 (N_16469,N_16047,N_16108);
and U16470 (N_16470,N_16030,N_16200);
xor U16471 (N_16471,N_16220,N_16045);
xor U16472 (N_16472,N_16211,N_16042);
or U16473 (N_16473,N_16193,N_16165);
and U16474 (N_16474,N_16225,N_16055);
and U16475 (N_16475,N_16008,N_16239);
and U16476 (N_16476,N_16221,N_16014);
nand U16477 (N_16477,N_16177,N_16020);
or U16478 (N_16478,N_16217,N_16136);
nand U16479 (N_16479,N_16147,N_16126);
and U16480 (N_16480,N_16095,N_16043);
xor U16481 (N_16481,N_16208,N_16161);
or U16482 (N_16482,N_16117,N_16021);
nand U16483 (N_16483,N_16009,N_16002);
nor U16484 (N_16484,N_16238,N_16135);
and U16485 (N_16485,N_16003,N_16011);
nor U16486 (N_16486,N_16199,N_16028);
xnor U16487 (N_16487,N_16218,N_16195);
nand U16488 (N_16488,N_16112,N_16031);
xor U16489 (N_16489,N_16128,N_16027);
nand U16490 (N_16490,N_16008,N_16101);
or U16491 (N_16491,N_16151,N_16119);
nor U16492 (N_16492,N_16193,N_16065);
and U16493 (N_16493,N_16021,N_16127);
nor U16494 (N_16494,N_16245,N_16170);
or U16495 (N_16495,N_16096,N_16177);
xor U16496 (N_16496,N_16189,N_16196);
xor U16497 (N_16497,N_16138,N_16017);
nand U16498 (N_16498,N_16167,N_16195);
and U16499 (N_16499,N_16242,N_16204);
xnor U16500 (N_16500,N_16315,N_16261);
nor U16501 (N_16501,N_16258,N_16477);
or U16502 (N_16502,N_16305,N_16356);
nor U16503 (N_16503,N_16293,N_16408);
xnor U16504 (N_16504,N_16371,N_16396);
and U16505 (N_16505,N_16351,N_16262);
xor U16506 (N_16506,N_16463,N_16487);
nor U16507 (N_16507,N_16479,N_16275);
nor U16508 (N_16508,N_16343,N_16439);
and U16509 (N_16509,N_16341,N_16354);
or U16510 (N_16510,N_16394,N_16296);
nand U16511 (N_16511,N_16347,N_16286);
xnor U16512 (N_16512,N_16272,N_16480);
nand U16513 (N_16513,N_16431,N_16337);
xor U16514 (N_16514,N_16367,N_16352);
nand U16515 (N_16515,N_16294,N_16457);
xor U16516 (N_16516,N_16357,N_16453);
nor U16517 (N_16517,N_16498,N_16342);
nand U16518 (N_16518,N_16464,N_16395);
and U16519 (N_16519,N_16376,N_16372);
nor U16520 (N_16520,N_16397,N_16414);
nor U16521 (N_16521,N_16329,N_16319);
xor U16522 (N_16522,N_16255,N_16361);
nor U16523 (N_16523,N_16322,N_16456);
nand U16524 (N_16524,N_16443,N_16270);
nor U16525 (N_16525,N_16393,N_16471);
xnor U16526 (N_16526,N_16484,N_16403);
nand U16527 (N_16527,N_16491,N_16475);
nor U16528 (N_16528,N_16425,N_16325);
nor U16529 (N_16529,N_16266,N_16476);
or U16530 (N_16530,N_16256,N_16497);
or U16531 (N_16531,N_16263,N_16360);
nand U16532 (N_16532,N_16432,N_16338);
and U16533 (N_16533,N_16427,N_16413);
nor U16534 (N_16534,N_16353,N_16318);
and U16535 (N_16535,N_16312,N_16459);
or U16536 (N_16536,N_16494,N_16276);
or U16537 (N_16537,N_16313,N_16374);
nand U16538 (N_16538,N_16451,N_16378);
nor U16539 (N_16539,N_16438,N_16369);
nand U16540 (N_16540,N_16303,N_16277);
nand U16541 (N_16541,N_16301,N_16274);
nand U16542 (N_16542,N_16482,N_16324);
and U16543 (N_16543,N_16271,N_16278);
or U16544 (N_16544,N_16254,N_16445);
nand U16545 (N_16545,N_16426,N_16265);
or U16546 (N_16546,N_16485,N_16469);
xor U16547 (N_16547,N_16365,N_16317);
or U16548 (N_16548,N_16268,N_16448);
or U16549 (N_16549,N_16444,N_16467);
or U16550 (N_16550,N_16348,N_16327);
and U16551 (N_16551,N_16380,N_16349);
nand U16552 (N_16552,N_16326,N_16346);
nor U16553 (N_16553,N_16492,N_16461);
nor U16554 (N_16554,N_16340,N_16295);
nand U16555 (N_16555,N_16437,N_16402);
nor U16556 (N_16556,N_16388,N_16412);
nor U16557 (N_16557,N_16385,N_16300);
and U16558 (N_16558,N_16405,N_16304);
xnor U16559 (N_16559,N_16355,N_16429);
xor U16560 (N_16560,N_16273,N_16259);
xnor U16561 (N_16561,N_16423,N_16363);
and U16562 (N_16562,N_16386,N_16302);
and U16563 (N_16563,N_16251,N_16489);
or U16564 (N_16564,N_16400,N_16350);
nor U16565 (N_16565,N_16499,N_16486);
nor U16566 (N_16566,N_16470,N_16260);
nor U16567 (N_16567,N_16428,N_16409);
and U16568 (N_16568,N_16335,N_16297);
and U16569 (N_16569,N_16288,N_16283);
nor U16570 (N_16570,N_16314,N_16379);
or U16571 (N_16571,N_16292,N_16344);
nand U16572 (N_16572,N_16460,N_16424);
nor U16573 (N_16573,N_16339,N_16488);
nand U16574 (N_16574,N_16267,N_16331);
nor U16575 (N_16575,N_16418,N_16377);
or U16576 (N_16576,N_16441,N_16364);
nor U16577 (N_16577,N_16481,N_16359);
nor U16578 (N_16578,N_16253,N_16373);
nand U16579 (N_16579,N_16328,N_16417);
or U16580 (N_16580,N_16398,N_16473);
and U16581 (N_16581,N_16495,N_16490);
nor U16582 (N_16582,N_16466,N_16311);
nor U16583 (N_16583,N_16472,N_16264);
xor U16584 (N_16584,N_16252,N_16307);
xnor U16585 (N_16585,N_16422,N_16269);
or U16586 (N_16586,N_16298,N_16446);
and U16587 (N_16587,N_16383,N_16435);
or U16588 (N_16588,N_16392,N_16452);
xor U16589 (N_16589,N_16391,N_16440);
or U16590 (N_16590,N_16330,N_16496);
or U16591 (N_16591,N_16345,N_16436);
nand U16592 (N_16592,N_16323,N_16291);
xor U16593 (N_16593,N_16309,N_16416);
or U16594 (N_16594,N_16334,N_16281);
xor U16595 (N_16595,N_16310,N_16447);
xor U16596 (N_16596,N_16401,N_16468);
xor U16597 (N_16597,N_16455,N_16454);
and U16598 (N_16598,N_16421,N_16336);
and U16599 (N_16599,N_16399,N_16419);
xnor U16600 (N_16600,N_16287,N_16279);
nor U16601 (N_16601,N_16407,N_16316);
nor U16602 (N_16602,N_16390,N_16358);
xor U16603 (N_16603,N_16384,N_16320);
and U16604 (N_16604,N_16366,N_16411);
xnor U16605 (N_16605,N_16375,N_16389);
nor U16606 (N_16606,N_16465,N_16493);
or U16607 (N_16607,N_16410,N_16257);
or U16608 (N_16608,N_16404,N_16368);
and U16609 (N_16609,N_16306,N_16450);
or U16610 (N_16610,N_16462,N_16290);
or U16611 (N_16611,N_16449,N_16370);
nor U16612 (N_16612,N_16299,N_16381);
nand U16613 (N_16613,N_16387,N_16382);
nand U16614 (N_16614,N_16474,N_16420);
nand U16615 (N_16615,N_16434,N_16282);
nand U16616 (N_16616,N_16362,N_16406);
xnor U16617 (N_16617,N_16280,N_16430);
or U16618 (N_16618,N_16478,N_16284);
nor U16619 (N_16619,N_16332,N_16321);
or U16620 (N_16620,N_16433,N_16289);
nor U16621 (N_16621,N_16333,N_16442);
and U16622 (N_16622,N_16415,N_16483);
xnor U16623 (N_16623,N_16250,N_16458);
and U16624 (N_16624,N_16308,N_16285);
nor U16625 (N_16625,N_16429,N_16321);
or U16626 (N_16626,N_16490,N_16427);
xnor U16627 (N_16627,N_16361,N_16381);
nand U16628 (N_16628,N_16444,N_16293);
nor U16629 (N_16629,N_16370,N_16409);
nand U16630 (N_16630,N_16253,N_16495);
nor U16631 (N_16631,N_16490,N_16432);
nand U16632 (N_16632,N_16343,N_16267);
nand U16633 (N_16633,N_16479,N_16252);
or U16634 (N_16634,N_16331,N_16293);
nand U16635 (N_16635,N_16266,N_16432);
xnor U16636 (N_16636,N_16412,N_16302);
or U16637 (N_16637,N_16293,N_16335);
xor U16638 (N_16638,N_16487,N_16329);
nor U16639 (N_16639,N_16490,N_16491);
and U16640 (N_16640,N_16436,N_16402);
xnor U16641 (N_16641,N_16498,N_16352);
or U16642 (N_16642,N_16324,N_16388);
xor U16643 (N_16643,N_16426,N_16387);
nor U16644 (N_16644,N_16493,N_16347);
and U16645 (N_16645,N_16461,N_16456);
and U16646 (N_16646,N_16478,N_16358);
xor U16647 (N_16647,N_16446,N_16451);
nand U16648 (N_16648,N_16389,N_16442);
xor U16649 (N_16649,N_16342,N_16353);
nor U16650 (N_16650,N_16340,N_16497);
nand U16651 (N_16651,N_16329,N_16356);
xor U16652 (N_16652,N_16386,N_16324);
xor U16653 (N_16653,N_16429,N_16400);
and U16654 (N_16654,N_16294,N_16313);
nor U16655 (N_16655,N_16343,N_16452);
nor U16656 (N_16656,N_16261,N_16328);
nand U16657 (N_16657,N_16451,N_16425);
xnor U16658 (N_16658,N_16251,N_16317);
nand U16659 (N_16659,N_16276,N_16441);
nand U16660 (N_16660,N_16288,N_16324);
xnor U16661 (N_16661,N_16380,N_16333);
or U16662 (N_16662,N_16367,N_16336);
nand U16663 (N_16663,N_16328,N_16345);
nor U16664 (N_16664,N_16345,N_16387);
xnor U16665 (N_16665,N_16265,N_16272);
nor U16666 (N_16666,N_16321,N_16495);
nand U16667 (N_16667,N_16267,N_16475);
and U16668 (N_16668,N_16409,N_16403);
nand U16669 (N_16669,N_16423,N_16473);
or U16670 (N_16670,N_16381,N_16443);
and U16671 (N_16671,N_16437,N_16371);
and U16672 (N_16672,N_16403,N_16366);
xnor U16673 (N_16673,N_16440,N_16374);
or U16674 (N_16674,N_16271,N_16489);
nand U16675 (N_16675,N_16419,N_16461);
or U16676 (N_16676,N_16415,N_16355);
nor U16677 (N_16677,N_16386,N_16299);
nor U16678 (N_16678,N_16416,N_16407);
xor U16679 (N_16679,N_16489,N_16345);
and U16680 (N_16680,N_16275,N_16264);
nor U16681 (N_16681,N_16328,N_16382);
nand U16682 (N_16682,N_16327,N_16344);
xnor U16683 (N_16683,N_16262,N_16308);
nor U16684 (N_16684,N_16477,N_16431);
xor U16685 (N_16685,N_16434,N_16304);
xor U16686 (N_16686,N_16329,N_16407);
and U16687 (N_16687,N_16399,N_16328);
nor U16688 (N_16688,N_16412,N_16378);
nor U16689 (N_16689,N_16372,N_16409);
and U16690 (N_16690,N_16482,N_16369);
or U16691 (N_16691,N_16403,N_16306);
or U16692 (N_16692,N_16280,N_16330);
nand U16693 (N_16693,N_16334,N_16445);
and U16694 (N_16694,N_16421,N_16261);
nand U16695 (N_16695,N_16410,N_16288);
nand U16696 (N_16696,N_16279,N_16435);
nor U16697 (N_16697,N_16291,N_16414);
xor U16698 (N_16698,N_16322,N_16287);
and U16699 (N_16699,N_16339,N_16300);
nand U16700 (N_16700,N_16328,N_16275);
nor U16701 (N_16701,N_16289,N_16321);
xor U16702 (N_16702,N_16413,N_16304);
nand U16703 (N_16703,N_16363,N_16435);
nand U16704 (N_16704,N_16277,N_16354);
xnor U16705 (N_16705,N_16474,N_16494);
nand U16706 (N_16706,N_16285,N_16479);
or U16707 (N_16707,N_16312,N_16375);
and U16708 (N_16708,N_16462,N_16440);
xor U16709 (N_16709,N_16446,N_16395);
and U16710 (N_16710,N_16339,N_16330);
or U16711 (N_16711,N_16339,N_16367);
or U16712 (N_16712,N_16321,N_16360);
nand U16713 (N_16713,N_16346,N_16366);
xor U16714 (N_16714,N_16479,N_16265);
and U16715 (N_16715,N_16438,N_16351);
nor U16716 (N_16716,N_16423,N_16494);
or U16717 (N_16717,N_16346,N_16265);
nand U16718 (N_16718,N_16327,N_16275);
xnor U16719 (N_16719,N_16341,N_16464);
and U16720 (N_16720,N_16251,N_16379);
nand U16721 (N_16721,N_16375,N_16413);
nor U16722 (N_16722,N_16317,N_16285);
and U16723 (N_16723,N_16255,N_16291);
or U16724 (N_16724,N_16315,N_16478);
nor U16725 (N_16725,N_16281,N_16276);
and U16726 (N_16726,N_16430,N_16457);
nor U16727 (N_16727,N_16459,N_16348);
and U16728 (N_16728,N_16416,N_16336);
nand U16729 (N_16729,N_16359,N_16453);
nor U16730 (N_16730,N_16344,N_16311);
or U16731 (N_16731,N_16486,N_16359);
xor U16732 (N_16732,N_16439,N_16360);
xnor U16733 (N_16733,N_16430,N_16254);
nand U16734 (N_16734,N_16354,N_16294);
and U16735 (N_16735,N_16483,N_16344);
and U16736 (N_16736,N_16308,N_16487);
nand U16737 (N_16737,N_16411,N_16278);
xnor U16738 (N_16738,N_16398,N_16341);
or U16739 (N_16739,N_16259,N_16268);
or U16740 (N_16740,N_16397,N_16255);
nor U16741 (N_16741,N_16421,N_16473);
and U16742 (N_16742,N_16259,N_16405);
and U16743 (N_16743,N_16433,N_16254);
nor U16744 (N_16744,N_16442,N_16403);
xnor U16745 (N_16745,N_16406,N_16267);
and U16746 (N_16746,N_16331,N_16261);
xor U16747 (N_16747,N_16468,N_16257);
nor U16748 (N_16748,N_16482,N_16318);
nand U16749 (N_16749,N_16425,N_16370);
xnor U16750 (N_16750,N_16530,N_16728);
or U16751 (N_16751,N_16634,N_16723);
or U16752 (N_16752,N_16520,N_16562);
nand U16753 (N_16753,N_16623,N_16616);
and U16754 (N_16754,N_16666,N_16517);
xnor U16755 (N_16755,N_16708,N_16629);
nor U16756 (N_16756,N_16555,N_16596);
xor U16757 (N_16757,N_16539,N_16516);
nor U16758 (N_16758,N_16542,N_16578);
nor U16759 (N_16759,N_16592,N_16696);
and U16760 (N_16760,N_16710,N_16613);
xnor U16761 (N_16761,N_16604,N_16677);
and U16762 (N_16762,N_16687,N_16577);
or U16763 (N_16763,N_16515,N_16587);
xor U16764 (N_16764,N_16675,N_16683);
nor U16765 (N_16765,N_16698,N_16511);
nand U16766 (N_16766,N_16618,N_16735);
nand U16767 (N_16767,N_16713,N_16615);
and U16768 (N_16768,N_16619,N_16660);
nor U16769 (N_16769,N_16681,N_16695);
or U16770 (N_16770,N_16513,N_16658);
or U16771 (N_16771,N_16664,N_16700);
or U16772 (N_16772,N_16525,N_16657);
nor U16773 (N_16773,N_16649,N_16575);
and U16774 (N_16774,N_16514,N_16565);
and U16775 (N_16775,N_16568,N_16746);
or U16776 (N_16776,N_16699,N_16504);
or U16777 (N_16777,N_16742,N_16557);
nand U16778 (N_16778,N_16741,N_16506);
and U16779 (N_16779,N_16680,N_16545);
xor U16780 (N_16780,N_16556,N_16685);
xor U16781 (N_16781,N_16673,N_16571);
nand U16782 (N_16782,N_16572,N_16548);
xnor U16783 (N_16783,N_16606,N_16653);
and U16784 (N_16784,N_16676,N_16648);
nand U16785 (N_16785,N_16724,N_16534);
nor U16786 (N_16786,N_16737,N_16652);
xor U16787 (N_16787,N_16720,N_16638);
xnor U16788 (N_16788,N_16684,N_16558);
or U16789 (N_16789,N_16704,N_16707);
or U16790 (N_16790,N_16636,N_16512);
nand U16791 (N_16791,N_16725,N_16612);
nor U16792 (N_16792,N_16627,N_16570);
xor U16793 (N_16793,N_16547,N_16559);
or U16794 (N_16794,N_16718,N_16553);
nand U16795 (N_16795,N_16549,N_16546);
xnor U16796 (N_16796,N_16607,N_16654);
xnor U16797 (N_16797,N_16691,N_16682);
xor U16798 (N_16798,N_16632,N_16608);
nand U16799 (N_16799,N_16591,N_16576);
and U16800 (N_16800,N_16583,N_16518);
nand U16801 (N_16801,N_16661,N_16602);
xnor U16802 (N_16802,N_16701,N_16538);
nor U16803 (N_16803,N_16533,N_16573);
nor U16804 (N_16804,N_16609,N_16597);
nor U16805 (N_16805,N_16635,N_16509);
nor U16806 (N_16806,N_16581,N_16738);
nand U16807 (N_16807,N_16605,N_16611);
or U16808 (N_16808,N_16719,N_16665);
nand U16809 (N_16809,N_16594,N_16650);
or U16810 (N_16810,N_16709,N_16643);
nor U16811 (N_16811,N_16736,N_16529);
nor U16812 (N_16812,N_16703,N_16730);
and U16813 (N_16813,N_16712,N_16543);
nand U16814 (N_16814,N_16519,N_16744);
and U16815 (N_16815,N_16552,N_16580);
or U16816 (N_16816,N_16579,N_16726);
and U16817 (N_16817,N_16540,N_16731);
nand U16818 (N_16818,N_16733,N_16510);
nand U16819 (N_16819,N_16689,N_16528);
or U16820 (N_16820,N_16531,N_16532);
nand U16821 (N_16821,N_16690,N_16715);
and U16822 (N_16822,N_16641,N_16745);
nor U16823 (N_16823,N_16706,N_16655);
and U16824 (N_16824,N_16586,N_16625);
and U16825 (N_16825,N_16717,N_16561);
nor U16826 (N_16826,N_16721,N_16523);
nor U16827 (N_16827,N_16659,N_16527);
or U16828 (N_16828,N_16574,N_16590);
nor U16829 (N_16829,N_16662,N_16729);
or U16830 (N_16830,N_16705,N_16656);
xor U16831 (N_16831,N_16614,N_16747);
nor U16832 (N_16832,N_16716,N_16631);
or U16833 (N_16833,N_16507,N_16630);
xnor U16834 (N_16834,N_16566,N_16567);
xor U16835 (N_16835,N_16651,N_16645);
xnor U16836 (N_16836,N_16593,N_16639);
nand U16837 (N_16837,N_16626,N_16694);
nor U16838 (N_16838,N_16501,N_16610);
and U16839 (N_16839,N_16622,N_16670);
xnor U16840 (N_16840,N_16617,N_16633);
and U16841 (N_16841,N_16727,N_16537);
nand U16842 (N_16842,N_16722,N_16624);
nor U16843 (N_16843,N_16505,N_16640);
nand U16844 (N_16844,N_16585,N_16672);
or U16845 (N_16845,N_16748,N_16564);
nand U16846 (N_16846,N_16544,N_16667);
and U16847 (N_16847,N_16550,N_16500);
nor U16848 (N_16848,N_16693,N_16620);
nand U16849 (N_16849,N_16588,N_16603);
xnor U16850 (N_16850,N_16668,N_16524);
or U16851 (N_16851,N_16688,N_16599);
or U16852 (N_16852,N_16734,N_16628);
xor U16853 (N_16853,N_16671,N_16601);
nand U16854 (N_16854,N_16595,N_16711);
nor U16855 (N_16855,N_16503,N_16663);
nand U16856 (N_16856,N_16536,N_16621);
xnor U16857 (N_16857,N_16678,N_16502);
xor U16858 (N_16858,N_16697,N_16560);
nand U16859 (N_16859,N_16582,N_16686);
and U16860 (N_16860,N_16740,N_16535);
nor U16861 (N_16861,N_16554,N_16589);
or U16862 (N_16862,N_16508,N_16598);
nand U16863 (N_16863,N_16749,N_16702);
nand U16864 (N_16864,N_16642,N_16647);
xor U16865 (N_16865,N_16669,N_16743);
and U16866 (N_16866,N_16584,N_16563);
xor U16867 (N_16867,N_16732,N_16522);
xnor U16868 (N_16868,N_16646,N_16526);
nor U16869 (N_16869,N_16692,N_16637);
or U16870 (N_16870,N_16521,N_16674);
and U16871 (N_16871,N_16714,N_16541);
and U16872 (N_16872,N_16569,N_16644);
nand U16873 (N_16873,N_16551,N_16679);
and U16874 (N_16874,N_16600,N_16739);
xnor U16875 (N_16875,N_16742,N_16736);
nor U16876 (N_16876,N_16665,N_16540);
xnor U16877 (N_16877,N_16526,N_16652);
or U16878 (N_16878,N_16745,N_16630);
xnor U16879 (N_16879,N_16659,N_16529);
nand U16880 (N_16880,N_16628,N_16691);
or U16881 (N_16881,N_16650,N_16504);
xor U16882 (N_16882,N_16526,N_16574);
and U16883 (N_16883,N_16626,N_16573);
xnor U16884 (N_16884,N_16520,N_16521);
nand U16885 (N_16885,N_16674,N_16568);
nor U16886 (N_16886,N_16578,N_16706);
nand U16887 (N_16887,N_16569,N_16523);
and U16888 (N_16888,N_16677,N_16668);
and U16889 (N_16889,N_16731,N_16739);
or U16890 (N_16890,N_16631,N_16557);
or U16891 (N_16891,N_16505,N_16588);
xnor U16892 (N_16892,N_16711,N_16691);
nand U16893 (N_16893,N_16642,N_16503);
or U16894 (N_16894,N_16672,N_16686);
nor U16895 (N_16895,N_16648,N_16543);
and U16896 (N_16896,N_16699,N_16561);
and U16897 (N_16897,N_16599,N_16523);
nand U16898 (N_16898,N_16680,N_16598);
and U16899 (N_16899,N_16636,N_16568);
nor U16900 (N_16900,N_16702,N_16648);
nor U16901 (N_16901,N_16737,N_16599);
or U16902 (N_16902,N_16735,N_16704);
or U16903 (N_16903,N_16659,N_16728);
nand U16904 (N_16904,N_16746,N_16667);
xnor U16905 (N_16905,N_16506,N_16693);
or U16906 (N_16906,N_16736,N_16744);
nand U16907 (N_16907,N_16593,N_16740);
or U16908 (N_16908,N_16616,N_16723);
nor U16909 (N_16909,N_16577,N_16643);
xor U16910 (N_16910,N_16664,N_16567);
nand U16911 (N_16911,N_16641,N_16551);
xnor U16912 (N_16912,N_16723,N_16548);
or U16913 (N_16913,N_16593,N_16738);
nand U16914 (N_16914,N_16532,N_16720);
and U16915 (N_16915,N_16655,N_16707);
or U16916 (N_16916,N_16672,N_16627);
xor U16917 (N_16917,N_16577,N_16627);
nor U16918 (N_16918,N_16580,N_16740);
nand U16919 (N_16919,N_16637,N_16586);
or U16920 (N_16920,N_16696,N_16702);
xnor U16921 (N_16921,N_16680,N_16736);
xor U16922 (N_16922,N_16609,N_16606);
xor U16923 (N_16923,N_16633,N_16524);
xor U16924 (N_16924,N_16740,N_16598);
and U16925 (N_16925,N_16600,N_16669);
and U16926 (N_16926,N_16597,N_16531);
nor U16927 (N_16927,N_16519,N_16570);
nor U16928 (N_16928,N_16580,N_16519);
nor U16929 (N_16929,N_16631,N_16728);
and U16930 (N_16930,N_16634,N_16679);
xnor U16931 (N_16931,N_16730,N_16749);
and U16932 (N_16932,N_16500,N_16553);
nor U16933 (N_16933,N_16666,N_16725);
nor U16934 (N_16934,N_16538,N_16716);
nand U16935 (N_16935,N_16637,N_16700);
nor U16936 (N_16936,N_16591,N_16532);
nor U16937 (N_16937,N_16526,N_16744);
or U16938 (N_16938,N_16581,N_16673);
xnor U16939 (N_16939,N_16508,N_16573);
nor U16940 (N_16940,N_16702,N_16528);
or U16941 (N_16941,N_16682,N_16612);
and U16942 (N_16942,N_16656,N_16688);
nor U16943 (N_16943,N_16660,N_16685);
and U16944 (N_16944,N_16562,N_16644);
or U16945 (N_16945,N_16508,N_16648);
nand U16946 (N_16946,N_16727,N_16680);
xor U16947 (N_16947,N_16658,N_16594);
and U16948 (N_16948,N_16708,N_16525);
nor U16949 (N_16949,N_16695,N_16646);
nor U16950 (N_16950,N_16557,N_16530);
xnor U16951 (N_16951,N_16744,N_16573);
nand U16952 (N_16952,N_16573,N_16512);
or U16953 (N_16953,N_16644,N_16738);
nand U16954 (N_16954,N_16619,N_16527);
nand U16955 (N_16955,N_16576,N_16670);
and U16956 (N_16956,N_16518,N_16696);
nand U16957 (N_16957,N_16580,N_16680);
or U16958 (N_16958,N_16663,N_16609);
and U16959 (N_16959,N_16703,N_16627);
and U16960 (N_16960,N_16540,N_16657);
nor U16961 (N_16961,N_16646,N_16693);
nand U16962 (N_16962,N_16705,N_16729);
xor U16963 (N_16963,N_16712,N_16648);
or U16964 (N_16964,N_16509,N_16684);
nand U16965 (N_16965,N_16743,N_16740);
and U16966 (N_16966,N_16583,N_16684);
or U16967 (N_16967,N_16580,N_16707);
xnor U16968 (N_16968,N_16691,N_16513);
and U16969 (N_16969,N_16515,N_16628);
and U16970 (N_16970,N_16708,N_16621);
nor U16971 (N_16971,N_16737,N_16512);
nand U16972 (N_16972,N_16657,N_16620);
xor U16973 (N_16973,N_16677,N_16687);
and U16974 (N_16974,N_16745,N_16696);
and U16975 (N_16975,N_16707,N_16694);
nand U16976 (N_16976,N_16710,N_16650);
and U16977 (N_16977,N_16642,N_16578);
or U16978 (N_16978,N_16575,N_16714);
or U16979 (N_16979,N_16719,N_16507);
nor U16980 (N_16980,N_16541,N_16603);
or U16981 (N_16981,N_16715,N_16661);
nand U16982 (N_16982,N_16569,N_16607);
nor U16983 (N_16983,N_16716,N_16717);
nand U16984 (N_16984,N_16672,N_16643);
xnor U16985 (N_16985,N_16628,N_16657);
nand U16986 (N_16986,N_16677,N_16591);
nand U16987 (N_16987,N_16569,N_16616);
and U16988 (N_16988,N_16597,N_16608);
nand U16989 (N_16989,N_16563,N_16673);
and U16990 (N_16990,N_16529,N_16727);
or U16991 (N_16991,N_16669,N_16618);
xor U16992 (N_16992,N_16691,N_16704);
nor U16993 (N_16993,N_16679,N_16552);
or U16994 (N_16994,N_16660,N_16591);
and U16995 (N_16995,N_16594,N_16559);
nand U16996 (N_16996,N_16530,N_16722);
and U16997 (N_16997,N_16632,N_16621);
nand U16998 (N_16998,N_16570,N_16533);
xnor U16999 (N_16999,N_16579,N_16574);
and U17000 (N_17000,N_16909,N_16820);
or U17001 (N_17001,N_16775,N_16889);
nor U17002 (N_17002,N_16761,N_16865);
nand U17003 (N_17003,N_16811,N_16930);
nor U17004 (N_17004,N_16933,N_16756);
nor U17005 (N_17005,N_16994,N_16784);
and U17006 (N_17006,N_16802,N_16814);
xnor U17007 (N_17007,N_16962,N_16827);
and U17008 (N_17008,N_16831,N_16763);
nand U17009 (N_17009,N_16760,N_16929);
nor U17010 (N_17010,N_16935,N_16970);
nand U17011 (N_17011,N_16984,N_16927);
nor U17012 (N_17012,N_16958,N_16950);
and U17013 (N_17013,N_16780,N_16982);
or U17014 (N_17014,N_16914,N_16836);
and U17015 (N_17015,N_16967,N_16995);
nand U17016 (N_17016,N_16875,N_16895);
nor U17017 (N_17017,N_16932,N_16871);
nor U17018 (N_17018,N_16826,N_16867);
or U17019 (N_17019,N_16953,N_16781);
and U17020 (N_17020,N_16808,N_16916);
xnor U17021 (N_17021,N_16908,N_16937);
nand U17022 (N_17022,N_16870,N_16860);
nand U17023 (N_17023,N_16806,N_16988);
nor U17024 (N_17024,N_16855,N_16766);
nand U17025 (N_17025,N_16825,N_16948);
or U17026 (N_17026,N_16900,N_16942);
or U17027 (N_17027,N_16877,N_16862);
nand U17028 (N_17028,N_16898,N_16846);
nor U17029 (N_17029,N_16949,N_16944);
and U17030 (N_17030,N_16754,N_16828);
or U17031 (N_17031,N_16985,N_16856);
and U17032 (N_17032,N_16829,N_16896);
nand U17033 (N_17033,N_16945,N_16818);
nor U17034 (N_17034,N_16920,N_16997);
or U17035 (N_17035,N_16750,N_16864);
nor U17036 (N_17036,N_16847,N_16922);
nor U17037 (N_17037,N_16803,N_16777);
xnor U17038 (N_17038,N_16892,N_16843);
and U17039 (N_17039,N_16790,N_16773);
nor U17040 (N_17040,N_16786,N_16854);
or U17041 (N_17041,N_16996,N_16897);
or U17042 (N_17042,N_16931,N_16963);
nand U17043 (N_17043,N_16800,N_16981);
or U17044 (N_17044,N_16793,N_16770);
xor U17045 (N_17045,N_16751,N_16753);
and U17046 (N_17046,N_16863,N_16907);
xor U17047 (N_17047,N_16762,N_16795);
nor U17048 (N_17048,N_16879,N_16835);
xnor U17049 (N_17049,N_16768,N_16926);
and U17050 (N_17050,N_16910,N_16921);
and U17051 (N_17051,N_16913,N_16817);
nand U17052 (N_17052,N_16964,N_16839);
or U17053 (N_17053,N_16960,N_16911);
nand U17054 (N_17054,N_16796,N_16974);
nand U17055 (N_17055,N_16801,N_16785);
and U17056 (N_17056,N_16901,N_16774);
nor U17057 (N_17057,N_16979,N_16906);
nor U17058 (N_17058,N_16805,N_16936);
nor U17059 (N_17059,N_16955,N_16853);
and U17060 (N_17060,N_16886,N_16788);
xor U17061 (N_17061,N_16815,N_16765);
nor U17062 (N_17062,N_16797,N_16833);
or U17063 (N_17063,N_16842,N_16983);
or U17064 (N_17064,N_16946,N_16961);
or U17065 (N_17065,N_16787,N_16965);
or U17066 (N_17066,N_16973,N_16776);
xor U17067 (N_17067,N_16872,N_16799);
nor U17068 (N_17068,N_16992,N_16903);
and U17069 (N_17069,N_16893,N_16923);
nor U17070 (N_17070,N_16940,N_16858);
or U17071 (N_17071,N_16852,N_16755);
xor U17072 (N_17072,N_16837,N_16758);
nand U17073 (N_17073,N_16759,N_16822);
and U17074 (N_17074,N_16959,N_16977);
and U17075 (N_17075,N_16838,N_16899);
nand U17076 (N_17076,N_16915,N_16824);
nor U17077 (N_17077,N_16832,N_16925);
nand U17078 (N_17078,N_16809,N_16885);
xor U17079 (N_17079,N_16989,N_16968);
xnor U17080 (N_17080,N_16873,N_16792);
nand U17081 (N_17081,N_16987,N_16868);
nor U17082 (N_17082,N_16840,N_16912);
nor U17083 (N_17083,N_16804,N_16998);
nand U17084 (N_17084,N_16807,N_16869);
nand U17085 (N_17085,N_16845,N_16918);
xor U17086 (N_17086,N_16859,N_16857);
and U17087 (N_17087,N_16993,N_16849);
or U17088 (N_17088,N_16991,N_16810);
nand U17089 (N_17089,N_16888,N_16999);
nand U17090 (N_17090,N_16816,N_16794);
or U17091 (N_17091,N_16894,N_16941);
nor U17092 (N_17092,N_16841,N_16769);
nand U17093 (N_17093,N_16813,N_16943);
or U17094 (N_17094,N_16851,N_16902);
nor U17095 (N_17095,N_16812,N_16767);
nand U17096 (N_17096,N_16971,N_16891);
xor U17097 (N_17097,N_16821,N_16772);
or U17098 (N_17098,N_16934,N_16905);
or U17099 (N_17099,N_16783,N_16952);
xnor U17100 (N_17100,N_16972,N_16938);
nand U17101 (N_17101,N_16887,N_16764);
nand U17102 (N_17102,N_16830,N_16917);
nand U17103 (N_17103,N_16844,N_16939);
and U17104 (N_17104,N_16834,N_16876);
or U17105 (N_17105,N_16771,N_16969);
nor U17106 (N_17106,N_16861,N_16976);
or U17107 (N_17107,N_16890,N_16947);
nor U17108 (N_17108,N_16819,N_16874);
nand U17109 (N_17109,N_16848,N_16978);
and U17110 (N_17110,N_16919,N_16954);
and U17111 (N_17111,N_16878,N_16823);
xor U17112 (N_17112,N_16778,N_16928);
nor U17113 (N_17113,N_16986,N_16904);
and U17114 (N_17114,N_16951,N_16884);
nand U17115 (N_17115,N_16882,N_16779);
or U17116 (N_17116,N_16980,N_16956);
nor U17117 (N_17117,N_16850,N_16798);
xor U17118 (N_17118,N_16957,N_16880);
nand U17119 (N_17119,N_16990,N_16752);
xor U17120 (N_17120,N_16782,N_16924);
and U17121 (N_17121,N_16789,N_16757);
nor U17122 (N_17122,N_16881,N_16791);
and U17123 (N_17123,N_16966,N_16975);
nor U17124 (N_17124,N_16866,N_16883);
xor U17125 (N_17125,N_16895,N_16815);
or U17126 (N_17126,N_16851,N_16970);
or U17127 (N_17127,N_16965,N_16756);
or U17128 (N_17128,N_16952,N_16767);
or U17129 (N_17129,N_16762,N_16846);
nand U17130 (N_17130,N_16754,N_16964);
nand U17131 (N_17131,N_16822,N_16870);
and U17132 (N_17132,N_16809,N_16839);
nor U17133 (N_17133,N_16946,N_16945);
nand U17134 (N_17134,N_16830,N_16954);
nor U17135 (N_17135,N_16918,N_16924);
nor U17136 (N_17136,N_16818,N_16925);
nand U17137 (N_17137,N_16870,N_16924);
xor U17138 (N_17138,N_16794,N_16835);
nor U17139 (N_17139,N_16787,N_16797);
or U17140 (N_17140,N_16904,N_16944);
or U17141 (N_17141,N_16981,N_16769);
xor U17142 (N_17142,N_16998,N_16904);
or U17143 (N_17143,N_16878,N_16817);
nand U17144 (N_17144,N_16953,N_16895);
and U17145 (N_17145,N_16895,N_16986);
or U17146 (N_17146,N_16750,N_16897);
and U17147 (N_17147,N_16777,N_16995);
and U17148 (N_17148,N_16863,N_16785);
and U17149 (N_17149,N_16935,N_16908);
and U17150 (N_17150,N_16942,N_16878);
or U17151 (N_17151,N_16776,N_16772);
or U17152 (N_17152,N_16923,N_16854);
nor U17153 (N_17153,N_16773,N_16771);
or U17154 (N_17154,N_16980,N_16996);
nor U17155 (N_17155,N_16870,N_16809);
nor U17156 (N_17156,N_16893,N_16935);
nand U17157 (N_17157,N_16866,N_16971);
xor U17158 (N_17158,N_16988,N_16836);
nor U17159 (N_17159,N_16955,N_16986);
or U17160 (N_17160,N_16902,N_16778);
nor U17161 (N_17161,N_16797,N_16992);
or U17162 (N_17162,N_16927,N_16905);
nand U17163 (N_17163,N_16919,N_16781);
nand U17164 (N_17164,N_16958,N_16805);
nor U17165 (N_17165,N_16845,N_16958);
nand U17166 (N_17166,N_16789,N_16793);
or U17167 (N_17167,N_16878,N_16886);
nor U17168 (N_17168,N_16990,N_16971);
nor U17169 (N_17169,N_16787,N_16872);
or U17170 (N_17170,N_16757,N_16918);
xor U17171 (N_17171,N_16987,N_16849);
xnor U17172 (N_17172,N_16959,N_16941);
nor U17173 (N_17173,N_16903,N_16947);
xnor U17174 (N_17174,N_16953,N_16975);
xnor U17175 (N_17175,N_16756,N_16964);
or U17176 (N_17176,N_16922,N_16938);
xor U17177 (N_17177,N_16944,N_16845);
and U17178 (N_17178,N_16896,N_16848);
and U17179 (N_17179,N_16917,N_16921);
nor U17180 (N_17180,N_16879,N_16979);
or U17181 (N_17181,N_16900,N_16940);
xor U17182 (N_17182,N_16752,N_16779);
xnor U17183 (N_17183,N_16770,N_16775);
xnor U17184 (N_17184,N_16840,N_16849);
nor U17185 (N_17185,N_16898,N_16824);
and U17186 (N_17186,N_16760,N_16871);
nand U17187 (N_17187,N_16820,N_16989);
nand U17188 (N_17188,N_16757,N_16829);
or U17189 (N_17189,N_16815,N_16776);
or U17190 (N_17190,N_16870,N_16946);
xor U17191 (N_17191,N_16931,N_16946);
and U17192 (N_17192,N_16883,N_16841);
nand U17193 (N_17193,N_16957,N_16906);
nor U17194 (N_17194,N_16771,N_16967);
xnor U17195 (N_17195,N_16902,N_16756);
and U17196 (N_17196,N_16872,N_16934);
and U17197 (N_17197,N_16934,N_16962);
and U17198 (N_17198,N_16761,N_16785);
nand U17199 (N_17199,N_16989,N_16927);
or U17200 (N_17200,N_16777,N_16960);
xor U17201 (N_17201,N_16914,N_16971);
nand U17202 (N_17202,N_16761,N_16884);
nand U17203 (N_17203,N_16793,N_16873);
xnor U17204 (N_17204,N_16775,N_16931);
nor U17205 (N_17205,N_16973,N_16750);
xnor U17206 (N_17206,N_16781,N_16882);
nor U17207 (N_17207,N_16819,N_16936);
xor U17208 (N_17208,N_16946,N_16770);
and U17209 (N_17209,N_16962,N_16837);
nor U17210 (N_17210,N_16752,N_16830);
or U17211 (N_17211,N_16907,N_16949);
nand U17212 (N_17212,N_16780,N_16957);
nand U17213 (N_17213,N_16905,N_16953);
and U17214 (N_17214,N_16839,N_16960);
nand U17215 (N_17215,N_16849,N_16768);
xor U17216 (N_17216,N_16957,N_16882);
xnor U17217 (N_17217,N_16862,N_16837);
nor U17218 (N_17218,N_16961,N_16960);
and U17219 (N_17219,N_16809,N_16806);
or U17220 (N_17220,N_16907,N_16855);
nor U17221 (N_17221,N_16891,N_16758);
and U17222 (N_17222,N_16904,N_16956);
or U17223 (N_17223,N_16790,N_16856);
nor U17224 (N_17224,N_16964,N_16969);
nor U17225 (N_17225,N_16906,N_16905);
or U17226 (N_17226,N_16980,N_16905);
or U17227 (N_17227,N_16851,N_16959);
and U17228 (N_17228,N_16910,N_16947);
and U17229 (N_17229,N_16834,N_16825);
nor U17230 (N_17230,N_16924,N_16769);
nand U17231 (N_17231,N_16932,N_16798);
nor U17232 (N_17232,N_16801,N_16796);
or U17233 (N_17233,N_16886,N_16777);
xnor U17234 (N_17234,N_16934,N_16786);
and U17235 (N_17235,N_16976,N_16827);
xor U17236 (N_17236,N_16950,N_16884);
and U17237 (N_17237,N_16853,N_16766);
nor U17238 (N_17238,N_16937,N_16864);
nor U17239 (N_17239,N_16801,N_16935);
nand U17240 (N_17240,N_16827,N_16793);
nand U17241 (N_17241,N_16821,N_16934);
nand U17242 (N_17242,N_16861,N_16783);
or U17243 (N_17243,N_16980,N_16904);
or U17244 (N_17244,N_16929,N_16805);
and U17245 (N_17245,N_16831,N_16891);
or U17246 (N_17246,N_16756,N_16993);
or U17247 (N_17247,N_16987,N_16871);
nor U17248 (N_17248,N_16914,N_16759);
xor U17249 (N_17249,N_16845,N_16976);
xnor U17250 (N_17250,N_17140,N_17212);
and U17251 (N_17251,N_17005,N_17168);
nand U17252 (N_17252,N_17178,N_17025);
nand U17253 (N_17253,N_17095,N_17017);
or U17254 (N_17254,N_17052,N_17021);
and U17255 (N_17255,N_17041,N_17231);
and U17256 (N_17256,N_17042,N_17000);
xnor U17257 (N_17257,N_17215,N_17228);
and U17258 (N_17258,N_17121,N_17176);
and U17259 (N_17259,N_17109,N_17039);
and U17260 (N_17260,N_17057,N_17242);
or U17261 (N_17261,N_17164,N_17125);
and U17262 (N_17262,N_17110,N_17193);
and U17263 (N_17263,N_17063,N_17093);
or U17264 (N_17264,N_17237,N_17236);
and U17265 (N_17265,N_17217,N_17013);
or U17266 (N_17266,N_17006,N_17122);
nor U17267 (N_17267,N_17081,N_17153);
xor U17268 (N_17268,N_17009,N_17015);
xor U17269 (N_17269,N_17221,N_17070);
nand U17270 (N_17270,N_17126,N_17055);
nand U17271 (N_17271,N_17019,N_17024);
nor U17272 (N_17272,N_17148,N_17112);
xnor U17273 (N_17273,N_17018,N_17048);
xor U17274 (N_17274,N_17056,N_17049);
nor U17275 (N_17275,N_17145,N_17249);
or U17276 (N_17276,N_17199,N_17062);
or U17277 (N_17277,N_17053,N_17181);
nor U17278 (N_17278,N_17031,N_17119);
xor U17279 (N_17279,N_17232,N_17149);
and U17280 (N_17280,N_17117,N_17129);
or U17281 (N_17281,N_17098,N_17034);
or U17282 (N_17282,N_17100,N_17014);
or U17283 (N_17283,N_17061,N_17083);
and U17284 (N_17284,N_17194,N_17162);
or U17285 (N_17285,N_17160,N_17043);
or U17286 (N_17286,N_17036,N_17209);
and U17287 (N_17287,N_17188,N_17071);
xnor U17288 (N_17288,N_17208,N_17045);
nand U17289 (N_17289,N_17084,N_17183);
xor U17290 (N_17290,N_17074,N_17127);
and U17291 (N_17291,N_17227,N_17218);
xor U17292 (N_17292,N_17147,N_17051);
nand U17293 (N_17293,N_17196,N_17174);
and U17294 (N_17294,N_17097,N_17244);
nor U17295 (N_17295,N_17115,N_17004);
and U17296 (N_17296,N_17046,N_17247);
nor U17297 (N_17297,N_17220,N_17152);
nand U17298 (N_17298,N_17184,N_17170);
xor U17299 (N_17299,N_17177,N_17230);
and U17300 (N_17300,N_17060,N_17202);
or U17301 (N_17301,N_17223,N_17066);
nand U17302 (N_17302,N_17191,N_17132);
nor U17303 (N_17303,N_17150,N_17204);
and U17304 (N_17304,N_17102,N_17225);
nand U17305 (N_17305,N_17107,N_17154);
or U17306 (N_17306,N_17101,N_17233);
and U17307 (N_17307,N_17085,N_17011);
nand U17308 (N_17308,N_17035,N_17136);
or U17309 (N_17309,N_17173,N_17141);
nor U17310 (N_17310,N_17038,N_17246);
and U17311 (N_17311,N_17167,N_17206);
xor U17312 (N_17312,N_17207,N_17026);
xor U17313 (N_17313,N_17216,N_17086);
xnor U17314 (N_17314,N_17108,N_17090);
xor U17315 (N_17315,N_17180,N_17075);
or U17316 (N_17316,N_17235,N_17187);
nor U17317 (N_17317,N_17158,N_17032);
xnor U17318 (N_17318,N_17128,N_17142);
and U17319 (N_17319,N_17137,N_17096);
nor U17320 (N_17320,N_17016,N_17205);
or U17321 (N_17321,N_17028,N_17088);
or U17322 (N_17322,N_17076,N_17171);
xnor U17323 (N_17323,N_17190,N_17003);
nand U17324 (N_17324,N_17106,N_17001);
and U17325 (N_17325,N_17224,N_17238);
nor U17326 (N_17326,N_17116,N_17118);
xor U17327 (N_17327,N_17058,N_17089);
nand U17328 (N_17328,N_17144,N_17213);
or U17329 (N_17329,N_17010,N_17033);
nand U17330 (N_17330,N_17064,N_17211);
nor U17331 (N_17331,N_17087,N_17134);
and U17332 (N_17332,N_17037,N_17091);
nor U17333 (N_17333,N_17186,N_17189);
nor U17334 (N_17334,N_17080,N_17007);
nor U17335 (N_17335,N_17114,N_17092);
and U17336 (N_17336,N_17226,N_17082);
or U17337 (N_17337,N_17040,N_17012);
and U17338 (N_17338,N_17192,N_17068);
nor U17339 (N_17339,N_17222,N_17094);
xor U17340 (N_17340,N_17104,N_17054);
and U17341 (N_17341,N_17241,N_17139);
nand U17342 (N_17342,N_17065,N_17023);
and U17343 (N_17343,N_17229,N_17203);
nor U17344 (N_17344,N_17077,N_17103);
xnor U17345 (N_17345,N_17197,N_17072);
xor U17346 (N_17346,N_17138,N_17185);
or U17347 (N_17347,N_17044,N_17111);
nand U17348 (N_17348,N_17133,N_17002);
xor U17349 (N_17349,N_17234,N_17008);
and U17350 (N_17350,N_17210,N_17155);
or U17351 (N_17351,N_17163,N_17050);
nand U17352 (N_17352,N_17157,N_17214);
xor U17353 (N_17353,N_17146,N_17143);
or U17354 (N_17354,N_17067,N_17047);
xor U17355 (N_17355,N_17248,N_17240);
nand U17356 (N_17356,N_17069,N_17156);
nand U17357 (N_17357,N_17172,N_17120);
nor U17358 (N_17358,N_17105,N_17165);
nand U17359 (N_17359,N_17175,N_17131);
or U17360 (N_17360,N_17079,N_17099);
xnor U17361 (N_17361,N_17239,N_17124);
xor U17362 (N_17362,N_17151,N_17135);
xnor U17363 (N_17363,N_17166,N_17179);
nand U17364 (N_17364,N_17130,N_17030);
xor U17365 (N_17365,N_17078,N_17201);
nand U17366 (N_17366,N_17022,N_17243);
and U17367 (N_17367,N_17195,N_17219);
and U17368 (N_17368,N_17169,N_17113);
or U17369 (N_17369,N_17059,N_17161);
or U17370 (N_17370,N_17198,N_17123);
nor U17371 (N_17371,N_17073,N_17182);
xor U17372 (N_17372,N_17027,N_17245);
xor U17373 (N_17373,N_17029,N_17159);
nor U17374 (N_17374,N_17020,N_17200);
or U17375 (N_17375,N_17142,N_17211);
nand U17376 (N_17376,N_17163,N_17122);
or U17377 (N_17377,N_17239,N_17089);
and U17378 (N_17378,N_17024,N_17205);
xor U17379 (N_17379,N_17205,N_17087);
xor U17380 (N_17380,N_17068,N_17169);
and U17381 (N_17381,N_17205,N_17153);
nand U17382 (N_17382,N_17072,N_17120);
nor U17383 (N_17383,N_17057,N_17225);
nor U17384 (N_17384,N_17080,N_17011);
or U17385 (N_17385,N_17241,N_17070);
xnor U17386 (N_17386,N_17041,N_17220);
nand U17387 (N_17387,N_17146,N_17130);
xnor U17388 (N_17388,N_17151,N_17220);
nor U17389 (N_17389,N_17230,N_17139);
or U17390 (N_17390,N_17107,N_17025);
and U17391 (N_17391,N_17019,N_17122);
nor U17392 (N_17392,N_17034,N_17025);
nand U17393 (N_17393,N_17235,N_17021);
or U17394 (N_17394,N_17227,N_17146);
xor U17395 (N_17395,N_17002,N_17052);
xor U17396 (N_17396,N_17243,N_17188);
or U17397 (N_17397,N_17160,N_17119);
or U17398 (N_17398,N_17194,N_17205);
nand U17399 (N_17399,N_17053,N_17103);
nor U17400 (N_17400,N_17175,N_17117);
nand U17401 (N_17401,N_17248,N_17175);
or U17402 (N_17402,N_17197,N_17052);
or U17403 (N_17403,N_17154,N_17026);
nand U17404 (N_17404,N_17148,N_17205);
nand U17405 (N_17405,N_17141,N_17157);
xor U17406 (N_17406,N_17005,N_17136);
nor U17407 (N_17407,N_17201,N_17075);
nand U17408 (N_17408,N_17248,N_17183);
or U17409 (N_17409,N_17214,N_17205);
nand U17410 (N_17410,N_17150,N_17152);
nand U17411 (N_17411,N_17125,N_17070);
or U17412 (N_17412,N_17205,N_17122);
or U17413 (N_17413,N_17058,N_17070);
and U17414 (N_17414,N_17247,N_17170);
and U17415 (N_17415,N_17174,N_17017);
nand U17416 (N_17416,N_17090,N_17058);
xnor U17417 (N_17417,N_17188,N_17205);
and U17418 (N_17418,N_17172,N_17245);
nand U17419 (N_17419,N_17238,N_17064);
nor U17420 (N_17420,N_17034,N_17188);
or U17421 (N_17421,N_17214,N_17120);
and U17422 (N_17422,N_17164,N_17195);
xnor U17423 (N_17423,N_17116,N_17035);
nand U17424 (N_17424,N_17056,N_17211);
and U17425 (N_17425,N_17179,N_17039);
nand U17426 (N_17426,N_17007,N_17020);
and U17427 (N_17427,N_17076,N_17044);
nor U17428 (N_17428,N_17073,N_17008);
nor U17429 (N_17429,N_17113,N_17237);
nor U17430 (N_17430,N_17215,N_17147);
and U17431 (N_17431,N_17184,N_17196);
and U17432 (N_17432,N_17030,N_17033);
nand U17433 (N_17433,N_17000,N_17244);
xnor U17434 (N_17434,N_17141,N_17153);
xnor U17435 (N_17435,N_17076,N_17118);
or U17436 (N_17436,N_17015,N_17131);
nor U17437 (N_17437,N_17073,N_17147);
nand U17438 (N_17438,N_17039,N_17201);
xor U17439 (N_17439,N_17181,N_17007);
nand U17440 (N_17440,N_17136,N_17061);
and U17441 (N_17441,N_17230,N_17095);
or U17442 (N_17442,N_17167,N_17179);
or U17443 (N_17443,N_17025,N_17069);
xnor U17444 (N_17444,N_17043,N_17063);
xnor U17445 (N_17445,N_17020,N_17150);
xnor U17446 (N_17446,N_17141,N_17065);
and U17447 (N_17447,N_17025,N_17143);
or U17448 (N_17448,N_17165,N_17002);
nand U17449 (N_17449,N_17060,N_17225);
or U17450 (N_17450,N_17049,N_17117);
and U17451 (N_17451,N_17237,N_17135);
nand U17452 (N_17452,N_17045,N_17108);
nor U17453 (N_17453,N_17042,N_17172);
nor U17454 (N_17454,N_17047,N_17194);
or U17455 (N_17455,N_17146,N_17096);
xor U17456 (N_17456,N_17043,N_17216);
or U17457 (N_17457,N_17189,N_17000);
nor U17458 (N_17458,N_17137,N_17004);
xor U17459 (N_17459,N_17030,N_17243);
and U17460 (N_17460,N_17115,N_17198);
nor U17461 (N_17461,N_17240,N_17034);
nand U17462 (N_17462,N_17208,N_17213);
xnor U17463 (N_17463,N_17050,N_17221);
or U17464 (N_17464,N_17142,N_17223);
and U17465 (N_17465,N_17008,N_17161);
nand U17466 (N_17466,N_17060,N_17092);
and U17467 (N_17467,N_17242,N_17108);
nand U17468 (N_17468,N_17032,N_17149);
and U17469 (N_17469,N_17248,N_17194);
xnor U17470 (N_17470,N_17073,N_17166);
xnor U17471 (N_17471,N_17158,N_17002);
nand U17472 (N_17472,N_17132,N_17084);
or U17473 (N_17473,N_17190,N_17124);
nor U17474 (N_17474,N_17019,N_17058);
and U17475 (N_17475,N_17030,N_17062);
nor U17476 (N_17476,N_17198,N_17073);
or U17477 (N_17477,N_17141,N_17124);
or U17478 (N_17478,N_17160,N_17233);
xnor U17479 (N_17479,N_17027,N_17135);
or U17480 (N_17480,N_17227,N_17151);
nand U17481 (N_17481,N_17143,N_17165);
nor U17482 (N_17482,N_17170,N_17148);
nor U17483 (N_17483,N_17119,N_17203);
nor U17484 (N_17484,N_17009,N_17165);
nand U17485 (N_17485,N_17214,N_17127);
nor U17486 (N_17486,N_17068,N_17230);
nor U17487 (N_17487,N_17095,N_17142);
nand U17488 (N_17488,N_17195,N_17139);
or U17489 (N_17489,N_17207,N_17181);
nor U17490 (N_17490,N_17005,N_17031);
nor U17491 (N_17491,N_17230,N_17200);
xnor U17492 (N_17492,N_17038,N_17178);
xor U17493 (N_17493,N_17118,N_17023);
or U17494 (N_17494,N_17038,N_17226);
nor U17495 (N_17495,N_17036,N_17002);
or U17496 (N_17496,N_17242,N_17079);
nor U17497 (N_17497,N_17100,N_17229);
and U17498 (N_17498,N_17221,N_17067);
or U17499 (N_17499,N_17004,N_17088);
and U17500 (N_17500,N_17274,N_17276);
and U17501 (N_17501,N_17319,N_17261);
xor U17502 (N_17502,N_17458,N_17372);
nand U17503 (N_17503,N_17471,N_17331);
and U17504 (N_17504,N_17295,N_17314);
and U17505 (N_17505,N_17491,N_17287);
and U17506 (N_17506,N_17288,N_17416);
nand U17507 (N_17507,N_17272,N_17452);
nor U17508 (N_17508,N_17353,N_17475);
nand U17509 (N_17509,N_17473,N_17489);
nand U17510 (N_17510,N_17270,N_17328);
nor U17511 (N_17511,N_17367,N_17482);
nor U17512 (N_17512,N_17398,N_17256);
and U17513 (N_17513,N_17459,N_17268);
xnor U17514 (N_17514,N_17356,N_17359);
nor U17515 (N_17515,N_17455,N_17321);
and U17516 (N_17516,N_17364,N_17439);
nand U17517 (N_17517,N_17376,N_17426);
or U17518 (N_17518,N_17349,N_17407);
nand U17519 (N_17519,N_17332,N_17454);
nor U17520 (N_17520,N_17291,N_17413);
and U17521 (N_17521,N_17290,N_17262);
and U17522 (N_17522,N_17487,N_17493);
nand U17523 (N_17523,N_17294,N_17365);
xnor U17524 (N_17524,N_17412,N_17438);
nand U17525 (N_17525,N_17307,N_17348);
nor U17526 (N_17526,N_17283,N_17345);
nor U17527 (N_17527,N_17476,N_17485);
and U17528 (N_17528,N_17440,N_17368);
and U17529 (N_17529,N_17460,N_17335);
xnor U17530 (N_17530,N_17255,N_17251);
xor U17531 (N_17531,N_17313,N_17496);
or U17532 (N_17532,N_17266,N_17343);
and U17533 (N_17533,N_17277,N_17379);
nand U17534 (N_17534,N_17263,N_17469);
and U17535 (N_17535,N_17380,N_17341);
xnor U17536 (N_17536,N_17339,N_17436);
nand U17537 (N_17537,N_17480,N_17453);
nand U17538 (N_17538,N_17435,N_17325);
nand U17539 (N_17539,N_17293,N_17405);
and U17540 (N_17540,N_17486,N_17378);
or U17541 (N_17541,N_17451,N_17479);
and U17542 (N_17542,N_17465,N_17468);
xor U17543 (N_17543,N_17397,N_17437);
xnor U17544 (N_17544,N_17267,N_17402);
nor U17545 (N_17545,N_17369,N_17415);
nand U17546 (N_17546,N_17420,N_17497);
and U17547 (N_17547,N_17279,N_17466);
or U17548 (N_17548,N_17389,N_17427);
nand U17549 (N_17549,N_17414,N_17252);
nand U17550 (N_17550,N_17396,N_17347);
or U17551 (N_17551,N_17474,N_17301);
nor U17552 (N_17552,N_17446,N_17334);
nand U17553 (N_17553,N_17271,N_17401);
and U17554 (N_17554,N_17385,N_17447);
and U17555 (N_17555,N_17406,N_17448);
nor U17556 (N_17556,N_17285,N_17442);
nand U17557 (N_17557,N_17377,N_17472);
nor U17558 (N_17558,N_17254,N_17352);
and U17559 (N_17559,N_17409,N_17302);
nand U17560 (N_17560,N_17375,N_17362);
xor U17561 (N_17561,N_17421,N_17417);
nor U17562 (N_17562,N_17400,N_17424);
xor U17563 (N_17563,N_17384,N_17269);
and U17564 (N_17564,N_17382,N_17445);
and U17565 (N_17565,N_17434,N_17253);
or U17566 (N_17566,N_17464,N_17483);
nand U17567 (N_17567,N_17373,N_17408);
nor U17568 (N_17568,N_17360,N_17296);
nor U17569 (N_17569,N_17257,N_17320);
nor U17570 (N_17570,N_17264,N_17383);
nor U17571 (N_17571,N_17284,N_17338);
nand U17572 (N_17572,N_17490,N_17404);
or U17573 (N_17573,N_17337,N_17333);
nor U17574 (N_17574,N_17392,N_17351);
xor U17575 (N_17575,N_17498,N_17323);
or U17576 (N_17576,N_17309,N_17278);
nand U17577 (N_17577,N_17258,N_17311);
nor U17578 (N_17578,N_17499,N_17327);
nor U17579 (N_17579,N_17428,N_17318);
nor U17580 (N_17580,N_17317,N_17342);
and U17581 (N_17581,N_17393,N_17456);
and U17582 (N_17582,N_17289,N_17322);
nor U17583 (N_17583,N_17336,N_17292);
nor U17584 (N_17584,N_17324,N_17273);
or U17585 (N_17585,N_17346,N_17403);
nor U17586 (N_17586,N_17488,N_17431);
nor U17587 (N_17587,N_17481,N_17363);
nand U17588 (N_17588,N_17250,N_17467);
xor U17589 (N_17589,N_17275,N_17361);
and U17590 (N_17590,N_17265,N_17441);
and U17591 (N_17591,N_17399,N_17316);
nor U17592 (N_17592,N_17304,N_17357);
and U17593 (N_17593,N_17388,N_17449);
and U17594 (N_17594,N_17450,N_17457);
and U17595 (N_17595,N_17330,N_17299);
or U17596 (N_17596,N_17366,N_17280);
and U17597 (N_17597,N_17430,N_17494);
nor U17598 (N_17598,N_17358,N_17390);
and U17599 (N_17599,N_17344,N_17298);
nand U17600 (N_17600,N_17418,N_17326);
and U17601 (N_17601,N_17419,N_17461);
nand U17602 (N_17602,N_17386,N_17300);
or U17603 (N_17603,N_17432,N_17395);
nand U17604 (N_17604,N_17286,N_17355);
nand U17605 (N_17605,N_17370,N_17306);
xnor U17606 (N_17606,N_17478,N_17297);
xor U17607 (N_17607,N_17312,N_17425);
nand U17608 (N_17608,N_17443,N_17282);
xor U17609 (N_17609,N_17423,N_17492);
and U17610 (N_17610,N_17354,N_17329);
nor U17611 (N_17611,N_17374,N_17340);
nand U17612 (N_17612,N_17462,N_17463);
and U17613 (N_17613,N_17422,N_17477);
or U17614 (N_17614,N_17371,N_17260);
or U17615 (N_17615,N_17381,N_17411);
or U17616 (N_17616,N_17305,N_17470);
nand U17617 (N_17617,N_17281,N_17387);
or U17618 (N_17618,N_17444,N_17308);
nand U17619 (N_17619,N_17303,N_17433);
xnor U17620 (N_17620,N_17391,N_17259);
and U17621 (N_17621,N_17429,N_17410);
nand U17622 (N_17622,N_17350,N_17315);
or U17623 (N_17623,N_17484,N_17394);
and U17624 (N_17624,N_17495,N_17310);
and U17625 (N_17625,N_17486,N_17268);
or U17626 (N_17626,N_17317,N_17454);
or U17627 (N_17627,N_17364,N_17309);
xnor U17628 (N_17628,N_17343,N_17272);
or U17629 (N_17629,N_17257,N_17463);
and U17630 (N_17630,N_17448,N_17386);
nand U17631 (N_17631,N_17481,N_17453);
xor U17632 (N_17632,N_17435,N_17371);
nor U17633 (N_17633,N_17496,N_17465);
or U17634 (N_17634,N_17486,N_17319);
and U17635 (N_17635,N_17417,N_17303);
nor U17636 (N_17636,N_17362,N_17437);
nand U17637 (N_17637,N_17257,N_17378);
nor U17638 (N_17638,N_17401,N_17263);
xnor U17639 (N_17639,N_17425,N_17322);
nor U17640 (N_17640,N_17403,N_17279);
or U17641 (N_17641,N_17464,N_17279);
or U17642 (N_17642,N_17430,N_17255);
xor U17643 (N_17643,N_17360,N_17495);
xor U17644 (N_17644,N_17412,N_17452);
and U17645 (N_17645,N_17490,N_17297);
or U17646 (N_17646,N_17320,N_17336);
nor U17647 (N_17647,N_17277,N_17294);
xor U17648 (N_17648,N_17358,N_17340);
and U17649 (N_17649,N_17267,N_17288);
xnor U17650 (N_17650,N_17256,N_17385);
nand U17651 (N_17651,N_17398,N_17304);
nor U17652 (N_17652,N_17400,N_17303);
and U17653 (N_17653,N_17302,N_17380);
xnor U17654 (N_17654,N_17277,N_17383);
nand U17655 (N_17655,N_17442,N_17344);
xor U17656 (N_17656,N_17490,N_17432);
nor U17657 (N_17657,N_17484,N_17439);
and U17658 (N_17658,N_17354,N_17469);
and U17659 (N_17659,N_17292,N_17258);
nand U17660 (N_17660,N_17424,N_17279);
or U17661 (N_17661,N_17391,N_17251);
or U17662 (N_17662,N_17358,N_17432);
nand U17663 (N_17663,N_17326,N_17299);
nor U17664 (N_17664,N_17361,N_17420);
or U17665 (N_17665,N_17308,N_17480);
nor U17666 (N_17666,N_17268,N_17350);
xnor U17667 (N_17667,N_17499,N_17494);
nand U17668 (N_17668,N_17471,N_17454);
nor U17669 (N_17669,N_17377,N_17312);
nor U17670 (N_17670,N_17446,N_17314);
and U17671 (N_17671,N_17319,N_17423);
or U17672 (N_17672,N_17261,N_17498);
nand U17673 (N_17673,N_17275,N_17325);
and U17674 (N_17674,N_17467,N_17440);
nor U17675 (N_17675,N_17397,N_17402);
and U17676 (N_17676,N_17465,N_17317);
or U17677 (N_17677,N_17472,N_17304);
xor U17678 (N_17678,N_17474,N_17333);
xor U17679 (N_17679,N_17373,N_17447);
or U17680 (N_17680,N_17394,N_17449);
and U17681 (N_17681,N_17321,N_17407);
and U17682 (N_17682,N_17300,N_17476);
nand U17683 (N_17683,N_17355,N_17283);
nor U17684 (N_17684,N_17375,N_17426);
nor U17685 (N_17685,N_17358,N_17310);
xor U17686 (N_17686,N_17301,N_17277);
or U17687 (N_17687,N_17468,N_17302);
xor U17688 (N_17688,N_17250,N_17299);
nor U17689 (N_17689,N_17297,N_17336);
and U17690 (N_17690,N_17391,N_17395);
xor U17691 (N_17691,N_17347,N_17471);
nor U17692 (N_17692,N_17304,N_17447);
and U17693 (N_17693,N_17449,N_17275);
xor U17694 (N_17694,N_17355,N_17317);
xnor U17695 (N_17695,N_17272,N_17331);
nand U17696 (N_17696,N_17283,N_17347);
xor U17697 (N_17697,N_17394,N_17413);
nor U17698 (N_17698,N_17496,N_17280);
and U17699 (N_17699,N_17309,N_17498);
nand U17700 (N_17700,N_17286,N_17390);
and U17701 (N_17701,N_17350,N_17275);
xor U17702 (N_17702,N_17329,N_17449);
xnor U17703 (N_17703,N_17483,N_17328);
and U17704 (N_17704,N_17435,N_17352);
and U17705 (N_17705,N_17395,N_17345);
nor U17706 (N_17706,N_17452,N_17332);
xor U17707 (N_17707,N_17264,N_17277);
nand U17708 (N_17708,N_17329,N_17352);
nand U17709 (N_17709,N_17255,N_17498);
xnor U17710 (N_17710,N_17254,N_17465);
or U17711 (N_17711,N_17311,N_17412);
and U17712 (N_17712,N_17309,N_17257);
or U17713 (N_17713,N_17292,N_17465);
xnor U17714 (N_17714,N_17338,N_17286);
xnor U17715 (N_17715,N_17483,N_17291);
or U17716 (N_17716,N_17479,N_17499);
or U17717 (N_17717,N_17481,N_17421);
or U17718 (N_17718,N_17327,N_17400);
or U17719 (N_17719,N_17398,N_17451);
or U17720 (N_17720,N_17338,N_17292);
and U17721 (N_17721,N_17422,N_17403);
and U17722 (N_17722,N_17438,N_17495);
and U17723 (N_17723,N_17426,N_17454);
xor U17724 (N_17724,N_17367,N_17304);
nand U17725 (N_17725,N_17374,N_17449);
or U17726 (N_17726,N_17482,N_17392);
nor U17727 (N_17727,N_17454,N_17444);
nand U17728 (N_17728,N_17323,N_17494);
nor U17729 (N_17729,N_17311,N_17422);
and U17730 (N_17730,N_17436,N_17461);
nand U17731 (N_17731,N_17439,N_17295);
xor U17732 (N_17732,N_17395,N_17328);
or U17733 (N_17733,N_17317,N_17387);
xnor U17734 (N_17734,N_17383,N_17346);
or U17735 (N_17735,N_17303,N_17311);
nor U17736 (N_17736,N_17331,N_17333);
and U17737 (N_17737,N_17309,N_17252);
xnor U17738 (N_17738,N_17490,N_17423);
xnor U17739 (N_17739,N_17263,N_17489);
or U17740 (N_17740,N_17267,N_17478);
or U17741 (N_17741,N_17457,N_17254);
or U17742 (N_17742,N_17277,N_17447);
xnor U17743 (N_17743,N_17325,N_17327);
and U17744 (N_17744,N_17278,N_17324);
nor U17745 (N_17745,N_17277,N_17435);
nor U17746 (N_17746,N_17325,N_17300);
and U17747 (N_17747,N_17438,N_17320);
nor U17748 (N_17748,N_17278,N_17297);
or U17749 (N_17749,N_17441,N_17376);
xnor U17750 (N_17750,N_17716,N_17585);
and U17751 (N_17751,N_17531,N_17602);
nand U17752 (N_17752,N_17623,N_17677);
xor U17753 (N_17753,N_17569,N_17596);
nor U17754 (N_17754,N_17699,N_17715);
nand U17755 (N_17755,N_17654,N_17719);
nor U17756 (N_17756,N_17624,N_17689);
xnor U17757 (N_17757,N_17705,N_17546);
nor U17758 (N_17758,N_17648,N_17685);
xor U17759 (N_17759,N_17671,N_17581);
nor U17760 (N_17760,N_17604,N_17527);
or U17761 (N_17761,N_17537,N_17698);
xnor U17762 (N_17762,N_17524,N_17579);
xor U17763 (N_17763,N_17574,N_17723);
and U17764 (N_17764,N_17506,N_17749);
xor U17765 (N_17765,N_17529,N_17707);
nand U17766 (N_17766,N_17739,N_17669);
xor U17767 (N_17767,N_17512,N_17678);
or U17768 (N_17768,N_17556,N_17712);
or U17769 (N_17769,N_17676,N_17727);
xor U17770 (N_17770,N_17608,N_17552);
and U17771 (N_17771,N_17570,N_17571);
and U17772 (N_17772,N_17639,N_17635);
nor U17773 (N_17773,N_17690,N_17728);
nor U17774 (N_17774,N_17706,N_17726);
nor U17775 (N_17775,N_17655,N_17652);
or U17776 (N_17776,N_17610,N_17734);
and U17777 (N_17777,N_17591,N_17516);
or U17778 (N_17778,N_17540,N_17566);
nor U17779 (N_17779,N_17643,N_17517);
or U17780 (N_17780,N_17600,N_17694);
nor U17781 (N_17781,N_17633,N_17651);
and U17782 (N_17782,N_17732,N_17733);
or U17783 (N_17783,N_17522,N_17586);
nor U17784 (N_17784,N_17684,N_17731);
xnor U17785 (N_17785,N_17553,N_17735);
or U17786 (N_17786,N_17644,N_17500);
and U17787 (N_17787,N_17704,N_17695);
and U17788 (N_17788,N_17597,N_17692);
nand U17789 (N_17789,N_17606,N_17557);
nor U17790 (N_17790,N_17621,N_17664);
nand U17791 (N_17791,N_17501,N_17673);
nand U17792 (N_17792,N_17642,N_17729);
or U17793 (N_17793,N_17550,N_17543);
nor U17794 (N_17794,N_17675,N_17658);
or U17795 (N_17795,N_17663,N_17555);
or U17796 (N_17796,N_17641,N_17584);
or U17797 (N_17797,N_17674,N_17708);
or U17798 (N_17798,N_17588,N_17737);
or U17799 (N_17799,N_17724,N_17554);
nand U17800 (N_17800,N_17713,N_17583);
nor U17801 (N_17801,N_17505,N_17587);
nand U17802 (N_17802,N_17741,N_17618);
nor U17803 (N_17803,N_17630,N_17525);
xnor U17804 (N_17804,N_17619,N_17509);
xor U17805 (N_17805,N_17541,N_17502);
nor U17806 (N_17806,N_17609,N_17535);
nor U17807 (N_17807,N_17738,N_17647);
nor U17808 (N_17808,N_17657,N_17665);
nand U17809 (N_17809,N_17565,N_17627);
nand U17810 (N_17810,N_17637,N_17598);
or U17811 (N_17811,N_17656,N_17526);
xor U17812 (N_17812,N_17701,N_17649);
xor U17813 (N_17813,N_17590,N_17616);
nand U17814 (N_17814,N_17575,N_17653);
nand U17815 (N_17815,N_17626,N_17717);
nor U17816 (N_17816,N_17612,N_17631);
or U17817 (N_17817,N_17672,N_17742);
nor U17818 (N_17818,N_17577,N_17686);
or U17819 (N_17819,N_17559,N_17528);
nor U17820 (N_17820,N_17746,N_17573);
nand U17821 (N_17821,N_17582,N_17564);
xor U17822 (N_17822,N_17634,N_17580);
or U17823 (N_17823,N_17613,N_17668);
and U17824 (N_17824,N_17520,N_17640);
and U17825 (N_17825,N_17576,N_17594);
nor U17826 (N_17826,N_17703,N_17518);
nor U17827 (N_17827,N_17681,N_17709);
nand U17828 (N_17828,N_17622,N_17725);
nand U17829 (N_17829,N_17660,N_17536);
or U17830 (N_17830,N_17691,N_17617);
nor U17831 (N_17831,N_17515,N_17693);
xnor U17832 (N_17832,N_17542,N_17603);
nor U17833 (N_17833,N_17504,N_17736);
xor U17834 (N_17834,N_17558,N_17625);
nand U17835 (N_17835,N_17547,N_17667);
and U17836 (N_17836,N_17514,N_17620);
nand U17837 (N_17837,N_17722,N_17539);
xor U17838 (N_17838,N_17567,N_17614);
and U17839 (N_17839,N_17538,N_17700);
or U17840 (N_17840,N_17650,N_17548);
or U17841 (N_17841,N_17611,N_17662);
and U17842 (N_17842,N_17551,N_17659);
or U17843 (N_17843,N_17682,N_17683);
or U17844 (N_17844,N_17720,N_17519);
or U17845 (N_17845,N_17562,N_17730);
and U17846 (N_17846,N_17544,N_17592);
and U17847 (N_17847,N_17628,N_17748);
xnor U17848 (N_17848,N_17666,N_17589);
nand U17849 (N_17849,N_17710,N_17605);
nand U17850 (N_17850,N_17632,N_17687);
nor U17851 (N_17851,N_17561,N_17534);
or U17852 (N_17852,N_17572,N_17523);
or U17853 (N_17853,N_17721,N_17513);
xnor U17854 (N_17854,N_17545,N_17711);
and U17855 (N_17855,N_17530,N_17646);
and U17856 (N_17856,N_17743,N_17638);
or U17857 (N_17857,N_17680,N_17645);
xnor U17858 (N_17858,N_17560,N_17718);
xnor U17859 (N_17859,N_17661,N_17578);
xor U17860 (N_17860,N_17563,N_17607);
and U17861 (N_17861,N_17702,N_17532);
and U17862 (N_17862,N_17679,N_17533);
nand U17863 (N_17863,N_17511,N_17745);
and U17864 (N_17864,N_17670,N_17696);
or U17865 (N_17865,N_17615,N_17595);
or U17866 (N_17866,N_17740,N_17508);
xnor U17867 (N_17867,N_17714,N_17507);
and U17868 (N_17868,N_17503,N_17568);
nand U17869 (N_17869,N_17629,N_17636);
nor U17870 (N_17870,N_17521,N_17747);
nand U17871 (N_17871,N_17510,N_17549);
xnor U17872 (N_17872,N_17688,N_17599);
or U17873 (N_17873,N_17697,N_17601);
nand U17874 (N_17874,N_17593,N_17744);
or U17875 (N_17875,N_17682,N_17634);
nor U17876 (N_17876,N_17624,N_17633);
or U17877 (N_17877,N_17639,N_17532);
nor U17878 (N_17878,N_17744,N_17606);
nor U17879 (N_17879,N_17587,N_17605);
nor U17880 (N_17880,N_17569,N_17680);
and U17881 (N_17881,N_17709,N_17733);
nor U17882 (N_17882,N_17642,N_17740);
nand U17883 (N_17883,N_17734,N_17666);
and U17884 (N_17884,N_17529,N_17518);
or U17885 (N_17885,N_17649,N_17573);
xnor U17886 (N_17886,N_17706,N_17500);
xnor U17887 (N_17887,N_17732,N_17707);
and U17888 (N_17888,N_17741,N_17566);
or U17889 (N_17889,N_17554,N_17565);
xnor U17890 (N_17890,N_17644,N_17557);
nor U17891 (N_17891,N_17690,N_17702);
nand U17892 (N_17892,N_17710,N_17533);
nor U17893 (N_17893,N_17572,N_17635);
nor U17894 (N_17894,N_17640,N_17745);
or U17895 (N_17895,N_17694,N_17602);
or U17896 (N_17896,N_17518,N_17571);
or U17897 (N_17897,N_17615,N_17670);
nand U17898 (N_17898,N_17668,N_17738);
or U17899 (N_17899,N_17622,N_17600);
and U17900 (N_17900,N_17704,N_17708);
nor U17901 (N_17901,N_17680,N_17737);
and U17902 (N_17902,N_17539,N_17617);
nor U17903 (N_17903,N_17747,N_17662);
nor U17904 (N_17904,N_17555,N_17561);
and U17905 (N_17905,N_17592,N_17559);
nor U17906 (N_17906,N_17501,N_17655);
nor U17907 (N_17907,N_17545,N_17594);
nand U17908 (N_17908,N_17552,N_17500);
and U17909 (N_17909,N_17563,N_17646);
and U17910 (N_17910,N_17673,N_17589);
nand U17911 (N_17911,N_17604,N_17563);
nand U17912 (N_17912,N_17639,N_17687);
or U17913 (N_17913,N_17723,N_17638);
nand U17914 (N_17914,N_17542,N_17746);
nand U17915 (N_17915,N_17662,N_17539);
or U17916 (N_17916,N_17611,N_17729);
and U17917 (N_17917,N_17502,N_17742);
or U17918 (N_17918,N_17618,N_17535);
and U17919 (N_17919,N_17632,N_17624);
and U17920 (N_17920,N_17724,N_17560);
and U17921 (N_17921,N_17680,N_17649);
and U17922 (N_17922,N_17637,N_17726);
and U17923 (N_17923,N_17733,N_17650);
and U17924 (N_17924,N_17508,N_17694);
xnor U17925 (N_17925,N_17694,N_17594);
xor U17926 (N_17926,N_17749,N_17617);
and U17927 (N_17927,N_17662,N_17535);
and U17928 (N_17928,N_17578,N_17575);
nand U17929 (N_17929,N_17639,N_17622);
nor U17930 (N_17930,N_17652,N_17623);
nor U17931 (N_17931,N_17543,N_17699);
or U17932 (N_17932,N_17552,N_17618);
or U17933 (N_17933,N_17540,N_17606);
nor U17934 (N_17934,N_17515,N_17615);
nor U17935 (N_17935,N_17520,N_17552);
xnor U17936 (N_17936,N_17677,N_17571);
and U17937 (N_17937,N_17590,N_17685);
and U17938 (N_17938,N_17509,N_17591);
nand U17939 (N_17939,N_17640,N_17541);
and U17940 (N_17940,N_17521,N_17729);
nand U17941 (N_17941,N_17686,N_17575);
nand U17942 (N_17942,N_17548,N_17579);
and U17943 (N_17943,N_17731,N_17530);
xnor U17944 (N_17944,N_17738,N_17664);
xnor U17945 (N_17945,N_17612,N_17604);
nand U17946 (N_17946,N_17661,N_17577);
and U17947 (N_17947,N_17673,N_17562);
and U17948 (N_17948,N_17665,N_17713);
nor U17949 (N_17949,N_17537,N_17541);
nor U17950 (N_17950,N_17674,N_17642);
or U17951 (N_17951,N_17677,N_17556);
or U17952 (N_17952,N_17574,N_17523);
xor U17953 (N_17953,N_17552,N_17728);
xnor U17954 (N_17954,N_17619,N_17622);
nand U17955 (N_17955,N_17534,N_17590);
and U17956 (N_17956,N_17560,N_17650);
nand U17957 (N_17957,N_17676,N_17653);
and U17958 (N_17958,N_17580,N_17529);
and U17959 (N_17959,N_17608,N_17537);
xor U17960 (N_17960,N_17539,N_17708);
nand U17961 (N_17961,N_17584,N_17629);
or U17962 (N_17962,N_17515,N_17623);
or U17963 (N_17963,N_17564,N_17630);
nand U17964 (N_17964,N_17551,N_17656);
nor U17965 (N_17965,N_17686,N_17701);
and U17966 (N_17966,N_17527,N_17506);
nand U17967 (N_17967,N_17547,N_17566);
or U17968 (N_17968,N_17526,N_17625);
nor U17969 (N_17969,N_17728,N_17634);
xor U17970 (N_17970,N_17547,N_17658);
xor U17971 (N_17971,N_17694,N_17521);
xnor U17972 (N_17972,N_17622,N_17515);
and U17973 (N_17973,N_17733,N_17734);
and U17974 (N_17974,N_17581,N_17599);
nor U17975 (N_17975,N_17522,N_17638);
and U17976 (N_17976,N_17590,N_17670);
or U17977 (N_17977,N_17681,N_17674);
xnor U17978 (N_17978,N_17531,N_17739);
or U17979 (N_17979,N_17744,N_17573);
or U17980 (N_17980,N_17566,N_17641);
or U17981 (N_17981,N_17653,N_17710);
nor U17982 (N_17982,N_17647,N_17610);
or U17983 (N_17983,N_17632,N_17583);
nor U17984 (N_17984,N_17632,N_17503);
nand U17985 (N_17985,N_17714,N_17743);
or U17986 (N_17986,N_17673,N_17704);
and U17987 (N_17987,N_17747,N_17579);
xnor U17988 (N_17988,N_17744,N_17506);
nand U17989 (N_17989,N_17593,N_17738);
xnor U17990 (N_17990,N_17696,N_17749);
or U17991 (N_17991,N_17638,N_17640);
nand U17992 (N_17992,N_17538,N_17684);
and U17993 (N_17993,N_17657,N_17608);
xor U17994 (N_17994,N_17733,N_17736);
nor U17995 (N_17995,N_17513,N_17595);
nand U17996 (N_17996,N_17660,N_17600);
nand U17997 (N_17997,N_17732,N_17672);
nor U17998 (N_17998,N_17735,N_17647);
nand U17999 (N_17999,N_17722,N_17586);
and U18000 (N_18000,N_17865,N_17912);
nor U18001 (N_18001,N_17875,N_17902);
nand U18002 (N_18002,N_17978,N_17815);
xnor U18003 (N_18003,N_17808,N_17974);
xnor U18004 (N_18004,N_17937,N_17946);
nor U18005 (N_18005,N_17931,N_17827);
or U18006 (N_18006,N_17909,N_17858);
xnor U18007 (N_18007,N_17955,N_17890);
or U18008 (N_18008,N_17926,N_17903);
and U18009 (N_18009,N_17973,N_17889);
nor U18010 (N_18010,N_17830,N_17940);
nor U18011 (N_18011,N_17873,N_17981);
or U18012 (N_18012,N_17755,N_17838);
and U18013 (N_18013,N_17753,N_17915);
xnor U18014 (N_18014,N_17866,N_17990);
or U18015 (N_18015,N_17862,N_17930);
or U18016 (N_18016,N_17919,N_17962);
nor U18017 (N_18017,N_17882,N_17952);
or U18018 (N_18018,N_17905,N_17906);
and U18019 (N_18019,N_17896,N_17789);
and U18020 (N_18020,N_17968,N_17798);
nor U18021 (N_18021,N_17831,N_17999);
nor U18022 (N_18022,N_17923,N_17871);
and U18023 (N_18023,N_17880,N_17975);
nand U18024 (N_18024,N_17939,N_17986);
xor U18025 (N_18025,N_17860,N_17996);
and U18026 (N_18026,N_17961,N_17886);
nand U18027 (N_18027,N_17960,N_17778);
and U18028 (N_18028,N_17754,N_17799);
or U18029 (N_18029,N_17944,N_17828);
xnor U18030 (N_18030,N_17760,N_17947);
xor U18031 (N_18031,N_17911,N_17966);
or U18032 (N_18032,N_17757,N_17956);
nand U18033 (N_18033,N_17872,N_17852);
nor U18034 (N_18034,N_17948,N_17985);
nand U18035 (N_18035,N_17984,N_17842);
nor U18036 (N_18036,N_17788,N_17997);
or U18037 (N_18037,N_17817,N_17797);
xnor U18038 (N_18038,N_17802,N_17795);
nor U18039 (N_18039,N_17979,N_17897);
nor U18040 (N_18040,N_17887,N_17811);
nor U18041 (N_18041,N_17777,N_17976);
and U18042 (N_18042,N_17806,N_17823);
nand U18043 (N_18043,N_17864,N_17989);
nand U18044 (N_18044,N_17980,N_17963);
or U18045 (N_18045,N_17837,N_17783);
xnor U18046 (N_18046,N_17950,N_17824);
nand U18047 (N_18047,N_17787,N_17868);
nand U18048 (N_18048,N_17921,N_17958);
xnor U18049 (N_18049,N_17899,N_17826);
or U18050 (N_18050,N_17987,N_17767);
xnor U18051 (N_18051,N_17907,N_17977);
nor U18052 (N_18052,N_17784,N_17917);
xnor U18053 (N_18053,N_17861,N_17764);
and U18054 (N_18054,N_17885,N_17949);
nand U18055 (N_18055,N_17800,N_17782);
and U18056 (N_18056,N_17771,N_17918);
and U18057 (N_18057,N_17769,N_17854);
nand U18058 (N_18058,N_17941,N_17957);
and U18059 (N_18059,N_17936,N_17879);
nor U18060 (N_18060,N_17943,N_17770);
nor U18061 (N_18061,N_17925,N_17779);
or U18062 (N_18062,N_17959,N_17874);
nand U18063 (N_18063,N_17821,N_17759);
or U18064 (N_18064,N_17801,N_17964);
and U18065 (N_18065,N_17859,N_17766);
or U18066 (N_18066,N_17792,N_17870);
nand U18067 (N_18067,N_17790,N_17867);
nand U18068 (N_18068,N_17869,N_17825);
nand U18069 (N_18069,N_17751,N_17983);
nor U18070 (N_18070,N_17796,N_17904);
nand U18071 (N_18071,N_17829,N_17791);
nor U18072 (N_18072,N_17851,N_17910);
or U18073 (N_18073,N_17992,N_17994);
or U18074 (N_18074,N_17850,N_17953);
or U18075 (N_18075,N_17818,N_17898);
nor U18076 (N_18076,N_17781,N_17835);
and U18077 (N_18077,N_17773,N_17793);
and U18078 (N_18078,N_17900,N_17846);
nand U18079 (N_18079,N_17935,N_17855);
xor U18080 (N_18080,N_17775,N_17933);
nand U18081 (N_18081,N_17991,N_17881);
and U18082 (N_18082,N_17929,N_17805);
nor U18083 (N_18083,N_17785,N_17847);
xnor U18084 (N_18084,N_17878,N_17932);
xnor U18085 (N_18085,N_17993,N_17942);
xnor U18086 (N_18086,N_17998,N_17807);
and U18087 (N_18087,N_17853,N_17863);
nand U18088 (N_18088,N_17970,N_17768);
or U18089 (N_18089,N_17967,N_17819);
nand U18090 (N_18090,N_17761,N_17914);
or U18091 (N_18091,N_17922,N_17988);
or U18092 (N_18092,N_17750,N_17794);
xor U18093 (N_18093,N_17776,N_17848);
nor U18094 (N_18094,N_17891,N_17833);
xnor U18095 (N_18095,N_17916,N_17908);
nor U18096 (N_18096,N_17844,N_17934);
xor U18097 (N_18097,N_17834,N_17756);
xnor U18098 (N_18098,N_17893,N_17845);
xnor U18099 (N_18099,N_17876,N_17892);
or U18100 (N_18100,N_17849,N_17995);
or U18101 (N_18101,N_17920,N_17816);
and U18102 (N_18102,N_17877,N_17803);
or U18103 (N_18103,N_17762,N_17839);
nand U18104 (N_18104,N_17945,N_17813);
nand U18105 (N_18105,N_17901,N_17812);
and U18106 (N_18106,N_17758,N_17786);
and U18107 (N_18107,N_17804,N_17951);
and U18108 (N_18108,N_17971,N_17780);
or U18109 (N_18109,N_17972,N_17969);
xnor U18110 (N_18110,N_17772,N_17822);
xnor U18111 (N_18111,N_17965,N_17888);
xnor U18112 (N_18112,N_17840,N_17895);
xnor U18113 (N_18113,N_17857,N_17774);
nor U18114 (N_18114,N_17982,N_17954);
nor U18115 (N_18115,N_17913,N_17832);
nor U18116 (N_18116,N_17820,N_17836);
xnor U18117 (N_18117,N_17927,N_17752);
and U18118 (N_18118,N_17928,N_17938);
nor U18119 (N_18119,N_17765,N_17884);
nand U18120 (N_18120,N_17763,N_17924);
nor U18121 (N_18121,N_17883,N_17894);
or U18122 (N_18122,N_17809,N_17843);
and U18123 (N_18123,N_17814,N_17841);
xor U18124 (N_18124,N_17856,N_17810);
nor U18125 (N_18125,N_17985,N_17863);
nor U18126 (N_18126,N_17908,N_17845);
and U18127 (N_18127,N_17822,N_17863);
nand U18128 (N_18128,N_17782,N_17966);
nand U18129 (N_18129,N_17822,N_17892);
nor U18130 (N_18130,N_17972,N_17929);
nor U18131 (N_18131,N_17933,N_17871);
nor U18132 (N_18132,N_17861,N_17830);
nand U18133 (N_18133,N_17840,N_17904);
or U18134 (N_18134,N_17975,N_17993);
xnor U18135 (N_18135,N_17824,N_17816);
and U18136 (N_18136,N_17771,N_17791);
and U18137 (N_18137,N_17867,N_17994);
xnor U18138 (N_18138,N_17825,N_17956);
and U18139 (N_18139,N_17961,N_17888);
or U18140 (N_18140,N_17899,N_17979);
nor U18141 (N_18141,N_17867,N_17975);
or U18142 (N_18142,N_17790,N_17966);
nor U18143 (N_18143,N_17893,N_17774);
xor U18144 (N_18144,N_17770,N_17786);
and U18145 (N_18145,N_17807,N_17994);
nand U18146 (N_18146,N_17888,N_17854);
and U18147 (N_18147,N_17762,N_17826);
xnor U18148 (N_18148,N_17965,N_17957);
xnor U18149 (N_18149,N_17768,N_17835);
nor U18150 (N_18150,N_17968,N_17761);
xnor U18151 (N_18151,N_17971,N_17968);
and U18152 (N_18152,N_17764,N_17795);
nand U18153 (N_18153,N_17847,N_17910);
or U18154 (N_18154,N_17942,N_17755);
or U18155 (N_18155,N_17761,N_17926);
nand U18156 (N_18156,N_17785,N_17997);
and U18157 (N_18157,N_17976,N_17804);
and U18158 (N_18158,N_17924,N_17931);
xor U18159 (N_18159,N_17981,N_17774);
or U18160 (N_18160,N_17828,N_17757);
nand U18161 (N_18161,N_17838,N_17861);
or U18162 (N_18162,N_17765,N_17931);
nor U18163 (N_18163,N_17911,N_17902);
nor U18164 (N_18164,N_17867,N_17992);
or U18165 (N_18165,N_17991,N_17843);
and U18166 (N_18166,N_17755,N_17790);
xnor U18167 (N_18167,N_17983,N_17864);
or U18168 (N_18168,N_17976,N_17904);
xor U18169 (N_18169,N_17875,N_17913);
or U18170 (N_18170,N_17857,N_17790);
and U18171 (N_18171,N_17795,N_17889);
nor U18172 (N_18172,N_17910,N_17978);
and U18173 (N_18173,N_17901,N_17847);
xnor U18174 (N_18174,N_17893,N_17833);
or U18175 (N_18175,N_17771,N_17817);
nor U18176 (N_18176,N_17947,N_17950);
nand U18177 (N_18177,N_17948,N_17991);
nand U18178 (N_18178,N_17758,N_17827);
and U18179 (N_18179,N_17755,N_17944);
nand U18180 (N_18180,N_17949,N_17791);
or U18181 (N_18181,N_17767,N_17864);
and U18182 (N_18182,N_17809,N_17803);
xnor U18183 (N_18183,N_17871,N_17932);
or U18184 (N_18184,N_17761,N_17999);
nand U18185 (N_18185,N_17987,N_17911);
and U18186 (N_18186,N_17874,N_17957);
nand U18187 (N_18187,N_17821,N_17804);
nor U18188 (N_18188,N_17944,N_17942);
nand U18189 (N_18189,N_17884,N_17874);
nand U18190 (N_18190,N_17952,N_17988);
or U18191 (N_18191,N_17921,N_17915);
and U18192 (N_18192,N_17911,N_17937);
nand U18193 (N_18193,N_17793,N_17974);
or U18194 (N_18194,N_17875,N_17860);
or U18195 (N_18195,N_17862,N_17981);
and U18196 (N_18196,N_17960,N_17988);
and U18197 (N_18197,N_17794,N_17939);
xor U18198 (N_18198,N_17870,N_17888);
xor U18199 (N_18199,N_17972,N_17998);
or U18200 (N_18200,N_17996,N_17914);
nor U18201 (N_18201,N_17945,N_17844);
or U18202 (N_18202,N_17833,N_17944);
nor U18203 (N_18203,N_17870,N_17883);
and U18204 (N_18204,N_17778,N_17827);
and U18205 (N_18205,N_17781,N_17905);
and U18206 (N_18206,N_17888,N_17949);
nand U18207 (N_18207,N_17970,N_17946);
or U18208 (N_18208,N_17849,N_17796);
xnor U18209 (N_18209,N_17927,N_17994);
nand U18210 (N_18210,N_17955,N_17821);
or U18211 (N_18211,N_17856,N_17948);
nor U18212 (N_18212,N_17979,N_17785);
nand U18213 (N_18213,N_17948,N_17886);
nand U18214 (N_18214,N_17826,N_17975);
and U18215 (N_18215,N_17757,N_17838);
or U18216 (N_18216,N_17945,N_17926);
or U18217 (N_18217,N_17986,N_17875);
nor U18218 (N_18218,N_17762,N_17972);
xnor U18219 (N_18219,N_17891,N_17813);
nor U18220 (N_18220,N_17847,N_17923);
nand U18221 (N_18221,N_17914,N_17910);
nor U18222 (N_18222,N_17822,N_17988);
or U18223 (N_18223,N_17952,N_17783);
nor U18224 (N_18224,N_17883,N_17785);
nor U18225 (N_18225,N_17760,N_17754);
nand U18226 (N_18226,N_17777,N_17980);
xnor U18227 (N_18227,N_17771,N_17782);
nor U18228 (N_18228,N_17856,N_17956);
and U18229 (N_18229,N_17780,N_17894);
nor U18230 (N_18230,N_17875,N_17823);
or U18231 (N_18231,N_17825,N_17969);
nor U18232 (N_18232,N_17903,N_17880);
xor U18233 (N_18233,N_17935,N_17772);
nand U18234 (N_18234,N_17836,N_17763);
or U18235 (N_18235,N_17790,N_17763);
or U18236 (N_18236,N_17960,N_17772);
nor U18237 (N_18237,N_17862,N_17768);
or U18238 (N_18238,N_17790,N_17885);
nand U18239 (N_18239,N_17835,N_17900);
xnor U18240 (N_18240,N_17779,N_17870);
nor U18241 (N_18241,N_17967,N_17918);
xnor U18242 (N_18242,N_17832,N_17876);
or U18243 (N_18243,N_17957,N_17906);
xnor U18244 (N_18244,N_17855,N_17834);
and U18245 (N_18245,N_17794,N_17759);
or U18246 (N_18246,N_17801,N_17969);
or U18247 (N_18247,N_17854,N_17809);
nor U18248 (N_18248,N_17968,N_17854);
nor U18249 (N_18249,N_17875,N_17905);
or U18250 (N_18250,N_18079,N_18248);
xnor U18251 (N_18251,N_18019,N_18140);
nand U18252 (N_18252,N_18071,N_18203);
and U18253 (N_18253,N_18062,N_18229);
xor U18254 (N_18254,N_18080,N_18135);
and U18255 (N_18255,N_18070,N_18075);
xor U18256 (N_18256,N_18205,N_18189);
nand U18257 (N_18257,N_18120,N_18178);
xnor U18258 (N_18258,N_18083,N_18162);
or U18259 (N_18259,N_18066,N_18169);
and U18260 (N_18260,N_18064,N_18133);
nand U18261 (N_18261,N_18008,N_18001);
nor U18262 (N_18262,N_18016,N_18240);
nand U18263 (N_18263,N_18085,N_18040);
or U18264 (N_18264,N_18047,N_18235);
and U18265 (N_18265,N_18111,N_18036);
and U18266 (N_18266,N_18226,N_18005);
and U18267 (N_18267,N_18215,N_18179);
and U18268 (N_18268,N_18065,N_18225);
or U18269 (N_18269,N_18220,N_18007);
and U18270 (N_18270,N_18216,N_18144);
nor U18271 (N_18271,N_18217,N_18227);
nor U18272 (N_18272,N_18043,N_18116);
nand U18273 (N_18273,N_18073,N_18190);
and U18274 (N_18274,N_18056,N_18078);
xor U18275 (N_18275,N_18011,N_18029);
nor U18276 (N_18276,N_18223,N_18018);
or U18277 (N_18277,N_18048,N_18241);
or U18278 (N_18278,N_18104,N_18233);
nand U18279 (N_18279,N_18055,N_18126);
or U18280 (N_18280,N_18035,N_18053);
nand U18281 (N_18281,N_18031,N_18157);
nor U18282 (N_18282,N_18000,N_18068);
and U18283 (N_18283,N_18171,N_18151);
nand U18284 (N_18284,N_18197,N_18173);
xnor U18285 (N_18285,N_18122,N_18050);
nand U18286 (N_18286,N_18054,N_18091);
nor U18287 (N_18287,N_18132,N_18209);
and U18288 (N_18288,N_18231,N_18167);
xor U18289 (N_18289,N_18159,N_18182);
nand U18290 (N_18290,N_18181,N_18097);
nor U18291 (N_18291,N_18187,N_18138);
nor U18292 (N_18292,N_18081,N_18023);
and U18293 (N_18293,N_18185,N_18152);
and U18294 (N_18294,N_18130,N_18088);
and U18295 (N_18295,N_18098,N_18245);
nor U18296 (N_18296,N_18172,N_18165);
nor U18297 (N_18297,N_18101,N_18117);
nand U18298 (N_18298,N_18030,N_18009);
or U18299 (N_18299,N_18163,N_18049);
xnor U18300 (N_18300,N_18058,N_18148);
or U18301 (N_18301,N_18090,N_18156);
nand U18302 (N_18302,N_18025,N_18014);
or U18303 (N_18303,N_18114,N_18191);
nand U18304 (N_18304,N_18067,N_18057);
xnor U18305 (N_18305,N_18200,N_18086);
xnor U18306 (N_18306,N_18180,N_18125);
xnor U18307 (N_18307,N_18143,N_18022);
and U18308 (N_18308,N_18017,N_18045);
nor U18309 (N_18309,N_18107,N_18202);
nand U18310 (N_18310,N_18141,N_18192);
or U18311 (N_18311,N_18224,N_18119);
xnor U18312 (N_18312,N_18027,N_18087);
xor U18313 (N_18313,N_18063,N_18129);
nor U18314 (N_18314,N_18033,N_18010);
or U18315 (N_18315,N_18006,N_18020);
nand U18316 (N_18316,N_18213,N_18204);
nor U18317 (N_18317,N_18124,N_18096);
and U18318 (N_18318,N_18243,N_18034);
xnor U18319 (N_18319,N_18059,N_18232);
xor U18320 (N_18320,N_18028,N_18242);
nor U18321 (N_18321,N_18222,N_18176);
nand U18322 (N_18322,N_18201,N_18150);
xor U18323 (N_18323,N_18089,N_18100);
and U18324 (N_18324,N_18155,N_18195);
nor U18325 (N_18325,N_18121,N_18032);
nand U18326 (N_18326,N_18039,N_18003);
or U18327 (N_18327,N_18188,N_18012);
nor U18328 (N_18328,N_18210,N_18024);
or U18329 (N_18329,N_18136,N_18153);
or U18330 (N_18330,N_18103,N_18002);
and U18331 (N_18331,N_18236,N_18084);
xnor U18332 (N_18332,N_18109,N_18099);
or U18333 (N_18333,N_18228,N_18060);
nand U18334 (N_18334,N_18094,N_18221);
or U18335 (N_18335,N_18131,N_18112);
nor U18336 (N_18336,N_18113,N_18093);
nand U18337 (N_18337,N_18106,N_18037);
nand U18338 (N_18338,N_18021,N_18015);
and U18339 (N_18339,N_18149,N_18147);
or U18340 (N_18340,N_18077,N_18118);
nor U18341 (N_18341,N_18168,N_18184);
xnor U18342 (N_18342,N_18183,N_18108);
nand U18343 (N_18343,N_18146,N_18142);
nor U18344 (N_18344,N_18249,N_18158);
and U18345 (N_18345,N_18069,N_18160);
and U18346 (N_18346,N_18198,N_18186);
xnor U18347 (N_18347,N_18042,N_18237);
or U18348 (N_18348,N_18175,N_18244);
nor U18349 (N_18349,N_18145,N_18230);
xnor U18350 (N_18350,N_18208,N_18041);
and U18351 (N_18351,N_18102,N_18074);
or U18352 (N_18352,N_18234,N_18214);
nand U18353 (N_18353,N_18004,N_18164);
or U18354 (N_18354,N_18026,N_18154);
nor U18355 (N_18355,N_18134,N_18218);
nand U18356 (N_18356,N_18219,N_18211);
nor U18357 (N_18357,N_18128,N_18239);
or U18358 (N_18358,N_18092,N_18194);
and U18359 (N_18359,N_18199,N_18105);
and U18360 (N_18360,N_18046,N_18061);
and U18361 (N_18361,N_18137,N_18095);
or U18362 (N_18362,N_18013,N_18207);
or U18363 (N_18363,N_18174,N_18206);
nor U18364 (N_18364,N_18082,N_18044);
nand U18365 (N_18365,N_18052,N_18038);
and U18366 (N_18366,N_18115,N_18161);
xor U18367 (N_18367,N_18076,N_18212);
nor U18368 (N_18368,N_18193,N_18170);
and U18369 (N_18369,N_18139,N_18247);
nand U18370 (N_18370,N_18123,N_18110);
xnor U18371 (N_18371,N_18246,N_18177);
nand U18372 (N_18372,N_18166,N_18127);
xnor U18373 (N_18373,N_18072,N_18051);
and U18374 (N_18374,N_18196,N_18238);
or U18375 (N_18375,N_18225,N_18043);
and U18376 (N_18376,N_18025,N_18224);
xnor U18377 (N_18377,N_18016,N_18069);
xor U18378 (N_18378,N_18028,N_18077);
or U18379 (N_18379,N_18209,N_18174);
and U18380 (N_18380,N_18135,N_18163);
or U18381 (N_18381,N_18105,N_18218);
nand U18382 (N_18382,N_18167,N_18034);
nand U18383 (N_18383,N_18015,N_18076);
and U18384 (N_18384,N_18085,N_18165);
nor U18385 (N_18385,N_18190,N_18121);
or U18386 (N_18386,N_18154,N_18011);
xor U18387 (N_18387,N_18029,N_18240);
nor U18388 (N_18388,N_18079,N_18117);
and U18389 (N_18389,N_18126,N_18000);
nand U18390 (N_18390,N_18165,N_18186);
xor U18391 (N_18391,N_18158,N_18228);
or U18392 (N_18392,N_18044,N_18069);
nor U18393 (N_18393,N_18042,N_18169);
and U18394 (N_18394,N_18240,N_18083);
nor U18395 (N_18395,N_18075,N_18193);
nand U18396 (N_18396,N_18177,N_18244);
and U18397 (N_18397,N_18169,N_18109);
and U18398 (N_18398,N_18158,N_18244);
nand U18399 (N_18399,N_18122,N_18231);
nor U18400 (N_18400,N_18234,N_18213);
nor U18401 (N_18401,N_18045,N_18176);
xor U18402 (N_18402,N_18153,N_18126);
nand U18403 (N_18403,N_18081,N_18209);
and U18404 (N_18404,N_18124,N_18201);
and U18405 (N_18405,N_18095,N_18077);
or U18406 (N_18406,N_18047,N_18247);
xor U18407 (N_18407,N_18004,N_18088);
or U18408 (N_18408,N_18065,N_18142);
nor U18409 (N_18409,N_18080,N_18195);
or U18410 (N_18410,N_18215,N_18109);
or U18411 (N_18411,N_18045,N_18066);
nor U18412 (N_18412,N_18168,N_18096);
or U18413 (N_18413,N_18169,N_18050);
and U18414 (N_18414,N_18182,N_18175);
xnor U18415 (N_18415,N_18007,N_18214);
and U18416 (N_18416,N_18168,N_18143);
and U18417 (N_18417,N_18140,N_18102);
and U18418 (N_18418,N_18180,N_18147);
xor U18419 (N_18419,N_18023,N_18094);
nand U18420 (N_18420,N_18018,N_18014);
nor U18421 (N_18421,N_18071,N_18003);
xor U18422 (N_18422,N_18021,N_18217);
and U18423 (N_18423,N_18203,N_18176);
and U18424 (N_18424,N_18184,N_18042);
nor U18425 (N_18425,N_18034,N_18053);
and U18426 (N_18426,N_18247,N_18022);
nor U18427 (N_18427,N_18217,N_18148);
nand U18428 (N_18428,N_18233,N_18022);
nor U18429 (N_18429,N_18022,N_18204);
nor U18430 (N_18430,N_18029,N_18093);
or U18431 (N_18431,N_18067,N_18227);
xor U18432 (N_18432,N_18031,N_18015);
or U18433 (N_18433,N_18196,N_18067);
nand U18434 (N_18434,N_18211,N_18065);
xor U18435 (N_18435,N_18189,N_18235);
and U18436 (N_18436,N_18243,N_18108);
and U18437 (N_18437,N_18007,N_18129);
or U18438 (N_18438,N_18097,N_18017);
and U18439 (N_18439,N_18242,N_18008);
xnor U18440 (N_18440,N_18086,N_18091);
xnor U18441 (N_18441,N_18173,N_18108);
nand U18442 (N_18442,N_18015,N_18024);
nor U18443 (N_18443,N_18001,N_18239);
or U18444 (N_18444,N_18067,N_18173);
nand U18445 (N_18445,N_18104,N_18163);
or U18446 (N_18446,N_18209,N_18166);
xnor U18447 (N_18447,N_18112,N_18211);
xnor U18448 (N_18448,N_18052,N_18122);
or U18449 (N_18449,N_18066,N_18051);
and U18450 (N_18450,N_18161,N_18246);
xor U18451 (N_18451,N_18214,N_18053);
and U18452 (N_18452,N_18093,N_18104);
or U18453 (N_18453,N_18234,N_18175);
nor U18454 (N_18454,N_18039,N_18207);
nand U18455 (N_18455,N_18172,N_18205);
or U18456 (N_18456,N_18015,N_18018);
nor U18457 (N_18457,N_18247,N_18049);
and U18458 (N_18458,N_18056,N_18191);
and U18459 (N_18459,N_18243,N_18143);
nor U18460 (N_18460,N_18227,N_18216);
and U18461 (N_18461,N_18006,N_18064);
and U18462 (N_18462,N_18093,N_18127);
nor U18463 (N_18463,N_18200,N_18195);
and U18464 (N_18464,N_18126,N_18176);
xor U18465 (N_18465,N_18114,N_18099);
xor U18466 (N_18466,N_18082,N_18114);
nand U18467 (N_18467,N_18210,N_18034);
xor U18468 (N_18468,N_18146,N_18016);
or U18469 (N_18469,N_18221,N_18149);
nand U18470 (N_18470,N_18141,N_18077);
or U18471 (N_18471,N_18103,N_18077);
xor U18472 (N_18472,N_18045,N_18076);
and U18473 (N_18473,N_18166,N_18032);
and U18474 (N_18474,N_18247,N_18118);
or U18475 (N_18475,N_18094,N_18211);
nand U18476 (N_18476,N_18182,N_18214);
xnor U18477 (N_18477,N_18081,N_18093);
nor U18478 (N_18478,N_18127,N_18176);
and U18479 (N_18479,N_18042,N_18079);
and U18480 (N_18480,N_18107,N_18236);
and U18481 (N_18481,N_18189,N_18214);
xnor U18482 (N_18482,N_18004,N_18234);
nand U18483 (N_18483,N_18150,N_18244);
xnor U18484 (N_18484,N_18099,N_18170);
xor U18485 (N_18485,N_18025,N_18090);
nand U18486 (N_18486,N_18065,N_18194);
xnor U18487 (N_18487,N_18103,N_18215);
nand U18488 (N_18488,N_18196,N_18007);
xnor U18489 (N_18489,N_18219,N_18198);
xnor U18490 (N_18490,N_18027,N_18052);
nor U18491 (N_18491,N_18211,N_18212);
and U18492 (N_18492,N_18197,N_18179);
xnor U18493 (N_18493,N_18239,N_18092);
nand U18494 (N_18494,N_18183,N_18118);
nor U18495 (N_18495,N_18183,N_18032);
nor U18496 (N_18496,N_18028,N_18036);
xor U18497 (N_18497,N_18119,N_18184);
xnor U18498 (N_18498,N_18213,N_18001);
or U18499 (N_18499,N_18029,N_18088);
nor U18500 (N_18500,N_18463,N_18316);
xnor U18501 (N_18501,N_18390,N_18284);
xnor U18502 (N_18502,N_18365,N_18472);
or U18503 (N_18503,N_18445,N_18326);
nand U18504 (N_18504,N_18392,N_18306);
and U18505 (N_18505,N_18469,N_18256);
and U18506 (N_18506,N_18263,N_18251);
nand U18507 (N_18507,N_18484,N_18279);
nor U18508 (N_18508,N_18489,N_18427);
nor U18509 (N_18509,N_18456,N_18267);
nand U18510 (N_18510,N_18368,N_18361);
nand U18511 (N_18511,N_18328,N_18317);
xnor U18512 (N_18512,N_18477,N_18337);
nor U18513 (N_18513,N_18367,N_18331);
nor U18514 (N_18514,N_18380,N_18264);
xor U18515 (N_18515,N_18372,N_18414);
and U18516 (N_18516,N_18266,N_18345);
or U18517 (N_18517,N_18354,N_18253);
nand U18518 (N_18518,N_18371,N_18418);
and U18519 (N_18519,N_18373,N_18307);
nor U18520 (N_18520,N_18313,N_18495);
or U18521 (N_18521,N_18433,N_18282);
xor U18522 (N_18522,N_18320,N_18357);
and U18523 (N_18523,N_18290,N_18301);
nor U18524 (N_18524,N_18274,N_18471);
and U18525 (N_18525,N_18482,N_18434);
and U18526 (N_18526,N_18397,N_18454);
nor U18527 (N_18527,N_18388,N_18483);
xor U18528 (N_18528,N_18449,N_18258);
and U18529 (N_18529,N_18499,N_18423);
and U18530 (N_18530,N_18448,N_18461);
or U18531 (N_18531,N_18323,N_18330);
nand U18532 (N_18532,N_18378,N_18322);
nand U18533 (N_18533,N_18492,N_18466);
and U18534 (N_18534,N_18362,N_18413);
or U18535 (N_18535,N_18281,N_18441);
nand U18536 (N_18536,N_18338,N_18339);
xor U18537 (N_18537,N_18415,N_18481);
xnor U18538 (N_18538,N_18341,N_18305);
and U18539 (N_18539,N_18476,N_18364);
or U18540 (N_18540,N_18447,N_18269);
or U18541 (N_18541,N_18470,N_18496);
xor U18542 (N_18542,N_18416,N_18324);
or U18543 (N_18543,N_18400,N_18366);
nor U18544 (N_18544,N_18292,N_18375);
and U18545 (N_18545,N_18298,N_18343);
and U18546 (N_18546,N_18485,N_18465);
nor U18547 (N_18547,N_18428,N_18321);
or U18548 (N_18548,N_18363,N_18382);
nor U18549 (N_18549,N_18488,N_18370);
and U18550 (N_18550,N_18406,N_18325);
xor U18551 (N_18551,N_18435,N_18391);
and U18552 (N_18552,N_18404,N_18405);
nand U18553 (N_18553,N_18389,N_18295);
xnor U18554 (N_18554,N_18276,N_18296);
nor U18555 (N_18555,N_18334,N_18257);
and U18556 (N_18556,N_18387,N_18459);
nor U18557 (N_18557,N_18261,N_18411);
xnor U18558 (N_18558,N_18310,N_18420);
and U18559 (N_18559,N_18285,N_18349);
and U18560 (N_18560,N_18344,N_18271);
xor U18561 (N_18561,N_18260,N_18342);
xor U18562 (N_18562,N_18304,N_18480);
nand U18563 (N_18563,N_18272,N_18430);
nand U18564 (N_18564,N_18302,N_18335);
or U18565 (N_18565,N_18451,N_18450);
xor U18566 (N_18566,N_18444,N_18315);
and U18567 (N_18567,N_18308,N_18312);
and U18568 (N_18568,N_18436,N_18452);
xnor U18569 (N_18569,N_18475,N_18395);
nor U18570 (N_18570,N_18309,N_18487);
nor U18571 (N_18571,N_18401,N_18376);
or U18572 (N_18572,N_18283,N_18280);
nor U18573 (N_18573,N_18297,N_18259);
and U18574 (N_18574,N_18396,N_18336);
nand U18575 (N_18575,N_18358,N_18473);
xor U18576 (N_18576,N_18369,N_18318);
or U18577 (N_18577,N_18303,N_18410);
xnor U18578 (N_18578,N_18408,N_18252);
nor U18579 (N_18579,N_18464,N_18467);
nor U18580 (N_18580,N_18491,N_18359);
nor U18581 (N_18581,N_18431,N_18494);
xor U18582 (N_18582,N_18409,N_18446);
and U18583 (N_18583,N_18497,N_18356);
and U18584 (N_18584,N_18439,N_18270);
nand U18585 (N_18585,N_18393,N_18314);
and U18586 (N_18586,N_18262,N_18377);
or U18587 (N_18587,N_18474,N_18398);
or U18588 (N_18588,N_18479,N_18384);
nand U18589 (N_18589,N_18468,N_18417);
or U18590 (N_18590,N_18462,N_18486);
xnor U18591 (N_18591,N_18268,N_18351);
or U18592 (N_18592,N_18287,N_18333);
and U18593 (N_18593,N_18327,N_18402);
nand U18594 (N_18594,N_18300,N_18374);
and U18595 (N_18595,N_18275,N_18407);
xnor U18596 (N_18596,N_18437,N_18291);
nor U18597 (N_18597,N_18379,N_18293);
nand U18598 (N_18598,N_18425,N_18255);
nand U18599 (N_18599,N_18286,N_18498);
nand U18600 (N_18600,N_18383,N_18348);
or U18601 (N_18601,N_18455,N_18289);
nand U18602 (N_18602,N_18443,N_18319);
and U18603 (N_18603,N_18453,N_18440);
nor U18604 (N_18604,N_18332,N_18347);
nand U18605 (N_18605,N_18350,N_18273);
xor U18606 (N_18606,N_18386,N_18294);
nor U18607 (N_18607,N_18458,N_18311);
and U18608 (N_18608,N_18299,N_18254);
nand U18609 (N_18609,N_18250,N_18360);
nand U18610 (N_18610,N_18381,N_18394);
or U18611 (N_18611,N_18288,N_18277);
xnor U18612 (N_18612,N_18385,N_18442);
and U18613 (N_18613,N_18490,N_18424);
nand U18614 (N_18614,N_18412,N_18399);
nor U18615 (N_18615,N_18478,N_18493);
and U18616 (N_18616,N_18346,N_18340);
and U18617 (N_18617,N_18278,N_18438);
and U18618 (N_18618,N_18265,N_18460);
nor U18619 (N_18619,N_18329,N_18421);
nand U18620 (N_18620,N_18352,N_18457);
nor U18621 (N_18621,N_18419,N_18403);
and U18622 (N_18622,N_18432,N_18429);
and U18623 (N_18623,N_18353,N_18426);
nor U18624 (N_18624,N_18422,N_18355);
or U18625 (N_18625,N_18354,N_18387);
xnor U18626 (N_18626,N_18380,N_18438);
nor U18627 (N_18627,N_18466,N_18282);
or U18628 (N_18628,N_18395,N_18449);
or U18629 (N_18629,N_18298,N_18316);
or U18630 (N_18630,N_18258,N_18414);
nor U18631 (N_18631,N_18476,N_18314);
and U18632 (N_18632,N_18462,N_18252);
nor U18633 (N_18633,N_18360,N_18478);
nand U18634 (N_18634,N_18318,N_18440);
nand U18635 (N_18635,N_18299,N_18257);
or U18636 (N_18636,N_18355,N_18476);
nand U18637 (N_18637,N_18414,N_18279);
nor U18638 (N_18638,N_18282,N_18327);
or U18639 (N_18639,N_18459,N_18281);
nand U18640 (N_18640,N_18314,N_18329);
nand U18641 (N_18641,N_18371,N_18314);
or U18642 (N_18642,N_18389,N_18262);
or U18643 (N_18643,N_18442,N_18471);
and U18644 (N_18644,N_18405,N_18427);
nand U18645 (N_18645,N_18480,N_18462);
nand U18646 (N_18646,N_18443,N_18467);
nand U18647 (N_18647,N_18374,N_18492);
nor U18648 (N_18648,N_18350,N_18349);
nor U18649 (N_18649,N_18259,N_18462);
xnor U18650 (N_18650,N_18391,N_18413);
xnor U18651 (N_18651,N_18253,N_18481);
xor U18652 (N_18652,N_18251,N_18382);
or U18653 (N_18653,N_18330,N_18440);
nand U18654 (N_18654,N_18433,N_18348);
or U18655 (N_18655,N_18433,N_18369);
or U18656 (N_18656,N_18424,N_18448);
or U18657 (N_18657,N_18472,N_18317);
and U18658 (N_18658,N_18467,N_18474);
nor U18659 (N_18659,N_18356,N_18299);
nand U18660 (N_18660,N_18496,N_18297);
nor U18661 (N_18661,N_18332,N_18360);
or U18662 (N_18662,N_18488,N_18409);
nor U18663 (N_18663,N_18296,N_18465);
xor U18664 (N_18664,N_18420,N_18488);
nor U18665 (N_18665,N_18334,N_18318);
nand U18666 (N_18666,N_18315,N_18420);
xor U18667 (N_18667,N_18274,N_18260);
nor U18668 (N_18668,N_18379,N_18435);
or U18669 (N_18669,N_18454,N_18469);
and U18670 (N_18670,N_18440,N_18425);
and U18671 (N_18671,N_18442,N_18288);
nor U18672 (N_18672,N_18389,N_18453);
nor U18673 (N_18673,N_18363,N_18431);
xor U18674 (N_18674,N_18400,N_18455);
xor U18675 (N_18675,N_18412,N_18353);
nand U18676 (N_18676,N_18336,N_18469);
or U18677 (N_18677,N_18405,N_18345);
nand U18678 (N_18678,N_18425,N_18337);
nor U18679 (N_18679,N_18372,N_18255);
or U18680 (N_18680,N_18428,N_18477);
nand U18681 (N_18681,N_18305,N_18363);
nor U18682 (N_18682,N_18338,N_18459);
xor U18683 (N_18683,N_18318,N_18298);
or U18684 (N_18684,N_18347,N_18391);
nor U18685 (N_18685,N_18427,N_18384);
or U18686 (N_18686,N_18305,N_18330);
nor U18687 (N_18687,N_18262,N_18406);
nor U18688 (N_18688,N_18269,N_18259);
nor U18689 (N_18689,N_18418,N_18355);
xnor U18690 (N_18690,N_18444,N_18461);
or U18691 (N_18691,N_18487,N_18250);
xor U18692 (N_18692,N_18354,N_18322);
and U18693 (N_18693,N_18391,N_18406);
nand U18694 (N_18694,N_18330,N_18326);
nor U18695 (N_18695,N_18296,N_18441);
xnor U18696 (N_18696,N_18476,N_18467);
xor U18697 (N_18697,N_18420,N_18400);
xnor U18698 (N_18698,N_18404,N_18333);
xor U18699 (N_18699,N_18303,N_18382);
or U18700 (N_18700,N_18380,N_18439);
nor U18701 (N_18701,N_18498,N_18277);
nor U18702 (N_18702,N_18485,N_18486);
xor U18703 (N_18703,N_18291,N_18433);
or U18704 (N_18704,N_18412,N_18286);
nor U18705 (N_18705,N_18451,N_18330);
or U18706 (N_18706,N_18416,N_18274);
xnor U18707 (N_18707,N_18328,N_18267);
nand U18708 (N_18708,N_18294,N_18348);
and U18709 (N_18709,N_18491,N_18258);
or U18710 (N_18710,N_18337,N_18308);
or U18711 (N_18711,N_18305,N_18251);
xnor U18712 (N_18712,N_18368,N_18311);
nor U18713 (N_18713,N_18336,N_18274);
nor U18714 (N_18714,N_18473,N_18378);
and U18715 (N_18715,N_18372,N_18469);
nand U18716 (N_18716,N_18478,N_18463);
nor U18717 (N_18717,N_18428,N_18376);
xor U18718 (N_18718,N_18288,N_18392);
and U18719 (N_18719,N_18312,N_18416);
or U18720 (N_18720,N_18398,N_18412);
or U18721 (N_18721,N_18281,N_18296);
nor U18722 (N_18722,N_18327,N_18281);
nor U18723 (N_18723,N_18268,N_18464);
or U18724 (N_18724,N_18257,N_18461);
and U18725 (N_18725,N_18424,N_18261);
and U18726 (N_18726,N_18413,N_18409);
nand U18727 (N_18727,N_18458,N_18472);
and U18728 (N_18728,N_18331,N_18471);
and U18729 (N_18729,N_18336,N_18363);
or U18730 (N_18730,N_18442,N_18499);
nand U18731 (N_18731,N_18458,N_18262);
nor U18732 (N_18732,N_18252,N_18323);
nand U18733 (N_18733,N_18277,N_18365);
and U18734 (N_18734,N_18451,N_18424);
and U18735 (N_18735,N_18388,N_18436);
nor U18736 (N_18736,N_18312,N_18293);
and U18737 (N_18737,N_18444,N_18455);
or U18738 (N_18738,N_18356,N_18370);
nand U18739 (N_18739,N_18252,N_18404);
nand U18740 (N_18740,N_18484,N_18359);
or U18741 (N_18741,N_18446,N_18443);
and U18742 (N_18742,N_18470,N_18269);
or U18743 (N_18743,N_18250,N_18474);
and U18744 (N_18744,N_18287,N_18439);
nand U18745 (N_18745,N_18442,N_18347);
nor U18746 (N_18746,N_18433,N_18469);
nand U18747 (N_18747,N_18272,N_18277);
or U18748 (N_18748,N_18264,N_18402);
nor U18749 (N_18749,N_18391,N_18323);
or U18750 (N_18750,N_18534,N_18667);
and U18751 (N_18751,N_18543,N_18612);
and U18752 (N_18752,N_18683,N_18620);
xor U18753 (N_18753,N_18560,N_18561);
nor U18754 (N_18754,N_18663,N_18725);
xnor U18755 (N_18755,N_18589,N_18528);
nand U18756 (N_18756,N_18711,N_18598);
nor U18757 (N_18757,N_18721,N_18697);
nand U18758 (N_18758,N_18614,N_18510);
and U18759 (N_18759,N_18553,N_18689);
or U18760 (N_18760,N_18719,N_18684);
or U18761 (N_18761,N_18690,N_18655);
and U18762 (N_18762,N_18502,N_18659);
xnor U18763 (N_18763,N_18657,N_18708);
nand U18764 (N_18764,N_18602,N_18610);
and U18765 (N_18765,N_18675,N_18664);
or U18766 (N_18766,N_18595,N_18578);
nand U18767 (N_18767,N_18660,N_18638);
and U18768 (N_18768,N_18681,N_18674);
nor U18769 (N_18769,N_18677,N_18642);
xor U18770 (N_18770,N_18525,N_18724);
or U18771 (N_18771,N_18590,N_18627);
nor U18772 (N_18772,N_18737,N_18630);
or U18773 (N_18773,N_18665,N_18713);
or U18774 (N_18774,N_18706,N_18701);
or U18775 (N_18775,N_18747,N_18732);
xor U18776 (N_18776,N_18524,N_18718);
nand U18777 (N_18777,N_18513,N_18714);
or U18778 (N_18778,N_18530,N_18507);
nor U18779 (N_18779,N_18717,N_18547);
nor U18780 (N_18780,N_18596,N_18519);
or U18781 (N_18781,N_18539,N_18694);
xnor U18782 (N_18782,N_18628,N_18639);
and U18783 (N_18783,N_18573,N_18535);
nand U18784 (N_18784,N_18552,N_18555);
xnor U18785 (N_18785,N_18640,N_18618);
or U18786 (N_18786,N_18575,N_18570);
xnor U18787 (N_18787,N_18647,N_18695);
or U18788 (N_18788,N_18532,N_18567);
or U18789 (N_18789,N_18529,N_18563);
xnor U18790 (N_18790,N_18641,N_18671);
xnor U18791 (N_18791,N_18545,N_18658);
or U18792 (N_18792,N_18691,N_18745);
nor U18793 (N_18793,N_18699,N_18669);
nor U18794 (N_18794,N_18738,N_18569);
nor U18795 (N_18795,N_18554,N_18599);
or U18796 (N_18796,N_18735,N_18716);
nand U18797 (N_18797,N_18582,N_18733);
or U18798 (N_18798,N_18601,N_18623);
and U18799 (N_18799,N_18604,N_18704);
or U18800 (N_18800,N_18741,N_18608);
and U18801 (N_18801,N_18603,N_18703);
or U18802 (N_18802,N_18593,N_18597);
and U18803 (N_18803,N_18637,N_18654);
nand U18804 (N_18804,N_18693,N_18729);
nand U18805 (N_18805,N_18526,N_18730);
nand U18806 (N_18806,N_18621,N_18523);
xnor U18807 (N_18807,N_18722,N_18509);
nor U18808 (N_18808,N_18583,N_18636);
or U18809 (N_18809,N_18615,N_18576);
nor U18810 (N_18810,N_18744,N_18562);
and U18811 (N_18811,N_18698,N_18505);
nor U18812 (N_18812,N_18629,N_18606);
and U18813 (N_18813,N_18586,N_18666);
and U18814 (N_18814,N_18653,N_18517);
and U18815 (N_18815,N_18670,N_18611);
nand U18816 (N_18816,N_18592,N_18688);
nand U18817 (N_18817,N_18679,N_18692);
nand U18818 (N_18818,N_18538,N_18672);
xor U18819 (N_18819,N_18515,N_18580);
nor U18820 (N_18820,N_18607,N_18727);
xnor U18821 (N_18821,N_18650,N_18726);
nor U18822 (N_18822,N_18619,N_18577);
and U18823 (N_18823,N_18546,N_18673);
or U18824 (N_18824,N_18522,N_18533);
or U18825 (N_18825,N_18696,N_18587);
xnor U18826 (N_18826,N_18503,N_18504);
nor U18827 (N_18827,N_18742,N_18668);
or U18828 (N_18828,N_18616,N_18702);
nand U18829 (N_18829,N_18712,N_18536);
and U18830 (N_18830,N_18501,N_18687);
xnor U18831 (N_18831,N_18736,N_18631);
xor U18832 (N_18832,N_18540,N_18743);
nand U18833 (N_18833,N_18521,N_18643);
nor U18834 (N_18834,N_18626,N_18574);
and U18835 (N_18835,N_18656,N_18746);
or U18836 (N_18836,N_18739,N_18565);
and U18837 (N_18837,N_18506,N_18720);
and U18838 (N_18838,N_18500,N_18705);
nand U18839 (N_18839,N_18748,N_18548);
or U18840 (N_18840,N_18564,N_18572);
nor U18841 (N_18841,N_18613,N_18609);
nand U18842 (N_18842,N_18676,N_18511);
xor U18843 (N_18843,N_18516,N_18644);
or U18844 (N_18844,N_18625,N_18520);
nand U18845 (N_18845,N_18556,N_18633);
xnor U18846 (N_18846,N_18514,N_18678);
or U18847 (N_18847,N_18709,N_18531);
nand U18848 (N_18848,N_18584,N_18594);
nor U18849 (N_18849,N_18549,N_18728);
nand U18850 (N_18850,N_18537,N_18700);
or U18851 (N_18851,N_18600,N_18617);
nor U18852 (N_18852,N_18686,N_18685);
nor U18853 (N_18853,N_18662,N_18648);
xor U18854 (N_18854,N_18558,N_18634);
nand U18855 (N_18855,N_18518,N_18680);
xnor U18856 (N_18856,N_18508,N_18591);
and U18857 (N_18857,N_18624,N_18571);
nand U18858 (N_18858,N_18710,N_18661);
or U18859 (N_18859,N_18588,N_18632);
nand U18860 (N_18860,N_18581,N_18566);
nor U18861 (N_18861,N_18622,N_18646);
and U18862 (N_18862,N_18734,N_18740);
nand U18863 (N_18863,N_18749,N_18568);
xnor U18864 (N_18864,N_18551,N_18635);
nand U18865 (N_18865,N_18707,N_18649);
nor U18866 (N_18866,N_18715,N_18585);
nand U18867 (N_18867,N_18682,N_18559);
xor U18868 (N_18868,N_18542,N_18645);
xor U18869 (N_18869,N_18723,N_18731);
nor U18870 (N_18870,N_18550,N_18527);
xnor U18871 (N_18871,N_18579,N_18544);
or U18872 (N_18872,N_18512,N_18652);
or U18873 (N_18873,N_18651,N_18541);
nand U18874 (N_18874,N_18605,N_18557);
or U18875 (N_18875,N_18540,N_18732);
and U18876 (N_18876,N_18678,N_18500);
or U18877 (N_18877,N_18740,N_18729);
and U18878 (N_18878,N_18524,N_18633);
or U18879 (N_18879,N_18557,N_18524);
xnor U18880 (N_18880,N_18622,N_18738);
or U18881 (N_18881,N_18743,N_18652);
nand U18882 (N_18882,N_18620,N_18637);
nand U18883 (N_18883,N_18723,N_18719);
nand U18884 (N_18884,N_18637,N_18630);
xnor U18885 (N_18885,N_18746,N_18643);
and U18886 (N_18886,N_18599,N_18711);
and U18887 (N_18887,N_18624,N_18703);
nor U18888 (N_18888,N_18590,N_18574);
or U18889 (N_18889,N_18678,N_18695);
nor U18890 (N_18890,N_18614,N_18625);
or U18891 (N_18891,N_18523,N_18532);
nor U18892 (N_18892,N_18558,N_18658);
and U18893 (N_18893,N_18637,N_18641);
xnor U18894 (N_18894,N_18620,N_18625);
or U18895 (N_18895,N_18510,N_18656);
or U18896 (N_18896,N_18674,N_18502);
nand U18897 (N_18897,N_18680,N_18612);
nor U18898 (N_18898,N_18622,N_18541);
and U18899 (N_18899,N_18580,N_18506);
or U18900 (N_18900,N_18595,N_18646);
xor U18901 (N_18901,N_18585,N_18548);
nand U18902 (N_18902,N_18635,N_18592);
xnor U18903 (N_18903,N_18588,N_18710);
xor U18904 (N_18904,N_18535,N_18615);
and U18905 (N_18905,N_18724,N_18634);
and U18906 (N_18906,N_18524,N_18669);
nand U18907 (N_18907,N_18624,N_18573);
xor U18908 (N_18908,N_18664,N_18740);
or U18909 (N_18909,N_18569,N_18686);
nor U18910 (N_18910,N_18501,N_18673);
nand U18911 (N_18911,N_18501,N_18644);
xor U18912 (N_18912,N_18689,N_18716);
xor U18913 (N_18913,N_18634,N_18611);
or U18914 (N_18914,N_18664,N_18579);
or U18915 (N_18915,N_18707,N_18524);
nand U18916 (N_18916,N_18539,N_18521);
or U18917 (N_18917,N_18580,N_18582);
and U18918 (N_18918,N_18611,N_18703);
nor U18919 (N_18919,N_18630,N_18586);
and U18920 (N_18920,N_18645,N_18603);
and U18921 (N_18921,N_18715,N_18725);
xnor U18922 (N_18922,N_18581,N_18605);
xnor U18923 (N_18923,N_18567,N_18665);
or U18924 (N_18924,N_18650,N_18662);
or U18925 (N_18925,N_18746,N_18589);
or U18926 (N_18926,N_18510,N_18581);
nand U18927 (N_18927,N_18535,N_18501);
xnor U18928 (N_18928,N_18601,N_18671);
or U18929 (N_18929,N_18588,N_18677);
and U18930 (N_18930,N_18730,N_18706);
and U18931 (N_18931,N_18631,N_18726);
or U18932 (N_18932,N_18586,N_18683);
and U18933 (N_18933,N_18504,N_18695);
xor U18934 (N_18934,N_18603,N_18558);
or U18935 (N_18935,N_18635,N_18618);
nand U18936 (N_18936,N_18583,N_18534);
xnor U18937 (N_18937,N_18606,N_18501);
and U18938 (N_18938,N_18685,N_18715);
nand U18939 (N_18939,N_18593,N_18724);
or U18940 (N_18940,N_18581,N_18678);
xor U18941 (N_18941,N_18649,N_18601);
nand U18942 (N_18942,N_18532,N_18749);
or U18943 (N_18943,N_18725,N_18528);
nand U18944 (N_18944,N_18719,N_18657);
and U18945 (N_18945,N_18656,N_18584);
nor U18946 (N_18946,N_18747,N_18696);
nand U18947 (N_18947,N_18673,N_18653);
nand U18948 (N_18948,N_18634,N_18683);
or U18949 (N_18949,N_18521,N_18686);
or U18950 (N_18950,N_18628,N_18591);
nor U18951 (N_18951,N_18695,N_18627);
nand U18952 (N_18952,N_18645,N_18631);
nor U18953 (N_18953,N_18584,N_18522);
or U18954 (N_18954,N_18551,N_18511);
nor U18955 (N_18955,N_18583,N_18527);
xor U18956 (N_18956,N_18707,N_18532);
xor U18957 (N_18957,N_18702,N_18663);
nand U18958 (N_18958,N_18737,N_18696);
or U18959 (N_18959,N_18530,N_18510);
nor U18960 (N_18960,N_18556,N_18739);
nor U18961 (N_18961,N_18632,N_18546);
nand U18962 (N_18962,N_18707,N_18589);
and U18963 (N_18963,N_18501,N_18604);
or U18964 (N_18964,N_18530,N_18709);
and U18965 (N_18965,N_18602,N_18644);
nand U18966 (N_18966,N_18594,N_18664);
nand U18967 (N_18967,N_18622,N_18736);
or U18968 (N_18968,N_18572,N_18580);
nand U18969 (N_18969,N_18653,N_18609);
nor U18970 (N_18970,N_18522,N_18543);
nor U18971 (N_18971,N_18687,N_18588);
or U18972 (N_18972,N_18702,N_18555);
and U18973 (N_18973,N_18724,N_18738);
or U18974 (N_18974,N_18542,N_18531);
xnor U18975 (N_18975,N_18532,N_18608);
nor U18976 (N_18976,N_18564,N_18503);
and U18977 (N_18977,N_18636,N_18521);
nand U18978 (N_18978,N_18615,N_18575);
nor U18979 (N_18979,N_18546,N_18601);
and U18980 (N_18980,N_18579,N_18504);
nor U18981 (N_18981,N_18606,N_18698);
nand U18982 (N_18982,N_18731,N_18642);
or U18983 (N_18983,N_18744,N_18587);
and U18984 (N_18984,N_18702,N_18642);
nor U18985 (N_18985,N_18728,N_18703);
and U18986 (N_18986,N_18686,N_18505);
or U18987 (N_18987,N_18634,N_18676);
xor U18988 (N_18988,N_18725,N_18692);
or U18989 (N_18989,N_18613,N_18629);
or U18990 (N_18990,N_18603,N_18564);
xnor U18991 (N_18991,N_18697,N_18739);
xnor U18992 (N_18992,N_18618,N_18601);
nor U18993 (N_18993,N_18504,N_18578);
or U18994 (N_18994,N_18642,N_18664);
nand U18995 (N_18995,N_18748,N_18725);
xnor U18996 (N_18996,N_18581,N_18742);
nor U18997 (N_18997,N_18657,N_18539);
nand U18998 (N_18998,N_18696,N_18711);
xor U18999 (N_18999,N_18553,N_18731);
nand U19000 (N_19000,N_18889,N_18831);
or U19001 (N_19001,N_18936,N_18909);
xor U19002 (N_19002,N_18856,N_18928);
nand U19003 (N_19003,N_18819,N_18849);
xnor U19004 (N_19004,N_18785,N_18790);
and U19005 (N_19005,N_18798,N_18767);
and U19006 (N_19006,N_18920,N_18836);
or U19007 (N_19007,N_18941,N_18838);
and U19008 (N_19008,N_18752,N_18977);
nand U19009 (N_19009,N_18773,N_18815);
nand U19010 (N_19010,N_18753,N_18884);
xor U19011 (N_19011,N_18963,N_18924);
xnor U19012 (N_19012,N_18929,N_18812);
xor U19013 (N_19013,N_18948,N_18876);
or U19014 (N_19014,N_18987,N_18829);
or U19015 (N_19015,N_18843,N_18821);
and U19016 (N_19016,N_18771,N_18908);
nand U19017 (N_19017,N_18768,N_18994);
nand U19018 (N_19018,N_18933,N_18806);
or U19019 (N_19019,N_18860,N_18765);
or U19020 (N_19020,N_18766,N_18844);
nor U19021 (N_19021,N_18841,N_18868);
or U19022 (N_19022,N_18960,N_18961);
nor U19023 (N_19023,N_18997,N_18760);
and U19024 (N_19024,N_18795,N_18754);
or U19025 (N_19025,N_18839,N_18947);
xnor U19026 (N_19026,N_18855,N_18750);
or U19027 (N_19027,N_18922,N_18899);
or U19028 (N_19028,N_18930,N_18890);
and U19029 (N_19029,N_18925,N_18923);
nor U19030 (N_19030,N_18916,N_18939);
and U19031 (N_19031,N_18793,N_18866);
nand U19032 (N_19032,N_18902,N_18896);
or U19033 (N_19033,N_18881,N_18917);
nand U19034 (N_19034,N_18776,N_18951);
and U19035 (N_19035,N_18833,N_18974);
xor U19036 (N_19036,N_18976,N_18932);
or U19037 (N_19037,N_18955,N_18956);
xnor U19038 (N_19038,N_18807,N_18891);
and U19039 (N_19039,N_18906,N_18938);
nor U19040 (N_19040,N_18864,N_18822);
or U19041 (N_19041,N_18847,N_18911);
or U19042 (N_19042,N_18910,N_18887);
nor U19043 (N_19043,N_18971,N_18969);
xor U19044 (N_19044,N_18931,N_18893);
nor U19045 (N_19045,N_18903,N_18772);
nor U19046 (N_19046,N_18787,N_18885);
and U19047 (N_19047,N_18981,N_18796);
xnor U19048 (N_19048,N_18888,N_18992);
or U19049 (N_19049,N_18804,N_18830);
nor U19050 (N_19050,N_18937,N_18781);
nor U19051 (N_19051,N_18805,N_18845);
or U19052 (N_19052,N_18770,N_18898);
nor U19053 (N_19053,N_18859,N_18826);
nand U19054 (N_19054,N_18802,N_18914);
nor U19055 (N_19055,N_18813,N_18820);
nor U19056 (N_19056,N_18799,N_18817);
or U19057 (N_19057,N_18962,N_18842);
and U19058 (N_19058,N_18763,N_18789);
nor U19059 (N_19059,N_18777,N_18854);
and U19060 (N_19060,N_18825,N_18999);
and U19061 (N_19061,N_18980,N_18861);
or U19062 (N_19062,N_18788,N_18949);
or U19063 (N_19063,N_18835,N_18823);
and U19064 (N_19064,N_18904,N_18975);
xor U19065 (N_19065,N_18983,N_18940);
nand U19066 (N_19066,N_18935,N_18791);
or U19067 (N_19067,N_18837,N_18784);
or U19068 (N_19068,N_18800,N_18945);
nor U19069 (N_19069,N_18900,N_18792);
and U19070 (N_19070,N_18946,N_18883);
nand U19071 (N_19071,N_18882,N_18897);
or U19072 (N_19072,N_18991,N_18848);
nand U19073 (N_19073,N_18985,N_18756);
or U19074 (N_19074,N_18959,N_18867);
nand U19075 (N_19075,N_18840,N_18886);
nand U19076 (N_19076,N_18775,N_18921);
and U19077 (N_19077,N_18942,N_18982);
or U19078 (N_19078,N_18895,N_18973);
nand U19079 (N_19079,N_18782,N_18912);
and U19080 (N_19080,N_18824,N_18783);
nor U19081 (N_19081,N_18852,N_18757);
nor U19082 (N_19082,N_18944,N_18873);
or U19083 (N_19083,N_18846,N_18778);
nand U19084 (N_19084,N_18797,N_18953);
or U19085 (N_19085,N_18943,N_18986);
or U19086 (N_19086,N_18979,N_18927);
nor U19087 (N_19087,N_18964,N_18869);
xor U19088 (N_19088,N_18863,N_18877);
nand U19089 (N_19089,N_18993,N_18915);
and U19090 (N_19090,N_18857,N_18834);
xnor U19091 (N_19091,N_18918,N_18816);
and U19092 (N_19092,N_18965,N_18871);
or U19093 (N_19093,N_18769,N_18984);
nand U19094 (N_19094,N_18762,N_18878);
xnor U19095 (N_19095,N_18901,N_18803);
nand U19096 (N_19096,N_18850,N_18759);
and U19097 (N_19097,N_18811,N_18958);
nand U19098 (N_19098,N_18801,N_18818);
nor U19099 (N_19099,N_18874,N_18755);
or U19100 (N_19100,N_18970,N_18894);
and U19101 (N_19101,N_18919,N_18978);
xor U19102 (N_19102,N_18814,N_18954);
or U19103 (N_19103,N_18774,N_18967);
nor U19104 (N_19104,N_18832,N_18966);
and U19105 (N_19105,N_18988,N_18758);
xor U19106 (N_19106,N_18905,N_18957);
nand U19107 (N_19107,N_18968,N_18879);
nand U19108 (N_19108,N_18865,N_18952);
nor U19109 (N_19109,N_18828,N_18998);
nand U19110 (N_19110,N_18972,N_18751);
and U19111 (N_19111,N_18794,N_18858);
and U19112 (N_19112,N_18872,N_18934);
nand U19113 (N_19113,N_18875,N_18827);
xor U19114 (N_19114,N_18764,N_18989);
xnor U19115 (N_19115,N_18851,N_18995);
nor U19116 (N_19116,N_18862,N_18907);
xnor U19117 (N_19117,N_18809,N_18810);
or U19118 (N_19118,N_18996,N_18808);
xor U19119 (N_19119,N_18779,N_18990);
or U19120 (N_19120,N_18950,N_18913);
nor U19121 (N_19121,N_18892,N_18761);
and U19122 (N_19122,N_18780,N_18786);
xor U19123 (N_19123,N_18880,N_18853);
nor U19124 (N_19124,N_18926,N_18870);
or U19125 (N_19125,N_18810,N_18871);
nor U19126 (N_19126,N_18928,N_18858);
or U19127 (N_19127,N_18929,N_18803);
nand U19128 (N_19128,N_18996,N_18777);
xnor U19129 (N_19129,N_18858,N_18884);
nand U19130 (N_19130,N_18947,N_18943);
nor U19131 (N_19131,N_18973,N_18775);
or U19132 (N_19132,N_18854,N_18847);
nand U19133 (N_19133,N_18903,N_18892);
nor U19134 (N_19134,N_18816,N_18771);
xnor U19135 (N_19135,N_18788,N_18996);
nor U19136 (N_19136,N_18784,N_18763);
nand U19137 (N_19137,N_18924,N_18881);
nor U19138 (N_19138,N_18836,N_18772);
or U19139 (N_19139,N_18782,N_18891);
or U19140 (N_19140,N_18890,N_18856);
or U19141 (N_19141,N_18847,N_18893);
xor U19142 (N_19142,N_18976,N_18949);
or U19143 (N_19143,N_18939,N_18899);
or U19144 (N_19144,N_18951,N_18965);
and U19145 (N_19145,N_18914,N_18843);
or U19146 (N_19146,N_18864,N_18820);
or U19147 (N_19147,N_18781,N_18811);
and U19148 (N_19148,N_18848,N_18841);
nor U19149 (N_19149,N_18862,N_18920);
or U19150 (N_19150,N_18957,N_18965);
nand U19151 (N_19151,N_18884,N_18783);
nand U19152 (N_19152,N_18947,N_18872);
nor U19153 (N_19153,N_18924,N_18807);
or U19154 (N_19154,N_18888,N_18901);
and U19155 (N_19155,N_18845,N_18910);
and U19156 (N_19156,N_18826,N_18895);
xor U19157 (N_19157,N_18848,N_18830);
xor U19158 (N_19158,N_18810,N_18837);
nor U19159 (N_19159,N_18850,N_18873);
nand U19160 (N_19160,N_18790,N_18961);
or U19161 (N_19161,N_18923,N_18772);
nand U19162 (N_19162,N_18816,N_18762);
nor U19163 (N_19163,N_18797,N_18841);
or U19164 (N_19164,N_18860,N_18874);
nand U19165 (N_19165,N_18857,N_18803);
nor U19166 (N_19166,N_18950,N_18917);
nand U19167 (N_19167,N_18919,N_18966);
nor U19168 (N_19168,N_18845,N_18946);
or U19169 (N_19169,N_18955,N_18945);
nor U19170 (N_19170,N_18852,N_18990);
xor U19171 (N_19171,N_18837,N_18972);
nor U19172 (N_19172,N_18778,N_18781);
nand U19173 (N_19173,N_18955,N_18878);
nor U19174 (N_19174,N_18790,N_18751);
or U19175 (N_19175,N_18989,N_18950);
nor U19176 (N_19176,N_18897,N_18862);
xnor U19177 (N_19177,N_18971,N_18935);
and U19178 (N_19178,N_18817,N_18888);
and U19179 (N_19179,N_18903,N_18857);
and U19180 (N_19180,N_18966,N_18945);
xor U19181 (N_19181,N_18861,N_18898);
nand U19182 (N_19182,N_18812,N_18754);
or U19183 (N_19183,N_18924,N_18849);
or U19184 (N_19184,N_18919,N_18928);
or U19185 (N_19185,N_18857,N_18814);
nor U19186 (N_19186,N_18885,N_18927);
and U19187 (N_19187,N_18950,N_18850);
nor U19188 (N_19188,N_18860,N_18959);
nor U19189 (N_19189,N_18819,N_18850);
nand U19190 (N_19190,N_18869,N_18886);
and U19191 (N_19191,N_18797,N_18965);
and U19192 (N_19192,N_18971,N_18898);
or U19193 (N_19193,N_18848,N_18896);
or U19194 (N_19194,N_18989,N_18850);
or U19195 (N_19195,N_18764,N_18901);
and U19196 (N_19196,N_18851,N_18868);
nand U19197 (N_19197,N_18757,N_18810);
nor U19198 (N_19198,N_18755,N_18779);
or U19199 (N_19199,N_18948,N_18960);
nand U19200 (N_19200,N_18891,N_18944);
or U19201 (N_19201,N_18886,N_18972);
nand U19202 (N_19202,N_18761,N_18876);
nor U19203 (N_19203,N_18753,N_18860);
nor U19204 (N_19204,N_18969,N_18798);
nand U19205 (N_19205,N_18990,N_18947);
nor U19206 (N_19206,N_18894,N_18991);
nand U19207 (N_19207,N_18995,N_18788);
xor U19208 (N_19208,N_18822,N_18989);
and U19209 (N_19209,N_18842,N_18753);
or U19210 (N_19210,N_18831,N_18914);
xnor U19211 (N_19211,N_18958,N_18796);
or U19212 (N_19212,N_18829,N_18836);
nand U19213 (N_19213,N_18843,N_18891);
or U19214 (N_19214,N_18956,N_18994);
nor U19215 (N_19215,N_18867,N_18875);
or U19216 (N_19216,N_18913,N_18921);
xnor U19217 (N_19217,N_18995,N_18920);
and U19218 (N_19218,N_18997,N_18796);
nor U19219 (N_19219,N_18928,N_18812);
and U19220 (N_19220,N_18858,N_18839);
xnor U19221 (N_19221,N_18938,N_18904);
nor U19222 (N_19222,N_18903,N_18828);
nand U19223 (N_19223,N_18996,N_18759);
or U19224 (N_19224,N_18978,N_18960);
or U19225 (N_19225,N_18921,N_18776);
xor U19226 (N_19226,N_18990,N_18876);
and U19227 (N_19227,N_18815,N_18921);
nor U19228 (N_19228,N_18788,N_18895);
nor U19229 (N_19229,N_18789,N_18875);
nor U19230 (N_19230,N_18850,N_18992);
and U19231 (N_19231,N_18914,N_18984);
xnor U19232 (N_19232,N_18940,N_18797);
nand U19233 (N_19233,N_18831,N_18868);
or U19234 (N_19234,N_18769,N_18817);
and U19235 (N_19235,N_18797,N_18941);
nand U19236 (N_19236,N_18884,N_18982);
and U19237 (N_19237,N_18787,N_18960);
xor U19238 (N_19238,N_18932,N_18781);
or U19239 (N_19239,N_18835,N_18878);
xor U19240 (N_19240,N_18931,N_18796);
nor U19241 (N_19241,N_18958,N_18867);
or U19242 (N_19242,N_18935,N_18984);
nor U19243 (N_19243,N_18867,N_18882);
nand U19244 (N_19244,N_18986,N_18769);
and U19245 (N_19245,N_18802,N_18841);
xor U19246 (N_19246,N_18814,N_18829);
nor U19247 (N_19247,N_18750,N_18998);
nand U19248 (N_19248,N_18798,N_18806);
and U19249 (N_19249,N_18906,N_18957);
and U19250 (N_19250,N_19127,N_19101);
xor U19251 (N_19251,N_19172,N_19075);
nand U19252 (N_19252,N_19020,N_19063);
nand U19253 (N_19253,N_19102,N_19081);
nor U19254 (N_19254,N_19079,N_19057);
and U19255 (N_19255,N_19227,N_19000);
nand U19256 (N_19256,N_19105,N_19166);
nand U19257 (N_19257,N_19206,N_19033);
nor U19258 (N_19258,N_19013,N_19224);
xor U19259 (N_19259,N_19204,N_19078);
or U19260 (N_19260,N_19168,N_19125);
xnor U19261 (N_19261,N_19199,N_19221);
or U19262 (N_19262,N_19178,N_19095);
xnor U19263 (N_19263,N_19119,N_19195);
or U19264 (N_19264,N_19086,N_19115);
and U19265 (N_19265,N_19175,N_19155);
and U19266 (N_19266,N_19183,N_19232);
and U19267 (N_19267,N_19117,N_19180);
xor U19268 (N_19268,N_19024,N_19233);
and U19269 (N_19269,N_19014,N_19005);
nand U19270 (N_19270,N_19062,N_19039);
nand U19271 (N_19271,N_19211,N_19110);
and U19272 (N_19272,N_19058,N_19149);
and U19273 (N_19273,N_19208,N_19114);
and U19274 (N_19274,N_19082,N_19192);
nand U19275 (N_19275,N_19070,N_19049);
xnor U19276 (N_19276,N_19093,N_19009);
and U19277 (N_19277,N_19006,N_19237);
or U19278 (N_19278,N_19076,N_19100);
or U19279 (N_19279,N_19123,N_19245);
xnor U19280 (N_19280,N_19174,N_19116);
nor U19281 (N_19281,N_19129,N_19152);
and U19282 (N_19282,N_19011,N_19069);
nand U19283 (N_19283,N_19176,N_19041);
nand U19284 (N_19284,N_19021,N_19084);
nand U19285 (N_19285,N_19177,N_19092);
or U19286 (N_19286,N_19001,N_19113);
nand U19287 (N_19287,N_19226,N_19243);
nor U19288 (N_19288,N_19036,N_19064);
xnor U19289 (N_19289,N_19098,N_19004);
or U19290 (N_19290,N_19225,N_19162);
or U19291 (N_19291,N_19094,N_19161);
or U19292 (N_19292,N_19173,N_19007);
or U19293 (N_19293,N_19133,N_19193);
nor U19294 (N_19294,N_19040,N_19203);
xor U19295 (N_19295,N_19061,N_19043);
xnor U19296 (N_19296,N_19128,N_19052);
nor U19297 (N_19297,N_19022,N_19207);
nand U19298 (N_19298,N_19025,N_19170);
and U19299 (N_19299,N_19141,N_19130);
nand U19300 (N_19300,N_19091,N_19201);
and U19301 (N_19301,N_19042,N_19028);
xnor U19302 (N_19302,N_19249,N_19003);
nand U19303 (N_19303,N_19072,N_19107);
nor U19304 (N_19304,N_19159,N_19090);
xnor U19305 (N_19305,N_19160,N_19214);
or U19306 (N_19306,N_19065,N_19147);
nor U19307 (N_19307,N_19066,N_19059);
nand U19308 (N_19308,N_19248,N_19118);
nor U19309 (N_19309,N_19104,N_19231);
or U19310 (N_19310,N_19038,N_19029);
nand U19311 (N_19311,N_19111,N_19015);
or U19312 (N_19312,N_19053,N_19145);
nor U19313 (N_19313,N_19055,N_19169);
nand U19314 (N_19314,N_19239,N_19150);
and U19315 (N_19315,N_19219,N_19136);
xnor U19316 (N_19316,N_19035,N_19045);
nand U19317 (N_19317,N_19151,N_19156);
and U19318 (N_19318,N_19074,N_19050);
nand U19319 (N_19319,N_19154,N_19012);
or U19320 (N_19320,N_19190,N_19167);
xor U19321 (N_19321,N_19108,N_19124);
nand U19322 (N_19322,N_19140,N_19077);
nand U19323 (N_19323,N_19034,N_19181);
nor U19324 (N_19324,N_19089,N_19158);
nor U19325 (N_19325,N_19085,N_19244);
or U19326 (N_19326,N_19080,N_19056);
xnor U19327 (N_19327,N_19213,N_19120);
xor U19328 (N_19328,N_19008,N_19048);
nor U19329 (N_19329,N_19131,N_19126);
nor U19330 (N_19330,N_19157,N_19026);
xnor U19331 (N_19331,N_19060,N_19247);
or U19332 (N_19332,N_19209,N_19184);
nand U19333 (N_19333,N_19179,N_19017);
or U19334 (N_19334,N_19210,N_19044);
and U19335 (N_19335,N_19241,N_19212);
or U19336 (N_19336,N_19139,N_19153);
nand U19337 (N_19337,N_19122,N_19073);
or U19338 (N_19338,N_19242,N_19216);
nand U19339 (N_19339,N_19197,N_19222);
xor U19340 (N_19340,N_19238,N_19023);
and U19341 (N_19341,N_19234,N_19121);
nor U19342 (N_19342,N_19240,N_19016);
xor U19343 (N_19343,N_19019,N_19137);
nor U19344 (N_19344,N_19202,N_19164);
and U19345 (N_19345,N_19112,N_19246);
nand U19346 (N_19346,N_19205,N_19217);
xnor U19347 (N_19347,N_19099,N_19071);
or U19348 (N_19348,N_19106,N_19163);
or U19349 (N_19349,N_19138,N_19196);
and U19350 (N_19350,N_19218,N_19109);
nor U19351 (N_19351,N_19146,N_19188);
xor U19352 (N_19352,N_19191,N_19067);
xor U19353 (N_19353,N_19046,N_19165);
nand U19354 (N_19354,N_19031,N_19047);
nand U19355 (N_19355,N_19200,N_19171);
or U19356 (N_19356,N_19032,N_19186);
nor U19357 (N_19357,N_19215,N_19051);
nor U19358 (N_19358,N_19148,N_19142);
and U19359 (N_19359,N_19182,N_19027);
nand U19360 (N_19360,N_19198,N_19054);
and U19361 (N_19361,N_19144,N_19220);
and U19362 (N_19362,N_19223,N_19010);
xnor U19363 (N_19363,N_19088,N_19235);
or U19364 (N_19364,N_19103,N_19002);
xor U19365 (N_19365,N_19097,N_19228);
xor U19366 (N_19366,N_19236,N_19030);
and U19367 (N_19367,N_19037,N_19143);
or U19368 (N_19368,N_19187,N_19068);
nand U19369 (N_19369,N_19185,N_19135);
nand U19370 (N_19370,N_19189,N_19230);
and U19371 (N_19371,N_19096,N_19083);
xor U19372 (N_19372,N_19134,N_19132);
or U19373 (N_19373,N_19229,N_19087);
nand U19374 (N_19374,N_19018,N_19194);
nor U19375 (N_19375,N_19228,N_19207);
xor U19376 (N_19376,N_19225,N_19070);
and U19377 (N_19377,N_19004,N_19010);
and U19378 (N_19378,N_19036,N_19245);
and U19379 (N_19379,N_19112,N_19185);
or U19380 (N_19380,N_19153,N_19202);
or U19381 (N_19381,N_19227,N_19001);
or U19382 (N_19382,N_19050,N_19109);
or U19383 (N_19383,N_19235,N_19193);
and U19384 (N_19384,N_19102,N_19139);
xnor U19385 (N_19385,N_19111,N_19105);
or U19386 (N_19386,N_19166,N_19200);
nor U19387 (N_19387,N_19083,N_19216);
or U19388 (N_19388,N_19069,N_19148);
nor U19389 (N_19389,N_19149,N_19043);
or U19390 (N_19390,N_19159,N_19152);
or U19391 (N_19391,N_19047,N_19058);
and U19392 (N_19392,N_19240,N_19160);
xor U19393 (N_19393,N_19178,N_19121);
nand U19394 (N_19394,N_19203,N_19033);
nand U19395 (N_19395,N_19053,N_19197);
xor U19396 (N_19396,N_19092,N_19157);
or U19397 (N_19397,N_19235,N_19205);
and U19398 (N_19398,N_19112,N_19029);
or U19399 (N_19399,N_19226,N_19040);
nand U19400 (N_19400,N_19100,N_19223);
xnor U19401 (N_19401,N_19128,N_19249);
xor U19402 (N_19402,N_19145,N_19074);
nor U19403 (N_19403,N_19160,N_19104);
or U19404 (N_19404,N_19240,N_19065);
and U19405 (N_19405,N_19068,N_19022);
and U19406 (N_19406,N_19168,N_19178);
nor U19407 (N_19407,N_19078,N_19213);
nand U19408 (N_19408,N_19219,N_19137);
nand U19409 (N_19409,N_19165,N_19064);
or U19410 (N_19410,N_19244,N_19078);
xor U19411 (N_19411,N_19104,N_19177);
nand U19412 (N_19412,N_19055,N_19098);
nor U19413 (N_19413,N_19192,N_19202);
xor U19414 (N_19414,N_19248,N_19080);
nor U19415 (N_19415,N_19195,N_19142);
xnor U19416 (N_19416,N_19087,N_19246);
nand U19417 (N_19417,N_19107,N_19080);
and U19418 (N_19418,N_19033,N_19167);
xnor U19419 (N_19419,N_19116,N_19232);
or U19420 (N_19420,N_19170,N_19117);
nand U19421 (N_19421,N_19014,N_19082);
and U19422 (N_19422,N_19079,N_19163);
nand U19423 (N_19423,N_19201,N_19167);
nor U19424 (N_19424,N_19008,N_19196);
nand U19425 (N_19425,N_19093,N_19019);
nand U19426 (N_19426,N_19079,N_19204);
or U19427 (N_19427,N_19062,N_19163);
nand U19428 (N_19428,N_19017,N_19235);
or U19429 (N_19429,N_19215,N_19068);
nor U19430 (N_19430,N_19090,N_19116);
and U19431 (N_19431,N_19078,N_19191);
and U19432 (N_19432,N_19161,N_19024);
nand U19433 (N_19433,N_19133,N_19216);
nand U19434 (N_19434,N_19223,N_19117);
nand U19435 (N_19435,N_19181,N_19207);
nor U19436 (N_19436,N_19015,N_19226);
xor U19437 (N_19437,N_19193,N_19015);
or U19438 (N_19438,N_19097,N_19149);
or U19439 (N_19439,N_19147,N_19099);
xnor U19440 (N_19440,N_19009,N_19133);
or U19441 (N_19441,N_19174,N_19172);
xor U19442 (N_19442,N_19246,N_19174);
nor U19443 (N_19443,N_19147,N_19023);
nand U19444 (N_19444,N_19017,N_19103);
xnor U19445 (N_19445,N_19131,N_19052);
xor U19446 (N_19446,N_19187,N_19173);
and U19447 (N_19447,N_19042,N_19093);
and U19448 (N_19448,N_19243,N_19245);
and U19449 (N_19449,N_19076,N_19107);
xor U19450 (N_19450,N_19196,N_19068);
and U19451 (N_19451,N_19000,N_19229);
or U19452 (N_19452,N_19023,N_19150);
nand U19453 (N_19453,N_19026,N_19127);
xnor U19454 (N_19454,N_19149,N_19044);
xor U19455 (N_19455,N_19209,N_19195);
nand U19456 (N_19456,N_19061,N_19031);
or U19457 (N_19457,N_19246,N_19011);
xor U19458 (N_19458,N_19187,N_19079);
nor U19459 (N_19459,N_19136,N_19101);
nor U19460 (N_19460,N_19066,N_19031);
nor U19461 (N_19461,N_19030,N_19143);
and U19462 (N_19462,N_19195,N_19189);
nand U19463 (N_19463,N_19213,N_19028);
xor U19464 (N_19464,N_19026,N_19005);
xor U19465 (N_19465,N_19222,N_19045);
nor U19466 (N_19466,N_19170,N_19101);
or U19467 (N_19467,N_19003,N_19028);
nor U19468 (N_19468,N_19232,N_19178);
xor U19469 (N_19469,N_19040,N_19054);
nand U19470 (N_19470,N_19028,N_19005);
nor U19471 (N_19471,N_19205,N_19212);
nand U19472 (N_19472,N_19196,N_19137);
and U19473 (N_19473,N_19027,N_19197);
nor U19474 (N_19474,N_19037,N_19238);
and U19475 (N_19475,N_19200,N_19175);
nor U19476 (N_19476,N_19144,N_19105);
or U19477 (N_19477,N_19187,N_19228);
and U19478 (N_19478,N_19246,N_19132);
nor U19479 (N_19479,N_19249,N_19101);
nand U19480 (N_19480,N_19225,N_19048);
nand U19481 (N_19481,N_19065,N_19172);
nand U19482 (N_19482,N_19222,N_19132);
nand U19483 (N_19483,N_19217,N_19103);
nand U19484 (N_19484,N_19139,N_19026);
or U19485 (N_19485,N_19235,N_19189);
or U19486 (N_19486,N_19018,N_19048);
or U19487 (N_19487,N_19034,N_19179);
nand U19488 (N_19488,N_19073,N_19190);
nor U19489 (N_19489,N_19239,N_19038);
and U19490 (N_19490,N_19189,N_19159);
nand U19491 (N_19491,N_19026,N_19029);
and U19492 (N_19492,N_19122,N_19095);
nand U19493 (N_19493,N_19245,N_19235);
nor U19494 (N_19494,N_19182,N_19028);
and U19495 (N_19495,N_19085,N_19062);
and U19496 (N_19496,N_19148,N_19137);
xnor U19497 (N_19497,N_19069,N_19010);
nor U19498 (N_19498,N_19237,N_19189);
nand U19499 (N_19499,N_19039,N_19169);
xnor U19500 (N_19500,N_19489,N_19342);
and U19501 (N_19501,N_19407,N_19394);
and U19502 (N_19502,N_19441,N_19393);
and U19503 (N_19503,N_19308,N_19424);
or U19504 (N_19504,N_19434,N_19472);
nand U19505 (N_19505,N_19495,N_19476);
xor U19506 (N_19506,N_19259,N_19277);
or U19507 (N_19507,N_19387,N_19483);
nor U19508 (N_19508,N_19400,N_19296);
or U19509 (N_19509,N_19297,N_19498);
nand U19510 (N_19510,N_19363,N_19492);
and U19511 (N_19511,N_19262,N_19401);
or U19512 (N_19512,N_19357,N_19285);
nand U19513 (N_19513,N_19250,N_19331);
nor U19514 (N_19514,N_19328,N_19344);
nand U19515 (N_19515,N_19300,N_19379);
or U19516 (N_19516,N_19366,N_19444);
nor U19517 (N_19517,N_19390,N_19372);
or U19518 (N_19518,N_19327,N_19337);
xor U19519 (N_19519,N_19384,N_19375);
or U19520 (N_19520,N_19257,N_19431);
xor U19521 (N_19521,N_19332,N_19399);
xor U19522 (N_19522,N_19486,N_19360);
nand U19523 (N_19523,N_19348,N_19382);
and U19524 (N_19524,N_19345,N_19406);
and U19525 (N_19525,N_19352,N_19349);
nand U19526 (N_19526,N_19474,N_19397);
nand U19527 (N_19527,N_19252,N_19282);
and U19528 (N_19528,N_19435,N_19450);
nor U19529 (N_19529,N_19370,N_19485);
or U19530 (N_19530,N_19283,N_19267);
nand U19531 (N_19531,N_19288,N_19364);
xor U19532 (N_19532,N_19254,N_19494);
nand U19533 (N_19533,N_19471,N_19361);
or U19534 (N_19534,N_19430,N_19405);
and U19535 (N_19535,N_19323,N_19335);
nand U19536 (N_19536,N_19478,N_19266);
nor U19537 (N_19537,N_19278,N_19313);
and U19538 (N_19538,N_19449,N_19272);
nand U19539 (N_19539,N_19388,N_19301);
nor U19540 (N_19540,N_19263,N_19462);
xnor U19541 (N_19541,N_19341,N_19417);
and U19542 (N_19542,N_19420,N_19421);
or U19543 (N_19543,N_19460,N_19487);
or U19544 (N_19544,N_19355,N_19322);
and U19545 (N_19545,N_19347,N_19311);
xor U19546 (N_19546,N_19412,N_19351);
nand U19547 (N_19547,N_19496,N_19446);
nor U19548 (N_19548,N_19287,N_19423);
and U19549 (N_19549,N_19383,N_19398);
or U19550 (N_19550,N_19378,N_19426);
or U19551 (N_19551,N_19251,N_19289);
nand U19552 (N_19552,N_19330,N_19261);
or U19553 (N_19553,N_19353,N_19447);
xnor U19554 (N_19554,N_19377,N_19481);
or U19555 (N_19555,N_19437,N_19359);
or U19556 (N_19556,N_19368,N_19350);
xnor U19557 (N_19557,N_19461,N_19310);
nor U19558 (N_19558,N_19376,N_19336);
and U19559 (N_19559,N_19281,N_19291);
nand U19560 (N_19560,N_19258,N_19438);
nor U19561 (N_19561,N_19373,N_19318);
nand U19562 (N_19562,N_19326,N_19292);
or U19563 (N_19563,N_19455,N_19454);
nor U19564 (N_19564,N_19419,N_19451);
or U19565 (N_19565,N_19395,N_19439);
and U19566 (N_19566,N_19403,N_19470);
and U19567 (N_19567,N_19429,N_19271);
nand U19568 (N_19568,N_19414,N_19428);
or U19569 (N_19569,N_19380,N_19443);
xor U19570 (N_19570,N_19365,N_19367);
nand U19571 (N_19571,N_19298,N_19409);
nor U19572 (N_19572,N_19309,N_19427);
nor U19573 (N_19573,N_19402,N_19491);
nor U19574 (N_19574,N_19416,N_19269);
or U19575 (N_19575,N_19410,N_19415);
xor U19576 (N_19576,N_19457,N_19276);
or U19577 (N_19577,N_19480,N_19404);
and U19578 (N_19578,N_19264,N_19280);
nor U19579 (N_19579,N_19303,N_19268);
and U19580 (N_19580,N_19468,N_19466);
xor U19581 (N_19581,N_19334,N_19381);
nor U19582 (N_19582,N_19343,N_19293);
nor U19583 (N_19583,N_19473,N_19315);
nand U19584 (N_19584,N_19445,N_19294);
or U19585 (N_19585,N_19385,N_19340);
nor U19586 (N_19586,N_19433,N_19255);
xnor U19587 (N_19587,N_19463,N_19452);
nor U19588 (N_19588,N_19354,N_19490);
and U19589 (N_19589,N_19392,N_19339);
nand U19590 (N_19590,N_19456,N_19346);
nand U19591 (N_19591,N_19493,N_19448);
or U19592 (N_19592,N_19418,N_19432);
or U19593 (N_19593,N_19464,N_19273);
nor U19594 (N_19594,N_19411,N_19499);
nand U19595 (N_19595,N_19302,N_19307);
and U19596 (N_19596,N_19319,N_19358);
xor U19597 (N_19597,N_19479,N_19274);
nand U19598 (N_19598,N_19270,N_19482);
xnor U19599 (N_19599,N_19275,N_19484);
xnor U19600 (N_19600,N_19436,N_19316);
xor U19601 (N_19601,N_19290,N_19459);
xor U19602 (N_19602,N_19362,N_19413);
nand U19603 (N_19603,N_19425,N_19333);
and U19604 (N_19604,N_19465,N_19253);
and U19605 (N_19605,N_19304,N_19325);
or U19606 (N_19606,N_19467,N_19295);
nor U19607 (N_19607,N_19386,N_19312);
xnor U19608 (N_19608,N_19408,N_19306);
and U19609 (N_19609,N_19314,N_19389);
or U19610 (N_19610,N_19391,N_19453);
nor U19611 (N_19611,N_19469,N_19497);
nor U19612 (N_19612,N_19324,N_19422);
nor U19613 (N_19613,N_19320,N_19305);
or U19614 (N_19614,N_19356,N_19286);
and U19615 (N_19615,N_19442,N_19458);
xor U19616 (N_19616,N_19396,N_19299);
nor U19617 (N_19617,N_19317,N_19256);
xnor U19618 (N_19618,N_19321,N_19371);
and U19619 (N_19619,N_19475,N_19488);
nand U19620 (N_19620,N_19440,N_19374);
or U19621 (N_19621,N_19477,N_19279);
nor U19622 (N_19622,N_19284,N_19338);
nor U19623 (N_19623,N_19260,N_19265);
nand U19624 (N_19624,N_19329,N_19369);
xnor U19625 (N_19625,N_19302,N_19409);
nor U19626 (N_19626,N_19470,N_19280);
or U19627 (N_19627,N_19387,N_19326);
xor U19628 (N_19628,N_19353,N_19324);
or U19629 (N_19629,N_19307,N_19410);
nand U19630 (N_19630,N_19449,N_19478);
or U19631 (N_19631,N_19324,N_19359);
nand U19632 (N_19632,N_19473,N_19314);
nand U19633 (N_19633,N_19494,N_19460);
nand U19634 (N_19634,N_19438,N_19370);
nor U19635 (N_19635,N_19396,N_19494);
nor U19636 (N_19636,N_19295,N_19326);
or U19637 (N_19637,N_19457,N_19302);
xor U19638 (N_19638,N_19463,N_19496);
nor U19639 (N_19639,N_19312,N_19437);
or U19640 (N_19640,N_19352,N_19254);
and U19641 (N_19641,N_19379,N_19493);
xnor U19642 (N_19642,N_19442,N_19339);
or U19643 (N_19643,N_19384,N_19455);
nor U19644 (N_19644,N_19359,N_19275);
nand U19645 (N_19645,N_19467,N_19367);
nand U19646 (N_19646,N_19417,N_19489);
or U19647 (N_19647,N_19299,N_19371);
nor U19648 (N_19648,N_19257,N_19369);
nand U19649 (N_19649,N_19348,N_19468);
or U19650 (N_19650,N_19258,N_19283);
xor U19651 (N_19651,N_19419,N_19388);
or U19652 (N_19652,N_19323,N_19266);
nand U19653 (N_19653,N_19430,N_19461);
and U19654 (N_19654,N_19321,N_19364);
nand U19655 (N_19655,N_19478,N_19443);
xnor U19656 (N_19656,N_19262,N_19337);
nand U19657 (N_19657,N_19298,N_19399);
nand U19658 (N_19658,N_19446,N_19316);
and U19659 (N_19659,N_19330,N_19259);
nor U19660 (N_19660,N_19288,N_19291);
and U19661 (N_19661,N_19345,N_19297);
or U19662 (N_19662,N_19480,N_19266);
and U19663 (N_19663,N_19334,N_19291);
nor U19664 (N_19664,N_19333,N_19436);
and U19665 (N_19665,N_19279,N_19309);
xor U19666 (N_19666,N_19356,N_19306);
or U19667 (N_19667,N_19304,N_19343);
xor U19668 (N_19668,N_19270,N_19422);
or U19669 (N_19669,N_19291,N_19426);
nor U19670 (N_19670,N_19292,N_19435);
or U19671 (N_19671,N_19281,N_19353);
nand U19672 (N_19672,N_19271,N_19411);
or U19673 (N_19673,N_19472,N_19328);
nand U19674 (N_19674,N_19407,N_19418);
nand U19675 (N_19675,N_19426,N_19429);
nor U19676 (N_19676,N_19410,N_19339);
xor U19677 (N_19677,N_19473,N_19303);
or U19678 (N_19678,N_19313,N_19460);
nand U19679 (N_19679,N_19494,N_19481);
or U19680 (N_19680,N_19433,N_19422);
xnor U19681 (N_19681,N_19287,N_19349);
and U19682 (N_19682,N_19302,N_19420);
and U19683 (N_19683,N_19369,N_19462);
nor U19684 (N_19684,N_19314,N_19412);
or U19685 (N_19685,N_19497,N_19447);
or U19686 (N_19686,N_19466,N_19375);
xnor U19687 (N_19687,N_19408,N_19400);
or U19688 (N_19688,N_19298,N_19254);
nand U19689 (N_19689,N_19470,N_19346);
nand U19690 (N_19690,N_19432,N_19499);
xor U19691 (N_19691,N_19487,N_19499);
nand U19692 (N_19692,N_19462,N_19456);
nor U19693 (N_19693,N_19335,N_19299);
nor U19694 (N_19694,N_19317,N_19257);
nor U19695 (N_19695,N_19464,N_19473);
xor U19696 (N_19696,N_19364,N_19404);
or U19697 (N_19697,N_19264,N_19455);
nand U19698 (N_19698,N_19289,N_19407);
or U19699 (N_19699,N_19392,N_19440);
or U19700 (N_19700,N_19485,N_19425);
nand U19701 (N_19701,N_19379,N_19277);
and U19702 (N_19702,N_19325,N_19416);
nor U19703 (N_19703,N_19420,N_19493);
xor U19704 (N_19704,N_19381,N_19437);
nand U19705 (N_19705,N_19466,N_19491);
nor U19706 (N_19706,N_19262,N_19324);
or U19707 (N_19707,N_19412,N_19353);
nor U19708 (N_19708,N_19392,N_19475);
nor U19709 (N_19709,N_19454,N_19283);
xor U19710 (N_19710,N_19361,N_19306);
xnor U19711 (N_19711,N_19384,N_19293);
or U19712 (N_19712,N_19327,N_19312);
and U19713 (N_19713,N_19314,N_19399);
xnor U19714 (N_19714,N_19313,N_19256);
nor U19715 (N_19715,N_19255,N_19481);
and U19716 (N_19716,N_19492,N_19383);
nand U19717 (N_19717,N_19379,N_19252);
xnor U19718 (N_19718,N_19301,N_19355);
nor U19719 (N_19719,N_19377,N_19472);
nand U19720 (N_19720,N_19292,N_19479);
nor U19721 (N_19721,N_19475,N_19324);
xnor U19722 (N_19722,N_19386,N_19378);
nand U19723 (N_19723,N_19471,N_19294);
xnor U19724 (N_19724,N_19418,N_19448);
xnor U19725 (N_19725,N_19398,N_19481);
nor U19726 (N_19726,N_19336,N_19321);
and U19727 (N_19727,N_19482,N_19498);
and U19728 (N_19728,N_19447,N_19311);
xor U19729 (N_19729,N_19428,N_19416);
nor U19730 (N_19730,N_19395,N_19458);
nand U19731 (N_19731,N_19422,N_19316);
and U19732 (N_19732,N_19498,N_19291);
nand U19733 (N_19733,N_19310,N_19291);
xnor U19734 (N_19734,N_19357,N_19266);
nor U19735 (N_19735,N_19371,N_19495);
xnor U19736 (N_19736,N_19399,N_19455);
and U19737 (N_19737,N_19404,N_19397);
xnor U19738 (N_19738,N_19472,N_19368);
nand U19739 (N_19739,N_19498,N_19474);
nor U19740 (N_19740,N_19452,N_19320);
or U19741 (N_19741,N_19410,N_19370);
and U19742 (N_19742,N_19467,N_19449);
nand U19743 (N_19743,N_19449,N_19295);
and U19744 (N_19744,N_19296,N_19453);
xor U19745 (N_19745,N_19332,N_19270);
and U19746 (N_19746,N_19263,N_19435);
nand U19747 (N_19747,N_19374,N_19472);
xor U19748 (N_19748,N_19347,N_19310);
and U19749 (N_19749,N_19473,N_19460);
and U19750 (N_19750,N_19675,N_19668);
nand U19751 (N_19751,N_19591,N_19602);
xnor U19752 (N_19752,N_19710,N_19605);
or U19753 (N_19753,N_19533,N_19549);
xor U19754 (N_19754,N_19593,N_19665);
nor U19755 (N_19755,N_19679,N_19644);
or U19756 (N_19756,N_19589,N_19632);
nand U19757 (N_19757,N_19624,N_19596);
xnor U19758 (N_19758,N_19685,N_19625);
and U19759 (N_19759,N_19647,N_19555);
xor U19760 (N_19760,N_19699,N_19513);
or U19761 (N_19761,N_19671,N_19725);
xnor U19762 (N_19762,N_19515,N_19505);
xor U19763 (N_19763,N_19662,N_19709);
or U19764 (N_19764,N_19563,N_19693);
nand U19765 (N_19765,N_19580,N_19615);
or U19766 (N_19766,N_19733,N_19567);
or U19767 (N_19767,N_19546,N_19690);
nand U19768 (N_19768,N_19527,N_19538);
nand U19769 (N_19769,N_19528,N_19559);
nand U19770 (N_19770,N_19719,N_19748);
and U19771 (N_19771,N_19749,N_19557);
or U19772 (N_19772,N_19648,N_19734);
and U19773 (N_19773,N_19636,N_19548);
xnor U19774 (N_19774,N_19703,N_19728);
nor U19775 (N_19775,N_19518,N_19583);
or U19776 (N_19776,N_19740,N_19657);
nor U19777 (N_19777,N_19678,N_19697);
or U19778 (N_19778,N_19738,N_19623);
nand U19779 (N_19779,N_19638,N_19512);
and U19780 (N_19780,N_19627,N_19706);
xor U19781 (N_19781,N_19698,N_19715);
nor U19782 (N_19782,N_19726,N_19532);
xnor U19783 (N_19783,N_19658,N_19737);
nor U19784 (N_19784,N_19607,N_19611);
nand U19785 (N_19785,N_19552,N_19574);
nand U19786 (N_19786,N_19735,N_19556);
and U19787 (N_19787,N_19742,N_19634);
or U19788 (N_19788,N_19551,N_19521);
and U19789 (N_19789,N_19718,N_19650);
or U19790 (N_19790,N_19722,N_19641);
or U19791 (N_19791,N_19586,N_19585);
and U19792 (N_19792,N_19656,N_19674);
and U19793 (N_19793,N_19616,N_19629);
or U19794 (N_19794,N_19716,N_19731);
nand U19795 (N_19795,N_19603,N_19601);
and U19796 (N_19796,N_19542,N_19696);
or U19797 (N_19797,N_19536,N_19522);
nand U19798 (N_19798,N_19677,N_19570);
xor U19799 (N_19799,N_19577,N_19640);
or U19800 (N_19800,N_19621,N_19729);
and U19801 (N_19801,N_19507,N_19712);
and U19802 (N_19802,N_19573,N_19612);
and U19803 (N_19803,N_19565,N_19724);
or U19804 (N_19804,N_19687,N_19720);
xor U19805 (N_19805,N_19702,N_19592);
nor U19806 (N_19806,N_19526,N_19608);
nand U19807 (N_19807,N_19637,N_19587);
xnor U19808 (N_19808,N_19569,N_19584);
nand U19809 (N_19809,N_19689,N_19504);
or U19810 (N_19810,N_19721,N_19568);
and U19811 (N_19811,N_19550,N_19564);
and U19812 (N_19812,N_19561,N_19683);
xnor U19813 (N_19813,N_19649,N_19540);
nand U19814 (N_19814,N_19610,N_19705);
and U19815 (N_19815,N_19578,N_19654);
nor U19816 (N_19816,N_19520,N_19660);
and U19817 (N_19817,N_19597,N_19673);
and U19818 (N_19818,N_19743,N_19509);
xor U19819 (N_19819,N_19711,N_19713);
or U19820 (N_19820,N_19730,N_19708);
and U19821 (N_19821,N_19506,N_19562);
nand U19822 (N_19822,N_19579,N_19667);
or U19823 (N_19823,N_19739,N_19599);
nor U19824 (N_19824,N_19595,N_19723);
and U19825 (N_19825,N_19663,N_19736);
nor U19826 (N_19826,N_19745,N_19566);
or U19827 (N_19827,N_19501,N_19626);
and U19828 (N_19828,N_19516,N_19541);
xnor U19829 (N_19829,N_19620,N_19514);
and U19830 (N_19830,N_19553,N_19590);
xor U19831 (N_19831,N_19511,N_19628);
xor U19832 (N_19832,N_19717,N_19519);
nand U19833 (N_19833,N_19622,N_19682);
nor U19834 (N_19834,N_19670,N_19609);
or U19835 (N_19835,N_19571,N_19672);
nor U19836 (N_19836,N_19617,N_19664);
and U19837 (N_19837,N_19535,N_19545);
nor U19838 (N_19838,N_19686,N_19732);
nor U19839 (N_19839,N_19543,N_19695);
nand U19840 (N_19840,N_19714,N_19618);
or U19841 (N_19841,N_19529,N_19544);
or U19842 (N_19842,N_19500,N_19539);
or U19843 (N_19843,N_19508,N_19614);
nand U19844 (N_19844,N_19680,N_19534);
or U19845 (N_19845,N_19510,N_19704);
and U19846 (N_19846,N_19619,N_19502);
or U19847 (N_19847,N_19594,N_19701);
and U19848 (N_19848,N_19631,N_19531);
nand U19849 (N_19849,N_19524,N_19581);
nand U19850 (N_19850,N_19642,N_19659);
nand U19851 (N_19851,N_19694,N_19669);
nand U19852 (N_19852,N_19646,N_19630);
and U19853 (N_19853,N_19684,N_19588);
nand U19854 (N_19854,N_19681,N_19558);
xor U19855 (N_19855,N_19576,N_19744);
and U19856 (N_19856,N_19606,N_19517);
xor U19857 (N_19857,N_19547,N_19572);
and U19858 (N_19858,N_19741,N_19653);
nand U19859 (N_19859,N_19700,N_19613);
and U19860 (N_19860,N_19598,N_19600);
and U19861 (N_19861,N_19651,N_19666);
xor U19862 (N_19862,N_19575,N_19661);
or U19863 (N_19863,N_19639,N_19655);
xor U19864 (N_19864,N_19635,N_19523);
nand U19865 (N_19865,N_19746,N_19747);
and U19866 (N_19866,N_19652,N_19688);
nand U19867 (N_19867,N_19691,N_19554);
or U19868 (N_19868,N_19676,N_19633);
nand U19869 (N_19869,N_19692,N_19645);
xor U19870 (N_19870,N_19604,N_19560);
xnor U19871 (N_19871,N_19503,N_19727);
nor U19872 (N_19872,N_19643,N_19525);
or U19873 (N_19873,N_19707,N_19530);
xor U19874 (N_19874,N_19537,N_19582);
and U19875 (N_19875,N_19742,N_19717);
nand U19876 (N_19876,N_19653,N_19549);
nor U19877 (N_19877,N_19563,N_19729);
or U19878 (N_19878,N_19624,N_19646);
or U19879 (N_19879,N_19735,N_19647);
nor U19880 (N_19880,N_19601,N_19714);
or U19881 (N_19881,N_19673,N_19737);
xnor U19882 (N_19882,N_19666,N_19699);
or U19883 (N_19883,N_19731,N_19743);
or U19884 (N_19884,N_19734,N_19699);
or U19885 (N_19885,N_19509,N_19608);
nand U19886 (N_19886,N_19544,N_19532);
or U19887 (N_19887,N_19645,N_19548);
nand U19888 (N_19888,N_19630,N_19701);
or U19889 (N_19889,N_19663,N_19709);
xnor U19890 (N_19890,N_19560,N_19525);
or U19891 (N_19891,N_19550,N_19724);
nor U19892 (N_19892,N_19642,N_19579);
nand U19893 (N_19893,N_19574,N_19657);
nand U19894 (N_19894,N_19718,N_19647);
and U19895 (N_19895,N_19580,N_19730);
and U19896 (N_19896,N_19743,N_19661);
or U19897 (N_19897,N_19611,N_19687);
and U19898 (N_19898,N_19581,N_19578);
or U19899 (N_19899,N_19533,N_19739);
nor U19900 (N_19900,N_19662,N_19630);
nand U19901 (N_19901,N_19588,N_19652);
nor U19902 (N_19902,N_19581,N_19692);
nor U19903 (N_19903,N_19624,N_19643);
nor U19904 (N_19904,N_19728,N_19579);
nand U19905 (N_19905,N_19523,N_19651);
xor U19906 (N_19906,N_19608,N_19555);
nor U19907 (N_19907,N_19714,N_19572);
and U19908 (N_19908,N_19729,N_19503);
and U19909 (N_19909,N_19512,N_19564);
xnor U19910 (N_19910,N_19734,N_19552);
and U19911 (N_19911,N_19573,N_19524);
nand U19912 (N_19912,N_19692,N_19587);
and U19913 (N_19913,N_19732,N_19630);
xor U19914 (N_19914,N_19748,N_19675);
or U19915 (N_19915,N_19625,N_19551);
nor U19916 (N_19916,N_19563,N_19601);
or U19917 (N_19917,N_19532,N_19503);
nor U19918 (N_19918,N_19735,N_19661);
nand U19919 (N_19919,N_19523,N_19578);
nand U19920 (N_19920,N_19679,N_19633);
xnor U19921 (N_19921,N_19665,N_19575);
or U19922 (N_19922,N_19694,N_19603);
nand U19923 (N_19923,N_19601,N_19519);
or U19924 (N_19924,N_19513,N_19729);
or U19925 (N_19925,N_19730,N_19636);
and U19926 (N_19926,N_19606,N_19698);
nand U19927 (N_19927,N_19551,N_19726);
and U19928 (N_19928,N_19731,N_19556);
xor U19929 (N_19929,N_19629,N_19729);
or U19930 (N_19930,N_19683,N_19631);
xor U19931 (N_19931,N_19660,N_19564);
nor U19932 (N_19932,N_19508,N_19714);
xnor U19933 (N_19933,N_19667,N_19540);
nand U19934 (N_19934,N_19727,N_19722);
and U19935 (N_19935,N_19628,N_19575);
nand U19936 (N_19936,N_19597,N_19622);
or U19937 (N_19937,N_19575,N_19534);
nand U19938 (N_19938,N_19577,N_19563);
nor U19939 (N_19939,N_19501,N_19622);
xor U19940 (N_19940,N_19615,N_19644);
or U19941 (N_19941,N_19736,N_19538);
nor U19942 (N_19942,N_19692,N_19737);
nand U19943 (N_19943,N_19632,N_19646);
nand U19944 (N_19944,N_19557,N_19707);
or U19945 (N_19945,N_19567,N_19500);
xnor U19946 (N_19946,N_19632,N_19505);
or U19947 (N_19947,N_19722,N_19519);
xor U19948 (N_19948,N_19567,N_19626);
nor U19949 (N_19949,N_19557,N_19663);
nor U19950 (N_19950,N_19739,N_19629);
nor U19951 (N_19951,N_19593,N_19556);
and U19952 (N_19952,N_19689,N_19725);
nor U19953 (N_19953,N_19570,N_19662);
nor U19954 (N_19954,N_19514,N_19734);
xnor U19955 (N_19955,N_19628,N_19502);
or U19956 (N_19956,N_19736,N_19622);
xor U19957 (N_19957,N_19574,N_19672);
and U19958 (N_19958,N_19566,N_19662);
xnor U19959 (N_19959,N_19602,N_19501);
nand U19960 (N_19960,N_19602,N_19647);
or U19961 (N_19961,N_19698,N_19744);
nand U19962 (N_19962,N_19589,N_19563);
and U19963 (N_19963,N_19549,N_19525);
or U19964 (N_19964,N_19676,N_19622);
xnor U19965 (N_19965,N_19740,N_19613);
nand U19966 (N_19966,N_19565,N_19669);
and U19967 (N_19967,N_19714,N_19709);
and U19968 (N_19968,N_19706,N_19605);
nand U19969 (N_19969,N_19556,N_19720);
nor U19970 (N_19970,N_19603,N_19520);
and U19971 (N_19971,N_19608,N_19620);
nor U19972 (N_19972,N_19735,N_19676);
nor U19973 (N_19973,N_19641,N_19749);
nand U19974 (N_19974,N_19618,N_19539);
xnor U19975 (N_19975,N_19699,N_19546);
and U19976 (N_19976,N_19500,N_19704);
and U19977 (N_19977,N_19727,N_19652);
and U19978 (N_19978,N_19747,N_19636);
xor U19979 (N_19979,N_19532,N_19595);
nor U19980 (N_19980,N_19732,N_19525);
or U19981 (N_19981,N_19688,N_19612);
nand U19982 (N_19982,N_19651,N_19716);
or U19983 (N_19983,N_19712,N_19609);
nand U19984 (N_19984,N_19696,N_19682);
or U19985 (N_19985,N_19689,N_19514);
and U19986 (N_19986,N_19540,N_19738);
nor U19987 (N_19987,N_19599,N_19733);
or U19988 (N_19988,N_19604,N_19746);
nand U19989 (N_19989,N_19680,N_19504);
nand U19990 (N_19990,N_19675,N_19526);
and U19991 (N_19991,N_19625,N_19678);
and U19992 (N_19992,N_19643,N_19696);
or U19993 (N_19993,N_19582,N_19738);
nor U19994 (N_19994,N_19542,N_19716);
nand U19995 (N_19995,N_19742,N_19641);
nand U19996 (N_19996,N_19583,N_19554);
nand U19997 (N_19997,N_19592,N_19609);
nand U19998 (N_19998,N_19632,N_19640);
or U19999 (N_19999,N_19662,N_19619);
nand UO_0 (O_0,N_19837,N_19985);
and UO_1 (O_1,N_19804,N_19991);
and UO_2 (O_2,N_19949,N_19953);
nor UO_3 (O_3,N_19814,N_19931);
nor UO_4 (O_4,N_19973,N_19938);
nor UO_5 (O_5,N_19900,N_19848);
xnor UO_6 (O_6,N_19901,N_19936);
nor UO_7 (O_7,N_19779,N_19855);
nand UO_8 (O_8,N_19939,N_19959);
nand UO_9 (O_9,N_19849,N_19926);
and UO_10 (O_10,N_19917,N_19792);
nor UO_11 (O_11,N_19839,N_19961);
nand UO_12 (O_12,N_19971,N_19751);
or UO_13 (O_13,N_19811,N_19881);
or UO_14 (O_14,N_19913,N_19944);
nor UO_15 (O_15,N_19977,N_19907);
or UO_16 (O_16,N_19833,N_19873);
nand UO_17 (O_17,N_19951,N_19947);
nand UO_18 (O_18,N_19882,N_19864);
and UO_19 (O_19,N_19980,N_19797);
nor UO_20 (O_20,N_19821,N_19825);
nand UO_21 (O_21,N_19893,N_19834);
nand UO_22 (O_22,N_19762,N_19874);
nor UO_23 (O_23,N_19948,N_19851);
or UO_24 (O_24,N_19831,N_19754);
and UO_25 (O_25,N_19856,N_19803);
or UO_26 (O_26,N_19776,N_19924);
nor UO_27 (O_27,N_19880,N_19940);
and UO_28 (O_28,N_19784,N_19935);
or UO_29 (O_29,N_19927,N_19863);
and UO_30 (O_30,N_19807,N_19962);
and UO_31 (O_31,N_19758,N_19846);
or UO_32 (O_32,N_19889,N_19958);
xnor UO_33 (O_33,N_19918,N_19823);
and UO_34 (O_34,N_19755,N_19905);
nor UO_35 (O_35,N_19921,N_19794);
nor UO_36 (O_36,N_19995,N_19885);
xnor UO_37 (O_37,N_19795,N_19802);
nor UO_38 (O_38,N_19876,N_19812);
or UO_39 (O_39,N_19816,N_19820);
or UO_40 (O_40,N_19886,N_19916);
nor UO_41 (O_41,N_19950,N_19832);
nand UO_42 (O_42,N_19994,N_19999);
xor UO_43 (O_43,N_19860,N_19750);
and UO_44 (O_44,N_19857,N_19915);
or UO_45 (O_45,N_19978,N_19819);
or UO_46 (O_46,N_19796,N_19782);
and UO_47 (O_47,N_19898,N_19790);
or UO_48 (O_48,N_19909,N_19764);
or UO_49 (O_49,N_19967,N_19847);
nor UO_50 (O_50,N_19853,N_19810);
and UO_51 (O_51,N_19897,N_19968);
or UO_52 (O_52,N_19911,N_19791);
nor UO_53 (O_53,N_19761,N_19894);
nor UO_54 (O_54,N_19888,N_19861);
xnor UO_55 (O_55,N_19793,N_19982);
or UO_56 (O_56,N_19925,N_19786);
xor UO_57 (O_57,N_19989,N_19799);
xor UO_58 (O_58,N_19914,N_19941);
nor UO_59 (O_59,N_19870,N_19983);
nand UO_60 (O_60,N_19988,N_19840);
xnor UO_61 (O_61,N_19890,N_19970);
and UO_62 (O_62,N_19960,N_19932);
and UO_63 (O_63,N_19767,N_19878);
nand UO_64 (O_64,N_19867,N_19829);
nand UO_65 (O_65,N_19892,N_19929);
and UO_66 (O_66,N_19969,N_19923);
nor UO_67 (O_67,N_19800,N_19809);
and UO_68 (O_68,N_19906,N_19842);
or UO_69 (O_69,N_19843,N_19976);
nand UO_70 (O_70,N_19963,N_19763);
or UO_71 (O_71,N_19770,N_19818);
and UO_72 (O_72,N_19835,N_19928);
and UO_73 (O_73,N_19954,N_19753);
nor UO_74 (O_74,N_19805,N_19903);
nand UO_75 (O_75,N_19775,N_19788);
nand UO_76 (O_76,N_19752,N_19922);
xor UO_77 (O_77,N_19986,N_19854);
and UO_78 (O_78,N_19828,N_19964);
or UO_79 (O_79,N_19827,N_19992);
nor UO_80 (O_80,N_19930,N_19887);
nor UO_81 (O_81,N_19801,N_19824);
and UO_82 (O_82,N_19815,N_19822);
xor UO_83 (O_83,N_19912,N_19836);
nand UO_84 (O_84,N_19768,N_19757);
nor UO_85 (O_85,N_19841,N_19956);
and UO_86 (O_86,N_19875,N_19965);
and UO_87 (O_87,N_19896,N_19979);
nor UO_88 (O_88,N_19871,N_19780);
nor UO_89 (O_89,N_19883,N_19877);
and UO_90 (O_90,N_19765,N_19937);
or UO_91 (O_91,N_19879,N_19769);
xnor UO_92 (O_92,N_19984,N_19785);
nand UO_93 (O_93,N_19774,N_19902);
and UO_94 (O_94,N_19760,N_19899);
nor UO_95 (O_95,N_19996,N_19966);
or UO_96 (O_96,N_19838,N_19972);
and UO_97 (O_97,N_19981,N_19771);
nor UO_98 (O_98,N_19756,N_19993);
and UO_99 (O_99,N_19830,N_19952);
xor UO_100 (O_100,N_19808,N_19783);
nand UO_101 (O_101,N_19919,N_19895);
nand UO_102 (O_102,N_19934,N_19813);
or UO_103 (O_103,N_19987,N_19865);
nor UO_104 (O_104,N_19773,N_19759);
and UO_105 (O_105,N_19910,N_19974);
nor UO_106 (O_106,N_19858,N_19789);
nor UO_107 (O_107,N_19777,N_19798);
nand UO_108 (O_108,N_19957,N_19998);
and UO_109 (O_109,N_19766,N_19826);
nand UO_110 (O_110,N_19866,N_19946);
nand UO_111 (O_111,N_19904,N_19844);
nand UO_112 (O_112,N_19869,N_19772);
nor UO_113 (O_113,N_19850,N_19884);
xnor UO_114 (O_114,N_19942,N_19997);
nor UO_115 (O_115,N_19933,N_19778);
nor UO_116 (O_116,N_19859,N_19990);
or UO_117 (O_117,N_19817,N_19787);
and UO_118 (O_118,N_19891,N_19781);
and UO_119 (O_119,N_19975,N_19908);
nor UO_120 (O_120,N_19862,N_19845);
nor UO_121 (O_121,N_19945,N_19868);
nor UO_122 (O_122,N_19872,N_19852);
nor UO_123 (O_123,N_19955,N_19920);
xnor UO_124 (O_124,N_19806,N_19943);
nor UO_125 (O_125,N_19867,N_19785);
and UO_126 (O_126,N_19785,N_19927);
nor UO_127 (O_127,N_19929,N_19960);
nor UO_128 (O_128,N_19940,N_19783);
nand UO_129 (O_129,N_19956,N_19985);
xor UO_130 (O_130,N_19967,N_19800);
and UO_131 (O_131,N_19948,N_19789);
nand UO_132 (O_132,N_19897,N_19771);
and UO_133 (O_133,N_19956,N_19855);
xnor UO_134 (O_134,N_19833,N_19978);
nor UO_135 (O_135,N_19817,N_19917);
nand UO_136 (O_136,N_19978,N_19930);
xor UO_137 (O_137,N_19944,N_19762);
nor UO_138 (O_138,N_19904,N_19768);
xor UO_139 (O_139,N_19887,N_19844);
nand UO_140 (O_140,N_19847,N_19906);
and UO_141 (O_141,N_19899,N_19849);
xor UO_142 (O_142,N_19858,N_19964);
xnor UO_143 (O_143,N_19789,N_19937);
or UO_144 (O_144,N_19954,N_19983);
or UO_145 (O_145,N_19840,N_19890);
or UO_146 (O_146,N_19790,N_19909);
and UO_147 (O_147,N_19855,N_19998);
nor UO_148 (O_148,N_19769,N_19992);
xnor UO_149 (O_149,N_19861,N_19789);
xnor UO_150 (O_150,N_19772,N_19998);
and UO_151 (O_151,N_19975,N_19833);
xor UO_152 (O_152,N_19757,N_19863);
nor UO_153 (O_153,N_19992,N_19983);
xor UO_154 (O_154,N_19785,N_19779);
and UO_155 (O_155,N_19940,N_19752);
xnor UO_156 (O_156,N_19912,N_19958);
nor UO_157 (O_157,N_19943,N_19871);
or UO_158 (O_158,N_19915,N_19844);
and UO_159 (O_159,N_19839,N_19834);
nor UO_160 (O_160,N_19820,N_19915);
nor UO_161 (O_161,N_19914,N_19998);
or UO_162 (O_162,N_19988,N_19907);
and UO_163 (O_163,N_19935,N_19861);
nor UO_164 (O_164,N_19763,N_19960);
or UO_165 (O_165,N_19811,N_19838);
nand UO_166 (O_166,N_19846,N_19996);
nand UO_167 (O_167,N_19761,N_19915);
or UO_168 (O_168,N_19803,N_19898);
xor UO_169 (O_169,N_19907,N_19997);
xor UO_170 (O_170,N_19959,N_19819);
and UO_171 (O_171,N_19818,N_19797);
and UO_172 (O_172,N_19814,N_19825);
nand UO_173 (O_173,N_19996,N_19839);
and UO_174 (O_174,N_19875,N_19999);
and UO_175 (O_175,N_19805,N_19917);
xnor UO_176 (O_176,N_19763,N_19846);
nor UO_177 (O_177,N_19808,N_19776);
xor UO_178 (O_178,N_19854,N_19903);
and UO_179 (O_179,N_19795,N_19871);
xnor UO_180 (O_180,N_19980,N_19771);
nand UO_181 (O_181,N_19947,N_19755);
and UO_182 (O_182,N_19840,N_19991);
or UO_183 (O_183,N_19806,N_19900);
and UO_184 (O_184,N_19870,N_19814);
xnor UO_185 (O_185,N_19871,N_19884);
or UO_186 (O_186,N_19780,N_19999);
or UO_187 (O_187,N_19766,N_19847);
nand UO_188 (O_188,N_19860,N_19925);
nand UO_189 (O_189,N_19774,N_19848);
nand UO_190 (O_190,N_19813,N_19957);
nor UO_191 (O_191,N_19999,N_19879);
nor UO_192 (O_192,N_19897,N_19999);
or UO_193 (O_193,N_19986,N_19822);
nand UO_194 (O_194,N_19916,N_19754);
xnor UO_195 (O_195,N_19986,N_19873);
nor UO_196 (O_196,N_19835,N_19917);
nor UO_197 (O_197,N_19895,N_19768);
nand UO_198 (O_198,N_19842,N_19870);
nor UO_199 (O_199,N_19867,N_19870);
or UO_200 (O_200,N_19881,N_19752);
xor UO_201 (O_201,N_19778,N_19838);
or UO_202 (O_202,N_19955,N_19931);
or UO_203 (O_203,N_19901,N_19792);
nand UO_204 (O_204,N_19917,N_19880);
nor UO_205 (O_205,N_19806,N_19925);
nor UO_206 (O_206,N_19859,N_19915);
xor UO_207 (O_207,N_19878,N_19862);
nand UO_208 (O_208,N_19792,N_19797);
or UO_209 (O_209,N_19895,N_19909);
nor UO_210 (O_210,N_19866,N_19894);
xnor UO_211 (O_211,N_19753,N_19991);
and UO_212 (O_212,N_19834,N_19877);
nand UO_213 (O_213,N_19770,N_19913);
or UO_214 (O_214,N_19759,N_19840);
and UO_215 (O_215,N_19943,N_19780);
nand UO_216 (O_216,N_19916,N_19906);
nand UO_217 (O_217,N_19773,N_19873);
and UO_218 (O_218,N_19860,N_19879);
nor UO_219 (O_219,N_19784,N_19861);
xnor UO_220 (O_220,N_19955,N_19914);
and UO_221 (O_221,N_19789,N_19911);
nor UO_222 (O_222,N_19783,N_19974);
and UO_223 (O_223,N_19820,N_19897);
or UO_224 (O_224,N_19771,N_19890);
xnor UO_225 (O_225,N_19834,N_19820);
xor UO_226 (O_226,N_19975,N_19811);
xnor UO_227 (O_227,N_19878,N_19962);
nor UO_228 (O_228,N_19927,N_19766);
and UO_229 (O_229,N_19897,N_19827);
nor UO_230 (O_230,N_19979,N_19916);
and UO_231 (O_231,N_19957,N_19942);
and UO_232 (O_232,N_19948,N_19995);
xor UO_233 (O_233,N_19800,N_19862);
and UO_234 (O_234,N_19847,N_19960);
xnor UO_235 (O_235,N_19978,N_19788);
and UO_236 (O_236,N_19891,N_19801);
or UO_237 (O_237,N_19926,N_19937);
nand UO_238 (O_238,N_19907,N_19996);
and UO_239 (O_239,N_19810,N_19957);
xor UO_240 (O_240,N_19929,N_19932);
nand UO_241 (O_241,N_19921,N_19870);
nand UO_242 (O_242,N_19955,N_19814);
or UO_243 (O_243,N_19818,N_19939);
nand UO_244 (O_244,N_19829,N_19792);
nor UO_245 (O_245,N_19860,N_19840);
nand UO_246 (O_246,N_19983,N_19812);
xnor UO_247 (O_247,N_19896,N_19885);
xnor UO_248 (O_248,N_19844,N_19829);
xnor UO_249 (O_249,N_19968,N_19964);
or UO_250 (O_250,N_19756,N_19948);
and UO_251 (O_251,N_19959,N_19966);
xor UO_252 (O_252,N_19838,N_19952);
or UO_253 (O_253,N_19917,N_19980);
nor UO_254 (O_254,N_19761,N_19940);
nand UO_255 (O_255,N_19823,N_19794);
nand UO_256 (O_256,N_19982,N_19770);
and UO_257 (O_257,N_19978,N_19835);
or UO_258 (O_258,N_19981,N_19890);
xnor UO_259 (O_259,N_19897,N_19780);
xor UO_260 (O_260,N_19921,N_19977);
nor UO_261 (O_261,N_19913,N_19867);
nand UO_262 (O_262,N_19978,N_19851);
xor UO_263 (O_263,N_19967,N_19966);
xnor UO_264 (O_264,N_19910,N_19821);
nand UO_265 (O_265,N_19827,N_19791);
or UO_266 (O_266,N_19810,N_19822);
xor UO_267 (O_267,N_19924,N_19786);
and UO_268 (O_268,N_19969,N_19809);
or UO_269 (O_269,N_19821,N_19963);
nand UO_270 (O_270,N_19948,N_19917);
or UO_271 (O_271,N_19975,N_19967);
nor UO_272 (O_272,N_19827,N_19810);
nand UO_273 (O_273,N_19860,N_19807);
xor UO_274 (O_274,N_19974,N_19796);
or UO_275 (O_275,N_19789,N_19817);
xor UO_276 (O_276,N_19838,N_19791);
and UO_277 (O_277,N_19917,N_19908);
and UO_278 (O_278,N_19846,N_19891);
nor UO_279 (O_279,N_19797,N_19813);
xnor UO_280 (O_280,N_19916,N_19790);
nor UO_281 (O_281,N_19791,N_19872);
and UO_282 (O_282,N_19888,N_19962);
or UO_283 (O_283,N_19967,N_19790);
nand UO_284 (O_284,N_19904,N_19851);
nor UO_285 (O_285,N_19936,N_19981);
nor UO_286 (O_286,N_19798,N_19823);
xnor UO_287 (O_287,N_19976,N_19880);
nand UO_288 (O_288,N_19771,N_19913);
nand UO_289 (O_289,N_19821,N_19861);
or UO_290 (O_290,N_19810,N_19770);
nand UO_291 (O_291,N_19930,N_19882);
or UO_292 (O_292,N_19849,N_19930);
nand UO_293 (O_293,N_19968,N_19936);
nor UO_294 (O_294,N_19948,N_19787);
or UO_295 (O_295,N_19786,N_19893);
xnor UO_296 (O_296,N_19874,N_19980);
nand UO_297 (O_297,N_19838,N_19752);
or UO_298 (O_298,N_19887,N_19777);
xor UO_299 (O_299,N_19898,N_19860);
and UO_300 (O_300,N_19889,N_19768);
nand UO_301 (O_301,N_19926,N_19890);
and UO_302 (O_302,N_19794,N_19998);
or UO_303 (O_303,N_19864,N_19860);
nand UO_304 (O_304,N_19979,N_19944);
nand UO_305 (O_305,N_19866,N_19862);
xor UO_306 (O_306,N_19964,N_19865);
or UO_307 (O_307,N_19858,N_19907);
and UO_308 (O_308,N_19857,N_19903);
xor UO_309 (O_309,N_19997,N_19809);
or UO_310 (O_310,N_19964,N_19901);
nor UO_311 (O_311,N_19948,N_19845);
xnor UO_312 (O_312,N_19882,N_19821);
or UO_313 (O_313,N_19836,N_19826);
nor UO_314 (O_314,N_19914,N_19925);
and UO_315 (O_315,N_19973,N_19820);
nand UO_316 (O_316,N_19860,N_19801);
nor UO_317 (O_317,N_19848,N_19968);
nor UO_318 (O_318,N_19845,N_19817);
nand UO_319 (O_319,N_19883,N_19825);
xor UO_320 (O_320,N_19871,N_19925);
nor UO_321 (O_321,N_19917,N_19891);
nor UO_322 (O_322,N_19942,N_19812);
nor UO_323 (O_323,N_19797,N_19834);
or UO_324 (O_324,N_19984,N_19965);
xnor UO_325 (O_325,N_19984,N_19782);
nand UO_326 (O_326,N_19943,N_19961);
and UO_327 (O_327,N_19925,N_19897);
nand UO_328 (O_328,N_19943,N_19952);
and UO_329 (O_329,N_19823,N_19755);
nor UO_330 (O_330,N_19978,N_19957);
nand UO_331 (O_331,N_19971,N_19850);
xor UO_332 (O_332,N_19925,N_19898);
and UO_333 (O_333,N_19946,N_19952);
and UO_334 (O_334,N_19951,N_19956);
nor UO_335 (O_335,N_19839,N_19885);
nand UO_336 (O_336,N_19946,N_19813);
nor UO_337 (O_337,N_19924,N_19802);
and UO_338 (O_338,N_19782,N_19980);
nand UO_339 (O_339,N_19912,N_19768);
xor UO_340 (O_340,N_19810,N_19816);
xor UO_341 (O_341,N_19773,N_19874);
nand UO_342 (O_342,N_19828,N_19808);
xor UO_343 (O_343,N_19895,N_19755);
or UO_344 (O_344,N_19827,N_19776);
xnor UO_345 (O_345,N_19775,N_19773);
nand UO_346 (O_346,N_19972,N_19888);
and UO_347 (O_347,N_19988,N_19931);
nand UO_348 (O_348,N_19930,N_19873);
and UO_349 (O_349,N_19841,N_19847);
and UO_350 (O_350,N_19906,N_19931);
nor UO_351 (O_351,N_19815,N_19856);
nand UO_352 (O_352,N_19773,N_19818);
nor UO_353 (O_353,N_19852,N_19961);
and UO_354 (O_354,N_19962,N_19848);
nand UO_355 (O_355,N_19990,N_19852);
xnor UO_356 (O_356,N_19995,N_19773);
or UO_357 (O_357,N_19891,N_19829);
nand UO_358 (O_358,N_19977,N_19812);
or UO_359 (O_359,N_19947,N_19928);
or UO_360 (O_360,N_19876,N_19986);
xor UO_361 (O_361,N_19915,N_19875);
nor UO_362 (O_362,N_19915,N_19991);
or UO_363 (O_363,N_19831,N_19977);
xor UO_364 (O_364,N_19770,N_19932);
and UO_365 (O_365,N_19866,N_19758);
or UO_366 (O_366,N_19843,N_19757);
xor UO_367 (O_367,N_19836,N_19945);
or UO_368 (O_368,N_19829,N_19922);
or UO_369 (O_369,N_19967,N_19985);
or UO_370 (O_370,N_19827,N_19900);
xnor UO_371 (O_371,N_19938,N_19791);
nand UO_372 (O_372,N_19877,N_19805);
xor UO_373 (O_373,N_19888,N_19784);
or UO_374 (O_374,N_19904,N_19954);
or UO_375 (O_375,N_19826,N_19915);
xnor UO_376 (O_376,N_19906,N_19947);
nor UO_377 (O_377,N_19919,N_19766);
nor UO_378 (O_378,N_19807,N_19796);
or UO_379 (O_379,N_19772,N_19815);
or UO_380 (O_380,N_19782,N_19926);
or UO_381 (O_381,N_19800,N_19918);
nand UO_382 (O_382,N_19830,N_19750);
or UO_383 (O_383,N_19775,N_19938);
or UO_384 (O_384,N_19985,N_19774);
nand UO_385 (O_385,N_19908,N_19919);
xor UO_386 (O_386,N_19869,N_19985);
nand UO_387 (O_387,N_19792,N_19779);
nor UO_388 (O_388,N_19865,N_19811);
or UO_389 (O_389,N_19943,N_19975);
or UO_390 (O_390,N_19849,N_19777);
xor UO_391 (O_391,N_19854,N_19815);
and UO_392 (O_392,N_19900,N_19934);
xor UO_393 (O_393,N_19908,N_19810);
nand UO_394 (O_394,N_19828,N_19945);
nor UO_395 (O_395,N_19804,N_19807);
or UO_396 (O_396,N_19870,N_19923);
nand UO_397 (O_397,N_19995,N_19771);
and UO_398 (O_398,N_19809,N_19816);
nor UO_399 (O_399,N_19785,N_19881);
xor UO_400 (O_400,N_19992,N_19980);
nand UO_401 (O_401,N_19958,N_19992);
or UO_402 (O_402,N_19853,N_19930);
and UO_403 (O_403,N_19837,N_19973);
nor UO_404 (O_404,N_19886,N_19923);
nand UO_405 (O_405,N_19872,N_19897);
nor UO_406 (O_406,N_19877,N_19862);
nand UO_407 (O_407,N_19832,N_19940);
or UO_408 (O_408,N_19795,N_19872);
nand UO_409 (O_409,N_19777,N_19790);
nand UO_410 (O_410,N_19888,N_19995);
or UO_411 (O_411,N_19791,N_19819);
nand UO_412 (O_412,N_19988,N_19852);
nor UO_413 (O_413,N_19844,N_19969);
xor UO_414 (O_414,N_19870,N_19816);
xnor UO_415 (O_415,N_19934,N_19875);
nor UO_416 (O_416,N_19866,N_19960);
xor UO_417 (O_417,N_19969,N_19934);
nor UO_418 (O_418,N_19835,N_19855);
or UO_419 (O_419,N_19826,N_19778);
and UO_420 (O_420,N_19831,N_19839);
nand UO_421 (O_421,N_19998,N_19905);
xor UO_422 (O_422,N_19763,N_19766);
nor UO_423 (O_423,N_19944,N_19958);
and UO_424 (O_424,N_19875,N_19922);
xnor UO_425 (O_425,N_19936,N_19870);
or UO_426 (O_426,N_19941,N_19923);
and UO_427 (O_427,N_19903,N_19905);
nand UO_428 (O_428,N_19767,N_19785);
nor UO_429 (O_429,N_19803,N_19990);
nor UO_430 (O_430,N_19913,N_19768);
and UO_431 (O_431,N_19906,N_19975);
nand UO_432 (O_432,N_19757,N_19762);
and UO_433 (O_433,N_19817,N_19896);
nand UO_434 (O_434,N_19849,N_19933);
nand UO_435 (O_435,N_19994,N_19838);
or UO_436 (O_436,N_19786,N_19773);
or UO_437 (O_437,N_19789,N_19929);
and UO_438 (O_438,N_19910,N_19956);
nor UO_439 (O_439,N_19802,N_19976);
xor UO_440 (O_440,N_19758,N_19902);
xnor UO_441 (O_441,N_19996,N_19791);
nand UO_442 (O_442,N_19952,N_19756);
or UO_443 (O_443,N_19843,N_19923);
xor UO_444 (O_444,N_19934,N_19932);
xnor UO_445 (O_445,N_19822,N_19997);
and UO_446 (O_446,N_19989,N_19792);
or UO_447 (O_447,N_19772,N_19836);
and UO_448 (O_448,N_19878,N_19951);
nand UO_449 (O_449,N_19903,N_19787);
nand UO_450 (O_450,N_19871,N_19846);
nor UO_451 (O_451,N_19860,N_19773);
and UO_452 (O_452,N_19820,N_19854);
and UO_453 (O_453,N_19794,N_19760);
nand UO_454 (O_454,N_19999,N_19967);
xor UO_455 (O_455,N_19752,N_19750);
or UO_456 (O_456,N_19793,N_19945);
or UO_457 (O_457,N_19816,N_19944);
nor UO_458 (O_458,N_19972,N_19957);
xor UO_459 (O_459,N_19762,N_19994);
or UO_460 (O_460,N_19920,N_19831);
or UO_461 (O_461,N_19806,N_19914);
nor UO_462 (O_462,N_19838,N_19871);
and UO_463 (O_463,N_19915,N_19769);
or UO_464 (O_464,N_19855,N_19766);
nand UO_465 (O_465,N_19971,N_19900);
or UO_466 (O_466,N_19821,N_19991);
and UO_467 (O_467,N_19922,N_19971);
nor UO_468 (O_468,N_19899,N_19875);
or UO_469 (O_469,N_19995,N_19955);
nor UO_470 (O_470,N_19873,N_19848);
or UO_471 (O_471,N_19807,N_19988);
and UO_472 (O_472,N_19998,N_19826);
nor UO_473 (O_473,N_19869,N_19936);
nor UO_474 (O_474,N_19811,N_19780);
nand UO_475 (O_475,N_19955,N_19755);
or UO_476 (O_476,N_19807,N_19923);
xor UO_477 (O_477,N_19809,N_19932);
xnor UO_478 (O_478,N_19943,N_19840);
and UO_479 (O_479,N_19894,N_19835);
or UO_480 (O_480,N_19983,N_19864);
or UO_481 (O_481,N_19864,N_19923);
or UO_482 (O_482,N_19800,N_19820);
nand UO_483 (O_483,N_19860,N_19867);
or UO_484 (O_484,N_19866,N_19985);
and UO_485 (O_485,N_19799,N_19754);
or UO_486 (O_486,N_19931,N_19966);
and UO_487 (O_487,N_19859,N_19774);
and UO_488 (O_488,N_19931,N_19893);
or UO_489 (O_489,N_19938,N_19831);
nor UO_490 (O_490,N_19846,N_19999);
or UO_491 (O_491,N_19993,N_19909);
xor UO_492 (O_492,N_19771,N_19931);
nand UO_493 (O_493,N_19869,N_19884);
xor UO_494 (O_494,N_19994,N_19829);
nand UO_495 (O_495,N_19972,N_19992);
and UO_496 (O_496,N_19817,N_19810);
xnor UO_497 (O_497,N_19900,N_19989);
nand UO_498 (O_498,N_19875,N_19860);
nand UO_499 (O_499,N_19962,N_19777);
xnor UO_500 (O_500,N_19779,N_19795);
or UO_501 (O_501,N_19779,N_19927);
nor UO_502 (O_502,N_19785,N_19952);
nand UO_503 (O_503,N_19887,N_19761);
or UO_504 (O_504,N_19926,N_19865);
xor UO_505 (O_505,N_19946,N_19874);
nor UO_506 (O_506,N_19756,N_19766);
xnor UO_507 (O_507,N_19990,N_19930);
or UO_508 (O_508,N_19854,N_19964);
and UO_509 (O_509,N_19772,N_19934);
nand UO_510 (O_510,N_19798,N_19923);
nand UO_511 (O_511,N_19945,N_19990);
nor UO_512 (O_512,N_19881,N_19874);
nand UO_513 (O_513,N_19782,N_19890);
or UO_514 (O_514,N_19935,N_19952);
nand UO_515 (O_515,N_19875,N_19928);
nor UO_516 (O_516,N_19796,N_19874);
xor UO_517 (O_517,N_19765,N_19789);
or UO_518 (O_518,N_19789,N_19940);
or UO_519 (O_519,N_19769,N_19825);
nor UO_520 (O_520,N_19937,N_19794);
nor UO_521 (O_521,N_19845,N_19847);
nor UO_522 (O_522,N_19950,N_19956);
nor UO_523 (O_523,N_19851,N_19777);
nor UO_524 (O_524,N_19866,N_19858);
or UO_525 (O_525,N_19871,N_19886);
nor UO_526 (O_526,N_19769,N_19857);
or UO_527 (O_527,N_19812,N_19939);
xor UO_528 (O_528,N_19817,N_19989);
nor UO_529 (O_529,N_19874,N_19992);
or UO_530 (O_530,N_19912,N_19927);
nor UO_531 (O_531,N_19911,N_19796);
nand UO_532 (O_532,N_19836,N_19815);
xor UO_533 (O_533,N_19890,N_19962);
or UO_534 (O_534,N_19843,N_19767);
nor UO_535 (O_535,N_19788,N_19919);
and UO_536 (O_536,N_19941,N_19755);
and UO_537 (O_537,N_19982,N_19969);
or UO_538 (O_538,N_19866,N_19823);
and UO_539 (O_539,N_19872,N_19891);
or UO_540 (O_540,N_19756,N_19964);
xnor UO_541 (O_541,N_19847,N_19792);
nor UO_542 (O_542,N_19906,N_19918);
or UO_543 (O_543,N_19781,N_19774);
nand UO_544 (O_544,N_19762,N_19776);
xor UO_545 (O_545,N_19804,N_19893);
and UO_546 (O_546,N_19811,N_19834);
xor UO_547 (O_547,N_19954,N_19935);
nand UO_548 (O_548,N_19961,N_19798);
nor UO_549 (O_549,N_19804,N_19829);
xnor UO_550 (O_550,N_19833,N_19875);
xor UO_551 (O_551,N_19990,N_19941);
or UO_552 (O_552,N_19926,N_19909);
nand UO_553 (O_553,N_19968,N_19990);
nand UO_554 (O_554,N_19949,N_19783);
and UO_555 (O_555,N_19856,N_19891);
nand UO_556 (O_556,N_19803,N_19878);
and UO_557 (O_557,N_19945,N_19871);
nor UO_558 (O_558,N_19774,N_19770);
or UO_559 (O_559,N_19948,N_19959);
or UO_560 (O_560,N_19877,N_19885);
nor UO_561 (O_561,N_19793,N_19858);
or UO_562 (O_562,N_19783,N_19876);
and UO_563 (O_563,N_19864,N_19920);
or UO_564 (O_564,N_19864,N_19890);
and UO_565 (O_565,N_19856,N_19967);
or UO_566 (O_566,N_19849,N_19994);
or UO_567 (O_567,N_19763,N_19995);
or UO_568 (O_568,N_19914,N_19994);
nand UO_569 (O_569,N_19831,N_19836);
nor UO_570 (O_570,N_19872,N_19999);
xnor UO_571 (O_571,N_19952,N_19902);
nand UO_572 (O_572,N_19805,N_19771);
or UO_573 (O_573,N_19884,N_19943);
xor UO_574 (O_574,N_19989,N_19832);
xor UO_575 (O_575,N_19830,N_19906);
xnor UO_576 (O_576,N_19994,N_19778);
nor UO_577 (O_577,N_19846,N_19981);
or UO_578 (O_578,N_19892,N_19944);
and UO_579 (O_579,N_19774,N_19787);
nor UO_580 (O_580,N_19998,N_19939);
nor UO_581 (O_581,N_19812,N_19750);
xnor UO_582 (O_582,N_19880,N_19785);
xor UO_583 (O_583,N_19800,N_19935);
and UO_584 (O_584,N_19770,N_19861);
and UO_585 (O_585,N_19822,N_19836);
and UO_586 (O_586,N_19971,N_19787);
or UO_587 (O_587,N_19842,N_19756);
nand UO_588 (O_588,N_19847,N_19996);
nor UO_589 (O_589,N_19962,N_19904);
or UO_590 (O_590,N_19993,N_19921);
and UO_591 (O_591,N_19905,N_19912);
nand UO_592 (O_592,N_19929,N_19958);
and UO_593 (O_593,N_19849,N_19823);
and UO_594 (O_594,N_19802,N_19939);
or UO_595 (O_595,N_19949,N_19997);
xnor UO_596 (O_596,N_19866,N_19912);
nor UO_597 (O_597,N_19910,N_19855);
or UO_598 (O_598,N_19811,N_19863);
and UO_599 (O_599,N_19876,N_19959);
or UO_600 (O_600,N_19804,N_19976);
nand UO_601 (O_601,N_19932,N_19930);
or UO_602 (O_602,N_19860,N_19963);
nand UO_603 (O_603,N_19771,N_19946);
nand UO_604 (O_604,N_19981,N_19795);
and UO_605 (O_605,N_19818,N_19917);
nand UO_606 (O_606,N_19815,N_19803);
nand UO_607 (O_607,N_19932,N_19759);
xnor UO_608 (O_608,N_19904,N_19767);
and UO_609 (O_609,N_19888,N_19906);
nor UO_610 (O_610,N_19906,N_19894);
or UO_611 (O_611,N_19769,N_19884);
nor UO_612 (O_612,N_19897,N_19952);
or UO_613 (O_613,N_19833,N_19798);
and UO_614 (O_614,N_19896,N_19991);
or UO_615 (O_615,N_19956,N_19850);
nand UO_616 (O_616,N_19918,N_19837);
or UO_617 (O_617,N_19943,N_19902);
and UO_618 (O_618,N_19797,N_19948);
or UO_619 (O_619,N_19986,N_19787);
or UO_620 (O_620,N_19784,N_19950);
and UO_621 (O_621,N_19902,N_19854);
nand UO_622 (O_622,N_19906,N_19948);
or UO_623 (O_623,N_19951,N_19984);
or UO_624 (O_624,N_19875,N_19930);
xnor UO_625 (O_625,N_19957,N_19983);
and UO_626 (O_626,N_19880,N_19904);
xnor UO_627 (O_627,N_19861,N_19751);
xnor UO_628 (O_628,N_19799,N_19881);
or UO_629 (O_629,N_19882,N_19938);
nand UO_630 (O_630,N_19975,N_19969);
xnor UO_631 (O_631,N_19791,N_19836);
xnor UO_632 (O_632,N_19823,N_19987);
and UO_633 (O_633,N_19824,N_19795);
and UO_634 (O_634,N_19881,N_19944);
nor UO_635 (O_635,N_19794,N_19948);
or UO_636 (O_636,N_19982,N_19948);
xor UO_637 (O_637,N_19907,N_19891);
or UO_638 (O_638,N_19891,N_19761);
or UO_639 (O_639,N_19992,N_19934);
nor UO_640 (O_640,N_19905,N_19770);
nand UO_641 (O_641,N_19993,N_19771);
xnor UO_642 (O_642,N_19946,N_19758);
and UO_643 (O_643,N_19995,N_19825);
nand UO_644 (O_644,N_19928,N_19846);
xor UO_645 (O_645,N_19939,N_19764);
xnor UO_646 (O_646,N_19839,N_19842);
xnor UO_647 (O_647,N_19951,N_19958);
xnor UO_648 (O_648,N_19974,N_19833);
nand UO_649 (O_649,N_19886,N_19966);
nor UO_650 (O_650,N_19920,N_19957);
or UO_651 (O_651,N_19762,N_19900);
nand UO_652 (O_652,N_19809,N_19970);
xnor UO_653 (O_653,N_19783,N_19899);
nand UO_654 (O_654,N_19933,N_19938);
nand UO_655 (O_655,N_19940,N_19793);
or UO_656 (O_656,N_19998,N_19887);
nand UO_657 (O_657,N_19901,N_19806);
and UO_658 (O_658,N_19843,N_19782);
and UO_659 (O_659,N_19774,N_19906);
or UO_660 (O_660,N_19909,N_19814);
nor UO_661 (O_661,N_19925,N_19991);
xor UO_662 (O_662,N_19772,N_19966);
and UO_663 (O_663,N_19927,N_19967);
or UO_664 (O_664,N_19835,N_19926);
and UO_665 (O_665,N_19882,N_19781);
and UO_666 (O_666,N_19903,N_19785);
nor UO_667 (O_667,N_19874,N_19999);
nor UO_668 (O_668,N_19771,N_19852);
xnor UO_669 (O_669,N_19854,N_19800);
and UO_670 (O_670,N_19778,N_19832);
or UO_671 (O_671,N_19924,N_19908);
or UO_672 (O_672,N_19803,N_19805);
or UO_673 (O_673,N_19806,N_19832);
xnor UO_674 (O_674,N_19940,N_19851);
nor UO_675 (O_675,N_19826,N_19863);
or UO_676 (O_676,N_19926,N_19919);
nand UO_677 (O_677,N_19942,N_19973);
xor UO_678 (O_678,N_19909,N_19903);
xor UO_679 (O_679,N_19829,N_19984);
or UO_680 (O_680,N_19764,N_19811);
and UO_681 (O_681,N_19929,N_19763);
and UO_682 (O_682,N_19783,N_19959);
and UO_683 (O_683,N_19856,N_19823);
xnor UO_684 (O_684,N_19813,N_19822);
xnor UO_685 (O_685,N_19833,N_19895);
or UO_686 (O_686,N_19819,N_19781);
nand UO_687 (O_687,N_19855,N_19797);
or UO_688 (O_688,N_19910,N_19803);
xor UO_689 (O_689,N_19869,N_19787);
nand UO_690 (O_690,N_19778,N_19943);
nand UO_691 (O_691,N_19836,N_19800);
or UO_692 (O_692,N_19896,N_19971);
and UO_693 (O_693,N_19814,N_19766);
nand UO_694 (O_694,N_19950,N_19998);
or UO_695 (O_695,N_19890,N_19851);
or UO_696 (O_696,N_19923,N_19948);
xor UO_697 (O_697,N_19834,N_19750);
nand UO_698 (O_698,N_19797,N_19844);
nor UO_699 (O_699,N_19778,N_19813);
nand UO_700 (O_700,N_19911,N_19907);
nand UO_701 (O_701,N_19786,N_19838);
nor UO_702 (O_702,N_19828,N_19907);
or UO_703 (O_703,N_19783,N_19790);
xnor UO_704 (O_704,N_19923,N_19767);
xor UO_705 (O_705,N_19917,N_19924);
nor UO_706 (O_706,N_19968,N_19917);
and UO_707 (O_707,N_19962,N_19920);
xor UO_708 (O_708,N_19985,N_19851);
nor UO_709 (O_709,N_19912,N_19807);
or UO_710 (O_710,N_19772,N_19776);
and UO_711 (O_711,N_19763,N_19858);
or UO_712 (O_712,N_19973,N_19936);
and UO_713 (O_713,N_19885,N_19938);
or UO_714 (O_714,N_19909,N_19774);
nand UO_715 (O_715,N_19874,N_19844);
or UO_716 (O_716,N_19967,N_19759);
xnor UO_717 (O_717,N_19896,N_19794);
or UO_718 (O_718,N_19846,N_19828);
nand UO_719 (O_719,N_19876,N_19974);
xor UO_720 (O_720,N_19990,N_19837);
nor UO_721 (O_721,N_19999,N_19849);
xnor UO_722 (O_722,N_19766,N_19782);
nor UO_723 (O_723,N_19971,N_19879);
nor UO_724 (O_724,N_19803,N_19811);
nand UO_725 (O_725,N_19835,N_19960);
nor UO_726 (O_726,N_19950,N_19984);
xnor UO_727 (O_727,N_19961,N_19833);
xor UO_728 (O_728,N_19841,N_19812);
nand UO_729 (O_729,N_19930,N_19753);
nand UO_730 (O_730,N_19950,N_19878);
and UO_731 (O_731,N_19896,N_19803);
nor UO_732 (O_732,N_19879,N_19797);
and UO_733 (O_733,N_19809,N_19845);
or UO_734 (O_734,N_19952,N_19998);
nand UO_735 (O_735,N_19818,N_19812);
or UO_736 (O_736,N_19889,N_19857);
or UO_737 (O_737,N_19981,N_19797);
and UO_738 (O_738,N_19818,N_19950);
xor UO_739 (O_739,N_19823,N_19861);
xor UO_740 (O_740,N_19771,N_19903);
nor UO_741 (O_741,N_19754,N_19818);
nand UO_742 (O_742,N_19761,N_19879);
or UO_743 (O_743,N_19997,N_19837);
and UO_744 (O_744,N_19894,N_19922);
xor UO_745 (O_745,N_19798,N_19801);
nand UO_746 (O_746,N_19906,N_19757);
nand UO_747 (O_747,N_19968,N_19798);
or UO_748 (O_748,N_19899,N_19785);
nor UO_749 (O_749,N_19759,N_19965);
nand UO_750 (O_750,N_19943,N_19926);
xor UO_751 (O_751,N_19814,N_19954);
xnor UO_752 (O_752,N_19954,N_19879);
xnor UO_753 (O_753,N_19781,N_19975);
nand UO_754 (O_754,N_19816,N_19751);
or UO_755 (O_755,N_19968,N_19959);
and UO_756 (O_756,N_19863,N_19874);
nand UO_757 (O_757,N_19888,N_19983);
or UO_758 (O_758,N_19833,N_19926);
xor UO_759 (O_759,N_19891,N_19979);
or UO_760 (O_760,N_19867,N_19807);
nor UO_761 (O_761,N_19867,N_19998);
nand UO_762 (O_762,N_19913,N_19818);
nor UO_763 (O_763,N_19965,N_19853);
and UO_764 (O_764,N_19756,N_19823);
and UO_765 (O_765,N_19868,N_19785);
nor UO_766 (O_766,N_19767,N_19928);
xnor UO_767 (O_767,N_19828,N_19909);
nor UO_768 (O_768,N_19866,N_19899);
nor UO_769 (O_769,N_19968,N_19778);
and UO_770 (O_770,N_19750,N_19877);
nand UO_771 (O_771,N_19775,N_19751);
nand UO_772 (O_772,N_19846,N_19877);
or UO_773 (O_773,N_19901,N_19790);
xnor UO_774 (O_774,N_19814,N_19963);
nor UO_775 (O_775,N_19887,N_19889);
and UO_776 (O_776,N_19795,N_19980);
xnor UO_777 (O_777,N_19956,N_19840);
nand UO_778 (O_778,N_19803,N_19797);
nor UO_779 (O_779,N_19752,N_19894);
or UO_780 (O_780,N_19969,N_19799);
nand UO_781 (O_781,N_19998,N_19961);
nor UO_782 (O_782,N_19971,N_19756);
nor UO_783 (O_783,N_19817,N_19979);
or UO_784 (O_784,N_19750,N_19937);
or UO_785 (O_785,N_19940,N_19952);
xor UO_786 (O_786,N_19933,N_19819);
xor UO_787 (O_787,N_19888,N_19827);
nand UO_788 (O_788,N_19801,N_19877);
nand UO_789 (O_789,N_19968,N_19989);
or UO_790 (O_790,N_19939,N_19832);
nor UO_791 (O_791,N_19818,N_19868);
or UO_792 (O_792,N_19870,N_19987);
or UO_793 (O_793,N_19878,N_19885);
or UO_794 (O_794,N_19896,N_19934);
and UO_795 (O_795,N_19972,N_19781);
or UO_796 (O_796,N_19763,N_19944);
and UO_797 (O_797,N_19931,N_19925);
nor UO_798 (O_798,N_19949,N_19928);
nor UO_799 (O_799,N_19966,N_19891);
nand UO_800 (O_800,N_19908,N_19824);
nand UO_801 (O_801,N_19753,N_19931);
xnor UO_802 (O_802,N_19901,N_19755);
nor UO_803 (O_803,N_19855,N_19889);
xor UO_804 (O_804,N_19933,N_19833);
nand UO_805 (O_805,N_19862,N_19829);
nand UO_806 (O_806,N_19777,N_19963);
or UO_807 (O_807,N_19797,N_19977);
xnor UO_808 (O_808,N_19766,N_19764);
xor UO_809 (O_809,N_19894,N_19756);
xnor UO_810 (O_810,N_19759,N_19883);
xor UO_811 (O_811,N_19991,N_19777);
and UO_812 (O_812,N_19815,N_19830);
or UO_813 (O_813,N_19903,N_19915);
nor UO_814 (O_814,N_19827,N_19839);
xnor UO_815 (O_815,N_19956,N_19932);
nor UO_816 (O_816,N_19750,N_19773);
and UO_817 (O_817,N_19925,N_19905);
or UO_818 (O_818,N_19832,N_19777);
nand UO_819 (O_819,N_19821,N_19797);
nor UO_820 (O_820,N_19856,N_19871);
nand UO_821 (O_821,N_19776,N_19963);
nor UO_822 (O_822,N_19854,N_19822);
or UO_823 (O_823,N_19948,N_19886);
nor UO_824 (O_824,N_19920,N_19964);
nand UO_825 (O_825,N_19955,N_19784);
nand UO_826 (O_826,N_19968,N_19997);
nor UO_827 (O_827,N_19807,N_19765);
nor UO_828 (O_828,N_19965,N_19813);
xor UO_829 (O_829,N_19909,N_19977);
xor UO_830 (O_830,N_19929,N_19884);
and UO_831 (O_831,N_19822,N_19844);
xor UO_832 (O_832,N_19927,N_19889);
nand UO_833 (O_833,N_19969,N_19762);
xor UO_834 (O_834,N_19851,N_19753);
nand UO_835 (O_835,N_19943,N_19971);
and UO_836 (O_836,N_19898,N_19965);
xnor UO_837 (O_837,N_19863,N_19944);
nand UO_838 (O_838,N_19814,N_19820);
or UO_839 (O_839,N_19814,N_19876);
and UO_840 (O_840,N_19974,N_19866);
or UO_841 (O_841,N_19860,N_19971);
nand UO_842 (O_842,N_19993,N_19828);
or UO_843 (O_843,N_19902,N_19944);
or UO_844 (O_844,N_19873,N_19858);
and UO_845 (O_845,N_19880,N_19826);
xnor UO_846 (O_846,N_19943,N_19955);
nor UO_847 (O_847,N_19969,N_19852);
nand UO_848 (O_848,N_19985,N_19830);
or UO_849 (O_849,N_19805,N_19931);
or UO_850 (O_850,N_19800,N_19971);
xor UO_851 (O_851,N_19791,N_19782);
nor UO_852 (O_852,N_19921,N_19821);
nor UO_853 (O_853,N_19830,N_19873);
or UO_854 (O_854,N_19878,N_19965);
xor UO_855 (O_855,N_19919,N_19922);
xor UO_856 (O_856,N_19772,N_19771);
xor UO_857 (O_857,N_19973,N_19855);
nor UO_858 (O_858,N_19804,N_19878);
and UO_859 (O_859,N_19978,N_19812);
and UO_860 (O_860,N_19977,N_19902);
xnor UO_861 (O_861,N_19933,N_19883);
nand UO_862 (O_862,N_19875,N_19812);
nand UO_863 (O_863,N_19888,N_19866);
nand UO_864 (O_864,N_19869,N_19785);
and UO_865 (O_865,N_19943,N_19846);
nand UO_866 (O_866,N_19888,N_19849);
or UO_867 (O_867,N_19898,N_19846);
and UO_868 (O_868,N_19956,N_19896);
xnor UO_869 (O_869,N_19989,N_19927);
and UO_870 (O_870,N_19891,N_19967);
and UO_871 (O_871,N_19963,N_19978);
nor UO_872 (O_872,N_19974,N_19803);
nor UO_873 (O_873,N_19791,N_19897);
nand UO_874 (O_874,N_19892,N_19757);
nor UO_875 (O_875,N_19798,N_19839);
and UO_876 (O_876,N_19758,N_19954);
nand UO_877 (O_877,N_19961,N_19854);
nand UO_878 (O_878,N_19837,N_19760);
nand UO_879 (O_879,N_19804,N_19832);
nor UO_880 (O_880,N_19936,N_19808);
and UO_881 (O_881,N_19763,N_19821);
xnor UO_882 (O_882,N_19917,N_19832);
and UO_883 (O_883,N_19837,N_19978);
nor UO_884 (O_884,N_19951,N_19962);
or UO_885 (O_885,N_19863,N_19912);
or UO_886 (O_886,N_19802,N_19998);
xnor UO_887 (O_887,N_19977,N_19945);
or UO_888 (O_888,N_19790,N_19811);
or UO_889 (O_889,N_19995,N_19916);
or UO_890 (O_890,N_19843,N_19829);
nor UO_891 (O_891,N_19760,N_19850);
or UO_892 (O_892,N_19907,N_19815);
nor UO_893 (O_893,N_19888,N_19752);
nand UO_894 (O_894,N_19820,N_19891);
and UO_895 (O_895,N_19929,N_19886);
or UO_896 (O_896,N_19964,N_19987);
and UO_897 (O_897,N_19916,N_19780);
or UO_898 (O_898,N_19766,N_19977);
or UO_899 (O_899,N_19794,N_19976);
nor UO_900 (O_900,N_19827,N_19757);
xnor UO_901 (O_901,N_19751,N_19938);
or UO_902 (O_902,N_19931,N_19990);
nor UO_903 (O_903,N_19818,N_19929);
xnor UO_904 (O_904,N_19797,N_19830);
and UO_905 (O_905,N_19839,N_19978);
xor UO_906 (O_906,N_19999,N_19814);
nor UO_907 (O_907,N_19834,N_19755);
or UO_908 (O_908,N_19846,N_19880);
nand UO_909 (O_909,N_19838,N_19858);
nor UO_910 (O_910,N_19918,N_19878);
xnor UO_911 (O_911,N_19861,N_19931);
or UO_912 (O_912,N_19757,N_19816);
or UO_913 (O_913,N_19873,N_19905);
nand UO_914 (O_914,N_19820,N_19751);
xnor UO_915 (O_915,N_19844,N_19769);
nand UO_916 (O_916,N_19850,N_19801);
and UO_917 (O_917,N_19797,N_19753);
and UO_918 (O_918,N_19908,N_19831);
xor UO_919 (O_919,N_19967,N_19768);
nand UO_920 (O_920,N_19922,N_19904);
xor UO_921 (O_921,N_19803,N_19887);
xor UO_922 (O_922,N_19971,N_19827);
or UO_923 (O_923,N_19874,N_19864);
or UO_924 (O_924,N_19929,N_19872);
nand UO_925 (O_925,N_19824,N_19869);
or UO_926 (O_926,N_19901,N_19866);
and UO_927 (O_927,N_19815,N_19821);
xor UO_928 (O_928,N_19973,N_19920);
and UO_929 (O_929,N_19842,N_19790);
and UO_930 (O_930,N_19906,N_19773);
or UO_931 (O_931,N_19826,N_19799);
xnor UO_932 (O_932,N_19840,N_19765);
nand UO_933 (O_933,N_19960,N_19900);
and UO_934 (O_934,N_19883,N_19774);
nand UO_935 (O_935,N_19757,N_19819);
and UO_936 (O_936,N_19904,N_19836);
nand UO_937 (O_937,N_19778,N_19850);
and UO_938 (O_938,N_19762,N_19806);
and UO_939 (O_939,N_19836,N_19771);
xor UO_940 (O_940,N_19968,N_19982);
xor UO_941 (O_941,N_19925,N_19874);
xnor UO_942 (O_942,N_19760,N_19826);
or UO_943 (O_943,N_19754,N_19907);
nand UO_944 (O_944,N_19881,N_19884);
nand UO_945 (O_945,N_19859,N_19773);
xor UO_946 (O_946,N_19773,N_19865);
xnor UO_947 (O_947,N_19973,N_19875);
and UO_948 (O_948,N_19951,N_19837);
xor UO_949 (O_949,N_19969,N_19893);
and UO_950 (O_950,N_19768,N_19943);
nand UO_951 (O_951,N_19935,N_19815);
and UO_952 (O_952,N_19876,N_19906);
and UO_953 (O_953,N_19970,N_19786);
nand UO_954 (O_954,N_19978,N_19778);
nor UO_955 (O_955,N_19929,N_19855);
xnor UO_956 (O_956,N_19936,N_19961);
nand UO_957 (O_957,N_19923,N_19966);
or UO_958 (O_958,N_19764,N_19918);
and UO_959 (O_959,N_19963,N_19781);
and UO_960 (O_960,N_19947,N_19945);
and UO_961 (O_961,N_19952,N_19927);
nor UO_962 (O_962,N_19839,N_19872);
or UO_963 (O_963,N_19923,N_19889);
nand UO_964 (O_964,N_19938,N_19796);
and UO_965 (O_965,N_19775,N_19861);
xor UO_966 (O_966,N_19990,N_19850);
xor UO_967 (O_967,N_19869,N_19865);
or UO_968 (O_968,N_19753,N_19782);
or UO_969 (O_969,N_19866,N_19814);
nand UO_970 (O_970,N_19972,N_19911);
and UO_971 (O_971,N_19990,N_19765);
nor UO_972 (O_972,N_19768,N_19992);
nand UO_973 (O_973,N_19787,N_19778);
nor UO_974 (O_974,N_19992,N_19810);
and UO_975 (O_975,N_19956,N_19954);
nand UO_976 (O_976,N_19934,N_19881);
xor UO_977 (O_977,N_19995,N_19892);
nand UO_978 (O_978,N_19762,N_19804);
nand UO_979 (O_979,N_19842,N_19789);
or UO_980 (O_980,N_19859,N_19807);
nand UO_981 (O_981,N_19825,N_19755);
and UO_982 (O_982,N_19956,N_19945);
xnor UO_983 (O_983,N_19880,N_19761);
nor UO_984 (O_984,N_19809,N_19918);
or UO_985 (O_985,N_19836,N_19781);
or UO_986 (O_986,N_19975,N_19984);
nand UO_987 (O_987,N_19846,N_19978);
xor UO_988 (O_988,N_19923,N_19949);
nor UO_989 (O_989,N_19852,N_19986);
and UO_990 (O_990,N_19886,N_19785);
and UO_991 (O_991,N_19790,N_19830);
and UO_992 (O_992,N_19957,N_19951);
nand UO_993 (O_993,N_19965,N_19838);
nor UO_994 (O_994,N_19844,N_19973);
and UO_995 (O_995,N_19801,N_19895);
nand UO_996 (O_996,N_19871,N_19916);
or UO_997 (O_997,N_19759,N_19959);
nor UO_998 (O_998,N_19926,N_19765);
or UO_999 (O_999,N_19898,N_19869);
or UO_1000 (O_1000,N_19780,N_19866);
nand UO_1001 (O_1001,N_19857,N_19774);
nand UO_1002 (O_1002,N_19948,N_19965);
nand UO_1003 (O_1003,N_19968,N_19921);
and UO_1004 (O_1004,N_19896,N_19970);
or UO_1005 (O_1005,N_19912,N_19808);
and UO_1006 (O_1006,N_19807,N_19945);
nand UO_1007 (O_1007,N_19950,N_19776);
and UO_1008 (O_1008,N_19893,N_19947);
xor UO_1009 (O_1009,N_19868,N_19750);
nand UO_1010 (O_1010,N_19784,N_19870);
or UO_1011 (O_1011,N_19952,N_19969);
nand UO_1012 (O_1012,N_19950,N_19922);
and UO_1013 (O_1013,N_19910,N_19816);
nand UO_1014 (O_1014,N_19995,N_19782);
nand UO_1015 (O_1015,N_19790,N_19918);
nor UO_1016 (O_1016,N_19829,N_19905);
nor UO_1017 (O_1017,N_19776,N_19758);
nand UO_1018 (O_1018,N_19921,N_19978);
xor UO_1019 (O_1019,N_19801,N_19846);
or UO_1020 (O_1020,N_19951,N_19895);
xor UO_1021 (O_1021,N_19945,N_19887);
and UO_1022 (O_1022,N_19946,N_19823);
nand UO_1023 (O_1023,N_19959,N_19864);
or UO_1024 (O_1024,N_19934,N_19953);
and UO_1025 (O_1025,N_19891,N_19811);
or UO_1026 (O_1026,N_19939,N_19957);
nand UO_1027 (O_1027,N_19863,N_19800);
and UO_1028 (O_1028,N_19951,N_19800);
nand UO_1029 (O_1029,N_19964,N_19989);
xor UO_1030 (O_1030,N_19924,N_19984);
xnor UO_1031 (O_1031,N_19816,N_19891);
nand UO_1032 (O_1032,N_19997,N_19829);
or UO_1033 (O_1033,N_19966,N_19813);
nand UO_1034 (O_1034,N_19820,N_19771);
nand UO_1035 (O_1035,N_19966,N_19842);
or UO_1036 (O_1036,N_19856,N_19832);
nand UO_1037 (O_1037,N_19794,N_19904);
nand UO_1038 (O_1038,N_19992,N_19883);
or UO_1039 (O_1039,N_19765,N_19776);
or UO_1040 (O_1040,N_19872,N_19854);
and UO_1041 (O_1041,N_19966,N_19818);
or UO_1042 (O_1042,N_19832,N_19760);
or UO_1043 (O_1043,N_19851,N_19830);
and UO_1044 (O_1044,N_19829,N_19934);
xnor UO_1045 (O_1045,N_19765,N_19920);
nor UO_1046 (O_1046,N_19925,N_19902);
nand UO_1047 (O_1047,N_19838,N_19775);
and UO_1048 (O_1048,N_19850,N_19958);
nand UO_1049 (O_1049,N_19960,N_19966);
xor UO_1050 (O_1050,N_19964,N_19786);
nand UO_1051 (O_1051,N_19779,N_19891);
xnor UO_1052 (O_1052,N_19980,N_19898);
or UO_1053 (O_1053,N_19912,N_19776);
nor UO_1054 (O_1054,N_19750,N_19757);
xnor UO_1055 (O_1055,N_19842,N_19996);
nor UO_1056 (O_1056,N_19755,N_19865);
and UO_1057 (O_1057,N_19777,N_19874);
nor UO_1058 (O_1058,N_19856,N_19987);
xnor UO_1059 (O_1059,N_19803,N_19870);
and UO_1060 (O_1060,N_19750,N_19962);
nor UO_1061 (O_1061,N_19838,N_19788);
xnor UO_1062 (O_1062,N_19838,N_19851);
nor UO_1063 (O_1063,N_19883,N_19972);
nor UO_1064 (O_1064,N_19977,N_19778);
and UO_1065 (O_1065,N_19889,N_19879);
xnor UO_1066 (O_1066,N_19821,N_19776);
and UO_1067 (O_1067,N_19931,N_19758);
and UO_1068 (O_1068,N_19859,N_19864);
xor UO_1069 (O_1069,N_19890,N_19868);
nor UO_1070 (O_1070,N_19774,N_19856);
nand UO_1071 (O_1071,N_19803,N_19902);
xor UO_1072 (O_1072,N_19770,N_19915);
or UO_1073 (O_1073,N_19851,N_19839);
or UO_1074 (O_1074,N_19813,N_19829);
nor UO_1075 (O_1075,N_19801,N_19842);
or UO_1076 (O_1076,N_19751,N_19873);
or UO_1077 (O_1077,N_19806,N_19767);
nand UO_1078 (O_1078,N_19823,N_19976);
nor UO_1079 (O_1079,N_19765,N_19863);
or UO_1080 (O_1080,N_19755,N_19991);
and UO_1081 (O_1081,N_19762,N_19890);
or UO_1082 (O_1082,N_19961,N_19898);
nand UO_1083 (O_1083,N_19902,N_19767);
or UO_1084 (O_1084,N_19924,N_19976);
nor UO_1085 (O_1085,N_19846,N_19966);
nand UO_1086 (O_1086,N_19932,N_19813);
xor UO_1087 (O_1087,N_19896,N_19872);
nor UO_1088 (O_1088,N_19943,N_19939);
nand UO_1089 (O_1089,N_19944,N_19759);
nor UO_1090 (O_1090,N_19909,N_19818);
or UO_1091 (O_1091,N_19775,N_19899);
or UO_1092 (O_1092,N_19937,N_19921);
and UO_1093 (O_1093,N_19912,N_19760);
or UO_1094 (O_1094,N_19750,N_19793);
and UO_1095 (O_1095,N_19856,N_19818);
or UO_1096 (O_1096,N_19825,N_19910);
xnor UO_1097 (O_1097,N_19997,N_19787);
xnor UO_1098 (O_1098,N_19898,N_19779);
or UO_1099 (O_1099,N_19911,N_19991);
xnor UO_1100 (O_1100,N_19833,N_19762);
or UO_1101 (O_1101,N_19935,N_19803);
nand UO_1102 (O_1102,N_19755,N_19918);
and UO_1103 (O_1103,N_19936,N_19871);
nand UO_1104 (O_1104,N_19883,N_19908);
nand UO_1105 (O_1105,N_19941,N_19919);
nor UO_1106 (O_1106,N_19965,N_19910);
or UO_1107 (O_1107,N_19794,N_19856);
and UO_1108 (O_1108,N_19926,N_19894);
xor UO_1109 (O_1109,N_19860,N_19815);
xnor UO_1110 (O_1110,N_19832,N_19966);
xnor UO_1111 (O_1111,N_19813,N_19980);
or UO_1112 (O_1112,N_19776,N_19835);
and UO_1113 (O_1113,N_19762,N_19882);
nor UO_1114 (O_1114,N_19948,N_19824);
or UO_1115 (O_1115,N_19993,N_19998);
and UO_1116 (O_1116,N_19856,N_19977);
nor UO_1117 (O_1117,N_19861,N_19962);
xnor UO_1118 (O_1118,N_19852,N_19822);
nor UO_1119 (O_1119,N_19917,N_19962);
or UO_1120 (O_1120,N_19894,N_19837);
or UO_1121 (O_1121,N_19993,N_19808);
and UO_1122 (O_1122,N_19991,N_19758);
nand UO_1123 (O_1123,N_19875,N_19951);
nor UO_1124 (O_1124,N_19941,N_19901);
xnor UO_1125 (O_1125,N_19774,N_19756);
or UO_1126 (O_1126,N_19932,N_19946);
xor UO_1127 (O_1127,N_19798,N_19882);
or UO_1128 (O_1128,N_19891,N_19754);
and UO_1129 (O_1129,N_19804,N_19950);
nand UO_1130 (O_1130,N_19949,N_19973);
nor UO_1131 (O_1131,N_19774,N_19959);
or UO_1132 (O_1132,N_19875,N_19880);
and UO_1133 (O_1133,N_19928,N_19896);
nand UO_1134 (O_1134,N_19849,N_19955);
or UO_1135 (O_1135,N_19823,N_19876);
or UO_1136 (O_1136,N_19919,N_19977);
xor UO_1137 (O_1137,N_19956,N_19887);
and UO_1138 (O_1138,N_19963,N_19890);
nor UO_1139 (O_1139,N_19770,N_19840);
nand UO_1140 (O_1140,N_19752,N_19930);
xor UO_1141 (O_1141,N_19764,N_19845);
and UO_1142 (O_1142,N_19760,N_19823);
xnor UO_1143 (O_1143,N_19881,N_19762);
xnor UO_1144 (O_1144,N_19958,N_19976);
nand UO_1145 (O_1145,N_19927,N_19956);
nand UO_1146 (O_1146,N_19800,N_19808);
nor UO_1147 (O_1147,N_19753,N_19769);
nand UO_1148 (O_1148,N_19801,N_19879);
nand UO_1149 (O_1149,N_19751,N_19881);
or UO_1150 (O_1150,N_19953,N_19852);
or UO_1151 (O_1151,N_19918,N_19895);
xor UO_1152 (O_1152,N_19839,N_19925);
xnor UO_1153 (O_1153,N_19875,N_19883);
and UO_1154 (O_1154,N_19933,N_19783);
xor UO_1155 (O_1155,N_19929,N_19799);
nand UO_1156 (O_1156,N_19929,N_19777);
nor UO_1157 (O_1157,N_19776,N_19880);
and UO_1158 (O_1158,N_19970,N_19768);
nand UO_1159 (O_1159,N_19970,N_19905);
and UO_1160 (O_1160,N_19993,N_19835);
or UO_1161 (O_1161,N_19909,N_19812);
xor UO_1162 (O_1162,N_19789,N_19867);
xor UO_1163 (O_1163,N_19867,N_19955);
and UO_1164 (O_1164,N_19834,N_19962);
nand UO_1165 (O_1165,N_19873,N_19761);
or UO_1166 (O_1166,N_19946,N_19966);
nand UO_1167 (O_1167,N_19942,N_19857);
and UO_1168 (O_1168,N_19966,N_19861);
nor UO_1169 (O_1169,N_19921,N_19847);
nor UO_1170 (O_1170,N_19964,N_19875);
xor UO_1171 (O_1171,N_19916,N_19869);
or UO_1172 (O_1172,N_19802,N_19867);
xor UO_1173 (O_1173,N_19783,N_19976);
nor UO_1174 (O_1174,N_19900,N_19843);
nor UO_1175 (O_1175,N_19952,N_19880);
xor UO_1176 (O_1176,N_19978,N_19763);
nand UO_1177 (O_1177,N_19797,N_19777);
nand UO_1178 (O_1178,N_19794,N_19958);
and UO_1179 (O_1179,N_19935,N_19982);
nand UO_1180 (O_1180,N_19971,N_19815);
nor UO_1181 (O_1181,N_19951,N_19990);
or UO_1182 (O_1182,N_19920,N_19808);
xnor UO_1183 (O_1183,N_19887,N_19750);
nand UO_1184 (O_1184,N_19978,N_19886);
or UO_1185 (O_1185,N_19896,N_19944);
nand UO_1186 (O_1186,N_19804,N_19921);
or UO_1187 (O_1187,N_19956,N_19754);
nand UO_1188 (O_1188,N_19945,N_19750);
nor UO_1189 (O_1189,N_19992,N_19912);
xor UO_1190 (O_1190,N_19960,N_19926);
nand UO_1191 (O_1191,N_19841,N_19995);
xnor UO_1192 (O_1192,N_19843,N_19845);
nand UO_1193 (O_1193,N_19938,N_19822);
or UO_1194 (O_1194,N_19758,N_19886);
nand UO_1195 (O_1195,N_19927,N_19983);
nand UO_1196 (O_1196,N_19940,N_19890);
nand UO_1197 (O_1197,N_19755,N_19812);
xnor UO_1198 (O_1198,N_19781,N_19923);
nand UO_1199 (O_1199,N_19953,N_19909);
xnor UO_1200 (O_1200,N_19824,N_19814);
nand UO_1201 (O_1201,N_19872,N_19821);
and UO_1202 (O_1202,N_19814,N_19998);
nand UO_1203 (O_1203,N_19856,N_19788);
nor UO_1204 (O_1204,N_19861,N_19827);
xnor UO_1205 (O_1205,N_19752,N_19906);
xnor UO_1206 (O_1206,N_19846,N_19950);
and UO_1207 (O_1207,N_19980,N_19901);
xor UO_1208 (O_1208,N_19789,N_19913);
nor UO_1209 (O_1209,N_19751,N_19848);
xor UO_1210 (O_1210,N_19888,N_19832);
and UO_1211 (O_1211,N_19917,N_19862);
nand UO_1212 (O_1212,N_19874,N_19986);
nand UO_1213 (O_1213,N_19872,N_19773);
or UO_1214 (O_1214,N_19903,N_19791);
and UO_1215 (O_1215,N_19758,N_19785);
xor UO_1216 (O_1216,N_19885,N_19905);
xnor UO_1217 (O_1217,N_19976,N_19750);
and UO_1218 (O_1218,N_19918,N_19760);
xor UO_1219 (O_1219,N_19990,N_19890);
nand UO_1220 (O_1220,N_19895,N_19985);
and UO_1221 (O_1221,N_19783,N_19758);
and UO_1222 (O_1222,N_19908,N_19970);
nand UO_1223 (O_1223,N_19795,N_19878);
xnor UO_1224 (O_1224,N_19990,N_19997);
nand UO_1225 (O_1225,N_19861,N_19757);
nand UO_1226 (O_1226,N_19867,N_19932);
or UO_1227 (O_1227,N_19934,N_19929);
and UO_1228 (O_1228,N_19767,N_19999);
and UO_1229 (O_1229,N_19929,N_19990);
nand UO_1230 (O_1230,N_19791,N_19756);
and UO_1231 (O_1231,N_19918,N_19994);
and UO_1232 (O_1232,N_19907,N_19885);
nand UO_1233 (O_1233,N_19906,N_19792);
and UO_1234 (O_1234,N_19998,N_19970);
and UO_1235 (O_1235,N_19971,N_19779);
xnor UO_1236 (O_1236,N_19861,N_19780);
nor UO_1237 (O_1237,N_19948,N_19815);
nor UO_1238 (O_1238,N_19758,N_19980);
nor UO_1239 (O_1239,N_19758,N_19784);
nand UO_1240 (O_1240,N_19881,N_19842);
and UO_1241 (O_1241,N_19953,N_19948);
xor UO_1242 (O_1242,N_19835,N_19990);
xor UO_1243 (O_1243,N_19947,N_19849);
nor UO_1244 (O_1244,N_19836,N_19851);
nor UO_1245 (O_1245,N_19802,N_19877);
xnor UO_1246 (O_1246,N_19938,N_19994);
or UO_1247 (O_1247,N_19838,N_19940);
nand UO_1248 (O_1248,N_19980,N_19969);
or UO_1249 (O_1249,N_19998,N_19785);
xor UO_1250 (O_1250,N_19754,N_19823);
xor UO_1251 (O_1251,N_19962,N_19847);
xnor UO_1252 (O_1252,N_19944,N_19778);
nor UO_1253 (O_1253,N_19967,N_19779);
xor UO_1254 (O_1254,N_19808,N_19972);
or UO_1255 (O_1255,N_19895,N_19922);
nor UO_1256 (O_1256,N_19879,N_19770);
or UO_1257 (O_1257,N_19961,N_19792);
and UO_1258 (O_1258,N_19799,N_19894);
xnor UO_1259 (O_1259,N_19826,N_19829);
nand UO_1260 (O_1260,N_19775,N_19778);
nand UO_1261 (O_1261,N_19867,N_19975);
nor UO_1262 (O_1262,N_19996,N_19836);
or UO_1263 (O_1263,N_19970,N_19964);
nand UO_1264 (O_1264,N_19923,N_19838);
nand UO_1265 (O_1265,N_19988,N_19987);
or UO_1266 (O_1266,N_19897,N_19985);
and UO_1267 (O_1267,N_19955,N_19890);
nor UO_1268 (O_1268,N_19904,N_19974);
nand UO_1269 (O_1269,N_19829,N_19930);
nand UO_1270 (O_1270,N_19807,N_19998);
nand UO_1271 (O_1271,N_19771,N_19955);
xor UO_1272 (O_1272,N_19923,N_19955);
nor UO_1273 (O_1273,N_19987,N_19933);
nor UO_1274 (O_1274,N_19994,N_19758);
nand UO_1275 (O_1275,N_19962,N_19941);
or UO_1276 (O_1276,N_19956,N_19883);
xor UO_1277 (O_1277,N_19930,N_19836);
nor UO_1278 (O_1278,N_19859,N_19772);
or UO_1279 (O_1279,N_19876,N_19782);
or UO_1280 (O_1280,N_19950,N_19907);
nor UO_1281 (O_1281,N_19916,N_19796);
nor UO_1282 (O_1282,N_19968,N_19844);
nor UO_1283 (O_1283,N_19962,N_19981);
xor UO_1284 (O_1284,N_19850,N_19807);
and UO_1285 (O_1285,N_19958,N_19761);
nor UO_1286 (O_1286,N_19767,N_19840);
xor UO_1287 (O_1287,N_19794,N_19923);
nor UO_1288 (O_1288,N_19932,N_19968);
xor UO_1289 (O_1289,N_19870,N_19891);
xnor UO_1290 (O_1290,N_19864,N_19760);
xnor UO_1291 (O_1291,N_19757,N_19990);
or UO_1292 (O_1292,N_19979,N_19913);
xnor UO_1293 (O_1293,N_19956,N_19750);
and UO_1294 (O_1294,N_19968,N_19972);
and UO_1295 (O_1295,N_19846,N_19759);
and UO_1296 (O_1296,N_19933,N_19893);
and UO_1297 (O_1297,N_19805,N_19838);
xor UO_1298 (O_1298,N_19913,N_19820);
nor UO_1299 (O_1299,N_19758,N_19971);
and UO_1300 (O_1300,N_19801,N_19815);
nor UO_1301 (O_1301,N_19952,N_19853);
nand UO_1302 (O_1302,N_19948,N_19821);
xor UO_1303 (O_1303,N_19931,N_19894);
or UO_1304 (O_1304,N_19873,N_19802);
or UO_1305 (O_1305,N_19805,N_19797);
nor UO_1306 (O_1306,N_19915,N_19966);
and UO_1307 (O_1307,N_19753,N_19975);
nand UO_1308 (O_1308,N_19810,N_19961);
nor UO_1309 (O_1309,N_19795,N_19771);
nor UO_1310 (O_1310,N_19983,N_19973);
nor UO_1311 (O_1311,N_19822,N_19751);
xor UO_1312 (O_1312,N_19807,N_19814);
and UO_1313 (O_1313,N_19858,N_19791);
nand UO_1314 (O_1314,N_19824,N_19792);
and UO_1315 (O_1315,N_19883,N_19984);
and UO_1316 (O_1316,N_19858,N_19820);
and UO_1317 (O_1317,N_19905,N_19999);
and UO_1318 (O_1318,N_19769,N_19935);
nand UO_1319 (O_1319,N_19770,N_19875);
xor UO_1320 (O_1320,N_19871,N_19897);
nor UO_1321 (O_1321,N_19952,N_19860);
nand UO_1322 (O_1322,N_19909,N_19837);
and UO_1323 (O_1323,N_19768,N_19835);
or UO_1324 (O_1324,N_19883,N_19848);
and UO_1325 (O_1325,N_19875,N_19815);
or UO_1326 (O_1326,N_19956,N_19835);
nor UO_1327 (O_1327,N_19863,N_19955);
nor UO_1328 (O_1328,N_19973,N_19859);
xor UO_1329 (O_1329,N_19793,N_19972);
or UO_1330 (O_1330,N_19821,N_19957);
and UO_1331 (O_1331,N_19753,N_19879);
or UO_1332 (O_1332,N_19867,N_19917);
nand UO_1333 (O_1333,N_19980,N_19804);
or UO_1334 (O_1334,N_19858,N_19969);
and UO_1335 (O_1335,N_19994,N_19840);
xnor UO_1336 (O_1336,N_19879,N_19878);
and UO_1337 (O_1337,N_19826,N_19966);
nor UO_1338 (O_1338,N_19840,N_19939);
or UO_1339 (O_1339,N_19888,N_19930);
xor UO_1340 (O_1340,N_19811,N_19876);
and UO_1341 (O_1341,N_19825,N_19962);
or UO_1342 (O_1342,N_19954,N_19866);
or UO_1343 (O_1343,N_19829,N_19785);
or UO_1344 (O_1344,N_19929,N_19956);
nor UO_1345 (O_1345,N_19769,N_19795);
or UO_1346 (O_1346,N_19959,N_19956);
and UO_1347 (O_1347,N_19828,N_19767);
nand UO_1348 (O_1348,N_19860,N_19961);
nand UO_1349 (O_1349,N_19860,N_19819);
nor UO_1350 (O_1350,N_19784,N_19800);
xor UO_1351 (O_1351,N_19905,N_19923);
nand UO_1352 (O_1352,N_19772,N_19997);
and UO_1353 (O_1353,N_19803,N_19789);
nor UO_1354 (O_1354,N_19848,N_19776);
and UO_1355 (O_1355,N_19957,N_19965);
xnor UO_1356 (O_1356,N_19988,N_19941);
nand UO_1357 (O_1357,N_19829,N_19969);
and UO_1358 (O_1358,N_19799,N_19986);
nor UO_1359 (O_1359,N_19864,N_19765);
or UO_1360 (O_1360,N_19781,N_19949);
nand UO_1361 (O_1361,N_19932,N_19799);
and UO_1362 (O_1362,N_19795,N_19805);
nor UO_1363 (O_1363,N_19949,N_19800);
or UO_1364 (O_1364,N_19814,N_19779);
and UO_1365 (O_1365,N_19961,N_19937);
or UO_1366 (O_1366,N_19871,N_19971);
and UO_1367 (O_1367,N_19999,N_19895);
or UO_1368 (O_1368,N_19793,N_19999);
or UO_1369 (O_1369,N_19878,N_19778);
nor UO_1370 (O_1370,N_19822,N_19805);
nand UO_1371 (O_1371,N_19783,N_19936);
xor UO_1372 (O_1372,N_19750,N_19794);
nand UO_1373 (O_1373,N_19864,N_19893);
nand UO_1374 (O_1374,N_19915,N_19902);
nand UO_1375 (O_1375,N_19862,N_19923);
nand UO_1376 (O_1376,N_19936,N_19903);
xor UO_1377 (O_1377,N_19833,N_19787);
xnor UO_1378 (O_1378,N_19986,N_19845);
or UO_1379 (O_1379,N_19918,N_19896);
or UO_1380 (O_1380,N_19796,N_19910);
nor UO_1381 (O_1381,N_19758,N_19829);
nand UO_1382 (O_1382,N_19796,N_19951);
nand UO_1383 (O_1383,N_19996,N_19982);
xor UO_1384 (O_1384,N_19958,N_19915);
nor UO_1385 (O_1385,N_19954,N_19897);
xor UO_1386 (O_1386,N_19863,N_19990);
xor UO_1387 (O_1387,N_19924,N_19803);
xor UO_1388 (O_1388,N_19887,N_19948);
or UO_1389 (O_1389,N_19838,N_19751);
or UO_1390 (O_1390,N_19765,N_19798);
nand UO_1391 (O_1391,N_19802,N_19779);
nor UO_1392 (O_1392,N_19824,N_19955);
xor UO_1393 (O_1393,N_19897,N_19941);
xnor UO_1394 (O_1394,N_19815,N_19809);
or UO_1395 (O_1395,N_19962,N_19932);
xnor UO_1396 (O_1396,N_19828,N_19827);
xor UO_1397 (O_1397,N_19881,N_19852);
nand UO_1398 (O_1398,N_19913,N_19921);
or UO_1399 (O_1399,N_19784,N_19892);
nand UO_1400 (O_1400,N_19865,N_19990);
nand UO_1401 (O_1401,N_19811,N_19851);
and UO_1402 (O_1402,N_19935,N_19871);
xnor UO_1403 (O_1403,N_19839,N_19998);
nor UO_1404 (O_1404,N_19945,N_19845);
nand UO_1405 (O_1405,N_19983,N_19953);
xor UO_1406 (O_1406,N_19949,N_19771);
and UO_1407 (O_1407,N_19901,N_19954);
xnor UO_1408 (O_1408,N_19952,N_19879);
nor UO_1409 (O_1409,N_19821,N_19916);
and UO_1410 (O_1410,N_19960,N_19892);
nor UO_1411 (O_1411,N_19823,N_19979);
nand UO_1412 (O_1412,N_19903,N_19957);
xor UO_1413 (O_1413,N_19774,N_19858);
xnor UO_1414 (O_1414,N_19772,N_19779);
xor UO_1415 (O_1415,N_19907,N_19989);
nand UO_1416 (O_1416,N_19949,N_19851);
nand UO_1417 (O_1417,N_19969,N_19936);
or UO_1418 (O_1418,N_19988,N_19820);
and UO_1419 (O_1419,N_19813,N_19950);
or UO_1420 (O_1420,N_19976,N_19916);
nand UO_1421 (O_1421,N_19989,N_19983);
and UO_1422 (O_1422,N_19863,N_19907);
xor UO_1423 (O_1423,N_19867,N_19795);
and UO_1424 (O_1424,N_19808,N_19766);
nor UO_1425 (O_1425,N_19957,N_19986);
nand UO_1426 (O_1426,N_19780,N_19754);
nand UO_1427 (O_1427,N_19823,N_19857);
xnor UO_1428 (O_1428,N_19777,N_19788);
or UO_1429 (O_1429,N_19999,N_19989);
nand UO_1430 (O_1430,N_19880,N_19999);
or UO_1431 (O_1431,N_19760,N_19818);
or UO_1432 (O_1432,N_19887,N_19873);
xor UO_1433 (O_1433,N_19959,N_19936);
nor UO_1434 (O_1434,N_19956,N_19757);
xor UO_1435 (O_1435,N_19792,N_19974);
and UO_1436 (O_1436,N_19932,N_19928);
nand UO_1437 (O_1437,N_19989,N_19790);
xnor UO_1438 (O_1438,N_19763,N_19778);
xor UO_1439 (O_1439,N_19986,N_19816);
xnor UO_1440 (O_1440,N_19910,N_19761);
nor UO_1441 (O_1441,N_19918,N_19775);
and UO_1442 (O_1442,N_19885,N_19855);
xor UO_1443 (O_1443,N_19958,N_19891);
or UO_1444 (O_1444,N_19918,N_19899);
xnor UO_1445 (O_1445,N_19926,N_19775);
or UO_1446 (O_1446,N_19941,N_19826);
and UO_1447 (O_1447,N_19899,N_19903);
or UO_1448 (O_1448,N_19756,N_19906);
nand UO_1449 (O_1449,N_19958,N_19787);
xor UO_1450 (O_1450,N_19921,N_19851);
nand UO_1451 (O_1451,N_19835,N_19844);
xnor UO_1452 (O_1452,N_19968,N_19754);
or UO_1453 (O_1453,N_19763,N_19893);
and UO_1454 (O_1454,N_19878,N_19927);
or UO_1455 (O_1455,N_19952,N_19759);
xor UO_1456 (O_1456,N_19995,N_19965);
or UO_1457 (O_1457,N_19769,N_19946);
and UO_1458 (O_1458,N_19973,N_19919);
or UO_1459 (O_1459,N_19949,N_19760);
or UO_1460 (O_1460,N_19880,N_19812);
xnor UO_1461 (O_1461,N_19864,N_19855);
and UO_1462 (O_1462,N_19963,N_19916);
nor UO_1463 (O_1463,N_19864,N_19773);
nand UO_1464 (O_1464,N_19886,N_19884);
nor UO_1465 (O_1465,N_19758,N_19800);
and UO_1466 (O_1466,N_19903,N_19792);
nand UO_1467 (O_1467,N_19971,N_19992);
and UO_1468 (O_1468,N_19778,N_19987);
xnor UO_1469 (O_1469,N_19928,N_19943);
nand UO_1470 (O_1470,N_19834,N_19837);
xor UO_1471 (O_1471,N_19938,N_19800);
xor UO_1472 (O_1472,N_19934,N_19886);
or UO_1473 (O_1473,N_19850,N_19861);
xor UO_1474 (O_1474,N_19977,N_19916);
nand UO_1475 (O_1475,N_19969,N_19756);
nor UO_1476 (O_1476,N_19786,N_19833);
or UO_1477 (O_1477,N_19857,N_19787);
and UO_1478 (O_1478,N_19838,N_19770);
or UO_1479 (O_1479,N_19812,N_19984);
xnor UO_1480 (O_1480,N_19898,N_19984);
nand UO_1481 (O_1481,N_19960,N_19967);
xnor UO_1482 (O_1482,N_19985,N_19871);
or UO_1483 (O_1483,N_19810,N_19980);
nor UO_1484 (O_1484,N_19856,N_19975);
nand UO_1485 (O_1485,N_19799,N_19931);
xor UO_1486 (O_1486,N_19926,N_19846);
nor UO_1487 (O_1487,N_19956,N_19808);
or UO_1488 (O_1488,N_19883,N_19902);
or UO_1489 (O_1489,N_19963,N_19785);
nand UO_1490 (O_1490,N_19776,N_19820);
nand UO_1491 (O_1491,N_19976,N_19952);
or UO_1492 (O_1492,N_19855,N_19924);
and UO_1493 (O_1493,N_19819,N_19777);
nand UO_1494 (O_1494,N_19956,N_19807);
nand UO_1495 (O_1495,N_19870,N_19845);
nand UO_1496 (O_1496,N_19799,N_19876);
or UO_1497 (O_1497,N_19960,N_19828);
xor UO_1498 (O_1498,N_19863,N_19799);
xor UO_1499 (O_1499,N_19781,N_19858);
nand UO_1500 (O_1500,N_19838,N_19948);
nand UO_1501 (O_1501,N_19885,N_19865);
or UO_1502 (O_1502,N_19797,N_19846);
nand UO_1503 (O_1503,N_19813,N_19859);
nand UO_1504 (O_1504,N_19807,N_19805);
xor UO_1505 (O_1505,N_19775,N_19812);
and UO_1506 (O_1506,N_19920,N_19802);
or UO_1507 (O_1507,N_19783,N_19872);
and UO_1508 (O_1508,N_19798,N_19781);
xor UO_1509 (O_1509,N_19986,N_19901);
and UO_1510 (O_1510,N_19772,N_19803);
xnor UO_1511 (O_1511,N_19819,N_19853);
nor UO_1512 (O_1512,N_19909,N_19979);
nand UO_1513 (O_1513,N_19942,N_19881);
or UO_1514 (O_1514,N_19816,N_19851);
and UO_1515 (O_1515,N_19937,N_19845);
xor UO_1516 (O_1516,N_19898,N_19903);
nor UO_1517 (O_1517,N_19811,N_19934);
or UO_1518 (O_1518,N_19832,N_19849);
xor UO_1519 (O_1519,N_19960,N_19848);
nor UO_1520 (O_1520,N_19772,N_19780);
nor UO_1521 (O_1521,N_19954,N_19873);
and UO_1522 (O_1522,N_19854,N_19944);
xnor UO_1523 (O_1523,N_19946,N_19980);
nor UO_1524 (O_1524,N_19904,N_19876);
nor UO_1525 (O_1525,N_19825,N_19988);
and UO_1526 (O_1526,N_19936,N_19919);
or UO_1527 (O_1527,N_19898,N_19759);
and UO_1528 (O_1528,N_19827,N_19768);
or UO_1529 (O_1529,N_19798,N_19846);
nor UO_1530 (O_1530,N_19807,N_19769);
and UO_1531 (O_1531,N_19940,N_19886);
nor UO_1532 (O_1532,N_19864,N_19786);
nor UO_1533 (O_1533,N_19878,N_19769);
nor UO_1534 (O_1534,N_19823,N_19784);
xor UO_1535 (O_1535,N_19827,N_19964);
xnor UO_1536 (O_1536,N_19984,N_19930);
xor UO_1537 (O_1537,N_19834,N_19870);
and UO_1538 (O_1538,N_19944,N_19919);
nand UO_1539 (O_1539,N_19831,N_19923);
or UO_1540 (O_1540,N_19990,N_19794);
xnor UO_1541 (O_1541,N_19831,N_19770);
or UO_1542 (O_1542,N_19825,N_19991);
nand UO_1543 (O_1543,N_19974,N_19949);
xnor UO_1544 (O_1544,N_19936,N_19993);
and UO_1545 (O_1545,N_19890,N_19931);
or UO_1546 (O_1546,N_19894,N_19779);
or UO_1547 (O_1547,N_19975,N_19813);
nor UO_1548 (O_1548,N_19965,N_19837);
nor UO_1549 (O_1549,N_19900,N_19756);
and UO_1550 (O_1550,N_19989,N_19772);
or UO_1551 (O_1551,N_19790,N_19822);
and UO_1552 (O_1552,N_19765,N_19766);
xnor UO_1553 (O_1553,N_19969,N_19813);
nor UO_1554 (O_1554,N_19873,N_19849);
or UO_1555 (O_1555,N_19838,N_19928);
and UO_1556 (O_1556,N_19808,N_19838);
nor UO_1557 (O_1557,N_19952,N_19833);
nand UO_1558 (O_1558,N_19907,N_19890);
xor UO_1559 (O_1559,N_19951,N_19980);
xnor UO_1560 (O_1560,N_19756,N_19956);
xnor UO_1561 (O_1561,N_19888,N_19768);
or UO_1562 (O_1562,N_19972,N_19914);
nor UO_1563 (O_1563,N_19828,N_19805);
or UO_1564 (O_1564,N_19895,N_19897);
nand UO_1565 (O_1565,N_19902,N_19787);
or UO_1566 (O_1566,N_19957,N_19862);
or UO_1567 (O_1567,N_19804,N_19966);
or UO_1568 (O_1568,N_19781,N_19790);
nor UO_1569 (O_1569,N_19870,N_19960);
xnor UO_1570 (O_1570,N_19935,N_19946);
xnor UO_1571 (O_1571,N_19797,N_19849);
nand UO_1572 (O_1572,N_19813,N_19825);
or UO_1573 (O_1573,N_19832,N_19865);
or UO_1574 (O_1574,N_19954,N_19884);
xor UO_1575 (O_1575,N_19981,N_19928);
xnor UO_1576 (O_1576,N_19967,N_19795);
xor UO_1577 (O_1577,N_19921,N_19846);
nor UO_1578 (O_1578,N_19770,N_19942);
and UO_1579 (O_1579,N_19810,N_19778);
nand UO_1580 (O_1580,N_19766,N_19946);
nand UO_1581 (O_1581,N_19960,N_19865);
nor UO_1582 (O_1582,N_19904,N_19920);
and UO_1583 (O_1583,N_19872,N_19961);
and UO_1584 (O_1584,N_19801,N_19997);
or UO_1585 (O_1585,N_19954,N_19874);
xor UO_1586 (O_1586,N_19762,N_19780);
or UO_1587 (O_1587,N_19984,N_19858);
nor UO_1588 (O_1588,N_19758,N_19989);
nand UO_1589 (O_1589,N_19848,N_19783);
and UO_1590 (O_1590,N_19787,N_19926);
and UO_1591 (O_1591,N_19772,N_19907);
nand UO_1592 (O_1592,N_19975,N_19832);
xnor UO_1593 (O_1593,N_19828,N_19884);
nand UO_1594 (O_1594,N_19838,N_19971);
nand UO_1595 (O_1595,N_19992,N_19754);
xor UO_1596 (O_1596,N_19878,N_19761);
and UO_1597 (O_1597,N_19755,N_19827);
or UO_1598 (O_1598,N_19869,N_19781);
and UO_1599 (O_1599,N_19926,N_19920);
nand UO_1600 (O_1600,N_19764,N_19882);
nor UO_1601 (O_1601,N_19872,N_19935);
and UO_1602 (O_1602,N_19853,N_19868);
nand UO_1603 (O_1603,N_19931,N_19804);
nand UO_1604 (O_1604,N_19967,N_19949);
xnor UO_1605 (O_1605,N_19885,N_19903);
and UO_1606 (O_1606,N_19769,N_19870);
nor UO_1607 (O_1607,N_19948,N_19844);
xor UO_1608 (O_1608,N_19932,N_19787);
xnor UO_1609 (O_1609,N_19774,N_19775);
nor UO_1610 (O_1610,N_19986,N_19975);
nor UO_1611 (O_1611,N_19822,N_19964);
xnor UO_1612 (O_1612,N_19954,N_19859);
or UO_1613 (O_1613,N_19991,N_19863);
xor UO_1614 (O_1614,N_19801,N_19911);
xnor UO_1615 (O_1615,N_19766,N_19995);
xnor UO_1616 (O_1616,N_19757,N_19865);
or UO_1617 (O_1617,N_19799,N_19813);
and UO_1618 (O_1618,N_19945,N_19853);
xnor UO_1619 (O_1619,N_19928,N_19851);
or UO_1620 (O_1620,N_19806,N_19781);
nand UO_1621 (O_1621,N_19826,N_19827);
xnor UO_1622 (O_1622,N_19845,N_19801);
nor UO_1623 (O_1623,N_19806,N_19778);
or UO_1624 (O_1624,N_19836,N_19911);
or UO_1625 (O_1625,N_19885,N_19860);
nand UO_1626 (O_1626,N_19939,N_19814);
xor UO_1627 (O_1627,N_19897,N_19918);
nand UO_1628 (O_1628,N_19877,N_19850);
nor UO_1629 (O_1629,N_19957,N_19919);
xor UO_1630 (O_1630,N_19767,N_19859);
nand UO_1631 (O_1631,N_19752,N_19794);
and UO_1632 (O_1632,N_19840,N_19965);
and UO_1633 (O_1633,N_19970,N_19814);
xnor UO_1634 (O_1634,N_19983,N_19866);
and UO_1635 (O_1635,N_19933,N_19926);
nor UO_1636 (O_1636,N_19754,N_19758);
nor UO_1637 (O_1637,N_19784,N_19967);
nor UO_1638 (O_1638,N_19834,N_19847);
nor UO_1639 (O_1639,N_19940,N_19947);
or UO_1640 (O_1640,N_19820,N_19936);
nand UO_1641 (O_1641,N_19783,N_19975);
nand UO_1642 (O_1642,N_19983,N_19919);
nand UO_1643 (O_1643,N_19774,N_19952);
or UO_1644 (O_1644,N_19940,N_19937);
and UO_1645 (O_1645,N_19805,N_19921);
nor UO_1646 (O_1646,N_19987,N_19890);
nand UO_1647 (O_1647,N_19787,N_19750);
and UO_1648 (O_1648,N_19929,N_19962);
nand UO_1649 (O_1649,N_19965,N_19811);
or UO_1650 (O_1650,N_19921,N_19772);
or UO_1651 (O_1651,N_19913,N_19853);
nand UO_1652 (O_1652,N_19771,N_19883);
nand UO_1653 (O_1653,N_19941,N_19983);
xor UO_1654 (O_1654,N_19878,N_19888);
xor UO_1655 (O_1655,N_19996,N_19930);
and UO_1656 (O_1656,N_19854,N_19906);
xor UO_1657 (O_1657,N_19780,N_19806);
and UO_1658 (O_1658,N_19789,N_19931);
xor UO_1659 (O_1659,N_19938,N_19979);
and UO_1660 (O_1660,N_19962,N_19837);
nor UO_1661 (O_1661,N_19837,N_19826);
or UO_1662 (O_1662,N_19757,N_19829);
nand UO_1663 (O_1663,N_19974,N_19751);
or UO_1664 (O_1664,N_19898,N_19899);
nor UO_1665 (O_1665,N_19767,N_19962);
xor UO_1666 (O_1666,N_19916,N_19907);
or UO_1667 (O_1667,N_19978,N_19822);
nor UO_1668 (O_1668,N_19986,N_19815);
and UO_1669 (O_1669,N_19861,N_19928);
and UO_1670 (O_1670,N_19810,N_19776);
nand UO_1671 (O_1671,N_19914,N_19755);
and UO_1672 (O_1672,N_19858,N_19877);
and UO_1673 (O_1673,N_19947,N_19932);
nor UO_1674 (O_1674,N_19824,N_19906);
and UO_1675 (O_1675,N_19954,N_19806);
or UO_1676 (O_1676,N_19963,N_19880);
nand UO_1677 (O_1677,N_19750,N_19989);
or UO_1678 (O_1678,N_19750,N_19910);
nand UO_1679 (O_1679,N_19830,N_19800);
and UO_1680 (O_1680,N_19782,N_19802);
xnor UO_1681 (O_1681,N_19822,N_19759);
xor UO_1682 (O_1682,N_19835,N_19816);
nand UO_1683 (O_1683,N_19971,N_19872);
or UO_1684 (O_1684,N_19919,N_19901);
or UO_1685 (O_1685,N_19886,N_19800);
nor UO_1686 (O_1686,N_19845,N_19832);
or UO_1687 (O_1687,N_19894,N_19900);
xor UO_1688 (O_1688,N_19831,N_19916);
xor UO_1689 (O_1689,N_19940,N_19843);
or UO_1690 (O_1690,N_19822,N_19858);
and UO_1691 (O_1691,N_19796,N_19983);
and UO_1692 (O_1692,N_19835,N_19760);
nor UO_1693 (O_1693,N_19760,N_19843);
nor UO_1694 (O_1694,N_19846,N_19779);
xor UO_1695 (O_1695,N_19903,N_19895);
xor UO_1696 (O_1696,N_19939,N_19991);
or UO_1697 (O_1697,N_19985,N_19890);
or UO_1698 (O_1698,N_19873,N_19935);
or UO_1699 (O_1699,N_19865,N_19969);
or UO_1700 (O_1700,N_19886,N_19883);
nand UO_1701 (O_1701,N_19810,N_19936);
and UO_1702 (O_1702,N_19880,N_19882);
or UO_1703 (O_1703,N_19998,N_19918);
xor UO_1704 (O_1704,N_19932,N_19785);
xor UO_1705 (O_1705,N_19965,N_19985);
and UO_1706 (O_1706,N_19988,N_19943);
nand UO_1707 (O_1707,N_19963,N_19769);
or UO_1708 (O_1708,N_19958,N_19938);
or UO_1709 (O_1709,N_19765,N_19884);
or UO_1710 (O_1710,N_19898,N_19782);
and UO_1711 (O_1711,N_19890,N_19904);
nor UO_1712 (O_1712,N_19975,N_19773);
and UO_1713 (O_1713,N_19993,N_19918);
nand UO_1714 (O_1714,N_19947,N_19790);
nand UO_1715 (O_1715,N_19995,N_19904);
or UO_1716 (O_1716,N_19984,N_19828);
or UO_1717 (O_1717,N_19867,N_19981);
xnor UO_1718 (O_1718,N_19786,N_19981);
nand UO_1719 (O_1719,N_19946,N_19822);
and UO_1720 (O_1720,N_19870,N_19910);
or UO_1721 (O_1721,N_19853,N_19869);
nor UO_1722 (O_1722,N_19750,N_19876);
nand UO_1723 (O_1723,N_19805,N_19775);
nor UO_1724 (O_1724,N_19828,N_19895);
nor UO_1725 (O_1725,N_19946,N_19821);
nand UO_1726 (O_1726,N_19795,N_19946);
or UO_1727 (O_1727,N_19904,N_19853);
or UO_1728 (O_1728,N_19891,N_19757);
or UO_1729 (O_1729,N_19828,N_19965);
nor UO_1730 (O_1730,N_19903,N_19934);
xnor UO_1731 (O_1731,N_19924,N_19830);
nor UO_1732 (O_1732,N_19976,N_19837);
and UO_1733 (O_1733,N_19939,N_19885);
xnor UO_1734 (O_1734,N_19752,N_19841);
and UO_1735 (O_1735,N_19772,N_19784);
and UO_1736 (O_1736,N_19822,N_19931);
nand UO_1737 (O_1737,N_19788,N_19888);
and UO_1738 (O_1738,N_19977,N_19959);
xor UO_1739 (O_1739,N_19823,N_19852);
xor UO_1740 (O_1740,N_19999,N_19777);
nand UO_1741 (O_1741,N_19972,N_19908);
and UO_1742 (O_1742,N_19806,N_19876);
nor UO_1743 (O_1743,N_19853,N_19801);
nand UO_1744 (O_1744,N_19927,N_19897);
nand UO_1745 (O_1745,N_19853,N_19979);
or UO_1746 (O_1746,N_19817,N_19934);
or UO_1747 (O_1747,N_19815,N_19997);
nand UO_1748 (O_1748,N_19902,N_19908);
or UO_1749 (O_1749,N_19970,N_19892);
and UO_1750 (O_1750,N_19859,N_19842);
nor UO_1751 (O_1751,N_19951,N_19789);
xor UO_1752 (O_1752,N_19795,N_19834);
nor UO_1753 (O_1753,N_19911,N_19971);
xor UO_1754 (O_1754,N_19963,N_19930);
nand UO_1755 (O_1755,N_19759,N_19987);
nand UO_1756 (O_1756,N_19770,N_19809);
or UO_1757 (O_1757,N_19820,N_19875);
and UO_1758 (O_1758,N_19804,N_19791);
and UO_1759 (O_1759,N_19936,N_19768);
or UO_1760 (O_1760,N_19787,N_19860);
or UO_1761 (O_1761,N_19993,N_19902);
or UO_1762 (O_1762,N_19950,N_19927);
and UO_1763 (O_1763,N_19768,N_19937);
xnor UO_1764 (O_1764,N_19826,N_19769);
xnor UO_1765 (O_1765,N_19821,N_19801);
nor UO_1766 (O_1766,N_19808,N_19951);
and UO_1767 (O_1767,N_19890,N_19811);
nor UO_1768 (O_1768,N_19956,N_19953);
xor UO_1769 (O_1769,N_19939,N_19861);
nor UO_1770 (O_1770,N_19806,N_19896);
and UO_1771 (O_1771,N_19954,N_19925);
or UO_1772 (O_1772,N_19855,N_19883);
and UO_1773 (O_1773,N_19868,N_19973);
and UO_1774 (O_1774,N_19843,N_19889);
xor UO_1775 (O_1775,N_19773,N_19958);
nand UO_1776 (O_1776,N_19846,N_19811);
and UO_1777 (O_1777,N_19836,N_19751);
or UO_1778 (O_1778,N_19874,N_19997);
nor UO_1779 (O_1779,N_19989,N_19881);
or UO_1780 (O_1780,N_19794,N_19880);
and UO_1781 (O_1781,N_19757,N_19853);
nand UO_1782 (O_1782,N_19841,N_19904);
and UO_1783 (O_1783,N_19935,N_19859);
or UO_1784 (O_1784,N_19840,N_19958);
and UO_1785 (O_1785,N_19940,N_19898);
nor UO_1786 (O_1786,N_19857,N_19949);
or UO_1787 (O_1787,N_19930,N_19816);
nor UO_1788 (O_1788,N_19895,N_19944);
nor UO_1789 (O_1789,N_19955,N_19835);
xor UO_1790 (O_1790,N_19855,N_19862);
or UO_1791 (O_1791,N_19876,N_19994);
nor UO_1792 (O_1792,N_19925,N_19772);
nor UO_1793 (O_1793,N_19996,N_19786);
xnor UO_1794 (O_1794,N_19911,N_19822);
nor UO_1795 (O_1795,N_19947,N_19856);
xnor UO_1796 (O_1796,N_19975,N_19842);
xor UO_1797 (O_1797,N_19908,N_19782);
and UO_1798 (O_1798,N_19761,N_19780);
or UO_1799 (O_1799,N_19973,N_19960);
or UO_1800 (O_1800,N_19943,N_19815);
and UO_1801 (O_1801,N_19885,N_19886);
nor UO_1802 (O_1802,N_19766,N_19830);
or UO_1803 (O_1803,N_19806,N_19839);
nand UO_1804 (O_1804,N_19848,N_19986);
and UO_1805 (O_1805,N_19965,N_19841);
xnor UO_1806 (O_1806,N_19882,N_19959);
xnor UO_1807 (O_1807,N_19752,N_19795);
xor UO_1808 (O_1808,N_19794,N_19870);
xnor UO_1809 (O_1809,N_19767,N_19911);
and UO_1810 (O_1810,N_19859,N_19850);
xnor UO_1811 (O_1811,N_19952,N_19922);
and UO_1812 (O_1812,N_19796,N_19752);
and UO_1813 (O_1813,N_19795,N_19870);
and UO_1814 (O_1814,N_19868,N_19807);
nor UO_1815 (O_1815,N_19887,N_19805);
nor UO_1816 (O_1816,N_19762,N_19777);
xnor UO_1817 (O_1817,N_19919,N_19943);
nor UO_1818 (O_1818,N_19866,N_19817);
nand UO_1819 (O_1819,N_19760,N_19960);
or UO_1820 (O_1820,N_19955,N_19978);
nor UO_1821 (O_1821,N_19755,N_19772);
and UO_1822 (O_1822,N_19845,N_19977);
xnor UO_1823 (O_1823,N_19764,N_19802);
nand UO_1824 (O_1824,N_19876,N_19895);
nor UO_1825 (O_1825,N_19978,N_19924);
and UO_1826 (O_1826,N_19820,N_19964);
nand UO_1827 (O_1827,N_19819,N_19752);
nand UO_1828 (O_1828,N_19765,N_19846);
or UO_1829 (O_1829,N_19923,N_19933);
and UO_1830 (O_1830,N_19785,N_19946);
nand UO_1831 (O_1831,N_19878,N_19828);
xor UO_1832 (O_1832,N_19835,N_19937);
xnor UO_1833 (O_1833,N_19941,N_19812);
nand UO_1834 (O_1834,N_19989,N_19993);
or UO_1835 (O_1835,N_19899,N_19948);
or UO_1836 (O_1836,N_19803,N_19773);
nand UO_1837 (O_1837,N_19786,N_19804);
or UO_1838 (O_1838,N_19885,N_19880);
nor UO_1839 (O_1839,N_19811,N_19921);
nor UO_1840 (O_1840,N_19773,N_19976);
nand UO_1841 (O_1841,N_19799,N_19809);
and UO_1842 (O_1842,N_19751,N_19936);
or UO_1843 (O_1843,N_19810,N_19779);
or UO_1844 (O_1844,N_19796,N_19925);
and UO_1845 (O_1845,N_19938,N_19925);
nor UO_1846 (O_1846,N_19770,N_19980);
or UO_1847 (O_1847,N_19756,N_19836);
and UO_1848 (O_1848,N_19906,N_19766);
nor UO_1849 (O_1849,N_19994,N_19906);
and UO_1850 (O_1850,N_19938,N_19876);
nor UO_1851 (O_1851,N_19891,N_19898);
nor UO_1852 (O_1852,N_19979,N_19829);
and UO_1853 (O_1853,N_19988,N_19921);
and UO_1854 (O_1854,N_19963,N_19771);
nor UO_1855 (O_1855,N_19999,N_19902);
nand UO_1856 (O_1856,N_19897,N_19862);
xnor UO_1857 (O_1857,N_19879,N_19832);
nand UO_1858 (O_1858,N_19940,N_19798);
nand UO_1859 (O_1859,N_19985,N_19819);
xor UO_1860 (O_1860,N_19779,N_19847);
xnor UO_1861 (O_1861,N_19937,N_19928);
xor UO_1862 (O_1862,N_19877,N_19784);
nor UO_1863 (O_1863,N_19940,N_19835);
xnor UO_1864 (O_1864,N_19787,N_19858);
xnor UO_1865 (O_1865,N_19913,N_19973);
nor UO_1866 (O_1866,N_19832,N_19919);
nand UO_1867 (O_1867,N_19773,N_19847);
or UO_1868 (O_1868,N_19873,N_19922);
or UO_1869 (O_1869,N_19959,N_19858);
and UO_1870 (O_1870,N_19881,N_19897);
nand UO_1871 (O_1871,N_19981,N_19820);
or UO_1872 (O_1872,N_19967,N_19911);
xor UO_1873 (O_1873,N_19773,N_19821);
nand UO_1874 (O_1874,N_19890,N_19775);
xnor UO_1875 (O_1875,N_19823,N_19971);
nand UO_1876 (O_1876,N_19913,N_19788);
nand UO_1877 (O_1877,N_19841,N_19953);
xor UO_1878 (O_1878,N_19827,N_19878);
or UO_1879 (O_1879,N_19867,N_19990);
or UO_1880 (O_1880,N_19878,N_19810);
or UO_1881 (O_1881,N_19902,N_19820);
or UO_1882 (O_1882,N_19994,N_19855);
nor UO_1883 (O_1883,N_19862,N_19781);
nor UO_1884 (O_1884,N_19837,N_19756);
nand UO_1885 (O_1885,N_19892,N_19934);
nor UO_1886 (O_1886,N_19897,N_19873);
xnor UO_1887 (O_1887,N_19992,N_19906);
or UO_1888 (O_1888,N_19761,N_19853);
and UO_1889 (O_1889,N_19904,N_19824);
nor UO_1890 (O_1890,N_19902,N_19945);
nand UO_1891 (O_1891,N_19936,N_19890);
nand UO_1892 (O_1892,N_19817,N_19842);
xor UO_1893 (O_1893,N_19900,N_19953);
nand UO_1894 (O_1894,N_19821,N_19911);
nand UO_1895 (O_1895,N_19770,N_19912);
xor UO_1896 (O_1896,N_19845,N_19803);
nor UO_1897 (O_1897,N_19858,N_19962);
nand UO_1898 (O_1898,N_19948,N_19891);
nand UO_1899 (O_1899,N_19817,N_19972);
or UO_1900 (O_1900,N_19995,N_19849);
or UO_1901 (O_1901,N_19779,N_19941);
or UO_1902 (O_1902,N_19875,N_19777);
and UO_1903 (O_1903,N_19898,N_19954);
xor UO_1904 (O_1904,N_19959,N_19892);
nor UO_1905 (O_1905,N_19825,N_19963);
xor UO_1906 (O_1906,N_19841,N_19774);
and UO_1907 (O_1907,N_19832,N_19822);
or UO_1908 (O_1908,N_19905,N_19922);
nand UO_1909 (O_1909,N_19880,N_19854);
or UO_1910 (O_1910,N_19906,N_19770);
or UO_1911 (O_1911,N_19999,N_19852);
nand UO_1912 (O_1912,N_19801,N_19810);
or UO_1913 (O_1913,N_19755,N_19915);
xnor UO_1914 (O_1914,N_19902,N_19911);
nor UO_1915 (O_1915,N_19753,N_19965);
xor UO_1916 (O_1916,N_19765,N_19887);
nor UO_1917 (O_1917,N_19893,N_19814);
or UO_1918 (O_1918,N_19936,N_19977);
or UO_1919 (O_1919,N_19886,N_19813);
or UO_1920 (O_1920,N_19933,N_19797);
xor UO_1921 (O_1921,N_19867,N_19773);
nor UO_1922 (O_1922,N_19785,N_19885);
xnor UO_1923 (O_1923,N_19807,N_19750);
and UO_1924 (O_1924,N_19761,N_19795);
nor UO_1925 (O_1925,N_19994,N_19773);
and UO_1926 (O_1926,N_19822,N_19752);
nand UO_1927 (O_1927,N_19818,N_19766);
and UO_1928 (O_1928,N_19902,N_19896);
xnor UO_1929 (O_1929,N_19824,N_19825);
and UO_1930 (O_1930,N_19821,N_19750);
nor UO_1931 (O_1931,N_19999,N_19834);
nor UO_1932 (O_1932,N_19888,N_19948);
or UO_1933 (O_1933,N_19757,N_19760);
and UO_1934 (O_1934,N_19951,N_19953);
nor UO_1935 (O_1935,N_19753,N_19917);
nand UO_1936 (O_1936,N_19931,N_19937);
and UO_1937 (O_1937,N_19914,N_19797);
nor UO_1938 (O_1938,N_19809,N_19937);
and UO_1939 (O_1939,N_19974,N_19947);
xnor UO_1940 (O_1940,N_19854,N_19868);
nand UO_1941 (O_1941,N_19805,N_19791);
or UO_1942 (O_1942,N_19772,N_19922);
nor UO_1943 (O_1943,N_19894,N_19764);
xor UO_1944 (O_1944,N_19976,N_19899);
or UO_1945 (O_1945,N_19918,N_19807);
nor UO_1946 (O_1946,N_19935,N_19937);
xor UO_1947 (O_1947,N_19936,N_19757);
and UO_1948 (O_1948,N_19969,N_19943);
and UO_1949 (O_1949,N_19955,N_19831);
xnor UO_1950 (O_1950,N_19792,N_19837);
xor UO_1951 (O_1951,N_19762,N_19957);
nor UO_1952 (O_1952,N_19946,N_19845);
xnor UO_1953 (O_1953,N_19869,N_19791);
or UO_1954 (O_1954,N_19937,N_19920);
nand UO_1955 (O_1955,N_19997,N_19957);
xnor UO_1956 (O_1956,N_19959,N_19962);
or UO_1957 (O_1957,N_19947,N_19890);
or UO_1958 (O_1958,N_19951,N_19988);
xnor UO_1959 (O_1959,N_19750,N_19838);
xnor UO_1960 (O_1960,N_19880,N_19797);
or UO_1961 (O_1961,N_19926,N_19822);
nor UO_1962 (O_1962,N_19754,N_19868);
and UO_1963 (O_1963,N_19784,N_19901);
and UO_1964 (O_1964,N_19949,N_19898);
and UO_1965 (O_1965,N_19830,N_19895);
and UO_1966 (O_1966,N_19866,N_19950);
nor UO_1967 (O_1967,N_19914,N_19881);
and UO_1968 (O_1968,N_19874,N_19791);
xnor UO_1969 (O_1969,N_19820,N_19852);
or UO_1970 (O_1970,N_19884,N_19858);
or UO_1971 (O_1971,N_19942,N_19837);
xor UO_1972 (O_1972,N_19858,N_19936);
xor UO_1973 (O_1973,N_19765,N_19862);
nand UO_1974 (O_1974,N_19973,N_19753);
nor UO_1975 (O_1975,N_19752,N_19854);
nor UO_1976 (O_1976,N_19844,N_19818);
xnor UO_1977 (O_1977,N_19878,N_19752);
or UO_1978 (O_1978,N_19940,N_19873);
xnor UO_1979 (O_1979,N_19977,N_19938);
nor UO_1980 (O_1980,N_19994,N_19953);
xor UO_1981 (O_1981,N_19956,N_19878);
xor UO_1982 (O_1982,N_19771,N_19930);
nor UO_1983 (O_1983,N_19762,N_19867);
and UO_1984 (O_1984,N_19930,N_19794);
nor UO_1985 (O_1985,N_19920,N_19756);
nand UO_1986 (O_1986,N_19780,N_19997);
nand UO_1987 (O_1987,N_19913,N_19919);
nand UO_1988 (O_1988,N_19994,N_19904);
or UO_1989 (O_1989,N_19885,N_19931);
xnor UO_1990 (O_1990,N_19848,N_19831);
nand UO_1991 (O_1991,N_19838,N_19856);
xor UO_1992 (O_1992,N_19975,N_19875);
or UO_1993 (O_1993,N_19941,N_19891);
or UO_1994 (O_1994,N_19833,N_19925);
nand UO_1995 (O_1995,N_19910,N_19901);
or UO_1996 (O_1996,N_19956,N_19919);
nand UO_1997 (O_1997,N_19997,N_19753);
and UO_1998 (O_1998,N_19906,N_19844);
or UO_1999 (O_1999,N_19805,N_19938);
and UO_2000 (O_2000,N_19785,N_19819);
nor UO_2001 (O_2001,N_19806,N_19787);
nor UO_2002 (O_2002,N_19915,N_19853);
xnor UO_2003 (O_2003,N_19988,N_19847);
xor UO_2004 (O_2004,N_19770,N_19966);
nand UO_2005 (O_2005,N_19824,N_19800);
nand UO_2006 (O_2006,N_19816,N_19961);
nor UO_2007 (O_2007,N_19762,N_19783);
nand UO_2008 (O_2008,N_19956,N_19938);
and UO_2009 (O_2009,N_19984,N_19848);
and UO_2010 (O_2010,N_19955,N_19794);
or UO_2011 (O_2011,N_19983,N_19991);
and UO_2012 (O_2012,N_19941,N_19771);
nand UO_2013 (O_2013,N_19853,N_19958);
and UO_2014 (O_2014,N_19896,N_19912);
and UO_2015 (O_2015,N_19775,N_19989);
and UO_2016 (O_2016,N_19812,N_19989);
nor UO_2017 (O_2017,N_19971,N_19856);
and UO_2018 (O_2018,N_19914,N_19750);
nand UO_2019 (O_2019,N_19989,N_19849);
nor UO_2020 (O_2020,N_19868,N_19878);
or UO_2021 (O_2021,N_19980,N_19889);
nor UO_2022 (O_2022,N_19969,N_19929);
nand UO_2023 (O_2023,N_19898,N_19767);
nor UO_2024 (O_2024,N_19913,N_19833);
xnor UO_2025 (O_2025,N_19864,N_19829);
and UO_2026 (O_2026,N_19815,N_19810);
xnor UO_2027 (O_2027,N_19931,N_19922);
xnor UO_2028 (O_2028,N_19993,N_19938);
and UO_2029 (O_2029,N_19778,N_19764);
nor UO_2030 (O_2030,N_19881,N_19827);
nand UO_2031 (O_2031,N_19768,N_19767);
nor UO_2032 (O_2032,N_19880,N_19886);
nand UO_2033 (O_2033,N_19849,N_19853);
xor UO_2034 (O_2034,N_19765,N_19983);
nor UO_2035 (O_2035,N_19930,N_19864);
xor UO_2036 (O_2036,N_19978,N_19793);
nand UO_2037 (O_2037,N_19854,N_19783);
and UO_2038 (O_2038,N_19828,N_19930);
nand UO_2039 (O_2039,N_19991,N_19859);
nand UO_2040 (O_2040,N_19774,N_19880);
and UO_2041 (O_2041,N_19884,N_19896);
xor UO_2042 (O_2042,N_19876,N_19909);
nand UO_2043 (O_2043,N_19876,N_19789);
or UO_2044 (O_2044,N_19777,N_19892);
or UO_2045 (O_2045,N_19841,N_19808);
nor UO_2046 (O_2046,N_19906,N_19934);
or UO_2047 (O_2047,N_19780,N_19826);
or UO_2048 (O_2048,N_19902,N_19970);
or UO_2049 (O_2049,N_19957,N_19777);
nand UO_2050 (O_2050,N_19963,N_19887);
xnor UO_2051 (O_2051,N_19779,N_19755);
nor UO_2052 (O_2052,N_19874,N_19962);
xnor UO_2053 (O_2053,N_19972,N_19915);
nand UO_2054 (O_2054,N_19933,N_19974);
xnor UO_2055 (O_2055,N_19793,N_19863);
or UO_2056 (O_2056,N_19923,N_19910);
nor UO_2057 (O_2057,N_19904,N_19766);
and UO_2058 (O_2058,N_19964,N_19957);
xor UO_2059 (O_2059,N_19927,N_19917);
nand UO_2060 (O_2060,N_19926,N_19810);
or UO_2061 (O_2061,N_19880,N_19916);
and UO_2062 (O_2062,N_19791,N_19940);
xor UO_2063 (O_2063,N_19912,N_19962);
nor UO_2064 (O_2064,N_19766,N_19785);
nand UO_2065 (O_2065,N_19943,N_19771);
xor UO_2066 (O_2066,N_19860,N_19899);
xor UO_2067 (O_2067,N_19888,N_19903);
nor UO_2068 (O_2068,N_19800,N_19850);
nor UO_2069 (O_2069,N_19919,N_19937);
or UO_2070 (O_2070,N_19831,N_19820);
or UO_2071 (O_2071,N_19779,N_19899);
xor UO_2072 (O_2072,N_19832,N_19923);
or UO_2073 (O_2073,N_19920,N_19868);
and UO_2074 (O_2074,N_19795,N_19886);
nor UO_2075 (O_2075,N_19851,N_19902);
nand UO_2076 (O_2076,N_19804,N_19812);
or UO_2077 (O_2077,N_19934,N_19802);
nand UO_2078 (O_2078,N_19943,N_19760);
nor UO_2079 (O_2079,N_19885,N_19775);
or UO_2080 (O_2080,N_19974,N_19989);
or UO_2081 (O_2081,N_19884,N_19778);
or UO_2082 (O_2082,N_19901,N_19966);
xor UO_2083 (O_2083,N_19814,N_19804);
or UO_2084 (O_2084,N_19989,N_19879);
nand UO_2085 (O_2085,N_19750,N_19826);
xnor UO_2086 (O_2086,N_19877,N_19797);
nand UO_2087 (O_2087,N_19817,N_19828);
or UO_2088 (O_2088,N_19772,N_19874);
and UO_2089 (O_2089,N_19901,N_19960);
or UO_2090 (O_2090,N_19931,N_19915);
and UO_2091 (O_2091,N_19754,N_19973);
and UO_2092 (O_2092,N_19792,N_19752);
nor UO_2093 (O_2093,N_19867,N_19841);
and UO_2094 (O_2094,N_19823,N_19883);
xnor UO_2095 (O_2095,N_19982,N_19881);
or UO_2096 (O_2096,N_19843,N_19937);
or UO_2097 (O_2097,N_19912,N_19786);
and UO_2098 (O_2098,N_19922,N_19918);
nor UO_2099 (O_2099,N_19815,N_19793);
or UO_2100 (O_2100,N_19996,N_19873);
or UO_2101 (O_2101,N_19776,N_19767);
nand UO_2102 (O_2102,N_19830,N_19979);
nor UO_2103 (O_2103,N_19940,N_19792);
nand UO_2104 (O_2104,N_19874,N_19856);
xnor UO_2105 (O_2105,N_19761,N_19972);
and UO_2106 (O_2106,N_19805,N_19804);
nand UO_2107 (O_2107,N_19837,N_19920);
nor UO_2108 (O_2108,N_19812,N_19787);
and UO_2109 (O_2109,N_19765,N_19858);
nor UO_2110 (O_2110,N_19816,N_19935);
or UO_2111 (O_2111,N_19858,N_19921);
nand UO_2112 (O_2112,N_19893,N_19757);
or UO_2113 (O_2113,N_19941,N_19787);
or UO_2114 (O_2114,N_19781,N_19979);
or UO_2115 (O_2115,N_19809,N_19958);
nor UO_2116 (O_2116,N_19827,N_19994);
xnor UO_2117 (O_2117,N_19976,N_19780);
or UO_2118 (O_2118,N_19933,N_19998);
xnor UO_2119 (O_2119,N_19999,N_19868);
xnor UO_2120 (O_2120,N_19960,N_19801);
nor UO_2121 (O_2121,N_19785,N_19956);
and UO_2122 (O_2122,N_19849,N_19977);
or UO_2123 (O_2123,N_19813,N_19939);
and UO_2124 (O_2124,N_19804,N_19940);
nand UO_2125 (O_2125,N_19965,N_19953);
xor UO_2126 (O_2126,N_19969,N_19857);
and UO_2127 (O_2127,N_19821,N_19847);
xnor UO_2128 (O_2128,N_19913,N_19998);
nand UO_2129 (O_2129,N_19825,N_19865);
nor UO_2130 (O_2130,N_19952,N_19932);
xnor UO_2131 (O_2131,N_19956,N_19966);
and UO_2132 (O_2132,N_19882,N_19867);
nand UO_2133 (O_2133,N_19882,N_19841);
xor UO_2134 (O_2134,N_19766,N_19990);
xnor UO_2135 (O_2135,N_19859,N_19886);
or UO_2136 (O_2136,N_19832,N_19803);
or UO_2137 (O_2137,N_19803,N_19822);
nand UO_2138 (O_2138,N_19752,N_19899);
or UO_2139 (O_2139,N_19952,N_19907);
nor UO_2140 (O_2140,N_19828,N_19892);
or UO_2141 (O_2141,N_19826,N_19787);
xor UO_2142 (O_2142,N_19901,N_19777);
or UO_2143 (O_2143,N_19927,N_19881);
or UO_2144 (O_2144,N_19852,N_19978);
or UO_2145 (O_2145,N_19824,N_19833);
nor UO_2146 (O_2146,N_19777,N_19844);
and UO_2147 (O_2147,N_19892,N_19771);
nor UO_2148 (O_2148,N_19951,N_19934);
or UO_2149 (O_2149,N_19795,N_19823);
and UO_2150 (O_2150,N_19860,N_19816);
nand UO_2151 (O_2151,N_19871,N_19760);
nor UO_2152 (O_2152,N_19925,N_19752);
and UO_2153 (O_2153,N_19965,N_19771);
and UO_2154 (O_2154,N_19986,N_19987);
and UO_2155 (O_2155,N_19971,N_19757);
nor UO_2156 (O_2156,N_19796,N_19755);
nor UO_2157 (O_2157,N_19918,N_19944);
or UO_2158 (O_2158,N_19824,N_19945);
or UO_2159 (O_2159,N_19877,N_19844);
and UO_2160 (O_2160,N_19832,N_19843);
or UO_2161 (O_2161,N_19775,N_19839);
and UO_2162 (O_2162,N_19990,N_19924);
nor UO_2163 (O_2163,N_19913,N_19852);
nand UO_2164 (O_2164,N_19851,N_19800);
and UO_2165 (O_2165,N_19790,N_19931);
xnor UO_2166 (O_2166,N_19811,N_19894);
nor UO_2167 (O_2167,N_19908,N_19927);
nand UO_2168 (O_2168,N_19771,N_19950);
and UO_2169 (O_2169,N_19900,N_19957);
or UO_2170 (O_2170,N_19968,N_19931);
nand UO_2171 (O_2171,N_19891,N_19780);
xor UO_2172 (O_2172,N_19872,N_19782);
or UO_2173 (O_2173,N_19885,N_19900);
nor UO_2174 (O_2174,N_19838,N_19886);
nand UO_2175 (O_2175,N_19872,N_19817);
nand UO_2176 (O_2176,N_19846,N_19944);
xnor UO_2177 (O_2177,N_19991,N_19959);
xor UO_2178 (O_2178,N_19947,N_19997);
and UO_2179 (O_2179,N_19957,N_19756);
nand UO_2180 (O_2180,N_19945,N_19861);
nand UO_2181 (O_2181,N_19936,N_19911);
xor UO_2182 (O_2182,N_19842,N_19948);
xnor UO_2183 (O_2183,N_19848,N_19759);
or UO_2184 (O_2184,N_19788,N_19848);
and UO_2185 (O_2185,N_19780,N_19839);
and UO_2186 (O_2186,N_19846,N_19816);
or UO_2187 (O_2187,N_19823,N_19843);
nand UO_2188 (O_2188,N_19813,N_19875);
nand UO_2189 (O_2189,N_19929,N_19775);
and UO_2190 (O_2190,N_19771,N_19935);
nand UO_2191 (O_2191,N_19769,N_19867);
and UO_2192 (O_2192,N_19825,N_19928);
nand UO_2193 (O_2193,N_19945,N_19920);
nor UO_2194 (O_2194,N_19917,N_19935);
and UO_2195 (O_2195,N_19879,N_19997);
or UO_2196 (O_2196,N_19846,N_19768);
xnor UO_2197 (O_2197,N_19969,N_19772);
xor UO_2198 (O_2198,N_19809,N_19993);
nor UO_2199 (O_2199,N_19860,N_19805);
xor UO_2200 (O_2200,N_19829,N_19913);
nor UO_2201 (O_2201,N_19756,N_19992);
or UO_2202 (O_2202,N_19802,N_19919);
nor UO_2203 (O_2203,N_19800,N_19931);
nand UO_2204 (O_2204,N_19897,N_19759);
nor UO_2205 (O_2205,N_19764,N_19962);
nor UO_2206 (O_2206,N_19986,N_19943);
xnor UO_2207 (O_2207,N_19983,N_19923);
xnor UO_2208 (O_2208,N_19990,N_19985);
nor UO_2209 (O_2209,N_19927,N_19833);
nand UO_2210 (O_2210,N_19915,N_19945);
xor UO_2211 (O_2211,N_19820,N_19824);
or UO_2212 (O_2212,N_19950,N_19891);
xnor UO_2213 (O_2213,N_19882,N_19915);
or UO_2214 (O_2214,N_19844,N_19823);
nand UO_2215 (O_2215,N_19975,N_19806);
nor UO_2216 (O_2216,N_19894,N_19962);
nand UO_2217 (O_2217,N_19976,N_19934);
or UO_2218 (O_2218,N_19840,N_19776);
or UO_2219 (O_2219,N_19874,N_19846);
or UO_2220 (O_2220,N_19893,N_19935);
xor UO_2221 (O_2221,N_19799,N_19855);
or UO_2222 (O_2222,N_19923,N_19919);
xor UO_2223 (O_2223,N_19913,N_19872);
or UO_2224 (O_2224,N_19923,N_19884);
or UO_2225 (O_2225,N_19907,N_19781);
and UO_2226 (O_2226,N_19819,N_19873);
and UO_2227 (O_2227,N_19982,N_19804);
or UO_2228 (O_2228,N_19985,N_19901);
xor UO_2229 (O_2229,N_19988,N_19828);
and UO_2230 (O_2230,N_19927,N_19803);
nand UO_2231 (O_2231,N_19839,N_19896);
nand UO_2232 (O_2232,N_19880,N_19966);
or UO_2233 (O_2233,N_19956,N_19939);
nor UO_2234 (O_2234,N_19929,N_19939);
xor UO_2235 (O_2235,N_19796,N_19829);
and UO_2236 (O_2236,N_19873,N_19758);
nand UO_2237 (O_2237,N_19963,N_19868);
and UO_2238 (O_2238,N_19976,N_19894);
nand UO_2239 (O_2239,N_19802,N_19835);
xor UO_2240 (O_2240,N_19997,N_19783);
and UO_2241 (O_2241,N_19810,N_19989);
or UO_2242 (O_2242,N_19772,N_19816);
nand UO_2243 (O_2243,N_19899,N_19761);
nand UO_2244 (O_2244,N_19958,N_19862);
nand UO_2245 (O_2245,N_19793,N_19881);
or UO_2246 (O_2246,N_19897,N_19831);
nand UO_2247 (O_2247,N_19761,N_19872);
nor UO_2248 (O_2248,N_19967,N_19806);
nand UO_2249 (O_2249,N_19812,N_19844);
xnor UO_2250 (O_2250,N_19856,N_19998);
nor UO_2251 (O_2251,N_19862,N_19756);
xor UO_2252 (O_2252,N_19951,N_19959);
xnor UO_2253 (O_2253,N_19937,N_19916);
nand UO_2254 (O_2254,N_19995,N_19820);
nor UO_2255 (O_2255,N_19967,N_19968);
and UO_2256 (O_2256,N_19849,N_19961);
xor UO_2257 (O_2257,N_19775,N_19948);
nand UO_2258 (O_2258,N_19990,N_19959);
nand UO_2259 (O_2259,N_19789,N_19839);
nor UO_2260 (O_2260,N_19831,N_19978);
and UO_2261 (O_2261,N_19997,N_19770);
xnor UO_2262 (O_2262,N_19773,N_19901);
nand UO_2263 (O_2263,N_19783,N_19926);
xnor UO_2264 (O_2264,N_19752,N_19784);
nand UO_2265 (O_2265,N_19763,N_19768);
xor UO_2266 (O_2266,N_19970,N_19847);
xnor UO_2267 (O_2267,N_19819,N_19965);
xor UO_2268 (O_2268,N_19793,N_19868);
nor UO_2269 (O_2269,N_19770,N_19874);
or UO_2270 (O_2270,N_19990,N_19875);
nor UO_2271 (O_2271,N_19925,N_19862);
nand UO_2272 (O_2272,N_19952,N_19818);
or UO_2273 (O_2273,N_19786,N_19837);
or UO_2274 (O_2274,N_19752,N_19958);
nand UO_2275 (O_2275,N_19778,N_19958);
or UO_2276 (O_2276,N_19942,N_19966);
or UO_2277 (O_2277,N_19978,N_19966);
and UO_2278 (O_2278,N_19859,N_19948);
or UO_2279 (O_2279,N_19905,N_19858);
or UO_2280 (O_2280,N_19959,N_19806);
xnor UO_2281 (O_2281,N_19758,N_19851);
and UO_2282 (O_2282,N_19871,N_19872);
nor UO_2283 (O_2283,N_19965,N_19938);
and UO_2284 (O_2284,N_19812,N_19981);
xnor UO_2285 (O_2285,N_19777,N_19852);
and UO_2286 (O_2286,N_19768,N_19914);
nor UO_2287 (O_2287,N_19805,N_19796);
nor UO_2288 (O_2288,N_19879,N_19959);
nor UO_2289 (O_2289,N_19874,N_19947);
or UO_2290 (O_2290,N_19967,N_19916);
nor UO_2291 (O_2291,N_19830,N_19948);
nand UO_2292 (O_2292,N_19897,N_19809);
nand UO_2293 (O_2293,N_19889,N_19890);
and UO_2294 (O_2294,N_19977,N_19950);
xor UO_2295 (O_2295,N_19897,N_19861);
or UO_2296 (O_2296,N_19808,N_19771);
nor UO_2297 (O_2297,N_19783,N_19799);
nor UO_2298 (O_2298,N_19929,N_19964);
or UO_2299 (O_2299,N_19995,N_19939);
xnor UO_2300 (O_2300,N_19906,N_19908);
nand UO_2301 (O_2301,N_19898,N_19989);
and UO_2302 (O_2302,N_19915,N_19847);
nor UO_2303 (O_2303,N_19993,N_19847);
nand UO_2304 (O_2304,N_19775,N_19849);
xnor UO_2305 (O_2305,N_19939,N_19833);
and UO_2306 (O_2306,N_19803,N_19795);
nor UO_2307 (O_2307,N_19890,N_19808);
nand UO_2308 (O_2308,N_19982,N_19803);
nand UO_2309 (O_2309,N_19966,N_19885);
nand UO_2310 (O_2310,N_19752,N_19766);
nand UO_2311 (O_2311,N_19959,N_19869);
nor UO_2312 (O_2312,N_19968,N_19947);
nor UO_2313 (O_2313,N_19931,N_19918);
xnor UO_2314 (O_2314,N_19926,N_19795);
or UO_2315 (O_2315,N_19848,N_19999);
or UO_2316 (O_2316,N_19982,N_19940);
nor UO_2317 (O_2317,N_19785,N_19973);
nor UO_2318 (O_2318,N_19996,N_19895);
nand UO_2319 (O_2319,N_19997,N_19796);
nand UO_2320 (O_2320,N_19824,N_19963);
and UO_2321 (O_2321,N_19779,N_19987);
and UO_2322 (O_2322,N_19812,N_19913);
and UO_2323 (O_2323,N_19768,N_19842);
or UO_2324 (O_2324,N_19970,N_19778);
xnor UO_2325 (O_2325,N_19821,N_19884);
nor UO_2326 (O_2326,N_19787,N_19962);
xor UO_2327 (O_2327,N_19941,N_19955);
or UO_2328 (O_2328,N_19880,N_19965);
nand UO_2329 (O_2329,N_19842,N_19955);
and UO_2330 (O_2330,N_19853,N_19963);
nor UO_2331 (O_2331,N_19774,N_19828);
xnor UO_2332 (O_2332,N_19791,N_19925);
nor UO_2333 (O_2333,N_19958,N_19764);
or UO_2334 (O_2334,N_19867,N_19763);
xnor UO_2335 (O_2335,N_19891,N_19932);
and UO_2336 (O_2336,N_19914,N_19824);
or UO_2337 (O_2337,N_19782,N_19986);
or UO_2338 (O_2338,N_19788,N_19780);
or UO_2339 (O_2339,N_19876,N_19766);
xnor UO_2340 (O_2340,N_19779,N_19751);
nand UO_2341 (O_2341,N_19856,N_19962);
or UO_2342 (O_2342,N_19838,N_19863);
nand UO_2343 (O_2343,N_19779,N_19939);
xor UO_2344 (O_2344,N_19896,N_19774);
nand UO_2345 (O_2345,N_19862,N_19795);
nor UO_2346 (O_2346,N_19880,N_19881);
and UO_2347 (O_2347,N_19858,N_19945);
nor UO_2348 (O_2348,N_19832,N_19933);
xor UO_2349 (O_2349,N_19813,N_19760);
xor UO_2350 (O_2350,N_19764,N_19944);
nand UO_2351 (O_2351,N_19879,N_19779);
or UO_2352 (O_2352,N_19802,N_19886);
nand UO_2353 (O_2353,N_19862,N_19847);
or UO_2354 (O_2354,N_19986,N_19806);
nand UO_2355 (O_2355,N_19906,N_19865);
xnor UO_2356 (O_2356,N_19834,N_19948);
nand UO_2357 (O_2357,N_19806,N_19848);
nor UO_2358 (O_2358,N_19800,N_19831);
and UO_2359 (O_2359,N_19885,N_19929);
nor UO_2360 (O_2360,N_19836,N_19975);
nor UO_2361 (O_2361,N_19826,N_19948);
xor UO_2362 (O_2362,N_19842,N_19897);
nand UO_2363 (O_2363,N_19859,N_19904);
xor UO_2364 (O_2364,N_19934,N_19848);
and UO_2365 (O_2365,N_19820,N_19978);
nor UO_2366 (O_2366,N_19990,N_19763);
nand UO_2367 (O_2367,N_19788,N_19945);
xor UO_2368 (O_2368,N_19851,N_19801);
nor UO_2369 (O_2369,N_19881,N_19846);
nor UO_2370 (O_2370,N_19810,N_19962);
nand UO_2371 (O_2371,N_19782,N_19985);
or UO_2372 (O_2372,N_19826,N_19821);
or UO_2373 (O_2373,N_19964,N_19975);
xor UO_2374 (O_2374,N_19766,N_19871);
and UO_2375 (O_2375,N_19788,N_19977);
nand UO_2376 (O_2376,N_19912,N_19818);
and UO_2377 (O_2377,N_19805,N_19846);
and UO_2378 (O_2378,N_19914,N_19894);
nand UO_2379 (O_2379,N_19989,N_19763);
nand UO_2380 (O_2380,N_19821,N_19827);
and UO_2381 (O_2381,N_19893,N_19943);
or UO_2382 (O_2382,N_19769,N_19894);
and UO_2383 (O_2383,N_19950,N_19999);
and UO_2384 (O_2384,N_19802,N_19905);
or UO_2385 (O_2385,N_19780,N_19870);
or UO_2386 (O_2386,N_19933,N_19978);
nor UO_2387 (O_2387,N_19996,N_19757);
and UO_2388 (O_2388,N_19765,N_19896);
nand UO_2389 (O_2389,N_19810,N_19795);
nand UO_2390 (O_2390,N_19768,N_19862);
nor UO_2391 (O_2391,N_19831,N_19882);
nand UO_2392 (O_2392,N_19840,N_19844);
xnor UO_2393 (O_2393,N_19862,N_19889);
nor UO_2394 (O_2394,N_19750,N_19905);
and UO_2395 (O_2395,N_19790,N_19798);
nor UO_2396 (O_2396,N_19990,N_19832);
nor UO_2397 (O_2397,N_19820,N_19811);
nor UO_2398 (O_2398,N_19942,N_19949);
nor UO_2399 (O_2399,N_19857,N_19990);
nand UO_2400 (O_2400,N_19975,N_19791);
or UO_2401 (O_2401,N_19837,N_19810);
and UO_2402 (O_2402,N_19765,N_19886);
xor UO_2403 (O_2403,N_19961,N_19836);
xor UO_2404 (O_2404,N_19899,N_19932);
xor UO_2405 (O_2405,N_19992,N_19811);
and UO_2406 (O_2406,N_19753,N_19853);
nand UO_2407 (O_2407,N_19983,N_19769);
or UO_2408 (O_2408,N_19927,N_19906);
nor UO_2409 (O_2409,N_19802,N_19853);
or UO_2410 (O_2410,N_19841,N_19836);
xnor UO_2411 (O_2411,N_19829,N_19956);
nor UO_2412 (O_2412,N_19973,N_19767);
nand UO_2413 (O_2413,N_19998,N_19927);
and UO_2414 (O_2414,N_19815,N_19950);
nand UO_2415 (O_2415,N_19848,N_19785);
xnor UO_2416 (O_2416,N_19817,N_19951);
nand UO_2417 (O_2417,N_19760,N_19927);
nor UO_2418 (O_2418,N_19804,N_19944);
or UO_2419 (O_2419,N_19887,N_19851);
nor UO_2420 (O_2420,N_19973,N_19814);
nand UO_2421 (O_2421,N_19971,N_19999);
xor UO_2422 (O_2422,N_19962,N_19954);
nor UO_2423 (O_2423,N_19802,N_19926);
xnor UO_2424 (O_2424,N_19879,N_19814);
or UO_2425 (O_2425,N_19795,N_19846);
or UO_2426 (O_2426,N_19861,N_19830);
xor UO_2427 (O_2427,N_19893,N_19853);
and UO_2428 (O_2428,N_19975,N_19797);
nand UO_2429 (O_2429,N_19786,N_19950);
nand UO_2430 (O_2430,N_19975,N_19787);
and UO_2431 (O_2431,N_19763,N_19988);
xor UO_2432 (O_2432,N_19938,N_19832);
and UO_2433 (O_2433,N_19772,N_19948);
or UO_2434 (O_2434,N_19762,N_19760);
or UO_2435 (O_2435,N_19937,N_19884);
xor UO_2436 (O_2436,N_19800,N_19753);
or UO_2437 (O_2437,N_19880,N_19894);
nand UO_2438 (O_2438,N_19825,N_19990);
xor UO_2439 (O_2439,N_19937,N_19883);
and UO_2440 (O_2440,N_19829,N_19811);
nand UO_2441 (O_2441,N_19831,N_19877);
or UO_2442 (O_2442,N_19898,N_19920);
nor UO_2443 (O_2443,N_19936,N_19774);
nor UO_2444 (O_2444,N_19971,N_19902);
xnor UO_2445 (O_2445,N_19842,N_19934);
xnor UO_2446 (O_2446,N_19787,N_19927);
xnor UO_2447 (O_2447,N_19846,N_19757);
or UO_2448 (O_2448,N_19795,N_19895);
nor UO_2449 (O_2449,N_19930,N_19946);
and UO_2450 (O_2450,N_19820,N_19994);
nand UO_2451 (O_2451,N_19882,N_19962);
or UO_2452 (O_2452,N_19989,N_19882);
and UO_2453 (O_2453,N_19877,N_19851);
and UO_2454 (O_2454,N_19847,N_19990);
and UO_2455 (O_2455,N_19875,N_19767);
and UO_2456 (O_2456,N_19788,N_19964);
or UO_2457 (O_2457,N_19825,N_19889);
or UO_2458 (O_2458,N_19973,N_19871);
nor UO_2459 (O_2459,N_19983,N_19797);
and UO_2460 (O_2460,N_19751,N_19965);
xnor UO_2461 (O_2461,N_19955,N_19961);
or UO_2462 (O_2462,N_19765,N_19857);
and UO_2463 (O_2463,N_19989,N_19798);
nand UO_2464 (O_2464,N_19890,N_19966);
nor UO_2465 (O_2465,N_19894,N_19998);
nand UO_2466 (O_2466,N_19883,N_19880);
and UO_2467 (O_2467,N_19750,N_19921);
or UO_2468 (O_2468,N_19848,N_19816);
or UO_2469 (O_2469,N_19904,N_19849);
nand UO_2470 (O_2470,N_19921,N_19755);
or UO_2471 (O_2471,N_19986,N_19880);
xor UO_2472 (O_2472,N_19884,N_19998);
nand UO_2473 (O_2473,N_19772,N_19884);
nand UO_2474 (O_2474,N_19863,N_19852);
xnor UO_2475 (O_2475,N_19788,N_19905);
nand UO_2476 (O_2476,N_19765,N_19867);
or UO_2477 (O_2477,N_19926,N_19956);
or UO_2478 (O_2478,N_19894,N_19759);
and UO_2479 (O_2479,N_19813,N_19951);
nand UO_2480 (O_2480,N_19830,N_19908);
or UO_2481 (O_2481,N_19891,N_19847);
or UO_2482 (O_2482,N_19751,N_19949);
xor UO_2483 (O_2483,N_19868,N_19792);
xor UO_2484 (O_2484,N_19991,N_19867);
xor UO_2485 (O_2485,N_19851,N_19815);
and UO_2486 (O_2486,N_19994,N_19780);
or UO_2487 (O_2487,N_19828,N_19771);
nand UO_2488 (O_2488,N_19870,N_19752);
or UO_2489 (O_2489,N_19840,N_19849);
xnor UO_2490 (O_2490,N_19954,N_19783);
nor UO_2491 (O_2491,N_19944,N_19888);
or UO_2492 (O_2492,N_19864,N_19802);
and UO_2493 (O_2493,N_19972,N_19789);
xnor UO_2494 (O_2494,N_19768,N_19993);
xnor UO_2495 (O_2495,N_19858,N_19994);
nor UO_2496 (O_2496,N_19813,N_19852);
or UO_2497 (O_2497,N_19923,N_19811);
nand UO_2498 (O_2498,N_19925,N_19799);
or UO_2499 (O_2499,N_19799,N_19898);
endmodule