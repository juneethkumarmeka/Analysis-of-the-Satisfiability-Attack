module basic_500_3000_500_50_levels_10xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_106,In_18);
xnor U1 (N_1,In_425,In_240);
and U2 (N_2,In_144,In_377);
nor U3 (N_3,In_451,In_209);
nor U4 (N_4,In_66,In_181);
or U5 (N_5,In_338,In_271);
and U6 (N_6,In_252,In_440);
and U7 (N_7,In_41,In_237);
nor U8 (N_8,In_488,In_413);
and U9 (N_9,In_398,In_459);
xor U10 (N_10,In_169,In_487);
and U11 (N_11,In_184,In_369);
or U12 (N_12,In_37,In_311);
or U13 (N_13,In_485,In_443);
nor U14 (N_14,In_185,In_227);
or U15 (N_15,In_287,In_415);
and U16 (N_16,In_140,In_126);
xor U17 (N_17,In_216,In_180);
and U18 (N_18,In_420,In_94);
or U19 (N_19,In_375,In_177);
nor U20 (N_20,In_82,In_78);
nand U21 (N_21,In_238,In_173);
nand U22 (N_22,In_176,In_59);
nor U23 (N_23,In_444,In_164);
xnor U24 (N_24,In_42,In_482);
nand U25 (N_25,In_125,In_339);
xnor U26 (N_26,In_153,In_360);
or U27 (N_27,In_283,In_333);
and U28 (N_28,In_308,In_151);
or U29 (N_29,In_291,In_496);
nor U30 (N_30,In_53,In_267);
nor U31 (N_31,In_405,In_170);
or U32 (N_32,In_152,In_46);
or U33 (N_33,In_417,In_474);
nand U34 (N_34,In_211,In_92);
or U35 (N_35,In_162,In_483);
nand U36 (N_36,In_435,In_86);
and U37 (N_37,In_19,In_93);
and U38 (N_38,In_378,In_313);
xor U39 (N_39,In_103,In_498);
or U40 (N_40,In_77,In_255);
xor U41 (N_41,In_147,In_62);
and U42 (N_42,In_288,In_432);
or U43 (N_43,In_163,In_139);
and U44 (N_44,In_4,In_193);
xnor U45 (N_45,In_296,In_161);
and U46 (N_46,In_463,In_275);
nor U47 (N_47,In_259,In_225);
xnor U48 (N_48,In_118,In_71);
xor U49 (N_49,In_131,In_454);
nor U50 (N_50,In_129,In_198);
or U51 (N_51,In_457,In_402);
and U52 (N_52,In_316,In_433);
nand U53 (N_53,In_212,In_309);
nand U54 (N_54,In_69,In_419);
or U55 (N_55,In_335,In_245);
or U56 (N_56,In_494,In_351);
or U57 (N_57,In_325,In_328);
or U58 (N_58,In_290,In_213);
xnor U59 (N_59,In_88,In_136);
and U60 (N_60,In_90,In_421);
or U61 (N_61,In_124,In_231);
nor U62 (N_62,In_386,N_18);
nand U63 (N_63,In_430,In_358);
nor U64 (N_64,In_257,In_6);
nor U65 (N_65,In_95,In_9);
nor U66 (N_66,In_422,In_354);
nand U67 (N_67,N_19,In_168);
nand U68 (N_68,In_251,N_9);
nor U69 (N_69,In_426,In_171);
or U70 (N_70,In_280,N_6);
or U71 (N_71,In_408,In_324);
nand U72 (N_72,In_320,In_84);
nor U73 (N_73,In_337,In_206);
nor U74 (N_74,In_13,In_166);
nor U75 (N_75,In_133,In_76);
and U76 (N_76,N_14,In_22);
nand U77 (N_77,In_138,In_182);
nor U78 (N_78,In_74,N_46);
and U79 (N_79,In_465,In_468);
or U80 (N_80,N_37,In_391);
xnor U81 (N_81,In_233,In_8);
nand U82 (N_82,In_380,In_72);
xnor U83 (N_83,In_201,N_50);
nand U84 (N_84,In_146,In_300);
or U85 (N_85,N_34,In_302);
nand U86 (N_86,N_52,In_410);
or U87 (N_87,N_44,In_197);
and U88 (N_88,In_384,In_160);
and U89 (N_89,N_38,In_7);
xnor U90 (N_90,In_449,In_109);
and U91 (N_91,In_347,In_21);
nand U92 (N_92,N_54,In_349);
nand U93 (N_93,In_295,In_330);
nor U94 (N_94,In_98,In_234);
nand U95 (N_95,In_471,In_149);
xnor U96 (N_96,In_230,N_28);
nand U97 (N_97,In_248,In_148);
nor U98 (N_98,In_190,In_228);
and U99 (N_99,N_2,In_246);
nand U100 (N_100,N_56,In_481);
nor U101 (N_101,In_381,In_269);
or U102 (N_102,In_47,N_24);
nor U103 (N_103,In_108,In_478);
nor U104 (N_104,In_205,In_236);
or U105 (N_105,In_458,In_141);
and U106 (N_106,In_279,N_11);
and U107 (N_107,In_376,In_15);
and U108 (N_108,In_429,In_235);
and U109 (N_109,In_194,In_355);
or U110 (N_110,In_464,In_16);
nor U111 (N_111,In_242,In_50);
xor U112 (N_112,In_452,N_16);
and U113 (N_113,In_127,In_31);
or U114 (N_114,In_442,In_107);
nor U115 (N_115,In_24,In_29);
nand U116 (N_116,In_495,In_493);
xnor U117 (N_117,In_25,In_155);
nor U118 (N_118,In_396,In_286);
and U119 (N_119,In_484,In_373);
and U120 (N_120,N_1,N_116);
xnor U121 (N_121,In_315,In_489);
nand U122 (N_122,N_17,N_55);
and U123 (N_123,In_322,In_145);
nand U124 (N_124,N_33,N_114);
xor U125 (N_125,In_407,In_289);
nor U126 (N_126,In_120,In_218);
nand U127 (N_127,In_219,N_101);
nand U128 (N_128,N_25,In_423);
xor U129 (N_129,In_307,In_401);
and U130 (N_130,In_75,N_92);
or U131 (N_131,In_412,N_59);
and U132 (N_132,In_249,N_5);
nor U133 (N_133,In_297,In_264);
and U134 (N_134,N_76,In_359);
nand U135 (N_135,In_350,In_363);
nand U136 (N_136,In_438,In_372);
and U137 (N_137,In_111,N_10);
xnor U138 (N_138,N_51,In_154);
xor U139 (N_139,In_208,N_3);
xnor U140 (N_140,N_78,In_312);
and U141 (N_141,In_281,In_199);
xor U142 (N_142,N_96,N_15);
or U143 (N_143,In_374,In_310);
nand U144 (N_144,In_117,In_477);
xnor U145 (N_145,In_250,In_305);
nor U146 (N_146,In_357,In_390);
or U147 (N_147,In_48,In_455);
or U148 (N_148,In_214,In_273);
or U149 (N_149,In_2,N_27);
nand U150 (N_150,In_187,In_301);
and U151 (N_151,In_368,N_64);
nor U152 (N_152,In_314,N_0);
and U153 (N_153,In_96,In_292);
and U154 (N_154,In_370,In_244);
nor U155 (N_155,N_35,N_49);
or U156 (N_156,N_32,In_165);
or U157 (N_157,In_110,In_323);
nand U158 (N_158,In_30,In_456);
nand U159 (N_159,In_473,N_74);
nand U160 (N_160,In_352,In_55);
nor U161 (N_161,In_121,N_86);
and U162 (N_162,In_1,In_32);
xor U163 (N_163,N_36,In_362);
or U164 (N_164,In_61,In_348);
and U165 (N_165,In_183,In_116);
and U166 (N_166,In_89,In_33);
xor U167 (N_167,In_416,N_119);
nand U168 (N_168,In_14,N_39);
nor U169 (N_169,In_476,In_132);
xor U170 (N_170,In_393,N_69);
and U171 (N_171,In_65,In_434);
and U172 (N_172,N_70,N_113);
and U173 (N_173,N_106,In_353);
nor U174 (N_174,N_93,In_23);
xnor U175 (N_175,In_278,In_397);
nand U176 (N_176,In_406,N_66);
nand U177 (N_177,In_203,N_109);
nor U178 (N_178,In_293,N_26);
or U179 (N_179,In_399,In_56);
or U180 (N_180,In_27,N_80);
or U181 (N_181,In_467,In_331);
nand U182 (N_182,In_39,In_365);
nor U183 (N_183,In_207,In_400);
nand U184 (N_184,In_491,In_446);
nor U185 (N_185,In_385,In_122);
or U186 (N_186,N_68,In_441);
xor U187 (N_187,In_51,In_43);
and U188 (N_188,N_47,In_26);
or U189 (N_189,N_84,In_298);
and U190 (N_190,In_388,In_261);
xnor U191 (N_191,In_263,N_82);
nor U192 (N_192,In_67,N_81);
or U193 (N_193,N_30,In_174);
xnor U194 (N_194,N_179,In_63);
nor U195 (N_195,N_139,N_79);
and U196 (N_196,N_145,N_177);
or U197 (N_197,N_159,In_445);
nor U198 (N_198,In_5,N_171);
nand U199 (N_199,N_152,In_99);
nand U200 (N_200,In_58,In_189);
xnor U201 (N_201,In_270,In_364);
xnor U202 (N_202,In_226,N_136);
and U203 (N_203,N_20,In_394);
and U204 (N_204,In_191,N_130);
or U205 (N_205,N_176,In_395);
nor U206 (N_206,N_48,N_88);
and U207 (N_207,In_159,N_149);
nand U208 (N_208,N_110,N_129);
nand U209 (N_209,N_123,In_475);
nor U210 (N_210,In_10,In_427);
xnor U211 (N_211,N_57,In_130);
nand U212 (N_212,In_262,N_61);
or U213 (N_213,In_253,In_276);
nand U214 (N_214,In_192,In_389);
and U215 (N_215,In_303,In_424);
nor U216 (N_216,In_340,In_461);
nor U217 (N_217,In_178,N_22);
and U218 (N_218,In_260,N_175);
xnor U219 (N_219,In_210,N_140);
or U220 (N_220,In_480,In_327);
and U221 (N_221,In_460,N_168);
nor U222 (N_222,N_65,N_107);
nor U223 (N_223,In_128,N_98);
nor U224 (N_224,In_97,N_156);
xor U225 (N_225,In_17,N_83);
nor U226 (N_226,In_382,In_284);
nand U227 (N_227,N_103,In_254);
nand U228 (N_228,N_141,In_490);
nor U229 (N_229,In_68,N_146);
nor U230 (N_230,In_418,In_479);
nor U231 (N_231,N_142,In_11);
xor U232 (N_232,In_486,In_414);
and U233 (N_233,N_100,In_470);
or U234 (N_234,In_239,N_178);
and U235 (N_235,N_165,In_285);
or U236 (N_236,N_148,N_164);
xnor U237 (N_237,In_204,In_341);
and U238 (N_238,In_115,In_448);
and U239 (N_239,N_121,In_268);
or U240 (N_240,In_258,N_181);
xor U241 (N_241,N_95,N_134);
nand U242 (N_242,In_3,In_83);
nand U243 (N_243,N_173,In_157);
nand U244 (N_244,N_132,N_194);
nand U245 (N_245,N_161,N_232);
nor U246 (N_246,N_126,In_217);
or U247 (N_247,In_453,N_208);
xnor U248 (N_248,In_344,N_238);
or U249 (N_249,N_43,N_236);
nor U250 (N_250,N_205,In_243);
or U251 (N_251,N_185,In_64);
nand U252 (N_252,N_163,N_45);
or U253 (N_253,In_57,N_206);
and U254 (N_254,In_366,In_272);
or U255 (N_255,N_231,In_326);
and U256 (N_256,N_118,N_157);
xor U257 (N_257,In_143,In_105);
xnor U258 (N_258,In_345,N_224);
nand U259 (N_259,In_342,N_180);
nor U260 (N_260,N_125,N_99);
nor U261 (N_261,In_80,N_172);
xnor U262 (N_262,In_437,N_214);
and U263 (N_263,In_403,N_202);
and U264 (N_264,N_200,In_202);
or U265 (N_265,In_79,In_195);
or U266 (N_266,N_135,In_38);
or U267 (N_267,N_225,N_31);
or U268 (N_268,In_241,In_222);
nor U269 (N_269,In_232,In_229);
or U270 (N_270,N_216,In_404);
xnor U271 (N_271,In_220,N_144);
and U272 (N_272,In_492,In_35);
nand U273 (N_273,N_23,N_62);
nand U274 (N_274,In_436,In_361);
and U275 (N_275,N_160,In_167);
xor U276 (N_276,In_28,In_100);
and U277 (N_277,N_234,In_34);
and U278 (N_278,In_294,N_230);
nor U279 (N_279,In_114,N_89);
nand U280 (N_280,In_497,In_45);
xnor U281 (N_281,N_21,In_306);
nand U282 (N_282,N_193,N_184);
and U283 (N_283,N_108,In_134);
nand U284 (N_284,In_142,N_63);
and U285 (N_285,N_29,In_299);
xor U286 (N_286,N_186,N_115);
nand U287 (N_287,In_112,N_218);
nor U288 (N_288,N_67,N_209);
nor U289 (N_289,N_182,In_265);
nor U290 (N_290,In_367,N_12);
nor U291 (N_291,N_169,N_195);
xor U292 (N_292,N_167,N_147);
xor U293 (N_293,In_274,N_75);
nor U294 (N_294,N_154,N_138);
nand U295 (N_295,In_472,N_150);
or U296 (N_296,N_207,N_41);
nand U297 (N_297,N_220,N_90);
or U298 (N_298,N_151,In_371);
and U299 (N_299,In_73,In_462);
nor U300 (N_300,N_77,N_155);
xnor U301 (N_301,N_124,N_245);
and U302 (N_302,N_223,N_131);
and U303 (N_303,N_263,N_127);
nand U304 (N_304,In_36,In_20);
or U305 (N_305,N_274,In_81);
or U306 (N_306,N_85,N_192);
or U307 (N_307,N_247,N_265);
nor U308 (N_308,In_196,In_186);
nor U309 (N_309,N_275,N_128);
or U310 (N_310,N_253,N_286);
nand U311 (N_311,N_276,N_111);
and U312 (N_312,N_278,N_246);
or U313 (N_313,N_122,N_273);
nand U314 (N_314,N_187,N_281);
xor U315 (N_315,N_120,N_213);
or U316 (N_316,N_174,N_4);
xor U317 (N_317,N_211,In_317);
nand U318 (N_318,N_117,N_229);
and U319 (N_319,N_269,N_191);
or U320 (N_320,In_156,N_296);
xnor U321 (N_321,N_284,In_336);
nand U322 (N_322,N_133,N_219);
and U323 (N_323,In_304,In_392);
nand U324 (N_324,N_162,In_119);
and U325 (N_325,N_7,N_257);
xnor U326 (N_326,N_248,In_60);
xor U327 (N_327,N_261,In_188);
nand U328 (N_328,N_270,In_334);
nand U329 (N_329,N_102,In_379);
nand U330 (N_330,In_0,N_203);
and U331 (N_331,In_282,N_268);
and U332 (N_332,N_292,N_239);
or U333 (N_333,N_215,N_58);
nor U334 (N_334,N_251,N_104);
xor U335 (N_335,In_450,N_143);
or U336 (N_336,N_241,N_183);
nor U337 (N_337,N_280,In_224);
nor U338 (N_338,N_264,In_256);
nand U339 (N_339,N_237,In_409);
nor U340 (N_340,N_272,In_49);
nor U341 (N_341,In_356,N_198);
and U342 (N_342,In_150,In_215);
nor U343 (N_343,In_266,In_135);
nand U344 (N_344,N_94,In_319);
or U345 (N_345,N_294,In_466);
xnor U346 (N_346,N_40,N_266);
nand U347 (N_347,N_196,In_346);
xnor U348 (N_348,N_290,N_262);
and U349 (N_349,N_199,N_8);
and U350 (N_350,N_244,N_267);
xnor U351 (N_351,N_293,N_242);
nor U352 (N_352,In_104,In_102);
or U353 (N_353,N_71,N_217);
or U354 (N_354,N_227,In_137);
nor U355 (N_355,N_42,N_258);
or U356 (N_356,N_256,In_85);
nand U357 (N_357,In_221,N_105);
xor U358 (N_358,N_299,In_332);
xnor U359 (N_359,N_279,N_73);
or U360 (N_360,N_307,N_255);
xor U361 (N_361,N_235,N_359);
nor U362 (N_362,In_158,N_332);
or U363 (N_363,N_228,In_70);
xnor U364 (N_364,N_112,N_166);
nor U365 (N_365,N_13,N_303);
nor U366 (N_366,N_356,In_383);
xnor U367 (N_367,N_226,N_344);
nand U368 (N_368,N_158,N_295);
nand U369 (N_369,N_324,N_333);
nor U370 (N_370,N_188,N_327);
xor U371 (N_371,N_323,N_249);
nor U372 (N_372,In_12,N_283);
and U373 (N_373,N_325,N_310);
or U374 (N_374,N_354,N_358);
nor U375 (N_375,In_175,N_210);
nand U376 (N_376,N_301,N_282);
nand U377 (N_377,N_331,In_200);
or U378 (N_378,N_316,N_319);
nand U379 (N_379,In_329,N_170);
or U380 (N_380,N_346,In_87);
xor U381 (N_381,N_352,In_223);
xnor U382 (N_382,N_201,N_351);
nand U383 (N_383,N_338,In_447);
nand U384 (N_384,N_309,N_254);
xor U385 (N_385,N_342,N_243);
nand U386 (N_386,N_322,In_123);
or U387 (N_387,N_302,N_277);
nand U388 (N_388,N_91,N_60);
nor U389 (N_389,N_311,N_212);
nand U390 (N_390,N_330,N_259);
or U391 (N_391,N_321,In_113);
or U392 (N_392,In_321,N_314);
nor U393 (N_393,N_300,In_343);
nand U394 (N_394,N_313,In_277);
and U395 (N_395,N_328,N_347);
or U396 (N_396,N_304,N_87);
nand U397 (N_397,N_287,In_40);
xor U398 (N_398,N_345,In_44);
xor U399 (N_399,N_298,N_240);
and U400 (N_400,In_91,N_339);
nor U401 (N_401,In_431,N_349);
nor U402 (N_402,In_318,N_355);
nand U403 (N_403,N_297,N_197);
and U404 (N_404,N_271,N_53);
or U405 (N_405,N_289,In_428);
and U406 (N_406,In_469,In_101);
or U407 (N_407,N_353,N_336);
and U408 (N_408,N_317,N_326);
xnor U409 (N_409,N_72,N_348);
nor U410 (N_410,N_340,In_179);
nor U411 (N_411,N_341,N_204);
and U412 (N_412,N_320,N_335);
xor U413 (N_413,N_343,N_189);
and U414 (N_414,N_222,In_54);
xor U415 (N_415,N_250,In_499);
xor U416 (N_416,N_308,In_172);
nor U417 (N_417,N_315,In_52);
nor U418 (N_418,In_387,N_291);
nand U419 (N_419,N_252,N_334);
or U420 (N_420,N_412,In_439);
nor U421 (N_421,N_337,N_390);
or U422 (N_422,In_247,N_372);
nor U423 (N_423,N_388,N_368);
nor U424 (N_424,N_419,N_389);
nor U425 (N_425,N_377,N_397);
nand U426 (N_426,N_363,N_376);
or U427 (N_427,N_233,N_374);
nand U428 (N_428,N_416,N_305);
xor U429 (N_429,N_97,N_379);
and U430 (N_430,N_408,N_357);
or U431 (N_431,N_386,N_221);
xnor U432 (N_432,N_260,N_380);
nor U433 (N_433,N_418,N_410);
and U434 (N_434,N_399,N_378);
and U435 (N_435,N_417,N_409);
nor U436 (N_436,N_413,N_370);
nor U437 (N_437,N_366,N_306);
and U438 (N_438,N_365,N_398);
nand U439 (N_439,N_364,N_406);
nand U440 (N_440,N_395,N_285);
or U441 (N_441,N_400,N_396);
and U442 (N_442,N_137,N_153);
nand U443 (N_443,In_411,N_360);
xor U444 (N_444,N_402,N_414);
or U445 (N_445,N_393,N_387);
xor U446 (N_446,N_367,N_373);
xor U447 (N_447,N_381,N_288);
nor U448 (N_448,N_361,N_312);
nand U449 (N_449,N_362,N_401);
or U450 (N_450,N_385,N_371);
or U451 (N_451,N_375,N_190);
nor U452 (N_452,N_415,N_350);
and U453 (N_453,N_329,N_383);
nand U454 (N_454,N_382,N_404);
and U455 (N_455,N_318,N_394);
or U456 (N_456,N_403,N_407);
nor U457 (N_457,N_405,N_369);
and U458 (N_458,N_391,N_411);
nor U459 (N_459,N_384,N_392);
nand U460 (N_460,N_416,N_401);
xnor U461 (N_461,N_403,N_413);
or U462 (N_462,N_398,N_360);
or U463 (N_463,N_399,N_398);
or U464 (N_464,In_247,In_439);
nand U465 (N_465,N_392,N_395);
and U466 (N_466,N_403,N_370);
or U467 (N_467,N_400,N_371);
nand U468 (N_468,N_406,N_392);
or U469 (N_469,N_403,N_398);
or U470 (N_470,N_367,N_382);
or U471 (N_471,N_367,N_414);
and U472 (N_472,N_414,N_418);
nand U473 (N_473,N_404,N_377);
nor U474 (N_474,N_419,N_153);
and U475 (N_475,N_370,N_329);
xor U476 (N_476,N_285,N_409);
nor U477 (N_477,N_221,N_372);
nor U478 (N_478,N_404,N_360);
nand U479 (N_479,N_396,N_370);
and U480 (N_480,N_426,N_456);
or U481 (N_481,N_473,N_421);
xnor U482 (N_482,N_442,N_444);
or U483 (N_483,N_474,N_460);
nand U484 (N_484,N_423,N_479);
xor U485 (N_485,N_432,N_469);
or U486 (N_486,N_441,N_472);
or U487 (N_487,N_468,N_464);
xor U488 (N_488,N_446,N_430);
or U489 (N_489,N_463,N_436);
nor U490 (N_490,N_427,N_452);
nand U491 (N_491,N_420,N_453);
or U492 (N_492,N_445,N_458);
nand U493 (N_493,N_454,N_429);
nor U494 (N_494,N_466,N_455);
or U495 (N_495,N_449,N_461);
and U496 (N_496,N_451,N_443);
and U497 (N_497,N_422,N_450);
xor U498 (N_498,N_471,N_448);
nor U499 (N_499,N_465,N_434);
and U500 (N_500,N_467,N_438);
and U501 (N_501,N_437,N_435);
or U502 (N_502,N_476,N_440);
and U503 (N_503,N_470,N_457);
nor U504 (N_504,N_439,N_425);
xor U505 (N_505,N_431,N_475);
or U506 (N_506,N_428,N_477);
and U507 (N_507,N_424,N_459);
and U508 (N_508,N_447,N_462);
nor U509 (N_509,N_478,N_433);
and U510 (N_510,N_461,N_450);
and U511 (N_511,N_467,N_431);
xor U512 (N_512,N_427,N_475);
nor U513 (N_513,N_458,N_437);
xor U514 (N_514,N_457,N_453);
nand U515 (N_515,N_472,N_427);
nor U516 (N_516,N_461,N_469);
xor U517 (N_517,N_421,N_461);
xnor U518 (N_518,N_459,N_431);
nand U519 (N_519,N_443,N_449);
xnor U520 (N_520,N_456,N_433);
nor U521 (N_521,N_438,N_479);
and U522 (N_522,N_424,N_453);
xnor U523 (N_523,N_444,N_475);
nor U524 (N_524,N_473,N_422);
and U525 (N_525,N_446,N_462);
xor U526 (N_526,N_470,N_449);
or U527 (N_527,N_460,N_478);
nand U528 (N_528,N_462,N_454);
nor U529 (N_529,N_434,N_443);
and U530 (N_530,N_436,N_422);
nor U531 (N_531,N_479,N_458);
xnor U532 (N_532,N_444,N_462);
nand U533 (N_533,N_462,N_452);
nand U534 (N_534,N_476,N_459);
nand U535 (N_535,N_428,N_446);
xor U536 (N_536,N_456,N_431);
or U537 (N_537,N_442,N_457);
or U538 (N_538,N_456,N_423);
or U539 (N_539,N_460,N_467);
nor U540 (N_540,N_539,N_534);
xor U541 (N_541,N_492,N_530);
nor U542 (N_542,N_486,N_521);
nor U543 (N_543,N_499,N_490);
xor U544 (N_544,N_525,N_489);
nand U545 (N_545,N_535,N_498);
and U546 (N_546,N_481,N_512);
xnor U547 (N_547,N_538,N_518);
or U548 (N_548,N_522,N_533);
nor U549 (N_549,N_524,N_495);
or U550 (N_550,N_480,N_487);
nor U551 (N_551,N_496,N_511);
nand U552 (N_552,N_491,N_527);
and U553 (N_553,N_509,N_497);
nor U554 (N_554,N_483,N_493);
nand U555 (N_555,N_516,N_504);
nand U556 (N_556,N_506,N_514);
and U557 (N_557,N_517,N_520);
nand U558 (N_558,N_503,N_502);
or U559 (N_559,N_513,N_482);
and U560 (N_560,N_519,N_485);
nand U561 (N_561,N_529,N_523);
nand U562 (N_562,N_531,N_532);
xor U563 (N_563,N_528,N_507);
and U564 (N_564,N_494,N_505);
xor U565 (N_565,N_501,N_510);
nand U566 (N_566,N_515,N_488);
nand U567 (N_567,N_526,N_500);
nand U568 (N_568,N_536,N_484);
nor U569 (N_569,N_508,N_537);
nor U570 (N_570,N_535,N_508);
and U571 (N_571,N_522,N_510);
or U572 (N_572,N_518,N_484);
or U573 (N_573,N_505,N_516);
xnor U574 (N_574,N_514,N_505);
xnor U575 (N_575,N_506,N_538);
nand U576 (N_576,N_507,N_523);
or U577 (N_577,N_499,N_525);
xor U578 (N_578,N_536,N_526);
or U579 (N_579,N_516,N_495);
and U580 (N_580,N_536,N_525);
or U581 (N_581,N_521,N_483);
and U582 (N_582,N_487,N_499);
and U583 (N_583,N_518,N_501);
nor U584 (N_584,N_503,N_480);
nand U585 (N_585,N_522,N_496);
xor U586 (N_586,N_484,N_523);
and U587 (N_587,N_498,N_518);
and U588 (N_588,N_484,N_493);
or U589 (N_589,N_517,N_506);
or U590 (N_590,N_488,N_505);
nand U591 (N_591,N_527,N_481);
nand U592 (N_592,N_486,N_507);
xor U593 (N_593,N_536,N_480);
nand U594 (N_594,N_526,N_498);
nand U595 (N_595,N_512,N_495);
and U596 (N_596,N_488,N_507);
xnor U597 (N_597,N_495,N_538);
xor U598 (N_598,N_519,N_514);
xnor U599 (N_599,N_513,N_484);
nand U600 (N_600,N_585,N_553);
xnor U601 (N_601,N_575,N_540);
nand U602 (N_602,N_571,N_596);
nand U603 (N_603,N_555,N_590);
and U604 (N_604,N_582,N_541);
xor U605 (N_605,N_552,N_549);
nor U606 (N_606,N_588,N_576);
nand U607 (N_607,N_584,N_594);
nand U608 (N_608,N_595,N_544);
xor U609 (N_609,N_557,N_593);
xnor U610 (N_610,N_572,N_599);
xnor U611 (N_611,N_550,N_586);
or U612 (N_612,N_577,N_580);
xnor U613 (N_613,N_597,N_568);
nand U614 (N_614,N_569,N_574);
and U615 (N_615,N_542,N_543);
nand U616 (N_616,N_589,N_578);
nor U617 (N_617,N_562,N_551);
and U618 (N_618,N_579,N_566);
nor U619 (N_619,N_556,N_547);
and U620 (N_620,N_583,N_573);
nor U621 (N_621,N_558,N_548);
xnor U622 (N_622,N_570,N_567);
xnor U623 (N_623,N_561,N_598);
nor U624 (N_624,N_565,N_581);
and U625 (N_625,N_564,N_560);
and U626 (N_626,N_559,N_545);
or U627 (N_627,N_554,N_587);
nor U628 (N_628,N_591,N_592);
xor U629 (N_629,N_563,N_546);
and U630 (N_630,N_594,N_554);
and U631 (N_631,N_582,N_585);
xor U632 (N_632,N_593,N_556);
nand U633 (N_633,N_596,N_548);
xnor U634 (N_634,N_579,N_573);
nand U635 (N_635,N_571,N_546);
nor U636 (N_636,N_545,N_543);
or U637 (N_637,N_563,N_583);
xnor U638 (N_638,N_595,N_566);
and U639 (N_639,N_547,N_596);
nand U640 (N_640,N_552,N_550);
nand U641 (N_641,N_597,N_564);
nor U642 (N_642,N_581,N_578);
nor U643 (N_643,N_565,N_548);
xor U644 (N_644,N_569,N_555);
nor U645 (N_645,N_561,N_579);
or U646 (N_646,N_555,N_546);
nor U647 (N_647,N_562,N_567);
nand U648 (N_648,N_586,N_568);
and U649 (N_649,N_563,N_566);
and U650 (N_650,N_541,N_588);
and U651 (N_651,N_547,N_580);
xor U652 (N_652,N_594,N_542);
xor U653 (N_653,N_549,N_541);
or U654 (N_654,N_598,N_541);
or U655 (N_655,N_592,N_570);
xnor U656 (N_656,N_595,N_543);
and U657 (N_657,N_584,N_549);
and U658 (N_658,N_549,N_546);
nor U659 (N_659,N_573,N_560);
and U660 (N_660,N_635,N_644);
nand U661 (N_661,N_623,N_657);
or U662 (N_662,N_600,N_614);
or U663 (N_663,N_609,N_622);
nor U664 (N_664,N_649,N_602);
or U665 (N_665,N_627,N_629);
xnor U666 (N_666,N_640,N_648);
nor U667 (N_667,N_633,N_630);
nor U668 (N_668,N_645,N_643);
xnor U669 (N_669,N_608,N_652);
xnor U670 (N_670,N_658,N_615);
nand U671 (N_671,N_620,N_628);
xnor U672 (N_672,N_634,N_626);
and U673 (N_673,N_632,N_616);
xor U674 (N_674,N_604,N_641);
xor U675 (N_675,N_636,N_607);
nand U676 (N_676,N_613,N_646);
and U677 (N_677,N_655,N_612);
xor U678 (N_678,N_617,N_601);
xor U679 (N_679,N_606,N_651);
and U680 (N_680,N_653,N_639);
and U681 (N_681,N_619,N_603);
or U682 (N_682,N_638,N_631);
and U683 (N_683,N_642,N_624);
nor U684 (N_684,N_611,N_656);
and U685 (N_685,N_654,N_659);
and U686 (N_686,N_650,N_610);
nand U687 (N_687,N_605,N_625);
xnor U688 (N_688,N_647,N_618);
and U689 (N_689,N_621,N_637);
nand U690 (N_690,N_620,N_609);
nand U691 (N_691,N_622,N_603);
or U692 (N_692,N_636,N_604);
or U693 (N_693,N_644,N_611);
nor U694 (N_694,N_653,N_655);
nor U695 (N_695,N_613,N_649);
xor U696 (N_696,N_623,N_641);
xnor U697 (N_697,N_634,N_650);
xnor U698 (N_698,N_653,N_620);
and U699 (N_699,N_657,N_601);
xnor U700 (N_700,N_640,N_633);
and U701 (N_701,N_656,N_636);
nand U702 (N_702,N_610,N_632);
and U703 (N_703,N_645,N_634);
nand U704 (N_704,N_643,N_618);
and U705 (N_705,N_612,N_627);
and U706 (N_706,N_632,N_640);
nor U707 (N_707,N_632,N_618);
xor U708 (N_708,N_659,N_623);
nand U709 (N_709,N_620,N_639);
nand U710 (N_710,N_659,N_629);
and U711 (N_711,N_633,N_613);
nor U712 (N_712,N_632,N_629);
nor U713 (N_713,N_624,N_630);
nor U714 (N_714,N_644,N_655);
nor U715 (N_715,N_608,N_618);
or U716 (N_716,N_631,N_642);
or U717 (N_717,N_637,N_602);
or U718 (N_718,N_648,N_654);
xor U719 (N_719,N_618,N_620);
nor U720 (N_720,N_678,N_717);
nor U721 (N_721,N_692,N_714);
nor U722 (N_722,N_672,N_666);
or U723 (N_723,N_673,N_680);
xor U724 (N_724,N_682,N_670);
or U725 (N_725,N_689,N_686);
nand U726 (N_726,N_684,N_709);
nand U727 (N_727,N_702,N_687);
or U728 (N_728,N_708,N_715);
xnor U729 (N_729,N_701,N_704);
xnor U730 (N_730,N_664,N_668);
nand U731 (N_731,N_677,N_713);
nor U732 (N_732,N_710,N_681);
nand U733 (N_733,N_688,N_706);
xnor U734 (N_734,N_695,N_691);
and U735 (N_735,N_667,N_662);
nor U736 (N_736,N_698,N_716);
and U737 (N_737,N_712,N_700);
xor U738 (N_738,N_693,N_696);
xnor U739 (N_739,N_663,N_707);
or U740 (N_740,N_675,N_705);
or U741 (N_741,N_679,N_697);
xnor U742 (N_742,N_676,N_690);
xnor U743 (N_743,N_685,N_703);
xnor U744 (N_744,N_694,N_671);
xor U745 (N_745,N_719,N_718);
nor U746 (N_746,N_699,N_665);
nor U747 (N_747,N_660,N_711);
and U748 (N_748,N_683,N_661);
or U749 (N_749,N_669,N_674);
or U750 (N_750,N_660,N_707);
nand U751 (N_751,N_715,N_678);
nand U752 (N_752,N_696,N_701);
or U753 (N_753,N_711,N_670);
and U754 (N_754,N_697,N_694);
xnor U755 (N_755,N_665,N_684);
xor U756 (N_756,N_683,N_691);
nor U757 (N_757,N_702,N_682);
xnor U758 (N_758,N_711,N_705);
nor U759 (N_759,N_709,N_682);
or U760 (N_760,N_701,N_666);
xnor U761 (N_761,N_699,N_702);
xor U762 (N_762,N_702,N_661);
nor U763 (N_763,N_687,N_697);
and U764 (N_764,N_704,N_677);
xor U765 (N_765,N_704,N_698);
xor U766 (N_766,N_698,N_694);
nor U767 (N_767,N_696,N_713);
nor U768 (N_768,N_707,N_679);
nand U769 (N_769,N_704,N_676);
nor U770 (N_770,N_668,N_687);
or U771 (N_771,N_713,N_673);
xnor U772 (N_772,N_677,N_698);
and U773 (N_773,N_660,N_697);
and U774 (N_774,N_707,N_718);
nand U775 (N_775,N_661,N_717);
or U776 (N_776,N_664,N_682);
nand U777 (N_777,N_714,N_702);
nor U778 (N_778,N_685,N_667);
nor U779 (N_779,N_680,N_666);
nand U780 (N_780,N_775,N_757);
and U781 (N_781,N_746,N_747);
nand U782 (N_782,N_769,N_759);
or U783 (N_783,N_739,N_764);
xnor U784 (N_784,N_749,N_738);
xor U785 (N_785,N_734,N_770);
nand U786 (N_786,N_736,N_778);
or U787 (N_787,N_729,N_768);
nor U788 (N_788,N_732,N_766);
nor U789 (N_789,N_762,N_771);
xnor U790 (N_790,N_735,N_743);
and U791 (N_791,N_779,N_725);
xor U792 (N_792,N_767,N_772);
xor U793 (N_793,N_730,N_773);
nor U794 (N_794,N_723,N_774);
or U795 (N_795,N_765,N_742);
nor U796 (N_796,N_741,N_720);
xnor U797 (N_797,N_753,N_728);
nor U798 (N_798,N_750,N_755);
or U799 (N_799,N_752,N_744);
xnor U800 (N_800,N_724,N_733);
or U801 (N_801,N_761,N_754);
nand U802 (N_802,N_722,N_731);
or U803 (N_803,N_763,N_727);
nor U804 (N_804,N_777,N_776);
or U805 (N_805,N_748,N_737);
nand U806 (N_806,N_751,N_756);
nor U807 (N_807,N_726,N_758);
nand U808 (N_808,N_721,N_740);
nand U809 (N_809,N_745,N_760);
or U810 (N_810,N_771,N_761);
and U811 (N_811,N_753,N_773);
and U812 (N_812,N_740,N_759);
or U813 (N_813,N_737,N_778);
xnor U814 (N_814,N_773,N_737);
xor U815 (N_815,N_777,N_742);
nand U816 (N_816,N_740,N_728);
nand U817 (N_817,N_751,N_776);
nor U818 (N_818,N_766,N_731);
or U819 (N_819,N_755,N_749);
nand U820 (N_820,N_721,N_726);
and U821 (N_821,N_736,N_769);
and U822 (N_822,N_752,N_727);
nand U823 (N_823,N_748,N_738);
nor U824 (N_824,N_732,N_750);
nor U825 (N_825,N_723,N_777);
xor U826 (N_826,N_736,N_771);
and U827 (N_827,N_744,N_776);
or U828 (N_828,N_727,N_721);
nor U829 (N_829,N_721,N_746);
nor U830 (N_830,N_773,N_767);
nor U831 (N_831,N_770,N_733);
xor U832 (N_832,N_752,N_730);
nor U833 (N_833,N_757,N_770);
nand U834 (N_834,N_759,N_732);
and U835 (N_835,N_768,N_763);
nand U836 (N_836,N_722,N_723);
and U837 (N_837,N_757,N_760);
or U838 (N_838,N_766,N_771);
nand U839 (N_839,N_744,N_758);
nand U840 (N_840,N_836,N_829);
and U841 (N_841,N_790,N_803);
nand U842 (N_842,N_801,N_789);
and U843 (N_843,N_818,N_835);
nand U844 (N_844,N_802,N_806);
xor U845 (N_845,N_797,N_798);
or U846 (N_846,N_816,N_809);
nand U847 (N_847,N_833,N_783);
and U848 (N_848,N_837,N_832);
nand U849 (N_849,N_787,N_782);
and U850 (N_850,N_817,N_824);
xnor U851 (N_851,N_827,N_805);
xnor U852 (N_852,N_784,N_800);
and U853 (N_853,N_799,N_826);
or U854 (N_854,N_804,N_788);
or U855 (N_855,N_795,N_830);
or U856 (N_856,N_791,N_786);
and U857 (N_857,N_780,N_834);
or U858 (N_858,N_825,N_793);
and U859 (N_859,N_810,N_794);
and U860 (N_860,N_821,N_828);
nor U861 (N_861,N_785,N_808);
and U862 (N_862,N_820,N_781);
and U863 (N_863,N_814,N_819);
nand U864 (N_864,N_807,N_812);
nand U865 (N_865,N_823,N_831);
or U866 (N_866,N_822,N_811);
or U867 (N_867,N_838,N_815);
nor U868 (N_868,N_792,N_839);
or U869 (N_869,N_796,N_813);
nand U870 (N_870,N_808,N_839);
nand U871 (N_871,N_834,N_795);
and U872 (N_872,N_826,N_832);
xnor U873 (N_873,N_804,N_827);
nand U874 (N_874,N_830,N_825);
nor U875 (N_875,N_802,N_784);
nor U876 (N_876,N_839,N_807);
nor U877 (N_877,N_829,N_822);
xnor U878 (N_878,N_788,N_838);
nor U879 (N_879,N_814,N_805);
nand U880 (N_880,N_782,N_786);
or U881 (N_881,N_819,N_800);
and U882 (N_882,N_803,N_793);
and U883 (N_883,N_797,N_831);
or U884 (N_884,N_835,N_788);
xor U885 (N_885,N_797,N_830);
nor U886 (N_886,N_833,N_839);
xor U887 (N_887,N_819,N_784);
and U888 (N_888,N_784,N_807);
or U889 (N_889,N_782,N_814);
or U890 (N_890,N_791,N_785);
nor U891 (N_891,N_838,N_833);
nor U892 (N_892,N_791,N_793);
nor U893 (N_893,N_800,N_808);
xnor U894 (N_894,N_799,N_836);
nand U895 (N_895,N_822,N_792);
and U896 (N_896,N_821,N_829);
or U897 (N_897,N_781,N_793);
nand U898 (N_898,N_789,N_827);
and U899 (N_899,N_786,N_796);
and U900 (N_900,N_873,N_899);
or U901 (N_901,N_864,N_853);
nor U902 (N_902,N_892,N_857);
nor U903 (N_903,N_867,N_894);
or U904 (N_904,N_887,N_874);
or U905 (N_905,N_888,N_889);
xnor U906 (N_906,N_844,N_842);
and U907 (N_907,N_869,N_872);
and U908 (N_908,N_897,N_885);
nand U909 (N_909,N_886,N_840);
or U910 (N_910,N_882,N_841);
or U911 (N_911,N_855,N_876);
or U912 (N_912,N_893,N_863);
nand U913 (N_913,N_880,N_856);
nand U914 (N_914,N_895,N_851);
and U915 (N_915,N_878,N_879);
xor U916 (N_916,N_861,N_898);
nor U917 (N_917,N_846,N_884);
and U918 (N_918,N_848,N_849);
xor U919 (N_919,N_860,N_865);
xor U920 (N_920,N_866,N_852);
and U921 (N_921,N_896,N_891);
nor U922 (N_922,N_877,N_845);
nand U923 (N_923,N_847,N_843);
or U924 (N_924,N_890,N_871);
or U925 (N_925,N_868,N_870);
nand U926 (N_926,N_875,N_881);
nor U927 (N_927,N_859,N_858);
nor U928 (N_928,N_862,N_854);
nand U929 (N_929,N_883,N_850);
and U930 (N_930,N_843,N_864);
nand U931 (N_931,N_871,N_847);
or U932 (N_932,N_880,N_899);
nand U933 (N_933,N_887,N_881);
or U934 (N_934,N_894,N_864);
nor U935 (N_935,N_841,N_871);
nand U936 (N_936,N_888,N_850);
nor U937 (N_937,N_867,N_861);
and U938 (N_938,N_851,N_841);
xor U939 (N_939,N_850,N_860);
or U940 (N_940,N_859,N_877);
nor U941 (N_941,N_883,N_881);
nand U942 (N_942,N_845,N_879);
and U943 (N_943,N_870,N_857);
nor U944 (N_944,N_844,N_845);
and U945 (N_945,N_845,N_864);
xnor U946 (N_946,N_841,N_885);
or U947 (N_947,N_847,N_865);
or U948 (N_948,N_854,N_877);
and U949 (N_949,N_847,N_898);
nand U950 (N_950,N_871,N_877);
nand U951 (N_951,N_867,N_881);
xor U952 (N_952,N_850,N_879);
nand U953 (N_953,N_884,N_860);
xor U954 (N_954,N_878,N_865);
nor U955 (N_955,N_890,N_861);
xnor U956 (N_956,N_858,N_851);
or U957 (N_957,N_843,N_871);
and U958 (N_958,N_879,N_875);
nor U959 (N_959,N_889,N_881);
or U960 (N_960,N_911,N_901);
or U961 (N_961,N_933,N_917);
or U962 (N_962,N_953,N_942);
or U963 (N_963,N_920,N_921);
or U964 (N_964,N_919,N_958);
nand U965 (N_965,N_907,N_915);
and U966 (N_966,N_948,N_955);
and U967 (N_967,N_954,N_934);
nor U968 (N_968,N_956,N_913);
xnor U969 (N_969,N_938,N_940);
and U970 (N_970,N_957,N_922);
xnor U971 (N_971,N_904,N_950);
and U972 (N_972,N_902,N_935);
or U973 (N_973,N_943,N_951);
nand U974 (N_974,N_928,N_944);
and U975 (N_975,N_949,N_929);
nand U976 (N_976,N_910,N_947);
or U977 (N_977,N_916,N_906);
xor U978 (N_978,N_905,N_931);
xor U979 (N_979,N_926,N_912);
and U980 (N_980,N_903,N_936);
nor U981 (N_981,N_945,N_932);
nand U982 (N_982,N_941,N_939);
or U983 (N_983,N_909,N_946);
nand U984 (N_984,N_914,N_930);
xor U985 (N_985,N_923,N_900);
xnor U986 (N_986,N_927,N_908);
nand U987 (N_987,N_924,N_937);
and U988 (N_988,N_918,N_952);
and U989 (N_989,N_959,N_925);
nor U990 (N_990,N_924,N_908);
or U991 (N_991,N_910,N_932);
nor U992 (N_992,N_913,N_945);
and U993 (N_993,N_902,N_936);
nand U994 (N_994,N_958,N_925);
and U995 (N_995,N_920,N_905);
and U996 (N_996,N_906,N_905);
nand U997 (N_997,N_906,N_946);
and U998 (N_998,N_944,N_937);
nand U999 (N_999,N_957,N_916);
or U1000 (N_1000,N_954,N_902);
nand U1001 (N_1001,N_901,N_944);
xor U1002 (N_1002,N_902,N_956);
nand U1003 (N_1003,N_901,N_926);
or U1004 (N_1004,N_949,N_926);
or U1005 (N_1005,N_911,N_929);
xor U1006 (N_1006,N_912,N_906);
and U1007 (N_1007,N_913,N_914);
xnor U1008 (N_1008,N_941,N_959);
xor U1009 (N_1009,N_958,N_946);
and U1010 (N_1010,N_956,N_907);
nor U1011 (N_1011,N_932,N_913);
and U1012 (N_1012,N_935,N_917);
nand U1013 (N_1013,N_931,N_942);
and U1014 (N_1014,N_911,N_918);
xor U1015 (N_1015,N_925,N_946);
nor U1016 (N_1016,N_958,N_935);
nor U1017 (N_1017,N_944,N_902);
or U1018 (N_1018,N_945,N_901);
nor U1019 (N_1019,N_937,N_926);
or U1020 (N_1020,N_978,N_998);
and U1021 (N_1021,N_1011,N_974);
nor U1022 (N_1022,N_1016,N_963);
nand U1023 (N_1023,N_1017,N_973);
xnor U1024 (N_1024,N_990,N_1015);
or U1025 (N_1025,N_1007,N_1010);
xnor U1026 (N_1026,N_996,N_1019);
nor U1027 (N_1027,N_988,N_1000);
xnor U1028 (N_1028,N_972,N_991);
nor U1029 (N_1029,N_962,N_1012);
and U1030 (N_1030,N_981,N_997);
xor U1031 (N_1031,N_1014,N_977);
nor U1032 (N_1032,N_982,N_985);
and U1033 (N_1033,N_984,N_969);
xor U1034 (N_1034,N_989,N_1001);
nor U1035 (N_1035,N_964,N_961);
and U1036 (N_1036,N_1009,N_1003);
xor U1037 (N_1037,N_983,N_993);
nor U1038 (N_1038,N_1018,N_965);
nand U1039 (N_1039,N_987,N_966);
nand U1040 (N_1040,N_1005,N_992);
xor U1041 (N_1041,N_986,N_970);
or U1042 (N_1042,N_967,N_968);
xnor U1043 (N_1043,N_971,N_1008);
nand U1044 (N_1044,N_999,N_960);
and U1045 (N_1045,N_994,N_1006);
and U1046 (N_1046,N_1013,N_995);
xnor U1047 (N_1047,N_979,N_1002);
nor U1048 (N_1048,N_976,N_980);
and U1049 (N_1049,N_975,N_1004);
nand U1050 (N_1050,N_986,N_965);
nand U1051 (N_1051,N_962,N_989);
or U1052 (N_1052,N_992,N_983);
xnor U1053 (N_1053,N_995,N_1001);
and U1054 (N_1054,N_985,N_1010);
nor U1055 (N_1055,N_997,N_1005);
and U1056 (N_1056,N_1012,N_972);
nor U1057 (N_1057,N_997,N_963);
xor U1058 (N_1058,N_1003,N_986);
nor U1059 (N_1059,N_992,N_962);
and U1060 (N_1060,N_1010,N_966);
or U1061 (N_1061,N_989,N_1010);
and U1062 (N_1062,N_978,N_963);
xor U1063 (N_1063,N_961,N_1013);
and U1064 (N_1064,N_1009,N_963);
nor U1065 (N_1065,N_972,N_976);
nor U1066 (N_1066,N_996,N_979);
xnor U1067 (N_1067,N_988,N_987);
or U1068 (N_1068,N_1012,N_976);
or U1069 (N_1069,N_978,N_962);
and U1070 (N_1070,N_975,N_1006);
xor U1071 (N_1071,N_991,N_1006);
xnor U1072 (N_1072,N_972,N_1011);
nor U1073 (N_1073,N_1015,N_979);
xnor U1074 (N_1074,N_976,N_973);
nand U1075 (N_1075,N_994,N_996);
nor U1076 (N_1076,N_961,N_966);
or U1077 (N_1077,N_1019,N_988);
nand U1078 (N_1078,N_982,N_1009);
nor U1079 (N_1079,N_982,N_1006);
and U1080 (N_1080,N_1043,N_1070);
or U1081 (N_1081,N_1029,N_1040);
and U1082 (N_1082,N_1027,N_1075);
xnor U1083 (N_1083,N_1025,N_1061);
or U1084 (N_1084,N_1076,N_1063);
nand U1085 (N_1085,N_1057,N_1032);
xnor U1086 (N_1086,N_1078,N_1021);
nand U1087 (N_1087,N_1037,N_1044);
xnor U1088 (N_1088,N_1052,N_1041);
nand U1089 (N_1089,N_1047,N_1066);
nor U1090 (N_1090,N_1064,N_1071);
nand U1091 (N_1091,N_1050,N_1049);
xnor U1092 (N_1092,N_1033,N_1077);
nor U1093 (N_1093,N_1058,N_1056);
or U1094 (N_1094,N_1055,N_1038);
nor U1095 (N_1095,N_1020,N_1079);
xnor U1096 (N_1096,N_1039,N_1074);
nor U1097 (N_1097,N_1023,N_1062);
nand U1098 (N_1098,N_1031,N_1067);
xor U1099 (N_1099,N_1073,N_1069);
and U1100 (N_1100,N_1059,N_1022);
or U1101 (N_1101,N_1060,N_1048);
and U1102 (N_1102,N_1036,N_1046);
xor U1103 (N_1103,N_1072,N_1030);
nor U1104 (N_1104,N_1034,N_1028);
nand U1105 (N_1105,N_1042,N_1053);
and U1106 (N_1106,N_1035,N_1026);
and U1107 (N_1107,N_1051,N_1024);
xnor U1108 (N_1108,N_1054,N_1065);
nand U1109 (N_1109,N_1045,N_1068);
xor U1110 (N_1110,N_1048,N_1023);
or U1111 (N_1111,N_1025,N_1022);
xor U1112 (N_1112,N_1049,N_1063);
or U1113 (N_1113,N_1046,N_1024);
xnor U1114 (N_1114,N_1027,N_1024);
or U1115 (N_1115,N_1062,N_1057);
xor U1116 (N_1116,N_1067,N_1059);
xor U1117 (N_1117,N_1070,N_1048);
nand U1118 (N_1118,N_1034,N_1062);
or U1119 (N_1119,N_1066,N_1027);
or U1120 (N_1120,N_1036,N_1071);
nor U1121 (N_1121,N_1072,N_1065);
nor U1122 (N_1122,N_1021,N_1037);
and U1123 (N_1123,N_1027,N_1023);
or U1124 (N_1124,N_1069,N_1022);
or U1125 (N_1125,N_1075,N_1020);
and U1126 (N_1126,N_1028,N_1067);
xnor U1127 (N_1127,N_1022,N_1060);
nand U1128 (N_1128,N_1047,N_1071);
nor U1129 (N_1129,N_1047,N_1028);
nor U1130 (N_1130,N_1070,N_1063);
nor U1131 (N_1131,N_1059,N_1045);
or U1132 (N_1132,N_1051,N_1044);
or U1133 (N_1133,N_1023,N_1064);
nand U1134 (N_1134,N_1071,N_1072);
nor U1135 (N_1135,N_1046,N_1049);
and U1136 (N_1136,N_1073,N_1054);
xnor U1137 (N_1137,N_1055,N_1044);
or U1138 (N_1138,N_1032,N_1025);
or U1139 (N_1139,N_1030,N_1069);
nor U1140 (N_1140,N_1137,N_1107);
xor U1141 (N_1141,N_1103,N_1084);
nand U1142 (N_1142,N_1108,N_1129);
nand U1143 (N_1143,N_1097,N_1110);
and U1144 (N_1144,N_1138,N_1113);
nand U1145 (N_1145,N_1096,N_1080);
xnor U1146 (N_1146,N_1082,N_1101);
nand U1147 (N_1147,N_1139,N_1106);
or U1148 (N_1148,N_1135,N_1099);
nor U1149 (N_1149,N_1118,N_1127);
and U1150 (N_1150,N_1093,N_1121);
nand U1151 (N_1151,N_1119,N_1098);
xnor U1152 (N_1152,N_1115,N_1105);
nand U1153 (N_1153,N_1125,N_1109);
xnor U1154 (N_1154,N_1120,N_1132);
and U1155 (N_1155,N_1089,N_1133);
or U1156 (N_1156,N_1117,N_1136);
nor U1157 (N_1157,N_1114,N_1083);
xor U1158 (N_1158,N_1086,N_1090);
xnor U1159 (N_1159,N_1104,N_1124);
nor U1160 (N_1160,N_1123,N_1094);
or U1161 (N_1161,N_1085,N_1131);
xor U1162 (N_1162,N_1088,N_1126);
xnor U1163 (N_1163,N_1122,N_1112);
and U1164 (N_1164,N_1134,N_1081);
xor U1165 (N_1165,N_1100,N_1128);
xor U1166 (N_1166,N_1102,N_1091);
or U1167 (N_1167,N_1087,N_1116);
or U1168 (N_1168,N_1095,N_1092);
nand U1169 (N_1169,N_1111,N_1130);
xor U1170 (N_1170,N_1109,N_1106);
nor U1171 (N_1171,N_1129,N_1103);
nand U1172 (N_1172,N_1089,N_1114);
xor U1173 (N_1173,N_1126,N_1112);
and U1174 (N_1174,N_1114,N_1085);
nand U1175 (N_1175,N_1092,N_1083);
or U1176 (N_1176,N_1093,N_1116);
xor U1177 (N_1177,N_1118,N_1114);
and U1178 (N_1178,N_1137,N_1120);
nand U1179 (N_1179,N_1125,N_1089);
nor U1180 (N_1180,N_1132,N_1114);
or U1181 (N_1181,N_1112,N_1119);
and U1182 (N_1182,N_1112,N_1138);
xnor U1183 (N_1183,N_1119,N_1093);
xor U1184 (N_1184,N_1093,N_1107);
xor U1185 (N_1185,N_1108,N_1139);
and U1186 (N_1186,N_1123,N_1115);
or U1187 (N_1187,N_1116,N_1091);
nor U1188 (N_1188,N_1103,N_1137);
and U1189 (N_1189,N_1081,N_1123);
xor U1190 (N_1190,N_1118,N_1134);
xnor U1191 (N_1191,N_1117,N_1107);
and U1192 (N_1192,N_1116,N_1104);
nor U1193 (N_1193,N_1123,N_1135);
nor U1194 (N_1194,N_1119,N_1114);
nand U1195 (N_1195,N_1136,N_1092);
xnor U1196 (N_1196,N_1137,N_1104);
and U1197 (N_1197,N_1095,N_1113);
or U1198 (N_1198,N_1129,N_1135);
or U1199 (N_1199,N_1113,N_1102);
xnor U1200 (N_1200,N_1145,N_1146);
nand U1201 (N_1201,N_1175,N_1191);
or U1202 (N_1202,N_1186,N_1174);
xor U1203 (N_1203,N_1173,N_1177);
and U1204 (N_1204,N_1157,N_1192);
and U1205 (N_1205,N_1168,N_1189);
nor U1206 (N_1206,N_1140,N_1150);
and U1207 (N_1207,N_1181,N_1156);
nand U1208 (N_1208,N_1178,N_1199);
xnor U1209 (N_1209,N_1152,N_1143);
xor U1210 (N_1210,N_1180,N_1193);
nand U1211 (N_1211,N_1166,N_1176);
or U1212 (N_1212,N_1182,N_1159);
and U1213 (N_1213,N_1190,N_1164);
nand U1214 (N_1214,N_1170,N_1169);
and U1215 (N_1215,N_1167,N_1165);
xor U1216 (N_1216,N_1198,N_1160);
xnor U1217 (N_1217,N_1187,N_1147);
and U1218 (N_1218,N_1142,N_1141);
nand U1219 (N_1219,N_1154,N_1179);
xnor U1220 (N_1220,N_1148,N_1184);
and U1221 (N_1221,N_1197,N_1196);
and U1222 (N_1222,N_1172,N_1151);
or U1223 (N_1223,N_1162,N_1144);
nor U1224 (N_1224,N_1185,N_1161);
nor U1225 (N_1225,N_1149,N_1171);
nand U1226 (N_1226,N_1194,N_1155);
and U1227 (N_1227,N_1183,N_1188);
nor U1228 (N_1228,N_1195,N_1153);
and U1229 (N_1229,N_1163,N_1158);
nor U1230 (N_1230,N_1165,N_1170);
and U1231 (N_1231,N_1149,N_1168);
nor U1232 (N_1232,N_1177,N_1184);
or U1233 (N_1233,N_1157,N_1172);
and U1234 (N_1234,N_1162,N_1147);
and U1235 (N_1235,N_1161,N_1162);
and U1236 (N_1236,N_1164,N_1184);
xor U1237 (N_1237,N_1168,N_1180);
and U1238 (N_1238,N_1188,N_1195);
and U1239 (N_1239,N_1189,N_1195);
and U1240 (N_1240,N_1163,N_1174);
nor U1241 (N_1241,N_1147,N_1180);
xnor U1242 (N_1242,N_1147,N_1149);
or U1243 (N_1243,N_1166,N_1199);
and U1244 (N_1244,N_1146,N_1194);
and U1245 (N_1245,N_1174,N_1155);
nand U1246 (N_1246,N_1182,N_1167);
or U1247 (N_1247,N_1171,N_1142);
and U1248 (N_1248,N_1185,N_1178);
or U1249 (N_1249,N_1143,N_1185);
nand U1250 (N_1250,N_1156,N_1144);
nor U1251 (N_1251,N_1195,N_1167);
xnor U1252 (N_1252,N_1179,N_1192);
xor U1253 (N_1253,N_1159,N_1171);
or U1254 (N_1254,N_1194,N_1163);
or U1255 (N_1255,N_1140,N_1177);
nand U1256 (N_1256,N_1175,N_1199);
or U1257 (N_1257,N_1170,N_1151);
nor U1258 (N_1258,N_1152,N_1163);
xor U1259 (N_1259,N_1198,N_1190);
nor U1260 (N_1260,N_1244,N_1224);
xor U1261 (N_1261,N_1243,N_1251);
nor U1262 (N_1262,N_1213,N_1212);
xor U1263 (N_1263,N_1220,N_1219);
or U1264 (N_1264,N_1245,N_1210);
nor U1265 (N_1265,N_1200,N_1207);
and U1266 (N_1266,N_1221,N_1229);
nor U1267 (N_1267,N_1252,N_1206);
nand U1268 (N_1268,N_1250,N_1246);
and U1269 (N_1269,N_1259,N_1203);
nand U1270 (N_1270,N_1249,N_1255);
nor U1271 (N_1271,N_1253,N_1201);
nand U1272 (N_1272,N_1217,N_1242);
nand U1273 (N_1273,N_1256,N_1247);
and U1274 (N_1274,N_1228,N_1215);
or U1275 (N_1275,N_1225,N_1208);
and U1276 (N_1276,N_1254,N_1248);
and U1277 (N_1277,N_1222,N_1216);
or U1278 (N_1278,N_1226,N_1232);
nor U1279 (N_1279,N_1230,N_1218);
and U1280 (N_1280,N_1233,N_1205);
xor U1281 (N_1281,N_1231,N_1235);
nand U1282 (N_1282,N_1240,N_1214);
nor U1283 (N_1283,N_1202,N_1241);
or U1284 (N_1284,N_1236,N_1238);
xor U1285 (N_1285,N_1227,N_1239);
nor U1286 (N_1286,N_1258,N_1223);
and U1287 (N_1287,N_1257,N_1237);
or U1288 (N_1288,N_1234,N_1211);
xnor U1289 (N_1289,N_1204,N_1209);
nand U1290 (N_1290,N_1251,N_1247);
xnor U1291 (N_1291,N_1246,N_1251);
nand U1292 (N_1292,N_1218,N_1223);
nand U1293 (N_1293,N_1253,N_1207);
nor U1294 (N_1294,N_1238,N_1231);
xnor U1295 (N_1295,N_1227,N_1231);
and U1296 (N_1296,N_1246,N_1243);
and U1297 (N_1297,N_1219,N_1241);
and U1298 (N_1298,N_1239,N_1243);
or U1299 (N_1299,N_1255,N_1245);
or U1300 (N_1300,N_1258,N_1203);
xnor U1301 (N_1301,N_1206,N_1242);
xor U1302 (N_1302,N_1207,N_1249);
nand U1303 (N_1303,N_1241,N_1226);
nand U1304 (N_1304,N_1230,N_1214);
xor U1305 (N_1305,N_1209,N_1201);
or U1306 (N_1306,N_1238,N_1247);
nor U1307 (N_1307,N_1226,N_1238);
nor U1308 (N_1308,N_1255,N_1202);
xor U1309 (N_1309,N_1240,N_1210);
xnor U1310 (N_1310,N_1201,N_1222);
xor U1311 (N_1311,N_1204,N_1215);
and U1312 (N_1312,N_1229,N_1207);
xor U1313 (N_1313,N_1230,N_1223);
or U1314 (N_1314,N_1206,N_1258);
nand U1315 (N_1315,N_1208,N_1207);
and U1316 (N_1316,N_1213,N_1236);
nor U1317 (N_1317,N_1249,N_1218);
nor U1318 (N_1318,N_1215,N_1231);
or U1319 (N_1319,N_1238,N_1252);
nor U1320 (N_1320,N_1279,N_1302);
and U1321 (N_1321,N_1312,N_1274);
nand U1322 (N_1322,N_1261,N_1308);
or U1323 (N_1323,N_1300,N_1307);
xnor U1324 (N_1324,N_1303,N_1284);
xnor U1325 (N_1325,N_1294,N_1275);
nor U1326 (N_1326,N_1299,N_1314);
xnor U1327 (N_1327,N_1282,N_1273);
nor U1328 (N_1328,N_1306,N_1287);
or U1329 (N_1329,N_1301,N_1298);
or U1330 (N_1330,N_1309,N_1263);
nor U1331 (N_1331,N_1283,N_1292);
xnor U1332 (N_1332,N_1277,N_1269);
and U1333 (N_1333,N_1316,N_1315);
or U1334 (N_1334,N_1264,N_1311);
nor U1335 (N_1335,N_1318,N_1317);
and U1336 (N_1336,N_1281,N_1286);
xor U1337 (N_1337,N_1289,N_1260);
nor U1338 (N_1338,N_1304,N_1265);
or U1339 (N_1339,N_1290,N_1291);
nand U1340 (N_1340,N_1272,N_1297);
nor U1341 (N_1341,N_1319,N_1296);
nor U1342 (N_1342,N_1305,N_1313);
and U1343 (N_1343,N_1266,N_1271);
and U1344 (N_1344,N_1293,N_1262);
or U1345 (N_1345,N_1288,N_1295);
xnor U1346 (N_1346,N_1285,N_1278);
nand U1347 (N_1347,N_1268,N_1270);
or U1348 (N_1348,N_1276,N_1280);
xnor U1349 (N_1349,N_1267,N_1310);
or U1350 (N_1350,N_1266,N_1311);
or U1351 (N_1351,N_1296,N_1313);
or U1352 (N_1352,N_1315,N_1262);
nand U1353 (N_1353,N_1262,N_1284);
nor U1354 (N_1354,N_1304,N_1315);
or U1355 (N_1355,N_1296,N_1308);
xor U1356 (N_1356,N_1270,N_1291);
nor U1357 (N_1357,N_1317,N_1291);
or U1358 (N_1358,N_1312,N_1306);
and U1359 (N_1359,N_1290,N_1295);
nand U1360 (N_1360,N_1304,N_1309);
xor U1361 (N_1361,N_1286,N_1291);
and U1362 (N_1362,N_1308,N_1305);
and U1363 (N_1363,N_1318,N_1307);
nor U1364 (N_1364,N_1302,N_1281);
xor U1365 (N_1365,N_1261,N_1306);
or U1366 (N_1366,N_1287,N_1294);
or U1367 (N_1367,N_1317,N_1275);
or U1368 (N_1368,N_1278,N_1261);
nand U1369 (N_1369,N_1269,N_1265);
xnor U1370 (N_1370,N_1307,N_1298);
and U1371 (N_1371,N_1283,N_1265);
or U1372 (N_1372,N_1280,N_1286);
nor U1373 (N_1373,N_1286,N_1263);
xnor U1374 (N_1374,N_1317,N_1303);
nand U1375 (N_1375,N_1266,N_1290);
and U1376 (N_1376,N_1303,N_1292);
or U1377 (N_1377,N_1261,N_1309);
nand U1378 (N_1378,N_1297,N_1301);
nand U1379 (N_1379,N_1303,N_1315);
or U1380 (N_1380,N_1335,N_1359);
nand U1381 (N_1381,N_1344,N_1325);
and U1382 (N_1382,N_1368,N_1349);
and U1383 (N_1383,N_1355,N_1348);
nand U1384 (N_1384,N_1353,N_1338);
nor U1385 (N_1385,N_1378,N_1324);
xnor U1386 (N_1386,N_1361,N_1345);
nand U1387 (N_1387,N_1334,N_1375);
nor U1388 (N_1388,N_1377,N_1364);
and U1389 (N_1389,N_1371,N_1330);
or U1390 (N_1390,N_1358,N_1322);
xor U1391 (N_1391,N_1360,N_1336);
or U1392 (N_1392,N_1333,N_1379);
or U1393 (N_1393,N_1328,N_1340);
nand U1394 (N_1394,N_1332,N_1346);
nor U1395 (N_1395,N_1357,N_1321);
nand U1396 (N_1396,N_1326,N_1331);
nand U1397 (N_1397,N_1362,N_1373);
nand U1398 (N_1398,N_1367,N_1376);
nand U1399 (N_1399,N_1347,N_1341);
nand U1400 (N_1400,N_1343,N_1354);
and U1401 (N_1401,N_1356,N_1342);
nor U1402 (N_1402,N_1370,N_1365);
nand U1403 (N_1403,N_1351,N_1350);
or U1404 (N_1404,N_1372,N_1323);
xor U1405 (N_1405,N_1352,N_1366);
nor U1406 (N_1406,N_1329,N_1363);
and U1407 (N_1407,N_1337,N_1327);
or U1408 (N_1408,N_1339,N_1374);
nand U1409 (N_1409,N_1369,N_1320);
nor U1410 (N_1410,N_1357,N_1347);
nor U1411 (N_1411,N_1336,N_1370);
nand U1412 (N_1412,N_1328,N_1358);
or U1413 (N_1413,N_1341,N_1320);
and U1414 (N_1414,N_1325,N_1337);
nand U1415 (N_1415,N_1344,N_1366);
nor U1416 (N_1416,N_1373,N_1359);
xnor U1417 (N_1417,N_1338,N_1332);
xnor U1418 (N_1418,N_1331,N_1345);
xor U1419 (N_1419,N_1323,N_1360);
nor U1420 (N_1420,N_1326,N_1327);
and U1421 (N_1421,N_1329,N_1379);
and U1422 (N_1422,N_1329,N_1369);
xor U1423 (N_1423,N_1365,N_1373);
and U1424 (N_1424,N_1334,N_1363);
nor U1425 (N_1425,N_1373,N_1363);
xnor U1426 (N_1426,N_1360,N_1376);
or U1427 (N_1427,N_1369,N_1370);
and U1428 (N_1428,N_1330,N_1364);
and U1429 (N_1429,N_1338,N_1321);
xor U1430 (N_1430,N_1351,N_1340);
and U1431 (N_1431,N_1373,N_1335);
xnor U1432 (N_1432,N_1368,N_1339);
and U1433 (N_1433,N_1357,N_1343);
nand U1434 (N_1434,N_1343,N_1323);
or U1435 (N_1435,N_1337,N_1353);
and U1436 (N_1436,N_1335,N_1346);
xor U1437 (N_1437,N_1322,N_1346);
or U1438 (N_1438,N_1336,N_1347);
nand U1439 (N_1439,N_1333,N_1354);
or U1440 (N_1440,N_1385,N_1391);
nand U1441 (N_1441,N_1420,N_1390);
nand U1442 (N_1442,N_1395,N_1423);
nor U1443 (N_1443,N_1418,N_1387);
or U1444 (N_1444,N_1434,N_1439);
nor U1445 (N_1445,N_1436,N_1409);
or U1446 (N_1446,N_1405,N_1389);
or U1447 (N_1447,N_1414,N_1393);
nor U1448 (N_1448,N_1417,N_1431);
xnor U1449 (N_1449,N_1438,N_1402);
or U1450 (N_1450,N_1406,N_1386);
xor U1451 (N_1451,N_1419,N_1412);
nand U1452 (N_1452,N_1382,N_1411);
xnor U1453 (N_1453,N_1432,N_1429);
nor U1454 (N_1454,N_1433,N_1422);
or U1455 (N_1455,N_1384,N_1404);
nand U1456 (N_1456,N_1427,N_1407);
nand U1457 (N_1457,N_1383,N_1437);
xnor U1458 (N_1458,N_1413,N_1397);
nand U1459 (N_1459,N_1381,N_1415);
xor U1460 (N_1460,N_1401,N_1425);
xnor U1461 (N_1461,N_1403,N_1416);
xor U1462 (N_1462,N_1398,N_1426);
nor U1463 (N_1463,N_1435,N_1410);
nand U1464 (N_1464,N_1424,N_1400);
nand U1465 (N_1465,N_1388,N_1399);
nor U1466 (N_1466,N_1408,N_1421);
or U1467 (N_1467,N_1396,N_1392);
nand U1468 (N_1468,N_1394,N_1430);
or U1469 (N_1469,N_1380,N_1428);
or U1470 (N_1470,N_1399,N_1381);
nor U1471 (N_1471,N_1428,N_1381);
nor U1472 (N_1472,N_1404,N_1419);
and U1473 (N_1473,N_1414,N_1411);
or U1474 (N_1474,N_1438,N_1422);
nand U1475 (N_1475,N_1435,N_1401);
nor U1476 (N_1476,N_1382,N_1437);
nor U1477 (N_1477,N_1402,N_1415);
and U1478 (N_1478,N_1430,N_1439);
xor U1479 (N_1479,N_1391,N_1395);
nor U1480 (N_1480,N_1393,N_1434);
or U1481 (N_1481,N_1380,N_1399);
xor U1482 (N_1482,N_1426,N_1399);
nor U1483 (N_1483,N_1387,N_1424);
and U1484 (N_1484,N_1403,N_1436);
nor U1485 (N_1485,N_1386,N_1389);
nor U1486 (N_1486,N_1438,N_1421);
and U1487 (N_1487,N_1403,N_1417);
or U1488 (N_1488,N_1436,N_1407);
nor U1489 (N_1489,N_1416,N_1391);
nand U1490 (N_1490,N_1404,N_1383);
xor U1491 (N_1491,N_1408,N_1435);
xnor U1492 (N_1492,N_1412,N_1409);
and U1493 (N_1493,N_1391,N_1437);
and U1494 (N_1494,N_1429,N_1416);
or U1495 (N_1495,N_1434,N_1387);
or U1496 (N_1496,N_1439,N_1389);
nor U1497 (N_1497,N_1411,N_1401);
nand U1498 (N_1498,N_1407,N_1403);
and U1499 (N_1499,N_1436,N_1399);
nor U1500 (N_1500,N_1468,N_1475);
nor U1501 (N_1501,N_1498,N_1465);
nand U1502 (N_1502,N_1476,N_1446);
and U1503 (N_1503,N_1488,N_1491);
or U1504 (N_1504,N_1455,N_1452);
nand U1505 (N_1505,N_1444,N_1490);
and U1506 (N_1506,N_1449,N_1471);
nor U1507 (N_1507,N_1442,N_1457);
nor U1508 (N_1508,N_1484,N_1494);
nand U1509 (N_1509,N_1461,N_1473);
xnor U1510 (N_1510,N_1458,N_1479);
or U1511 (N_1511,N_1443,N_1453);
nor U1512 (N_1512,N_1451,N_1464);
nand U1513 (N_1513,N_1497,N_1489);
and U1514 (N_1514,N_1472,N_1496);
and U1515 (N_1515,N_1447,N_1478);
and U1516 (N_1516,N_1460,N_1492);
and U1517 (N_1517,N_1466,N_1467);
nand U1518 (N_1518,N_1495,N_1469);
nand U1519 (N_1519,N_1493,N_1450);
nand U1520 (N_1520,N_1456,N_1487);
or U1521 (N_1521,N_1459,N_1463);
and U1522 (N_1522,N_1441,N_1499);
or U1523 (N_1523,N_1462,N_1448);
nor U1524 (N_1524,N_1480,N_1482);
xnor U1525 (N_1525,N_1477,N_1474);
and U1526 (N_1526,N_1470,N_1486);
or U1527 (N_1527,N_1483,N_1485);
nand U1528 (N_1528,N_1454,N_1481);
xor U1529 (N_1529,N_1445,N_1440);
nand U1530 (N_1530,N_1458,N_1493);
nand U1531 (N_1531,N_1488,N_1451);
xnor U1532 (N_1532,N_1480,N_1453);
or U1533 (N_1533,N_1466,N_1445);
or U1534 (N_1534,N_1453,N_1490);
nand U1535 (N_1535,N_1453,N_1449);
nand U1536 (N_1536,N_1488,N_1499);
and U1537 (N_1537,N_1467,N_1495);
xnor U1538 (N_1538,N_1489,N_1462);
and U1539 (N_1539,N_1477,N_1489);
or U1540 (N_1540,N_1455,N_1468);
and U1541 (N_1541,N_1474,N_1498);
nor U1542 (N_1542,N_1444,N_1448);
and U1543 (N_1543,N_1479,N_1478);
xor U1544 (N_1544,N_1495,N_1470);
or U1545 (N_1545,N_1448,N_1454);
and U1546 (N_1546,N_1461,N_1494);
and U1547 (N_1547,N_1493,N_1483);
nor U1548 (N_1548,N_1477,N_1444);
or U1549 (N_1549,N_1486,N_1462);
nand U1550 (N_1550,N_1488,N_1445);
or U1551 (N_1551,N_1472,N_1443);
nand U1552 (N_1552,N_1494,N_1455);
nor U1553 (N_1553,N_1461,N_1480);
nor U1554 (N_1554,N_1487,N_1474);
xnor U1555 (N_1555,N_1440,N_1451);
nand U1556 (N_1556,N_1484,N_1445);
nand U1557 (N_1557,N_1462,N_1493);
or U1558 (N_1558,N_1461,N_1471);
nand U1559 (N_1559,N_1490,N_1446);
nand U1560 (N_1560,N_1523,N_1554);
nand U1561 (N_1561,N_1545,N_1533);
and U1562 (N_1562,N_1516,N_1542);
xnor U1563 (N_1563,N_1546,N_1550);
nand U1564 (N_1564,N_1514,N_1559);
and U1565 (N_1565,N_1553,N_1500);
nor U1566 (N_1566,N_1515,N_1518);
nand U1567 (N_1567,N_1510,N_1557);
xnor U1568 (N_1568,N_1535,N_1501);
nor U1569 (N_1569,N_1509,N_1525);
and U1570 (N_1570,N_1544,N_1555);
xnor U1571 (N_1571,N_1541,N_1522);
nand U1572 (N_1572,N_1539,N_1543);
xnor U1573 (N_1573,N_1504,N_1540);
nor U1574 (N_1574,N_1506,N_1538);
or U1575 (N_1575,N_1521,N_1532);
nor U1576 (N_1576,N_1537,N_1520);
or U1577 (N_1577,N_1558,N_1508);
xor U1578 (N_1578,N_1551,N_1531);
nor U1579 (N_1579,N_1517,N_1505);
nor U1580 (N_1580,N_1502,N_1529);
and U1581 (N_1581,N_1524,N_1536);
xnor U1582 (N_1582,N_1548,N_1552);
nand U1583 (N_1583,N_1507,N_1511);
or U1584 (N_1584,N_1549,N_1547);
or U1585 (N_1585,N_1556,N_1534);
nand U1586 (N_1586,N_1530,N_1527);
or U1587 (N_1587,N_1513,N_1512);
and U1588 (N_1588,N_1503,N_1519);
and U1589 (N_1589,N_1528,N_1526);
nand U1590 (N_1590,N_1537,N_1559);
nand U1591 (N_1591,N_1540,N_1514);
or U1592 (N_1592,N_1510,N_1508);
or U1593 (N_1593,N_1558,N_1537);
nand U1594 (N_1594,N_1515,N_1549);
xor U1595 (N_1595,N_1505,N_1547);
xnor U1596 (N_1596,N_1549,N_1502);
or U1597 (N_1597,N_1518,N_1542);
and U1598 (N_1598,N_1557,N_1530);
xor U1599 (N_1599,N_1503,N_1546);
and U1600 (N_1600,N_1509,N_1521);
and U1601 (N_1601,N_1526,N_1502);
nand U1602 (N_1602,N_1535,N_1523);
nand U1603 (N_1603,N_1552,N_1524);
nand U1604 (N_1604,N_1534,N_1503);
and U1605 (N_1605,N_1548,N_1555);
xnor U1606 (N_1606,N_1533,N_1528);
xor U1607 (N_1607,N_1541,N_1516);
nor U1608 (N_1608,N_1500,N_1556);
nor U1609 (N_1609,N_1520,N_1503);
or U1610 (N_1610,N_1527,N_1516);
nor U1611 (N_1611,N_1529,N_1546);
nor U1612 (N_1612,N_1531,N_1506);
nor U1613 (N_1613,N_1533,N_1511);
and U1614 (N_1614,N_1529,N_1528);
or U1615 (N_1615,N_1519,N_1545);
and U1616 (N_1616,N_1528,N_1515);
and U1617 (N_1617,N_1509,N_1546);
and U1618 (N_1618,N_1535,N_1550);
nand U1619 (N_1619,N_1541,N_1523);
or U1620 (N_1620,N_1604,N_1606);
xnor U1621 (N_1621,N_1580,N_1605);
and U1622 (N_1622,N_1567,N_1612);
or U1623 (N_1623,N_1594,N_1618);
xnor U1624 (N_1624,N_1592,N_1600);
nor U1625 (N_1625,N_1617,N_1581);
or U1626 (N_1626,N_1583,N_1599);
or U1627 (N_1627,N_1601,N_1602);
xnor U1628 (N_1628,N_1570,N_1609);
nand U1629 (N_1629,N_1582,N_1608);
xnor U1630 (N_1630,N_1571,N_1588);
nor U1631 (N_1631,N_1607,N_1564);
nand U1632 (N_1632,N_1560,N_1593);
xnor U1633 (N_1633,N_1591,N_1614);
nor U1634 (N_1634,N_1586,N_1578);
or U1635 (N_1635,N_1585,N_1579);
and U1636 (N_1636,N_1597,N_1561);
and U1637 (N_1637,N_1562,N_1603);
and U1638 (N_1638,N_1573,N_1566);
xnor U1639 (N_1639,N_1596,N_1610);
xnor U1640 (N_1640,N_1569,N_1568);
nor U1641 (N_1641,N_1587,N_1598);
nor U1642 (N_1642,N_1572,N_1576);
nor U1643 (N_1643,N_1574,N_1616);
and U1644 (N_1644,N_1584,N_1563);
and U1645 (N_1645,N_1589,N_1590);
or U1646 (N_1646,N_1611,N_1595);
nor U1647 (N_1647,N_1613,N_1565);
or U1648 (N_1648,N_1619,N_1615);
and U1649 (N_1649,N_1577,N_1575);
and U1650 (N_1650,N_1575,N_1607);
nand U1651 (N_1651,N_1593,N_1607);
xnor U1652 (N_1652,N_1596,N_1578);
nand U1653 (N_1653,N_1569,N_1579);
nor U1654 (N_1654,N_1586,N_1572);
and U1655 (N_1655,N_1615,N_1570);
nand U1656 (N_1656,N_1613,N_1560);
or U1657 (N_1657,N_1586,N_1607);
and U1658 (N_1658,N_1616,N_1603);
xnor U1659 (N_1659,N_1611,N_1592);
xor U1660 (N_1660,N_1592,N_1560);
nand U1661 (N_1661,N_1603,N_1596);
nor U1662 (N_1662,N_1581,N_1605);
and U1663 (N_1663,N_1590,N_1603);
or U1664 (N_1664,N_1598,N_1609);
nor U1665 (N_1665,N_1611,N_1615);
xnor U1666 (N_1666,N_1614,N_1596);
or U1667 (N_1667,N_1562,N_1567);
and U1668 (N_1668,N_1601,N_1567);
nor U1669 (N_1669,N_1599,N_1604);
nor U1670 (N_1670,N_1566,N_1608);
and U1671 (N_1671,N_1577,N_1611);
nor U1672 (N_1672,N_1619,N_1569);
nand U1673 (N_1673,N_1569,N_1567);
xor U1674 (N_1674,N_1594,N_1599);
nand U1675 (N_1675,N_1593,N_1617);
and U1676 (N_1676,N_1588,N_1609);
or U1677 (N_1677,N_1564,N_1563);
nand U1678 (N_1678,N_1572,N_1589);
or U1679 (N_1679,N_1614,N_1609);
nor U1680 (N_1680,N_1670,N_1648);
nor U1681 (N_1681,N_1661,N_1639);
or U1682 (N_1682,N_1677,N_1620);
and U1683 (N_1683,N_1638,N_1654);
or U1684 (N_1684,N_1676,N_1656);
and U1685 (N_1685,N_1640,N_1624);
and U1686 (N_1686,N_1631,N_1663);
xnor U1687 (N_1687,N_1622,N_1675);
nor U1688 (N_1688,N_1671,N_1627);
or U1689 (N_1689,N_1664,N_1672);
nand U1690 (N_1690,N_1621,N_1626);
nand U1691 (N_1691,N_1643,N_1674);
nor U1692 (N_1692,N_1655,N_1635);
or U1693 (N_1693,N_1628,N_1657);
and U1694 (N_1694,N_1641,N_1650);
nand U1695 (N_1695,N_1679,N_1653);
nor U1696 (N_1696,N_1630,N_1652);
or U1697 (N_1697,N_1649,N_1658);
nand U1698 (N_1698,N_1666,N_1642);
nor U1699 (N_1699,N_1623,N_1665);
and U1700 (N_1700,N_1646,N_1669);
xor U1701 (N_1701,N_1636,N_1659);
nand U1702 (N_1702,N_1662,N_1637);
or U1703 (N_1703,N_1678,N_1629);
and U1704 (N_1704,N_1647,N_1644);
and U1705 (N_1705,N_1634,N_1667);
or U1706 (N_1706,N_1660,N_1632);
nand U1707 (N_1707,N_1625,N_1668);
xor U1708 (N_1708,N_1633,N_1645);
nand U1709 (N_1709,N_1651,N_1673);
or U1710 (N_1710,N_1637,N_1666);
nor U1711 (N_1711,N_1664,N_1676);
and U1712 (N_1712,N_1677,N_1630);
or U1713 (N_1713,N_1643,N_1647);
or U1714 (N_1714,N_1621,N_1660);
or U1715 (N_1715,N_1625,N_1632);
nand U1716 (N_1716,N_1653,N_1660);
nand U1717 (N_1717,N_1657,N_1671);
nand U1718 (N_1718,N_1649,N_1661);
nand U1719 (N_1719,N_1642,N_1622);
nor U1720 (N_1720,N_1661,N_1660);
nor U1721 (N_1721,N_1678,N_1635);
nand U1722 (N_1722,N_1673,N_1626);
or U1723 (N_1723,N_1638,N_1668);
xnor U1724 (N_1724,N_1639,N_1664);
and U1725 (N_1725,N_1672,N_1648);
nand U1726 (N_1726,N_1642,N_1629);
or U1727 (N_1727,N_1645,N_1664);
and U1728 (N_1728,N_1664,N_1646);
and U1729 (N_1729,N_1672,N_1654);
or U1730 (N_1730,N_1674,N_1645);
nor U1731 (N_1731,N_1666,N_1623);
nand U1732 (N_1732,N_1638,N_1648);
nand U1733 (N_1733,N_1660,N_1641);
and U1734 (N_1734,N_1634,N_1656);
xor U1735 (N_1735,N_1640,N_1643);
nand U1736 (N_1736,N_1661,N_1652);
nor U1737 (N_1737,N_1665,N_1670);
or U1738 (N_1738,N_1651,N_1640);
and U1739 (N_1739,N_1625,N_1678);
nand U1740 (N_1740,N_1685,N_1691);
and U1741 (N_1741,N_1717,N_1683);
or U1742 (N_1742,N_1707,N_1710);
nand U1743 (N_1743,N_1693,N_1701);
and U1744 (N_1744,N_1720,N_1723);
nand U1745 (N_1745,N_1711,N_1688);
nand U1746 (N_1746,N_1715,N_1730);
nor U1747 (N_1747,N_1708,N_1719);
xnor U1748 (N_1748,N_1697,N_1726);
xor U1749 (N_1749,N_1692,N_1722);
xnor U1750 (N_1750,N_1729,N_1713);
and U1751 (N_1751,N_1680,N_1739);
or U1752 (N_1752,N_1738,N_1718);
nand U1753 (N_1753,N_1684,N_1706);
nor U1754 (N_1754,N_1734,N_1703);
nand U1755 (N_1755,N_1727,N_1698);
and U1756 (N_1756,N_1735,N_1716);
xnor U1757 (N_1757,N_1682,N_1686);
or U1758 (N_1758,N_1721,N_1705);
nor U1759 (N_1759,N_1704,N_1728);
or U1760 (N_1760,N_1731,N_1737);
and U1761 (N_1761,N_1689,N_1696);
and U1762 (N_1762,N_1714,N_1700);
nand U1763 (N_1763,N_1724,N_1681);
xor U1764 (N_1764,N_1736,N_1695);
xor U1765 (N_1765,N_1702,N_1709);
xnor U1766 (N_1766,N_1687,N_1733);
and U1767 (N_1767,N_1712,N_1699);
xor U1768 (N_1768,N_1690,N_1732);
or U1769 (N_1769,N_1694,N_1725);
and U1770 (N_1770,N_1736,N_1725);
nand U1771 (N_1771,N_1723,N_1721);
xor U1772 (N_1772,N_1736,N_1694);
xor U1773 (N_1773,N_1706,N_1716);
or U1774 (N_1774,N_1739,N_1697);
xnor U1775 (N_1775,N_1708,N_1711);
nand U1776 (N_1776,N_1685,N_1731);
and U1777 (N_1777,N_1712,N_1730);
nand U1778 (N_1778,N_1707,N_1732);
nand U1779 (N_1779,N_1731,N_1705);
nand U1780 (N_1780,N_1739,N_1685);
or U1781 (N_1781,N_1728,N_1691);
nand U1782 (N_1782,N_1704,N_1717);
xnor U1783 (N_1783,N_1727,N_1710);
nor U1784 (N_1784,N_1704,N_1731);
nor U1785 (N_1785,N_1703,N_1709);
or U1786 (N_1786,N_1698,N_1681);
nand U1787 (N_1787,N_1716,N_1738);
nor U1788 (N_1788,N_1713,N_1697);
and U1789 (N_1789,N_1720,N_1704);
or U1790 (N_1790,N_1720,N_1685);
nand U1791 (N_1791,N_1686,N_1716);
xor U1792 (N_1792,N_1685,N_1736);
and U1793 (N_1793,N_1739,N_1709);
or U1794 (N_1794,N_1682,N_1695);
and U1795 (N_1795,N_1697,N_1720);
or U1796 (N_1796,N_1731,N_1703);
xnor U1797 (N_1797,N_1731,N_1718);
or U1798 (N_1798,N_1718,N_1696);
xnor U1799 (N_1799,N_1689,N_1717);
or U1800 (N_1800,N_1770,N_1798);
or U1801 (N_1801,N_1777,N_1746);
nand U1802 (N_1802,N_1794,N_1781);
xor U1803 (N_1803,N_1747,N_1768);
nor U1804 (N_1804,N_1783,N_1766);
and U1805 (N_1805,N_1773,N_1771);
and U1806 (N_1806,N_1759,N_1740);
or U1807 (N_1807,N_1753,N_1760);
and U1808 (N_1808,N_1761,N_1755);
xor U1809 (N_1809,N_1792,N_1742);
or U1810 (N_1810,N_1790,N_1751);
or U1811 (N_1811,N_1752,N_1796);
xor U1812 (N_1812,N_1775,N_1793);
or U1813 (N_1813,N_1797,N_1787);
nand U1814 (N_1814,N_1757,N_1782);
and U1815 (N_1815,N_1799,N_1767);
or U1816 (N_1816,N_1764,N_1786);
or U1817 (N_1817,N_1785,N_1765);
and U1818 (N_1818,N_1788,N_1779);
nor U1819 (N_1819,N_1778,N_1743);
and U1820 (N_1820,N_1754,N_1784);
and U1821 (N_1821,N_1772,N_1744);
xnor U1822 (N_1822,N_1774,N_1758);
nand U1823 (N_1823,N_1749,N_1769);
and U1824 (N_1824,N_1776,N_1756);
or U1825 (N_1825,N_1750,N_1789);
or U1826 (N_1826,N_1762,N_1741);
xor U1827 (N_1827,N_1780,N_1763);
xor U1828 (N_1828,N_1795,N_1745);
nor U1829 (N_1829,N_1791,N_1748);
and U1830 (N_1830,N_1798,N_1780);
xnor U1831 (N_1831,N_1772,N_1755);
nand U1832 (N_1832,N_1793,N_1765);
xnor U1833 (N_1833,N_1745,N_1789);
and U1834 (N_1834,N_1747,N_1792);
nand U1835 (N_1835,N_1778,N_1771);
or U1836 (N_1836,N_1749,N_1798);
or U1837 (N_1837,N_1784,N_1747);
xor U1838 (N_1838,N_1786,N_1761);
or U1839 (N_1839,N_1741,N_1769);
xor U1840 (N_1840,N_1789,N_1746);
nand U1841 (N_1841,N_1781,N_1759);
and U1842 (N_1842,N_1778,N_1799);
nand U1843 (N_1843,N_1766,N_1751);
nor U1844 (N_1844,N_1793,N_1744);
nand U1845 (N_1845,N_1791,N_1772);
nor U1846 (N_1846,N_1775,N_1760);
xnor U1847 (N_1847,N_1780,N_1773);
nand U1848 (N_1848,N_1746,N_1758);
xor U1849 (N_1849,N_1761,N_1759);
and U1850 (N_1850,N_1783,N_1770);
and U1851 (N_1851,N_1758,N_1799);
nor U1852 (N_1852,N_1777,N_1773);
xnor U1853 (N_1853,N_1783,N_1795);
xnor U1854 (N_1854,N_1776,N_1792);
nand U1855 (N_1855,N_1767,N_1768);
and U1856 (N_1856,N_1769,N_1750);
xor U1857 (N_1857,N_1764,N_1742);
and U1858 (N_1858,N_1784,N_1751);
nand U1859 (N_1859,N_1751,N_1772);
and U1860 (N_1860,N_1827,N_1829);
or U1861 (N_1861,N_1819,N_1853);
or U1862 (N_1862,N_1816,N_1831);
and U1863 (N_1863,N_1802,N_1801);
and U1864 (N_1864,N_1840,N_1824);
nor U1865 (N_1865,N_1841,N_1825);
and U1866 (N_1866,N_1810,N_1805);
xnor U1867 (N_1867,N_1822,N_1848);
or U1868 (N_1868,N_1856,N_1804);
nor U1869 (N_1869,N_1823,N_1806);
xnor U1870 (N_1870,N_1812,N_1836);
and U1871 (N_1871,N_1844,N_1837);
nand U1872 (N_1872,N_1821,N_1814);
nand U1873 (N_1873,N_1855,N_1811);
and U1874 (N_1874,N_1859,N_1815);
xor U1875 (N_1875,N_1803,N_1832);
nor U1876 (N_1876,N_1843,N_1838);
and U1877 (N_1877,N_1851,N_1842);
or U1878 (N_1878,N_1833,N_1857);
nor U1879 (N_1879,N_1826,N_1813);
or U1880 (N_1880,N_1807,N_1830);
xnor U1881 (N_1881,N_1834,N_1817);
and U1882 (N_1882,N_1808,N_1847);
and U1883 (N_1883,N_1818,N_1846);
nand U1884 (N_1884,N_1820,N_1858);
nand U1885 (N_1885,N_1854,N_1852);
nor U1886 (N_1886,N_1828,N_1845);
or U1887 (N_1887,N_1809,N_1850);
nand U1888 (N_1888,N_1849,N_1835);
or U1889 (N_1889,N_1839,N_1800);
nor U1890 (N_1890,N_1844,N_1853);
or U1891 (N_1891,N_1811,N_1818);
nand U1892 (N_1892,N_1808,N_1840);
nand U1893 (N_1893,N_1844,N_1814);
nor U1894 (N_1894,N_1800,N_1829);
nand U1895 (N_1895,N_1840,N_1813);
and U1896 (N_1896,N_1822,N_1806);
nor U1897 (N_1897,N_1839,N_1815);
nor U1898 (N_1898,N_1859,N_1857);
nor U1899 (N_1899,N_1800,N_1811);
nand U1900 (N_1900,N_1856,N_1820);
or U1901 (N_1901,N_1810,N_1822);
and U1902 (N_1902,N_1859,N_1852);
nor U1903 (N_1903,N_1835,N_1807);
or U1904 (N_1904,N_1834,N_1806);
nand U1905 (N_1905,N_1820,N_1833);
and U1906 (N_1906,N_1823,N_1803);
and U1907 (N_1907,N_1820,N_1821);
xor U1908 (N_1908,N_1845,N_1859);
nor U1909 (N_1909,N_1846,N_1814);
xor U1910 (N_1910,N_1853,N_1800);
or U1911 (N_1911,N_1858,N_1804);
xor U1912 (N_1912,N_1845,N_1847);
or U1913 (N_1913,N_1844,N_1834);
nand U1914 (N_1914,N_1814,N_1852);
nand U1915 (N_1915,N_1834,N_1832);
nor U1916 (N_1916,N_1801,N_1839);
nor U1917 (N_1917,N_1813,N_1851);
nand U1918 (N_1918,N_1850,N_1842);
nor U1919 (N_1919,N_1848,N_1849);
xor U1920 (N_1920,N_1874,N_1902);
nand U1921 (N_1921,N_1914,N_1896);
nand U1922 (N_1922,N_1911,N_1870);
nand U1923 (N_1923,N_1897,N_1910);
nand U1924 (N_1924,N_1887,N_1881);
xnor U1925 (N_1925,N_1886,N_1869);
xor U1926 (N_1926,N_1891,N_1871);
or U1927 (N_1927,N_1862,N_1905);
nand U1928 (N_1928,N_1916,N_1912);
nand U1929 (N_1929,N_1861,N_1909);
and U1930 (N_1930,N_1898,N_1888);
or U1931 (N_1931,N_1892,N_1868);
xnor U1932 (N_1932,N_1913,N_1900);
nand U1933 (N_1933,N_1878,N_1873);
xnor U1934 (N_1934,N_1884,N_1893);
nor U1935 (N_1935,N_1882,N_1895);
and U1936 (N_1936,N_1894,N_1903);
and U1937 (N_1937,N_1907,N_1879);
and U1938 (N_1938,N_1908,N_1899);
xnor U1939 (N_1939,N_1901,N_1876);
nand U1940 (N_1940,N_1906,N_1883);
xor U1941 (N_1941,N_1915,N_1918);
xor U1942 (N_1942,N_1917,N_1865);
or U1943 (N_1943,N_1889,N_1866);
nor U1944 (N_1944,N_1890,N_1860);
nand U1945 (N_1945,N_1904,N_1919);
xnor U1946 (N_1946,N_1875,N_1864);
nand U1947 (N_1947,N_1863,N_1867);
or U1948 (N_1948,N_1880,N_1885);
or U1949 (N_1949,N_1877,N_1872);
nor U1950 (N_1950,N_1919,N_1863);
or U1951 (N_1951,N_1886,N_1885);
or U1952 (N_1952,N_1898,N_1875);
and U1953 (N_1953,N_1904,N_1908);
and U1954 (N_1954,N_1863,N_1888);
and U1955 (N_1955,N_1919,N_1898);
and U1956 (N_1956,N_1903,N_1896);
nand U1957 (N_1957,N_1880,N_1878);
nor U1958 (N_1958,N_1870,N_1900);
nor U1959 (N_1959,N_1893,N_1903);
nand U1960 (N_1960,N_1887,N_1865);
nor U1961 (N_1961,N_1898,N_1871);
nor U1962 (N_1962,N_1864,N_1907);
nand U1963 (N_1963,N_1908,N_1874);
and U1964 (N_1964,N_1868,N_1870);
and U1965 (N_1965,N_1906,N_1865);
xnor U1966 (N_1966,N_1887,N_1907);
and U1967 (N_1967,N_1893,N_1913);
and U1968 (N_1968,N_1878,N_1917);
nand U1969 (N_1969,N_1862,N_1861);
xnor U1970 (N_1970,N_1890,N_1914);
and U1971 (N_1971,N_1914,N_1866);
nand U1972 (N_1972,N_1896,N_1900);
or U1973 (N_1973,N_1908,N_1905);
xor U1974 (N_1974,N_1889,N_1902);
and U1975 (N_1975,N_1881,N_1861);
or U1976 (N_1976,N_1867,N_1870);
or U1977 (N_1977,N_1893,N_1911);
and U1978 (N_1978,N_1898,N_1896);
xnor U1979 (N_1979,N_1897,N_1888);
nand U1980 (N_1980,N_1958,N_1944);
nand U1981 (N_1981,N_1923,N_1946);
nand U1982 (N_1982,N_1976,N_1974);
and U1983 (N_1983,N_1948,N_1934);
nor U1984 (N_1984,N_1977,N_1975);
xor U1985 (N_1985,N_1969,N_1978);
xnor U1986 (N_1986,N_1964,N_1965);
nand U1987 (N_1987,N_1928,N_1941);
and U1988 (N_1988,N_1952,N_1956);
nor U1989 (N_1989,N_1935,N_1972);
and U1990 (N_1990,N_1945,N_1979);
or U1991 (N_1991,N_1943,N_1937);
nand U1992 (N_1992,N_1968,N_1921);
nor U1993 (N_1993,N_1925,N_1930);
nand U1994 (N_1994,N_1924,N_1966);
and U1995 (N_1995,N_1962,N_1920);
xor U1996 (N_1996,N_1971,N_1954);
xor U1997 (N_1997,N_1960,N_1957);
nand U1998 (N_1998,N_1953,N_1931);
nor U1999 (N_1999,N_1951,N_1947);
nand U2000 (N_2000,N_1959,N_1932);
and U2001 (N_2001,N_1967,N_1940);
nor U2002 (N_2002,N_1939,N_1970);
xnor U2003 (N_2003,N_1942,N_1950);
nand U2004 (N_2004,N_1949,N_1926);
or U2005 (N_2005,N_1933,N_1938);
and U2006 (N_2006,N_1922,N_1929);
xor U2007 (N_2007,N_1973,N_1961);
xnor U2008 (N_2008,N_1936,N_1955);
or U2009 (N_2009,N_1927,N_1963);
xor U2010 (N_2010,N_1946,N_1920);
nand U2011 (N_2011,N_1937,N_1967);
and U2012 (N_2012,N_1962,N_1933);
xor U2013 (N_2013,N_1977,N_1927);
or U2014 (N_2014,N_1929,N_1930);
or U2015 (N_2015,N_1957,N_1922);
or U2016 (N_2016,N_1971,N_1961);
nor U2017 (N_2017,N_1929,N_1953);
xnor U2018 (N_2018,N_1951,N_1935);
xor U2019 (N_2019,N_1953,N_1937);
or U2020 (N_2020,N_1957,N_1925);
and U2021 (N_2021,N_1953,N_1955);
nand U2022 (N_2022,N_1962,N_1923);
xnor U2023 (N_2023,N_1975,N_1953);
nor U2024 (N_2024,N_1952,N_1950);
nand U2025 (N_2025,N_1978,N_1972);
nor U2026 (N_2026,N_1950,N_1969);
xor U2027 (N_2027,N_1965,N_1979);
nor U2028 (N_2028,N_1928,N_1936);
or U2029 (N_2029,N_1949,N_1951);
nand U2030 (N_2030,N_1974,N_1950);
nor U2031 (N_2031,N_1973,N_1977);
or U2032 (N_2032,N_1929,N_1964);
and U2033 (N_2033,N_1957,N_1926);
or U2034 (N_2034,N_1933,N_1974);
and U2035 (N_2035,N_1955,N_1971);
nor U2036 (N_2036,N_1955,N_1939);
nor U2037 (N_2037,N_1969,N_1947);
nor U2038 (N_2038,N_1937,N_1932);
and U2039 (N_2039,N_1967,N_1944);
nand U2040 (N_2040,N_2014,N_1991);
or U2041 (N_2041,N_1985,N_2010);
and U2042 (N_2042,N_2027,N_1980);
and U2043 (N_2043,N_2018,N_1999);
nand U2044 (N_2044,N_2008,N_1981);
xnor U2045 (N_2045,N_2036,N_2023);
xnor U2046 (N_2046,N_1996,N_2009);
and U2047 (N_2047,N_1994,N_1989);
and U2048 (N_2048,N_2028,N_2004);
nand U2049 (N_2049,N_1986,N_2012);
xnor U2050 (N_2050,N_1982,N_2031);
xor U2051 (N_2051,N_2029,N_1988);
and U2052 (N_2052,N_2000,N_2003);
and U2053 (N_2053,N_2019,N_2035);
or U2054 (N_2054,N_2039,N_1998);
or U2055 (N_2055,N_1987,N_2017);
xnor U2056 (N_2056,N_1992,N_1990);
or U2057 (N_2057,N_2015,N_2026);
xnor U2058 (N_2058,N_2025,N_1995);
xor U2059 (N_2059,N_2032,N_2034);
nand U2060 (N_2060,N_2022,N_2038);
nor U2061 (N_2061,N_2005,N_2021);
nor U2062 (N_2062,N_2006,N_2016);
xor U2063 (N_2063,N_2037,N_2013);
xnor U2064 (N_2064,N_1993,N_2001);
xnor U2065 (N_2065,N_1984,N_1997);
or U2066 (N_2066,N_1983,N_2030);
nand U2067 (N_2067,N_2007,N_2020);
and U2068 (N_2068,N_2024,N_2011);
xnor U2069 (N_2069,N_2002,N_2033);
xnor U2070 (N_2070,N_2007,N_2028);
xor U2071 (N_2071,N_2008,N_2004);
nand U2072 (N_2072,N_2003,N_2013);
xor U2073 (N_2073,N_1996,N_2017);
or U2074 (N_2074,N_1986,N_2034);
or U2075 (N_2075,N_2027,N_1995);
nor U2076 (N_2076,N_2019,N_2018);
and U2077 (N_2077,N_2015,N_1983);
nand U2078 (N_2078,N_1991,N_2015);
xnor U2079 (N_2079,N_1982,N_2036);
nand U2080 (N_2080,N_1997,N_1989);
xor U2081 (N_2081,N_1981,N_2011);
and U2082 (N_2082,N_1998,N_2035);
xnor U2083 (N_2083,N_2011,N_2021);
xor U2084 (N_2084,N_1985,N_1987);
nand U2085 (N_2085,N_2014,N_1983);
and U2086 (N_2086,N_2012,N_2025);
or U2087 (N_2087,N_2025,N_1983);
xor U2088 (N_2088,N_1998,N_2005);
nand U2089 (N_2089,N_2016,N_1981);
and U2090 (N_2090,N_2022,N_2017);
nor U2091 (N_2091,N_1981,N_1999);
and U2092 (N_2092,N_1996,N_2039);
or U2093 (N_2093,N_1991,N_1999);
and U2094 (N_2094,N_1990,N_2023);
and U2095 (N_2095,N_2020,N_2029);
xnor U2096 (N_2096,N_1984,N_1980);
and U2097 (N_2097,N_2022,N_2034);
and U2098 (N_2098,N_1981,N_2009);
xor U2099 (N_2099,N_2012,N_1989);
nand U2100 (N_2100,N_2077,N_2070);
nand U2101 (N_2101,N_2096,N_2092);
or U2102 (N_2102,N_2043,N_2085);
or U2103 (N_2103,N_2055,N_2069);
xnor U2104 (N_2104,N_2044,N_2057);
or U2105 (N_2105,N_2050,N_2041);
nand U2106 (N_2106,N_2068,N_2079);
nor U2107 (N_2107,N_2058,N_2062);
nand U2108 (N_2108,N_2088,N_2098);
and U2109 (N_2109,N_2054,N_2082);
xor U2110 (N_2110,N_2087,N_2099);
or U2111 (N_2111,N_2076,N_2074);
and U2112 (N_2112,N_2046,N_2078);
nor U2113 (N_2113,N_2095,N_2042);
nor U2114 (N_2114,N_2056,N_2093);
nand U2115 (N_2115,N_2049,N_2045);
and U2116 (N_2116,N_2047,N_2090);
nor U2117 (N_2117,N_2052,N_2053);
xnor U2118 (N_2118,N_2064,N_2091);
xnor U2119 (N_2119,N_2073,N_2083);
nand U2120 (N_2120,N_2048,N_2060);
or U2121 (N_2121,N_2094,N_2097);
nand U2122 (N_2122,N_2086,N_2089);
or U2123 (N_2123,N_2061,N_2040);
and U2124 (N_2124,N_2066,N_2063);
nand U2125 (N_2125,N_2075,N_2071);
xnor U2126 (N_2126,N_2059,N_2067);
nand U2127 (N_2127,N_2072,N_2051);
nor U2128 (N_2128,N_2065,N_2084);
or U2129 (N_2129,N_2081,N_2080);
xnor U2130 (N_2130,N_2080,N_2042);
nor U2131 (N_2131,N_2096,N_2089);
or U2132 (N_2132,N_2043,N_2076);
nor U2133 (N_2133,N_2085,N_2099);
xor U2134 (N_2134,N_2098,N_2054);
or U2135 (N_2135,N_2048,N_2044);
and U2136 (N_2136,N_2089,N_2064);
nand U2137 (N_2137,N_2079,N_2064);
or U2138 (N_2138,N_2055,N_2084);
nor U2139 (N_2139,N_2083,N_2055);
nor U2140 (N_2140,N_2049,N_2050);
xnor U2141 (N_2141,N_2090,N_2050);
nor U2142 (N_2142,N_2040,N_2087);
nand U2143 (N_2143,N_2059,N_2076);
nor U2144 (N_2144,N_2055,N_2079);
or U2145 (N_2145,N_2077,N_2097);
nand U2146 (N_2146,N_2041,N_2040);
nor U2147 (N_2147,N_2070,N_2042);
nor U2148 (N_2148,N_2074,N_2077);
or U2149 (N_2149,N_2085,N_2088);
nand U2150 (N_2150,N_2047,N_2083);
nand U2151 (N_2151,N_2051,N_2067);
xor U2152 (N_2152,N_2093,N_2079);
xnor U2153 (N_2153,N_2069,N_2049);
nand U2154 (N_2154,N_2050,N_2076);
or U2155 (N_2155,N_2093,N_2054);
xnor U2156 (N_2156,N_2052,N_2043);
nor U2157 (N_2157,N_2079,N_2087);
or U2158 (N_2158,N_2045,N_2071);
xnor U2159 (N_2159,N_2083,N_2085);
nor U2160 (N_2160,N_2125,N_2123);
xor U2161 (N_2161,N_2127,N_2143);
and U2162 (N_2162,N_2140,N_2139);
nor U2163 (N_2163,N_2119,N_2122);
or U2164 (N_2164,N_2142,N_2155);
xor U2165 (N_2165,N_2103,N_2128);
or U2166 (N_2166,N_2151,N_2144);
or U2167 (N_2167,N_2115,N_2135);
nor U2168 (N_2168,N_2113,N_2137);
xnor U2169 (N_2169,N_2129,N_2141);
nor U2170 (N_2170,N_2105,N_2159);
xor U2171 (N_2171,N_2156,N_2118);
xor U2172 (N_2172,N_2117,N_2146);
nand U2173 (N_2173,N_2110,N_2107);
and U2174 (N_2174,N_2104,N_2111);
and U2175 (N_2175,N_2112,N_2130);
and U2176 (N_2176,N_2114,N_2138);
nand U2177 (N_2177,N_2101,N_2157);
nand U2178 (N_2178,N_2136,N_2108);
and U2179 (N_2179,N_2106,N_2132);
nand U2180 (N_2180,N_2148,N_2120);
xor U2181 (N_2181,N_2154,N_2124);
xnor U2182 (N_2182,N_2116,N_2149);
xnor U2183 (N_2183,N_2109,N_2153);
nor U2184 (N_2184,N_2102,N_2150);
and U2185 (N_2185,N_2158,N_2145);
or U2186 (N_2186,N_2131,N_2100);
xnor U2187 (N_2187,N_2126,N_2134);
nand U2188 (N_2188,N_2152,N_2133);
nand U2189 (N_2189,N_2147,N_2121);
and U2190 (N_2190,N_2130,N_2158);
or U2191 (N_2191,N_2137,N_2120);
and U2192 (N_2192,N_2159,N_2122);
and U2193 (N_2193,N_2145,N_2141);
and U2194 (N_2194,N_2115,N_2114);
or U2195 (N_2195,N_2135,N_2149);
and U2196 (N_2196,N_2120,N_2128);
or U2197 (N_2197,N_2152,N_2159);
nand U2198 (N_2198,N_2132,N_2139);
and U2199 (N_2199,N_2156,N_2115);
nand U2200 (N_2200,N_2134,N_2141);
nor U2201 (N_2201,N_2137,N_2157);
or U2202 (N_2202,N_2110,N_2140);
xnor U2203 (N_2203,N_2156,N_2144);
nor U2204 (N_2204,N_2150,N_2141);
or U2205 (N_2205,N_2101,N_2146);
and U2206 (N_2206,N_2122,N_2137);
nor U2207 (N_2207,N_2101,N_2136);
nand U2208 (N_2208,N_2136,N_2141);
or U2209 (N_2209,N_2138,N_2107);
and U2210 (N_2210,N_2154,N_2139);
or U2211 (N_2211,N_2104,N_2133);
xnor U2212 (N_2212,N_2157,N_2109);
xnor U2213 (N_2213,N_2112,N_2157);
nor U2214 (N_2214,N_2150,N_2103);
and U2215 (N_2215,N_2123,N_2159);
or U2216 (N_2216,N_2142,N_2111);
nand U2217 (N_2217,N_2135,N_2125);
xnor U2218 (N_2218,N_2102,N_2121);
and U2219 (N_2219,N_2155,N_2136);
or U2220 (N_2220,N_2208,N_2195);
and U2221 (N_2221,N_2201,N_2165);
nor U2222 (N_2222,N_2160,N_2209);
and U2223 (N_2223,N_2188,N_2210);
and U2224 (N_2224,N_2163,N_2211);
xor U2225 (N_2225,N_2170,N_2178);
nor U2226 (N_2226,N_2184,N_2202);
xnor U2227 (N_2227,N_2193,N_2200);
nor U2228 (N_2228,N_2179,N_2181);
or U2229 (N_2229,N_2186,N_2167);
or U2230 (N_2230,N_2171,N_2174);
xnor U2231 (N_2231,N_2176,N_2198);
xor U2232 (N_2232,N_2187,N_2215);
nand U2233 (N_2233,N_2204,N_2207);
or U2234 (N_2234,N_2216,N_2197);
nand U2235 (N_2235,N_2203,N_2166);
nor U2236 (N_2236,N_2199,N_2190);
or U2237 (N_2237,N_2189,N_2194);
nand U2238 (N_2238,N_2191,N_2213);
or U2239 (N_2239,N_2183,N_2175);
nor U2240 (N_2240,N_2185,N_2219);
or U2241 (N_2241,N_2172,N_2180);
nor U2242 (N_2242,N_2212,N_2217);
or U2243 (N_2243,N_2164,N_2218);
xnor U2244 (N_2244,N_2192,N_2168);
xor U2245 (N_2245,N_2214,N_2173);
nor U2246 (N_2246,N_2169,N_2205);
nand U2247 (N_2247,N_2196,N_2177);
or U2248 (N_2248,N_2206,N_2162);
and U2249 (N_2249,N_2161,N_2182);
or U2250 (N_2250,N_2200,N_2186);
nand U2251 (N_2251,N_2173,N_2211);
xnor U2252 (N_2252,N_2210,N_2189);
xor U2253 (N_2253,N_2170,N_2194);
nand U2254 (N_2254,N_2208,N_2199);
or U2255 (N_2255,N_2171,N_2161);
nand U2256 (N_2256,N_2201,N_2175);
nor U2257 (N_2257,N_2185,N_2210);
or U2258 (N_2258,N_2199,N_2212);
or U2259 (N_2259,N_2193,N_2197);
and U2260 (N_2260,N_2189,N_2162);
or U2261 (N_2261,N_2214,N_2216);
nor U2262 (N_2262,N_2205,N_2185);
or U2263 (N_2263,N_2162,N_2213);
nand U2264 (N_2264,N_2197,N_2160);
and U2265 (N_2265,N_2175,N_2161);
and U2266 (N_2266,N_2170,N_2161);
or U2267 (N_2267,N_2201,N_2212);
and U2268 (N_2268,N_2163,N_2193);
xor U2269 (N_2269,N_2178,N_2198);
nand U2270 (N_2270,N_2176,N_2197);
nor U2271 (N_2271,N_2176,N_2160);
xnor U2272 (N_2272,N_2166,N_2176);
or U2273 (N_2273,N_2187,N_2217);
and U2274 (N_2274,N_2168,N_2176);
nand U2275 (N_2275,N_2176,N_2202);
or U2276 (N_2276,N_2174,N_2180);
nor U2277 (N_2277,N_2186,N_2197);
nor U2278 (N_2278,N_2196,N_2215);
xnor U2279 (N_2279,N_2211,N_2189);
nand U2280 (N_2280,N_2243,N_2275);
nand U2281 (N_2281,N_2274,N_2263);
nand U2282 (N_2282,N_2276,N_2236);
nor U2283 (N_2283,N_2262,N_2251);
and U2284 (N_2284,N_2278,N_2220);
nand U2285 (N_2285,N_2268,N_2258);
nor U2286 (N_2286,N_2272,N_2230);
nand U2287 (N_2287,N_2250,N_2273);
xor U2288 (N_2288,N_2223,N_2247);
or U2289 (N_2289,N_2253,N_2226);
and U2290 (N_2290,N_2241,N_2269);
xor U2291 (N_2291,N_2237,N_2249);
xor U2292 (N_2292,N_2261,N_2225);
xor U2293 (N_2293,N_2232,N_2246);
nor U2294 (N_2294,N_2270,N_2227);
and U2295 (N_2295,N_2234,N_2245);
nor U2296 (N_2296,N_2277,N_2233);
nor U2297 (N_2297,N_2267,N_2231);
nand U2298 (N_2298,N_2254,N_2228);
nand U2299 (N_2299,N_2240,N_2279);
or U2300 (N_2300,N_2256,N_2252);
xor U2301 (N_2301,N_2235,N_2264);
or U2302 (N_2302,N_2239,N_2222);
nor U2303 (N_2303,N_2221,N_2242);
nor U2304 (N_2304,N_2265,N_2257);
xnor U2305 (N_2305,N_2244,N_2255);
xor U2306 (N_2306,N_2224,N_2238);
and U2307 (N_2307,N_2229,N_2266);
and U2308 (N_2308,N_2248,N_2271);
nor U2309 (N_2309,N_2260,N_2259);
or U2310 (N_2310,N_2270,N_2239);
or U2311 (N_2311,N_2256,N_2254);
or U2312 (N_2312,N_2260,N_2242);
and U2313 (N_2313,N_2251,N_2250);
xor U2314 (N_2314,N_2278,N_2250);
and U2315 (N_2315,N_2277,N_2266);
nor U2316 (N_2316,N_2244,N_2242);
nor U2317 (N_2317,N_2259,N_2227);
nor U2318 (N_2318,N_2265,N_2274);
and U2319 (N_2319,N_2249,N_2251);
or U2320 (N_2320,N_2266,N_2275);
and U2321 (N_2321,N_2241,N_2220);
nand U2322 (N_2322,N_2256,N_2243);
nand U2323 (N_2323,N_2247,N_2251);
nand U2324 (N_2324,N_2238,N_2241);
nand U2325 (N_2325,N_2263,N_2243);
nor U2326 (N_2326,N_2232,N_2240);
and U2327 (N_2327,N_2270,N_2255);
and U2328 (N_2328,N_2261,N_2239);
nand U2329 (N_2329,N_2239,N_2245);
xnor U2330 (N_2330,N_2234,N_2264);
xor U2331 (N_2331,N_2234,N_2267);
and U2332 (N_2332,N_2253,N_2229);
nand U2333 (N_2333,N_2274,N_2252);
nor U2334 (N_2334,N_2223,N_2227);
xor U2335 (N_2335,N_2273,N_2275);
nor U2336 (N_2336,N_2241,N_2240);
nand U2337 (N_2337,N_2229,N_2240);
or U2338 (N_2338,N_2253,N_2251);
xor U2339 (N_2339,N_2261,N_2230);
xnor U2340 (N_2340,N_2306,N_2317);
or U2341 (N_2341,N_2289,N_2319);
nand U2342 (N_2342,N_2298,N_2335);
nor U2343 (N_2343,N_2281,N_2292);
nand U2344 (N_2344,N_2291,N_2325);
xnor U2345 (N_2345,N_2309,N_2300);
xnor U2346 (N_2346,N_2301,N_2307);
xnor U2347 (N_2347,N_2280,N_2312);
nor U2348 (N_2348,N_2324,N_2336);
nor U2349 (N_2349,N_2296,N_2327);
and U2350 (N_2350,N_2305,N_2293);
nor U2351 (N_2351,N_2334,N_2333);
xnor U2352 (N_2352,N_2304,N_2332);
or U2353 (N_2353,N_2338,N_2299);
and U2354 (N_2354,N_2286,N_2284);
or U2355 (N_2355,N_2294,N_2339);
xor U2356 (N_2356,N_2283,N_2320);
and U2357 (N_2357,N_2295,N_2314);
and U2358 (N_2358,N_2322,N_2331);
or U2359 (N_2359,N_2287,N_2318);
nand U2360 (N_2360,N_2311,N_2315);
and U2361 (N_2361,N_2302,N_2313);
or U2362 (N_2362,N_2323,N_2282);
nand U2363 (N_2363,N_2308,N_2288);
xnor U2364 (N_2364,N_2285,N_2297);
or U2365 (N_2365,N_2303,N_2337);
xor U2366 (N_2366,N_2329,N_2316);
xor U2367 (N_2367,N_2328,N_2310);
nand U2368 (N_2368,N_2330,N_2321);
nand U2369 (N_2369,N_2326,N_2290);
xor U2370 (N_2370,N_2335,N_2280);
and U2371 (N_2371,N_2281,N_2296);
and U2372 (N_2372,N_2285,N_2293);
or U2373 (N_2373,N_2336,N_2298);
nand U2374 (N_2374,N_2316,N_2292);
nand U2375 (N_2375,N_2327,N_2332);
nor U2376 (N_2376,N_2316,N_2287);
nand U2377 (N_2377,N_2314,N_2318);
xor U2378 (N_2378,N_2306,N_2339);
or U2379 (N_2379,N_2281,N_2319);
nor U2380 (N_2380,N_2289,N_2309);
and U2381 (N_2381,N_2311,N_2295);
and U2382 (N_2382,N_2286,N_2334);
and U2383 (N_2383,N_2304,N_2318);
nand U2384 (N_2384,N_2301,N_2318);
and U2385 (N_2385,N_2327,N_2311);
nor U2386 (N_2386,N_2293,N_2310);
nor U2387 (N_2387,N_2336,N_2329);
nor U2388 (N_2388,N_2289,N_2328);
or U2389 (N_2389,N_2320,N_2304);
xor U2390 (N_2390,N_2311,N_2302);
and U2391 (N_2391,N_2321,N_2339);
nor U2392 (N_2392,N_2334,N_2329);
nor U2393 (N_2393,N_2315,N_2297);
and U2394 (N_2394,N_2305,N_2283);
xnor U2395 (N_2395,N_2337,N_2290);
or U2396 (N_2396,N_2294,N_2322);
xor U2397 (N_2397,N_2321,N_2317);
nor U2398 (N_2398,N_2287,N_2292);
and U2399 (N_2399,N_2333,N_2330);
nor U2400 (N_2400,N_2375,N_2369);
and U2401 (N_2401,N_2342,N_2374);
nor U2402 (N_2402,N_2378,N_2357);
or U2403 (N_2403,N_2395,N_2388);
nand U2404 (N_2404,N_2345,N_2348);
and U2405 (N_2405,N_2382,N_2372);
xor U2406 (N_2406,N_2352,N_2367);
nor U2407 (N_2407,N_2384,N_2380);
xor U2408 (N_2408,N_2362,N_2381);
nand U2409 (N_2409,N_2398,N_2359);
and U2410 (N_2410,N_2394,N_2373);
and U2411 (N_2411,N_2344,N_2349);
xnor U2412 (N_2412,N_2354,N_2361);
xor U2413 (N_2413,N_2366,N_2389);
or U2414 (N_2414,N_2387,N_2386);
or U2415 (N_2415,N_2368,N_2393);
nor U2416 (N_2416,N_2397,N_2396);
xor U2417 (N_2417,N_2390,N_2341);
or U2418 (N_2418,N_2346,N_2392);
nand U2419 (N_2419,N_2363,N_2350);
or U2420 (N_2420,N_2379,N_2351);
nor U2421 (N_2421,N_2360,N_2376);
xnor U2422 (N_2422,N_2356,N_2355);
nand U2423 (N_2423,N_2347,N_2340);
nand U2424 (N_2424,N_2365,N_2358);
nand U2425 (N_2425,N_2371,N_2377);
or U2426 (N_2426,N_2383,N_2385);
nand U2427 (N_2427,N_2370,N_2399);
xnor U2428 (N_2428,N_2391,N_2343);
or U2429 (N_2429,N_2353,N_2364);
and U2430 (N_2430,N_2360,N_2354);
nand U2431 (N_2431,N_2397,N_2353);
xnor U2432 (N_2432,N_2383,N_2387);
nor U2433 (N_2433,N_2349,N_2382);
nor U2434 (N_2434,N_2368,N_2364);
nand U2435 (N_2435,N_2375,N_2362);
xnor U2436 (N_2436,N_2381,N_2368);
nand U2437 (N_2437,N_2368,N_2360);
xor U2438 (N_2438,N_2393,N_2341);
nand U2439 (N_2439,N_2358,N_2340);
xor U2440 (N_2440,N_2359,N_2389);
nor U2441 (N_2441,N_2386,N_2344);
and U2442 (N_2442,N_2358,N_2359);
nand U2443 (N_2443,N_2387,N_2385);
and U2444 (N_2444,N_2346,N_2396);
nor U2445 (N_2445,N_2396,N_2367);
xor U2446 (N_2446,N_2348,N_2366);
or U2447 (N_2447,N_2351,N_2397);
nand U2448 (N_2448,N_2371,N_2375);
nand U2449 (N_2449,N_2370,N_2376);
xor U2450 (N_2450,N_2342,N_2385);
nand U2451 (N_2451,N_2374,N_2389);
and U2452 (N_2452,N_2379,N_2372);
nor U2453 (N_2453,N_2374,N_2380);
nand U2454 (N_2454,N_2389,N_2355);
and U2455 (N_2455,N_2367,N_2348);
nor U2456 (N_2456,N_2352,N_2373);
nor U2457 (N_2457,N_2395,N_2357);
and U2458 (N_2458,N_2383,N_2340);
nor U2459 (N_2459,N_2390,N_2384);
xor U2460 (N_2460,N_2452,N_2417);
nor U2461 (N_2461,N_2423,N_2409);
nand U2462 (N_2462,N_2432,N_2415);
nand U2463 (N_2463,N_2431,N_2442);
and U2464 (N_2464,N_2419,N_2439);
xnor U2465 (N_2465,N_2455,N_2433);
nor U2466 (N_2466,N_2443,N_2437);
and U2467 (N_2467,N_2427,N_2425);
xnor U2468 (N_2468,N_2453,N_2429);
nor U2469 (N_2469,N_2420,N_2428);
nor U2470 (N_2470,N_2414,N_2456);
nor U2471 (N_2471,N_2408,N_2448);
and U2472 (N_2472,N_2404,N_2424);
or U2473 (N_2473,N_2418,N_2430);
nand U2474 (N_2474,N_2434,N_2440);
xor U2475 (N_2475,N_2401,N_2438);
and U2476 (N_2476,N_2403,N_2458);
or U2477 (N_2477,N_2405,N_2444);
nor U2478 (N_2478,N_2407,N_2406);
and U2479 (N_2479,N_2451,N_2454);
xor U2480 (N_2480,N_2445,N_2422);
and U2481 (N_2481,N_2410,N_2447);
xor U2482 (N_2482,N_2412,N_2457);
xor U2483 (N_2483,N_2402,N_2450);
or U2484 (N_2484,N_2413,N_2421);
nor U2485 (N_2485,N_2416,N_2426);
and U2486 (N_2486,N_2435,N_2459);
nor U2487 (N_2487,N_2441,N_2449);
and U2488 (N_2488,N_2411,N_2436);
xor U2489 (N_2489,N_2400,N_2446);
and U2490 (N_2490,N_2436,N_2459);
nand U2491 (N_2491,N_2400,N_2437);
and U2492 (N_2492,N_2419,N_2448);
and U2493 (N_2493,N_2408,N_2404);
nor U2494 (N_2494,N_2419,N_2432);
or U2495 (N_2495,N_2438,N_2459);
nand U2496 (N_2496,N_2443,N_2416);
and U2497 (N_2497,N_2450,N_2440);
or U2498 (N_2498,N_2402,N_2424);
nand U2499 (N_2499,N_2438,N_2445);
nor U2500 (N_2500,N_2455,N_2415);
nand U2501 (N_2501,N_2408,N_2424);
nor U2502 (N_2502,N_2443,N_2423);
and U2503 (N_2503,N_2448,N_2452);
or U2504 (N_2504,N_2429,N_2436);
and U2505 (N_2505,N_2400,N_2438);
and U2506 (N_2506,N_2457,N_2433);
xnor U2507 (N_2507,N_2452,N_2434);
nand U2508 (N_2508,N_2459,N_2430);
nand U2509 (N_2509,N_2458,N_2424);
xor U2510 (N_2510,N_2454,N_2421);
xor U2511 (N_2511,N_2435,N_2454);
nor U2512 (N_2512,N_2432,N_2417);
nor U2513 (N_2513,N_2446,N_2451);
nor U2514 (N_2514,N_2403,N_2410);
and U2515 (N_2515,N_2435,N_2443);
xor U2516 (N_2516,N_2449,N_2411);
nor U2517 (N_2517,N_2418,N_2437);
nand U2518 (N_2518,N_2403,N_2454);
nor U2519 (N_2519,N_2423,N_2416);
xor U2520 (N_2520,N_2481,N_2487);
nor U2521 (N_2521,N_2503,N_2489);
or U2522 (N_2522,N_2460,N_2499);
nor U2523 (N_2523,N_2504,N_2501);
and U2524 (N_2524,N_2492,N_2518);
nand U2525 (N_2525,N_2500,N_2463);
or U2526 (N_2526,N_2475,N_2506);
or U2527 (N_2527,N_2511,N_2478);
or U2528 (N_2528,N_2488,N_2494);
or U2529 (N_2529,N_2472,N_2505);
or U2530 (N_2530,N_2467,N_2464);
xnor U2531 (N_2531,N_2490,N_2482);
or U2532 (N_2532,N_2502,N_2476);
nor U2533 (N_2533,N_2509,N_2468);
and U2534 (N_2534,N_2495,N_2477);
nand U2535 (N_2535,N_2462,N_2479);
nand U2536 (N_2536,N_2516,N_2517);
xnor U2537 (N_2537,N_2515,N_2465);
nor U2538 (N_2538,N_2469,N_2514);
nor U2539 (N_2539,N_2496,N_2485);
and U2540 (N_2540,N_2493,N_2466);
xnor U2541 (N_2541,N_2480,N_2510);
nor U2542 (N_2542,N_2507,N_2512);
and U2543 (N_2543,N_2484,N_2491);
or U2544 (N_2544,N_2513,N_2497);
xnor U2545 (N_2545,N_2470,N_2483);
xor U2546 (N_2546,N_2508,N_2474);
xnor U2547 (N_2547,N_2486,N_2461);
xnor U2548 (N_2548,N_2498,N_2471);
nor U2549 (N_2549,N_2473,N_2519);
or U2550 (N_2550,N_2483,N_2479);
xor U2551 (N_2551,N_2480,N_2512);
and U2552 (N_2552,N_2470,N_2467);
or U2553 (N_2553,N_2502,N_2481);
xor U2554 (N_2554,N_2512,N_2485);
nor U2555 (N_2555,N_2490,N_2489);
and U2556 (N_2556,N_2471,N_2499);
xnor U2557 (N_2557,N_2461,N_2499);
or U2558 (N_2558,N_2497,N_2460);
xor U2559 (N_2559,N_2469,N_2472);
nor U2560 (N_2560,N_2474,N_2515);
nor U2561 (N_2561,N_2478,N_2481);
nor U2562 (N_2562,N_2496,N_2460);
or U2563 (N_2563,N_2501,N_2486);
nor U2564 (N_2564,N_2507,N_2486);
nor U2565 (N_2565,N_2475,N_2481);
xnor U2566 (N_2566,N_2519,N_2513);
and U2567 (N_2567,N_2465,N_2484);
xnor U2568 (N_2568,N_2503,N_2465);
nor U2569 (N_2569,N_2473,N_2518);
xnor U2570 (N_2570,N_2506,N_2483);
nand U2571 (N_2571,N_2499,N_2490);
nand U2572 (N_2572,N_2502,N_2485);
xnor U2573 (N_2573,N_2471,N_2491);
xnor U2574 (N_2574,N_2462,N_2472);
xor U2575 (N_2575,N_2494,N_2475);
nand U2576 (N_2576,N_2486,N_2464);
nand U2577 (N_2577,N_2465,N_2506);
xor U2578 (N_2578,N_2517,N_2488);
and U2579 (N_2579,N_2480,N_2496);
and U2580 (N_2580,N_2555,N_2574);
and U2581 (N_2581,N_2554,N_2563);
nand U2582 (N_2582,N_2567,N_2556);
or U2583 (N_2583,N_2541,N_2552);
xnor U2584 (N_2584,N_2551,N_2538);
and U2585 (N_2585,N_2525,N_2537);
xor U2586 (N_2586,N_2570,N_2557);
xor U2587 (N_2587,N_2546,N_2529);
xor U2588 (N_2588,N_2530,N_2526);
and U2589 (N_2589,N_2549,N_2568);
and U2590 (N_2590,N_2561,N_2531);
or U2591 (N_2591,N_2560,N_2575);
xor U2592 (N_2592,N_2532,N_2523);
or U2593 (N_2593,N_2573,N_2533);
and U2594 (N_2594,N_2576,N_2565);
nand U2595 (N_2595,N_2524,N_2564);
or U2596 (N_2596,N_2572,N_2539);
or U2597 (N_2597,N_2545,N_2528);
and U2598 (N_2598,N_2569,N_2540);
nor U2599 (N_2599,N_2543,N_2547);
nor U2600 (N_2600,N_2566,N_2577);
nand U2601 (N_2601,N_2521,N_2544);
or U2602 (N_2602,N_2571,N_2578);
nand U2603 (N_2603,N_2522,N_2562);
and U2604 (N_2604,N_2527,N_2536);
nand U2605 (N_2605,N_2550,N_2558);
nand U2606 (N_2606,N_2579,N_2553);
xnor U2607 (N_2607,N_2542,N_2520);
xor U2608 (N_2608,N_2559,N_2535);
nor U2609 (N_2609,N_2534,N_2548);
nor U2610 (N_2610,N_2521,N_2549);
or U2611 (N_2611,N_2538,N_2539);
xnor U2612 (N_2612,N_2528,N_2541);
or U2613 (N_2613,N_2568,N_2551);
and U2614 (N_2614,N_2520,N_2563);
nand U2615 (N_2615,N_2567,N_2558);
or U2616 (N_2616,N_2522,N_2572);
or U2617 (N_2617,N_2553,N_2563);
and U2618 (N_2618,N_2530,N_2520);
nand U2619 (N_2619,N_2578,N_2562);
nor U2620 (N_2620,N_2557,N_2572);
and U2621 (N_2621,N_2529,N_2561);
nor U2622 (N_2622,N_2547,N_2565);
and U2623 (N_2623,N_2529,N_2528);
nor U2624 (N_2624,N_2533,N_2541);
xnor U2625 (N_2625,N_2559,N_2533);
and U2626 (N_2626,N_2544,N_2522);
and U2627 (N_2627,N_2522,N_2523);
or U2628 (N_2628,N_2523,N_2550);
nand U2629 (N_2629,N_2526,N_2557);
nor U2630 (N_2630,N_2555,N_2575);
xnor U2631 (N_2631,N_2564,N_2541);
xnor U2632 (N_2632,N_2546,N_2578);
xor U2633 (N_2633,N_2560,N_2569);
nor U2634 (N_2634,N_2555,N_2551);
or U2635 (N_2635,N_2550,N_2534);
xnor U2636 (N_2636,N_2538,N_2530);
or U2637 (N_2637,N_2572,N_2551);
xnor U2638 (N_2638,N_2522,N_2545);
nor U2639 (N_2639,N_2556,N_2546);
xnor U2640 (N_2640,N_2625,N_2635);
nor U2641 (N_2641,N_2593,N_2607);
nor U2642 (N_2642,N_2618,N_2613);
nor U2643 (N_2643,N_2619,N_2622);
or U2644 (N_2644,N_2616,N_2621);
or U2645 (N_2645,N_2606,N_2636);
nor U2646 (N_2646,N_2582,N_2605);
or U2647 (N_2647,N_2585,N_2612);
and U2648 (N_2648,N_2608,N_2629);
nor U2649 (N_2649,N_2589,N_2592);
nor U2650 (N_2650,N_2638,N_2603);
and U2651 (N_2651,N_2610,N_2586);
or U2652 (N_2652,N_2590,N_2623);
nand U2653 (N_2653,N_2637,N_2598);
nor U2654 (N_2654,N_2630,N_2628);
nor U2655 (N_2655,N_2626,N_2601);
or U2656 (N_2656,N_2587,N_2611);
or U2657 (N_2657,N_2615,N_2588);
nor U2658 (N_2658,N_2627,N_2634);
nand U2659 (N_2659,N_2633,N_2595);
or U2660 (N_2660,N_2583,N_2617);
or U2661 (N_2661,N_2609,N_2599);
or U2662 (N_2662,N_2584,N_2614);
nand U2663 (N_2663,N_2602,N_2620);
or U2664 (N_2664,N_2639,N_2594);
and U2665 (N_2665,N_2600,N_2581);
nor U2666 (N_2666,N_2624,N_2597);
xnor U2667 (N_2667,N_2580,N_2631);
nand U2668 (N_2668,N_2604,N_2632);
or U2669 (N_2669,N_2591,N_2596);
nand U2670 (N_2670,N_2616,N_2581);
or U2671 (N_2671,N_2600,N_2634);
or U2672 (N_2672,N_2628,N_2626);
nor U2673 (N_2673,N_2639,N_2614);
nand U2674 (N_2674,N_2601,N_2597);
or U2675 (N_2675,N_2584,N_2600);
or U2676 (N_2676,N_2591,N_2624);
and U2677 (N_2677,N_2616,N_2627);
nand U2678 (N_2678,N_2637,N_2601);
or U2679 (N_2679,N_2605,N_2634);
nor U2680 (N_2680,N_2601,N_2636);
nand U2681 (N_2681,N_2591,N_2627);
and U2682 (N_2682,N_2607,N_2602);
xnor U2683 (N_2683,N_2633,N_2611);
nand U2684 (N_2684,N_2594,N_2590);
nor U2685 (N_2685,N_2626,N_2618);
and U2686 (N_2686,N_2584,N_2634);
nor U2687 (N_2687,N_2589,N_2619);
nor U2688 (N_2688,N_2584,N_2629);
and U2689 (N_2689,N_2587,N_2634);
nand U2690 (N_2690,N_2622,N_2606);
or U2691 (N_2691,N_2598,N_2600);
nand U2692 (N_2692,N_2625,N_2618);
or U2693 (N_2693,N_2611,N_2584);
xnor U2694 (N_2694,N_2593,N_2621);
and U2695 (N_2695,N_2635,N_2580);
xor U2696 (N_2696,N_2611,N_2608);
xnor U2697 (N_2697,N_2630,N_2613);
nand U2698 (N_2698,N_2628,N_2599);
or U2699 (N_2699,N_2600,N_2621);
xor U2700 (N_2700,N_2682,N_2690);
nor U2701 (N_2701,N_2640,N_2689);
or U2702 (N_2702,N_2693,N_2654);
xnor U2703 (N_2703,N_2666,N_2667);
xnor U2704 (N_2704,N_2649,N_2680);
and U2705 (N_2705,N_2650,N_2675);
or U2706 (N_2706,N_2678,N_2674);
nor U2707 (N_2707,N_2657,N_2672);
nor U2708 (N_2708,N_2668,N_2695);
or U2709 (N_2709,N_2683,N_2648);
nand U2710 (N_2710,N_2653,N_2681);
nor U2711 (N_2711,N_2660,N_2645);
nor U2712 (N_2712,N_2685,N_2641);
nand U2713 (N_2713,N_2677,N_2670);
and U2714 (N_2714,N_2652,N_2662);
or U2715 (N_2715,N_2664,N_2673);
and U2716 (N_2716,N_2679,N_2698);
xnor U2717 (N_2717,N_2643,N_2642);
or U2718 (N_2718,N_2697,N_2658);
nand U2719 (N_2719,N_2686,N_2684);
xor U2720 (N_2720,N_2687,N_2646);
nor U2721 (N_2721,N_2651,N_2655);
xor U2722 (N_2722,N_2669,N_2688);
nor U2723 (N_2723,N_2661,N_2647);
and U2724 (N_2724,N_2671,N_2694);
or U2725 (N_2725,N_2665,N_2663);
xnor U2726 (N_2726,N_2676,N_2691);
nor U2727 (N_2727,N_2644,N_2656);
and U2728 (N_2728,N_2696,N_2692);
xor U2729 (N_2729,N_2659,N_2699);
and U2730 (N_2730,N_2695,N_2662);
or U2731 (N_2731,N_2673,N_2670);
or U2732 (N_2732,N_2671,N_2679);
nand U2733 (N_2733,N_2645,N_2656);
or U2734 (N_2734,N_2654,N_2699);
and U2735 (N_2735,N_2664,N_2658);
or U2736 (N_2736,N_2655,N_2695);
or U2737 (N_2737,N_2676,N_2695);
nand U2738 (N_2738,N_2646,N_2692);
and U2739 (N_2739,N_2647,N_2687);
nor U2740 (N_2740,N_2666,N_2694);
nand U2741 (N_2741,N_2696,N_2682);
xor U2742 (N_2742,N_2685,N_2668);
and U2743 (N_2743,N_2654,N_2640);
nor U2744 (N_2744,N_2674,N_2677);
nand U2745 (N_2745,N_2691,N_2683);
or U2746 (N_2746,N_2661,N_2676);
xnor U2747 (N_2747,N_2650,N_2684);
and U2748 (N_2748,N_2677,N_2697);
and U2749 (N_2749,N_2667,N_2674);
and U2750 (N_2750,N_2653,N_2658);
xnor U2751 (N_2751,N_2658,N_2679);
xor U2752 (N_2752,N_2699,N_2644);
xor U2753 (N_2753,N_2643,N_2660);
nand U2754 (N_2754,N_2692,N_2651);
and U2755 (N_2755,N_2656,N_2670);
nand U2756 (N_2756,N_2693,N_2649);
nor U2757 (N_2757,N_2684,N_2661);
nor U2758 (N_2758,N_2652,N_2647);
xnor U2759 (N_2759,N_2672,N_2658);
xor U2760 (N_2760,N_2717,N_2743);
xor U2761 (N_2761,N_2708,N_2703);
nand U2762 (N_2762,N_2753,N_2722);
nor U2763 (N_2763,N_2710,N_2741);
nor U2764 (N_2764,N_2725,N_2745);
or U2765 (N_2765,N_2714,N_2726);
nor U2766 (N_2766,N_2715,N_2759);
nand U2767 (N_2767,N_2723,N_2718);
xnor U2768 (N_2768,N_2749,N_2727);
nand U2769 (N_2769,N_2729,N_2734);
and U2770 (N_2770,N_2709,N_2756);
nand U2771 (N_2771,N_2731,N_2733);
nor U2772 (N_2772,N_2739,N_2704);
nor U2773 (N_2773,N_2735,N_2721);
xor U2774 (N_2774,N_2732,N_2736);
xnor U2775 (N_2775,N_2728,N_2711);
nor U2776 (N_2776,N_2757,N_2747);
xor U2777 (N_2777,N_2740,N_2755);
or U2778 (N_2778,N_2720,N_2716);
and U2779 (N_2779,N_2744,N_2752);
xor U2780 (N_2780,N_2713,N_2705);
and U2781 (N_2781,N_2738,N_2700);
xor U2782 (N_2782,N_2712,N_2742);
and U2783 (N_2783,N_2754,N_2751);
xnor U2784 (N_2784,N_2750,N_2758);
nor U2785 (N_2785,N_2748,N_2746);
xor U2786 (N_2786,N_2702,N_2706);
xor U2787 (N_2787,N_2701,N_2724);
nor U2788 (N_2788,N_2737,N_2730);
xor U2789 (N_2789,N_2707,N_2719);
nor U2790 (N_2790,N_2707,N_2703);
nor U2791 (N_2791,N_2742,N_2702);
nand U2792 (N_2792,N_2735,N_2700);
nor U2793 (N_2793,N_2749,N_2750);
and U2794 (N_2794,N_2730,N_2736);
nor U2795 (N_2795,N_2722,N_2727);
or U2796 (N_2796,N_2734,N_2707);
xor U2797 (N_2797,N_2739,N_2751);
xor U2798 (N_2798,N_2755,N_2730);
or U2799 (N_2799,N_2721,N_2755);
nand U2800 (N_2800,N_2723,N_2730);
and U2801 (N_2801,N_2737,N_2704);
xor U2802 (N_2802,N_2720,N_2722);
or U2803 (N_2803,N_2723,N_2733);
and U2804 (N_2804,N_2741,N_2700);
nor U2805 (N_2805,N_2732,N_2724);
and U2806 (N_2806,N_2713,N_2744);
nand U2807 (N_2807,N_2711,N_2752);
nand U2808 (N_2808,N_2729,N_2717);
nor U2809 (N_2809,N_2730,N_2745);
nand U2810 (N_2810,N_2725,N_2712);
nand U2811 (N_2811,N_2716,N_2715);
nor U2812 (N_2812,N_2729,N_2711);
xnor U2813 (N_2813,N_2725,N_2719);
and U2814 (N_2814,N_2741,N_2728);
xor U2815 (N_2815,N_2707,N_2752);
nand U2816 (N_2816,N_2741,N_2704);
xnor U2817 (N_2817,N_2759,N_2702);
or U2818 (N_2818,N_2701,N_2705);
and U2819 (N_2819,N_2747,N_2745);
or U2820 (N_2820,N_2763,N_2780);
xor U2821 (N_2821,N_2797,N_2810);
nand U2822 (N_2822,N_2776,N_2812);
nor U2823 (N_2823,N_2789,N_2796);
and U2824 (N_2824,N_2761,N_2802);
xnor U2825 (N_2825,N_2806,N_2795);
nor U2826 (N_2826,N_2764,N_2794);
nand U2827 (N_2827,N_2791,N_2816);
nand U2828 (N_2828,N_2813,N_2777);
and U2829 (N_2829,N_2786,N_2790);
and U2830 (N_2830,N_2814,N_2817);
nand U2831 (N_2831,N_2792,N_2793);
and U2832 (N_2832,N_2783,N_2805);
nor U2833 (N_2833,N_2782,N_2807);
nand U2834 (N_2834,N_2775,N_2772);
nand U2835 (N_2835,N_2787,N_2778);
nor U2836 (N_2836,N_2800,N_2760);
nor U2837 (N_2837,N_2799,N_2769);
nor U2838 (N_2838,N_2781,N_2762);
nor U2839 (N_2839,N_2804,N_2808);
nor U2840 (N_2840,N_2785,N_2784);
nand U2841 (N_2841,N_2803,N_2818);
nor U2842 (N_2842,N_2766,N_2819);
nand U2843 (N_2843,N_2788,N_2774);
or U2844 (N_2844,N_2779,N_2801);
xor U2845 (N_2845,N_2773,N_2767);
nand U2846 (N_2846,N_2811,N_2768);
xnor U2847 (N_2847,N_2770,N_2798);
and U2848 (N_2848,N_2815,N_2765);
and U2849 (N_2849,N_2771,N_2809);
and U2850 (N_2850,N_2795,N_2778);
nand U2851 (N_2851,N_2792,N_2767);
nand U2852 (N_2852,N_2772,N_2817);
and U2853 (N_2853,N_2783,N_2786);
and U2854 (N_2854,N_2780,N_2807);
xnor U2855 (N_2855,N_2787,N_2786);
xor U2856 (N_2856,N_2809,N_2811);
nor U2857 (N_2857,N_2773,N_2790);
xor U2858 (N_2858,N_2816,N_2787);
and U2859 (N_2859,N_2797,N_2786);
xor U2860 (N_2860,N_2790,N_2791);
xor U2861 (N_2861,N_2802,N_2773);
nand U2862 (N_2862,N_2774,N_2806);
nor U2863 (N_2863,N_2799,N_2818);
nor U2864 (N_2864,N_2776,N_2775);
xor U2865 (N_2865,N_2776,N_2808);
xor U2866 (N_2866,N_2788,N_2790);
nand U2867 (N_2867,N_2763,N_2790);
nand U2868 (N_2868,N_2781,N_2778);
or U2869 (N_2869,N_2797,N_2762);
xor U2870 (N_2870,N_2789,N_2787);
nor U2871 (N_2871,N_2781,N_2783);
and U2872 (N_2872,N_2777,N_2810);
or U2873 (N_2873,N_2818,N_2815);
xnor U2874 (N_2874,N_2803,N_2816);
or U2875 (N_2875,N_2772,N_2769);
nor U2876 (N_2876,N_2783,N_2772);
and U2877 (N_2877,N_2775,N_2817);
nor U2878 (N_2878,N_2810,N_2812);
or U2879 (N_2879,N_2818,N_2781);
or U2880 (N_2880,N_2849,N_2858);
nand U2881 (N_2881,N_2853,N_2879);
and U2882 (N_2882,N_2829,N_2837);
and U2883 (N_2883,N_2852,N_2834);
nor U2884 (N_2884,N_2840,N_2836);
and U2885 (N_2885,N_2869,N_2872);
or U2886 (N_2886,N_2859,N_2860);
nand U2887 (N_2887,N_2845,N_2861);
xnor U2888 (N_2888,N_2874,N_2848);
or U2889 (N_2889,N_2830,N_2839);
nand U2890 (N_2890,N_2828,N_2846);
and U2891 (N_2891,N_2842,N_2825);
or U2892 (N_2892,N_2867,N_2877);
nor U2893 (N_2893,N_2857,N_2856);
or U2894 (N_2894,N_2843,N_2855);
nor U2895 (N_2895,N_2851,N_2831);
nand U2896 (N_2896,N_2854,N_2863);
and U2897 (N_2897,N_2821,N_2876);
or U2898 (N_2898,N_2875,N_2864);
xor U2899 (N_2899,N_2835,N_2865);
nand U2900 (N_2900,N_2820,N_2847);
or U2901 (N_2901,N_2862,N_2833);
xnor U2902 (N_2902,N_2844,N_2850);
or U2903 (N_2903,N_2873,N_2823);
xor U2904 (N_2904,N_2822,N_2838);
or U2905 (N_2905,N_2841,N_2827);
or U2906 (N_2906,N_2832,N_2870);
nor U2907 (N_2907,N_2871,N_2866);
nand U2908 (N_2908,N_2868,N_2826);
and U2909 (N_2909,N_2824,N_2878);
nand U2910 (N_2910,N_2847,N_2859);
nor U2911 (N_2911,N_2863,N_2862);
nand U2912 (N_2912,N_2867,N_2826);
nand U2913 (N_2913,N_2871,N_2825);
xnor U2914 (N_2914,N_2865,N_2860);
xnor U2915 (N_2915,N_2820,N_2839);
and U2916 (N_2916,N_2821,N_2853);
nand U2917 (N_2917,N_2872,N_2852);
nor U2918 (N_2918,N_2839,N_2821);
or U2919 (N_2919,N_2871,N_2874);
nor U2920 (N_2920,N_2857,N_2863);
nand U2921 (N_2921,N_2858,N_2865);
or U2922 (N_2922,N_2836,N_2860);
and U2923 (N_2923,N_2827,N_2859);
xor U2924 (N_2924,N_2867,N_2848);
xor U2925 (N_2925,N_2867,N_2873);
xnor U2926 (N_2926,N_2820,N_2824);
nor U2927 (N_2927,N_2849,N_2827);
and U2928 (N_2928,N_2846,N_2874);
nand U2929 (N_2929,N_2832,N_2879);
xor U2930 (N_2930,N_2846,N_2840);
xnor U2931 (N_2931,N_2867,N_2828);
nor U2932 (N_2932,N_2823,N_2835);
or U2933 (N_2933,N_2830,N_2861);
or U2934 (N_2934,N_2864,N_2843);
nand U2935 (N_2935,N_2836,N_2854);
and U2936 (N_2936,N_2825,N_2849);
nand U2937 (N_2937,N_2864,N_2832);
nor U2938 (N_2938,N_2833,N_2875);
or U2939 (N_2939,N_2830,N_2865);
xor U2940 (N_2940,N_2897,N_2913);
nor U2941 (N_2941,N_2881,N_2892);
or U2942 (N_2942,N_2929,N_2934);
or U2943 (N_2943,N_2909,N_2904);
nand U2944 (N_2944,N_2917,N_2883);
nor U2945 (N_2945,N_2930,N_2880);
or U2946 (N_2946,N_2926,N_2893);
or U2947 (N_2947,N_2920,N_2912);
xor U2948 (N_2948,N_2895,N_2900);
and U2949 (N_2949,N_2894,N_2924);
and U2950 (N_2950,N_2921,N_2919);
or U2951 (N_2951,N_2884,N_2882);
or U2952 (N_2952,N_2906,N_2918);
xor U2953 (N_2953,N_2907,N_2896);
nand U2954 (N_2954,N_2939,N_2890);
and U2955 (N_2955,N_2936,N_2887);
xnor U2956 (N_2956,N_2885,N_2927);
or U2957 (N_2957,N_2910,N_2928);
nor U2958 (N_2958,N_2925,N_2888);
nor U2959 (N_2959,N_2931,N_2903);
nor U2960 (N_2960,N_2902,N_2901);
and U2961 (N_2961,N_2922,N_2891);
nor U2962 (N_2962,N_2899,N_2905);
and U2963 (N_2963,N_2898,N_2933);
nor U2964 (N_2964,N_2938,N_2935);
nor U2965 (N_2965,N_2889,N_2916);
or U2966 (N_2966,N_2908,N_2911);
nor U2967 (N_2967,N_2915,N_2886);
nand U2968 (N_2968,N_2937,N_2923);
xnor U2969 (N_2969,N_2932,N_2914);
nor U2970 (N_2970,N_2922,N_2896);
or U2971 (N_2971,N_2910,N_2922);
nand U2972 (N_2972,N_2894,N_2884);
nand U2973 (N_2973,N_2884,N_2881);
and U2974 (N_2974,N_2890,N_2912);
and U2975 (N_2975,N_2931,N_2900);
nor U2976 (N_2976,N_2938,N_2916);
xor U2977 (N_2977,N_2890,N_2895);
nand U2978 (N_2978,N_2895,N_2893);
nor U2979 (N_2979,N_2909,N_2918);
nand U2980 (N_2980,N_2917,N_2936);
xnor U2981 (N_2981,N_2933,N_2926);
or U2982 (N_2982,N_2913,N_2881);
or U2983 (N_2983,N_2934,N_2909);
nand U2984 (N_2984,N_2911,N_2930);
nor U2985 (N_2985,N_2921,N_2913);
xnor U2986 (N_2986,N_2907,N_2887);
nor U2987 (N_2987,N_2906,N_2903);
nor U2988 (N_2988,N_2885,N_2898);
nand U2989 (N_2989,N_2932,N_2893);
xor U2990 (N_2990,N_2882,N_2895);
nand U2991 (N_2991,N_2933,N_2922);
nor U2992 (N_2992,N_2909,N_2930);
nor U2993 (N_2993,N_2923,N_2880);
nand U2994 (N_2994,N_2919,N_2892);
nor U2995 (N_2995,N_2890,N_2935);
and U2996 (N_2996,N_2892,N_2922);
nor U2997 (N_2997,N_2915,N_2888);
and U2998 (N_2998,N_2938,N_2922);
nor U2999 (N_2999,N_2913,N_2919);
nand UO_0 (O_0,N_2945,N_2954);
nor UO_1 (O_1,N_2981,N_2980);
and UO_2 (O_2,N_2965,N_2951);
nor UO_3 (O_3,N_2995,N_2959);
xnor UO_4 (O_4,N_2984,N_2993);
nand UO_5 (O_5,N_2991,N_2996);
nand UO_6 (O_6,N_2964,N_2971);
xnor UO_7 (O_7,N_2941,N_2961);
nor UO_8 (O_8,N_2943,N_2983);
nor UO_9 (O_9,N_2947,N_2948);
nor UO_10 (O_10,N_2977,N_2988);
or UO_11 (O_11,N_2953,N_2990);
or UO_12 (O_12,N_2967,N_2969);
nand UO_13 (O_13,N_2952,N_2950);
nand UO_14 (O_14,N_2946,N_2979);
nand UO_15 (O_15,N_2970,N_2968);
nand UO_16 (O_16,N_2999,N_2972);
or UO_17 (O_17,N_2998,N_2997);
nand UO_18 (O_18,N_2962,N_2978);
nand UO_19 (O_19,N_2955,N_2956);
nor UO_20 (O_20,N_2989,N_2974);
or UO_21 (O_21,N_2957,N_2973);
xnor UO_22 (O_22,N_2963,N_2942);
nor UO_23 (O_23,N_2940,N_2975);
nand UO_24 (O_24,N_2986,N_2982);
and UO_25 (O_25,N_2994,N_2985);
xor UO_26 (O_26,N_2958,N_2960);
and UO_27 (O_27,N_2992,N_2987);
or UO_28 (O_28,N_2949,N_2976);
nor UO_29 (O_29,N_2966,N_2944);
and UO_30 (O_30,N_2959,N_2951);
nor UO_31 (O_31,N_2993,N_2949);
nand UO_32 (O_32,N_2940,N_2988);
nor UO_33 (O_33,N_2948,N_2955);
and UO_34 (O_34,N_2940,N_2993);
nor UO_35 (O_35,N_2942,N_2953);
or UO_36 (O_36,N_2954,N_2976);
xnor UO_37 (O_37,N_2997,N_2940);
nand UO_38 (O_38,N_2987,N_2994);
xor UO_39 (O_39,N_2981,N_2972);
nand UO_40 (O_40,N_2993,N_2968);
nor UO_41 (O_41,N_2987,N_2972);
nor UO_42 (O_42,N_2960,N_2995);
or UO_43 (O_43,N_2941,N_2981);
nand UO_44 (O_44,N_2941,N_2989);
and UO_45 (O_45,N_2981,N_2961);
xor UO_46 (O_46,N_2979,N_2994);
or UO_47 (O_47,N_2948,N_2985);
xnor UO_48 (O_48,N_2963,N_2979);
xnor UO_49 (O_49,N_2967,N_2955);
or UO_50 (O_50,N_2990,N_2972);
xor UO_51 (O_51,N_2943,N_2989);
xor UO_52 (O_52,N_2953,N_2960);
nand UO_53 (O_53,N_2966,N_2942);
xnor UO_54 (O_54,N_2962,N_2985);
nand UO_55 (O_55,N_2983,N_2971);
nor UO_56 (O_56,N_2949,N_2983);
and UO_57 (O_57,N_2974,N_2957);
xnor UO_58 (O_58,N_2970,N_2993);
and UO_59 (O_59,N_2989,N_2998);
nand UO_60 (O_60,N_2974,N_2950);
or UO_61 (O_61,N_2945,N_2989);
xnor UO_62 (O_62,N_2968,N_2942);
and UO_63 (O_63,N_2995,N_2941);
nand UO_64 (O_64,N_2995,N_2953);
and UO_65 (O_65,N_2970,N_2965);
nor UO_66 (O_66,N_2982,N_2973);
and UO_67 (O_67,N_2940,N_2972);
nand UO_68 (O_68,N_2979,N_2962);
or UO_69 (O_69,N_2974,N_2946);
nor UO_70 (O_70,N_2951,N_2960);
xnor UO_71 (O_71,N_2993,N_2980);
nand UO_72 (O_72,N_2955,N_2985);
nor UO_73 (O_73,N_2987,N_2940);
or UO_74 (O_74,N_2951,N_2978);
or UO_75 (O_75,N_2941,N_2968);
nand UO_76 (O_76,N_2948,N_2956);
or UO_77 (O_77,N_2943,N_2968);
nand UO_78 (O_78,N_2974,N_2944);
nand UO_79 (O_79,N_2987,N_2999);
xnor UO_80 (O_80,N_2963,N_2967);
or UO_81 (O_81,N_2972,N_2977);
nor UO_82 (O_82,N_2976,N_2992);
nand UO_83 (O_83,N_2984,N_2948);
xnor UO_84 (O_84,N_2990,N_2940);
and UO_85 (O_85,N_2956,N_2966);
xnor UO_86 (O_86,N_2987,N_2978);
and UO_87 (O_87,N_2990,N_2947);
xor UO_88 (O_88,N_2974,N_2975);
nor UO_89 (O_89,N_2962,N_2942);
and UO_90 (O_90,N_2974,N_2960);
and UO_91 (O_91,N_2954,N_2986);
nor UO_92 (O_92,N_2947,N_2949);
nand UO_93 (O_93,N_2981,N_2986);
nor UO_94 (O_94,N_2971,N_2974);
or UO_95 (O_95,N_2953,N_2951);
and UO_96 (O_96,N_2956,N_2987);
xor UO_97 (O_97,N_2988,N_2957);
nor UO_98 (O_98,N_2954,N_2949);
and UO_99 (O_99,N_2952,N_2965);
and UO_100 (O_100,N_2950,N_2993);
and UO_101 (O_101,N_2941,N_2963);
and UO_102 (O_102,N_2948,N_2970);
and UO_103 (O_103,N_2971,N_2945);
nand UO_104 (O_104,N_2943,N_2975);
xor UO_105 (O_105,N_2958,N_2950);
or UO_106 (O_106,N_2949,N_2975);
and UO_107 (O_107,N_2998,N_2976);
and UO_108 (O_108,N_2940,N_2947);
and UO_109 (O_109,N_2952,N_2970);
xor UO_110 (O_110,N_2972,N_2973);
nor UO_111 (O_111,N_2989,N_2973);
or UO_112 (O_112,N_2965,N_2963);
nor UO_113 (O_113,N_2956,N_2965);
nor UO_114 (O_114,N_2982,N_2941);
xor UO_115 (O_115,N_2996,N_2979);
and UO_116 (O_116,N_2949,N_2953);
nand UO_117 (O_117,N_2990,N_2988);
or UO_118 (O_118,N_2989,N_2942);
xor UO_119 (O_119,N_2991,N_2968);
xor UO_120 (O_120,N_2993,N_2990);
xnor UO_121 (O_121,N_2994,N_2981);
nand UO_122 (O_122,N_2979,N_2990);
and UO_123 (O_123,N_2991,N_2967);
nor UO_124 (O_124,N_2943,N_2957);
and UO_125 (O_125,N_2997,N_2945);
or UO_126 (O_126,N_2984,N_2963);
xnor UO_127 (O_127,N_2982,N_2983);
nand UO_128 (O_128,N_2978,N_2964);
xor UO_129 (O_129,N_2957,N_2959);
xnor UO_130 (O_130,N_2986,N_2963);
or UO_131 (O_131,N_2987,N_2970);
or UO_132 (O_132,N_2978,N_2966);
or UO_133 (O_133,N_2980,N_2985);
or UO_134 (O_134,N_2962,N_2995);
nor UO_135 (O_135,N_2958,N_2998);
or UO_136 (O_136,N_2977,N_2954);
or UO_137 (O_137,N_2966,N_2995);
or UO_138 (O_138,N_2956,N_2974);
xnor UO_139 (O_139,N_2951,N_2964);
or UO_140 (O_140,N_2944,N_2962);
nor UO_141 (O_141,N_2950,N_2985);
nand UO_142 (O_142,N_2979,N_2958);
nand UO_143 (O_143,N_2960,N_2942);
or UO_144 (O_144,N_2982,N_2963);
nand UO_145 (O_145,N_2977,N_2941);
or UO_146 (O_146,N_2959,N_2942);
xnor UO_147 (O_147,N_2963,N_2945);
nor UO_148 (O_148,N_2977,N_2966);
or UO_149 (O_149,N_2993,N_2942);
or UO_150 (O_150,N_2949,N_2965);
xnor UO_151 (O_151,N_2972,N_2950);
and UO_152 (O_152,N_2960,N_2967);
nand UO_153 (O_153,N_2960,N_2990);
nor UO_154 (O_154,N_2951,N_2995);
nor UO_155 (O_155,N_2941,N_2964);
xnor UO_156 (O_156,N_2948,N_2943);
xor UO_157 (O_157,N_2976,N_2982);
nor UO_158 (O_158,N_2970,N_2957);
and UO_159 (O_159,N_2951,N_2944);
xnor UO_160 (O_160,N_2964,N_2992);
or UO_161 (O_161,N_2985,N_2987);
nor UO_162 (O_162,N_2960,N_2978);
and UO_163 (O_163,N_2965,N_2953);
or UO_164 (O_164,N_2996,N_2971);
nor UO_165 (O_165,N_2966,N_2952);
and UO_166 (O_166,N_2989,N_2965);
and UO_167 (O_167,N_2987,N_2997);
nor UO_168 (O_168,N_2962,N_2998);
xnor UO_169 (O_169,N_2966,N_2961);
xor UO_170 (O_170,N_2981,N_2969);
nand UO_171 (O_171,N_2968,N_2959);
or UO_172 (O_172,N_2993,N_2987);
nor UO_173 (O_173,N_2996,N_2980);
nand UO_174 (O_174,N_2960,N_2994);
xnor UO_175 (O_175,N_2994,N_2954);
or UO_176 (O_176,N_2987,N_2949);
and UO_177 (O_177,N_2963,N_2962);
or UO_178 (O_178,N_2969,N_2971);
xor UO_179 (O_179,N_2967,N_2964);
and UO_180 (O_180,N_2997,N_2957);
or UO_181 (O_181,N_2948,N_2987);
and UO_182 (O_182,N_2999,N_2941);
or UO_183 (O_183,N_2994,N_2964);
or UO_184 (O_184,N_2967,N_2946);
xnor UO_185 (O_185,N_2965,N_2969);
nand UO_186 (O_186,N_2977,N_2964);
nand UO_187 (O_187,N_2949,N_2972);
or UO_188 (O_188,N_2988,N_2994);
nand UO_189 (O_189,N_2977,N_2945);
or UO_190 (O_190,N_2968,N_2971);
nand UO_191 (O_191,N_2942,N_2970);
xor UO_192 (O_192,N_2986,N_2987);
nor UO_193 (O_193,N_2983,N_2954);
or UO_194 (O_194,N_2991,N_2960);
nand UO_195 (O_195,N_2967,N_2982);
and UO_196 (O_196,N_2983,N_2958);
and UO_197 (O_197,N_2983,N_2996);
and UO_198 (O_198,N_2986,N_2957);
and UO_199 (O_199,N_2948,N_2942);
or UO_200 (O_200,N_2990,N_2989);
nor UO_201 (O_201,N_2980,N_2954);
or UO_202 (O_202,N_2993,N_2961);
and UO_203 (O_203,N_2974,N_2996);
nand UO_204 (O_204,N_2990,N_2974);
and UO_205 (O_205,N_2994,N_2953);
and UO_206 (O_206,N_2975,N_2982);
or UO_207 (O_207,N_2980,N_2942);
nor UO_208 (O_208,N_2943,N_2956);
nand UO_209 (O_209,N_2978,N_2973);
nor UO_210 (O_210,N_2986,N_2964);
nand UO_211 (O_211,N_2943,N_2994);
nor UO_212 (O_212,N_2943,N_2992);
xor UO_213 (O_213,N_2987,N_2969);
nand UO_214 (O_214,N_2962,N_2948);
and UO_215 (O_215,N_2985,N_2986);
nor UO_216 (O_216,N_2948,N_2951);
xor UO_217 (O_217,N_2981,N_2958);
or UO_218 (O_218,N_2974,N_2959);
xor UO_219 (O_219,N_2970,N_2996);
nor UO_220 (O_220,N_2948,N_2957);
xor UO_221 (O_221,N_2998,N_2951);
nor UO_222 (O_222,N_2947,N_2963);
xnor UO_223 (O_223,N_2950,N_2964);
or UO_224 (O_224,N_2976,N_2985);
xor UO_225 (O_225,N_2950,N_2967);
nor UO_226 (O_226,N_2992,N_2986);
and UO_227 (O_227,N_2951,N_2954);
and UO_228 (O_228,N_2970,N_2984);
nand UO_229 (O_229,N_2955,N_2941);
and UO_230 (O_230,N_2971,N_2963);
and UO_231 (O_231,N_2976,N_2964);
nand UO_232 (O_232,N_2986,N_2971);
xor UO_233 (O_233,N_2970,N_2980);
nor UO_234 (O_234,N_2969,N_2945);
nor UO_235 (O_235,N_2952,N_2987);
nor UO_236 (O_236,N_2956,N_2995);
and UO_237 (O_237,N_2964,N_2961);
or UO_238 (O_238,N_2962,N_2996);
xnor UO_239 (O_239,N_2945,N_2965);
xnor UO_240 (O_240,N_2946,N_2952);
or UO_241 (O_241,N_2978,N_2983);
xor UO_242 (O_242,N_2978,N_2981);
nand UO_243 (O_243,N_2951,N_2997);
nand UO_244 (O_244,N_2949,N_2997);
or UO_245 (O_245,N_2996,N_2941);
and UO_246 (O_246,N_2992,N_2982);
and UO_247 (O_247,N_2963,N_2948);
xor UO_248 (O_248,N_2991,N_2985);
or UO_249 (O_249,N_2985,N_2995);
xnor UO_250 (O_250,N_2962,N_2961);
and UO_251 (O_251,N_2967,N_2970);
nor UO_252 (O_252,N_2990,N_2957);
and UO_253 (O_253,N_2956,N_2954);
and UO_254 (O_254,N_2979,N_2972);
or UO_255 (O_255,N_2985,N_2952);
xnor UO_256 (O_256,N_2942,N_2984);
nand UO_257 (O_257,N_2980,N_2998);
nor UO_258 (O_258,N_2989,N_2968);
or UO_259 (O_259,N_2963,N_2957);
or UO_260 (O_260,N_2983,N_2956);
nand UO_261 (O_261,N_2977,N_2967);
nand UO_262 (O_262,N_2991,N_2948);
and UO_263 (O_263,N_2942,N_2971);
and UO_264 (O_264,N_2961,N_2965);
nand UO_265 (O_265,N_2967,N_2942);
or UO_266 (O_266,N_2952,N_2992);
and UO_267 (O_267,N_2972,N_2959);
nor UO_268 (O_268,N_2970,N_2959);
nand UO_269 (O_269,N_2970,N_2979);
or UO_270 (O_270,N_2946,N_2966);
or UO_271 (O_271,N_2983,N_2979);
nand UO_272 (O_272,N_2999,N_2984);
xor UO_273 (O_273,N_2949,N_2970);
or UO_274 (O_274,N_2959,N_2998);
xor UO_275 (O_275,N_2954,N_2974);
or UO_276 (O_276,N_2992,N_2988);
or UO_277 (O_277,N_2945,N_2978);
and UO_278 (O_278,N_2976,N_2944);
or UO_279 (O_279,N_2995,N_2990);
and UO_280 (O_280,N_2951,N_2996);
and UO_281 (O_281,N_2952,N_2963);
nor UO_282 (O_282,N_2953,N_2971);
nor UO_283 (O_283,N_2983,N_2944);
and UO_284 (O_284,N_2951,N_2946);
and UO_285 (O_285,N_2994,N_2941);
or UO_286 (O_286,N_2946,N_2958);
nand UO_287 (O_287,N_2950,N_2966);
nand UO_288 (O_288,N_2989,N_2955);
nand UO_289 (O_289,N_2998,N_2956);
nor UO_290 (O_290,N_2944,N_2986);
or UO_291 (O_291,N_2948,N_2973);
or UO_292 (O_292,N_2978,N_2969);
or UO_293 (O_293,N_2969,N_2947);
nand UO_294 (O_294,N_2944,N_2965);
or UO_295 (O_295,N_2973,N_2969);
and UO_296 (O_296,N_2947,N_2980);
and UO_297 (O_297,N_2941,N_2945);
nand UO_298 (O_298,N_2979,N_2991);
nor UO_299 (O_299,N_2943,N_2947);
or UO_300 (O_300,N_2971,N_2948);
nand UO_301 (O_301,N_2972,N_2945);
nand UO_302 (O_302,N_2995,N_2948);
or UO_303 (O_303,N_2949,N_2973);
nor UO_304 (O_304,N_2997,N_2946);
nand UO_305 (O_305,N_2997,N_2985);
and UO_306 (O_306,N_2964,N_2966);
or UO_307 (O_307,N_2971,N_2967);
and UO_308 (O_308,N_2954,N_2946);
nor UO_309 (O_309,N_2982,N_2947);
or UO_310 (O_310,N_2984,N_2965);
xor UO_311 (O_311,N_2942,N_2987);
xnor UO_312 (O_312,N_2943,N_2964);
xnor UO_313 (O_313,N_2981,N_2997);
xor UO_314 (O_314,N_2979,N_2999);
or UO_315 (O_315,N_2946,N_2996);
or UO_316 (O_316,N_2960,N_2998);
or UO_317 (O_317,N_2956,N_2940);
xnor UO_318 (O_318,N_2999,N_2940);
xor UO_319 (O_319,N_2943,N_2949);
nand UO_320 (O_320,N_2996,N_2964);
nand UO_321 (O_321,N_2976,N_2945);
nand UO_322 (O_322,N_2999,N_2978);
nand UO_323 (O_323,N_2977,N_2989);
nand UO_324 (O_324,N_2985,N_2953);
nand UO_325 (O_325,N_2964,N_2962);
or UO_326 (O_326,N_2952,N_2956);
nor UO_327 (O_327,N_2989,N_2952);
xnor UO_328 (O_328,N_2961,N_2950);
or UO_329 (O_329,N_2998,N_2992);
nor UO_330 (O_330,N_2961,N_2946);
and UO_331 (O_331,N_2959,N_2996);
nand UO_332 (O_332,N_2973,N_2943);
and UO_333 (O_333,N_2968,N_2951);
nand UO_334 (O_334,N_2975,N_2952);
xnor UO_335 (O_335,N_2947,N_2998);
nor UO_336 (O_336,N_2987,N_2953);
nor UO_337 (O_337,N_2953,N_2992);
xor UO_338 (O_338,N_2987,N_2965);
and UO_339 (O_339,N_2976,N_2999);
nor UO_340 (O_340,N_2954,N_2987);
or UO_341 (O_341,N_2971,N_2947);
or UO_342 (O_342,N_2946,N_2972);
nand UO_343 (O_343,N_2940,N_2973);
nor UO_344 (O_344,N_2957,N_2951);
and UO_345 (O_345,N_2998,N_2991);
nand UO_346 (O_346,N_2955,N_2976);
or UO_347 (O_347,N_2974,N_2967);
and UO_348 (O_348,N_2945,N_2966);
nor UO_349 (O_349,N_2983,N_2970);
nor UO_350 (O_350,N_2985,N_2990);
and UO_351 (O_351,N_2945,N_2944);
or UO_352 (O_352,N_2976,N_2979);
and UO_353 (O_353,N_2976,N_2956);
xnor UO_354 (O_354,N_2986,N_2972);
and UO_355 (O_355,N_2952,N_2972);
or UO_356 (O_356,N_2989,N_2972);
or UO_357 (O_357,N_2940,N_2960);
nand UO_358 (O_358,N_2940,N_2985);
or UO_359 (O_359,N_2964,N_2985);
and UO_360 (O_360,N_2992,N_2967);
nor UO_361 (O_361,N_2984,N_2973);
nor UO_362 (O_362,N_2997,N_2991);
and UO_363 (O_363,N_2973,N_2991);
nor UO_364 (O_364,N_2973,N_2950);
nand UO_365 (O_365,N_2989,N_2954);
xor UO_366 (O_366,N_2952,N_2983);
or UO_367 (O_367,N_2982,N_2940);
nand UO_368 (O_368,N_2955,N_2972);
nand UO_369 (O_369,N_2977,N_2983);
and UO_370 (O_370,N_2977,N_2996);
nand UO_371 (O_371,N_2987,N_2966);
nand UO_372 (O_372,N_2978,N_2950);
nand UO_373 (O_373,N_2984,N_2987);
xnor UO_374 (O_374,N_2953,N_2975);
and UO_375 (O_375,N_2999,N_2958);
nor UO_376 (O_376,N_2989,N_2981);
nor UO_377 (O_377,N_2974,N_2948);
or UO_378 (O_378,N_2982,N_2966);
xnor UO_379 (O_379,N_2953,N_2958);
or UO_380 (O_380,N_2943,N_2988);
nand UO_381 (O_381,N_2958,N_2956);
xnor UO_382 (O_382,N_2945,N_2948);
or UO_383 (O_383,N_2979,N_2959);
nor UO_384 (O_384,N_2968,N_2953);
and UO_385 (O_385,N_2993,N_2952);
nor UO_386 (O_386,N_2970,N_2941);
nor UO_387 (O_387,N_2977,N_2946);
xnor UO_388 (O_388,N_2997,N_2992);
and UO_389 (O_389,N_2972,N_2994);
or UO_390 (O_390,N_2942,N_2940);
and UO_391 (O_391,N_2944,N_2950);
nor UO_392 (O_392,N_2944,N_2958);
nand UO_393 (O_393,N_2953,N_2955);
nand UO_394 (O_394,N_2990,N_2954);
and UO_395 (O_395,N_2952,N_2960);
and UO_396 (O_396,N_2982,N_2945);
xnor UO_397 (O_397,N_2995,N_2961);
or UO_398 (O_398,N_2968,N_2963);
nand UO_399 (O_399,N_2988,N_2965);
nand UO_400 (O_400,N_2971,N_2955);
nor UO_401 (O_401,N_2947,N_2999);
and UO_402 (O_402,N_2986,N_2991);
xnor UO_403 (O_403,N_2965,N_2964);
nand UO_404 (O_404,N_2988,N_2985);
and UO_405 (O_405,N_2996,N_2950);
nor UO_406 (O_406,N_2943,N_2972);
or UO_407 (O_407,N_2962,N_2991);
nand UO_408 (O_408,N_2959,N_2975);
nand UO_409 (O_409,N_2947,N_2944);
xor UO_410 (O_410,N_2956,N_2942);
or UO_411 (O_411,N_2953,N_2976);
xnor UO_412 (O_412,N_2994,N_2998);
and UO_413 (O_413,N_2990,N_2968);
xor UO_414 (O_414,N_2961,N_2942);
xnor UO_415 (O_415,N_2947,N_2953);
nor UO_416 (O_416,N_2967,N_2993);
or UO_417 (O_417,N_2956,N_2991);
xnor UO_418 (O_418,N_2947,N_2962);
nor UO_419 (O_419,N_2943,N_2962);
and UO_420 (O_420,N_2964,N_2970);
or UO_421 (O_421,N_2985,N_2946);
and UO_422 (O_422,N_2970,N_2956);
nor UO_423 (O_423,N_2955,N_2957);
nor UO_424 (O_424,N_2957,N_2962);
nand UO_425 (O_425,N_2945,N_2991);
nand UO_426 (O_426,N_2944,N_2972);
or UO_427 (O_427,N_2952,N_2940);
and UO_428 (O_428,N_2954,N_2965);
nor UO_429 (O_429,N_2990,N_2951);
nor UO_430 (O_430,N_2957,N_2994);
xnor UO_431 (O_431,N_2996,N_2997);
nand UO_432 (O_432,N_2950,N_2943);
xor UO_433 (O_433,N_2948,N_2952);
nand UO_434 (O_434,N_2989,N_2975);
nand UO_435 (O_435,N_2958,N_2988);
xnor UO_436 (O_436,N_2941,N_2976);
and UO_437 (O_437,N_2953,N_2999);
nand UO_438 (O_438,N_2974,N_2997);
and UO_439 (O_439,N_2984,N_2940);
xor UO_440 (O_440,N_2979,N_2986);
nand UO_441 (O_441,N_2991,N_2961);
nor UO_442 (O_442,N_2961,N_2978);
xor UO_443 (O_443,N_2947,N_2955);
or UO_444 (O_444,N_2943,N_2977);
nand UO_445 (O_445,N_2999,N_2957);
nor UO_446 (O_446,N_2981,N_2991);
or UO_447 (O_447,N_2972,N_2941);
nand UO_448 (O_448,N_2983,N_2980);
or UO_449 (O_449,N_2969,N_2958);
nor UO_450 (O_450,N_2993,N_2953);
xnor UO_451 (O_451,N_2971,N_2950);
nor UO_452 (O_452,N_2962,N_2970);
and UO_453 (O_453,N_2985,N_2958);
xor UO_454 (O_454,N_2997,N_2966);
nand UO_455 (O_455,N_2954,N_2995);
or UO_456 (O_456,N_2988,N_2968);
or UO_457 (O_457,N_2959,N_2940);
xor UO_458 (O_458,N_2946,N_2981);
or UO_459 (O_459,N_2954,N_2944);
xor UO_460 (O_460,N_2958,N_2955);
nand UO_461 (O_461,N_2961,N_2955);
and UO_462 (O_462,N_2984,N_2968);
and UO_463 (O_463,N_2951,N_2947);
nand UO_464 (O_464,N_2942,N_2951);
or UO_465 (O_465,N_2951,N_2963);
nor UO_466 (O_466,N_2989,N_2992);
nand UO_467 (O_467,N_2941,N_2985);
or UO_468 (O_468,N_2973,N_2964);
or UO_469 (O_469,N_2950,N_2979);
nor UO_470 (O_470,N_2960,N_2944);
nor UO_471 (O_471,N_2942,N_2958);
xnor UO_472 (O_472,N_2975,N_2970);
xor UO_473 (O_473,N_2975,N_2972);
or UO_474 (O_474,N_2983,N_2985);
or UO_475 (O_475,N_2958,N_2992);
nor UO_476 (O_476,N_2996,N_2999);
nand UO_477 (O_477,N_2983,N_2946);
xnor UO_478 (O_478,N_2970,N_2995);
and UO_479 (O_479,N_2975,N_2981);
or UO_480 (O_480,N_2989,N_2951);
or UO_481 (O_481,N_2991,N_2990);
or UO_482 (O_482,N_2954,N_2959);
and UO_483 (O_483,N_2980,N_2959);
nor UO_484 (O_484,N_2965,N_2999);
or UO_485 (O_485,N_2955,N_2988);
or UO_486 (O_486,N_2955,N_2979);
nand UO_487 (O_487,N_2984,N_2989);
nor UO_488 (O_488,N_2988,N_2971);
nand UO_489 (O_489,N_2962,N_2958);
or UO_490 (O_490,N_2944,N_2961);
nand UO_491 (O_491,N_2948,N_2941);
nand UO_492 (O_492,N_2976,N_2990);
nor UO_493 (O_493,N_2970,N_2978);
nand UO_494 (O_494,N_2945,N_2992);
nand UO_495 (O_495,N_2951,N_2976);
and UO_496 (O_496,N_2955,N_2940);
or UO_497 (O_497,N_2989,N_2960);
xnor UO_498 (O_498,N_2981,N_2954);
nand UO_499 (O_499,N_2974,N_2963);
endmodule