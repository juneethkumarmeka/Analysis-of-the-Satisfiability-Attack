module basic_500_3000_500_40_levels_1xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_253,In_462);
or U1 (N_1,In_125,In_307);
nor U2 (N_2,In_295,In_335);
or U3 (N_3,In_352,In_189);
or U4 (N_4,In_230,In_313);
or U5 (N_5,In_263,In_221);
nor U6 (N_6,In_225,In_424);
and U7 (N_7,In_116,In_278);
nand U8 (N_8,In_287,In_317);
nor U9 (N_9,In_403,In_249);
and U10 (N_10,In_224,In_162);
nand U11 (N_11,In_23,In_132);
or U12 (N_12,In_367,In_427);
and U13 (N_13,In_419,In_94);
and U14 (N_14,In_393,In_44);
nand U15 (N_15,In_145,In_61);
and U16 (N_16,In_1,In_106);
or U17 (N_17,In_337,In_192);
nor U18 (N_18,In_46,In_179);
nand U19 (N_19,In_330,In_164);
and U20 (N_20,In_444,In_381);
and U21 (N_21,In_89,In_67);
nor U22 (N_22,In_100,In_205);
nand U23 (N_23,In_277,In_37);
or U24 (N_24,In_377,In_396);
or U25 (N_25,In_4,In_341);
and U26 (N_26,In_451,In_402);
xnor U27 (N_27,In_443,In_475);
nor U28 (N_28,In_196,In_312);
or U29 (N_29,In_273,In_487);
nand U30 (N_30,In_104,In_372);
xor U31 (N_31,In_30,In_364);
or U32 (N_32,In_136,In_260);
and U33 (N_33,In_360,In_413);
or U34 (N_34,In_329,In_168);
or U35 (N_35,In_201,In_315);
or U36 (N_36,In_129,In_480);
nor U37 (N_37,In_181,In_430);
nand U38 (N_38,In_442,In_344);
nand U39 (N_39,In_256,In_157);
nor U40 (N_40,In_452,In_121);
nor U41 (N_41,In_169,In_27);
nor U42 (N_42,In_466,In_382);
and U43 (N_43,In_264,In_434);
and U44 (N_44,In_450,In_68);
nor U45 (N_45,In_332,In_423);
nand U46 (N_46,In_325,In_302);
nand U47 (N_47,In_361,In_47);
or U48 (N_48,In_180,In_75);
nor U49 (N_49,In_453,In_175);
nor U50 (N_50,In_216,In_353);
nor U51 (N_51,In_149,In_73);
nor U52 (N_52,In_62,In_463);
or U53 (N_53,In_394,In_316);
or U54 (N_54,In_18,In_446);
and U55 (N_55,In_398,In_178);
and U56 (N_56,In_69,In_187);
and U57 (N_57,In_228,In_31);
nand U58 (N_58,In_214,In_139);
nand U59 (N_59,In_327,In_107);
nor U60 (N_60,In_217,In_248);
nor U61 (N_61,In_343,In_265);
nor U62 (N_62,In_152,In_211);
or U63 (N_63,In_238,In_25);
and U64 (N_64,In_71,In_399);
nand U65 (N_65,In_99,In_90);
nor U66 (N_66,In_355,In_209);
or U67 (N_67,In_400,In_24);
xnor U68 (N_68,In_490,In_252);
and U69 (N_69,In_279,In_338);
xor U70 (N_70,In_479,In_231);
and U71 (N_71,In_28,In_153);
or U72 (N_72,In_191,In_17);
nor U73 (N_73,In_433,In_418);
and U74 (N_74,In_432,In_455);
and U75 (N_75,N_63,N_60);
nand U76 (N_76,In_86,In_274);
nor U77 (N_77,In_469,In_236);
or U78 (N_78,In_227,In_156);
nand U79 (N_79,In_10,In_166);
or U80 (N_80,In_134,N_45);
nor U81 (N_81,In_448,In_291);
nor U82 (N_82,In_392,In_460);
nand U83 (N_83,In_405,In_297);
or U84 (N_84,N_51,In_321);
or U85 (N_85,In_440,In_314);
or U86 (N_86,In_112,In_246);
nor U87 (N_87,In_117,In_207);
nor U88 (N_88,N_70,In_190);
and U89 (N_89,In_150,In_262);
nand U90 (N_90,In_105,In_135);
nor U91 (N_91,In_483,N_4);
and U92 (N_92,In_22,In_366);
xnor U93 (N_93,In_384,N_22);
nor U94 (N_94,In_284,In_375);
nand U95 (N_95,N_1,In_130);
nand U96 (N_96,N_13,N_46);
nor U97 (N_97,In_472,In_354);
nor U98 (N_98,In_223,In_144);
nor U99 (N_99,In_141,N_62);
nand U100 (N_100,N_64,In_138);
or U101 (N_101,In_477,In_486);
nor U102 (N_102,In_102,In_435);
nor U103 (N_103,In_296,In_436);
nor U104 (N_104,N_68,In_220);
and U105 (N_105,N_61,In_328);
or U106 (N_106,In_323,In_78);
nor U107 (N_107,In_456,In_242);
nand U108 (N_108,In_218,In_385);
or U109 (N_109,In_373,In_210);
nand U110 (N_110,In_148,In_76);
and U111 (N_111,N_18,In_8);
and U112 (N_112,In_66,In_203);
or U113 (N_113,In_159,In_63);
nand U114 (N_114,In_15,In_499);
nor U115 (N_115,In_53,In_300);
nor U116 (N_116,In_488,In_70);
and U117 (N_117,N_58,In_49);
and U118 (N_118,N_29,N_9);
nand U119 (N_119,In_208,In_206);
or U120 (N_120,In_142,N_17);
or U121 (N_121,In_176,N_7);
and U122 (N_122,In_240,In_416);
nor U123 (N_123,In_83,In_82);
nor U124 (N_124,In_378,In_408);
and U125 (N_125,In_174,In_350);
nand U126 (N_126,N_2,In_348);
and U127 (N_127,In_155,N_67);
or U128 (N_128,In_151,In_186);
or U129 (N_129,In_26,In_177);
or U130 (N_130,In_411,In_33);
and U131 (N_131,In_124,In_441);
nor U132 (N_132,In_380,In_457);
and U133 (N_133,In_351,N_15);
or U134 (N_134,In_255,In_184);
or U135 (N_135,In_92,In_103);
or U136 (N_136,In_383,N_69);
or U137 (N_137,In_294,In_454);
and U138 (N_138,N_54,In_303);
or U139 (N_139,In_74,In_16);
and U140 (N_140,N_74,In_48);
nor U141 (N_141,N_12,In_266);
nand U142 (N_142,In_133,In_213);
or U143 (N_143,In_261,N_53);
nor U144 (N_144,N_49,In_122);
nand U145 (N_145,In_356,In_172);
and U146 (N_146,In_0,In_369);
and U147 (N_147,In_391,In_14);
nor U148 (N_148,In_11,In_493);
nor U149 (N_149,In_461,In_299);
or U150 (N_150,In_492,In_215);
and U151 (N_151,In_146,N_108);
nor U152 (N_152,N_24,In_346);
nor U153 (N_153,In_199,In_447);
nor U154 (N_154,In_473,In_183);
nand U155 (N_155,N_33,In_345);
or U156 (N_156,In_96,In_478);
nand U157 (N_157,N_145,N_42);
and U158 (N_158,In_270,In_401);
or U159 (N_159,N_119,In_54);
and U160 (N_160,In_165,N_6);
and U161 (N_161,N_36,N_113);
or U162 (N_162,N_144,In_304);
or U163 (N_163,In_267,In_7);
and U164 (N_164,In_21,In_194);
nand U165 (N_165,N_37,In_160);
xnor U166 (N_166,In_29,In_320);
and U167 (N_167,In_42,In_494);
and U168 (N_168,N_129,In_286);
and U169 (N_169,In_147,N_89);
or U170 (N_170,In_458,N_3);
nand U171 (N_171,In_368,In_77);
nand U172 (N_172,N_141,N_52);
and U173 (N_173,N_20,In_484);
or U174 (N_174,In_154,N_39);
nor U175 (N_175,In_195,In_497);
and U176 (N_176,In_386,In_421);
or U177 (N_177,In_95,In_202);
nand U178 (N_178,N_75,In_34);
nor U179 (N_179,N_140,N_10);
nor U180 (N_180,In_91,In_158);
or U181 (N_181,N_104,In_204);
nand U182 (N_182,N_100,In_425);
and U183 (N_183,In_81,In_237);
or U184 (N_184,N_133,N_97);
nand U185 (N_185,N_110,N_143);
and U186 (N_186,In_241,In_359);
nand U187 (N_187,In_171,In_410);
nand U188 (N_188,In_498,N_116);
and U189 (N_189,In_140,In_482);
and U190 (N_190,In_485,N_99);
nor U191 (N_191,In_467,N_86);
nor U192 (N_192,N_130,In_407);
nand U193 (N_193,In_257,N_21);
and U194 (N_194,In_72,In_119);
nor U195 (N_195,N_134,N_30);
and U196 (N_196,N_72,N_28);
nand U197 (N_197,In_13,N_94);
or U198 (N_198,In_310,N_55);
nor U199 (N_199,N_142,In_471);
nor U200 (N_200,N_50,In_51);
nand U201 (N_201,In_362,N_26);
nand U202 (N_202,In_331,In_87);
and U203 (N_203,N_11,In_250);
nor U204 (N_204,In_491,In_374);
and U205 (N_205,N_56,In_397);
nand U206 (N_206,In_288,In_259);
or U207 (N_207,N_136,N_31);
nor U208 (N_208,N_59,In_193);
nand U209 (N_209,In_420,N_73);
nor U210 (N_210,In_113,In_376);
nor U211 (N_211,N_93,In_2);
and U212 (N_212,In_336,In_59);
nor U213 (N_213,In_131,In_41);
nand U214 (N_214,In_12,In_342);
nor U215 (N_215,In_85,In_20);
and U216 (N_216,In_232,In_108);
and U217 (N_217,In_406,In_57);
nand U218 (N_218,In_404,In_289);
nand U219 (N_219,In_426,In_3);
and U220 (N_220,In_318,In_334);
and U221 (N_221,N_40,N_128);
or U222 (N_222,In_93,In_185);
nor U223 (N_223,N_98,N_101);
or U224 (N_224,In_110,In_198);
and U225 (N_225,N_23,In_43);
nand U226 (N_226,In_36,In_229);
and U227 (N_227,In_45,In_79);
or U228 (N_228,In_415,In_167);
or U229 (N_229,N_204,N_8);
or U230 (N_230,In_347,N_121);
and U231 (N_231,In_311,In_39);
nor U232 (N_232,N_183,In_281);
or U233 (N_233,N_210,N_201);
nand U234 (N_234,In_449,N_215);
nor U235 (N_235,N_88,N_195);
nor U236 (N_236,N_81,In_50);
nor U237 (N_237,N_188,N_78);
nand U238 (N_238,N_191,In_388);
nor U239 (N_239,In_137,N_214);
nor U240 (N_240,In_251,In_5);
nand U241 (N_241,N_109,In_437);
nor U242 (N_242,N_162,N_178);
or U243 (N_243,N_43,N_172);
nand U244 (N_244,N_181,N_212);
nand U245 (N_245,In_126,N_157);
and U246 (N_246,In_324,In_65);
nand U247 (N_247,N_165,In_389);
nand U248 (N_248,N_85,N_208);
nor U249 (N_249,N_95,N_77);
and U250 (N_250,N_200,In_19);
nor U251 (N_251,In_275,N_199);
or U252 (N_252,In_243,N_196);
or U253 (N_253,N_198,In_118);
nor U254 (N_254,In_128,N_167);
nor U255 (N_255,In_9,N_146);
nand U256 (N_256,N_115,In_98);
nand U257 (N_257,N_139,In_459);
xnor U258 (N_258,In_88,N_185);
nor U259 (N_259,N_122,In_173);
nand U260 (N_260,N_164,N_80);
nand U261 (N_261,In_244,N_44);
nor U262 (N_262,In_357,In_56);
nand U263 (N_263,N_211,In_308);
xnor U264 (N_264,In_163,In_258);
nor U265 (N_265,In_370,In_84);
nand U266 (N_266,N_174,N_153);
nand U267 (N_267,N_92,In_285);
nand U268 (N_268,In_496,In_219);
nor U269 (N_269,N_124,In_390);
nand U270 (N_270,In_109,In_322);
or U271 (N_271,N_206,N_163);
nand U272 (N_272,N_155,In_111);
nand U273 (N_273,N_125,In_200);
nand U274 (N_274,In_188,In_280);
nor U275 (N_275,In_292,N_90);
nand U276 (N_276,In_115,N_170);
nor U277 (N_277,N_103,N_117);
nand U278 (N_278,N_176,N_168);
or U279 (N_279,In_143,In_422);
and U280 (N_280,N_106,In_120);
nor U281 (N_281,N_179,In_114);
or U282 (N_282,In_254,N_216);
nand U283 (N_283,N_151,In_55);
nor U284 (N_284,In_101,In_97);
nor U285 (N_285,N_41,N_84);
or U286 (N_286,In_481,In_306);
or U287 (N_287,N_34,In_245);
or U288 (N_288,In_429,N_156);
nand U289 (N_289,N_83,In_333);
and U290 (N_290,N_57,In_414);
nand U291 (N_291,N_71,N_138);
and U292 (N_292,N_65,In_170);
nand U293 (N_293,In_271,In_64);
nor U294 (N_294,N_25,In_269);
nor U295 (N_295,N_147,N_105);
nor U296 (N_296,N_5,N_220);
and U297 (N_297,In_395,N_14);
nor U298 (N_298,In_417,N_107);
and U299 (N_299,In_305,N_193);
or U300 (N_300,N_47,N_272);
nor U301 (N_301,In_309,N_262);
nor U302 (N_302,N_274,N_263);
nor U303 (N_303,N_294,In_438);
and U304 (N_304,In_339,In_489);
and U305 (N_305,N_158,N_260);
and U306 (N_306,N_0,N_152);
nand U307 (N_307,N_223,N_82);
nand U308 (N_308,In_349,N_186);
nand U309 (N_309,In_283,In_439);
or U310 (N_310,N_226,N_102);
nor U311 (N_311,In_465,N_160);
nor U312 (N_312,N_269,In_412);
nand U313 (N_313,N_232,In_363);
nand U314 (N_314,In_326,N_286);
nor U315 (N_315,N_241,N_150);
nand U316 (N_316,N_218,N_173);
nor U317 (N_317,N_171,N_19);
nand U318 (N_318,N_190,In_282);
or U319 (N_319,N_253,N_114);
and U320 (N_320,N_166,N_229);
nor U321 (N_321,N_295,In_276);
or U322 (N_322,In_197,N_261);
and U323 (N_323,N_35,N_205);
nor U324 (N_324,In_365,In_226);
or U325 (N_325,N_227,N_213);
and U326 (N_326,N_221,In_340);
and U327 (N_327,In_233,N_268);
and U328 (N_328,N_264,N_248);
nand U329 (N_329,N_266,N_280);
nor U330 (N_330,N_127,In_6);
nor U331 (N_331,N_265,N_284);
nand U332 (N_332,N_203,In_298);
nor U333 (N_333,In_379,In_58);
nand U334 (N_334,N_255,N_252);
nand U335 (N_335,N_240,N_184);
nor U336 (N_336,In_319,In_464);
and U337 (N_337,N_267,N_291);
nand U338 (N_338,In_268,In_182);
and U339 (N_339,N_123,N_66);
or U340 (N_340,N_251,N_273);
nand U341 (N_341,In_239,N_161);
or U342 (N_342,N_250,N_243);
nor U343 (N_343,In_123,In_431);
or U344 (N_344,N_159,N_231);
and U345 (N_345,N_32,N_189);
and U346 (N_346,N_96,In_301);
and U347 (N_347,In_387,N_290);
nor U348 (N_348,N_120,N_112);
and U349 (N_349,N_257,N_118);
nor U350 (N_350,In_470,N_299);
nand U351 (N_351,In_127,N_287);
nor U352 (N_352,N_135,N_245);
and U353 (N_353,N_278,N_87);
or U354 (N_354,N_27,N_258);
or U355 (N_355,N_244,N_132);
nor U356 (N_356,N_202,N_239);
or U357 (N_357,N_217,N_234);
or U358 (N_358,In_293,N_224);
nand U359 (N_359,N_259,N_249);
nand U360 (N_360,N_91,N_281);
and U361 (N_361,N_222,N_238);
or U362 (N_362,N_288,N_225);
nand U363 (N_363,In_235,N_16);
or U364 (N_364,N_126,In_468);
nor U365 (N_365,In_38,N_254);
nand U366 (N_366,In_161,N_235);
nand U367 (N_367,N_79,N_219);
nor U368 (N_368,N_169,In_476);
nand U369 (N_369,N_297,In_371);
or U370 (N_370,In_35,N_236);
or U371 (N_371,In_52,N_192);
nor U372 (N_372,N_230,In_212);
and U373 (N_373,In_40,N_131);
nand U374 (N_374,N_149,In_445);
nand U375 (N_375,N_366,N_346);
xor U376 (N_376,N_331,N_357);
nand U377 (N_377,N_362,In_222);
and U378 (N_378,N_354,N_344);
and U379 (N_379,N_374,N_322);
and U380 (N_380,N_154,N_329);
or U381 (N_381,In_247,N_282);
or U382 (N_382,N_342,N_289);
and U383 (N_383,N_356,N_180);
nor U384 (N_384,In_272,In_60);
nand U385 (N_385,N_296,In_428);
and U386 (N_386,In_409,N_323);
and U387 (N_387,N_182,N_349);
nor U388 (N_388,N_148,N_332);
nor U389 (N_389,N_279,N_341);
or U390 (N_390,N_358,N_335);
nor U391 (N_391,N_317,In_358);
and U392 (N_392,N_326,N_275);
or U393 (N_393,N_369,N_312);
and U394 (N_394,N_321,N_247);
and U395 (N_395,N_197,N_270);
nor U396 (N_396,N_175,N_276);
nand U397 (N_397,N_338,In_495);
or U398 (N_398,In_290,N_370);
and U399 (N_399,N_340,N_137);
nand U400 (N_400,N_111,N_360);
nor U401 (N_401,N_38,N_301);
nand U402 (N_402,N_371,N_237);
nand U403 (N_403,N_334,N_307);
nand U404 (N_404,N_177,N_325);
and U405 (N_405,N_228,N_316);
and U406 (N_406,N_365,N_76);
or U407 (N_407,N_302,N_368);
nor U408 (N_408,N_309,N_303);
and U409 (N_409,N_283,N_194);
nand U410 (N_410,N_315,N_318);
or U411 (N_411,N_233,N_350);
nand U412 (N_412,N_348,N_187);
nand U413 (N_413,N_271,N_327);
nand U414 (N_414,N_305,N_352);
nor U415 (N_415,N_339,N_355);
or U416 (N_416,N_364,N_207);
and U417 (N_417,In_80,N_373);
nor U418 (N_418,N_330,N_324);
xnor U419 (N_419,In_234,N_363);
or U420 (N_420,N_246,N_256);
nand U421 (N_421,N_337,N_298);
or U422 (N_422,N_367,N_353);
nand U423 (N_423,N_314,N_361);
and U424 (N_424,N_308,N_351);
and U425 (N_425,N_311,N_242);
and U426 (N_426,N_306,N_359);
or U427 (N_427,N_345,N_209);
nor U428 (N_428,N_347,N_48);
or U429 (N_429,N_292,N_313);
or U430 (N_430,N_285,N_328);
nor U431 (N_431,N_319,N_320);
and U432 (N_432,N_333,In_32);
and U433 (N_433,N_372,N_343);
or U434 (N_434,N_336,In_474);
and U435 (N_435,N_277,N_310);
and U436 (N_436,N_300,N_304);
nand U437 (N_437,N_293,N_303);
nor U438 (N_438,N_330,N_207);
nand U439 (N_439,In_222,N_315);
nand U440 (N_440,N_38,N_276);
and U441 (N_441,N_364,N_237);
and U442 (N_442,N_308,N_368);
nand U443 (N_443,N_364,In_222);
and U444 (N_444,N_175,N_303);
or U445 (N_445,N_233,N_276);
or U446 (N_446,N_148,N_360);
nand U447 (N_447,N_332,N_111);
nand U448 (N_448,N_346,N_332);
nand U449 (N_449,N_338,N_308);
nor U450 (N_450,N_382,N_446);
and U451 (N_451,N_402,N_419);
and U452 (N_452,N_435,N_443);
or U453 (N_453,N_412,N_401);
nand U454 (N_454,N_391,N_448);
nor U455 (N_455,N_432,N_379);
nor U456 (N_456,N_398,N_433);
nand U457 (N_457,N_444,N_425);
nor U458 (N_458,N_427,N_434);
or U459 (N_459,N_424,N_405);
or U460 (N_460,N_409,N_396);
or U461 (N_461,N_406,N_421);
or U462 (N_462,N_385,N_418);
nand U463 (N_463,N_384,N_441);
nand U464 (N_464,N_381,N_389);
or U465 (N_465,N_417,N_439);
nor U466 (N_466,N_442,N_395);
and U467 (N_467,N_377,N_440);
and U468 (N_468,N_420,N_376);
nor U469 (N_469,N_449,N_383);
and U470 (N_470,N_400,N_408);
or U471 (N_471,N_407,N_378);
or U472 (N_472,N_387,N_393);
and U473 (N_473,N_388,N_390);
nor U474 (N_474,N_438,N_414);
and U475 (N_475,N_431,N_422);
or U476 (N_476,N_392,N_380);
nor U477 (N_477,N_411,N_447);
nor U478 (N_478,N_428,N_403);
nand U479 (N_479,N_437,N_415);
nand U480 (N_480,N_386,N_399);
and U481 (N_481,N_375,N_429);
nor U482 (N_482,N_416,N_423);
or U483 (N_483,N_436,N_404);
nor U484 (N_484,N_445,N_430);
and U485 (N_485,N_410,N_426);
nor U486 (N_486,N_397,N_394);
nand U487 (N_487,N_413,N_384);
and U488 (N_488,N_401,N_399);
nand U489 (N_489,N_430,N_437);
nand U490 (N_490,N_427,N_389);
nor U491 (N_491,N_388,N_394);
and U492 (N_492,N_431,N_414);
nand U493 (N_493,N_379,N_376);
nor U494 (N_494,N_399,N_419);
nand U495 (N_495,N_390,N_411);
nand U496 (N_496,N_400,N_380);
or U497 (N_497,N_394,N_448);
nor U498 (N_498,N_425,N_404);
nand U499 (N_499,N_436,N_385);
nand U500 (N_500,N_414,N_386);
nand U501 (N_501,N_412,N_395);
or U502 (N_502,N_423,N_377);
nor U503 (N_503,N_430,N_449);
or U504 (N_504,N_410,N_444);
and U505 (N_505,N_385,N_381);
nor U506 (N_506,N_397,N_434);
nand U507 (N_507,N_404,N_449);
nor U508 (N_508,N_438,N_444);
and U509 (N_509,N_394,N_396);
or U510 (N_510,N_435,N_433);
nand U511 (N_511,N_409,N_399);
nor U512 (N_512,N_429,N_383);
nand U513 (N_513,N_418,N_413);
and U514 (N_514,N_449,N_378);
nor U515 (N_515,N_407,N_383);
nor U516 (N_516,N_380,N_402);
or U517 (N_517,N_382,N_397);
nand U518 (N_518,N_404,N_437);
and U519 (N_519,N_422,N_415);
nand U520 (N_520,N_424,N_385);
nand U521 (N_521,N_425,N_381);
or U522 (N_522,N_380,N_404);
and U523 (N_523,N_422,N_414);
nand U524 (N_524,N_435,N_437);
nor U525 (N_525,N_459,N_478);
nor U526 (N_526,N_472,N_473);
and U527 (N_527,N_513,N_488);
nand U528 (N_528,N_512,N_468);
and U529 (N_529,N_463,N_523);
or U530 (N_530,N_454,N_509);
and U531 (N_531,N_486,N_496);
nor U532 (N_532,N_452,N_505);
or U533 (N_533,N_475,N_487);
or U534 (N_534,N_503,N_469);
and U535 (N_535,N_516,N_471);
nand U536 (N_536,N_502,N_479);
nand U537 (N_537,N_467,N_484);
and U538 (N_538,N_490,N_485);
or U539 (N_539,N_458,N_489);
nor U540 (N_540,N_494,N_457);
nor U541 (N_541,N_517,N_480);
or U542 (N_542,N_451,N_492);
nor U543 (N_543,N_499,N_477);
nor U544 (N_544,N_481,N_460);
nor U545 (N_545,N_455,N_511);
nand U546 (N_546,N_464,N_461);
and U547 (N_547,N_521,N_456);
or U548 (N_548,N_465,N_518);
or U549 (N_549,N_500,N_506);
or U550 (N_550,N_504,N_466);
and U551 (N_551,N_524,N_495);
and U552 (N_552,N_522,N_450);
and U553 (N_553,N_474,N_470);
and U554 (N_554,N_498,N_497);
nand U555 (N_555,N_493,N_482);
or U556 (N_556,N_483,N_510);
or U557 (N_557,N_514,N_519);
nand U558 (N_558,N_491,N_476);
or U559 (N_559,N_501,N_507);
nand U560 (N_560,N_453,N_508);
nand U561 (N_561,N_462,N_515);
nor U562 (N_562,N_520,N_450);
nor U563 (N_563,N_462,N_493);
nor U564 (N_564,N_504,N_470);
and U565 (N_565,N_512,N_465);
and U566 (N_566,N_501,N_455);
or U567 (N_567,N_462,N_484);
nand U568 (N_568,N_476,N_511);
and U569 (N_569,N_501,N_478);
and U570 (N_570,N_495,N_503);
or U571 (N_571,N_506,N_457);
nor U572 (N_572,N_473,N_488);
nand U573 (N_573,N_459,N_471);
and U574 (N_574,N_471,N_482);
nor U575 (N_575,N_495,N_506);
or U576 (N_576,N_480,N_462);
nand U577 (N_577,N_479,N_487);
and U578 (N_578,N_473,N_514);
or U579 (N_579,N_465,N_506);
nor U580 (N_580,N_489,N_496);
nand U581 (N_581,N_501,N_484);
and U582 (N_582,N_457,N_482);
nand U583 (N_583,N_489,N_506);
and U584 (N_584,N_473,N_495);
and U585 (N_585,N_470,N_464);
or U586 (N_586,N_521,N_481);
and U587 (N_587,N_476,N_490);
or U588 (N_588,N_523,N_452);
and U589 (N_589,N_509,N_521);
or U590 (N_590,N_488,N_464);
or U591 (N_591,N_478,N_469);
or U592 (N_592,N_522,N_493);
or U593 (N_593,N_522,N_492);
or U594 (N_594,N_510,N_514);
and U595 (N_595,N_477,N_491);
or U596 (N_596,N_483,N_472);
and U597 (N_597,N_468,N_476);
nand U598 (N_598,N_488,N_511);
nand U599 (N_599,N_511,N_458);
nor U600 (N_600,N_581,N_543);
and U601 (N_601,N_547,N_527);
or U602 (N_602,N_598,N_576);
or U603 (N_603,N_539,N_552);
or U604 (N_604,N_556,N_550);
and U605 (N_605,N_583,N_569);
nor U606 (N_606,N_546,N_596);
nor U607 (N_607,N_595,N_590);
nor U608 (N_608,N_532,N_558);
nor U609 (N_609,N_588,N_597);
nand U610 (N_610,N_529,N_549);
nor U611 (N_611,N_530,N_535);
and U612 (N_612,N_593,N_551);
nor U613 (N_613,N_572,N_567);
nand U614 (N_614,N_542,N_579);
or U615 (N_615,N_553,N_554);
or U616 (N_616,N_575,N_562);
or U617 (N_617,N_570,N_582);
nand U618 (N_618,N_561,N_594);
and U619 (N_619,N_548,N_577);
nor U620 (N_620,N_574,N_585);
or U621 (N_621,N_526,N_568);
nand U622 (N_622,N_587,N_566);
nand U623 (N_623,N_559,N_592);
nand U624 (N_624,N_573,N_537);
and U625 (N_625,N_545,N_555);
nor U626 (N_626,N_589,N_578);
and U627 (N_627,N_528,N_563);
or U628 (N_628,N_565,N_580);
nand U629 (N_629,N_525,N_571);
nor U630 (N_630,N_564,N_540);
or U631 (N_631,N_557,N_584);
or U632 (N_632,N_534,N_536);
or U633 (N_633,N_538,N_591);
nand U634 (N_634,N_531,N_544);
nand U635 (N_635,N_586,N_533);
and U636 (N_636,N_541,N_560);
and U637 (N_637,N_599,N_580);
or U638 (N_638,N_593,N_538);
nor U639 (N_639,N_595,N_561);
or U640 (N_640,N_532,N_557);
and U641 (N_641,N_597,N_532);
nand U642 (N_642,N_579,N_575);
or U643 (N_643,N_542,N_547);
and U644 (N_644,N_595,N_546);
nand U645 (N_645,N_581,N_576);
and U646 (N_646,N_534,N_592);
nor U647 (N_647,N_549,N_528);
nand U648 (N_648,N_571,N_570);
and U649 (N_649,N_552,N_559);
and U650 (N_650,N_532,N_549);
and U651 (N_651,N_528,N_531);
nor U652 (N_652,N_538,N_534);
and U653 (N_653,N_599,N_528);
and U654 (N_654,N_590,N_567);
nand U655 (N_655,N_566,N_573);
or U656 (N_656,N_569,N_590);
or U657 (N_657,N_540,N_526);
and U658 (N_658,N_571,N_599);
nand U659 (N_659,N_565,N_571);
nor U660 (N_660,N_539,N_535);
or U661 (N_661,N_530,N_532);
nand U662 (N_662,N_576,N_531);
nand U663 (N_663,N_550,N_592);
nor U664 (N_664,N_560,N_550);
or U665 (N_665,N_549,N_598);
nor U666 (N_666,N_571,N_543);
nand U667 (N_667,N_571,N_556);
or U668 (N_668,N_585,N_583);
and U669 (N_669,N_592,N_561);
nor U670 (N_670,N_580,N_568);
and U671 (N_671,N_544,N_575);
nor U672 (N_672,N_578,N_593);
or U673 (N_673,N_597,N_578);
and U674 (N_674,N_531,N_573);
and U675 (N_675,N_674,N_620);
or U676 (N_676,N_650,N_673);
and U677 (N_677,N_609,N_636);
xnor U678 (N_678,N_671,N_600);
nand U679 (N_679,N_647,N_667);
nor U680 (N_680,N_639,N_619);
and U681 (N_681,N_652,N_630);
nand U682 (N_682,N_616,N_658);
nor U683 (N_683,N_611,N_628);
nor U684 (N_684,N_670,N_663);
nor U685 (N_685,N_645,N_626);
nor U686 (N_686,N_617,N_627);
or U687 (N_687,N_612,N_655);
nor U688 (N_688,N_633,N_607);
nor U689 (N_689,N_661,N_622);
nor U690 (N_690,N_666,N_629);
and U691 (N_691,N_642,N_672);
or U692 (N_692,N_654,N_624);
nor U693 (N_693,N_644,N_643);
nand U694 (N_694,N_603,N_602);
or U695 (N_695,N_634,N_653);
and U696 (N_696,N_632,N_646);
nand U697 (N_697,N_608,N_657);
nand U698 (N_698,N_637,N_669);
nor U699 (N_699,N_623,N_638);
nor U700 (N_700,N_648,N_651);
nand U701 (N_701,N_631,N_604);
nor U702 (N_702,N_606,N_659);
nor U703 (N_703,N_605,N_613);
or U704 (N_704,N_665,N_641);
or U705 (N_705,N_635,N_649);
and U706 (N_706,N_640,N_664);
nor U707 (N_707,N_656,N_610);
or U708 (N_708,N_621,N_662);
and U709 (N_709,N_601,N_618);
nor U710 (N_710,N_614,N_625);
nor U711 (N_711,N_660,N_668);
nor U712 (N_712,N_615,N_607);
and U713 (N_713,N_655,N_619);
nor U714 (N_714,N_666,N_655);
and U715 (N_715,N_632,N_638);
nor U716 (N_716,N_626,N_627);
nand U717 (N_717,N_629,N_672);
and U718 (N_718,N_631,N_659);
xnor U719 (N_719,N_635,N_671);
and U720 (N_720,N_662,N_614);
or U721 (N_721,N_641,N_630);
and U722 (N_722,N_630,N_672);
and U723 (N_723,N_653,N_666);
nand U724 (N_724,N_631,N_618);
and U725 (N_725,N_607,N_648);
or U726 (N_726,N_645,N_660);
nand U727 (N_727,N_640,N_638);
nand U728 (N_728,N_660,N_631);
and U729 (N_729,N_602,N_637);
or U730 (N_730,N_656,N_624);
or U731 (N_731,N_622,N_671);
nor U732 (N_732,N_651,N_666);
nand U733 (N_733,N_615,N_658);
and U734 (N_734,N_619,N_674);
or U735 (N_735,N_667,N_663);
and U736 (N_736,N_670,N_629);
nand U737 (N_737,N_633,N_627);
nor U738 (N_738,N_634,N_609);
nor U739 (N_739,N_641,N_637);
nand U740 (N_740,N_610,N_607);
nand U741 (N_741,N_670,N_650);
nand U742 (N_742,N_659,N_620);
nand U743 (N_743,N_611,N_622);
nor U744 (N_744,N_660,N_674);
or U745 (N_745,N_631,N_622);
or U746 (N_746,N_602,N_614);
xnor U747 (N_747,N_644,N_663);
nand U748 (N_748,N_633,N_662);
or U749 (N_749,N_609,N_605);
nor U750 (N_750,N_712,N_746);
nand U751 (N_751,N_687,N_688);
and U752 (N_752,N_708,N_743);
nand U753 (N_753,N_722,N_677);
nor U754 (N_754,N_706,N_690);
nand U755 (N_755,N_729,N_703);
nand U756 (N_756,N_714,N_733);
or U757 (N_757,N_698,N_721);
nor U758 (N_758,N_716,N_681);
and U759 (N_759,N_740,N_683);
nor U760 (N_760,N_699,N_715);
and U761 (N_761,N_747,N_713);
or U762 (N_762,N_738,N_739);
or U763 (N_763,N_749,N_696);
nand U764 (N_764,N_728,N_689);
and U765 (N_765,N_725,N_702);
nor U766 (N_766,N_727,N_705);
nand U767 (N_767,N_691,N_719);
nor U768 (N_768,N_718,N_745);
or U769 (N_769,N_742,N_726);
nor U770 (N_770,N_732,N_717);
nor U771 (N_771,N_734,N_686);
nand U772 (N_772,N_678,N_694);
nor U773 (N_773,N_704,N_744);
and U774 (N_774,N_692,N_693);
and U775 (N_775,N_735,N_695);
nor U776 (N_776,N_675,N_731);
and U777 (N_777,N_724,N_697);
nor U778 (N_778,N_709,N_676);
nand U779 (N_779,N_723,N_748);
nand U780 (N_780,N_741,N_685);
and U781 (N_781,N_679,N_720);
nor U782 (N_782,N_700,N_737);
nor U783 (N_783,N_680,N_730);
and U784 (N_784,N_701,N_736);
or U785 (N_785,N_710,N_707);
nor U786 (N_786,N_682,N_684);
nor U787 (N_787,N_711,N_747);
and U788 (N_788,N_723,N_707);
or U789 (N_789,N_675,N_730);
nor U790 (N_790,N_724,N_744);
or U791 (N_791,N_713,N_680);
nor U792 (N_792,N_741,N_695);
and U793 (N_793,N_697,N_734);
or U794 (N_794,N_708,N_724);
and U795 (N_795,N_728,N_682);
nand U796 (N_796,N_706,N_745);
and U797 (N_797,N_691,N_681);
and U798 (N_798,N_676,N_726);
nand U799 (N_799,N_715,N_732);
or U800 (N_800,N_697,N_689);
or U801 (N_801,N_675,N_710);
nand U802 (N_802,N_721,N_680);
and U803 (N_803,N_741,N_713);
nor U804 (N_804,N_729,N_730);
and U805 (N_805,N_693,N_730);
nand U806 (N_806,N_680,N_686);
and U807 (N_807,N_708,N_723);
and U808 (N_808,N_734,N_687);
or U809 (N_809,N_709,N_695);
nor U810 (N_810,N_719,N_698);
or U811 (N_811,N_732,N_691);
or U812 (N_812,N_687,N_742);
nand U813 (N_813,N_677,N_725);
or U814 (N_814,N_745,N_710);
nand U815 (N_815,N_703,N_731);
and U816 (N_816,N_689,N_703);
nand U817 (N_817,N_696,N_702);
nand U818 (N_818,N_730,N_713);
and U819 (N_819,N_721,N_703);
or U820 (N_820,N_682,N_675);
and U821 (N_821,N_745,N_701);
nor U822 (N_822,N_749,N_739);
nand U823 (N_823,N_692,N_696);
and U824 (N_824,N_719,N_675);
and U825 (N_825,N_778,N_780);
nor U826 (N_826,N_787,N_815);
nor U827 (N_827,N_796,N_797);
and U828 (N_828,N_819,N_755);
or U829 (N_829,N_800,N_767);
or U830 (N_830,N_774,N_786);
nand U831 (N_831,N_775,N_788);
or U832 (N_832,N_813,N_770);
nor U833 (N_833,N_804,N_809);
and U834 (N_834,N_758,N_803);
nor U835 (N_835,N_824,N_773);
nor U836 (N_836,N_792,N_769);
nor U837 (N_837,N_794,N_772);
or U838 (N_838,N_817,N_771);
and U839 (N_839,N_752,N_765);
nand U840 (N_840,N_761,N_753);
and U841 (N_841,N_781,N_811);
nand U842 (N_842,N_801,N_785);
nand U843 (N_843,N_757,N_782);
and U844 (N_844,N_790,N_779);
and U845 (N_845,N_760,N_820);
nor U846 (N_846,N_768,N_822);
or U847 (N_847,N_791,N_814);
nor U848 (N_848,N_756,N_764);
or U849 (N_849,N_821,N_799);
or U850 (N_850,N_795,N_807);
nand U851 (N_851,N_806,N_759);
or U852 (N_852,N_751,N_784);
nand U853 (N_853,N_776,N_805);
nor U854 (N_854,N_783,N_762);
and U855 (N_855,N_810,N_802);
nor U856 (N_856,N_777,N_818);
nand U857 (N_857,N_798,N_789);
nand U858 (N_858,N_763,N_766);
or U859 (N_859,N_750,N_793);
or U860 (N_860,N_808,N_754);
and U861 (N_861,N_816,N_823);
xor U862 (N_862,N_812,N_795);
or U863 (N_863,N_785,N_772);
nand U864 (N_864,N_798,N_764);
and U865 (N_865,N_758,N_778);
xnor U866 (N_866,N_784,N_760);
nand U867 (N_867,N_795,N_766);
or U868 (N_868,N_753,N_785);
nand U869 (N_869,N_804,N_817);
nand U870 (N_870,N_784,N_786);
nand U871 (N_871,N_758,N_792);
or U872 (N_872,N_776,N_808);
and U873 (N_873,N_757,N_797);
nand U874 (N_874,N_773,N_756);
nor U875 (N_875,N_753,N_815);
or U876 (N_876,N_805,N_802);
nor U877 (N_877,N_777,N_769);
nor U878 (N_878,N_772,N_799);
xor U879 (N_879,N_779,N_795);
nand U880 (N_880,N_799,N_812);
or U881 (N_881,N_818,N_814);
nor U882 (N_882,N_778,N_764);
or U883 (N_883,N_782,N_814);
and U884 (N_884,N_801,N_810);
nor U885 (N_885,N_801,N_819);
nand U886 (N_886,N_799,N_792);
nand U887 (N_887,N_813,N_823);
nor U888 (N_888,N_780,N_793);
or U889 (N_889,N_767,N_750);
and U890 (N_890,N_767,N_787);
nand U891 (N_891,N_754,N_805);
and U892 (N_892,N_815,N_781);
or U893 (N_893,N_753,N_804);
nand U894 (N_894,N_764,N_800);
nor U895 (N_895,N_775,N_783);
nand U896 (N_896,N_757,N_787);
and U897 (N_897,N_822,N_750);
or U898 (N_898,N_754,N_803);
nand U899 (N_899,N_760,N_750);
or U900 (N_900,N_839,N_836);
and U901 (N_901,N_825,N_861);
nand U902 (N_902,N_827,N_890);
and U903 (N_903,N_857,N_883);
or U904 (N_904,N_881,N_856);
or U905 (N_905,N_872,N_862);
nand U906 (N_906,N_850,N_886);
or U907 (N_907,N_863,N_830);
and U908 (N_908,N_875,N_864);
nor U909 (N_909,N_841,N_898);
nand U910 (N_910,N_897,N_873);
nor U911 (N_911,N_828,N_853);
nor U912 (N_912,N_895,N_888);
nand U913 (N_913,N_891,N_884);
nand U914 (N_914,N_894,N_846);
or U915 (N_915,N_867,N_869);
nor U916 (N_916,N_865,N_868);
and U917 (N_917,N_837,N_848);
nor U918 (N_918,N_852,N_847);
and U919 (N_919,N_874,N_878);
nor U920 (N_920,N_854,N_882);
nor U921 (N_921,N_860,N_870);
nand U922 (N_922,N_835,N_849);
and U923 (N_923,N_859,N_899);
nand U924 (N_924,N_829,N_892);
nor U925 (N_925,N_876,N_880);
or U926 (N_926,N_832,N_851);
or U927 (N_927,N_831,N_855);
or U928 (N_928,N_833,N_843);
nor U929 (N_929,N_896,N_866);
nor U930 (N_930,N_885,N_845);
or U931 (N_931,N_889,N_858);
or U932 (N_932,N_842,N_838);
or U933 (N_933,N_844,N_840);
nand U934 (N_934,N_834,N_887);
nor U935 (N_935,N_879,N_877);
or U936 (N_936,N_871,N_826);
and U937 (N_937,N_893,N_895);
or U938 (N_938,N_859,N_829);
nor U939 (N_939,N_829,N_846);
nor U940 (N_940,N_839,N_848);
or U941 (N_941,N_886,N_869);
nand U942 (N_942,N_891,N_848);
and U943 (N_943,N_862,N_848);
nand U944 (N_944,N_845,N_840);
or U945 (N_945,N_835,N_882);
nor U946 (N_946,N_852,N_866);
nor U947 (N_947,N_876,N_862);
nand U948 (N_948,N_884,N_849);
nor U949 (N_949,N_848,N_894);
or U950 (N_950,N_895,N_896);
nor U951 (N_951,N_890,N_886);
or U952 (N_952,N_847,N_844);
and U953 (N_953,N_857,N_892);
or U954 (N_954,N_859,N_830);
and U955 (N_955,N_827,N_857);
nor U956 (N_956,N_874,N_869);
nand U957 (N_957,N_850,N_887);
and U958 (N_958,N_872,N_850);
nor U959 (N_959,N_894,N_886);
nand U960 (N_960,N_854,N_877);
nand U961 (N_961,N_867,N_872);
nor U962 (N_962,N_889,N_832);
and U963 (N_963,N_864,N_829);
nor U964 (N_964,N_864,N_861);
or U965 (N_965,N_874,N_894);
nor U966 (N_966,N_825,N_897);
nand U967 (N_967,N_892,N_886);
nand U968 (N_968,N_858,N_891);
nor U969 (N_969,N_840,N_884);
or U970 (N_970,N_872,N_845);
and U971 (N_971,N_885,N_868);
and U972 (N_972,N_888,N_894);
nand U973 (N_973,N_856,N_838);
nor U974 (N_974,N_830,N_896);
nor U975 (N_975,N_931,N_941);
or U976 (N_976,N_908,N_906);
nand U977 (N_977,N_935,N_955);
nor U978 (N_978,N_956,N_954);
nand U979 (N_979,N_943,N_947);
nor U980 (N_980,N_934,N_926);
nand U981 (N_981,N_958,N_974);
or U982 (N_982,N_960,N_916);
or U983 (N_983,N_963,N_959);
or U984 (N_984,N_967,N_913);
nor U985 (N_985,N_927,N_921);
nor U986 (N_986,N_904,N_948);
or U987 (N_987,N_900,N_973);
or U988 (N_988,N_957,N_937);
or U989 (N_989,N_914,N_938);
and U990 (N_990,N_951,N_910);
nand U991 (N_991,N_946,N_901);
and U992 (N_992,N_928,N_968);
or U993 (N_993,N_932,N_949);
nor U994 (N_994,N_950,N_923);
nor U995 (N_995,N_970,N_915);
nand U996 (N_996,N_962,N_925);
or U997 (N_997,N_965,N_942);
nand U998 (N_998,N_912,N_966);
and U999 (N_999,N_972,N_945);
or U1000 (N_1000,N_952,N_961);
nand U1001 (N_1001,N_936,N_903);
and U1002 (N_1002,N_944,N_909);
nor U1003 (N_1003,N_940,N_917);
or U1004 (N_1004,N_933,N_905);
or U1005 (N_1005,N_919,N_911);
or U1006 (N_1006,N_907,N_918);
and U1007 (N_1007,N_964,N_902);
xor U1008 (N_1008,N_924,N_929);
nand U1009 (N_1009,N_969,N_930);
or U1010 (N_1010,N_922,N_953);
nand U1011 (N_1011,N_939,N_920);
and U1012 (N_1012,N_971,N_915);
nor U1013 (N_1013,N_900,N_941);
and U1014 (N_1014,N_948,N_943);
nor U1015 (N_1015,N_909,N_954);
nor U1016 (N_1016,N_917,N_971);
or U1017 (N_1017,N_930,N_929);
and U1018 (N_1018,N_947,N_904);
or U1019 (N_1019,N_916,N_909);
xor U1020 (N_1020,N_947,N_963);
nor U1021 (N_1021,N_931,N_959);
nor U1022 (N_1022,N_925,N_909);
and U1023 (N_1023,N_958,N_931);
nor U1024 (N_1024,N_968,N_902);
and U1025 (N_1025,N_964,N_923);
nor U1026 (N_1026,N_974,N_930);
and U1027 (N_1027,N_929,N_927);
and U1028 (N_1028,N_939,N_970);
or U1029 (N_1029,N_937,N_962);
nor U1030 (N_1030,N_925,N_927);
nand U1031 (N_1031,N_964,N_970);
or U1032 (N_1032,N_939,N_974);
nor U1033 (N_1033,N_932,N_944);
nand U1034 (N_1034,N_945,N_959);
and U1035 (N_1035,N_964,N_927);
nor U1036 (N_1036,N_951,N_942);
nand U1037 (N_1037,N_922,N_942);
nand U1038 (N_1038,N_956,N_904);
nand U1039 (N_1039,N_914,N_916);
nor U1040 (N_1040,N_945,N_948);
nor U1041 (N_1041,N_956,N_964);
nand U1042 (N_1042,N_925,N_908);
or U1043 (N_1043,N_933,N_950);
nor U1044 (N_1044,N_929,N_945);
nand U1045 (N_1045,N_966,N_911);
nand U1046 (N_1046,N_922,N_943);
nor U1047 (N_1047,N_961,N_905);
nor U1048 (N_1048,N_963,N_946);
nor U1049 (N_1049,N_951,N_939);
and U1050 (N_1050,N_1003,N_1041);
or U1051 (N_1051,N_1024,N_988);
or U1052 (N_1052,N_1025,N_1036);
and U1053 (N_1053,N_984,N_1040);
nand U1054 (N_1054,N_1042,N_980);
and U1055 (N_1055,N_1015,N_1019);
nand U1056 (N_1056,N_1038,N_981);
or U1057 (N_1057,N_994,N_975);
nor U1058 (N_1058,N_1016,N_1017);
nor U1059 (N_1059,N_999,N_1013);
and U1060 (N_1060,N_990,N_1043);
and U1061 (N_1061,N_987,N_1030);
and U1062 (N_1062,N_1006,N_1008);
nand U1063 (N_1063,N_1039,N_1002);
or U1064 (N_1064,N_1049,N_976);
nor U1065 (N_1065,N_1023,N_998);
nor U1066 (N_1066,N_996,N_1009);
or U1067 (N_1067,N_1000,N_977);
nor U1068 (N_1068,N_1048,N_1011);
nor U1069 (N_1069,N_1044,N_1026);
and U1070 (N_1070,N_989,N_1028);
nor U1071 (N_1071,N_1046,N_978);
nor U1072 (N_1072,N_1018,N_1005);
nand U1073 (N_1073,N_1032,N_1014);
nor U1074 (N_1074,N_1035,N_1034);
or U1075 (N_1075,N_1020,N_986);
and U1076 (N_1076,N_983,N_985);
and U1077 (N_1077,N_1037,N_997);
and U1078 (N_1078,N_1021,N_1022);
or U1079 (N_1079,N_992,N_1004);
nor U1080 (N_1080,N_991,N_1027);
nor U1081 (N_1081,N_982,N_1033);
nor U1082 (N_1082,N_1029,N_1031);
or U1083 (N_1083,N_979,N_1001);
or U1084 (N_1084,N_1012,N_993);
and U1085 (N_1085,N_1007,N_1045);
and U1086 (N_1086,N_1047,N_995);
and U1087 (N_1087,N_1010,N_1030);
nand U1088 (N_1088,N_1029,N_1047);
nor U1089 (N_1089,N_1022,N_1047);
nand U1090 (N_1090,N_1046,N_1016);
and U1091 (N_1091,N_985,N_981);
and U1092 (N_1092,N_1027,N_1043);
or U1093 (N_1093,N_1045,N_1036);
or U1094 (N_1094,N_991,N_993);
nand U1095 (N_1095,N_980,N_1048);
nor U1096 (N_1096,N_1028,N_1031);
or U1097 (N_1097,N_1029,N_993);
or U1098 (N_1098,N_1030,N_990);
and U1099 (N_1099,N_1026,N_998);
or U1100 (N_1100,N_995,N_991);
nor U1101 (N_1101,N_1003,N_1032);
or U1102 (N_1102,N_994,N_1000);
nand U1103 (N_1103,N_1045,N_1010);
nor U1104 (N_1104,N_1042,N_1046);
nor U1105 (N_1105,N_997,N_988);
nand U1106 (N_1106,N_1024,N_1021);
and U1107 (N_1107,N_1049,N_995);
and U1108 (N_1108,N_999,N_992);
nand U1109 (N_1109,N_1027,N_1001);
and U1110 (N_1110,N_989,N_1012);
nor U1111 (N_1111,N_1009,N_981);
and U1112 (N_1112,N_1007,N_1014);
nand U1113 (N_1113,N_994,N_1044);
nand U1114 (N_1114,N_1025,N_977);
nand U1115 (N_1115,N_1041,N_1027);
nand U1116 (N_1116,N_1037,N_1040);
nor U1117 (N_1117,N_1038,N_991);
or U1118 (N_1118,N_1009,N_979);
or U1119 (N_1119,N_1021,N_1011);
nand U1120 (N_1120,N_998,N_1002);
or U1121 (N_1121,N_999,N_1047);
or U1122 (N_1122,N_1019,N_997);
or U1123 (N_1123,N_1016,N_1045);
and U1124 (N_1124,N_1041,N_993);
or U1125 (N_1125,N_1066,N_1087);
nand U1126 (N_1126,N_1093,N_1070);
nand U1127 (N_1127,N_1111,N_1084);
nand U1128 (N_1128,N_1100,N_1057);
or U1129 (N_1129,N_1086,N_1077);
nor U1130 (N_1130,N_1109,N_1116);
and U1131 (N_1131,N_1076,N_1061);
and U1132 (N_1132,N_1092,N_1123);
or U1133 (N_1133,N_1053,N_1113);
nor U1134 (N_1134,N_1085,N_1068);
or U1135 (N_1135,N_1099,N_1107);
or U1136 (N_1136,N_1058,N_1056);
nand U1137 (N_1137,N_1078,N_1102);
and U1138 (N_1138,N_1063,N_1097);
nor U1139 (N_1139,N_1110,N_1089);
and U1140 (N_1140,N_1060,N_1082);
nand U1141 (N_1141,N_1094,N_1081);
or U1142 (N_1142,N_1095,N_1075);
and U1143 (N_1143,N_1104,N_1072);
or U1144 (N_1144,N_1059,N_1117);
nand U1145 (N_1145,N_1079,N_1055);
xnor U1146 (N_1146,N_1073,N_1115);
nor U1147 (N_1147,N_1074,N_1090);
xnor U1148 (N_1148,N_1080,N_1069);
and U1149 (N_1149,N_1103,N_1054);
or U1150 (N_1150,N_1051,N_1114);
or U1151 (N_1151,N_1120,N_1121);
or U1152 (N_1152,N_1122,N_1067);
nand U1153 (N_1153,N_1119,N_1124);
or U1154 (N_1154,N_1112,N_1108);
nand U1155 (N_1155,N_1062,N_1118);
and U1156 (N_1156,N_1052,N_1106);
and U1157 (N_1157,N_1071,N_1096);
and U1158 (N_1158,N_1064,N_1101);
or U1159 (N_1159,N_1083,N_1098);
and U1160 (N_1160,N_1065,N_1091);
and U1161 (N_1161,N_1050,N_1088);
nor U1162 (N_1162,N_1105,N_1118);
nor U1163 (N_1163,N_1096,N_1073);
nand U1164 (N_1164,N_1122,N_1100);
or U1165 (N_1165,N_1064,N_1070);
nor U1166 (N_1166,N_1065,N_1084);
nor U1167 (N_1167,N_1108,N_1078);
or U1168 (N_1168,N_1105,N_1080);
and U1169 (N_1169,N_1053,N_1058);
or U1170 (N_1170,N_1095,N_1076);
and U1171 (N_1171,N_1090,N_1115);
nor U1172 (N_1172,N_1079,N_1062);
and U1173 (N_1173,N_1056,N_1093);
nor U1174 (N_1174,N_1091,N_1110);
nor U1175 (N_1175,N_1123,N_1080);
nor U1176 (N_1176,N_1106,N_1069);
or U1177 (N_1177,N_1109,N_1059);
nor U1178 (N_1178,N_1099,N_1078);
nor U1179 (N_1179,N_1093,N_1092);
and U1180 (N_1180,N_1121,N_1081);
nor U1181 (N_1181,N_1085,N_1067);
or U1182 (N_1182,N_1124,N_1099);
nor U1183 (N_1183,N_1118,N_1056);
or U1184 (N_1184,N_1117,N_1067);
nor U1185 (N_1185,N_1075,N_1119);
nand U1186 (N_1186,N_1080,N_1066);
and U1187 (N_1187,N_1122,N_1074);
nor U1188 (N_1188,N_1104,N_1116);
and U1189 (N_1189,N_1082,N_1086);
and U1190 (N_1190,N_1062,N_1074);
nor U1191 (N_1191,N_1122,N_1077);
and U1192 (N_1192,N_1122,N_1066);
or U1193 (N_1193,N_1115,N_1094);
or U1194 (N_1194,N_1090,N_1056);
and U1195 (N_1195,N_1076,N_1065);
nor U1196 (N_1196,N_1090,N_1118);
nor U1197 (N_1197,N_1091,N_1117);
nand U1198 (N_1198,N_1061,N_1117);
nand U1199 (N_1199,N_1051,N_1058);
and U1200 (N_1200,N_1174,N_1180);
nor U1201 (N_1201,N_1187,N_1172);
nand U1202 (N_1202,N_1179,N_1188);
or U1203 (N_1203,N_1152,N_1175);
and U1204 (N_1204,N_1166,N_1154);
nand U1205 (N_1205,N_1182,N_1190);
nand U1206 (N_1206,N_1153,N_1181);
nand U1207 (N_1207,N_1135,N_1165);
and U1208 (N_1208,N_1127,N_1164);
nand U1209 (N_1209,N_1196,N_1160);
nor U1210 (N_1210,N_1147,N_1146);
and U1211 (N_1211,N_1145,N_1134);
nand U1212 (N_1212,N_1198,N_1163);
and U1213 (N_1213,N_1197,N_1126);
nor U1214 (N_1214,N_1125,N_1171);
nor U1215 (N_1215,N_1142,N_1162);
or U1216 (N_1216,N_1138,N_1159);
and U1217 (N_1217,N_1143,N_1177);
nand U1218 (N_1218,N_1191,N_1149);
nand U1219 (N_1219,N_1133,N_1132);
or U1220 (N_1220,N_1140,N_1129);
and U1221 (N_1221,N_1167,N_1148);
or U1222 (N_1222,N_1128,N_1192);
and U1223 (N_1223,N_1168,N_1194);
and U1224 (N_1224,N_1151,N_1186);
and U1225 (N_1225,N_1137,N_1173);
and U1226 (N_1226,N_1176,N_1189);
and U1227 (N_1227,N_1195,N_1158);
nand U1228 (N_1228,N_1185,N_1183);
or U1229 (N_1229,N_1193,N_1178);
or U1230 (N_1230,N_1130,N_1157);
and U1231 (N_1231,N_1155,N_1184);
xor U1232 (N_1232,N_1156,N_1161);
and U1233 (N_1233,N_1150,N_1170);
and U1234 (N_1234,N_1169,N_1144);
and U1235 (N_1235,N_1139,N_1136);
and U1236 (N_1236,N_1141,N_1131);
and U1237 (N_1237,N_1199,N_1195);
or U1238 (N_1238,N_1192,N_1156);
or U1239 (N_1239,N_1146,N_1198);
xor U1240 (N_1240,N_1152,N_1146);
nor U1241 (N_1241,N_1176,N_1193);
and U1242 (N_1242,N_1191,N_1193);
and U1243 (N_1243,N_1133,N_1172);
nand U1244 (N_1244,N_1193,N_1172);
or U1245 (N_1245,N_1141,N_1165);
nor U1246 (N_1246,N_1197,N_1129);
and U1247 (N_1247,N_1142,N_1177);
nor U1248 (N_1248,N_1159,N_1127);
or U1249 (N_1249,N_1172,N_1151);
nor U1250 (N_1250,N_1163,N_1134);
nor U1251 (N_1251,N_1152,N_1194);
nor U1252 (N_1252,N_1170,N_1187);
nor U1253 (N_1253,N_1155,N_1189);
and U1254 (N_1254,N_1134,N_1192);
nor U1255 (N_1255,N_1188,N_1170);
or U1256 (N_1256,N_1146,N_1134);
and U1257 (N_1257,N_1179,N_1150);
or U1258 (N_1258,N_1197,N_1175);
and U1259 (N_1259,N_1198,N_1166);
nand U1260 (N_1260,N_1186,N_1179);
nand U1261 (N_1261,N_1181,N_1194);
or U1262 (N_1262,N_1135,N_1184);
nor U1263 (N_1263,N_1170,N_1176);
nand U1264 (N_1264,N_1134,N_1197);
and U1265 (N_1265,N_1195,N_1191);
nor U1266 (N_1266,N_1139,N_1164);
and U1267 (N_1267,N_1171,N_1149);
and U1268 (N_1268,N_1179,N_1199);
and U1269 (N_1269,N_1192,N_1180);
and U1270 (N_1270,N_1179,N_1178);
or U1271 (N_1271,N_1139,N_1191);
or U1272 (N_1272,N_1194,N_1138);
and U1273 (N_1273,N_1153,N_1129);
or U1274 (N_1274,N_1136,N_1189);
and U1275 (N_1275,N_1252,N_1246);
or U1276 (N_1276,N_1250,N_1207);
or U1277 (N_1277,N_1230,N_1239);
nand U1278 (N_1278,N_1208,N_1211);
nand U1279 (N_1279,N_1270,N_1214);
nand U1280 (N_1280,N_1267,N_1272);
or U1281 (N_1281,N_1225,N_1259);
nand U1282 (N_1282,N_1234,N_1254);
or U1283 (N_1283,N_1247,N_1274);
nand U1284 (N_1284,N_1256,N_1237);
nor U1285 (N_1285,N_1258,N_1242);
nand U1286 (N_1286,N_1243,N_1248);
or U1287 (N_1287,N_1210,N_1269);
nor U1288 (N_1288,N_1229,N_1264);
or U1289 (N_1289,N_1261,N_1226);
nor U1290 (N_1290,N_1203,N_1236);
and U1291 (N_1291,N_1268,N_1212);
or U1292 (N_1292,N_1265,N_1201);
and U1293 (N_1293,N_1233,N_1257);
or U1294 (N_1294,N_1202,N_1260);
nand U1295 (N_1295,N_1245,N_1266);
nand U1296 (N_1296,N_1231,N_1205);
and U1297 (N_1297,N_1213,N_1240);
or U1298 (N_1298,N_1232,N_1228);
nand U1299 (N_1299,N_1204,N_1218);
nand U1300 (N_1300,N_1263,N_1215);
nand U1301 (N_1301,N_1222,N_1209);
nor U1302 (N_1302,N_1255,N_1235);
nand U1303 (N_1303,N_1262,N_1253);
nand U1304 (N_1304,N_1224,N_1216);
and U1305 (N_1305,N_1251,N_1223);
or U1306 (N_1306,N_1219,N_1244);
nor U1307 (N_1307,N_1221,N_1227);
or U1308 (N_1308,N_1206,N_1241);
or U1309 (N_1309,N_1200,N_1271);
nand U1310 (N_1310,N_1217,N_1249);
nor U1311 (N_1311,N_1220,N_1238);
or U1312 (N_1312,N_1273,N_1251);
or U1313 (N_1313,N_1239,N_1245);
or U1314 (N_1314,N_1210,N_1238);
or U1315 (N_1315,N_1224,N_1274);
or U1316 (N_1316,N_1206,N_1201);
and U1317 (N_1317,N_1202,N_1224);
nor U1318 (N_1318,N_1267,N_1224);
nand U1319 (N_1319,N_1267,N_1223);
nor U1320 (N_1320,N_1229,N_1266);
nand U1321 (N_1321,N_1274,N_1270);
and U1322 (N_1322,N_1225,N_1208);
and U1323 (N_1323,N_1218,N_1203);
nand U1324 (N_1324,N_1226,N_1267);
and U1325 (N_1325,N_1215,N_1228);
and U1326 (N_1326,N_1211,N_1238);
or U1327 (N_1327,N_1246,N_1200);
or U1328 (N_1328,N_1207,N_1230);
nor U1329 (N_1329,N_1244,N_1266);
nand U1330 (N_1330,N_1245,N_1249);
and U1331 (N_1331,N_1225,N_1233);
and U1332 (N_1332,N_1263,N_1209);
nor U1333 (N_1333,N_1211,N_1201);
or U1334 (N_1334,N_1201,N_1246);
and U1335 (N_1335,N_1203,N_1273);
nor U1336 (N_1336,N_1206,N_1233);
nor U1337 (N_1337,N_1242,N_1252);
or U1338 (N_1338,N_1242,N_1217);
and U1339 (N_1339,N_1218,N_1267);
nand U1340 (N_1340,N_1238,N_1222);
nor U1341 (N_1341,N_1229,N_1223);
or U1342 (N_1342,N_1230,N_1227);
nand U1343 (N_1343,N_1204,N_1219);
nand U1344 (N_1344,N_1250,N_1265);
and U1345 (N_1345,N_1237,N_1253);
or U1346 (N_1346,N_1205,N_1248);
nand U1347 (N_1347,N_1268,N_1216);
nor U1348 (N_1348,N_1219,N_1243);
and U1349 (N_1349,N_1270,N_1207);
or U1350 (N_1350,N_1311,N_1315);
nor U1351 (N_1351,N_1305,N_1327);
nor U1352 (N_1352,N_1286,N_1336);
and U1353 (N_1353,N_1340,N_1320);
and U1354 (N_1354,N_1343,N_1275);
or U1355 (N_1355,N_1347,N_1301);
nor U1356 (N_1356,N_1283,N_1285);
and U1357 (N_1357,N_1280,N_1299);
or U1358 (N_1358,N_1338,N_1323);
and U1359 (N_1359,N_1276,N_1335);
nand U1360 (N_1360,N_1328,N_1317);
and U1361 (N_1361,N_1304,N_1284);
and U1362 (N_1362,N_1331,N_1298);
or U1363 (N_1363,N_1341,N_1308);
and U1364 (N_1364,N_1310,N_1289);
nor U1365 (N_1365,N_1307,N_1291);
or U1366 (N_1366,N_1316,N_1334);
and U1367 (N_1367,N_1344,N_1313);
nor U1368 (N_1368,N_1303,N_1296);
nor U1369 (N_1369,N_1321,N_1325);
and U1370 (N_1370,N_1337,N_1306);
and U1371 (N_1371,N_1281,N_1339);
nor U1372 (N_1372,N_1302,N_1332);
and U1373 (N_1373,N_1348,N_1312);
nand U1374 (N_1374,N_1282,N_1319);
nor U1375 (N_1375,N_1279,N_1322);
nand U1376 (N_1376,N_1346,N_1326);
or U1377 (N_1377,N_1342,N_1293);
nor U1378 (N_1378,N_1318,N_1333);
and U1379 (N_1379,N_1295,N_1278);
and U1380 (N_1380,N_1292,N_1287);
and U1381 (N_1381,N_1277,N_1324);
nor U1382 (N_1382,N_1297,N_1288);
or U1383 (N_1383,N_1314,N_1345);
nand U1384 (N_1384,N_1300,N_1294);
nor U1385 (N_1385,N_1349,N_1329);
nand U1386 (N_1386,N_1290,N_1330);
or U1387 (N_1387,N_1309,N_1317);
nand U1388 (N_1388,N_1288,N_1289);
nand U1389 (N_1389,N_1333,N_1302);
nand U1390 (N_1390,N_1314,N_1278);
or U1391 (N_1391,N_1322,N_1334);
nand U1392 (N_1392,N_1294,N_1291);
or U1393 (N_1393,N_1337,N_1323);
or U1394 (N_1394,N_1304,N_1283);
or U1395 (N_1395,N_1303,N_1333);
and U1396 (N_1396,N_1316,N_1311);
or U1397 (N_1397,N_1304,N_1308);
nand U1398 (N_1398,N_1304,N_1316);
nor U1399 (N_1399,N_1327,N_1338);
or U1400 (N_1400,N_1332,N_1310);
or U1401 (N_1401,N_1275,N_1283);
or U1402 (N_1402,N_1324,N_1347);
and U1403 (N_1403,N_1338,N_1340);
nand U1404 (N_1404,N_1337,N_1300);
nor U1405 (N_1405,N_1277,N_1328);
or U1406 (N_1406,N_1283,N_1345);
nor U1407 (N_1407,N_1287,N_1282);
nand U1408 (N_1408,N_1330,N_1335);
or U1409 (N_1409,N_1327,N_1346);
nor U1410 (N_1410,N_1337,N_1286);
nor U1411 (N_1411,N_1314,N_1293);
nor U1412 (N_1412,N_1333,N_1319);
or U1413 (N_1413,N_1287,N_1325);
nor U1414 (N_1414,N_1344,N_1299);
or U1415 (N_1415,N_1329,N_1312);
nand U1416 (N_1416,N_1305,N_1333);
nor U1417 (N_1417,N_1280,N_1282);
nand U1418 (N_1418,N_1281,N_1340);
nor U1419 (N_1419,N_1308,N_1297);
nand U1420 (N_1420,N_1283,N_1322);
nand U1421 (N_1421,N_1342,N_1347);
nor U1422 (N_1422,N_1320,N_1334);
nor U1423 (N_1423,N_1288,N_1311);
and U1424 (N_1424,N_1289,N_1338);
nand U1425 (N_1425,N_1364,N_1357);
or U1426 (N_1426,N_1393,N_1422);
or U1427 (N_1427,N_1385,N_1352);
and U1428 (N_1428,N_1374,N_1424);
or U1429 (N_1429,N_1367,N_1376);
nor U1430 (N_1430,N_1363,N_1396);
nor U1431 (N_1431,N_1414,N_1401);
nand U1432 (N_1432,N_1377,N_1366);
nor U1433 (N_1433,N_1388,N_1353);
nor U1434 (N_1434,N_1407,N_1409);
nor U1435 (N_1435,N_1423,N_1413);
and U1436 (N_1436,N_1380,N_1359);
and U1437 (N_1437,N_1408,N_1403);
and U1438 (N_1438,N_1356,N_1389);
nor U1439 (N_1439,N_1382,N_1369);
or U1440 (N_1440,N_1412,N_1383);
nor U1441 (N_1441,N_1420,N_1417);
nand U1442 (N_1442,N_1370,N_1371);
nand U1443 (N_1443,N_1394,N_1418);
and U1444 (N_1444,N_1368,N_1354);
and U1445 (N_1445,N_1379,N_1421);
or U1446 (N_1446,N_1378,N_1386);
nor U1447 (N_1447,N_1399,N_1406);
nand U1448 (N_1448,N_1375,N_1381);
or U1449 (N_1449,N_1402,N_1372);
and U1450 (N_1450,N_1404,N_1365);
or U1451 (N_1451,N_1384,N_1361);
nand U1452 (N_1452,N_1398,N_1387);
nand U1453 (N_1453,N_1400,N_1360);
and U1454 (N_1454,N_1355,N_1411);
nand U1455 (N_1455,N_1416,N_1390);
and U1456 (N_1456,N_1351,N_1405);
nand U1457 (N_1457,N_1350,N_1391);
nor U1458 (N_1458,N_1419,N_1392);
and U1459 (N_1459,N_1395,N_1397);
nand U1460 (N_1460,N_1415,N_1410);
or U1461 (N_1461,N_1362,N_1373);
nor U1462 (N_1462,N_1358,N_1392);
nand U1463 (N_1463,N_1417,N_1351);
nor U1464 (N_1464,N_1387,N_1379);
nand U1465 (N_1465,N_1359,N_1391);
or U1466 (N_1466,N_1371,N_1379);
or U1467 (N_1467,N_1357,N_1421);
or U1468 (N_1468,N_1366,N_1418);
and U1469 (N_1469,N_1415,N_1421);
and U1470 (N_1470,N_1378,N_1396);
nor U1471 (N_1471,N_1395,N_1413);
nand U1472 (N_1472,N_1421,N_1380);
nand U1473 (N_1473,N_1411,N_1352);
and U1474 (N_1474,N_1357,N_1361);
or U1475 (N_1475,N_1397,N_1421);
nand U1476 (N_1476,N_1408,N_1378);
nand U1477 (N_1477,N_1387,N_1409);
nand U1478 (N_1478,N_1358,N_1424);
or U1479 (N_1479,N_1405,N_1375);
nand U1480 (N_1480,N_1416,N_1362);
nand U1481 (N_1481,N_1353,N_1408);
or U1482 (N_1482,N_1400,N_1396);
and U1483 (N_1483,N_1374,N_1368);
nand U1484 (N_1484,N_1355,N_1373);
nand U1485 (N_1485,N_1388,N_1371);
or U1486 (N_1486,N_1376,N_1362);
and U1487 (N_1487,N_1406,N_1389);
and U1488 (N_1488,N_1354,N_1378);
and U1489 (N_1489,N_1354,N_1391);
nor U1490 (N_1490,N_1381,N_1360);
and U1491 (N_1491,N_1409,N_1404);
nand U1492 (N_1492,N_1410,N_1391);
or U1493 (N_1493,N_1381,N_1369);
and U1494 (N_1494,N_1421,N_1367);
or U1495 (N_1495,N_1422,N_1414);
nand U1496 (N_1496,N_1421,N_1375);
nand U1497 (N_1497,N_1417,N_1382);
or U1498 (N_1498,N_1361,N_1387);
nand U1499 (N_1499,N_1403,N_1367);
nor U1500 (N_1500,N_1451,N_1497);
and U1501 (N_1501,N_1486,N_1456);
or U1502 (N_1502,N_1446,N_1458);
nor U1503 (N_1503,N_1481,N_1485);
and U1504 (N_1504,N_1496,N_1487);
or U1505 (N_1505,N_1474,N_1489);
nand U1506 (N_1506,N_1453,N_1444);
nor U1507 (N_1507,N_1478,N_1429);
or U1508 (N_1508,N_1435,N_1493);
nand U1509 (N_1509,N_1498,N_1459);
nor U1510 (N_1510,N_1436,N_1491);
or U1511 (N_1511,N_1438,N_1440);
or U1512 (N_1512,N_1442,N_1472);
and U1513 (N_1513,N_1462,N_1476);
nor U1514 (N_1514,N_1466,N_1431);
nor U1515 (N_1515,N_1477,N_1482);
nor U1516 (N_1516,N_1432,N_1441);
nor U1517 (N_1517,N_1484,N_1465);
nor U1518 (N_1518,N_1426,N_1470);
or U1519 (N_1519,N_1471,N_1475);
nor U1520 (N_1520,N_1430,N_1499);
xnor U1521 (N_1521,N_1463,N_1488);
or U1522 (N_1522,N_1461,N_1437);
and U1523 (N_1523,N_1448,N_1445);
nor U1524 (N_1524,N_1464,N_1450);
nor U1525 (N_1525,N_1490,N_1495);
or U1526 (N_1526,N_1479,N_1434);
and U1527 (N_1527,N_1433,N_1443);
or U1528 (N_1528,N_1473,N_1494);
nor U1529 (N_1529,N_1428,N_1483);
nor U1530 (N_1530,N_1468,N_1469);
nor U1531 (N_1531,N_1467,N_1447);
xor U1532 (N_1532,N_1455,N_1460);
and U1533 (N_1533,N_1492,N_1425);
and U1534 (N_1534,N_1439,N_1427);
or U1535 (N_1535,N_1454,N_1457);
nor U1536 (N_1536,N_1449,N_1480);
nor U1537 (N_1537,N_1452,N_1425);
nand U1538 (N_1538,N_1488,N_1430);
or U1539 (N_1539,N_1480,N_1485);
nand U1540 (N_1540,N_1476,N_1431);
xnor U1541 (N_1541,N_1440,N_1477);
nand U1542 (N_1542,N_1492,N_1496);
nand U1543 (N_1543,N_1480,N_1487);
nand U1544 (N_1544,N_1459,N_1467);
nor U1545 (N_1545,N_1469,N_1488);
nand U1546 (N_1546,N_1471,N_1455);
or U1547 (N_1547,N_1495,N_1480);
nand U1548 (N_1548,N_1470,N_1495);
and U1549 (N_1549,N_1494,N_1438);
and U1550 (N_1550,N_1434,N_1488);
nand U1551 (N_1551,N_1490,N_1462);
or U1552 (N_1552,N_1426,N_1435);
nor U1553 (N_1553,N_1499,N_1441);
nand U1554 (N_1554,N_1469,N_1464);
or U1555 (N_1555,N_1447,N_1466);
and U1556 (N_1556,N_1467,N_1480);
and U1557 (N_1557,N_1491,N_1486);
nand U1558 (N_1558,N_1483,N_1482);
nor U1559 (N_1559,N_1450,N_1461);
or U1560 (N_1560,N_1460,N_1486);
nor U1561 (N_1561,N_1498,N_1436);
or U1562 (N_1562,N_1450,N_1460);
nand U1563 (N_1563,N_1451,N_1442);
or U1564 (N_1564,N_1493,N_1487);
nor U1565 (N_1565,N_1457,N_1479);
or U1566 (N_1566,N_1459,N_1427);
and U1567 (N_1567,N_1485,N_1464);
nor U1568 (N_1568,N_1468,N_1470);
and U1569 (N_1569,N_1464,N_1458);
nor U1570 (N_1570,N_1435,N_1437);
nand U1571 (N_1571,N_1442,N_1436);
nand U1572 (N_1572,N_1499,N_1495);
nand U1573 (N_1573,N_1486,N_1461);
or U1574 (N_1574,N_1433,N_1455);
nand U1575 (N_1575,N_1524,N_1547);
or U1576 (N_1576,N_1514,N_1566);
xnor U1577 (N_1577,N_1549,N_1507);
nand U1578 (N_1578,N_1546,N_1518);
and U1579 (N_1579,N_1517,N_1567);
or U1580 (N_1580,N_1569,N_1557);
or U1581 (N_1581,N_1564,N_1541);
or U1582 (N_1582,N_1553,N_1538);
nor U1583 (N_1583,N_1555,N_1565);
and U1584 (N_1584,N_1537,N_1563);
nand U1585 (N_1585,N_1502,N_1571);
or U1586 (N_1586,N_1520,N_1523);
xnor U1587 (N_1587,N_1534,N_1521);
nor U1588 (N_1588,N_1568,N_1505);
nand U1589 (N_1589,N_1526,N_1551);
nand U1590 (N_1590,N_1554,N_1550);
nor U1591 (N_1591,N_1570,N_1515);
nand U1592 (N_1592,N_1516,N_1530);
or U1593 (N_1593,N_1529,N_1558);
or U1594 (N_1594,N_1504,N_1532);
nor U1595 (N_1595,N_1542,N_1562);
nor U1596 (N_1596,N_1508,N_1556);
nand U1597 (N_1597,N_1533,N_1548);
and U1598 (N_1598,N_1510,N_1544);
and U1599 (N_1599,N_1574,N_1528);
nand U1600 (N_1600,N_1573,N_1561);
and U1601 (N_1601,N_1513,N_1559);
nand U1602 (N_1602,N_1540,N_1535);
nand U1603 (N_1603,N_1527,N_1543);
nand U1604 (N_1604,N_1531,N_1560);
or U1605 (N_1605,N_1545,N_1503);
and U1606 (N_1606,N_1500,N_1552);
and U1607 (N_1607,N_1511,N_1522);
nor U1608 (N_1608,N_1572,N_1501);
nor U1609 (N_1609,N_1536,N_1506);
nor U1610 (N_1610,N_1539,N_1525);
or U1611 (N_1611,N_1512,N_1519);
nor U1612 (N_1612,N_1509,N_1544);
or U1613 (N_1613,N_1502,N_1569);
and U1614 (N_1614,N_1517,N_1515);
nor U1615 (N_1615,N_1567,N_1536);
or U1616 (N_1616,N_1535,N_1510);
nor U1617 (N_1617,N_1556,N_1543);
and U1618 (N_1618,N_1573,N_1574);
nor U1619 (N_1619,N_1551,N_1566);
nand U1620 (N_1620,N_1561,N_1564);
and U1621 (N_1621,N_1564,N_1530);
and U1622 (N_1622,N_1520,N_1571);
and U1623 (N_1623,N_1511,N_1521);
or U1624 (N_1624,N_1555,N_1539);
nor U1625 (N_1625,N_1561,N_1515);
nor U1626 (N_1626,N_1552,N_1567);
nor U1627 (N_1627,N_1530,N_1513);
nand U1628 (N_1628,N_1549,N_1529);
nand U1629 (N_1629,N_1527,N_1542);
and U1630 (N_1630,N_1554,N_1508);
nor U1631 (N_1631,N_1509,N_1515);
and U1632 (N_1632,N_1566,N_1500);
nor U1633 (N_1633,N_1567,N_1521);
or U1634 (N_1634,N_1541,N_1512);
and U1635 (N_1635,N_1560,N_1519);
nor U1636 (N_1636,N_1517,N_1550);
nand U1637 (N_1637,N_1534,N_1574);
and U1638 (N_1638,N_1558,N_1554);
nor U1639 (N_1639,N_1537,N_1560);
and U1640 (N_1640,N_1514,N_1519);
and U1641 (N_1641,N_1543,N_1561);
nand U1642 (N_1642,N_1542,N_1573);
or U1643 (N_1643,N_1513,N_1574);
nor U1644 (N_1644,N_1561,N_1521);
nor U1645 (N_1645,N_1556,N_1515);
or U1646 (N_1646,N_1565,N_1543);
and U1647 (N_1647,N_1501,N_1555);
or U1648 (N_1648,N_1529,N_1563);
nor U1649 (N_1649,N_1500,N_1548);
nand U1650 (N_1650,N_1622,N_1609);
nand U1651 (N_1651,N_1586,N_1633);
or U1652 (N_1652,N_1589,N_1604);
nor U1653 (N_1653,N_1614,N_1642);
nor U1654 (N_1654,N_1587,N_1644);
and U1655 (N_1655,N_1634,N_1635);
nand U1656 (N_1656,N_1582,N_1619);
nor U1657 (N_1657,N_1583,N_1643);
and U1658 (N_1658,N_1646,N_1623);
or U1659 (N_1659,N_1600,N_1641);
nor U1660 (N_1660,N_1597,N_1649);
nand U1661 (N_1661,N_1618,N_1610);
or U1662 (N_1662,N_1601,N_1645);
or U1663 (N_1663,N_1599,N_1588);
nand U1664 (N_1664,N_1607,N_1637);
and U1665 (N_1665,N_1640,N_1580);
nand U1666 (N_1666,N_1603,N_1581);
or U1667 (N_1667,N_1579,N_1590);
nor U1668 (N_1668,N_1632,N_1611);
nor U1669 (N_1669,N_1596,N_1575);
nor U1670 (N_1670,N_1605,N_1598);
nor U1671 (N_1671,N_1647,N_1636);
nor U1672 (N_1672,N_1584,N_1578);
and U1673 (N_1673,N_1576,N_1577);
nor U1674 (N_1674,N_1608,N_1594);
and U1675 (N_1675,N_1592,N_1648);
and U1676 (N_1676,N_1616,N_1629);
nand U1677 (N_1677,N_1628,N_1585);
and U1678 (N_1678,N_1593,N_1620);
nor U1679 (N_1679,N_1602,N_1630);
nor U1680 (N_1680,N_1621,N_1625);
and U1681 (N_1681,N_1606,N_1631);
nor U1682 (N_1682,N_1615,N_1612);
or U1683 (N_1683,N_1617,N_1613);
or U1684 (N_1684,N_1627,N_1639);
or U1685 (N_1685,N_1638,N_1626);
nor U1686 (N_1686,N_1595,N_1591);
nand U1687 (N_1687,N_1624,N_1595);
nor U1688 (N_1688,N_1600,N_1581);
or U1689 (N_1689,N_1648,N_1636);
or U1690 (N_1690,N_1596,N_1590);
or U1691 (N_1691,N_1646,N_1607);
nand U1692 (N_1692,N_1610,N_1622);
nand U1693 (N_1693,N_1644,N_1617);
or U1694 (N_1694,N_1635,N_1621);
nand U1695 (N_1695,N_1617,N_1615);
and U1696 (N_1696,N_1615,N_1597);
or U1697 (N_1697,N_1602,N_1582);
xnor U1698 (N_1698,N_1624,N_1588);
nand U1699 (N_1699,N_1637,N_1583);
nor U1700 (N_1700,N_1602,N_1643);
nor U1701 (N_1701,N_1616,N_1599);
xnor U1702 (N_1702,N_1619,N_1589);
or U1703 (N_1703,N_1580,N_1596);
nand U1704 (N_1704,N_1646,N_1582);
nand U1705 (N_1705,N_1617,N_1607);
or U1706 (N_1706,N_1633,N_1600);
nand U1707 (N_1707,N_1628,N_1637);
nand U1708 (N_1708,N_1637,N_1612);
nand U1709 (N_1709,N_1615,N_1599);
nand U1710 (N_1710,N_1583,N_1585);
nor U1711 (N_1711,N_1608,N_1634);
or U1712 (N_1712,N_1637,N_1620);
nor U1713 (N_1713,N_1643,N_1611);
and U1714 (N_1714,N_1585,N_1616);
nand U1715 (N_1715,N_1620,N_1594);
nand U1716 (N_1716,N_1603,N_1637);
or U1717 (N_1717,N_1614,N_1583);
nor U1718 (N_1718,N_1592,N_1623);
and U1719 (N_1719,N_1639,N_1598);
or U1720 (N_1720,N_1584,N_1605);
nand U1721 (N_1721,N_1580,N_1606);
nor U1722 (N_1722,N_1581,N_1648);
nand U1723 (N_1723,N_1622,N_1624);
nor U1724 (N_1724,N_1591,N_1622);
nand U1725 (N_1725,N_1700,N_1666);
and U1726 (N_1726,N_1652,N_1665);
and U1727 (N_1727,N_1679,N_1704);
nand U1728 (N_1728,N_1718,N_1702);
nand U1729 (N_1729,N_1717,N_1721);
and U1730 (N_1730,N_1654,N_1691);
nand U1731 (N_1731,N_1663,N_1664);
nand U1732 (N_1732,N_1694,N_1667);
and U1733 (N_1733,N_1687,N_1705);
nand U1734 (N_1734,N_1707,N_1675);
and U1735 (N_1735,N_1678,N_1713);
nor U1736 (N_1736,N_1703,N_1681);
or U1737 (N_1737,N_1670,N_1716);
nand U1738 (N_1738,N_1708,N_1661);
and U1739 (N_1739,N_1680,N_1651);
or U1740 (N_1740,N_1697,N_1690);
nor U1741 (N_1741,N_1698,N_1706);
nor U1742 (N_1742,N_1673,N_1709);
nand U1743 (N_1743,N_1701,N_1671);
and U1744 (N_1744,N_1699,N_1696);
or U1745 (N_1745,N_1722,N_1685);
nand U1746 (N_1746,N_1719,N_1688);
nand U1747 (N_1747,N_1659,N_1658);
or U1748 (N_1748,N_1668,N_1683);
or U1749 (N_1749,N_1711,N_1712);
nor U1750 (N_1750,N_1672,N_1662);
nor U1751 (N_1751,N_1692,N_1723);
and U1752 (N_1752,N_1660,N_1650);
or U1753 (N_1753,N_1710,N_1677);
nor U1754 (N_1754,N_1724,N_1656);
nor U1755 (N_1755,N_1655,N_1714);
nor U1756 (N_1756,N_1676,N_1669);
nor U1757 (N_1757,N_1686,N_1695);
and U1758 (N_1758,N_1653,N_1720);
nor U1759 (N_1759,N_1689,N_1693);
or U1760 (N_1760,N_1715,N_1674);
nand U1761 (N_1761,N_1684,N_1657);
and U1762 (N_1762,N_1682,N_1675);
and U1763 (N_1763,N_1724,N_1670);
nand U1764 (N_1764,N_1670,N_1697);
nor U1765 (N_1765,N_1703,N_1685);
nand U1766 (N_1766,N_1697,N_1666);
nand U1767 (N_1767,N_1661,N_1679);
and U1768 (N_1768,N_1669,N_1667);
nand U1769 (N_1769,N_1699,N_1702);
nor U1770 (N_1770,N_1690,N_1715);
or U1771 (N_1771,N_1703,N_1701);
nand U1772 (N_1772,N_1709,N_1711);
xor U1773 (N_1773,N_1668,N_1691);
and U1774 (N_1774,N_1676,N_1678);
or U1775 (N_1775,N_1709,N_1681);
or U1776 (N_1776,N_1714,N_1693);
nand U1777 (N_1777,N_1651,N_1686);
nand U1778 (N_1778,N_1709,N_1670);
and U1779 (N_1779,N_1687,N_1685);
and U1780 (N_1780,N_1720,N_1676);
nor U1781 (N_1781,N_1677,N_1683);
nor U1782 (N_1782,N_1710,N_1708);
or U1783 (N_1783,N_1696,N_1695);
or U1784 (N_1784,N_1698,N_1696);
or U1785 (N_1785,N_1658,N_1699);
or U1786 (N_1786,N_1689,N_1722);
nand U1787 (N_1787,N_1713,N_1720);
nand U1788 (N_1788,N_1687,N_1651);
and U1789 (N_1789,N_1675,N_1698);
or U1790 (N_1790,N_1687,N_1708);
and U1791 (N_1791,N_1698,N_1714);
or U1792 (N_1792,N_1666,N_1699);
and U1793 (N_1793,N_1662,N_1714);
or U1794 (N_1794,N_1676,N_1697);
or U1795 (N_1795,N_1655,N_1674);
or U1796 (N_1796,N_1672,N_1679);
and U1797 (N_1797,N_1662,N_1669);
or U1798 (N_1798,N_1679,N_1692);
xnor U1799 (N_1799,N_1697,N_1669);
nand U1800 (N_1800,N_1773,N_1798);
nor U1801 (N_1801,N_1774,N_1776);
or U1802 (N_1802,N_1786,N_1756);
nand U1803 (N_1803,N_1779,N_1769);
nor U1804 (N_1804,N_1797,N_1772);
and U1805 (N_1805,N_1759,N_1780);
and U1806 (N_1806,N_1754,N_1745);
or U1807 (N_1807,N_1738,N_1770);
nor U1808 (N_1808,N_1741,N_1755);
and U1809 (N_1809,N_1758,N_1733);
or U1810 (N_1810,N_1775,N_1761);
nor U1811 (N_1811,N_1732,N_1746);
nand U1812 (N_1812,N_1760,N_1729);
xnor U1813 (N_1813,N_1739,N_1793);
and U1814 (N_1814,N_1791,N_1734);
and U1815 (N_1815,N_1743,N_1744);
nor U1816 (N_1816,N_1777,N_1790);
nor U1817 (N_1817,N_1768,N_1787);
and U1818 (N_1818,N_1767,N_1789);
nand U1819 (N_1819,N_1783,N_1725);
and U1820 (N_1820,N_1792,N_1765);
or U1821 (N_1821,N_1749,N_1751);
nand U1822 (N_1822,N_1764,N_1735);
nor U1823 (N_1823,N_1736,N_1771);
nor U1824 (N_1824,N_1796,N_1752);
nor U1825 (N_1825,N_1747,N_1757);
or U1826 (N_1826,N_1784,N_1728);
nor U1827 (N_1827,N_1748,N_1781);
and U1828 (N_1828,N_1799,N_1766);
nand U1829 (N_1829,N_1794,N_1726);
and U1830 (N_1830,N_1795,N_1788);
or U1831 (N_1831,N_1737,N_1782);
and U1832 (N_1832,N_1750,N_1778);
nand U1833 (N_1833,N_1730,N_1740);
and U1834 (N_1834,N_1727,N_1762);
nor U1835 (N_1835,N_1731,N_1763);
and U1836 (N_1836,N_1753,N_1785);
and U1837 (N_1837,N_1742,N_1760);
nor U1838 (N_1838,N_1732,N_1755);
and U1839 (N_1839,N_1782,N_1764);
or U1840 (N_1840,N_1779,N_1734);
nor U1841 (N_1841,N_1765,N_1764);
and U1842 (N_1842,N_1796,N_1739);
and U1843 (N_1843,N_1751,N_1784);
nor U1844 (N_1844,N_1791,N_1794);
nand U1845 (N_1845,N_1731,N_1742);
or U1846 (N_1846,N_1767,N_1775);
and U1847 (N_1847,N_1741,N_1757);
xnor U1848 (N_1848,N_1774,N_1761);
or U1849 (N_1849,N_1795,N_1754);
and U1850 (N_1850,N_1750,N_1760);
or U1851 (N_1851,N_1743,N_1738);
and U1852 (N_1852,N_1788,N_1729);
nand U1853 (N_1853,N_1725,N_1765);
and U1854 (N_1854,N_1777,N_1787);
nor U1855 (N_1855,N_1777,N_1740);
and U1856 (N_1856,N_1797,N_1760);
and U1857 (N_1857,N_1782,N_1777);
nor U1858 (N_1858,N_1788,N_1761);
nor U1859 (N_1859,N_1769,N_1784);
and U1860 (N_1860,N_1764,N_1729);
and U1861 (N_1861,N_1753,N_1784);
or U1862 (N_1862,N_1784,N_1736);
or U1863 (N_1863,N_1759,N_1776);
or U1864 (N_1864,N_1795,N_1777);
nor U1865 (N_1865,N_1797,N_1737);
nor U1866 (N_1866,N_1772,N_1730);
and U1867 (N_1867,N_1778,N_1793);
and U1868 (N_1868,N_1761,N_1770);
nand U1869 (N_1869,N_1743,N_1791);
and U1870 (N_1870,N_1735,N_1760);
or U1871 (N_1871,N_1731,N_1758);
nand U1872 (N_1872,N_1729,N_1774);
or U1873 (N_1873,N_1783,N_1732);
nor U1874 (N_1874,N_1728,N_1776);
nand U1875 (N_1875,N_1848,N_1820);
nand U1876 (N_1876,N_1865,N_1858);
nor U1877 (N_1877,N_1853,N_1839);
nor U1878 (N_1878,N_1857,N_1836);
or U1879 (N_1879,N_1849,N_1822);
nand U1880 (N_1880,N_1870,N_1826);
nand U1881 (N_1881,N_1808,N_1812);
and U1882 (N_1882,N_1827,N_1840);
and U1883 (N_1883,N_1855,N_1809);
and U1884 (N_1884,N_1852,N_1801);
and U1885 (N_1885,N_1872,N_1837);
nand U1886 (N_1886,N_1825,N_1811);
or U1887 (N_1887,N_1819,N_1805);
nor U1888 (N_1888,N_1873,N_1830);
or U1889 (N_1889,N_1844,N_1829);
or U1890 (N_1890,N_1847,N_1868);
and U1891 (N_1891,N_1862,N_1851);
nor U1892 (N_1892,N_1860,N_1859);
nor U1893 (N_1893,N_1835,N_1813);
nand U1894 (N_1894,N_1833,N_1823);
or U1895 (N_1895,N_1864,N_1841);
and U1896 (N_1896,N_1828,N_1856);
and U1897 (N_1897,N_1815,N_1861);
or U1898 (N_1898,N_1817,N_1842);
nand U1899 (N_1899,N_1810,N_1804);
xnor U1900 (N_1900,N_1866,N_1834);
nand U1901 (N_1901,N_1831,N_1838);
or U1902 (N_1902,N_1854,N_1832);
or U1903 (N_1903,N_1807,N_1816);
or U1904 (N_1904,N_1867,N_1818);
or U1905 (N_1905,N_1871,N_1843);
and U1906 (N_1906,N_1800,N_1806);
nor U1907 (N_1907,N_1850,N_1869);
nand U1908 (N_1908,N_1803,N_1846);
xnor U1909 (N_1909,N_1802,N_1845);
nor U1910 (N_1910,N_1863,N_1814);
nand U1911 (N_1911,N_1821,N_1874);
nand U1912 (N_1912,N_1824,N_1823);
nand U1913 (N_1913,N_1810,N_1869);
and U1914 (N_1914,N_1820,N_1851);
nor U1915 (N_1915,N_1815,N_1831);
or U1916 (N_1916,N_1819,N_1828);
or U1917 (N_1917,N_1857,N_1804);
nand U1918 (N_1918,N_1828,N_1822);
and U1919 (N_1919,N_1862,N_1861);
and U1920 (N_1920,N_1817,N_1837);
nand U1921 (N_1921,N_1874,N_1817);
nand U1922 (N_1922,N_1809,N_1815);
or U1923 (N_1923,N_1809,N_1856);
and U1924 (N_1924,N_1859,N_1868);
nor U1925 (N_1925,N_1861,N_1867);
and U1926 (N_1926,N_1845,N_1829);
nor U1927 (N_1927,N_1826,N_1802);
nand U1928 (N_1928,N_1862,N_1839);
nor U1929 (N_1929,N_1822,N_1814);
or U1930 (N_1930,N_1823,N_1853);
nor U1931 (N_1931,N_1870,N_1811);
or U1932 (N_1932,N_1834,N_1839);
nand U1933 (N_1933,N_1843,N_1831);
or U1934 (N_1934,N_1824,N_1857);
and U1935 (N_1935,N_1805,N_1846);
nand U1936 (N_1936,N_1808,N_1827);
nor U1937 (N_1937,N_1841,N_1843);
or U1938 (N_1938,N_1803,N_1840);
or U1939 (N_1939,N_1830,N_1817);
nand U1940 (N_1940,N_1827,N_1871);
nand U1941 (N_1941,N_1865,N_1857);
or U1942 (N_1942,N_1861,N_1851);
and U1943 (N_1943,N_1847,N_1859);
or U1944 (N_1944,N_1864,N_1867);
or U1945 (N_1945,N_1817,N_1855);
nor U1946 (N_1946,N_1810,N_1818);
and U1947 (N_1947,N_1828,N_1857);
nand U1948 (N_1948,N_1800,N_1853);
or U1949 (N_1949,N_1837,N_1830);
and U1950 (N_1950,N_1906,N_1903);
or U1951 (N_1951,N_1905,N_1902);
nand U1952 (N_1952,N_1895,N_1892);
and U1953 (N_1953,N_1916,N_1884);
nand U1954 (N_1954,N_1891,N_1918);
or U1955 (N_1955,N_1940,N_1936);
nand U1956 (N_1956,N_1943,N_1927);
nor U1957 (N_1957,N_1946,N_1901);
nand U1958 (N_1958,N_1882,N_1947);
nand U1959 (N_1959,N_1937,N_1910);
or U1960 (N_1960,N_1928,N_1899);
and U1961 (N_1961,N_1939,N_1877);
nand U1962 (N_1962,N_1923,N_1883);
and U1963 (N_1963,N_1889,N_1885);
and U1964 (N_1964,N_1887,N_1890);
nand U1965 (N_1965,N_1912,N_1933);
nor U1966 (N_1966,N_1908,N_1907);
or U1967 (N_1967,N_1878,N_1888);
nand U1968 (N_1968,N_1876,N_1917);
nor U1969 (N_1969,N_1909,N_1926);
nand U1970 (N_1970,N_1904,N_1935);
nor U1971 (N_1971,N_1886,N_1949);
nor U1972 (N_1972,N_1893,N_1919);
and U1973 (N_1973,N_1932,N_1948);
nand U1974 (N_1974,N_1911,N_1929);
or U1975 (N_1975,N_1898,N_1925);
nor U1976 (N_1976,N_1875,N_1914);
nand U1977 (N_1977,N_1930,N_1945);
nor U1978 (N_1978,N_1900,N_1880);
nor U1979 (N_1979,N_1915,N_1897);
nand U1980 (N_1980,N_1921,N_1944);
and U1981 (N_1981,N_1894,N_1913);
nand U1982 (N_1982,N_1924,N_1934);
nor U1983 (N_1983,N_1896,N_1881);
and U1984 (N_1984,N_1941,N_1922);
nand U1985 (N_1985,N_1938,N_1920);
xor U1986 (N_1986,N_1942,N_1931);
nand U1987 (N_1987,N_1879,N_1918);
or U1988 (N_1988,N_1946,N_1926);
nand U1989 (N_1989,N_1919,N_1902);
and U1990 (N_1990,N_1929,N_1943);
nand U1991 (N_1991,N_1929,N_1897);
nor U1992 (N_1992,N_1923,N_1891);
and U1993 (N_1993,N_1917,N_1948);
or U1994 (N_1994,N_1903,N_1895);
and U1995 (N_1995,N_1889,N_1883);
nor U1996 (N_1996,N_1890,N_1908);
and U1997 (N_1997,N_1934,N_1939);
nand U1998 (N_1998,N_1936,N_1939);
nand U1999 (N_1999,N_1917,N_1931);
or U2000 (N_2000,N_1887,N_1936);
nor U2001 (N_2001,N_1929,N_1938);
and U2002 (N_2002,N_1878,N_1876);
nand U2003 (N_2003,N_1928,N_1875);
or U2004 (N_2004,N_1893,N_1884);
and U2005 (N_2005,N_1906,N_1881);
nor U2006 (N_2006,N_1919,N_1946);
nand U2007 (N_2007,N_1891,N_1931);
nand U2008 (N_2008,N_1917,N_1940);
and U2009 (N_2009,N_1915,N_1932);
nor U2010 (N_2010,N_1887,N_1944);
xor U2011 (N_2011,N_1932,N_1947);
or U2012 (N_2012,N_1900,N_1915);
nor U2013 (N_2013,N_1888,N_1931);
nor U2014 (N_2014,N_1935,N_1934);
nand U2015 (N_2015,N_1920,N_1948);
or U2016 (N_2016,N_1894,N_1882);
nand U2017 (N_2017,N_1914,N_1908);
nor U2018 (N_2018,N_1885,N_1895);
and U2019 (N_2019,N_1942,N_1937);
and U2020 (N_2020,N_1915,N_1939);
and U2021 (N_2021,N_1908,N_1885);
and U2022 (N_2022,N_1876,N_1899);
nand U2023 (N_2023,N_1878,N_1880);
nand U2024 (N_2024,N_1930,N_1929);
nor U2025 (N_2025,N_1972,N_1978);
nand U2026 (N_2026,N_2023,N_2010);
nand U2027 (N_2027,N_2018,N_1994);
or U2028 (N_2028,N_1986,N_2005);
nor U2029 (N_2029,N_1997,N_1951);
and U2030 (N_2030,N_1981,N_1950);
nand U2031 (N_2031,N_2009,N_1984);
nor U2032 (N_2032,N_2011,N_1969);
or U2033 (N_2033,N_1957,N_1955);
nand U2034 (N_2034,N_1976,N_1971);
nor U2035 (N_2035,N_1979,N_1974);
or U2036 (N_2036,N_1996,N_1980);
and U2037 (N_2037,N_1985,N_2022);
or U2038 (N_2038,N_1988,N_1973);
and U2039 (N_2039,N_2002,N_1991);
nand U2040 (N_2040,N_2007,N_1968);
nor U2041 (N_2041,N_1983,N_2012);
and U2042 (N_2042,N_2016,N_1982);
nand U2043 (N_2043,N_1961,N_2017);
and U2044 (N_2044,N_1975,N_1959);
nand U2045 (N_2045,N_1995,N_1966);
nor U2046 (N_2046,N_2003,N_1989);
and U2047 (N_2047,N_1954,N_2019);
or U2048 (N_2048,N_1953,N_2020);
nand U2049 (N_2049,N_2014,N_1999);
nor U2050 (N_2050,N_2013,N_2015);
and U2051 (N_2051,N_2006,N_1970);
nand U2052 (N_2052,N_2008,N_1963);
nor U2053 (N_2053,N_1962,N_2021);
nor U2054 (N_2054,N_1993,N_1967);
and U2055 (N_2055,N_2004,N_1960);
nor U2056 (N_2056,N_1965,N_1952);
and U2057 (N_2057,N_2001,N_2024);
or U2058 (N_2058,N_1990,N_1964);
and U2059 (N_2059,N_1958,N_2000);
or U2060 (N_2060,N_1977,N_1987);
nand U2061 (N_2061,N_1998,N_1992);
nand U2062 (N_2062,N_1956,N_2013);
or U2063 (N_2063,N_2003,N_2012);
nand U2064 (N_2064,N_1971,N_2016);
nor U2065 (N_2065,N_2016,N_1996);
nor U2066 (N_2066,N_1999,N_1997);
nand U2067 (N_2067,N_1990,N_1956);
and U2068 (N_2068,N_2009,N_1989);
and U2069 (N_2069,N_1999,N_1979);
and U2070 (N_2070,N_1999,N_2008);
nor U2071 (N_2071,N_1964,N_2003);
nor U2072 (N_2072,N_1954,N_1998);
or U2073 (N_2073,N_1954,N_1952);
nand U2074 (N_2074,N_2006,N_2001);
nand U2075 (N_2075,N_2018,N_1984);
or U2076 (N_2076,N_2022,N_2011);
nor U2077 (N_2077,N_2015,N_1996);
and U2078 (N_2078,N_1966,N_1999);
nand U2079 (N_2079,N_2014,N_1981);
or U2080 (N_2080,N_1976,N_1985);
nor U2081 (N_2081,N_1957,N_2013);
nand U2082 (N_2082,N_1957,N_2011);
nor U2083 (N_2083,N_1952,N_1992);
and U2084 (N_2084,N_1972,N_1983);
and U2085 (N_2085,N_2016,N_2008);
nand U2086 (N_2086,N_2010,N_1977);
nor U2087 (N_2087,N_1966,N_1984);
or U2088 (N_2088,N_2000,N_2015);
nor U2089 (N_2089,N_1974,N_1966);
and U2090 (N_2090,N_1950,N_1985);
or U2091 (N_2091,N_1996,N_2021);
xor U2092 (N_2092,N_1977,N_2006);
nor U2093 (N_2093,N_1994,N_1970);
and U2094 (N_2094,N_1987,N_1999);
nand U2095 (N_2095,N_1955,N_1981);
nor U2096 (N_2096,N_1997,N_1976);
or U2097 (N_2097,N_1975,N_1971);
or U2098 (N_2098,N_2004,N_1971);
or U2099 (N_2099,N_2024,N_1986);
nand U2100 (N_2100,N_2096,N_2085);
and U2101 (N_2101,N_2088,N_2097);
nand U2102 (N_2102,N_2094,N_2061);
or U2103 (N_2103,N_2033,N_2048);
and U2104 (N_2104,N_2038,N_2071);
or U2105 (N_2105,N_2090,N_2078);
nand U2106 (N_2106,N_2058,N_2084);
nor U2107 (N_2107,N_2077,N_2079);
or U2108 (N_2108,N_2083,N_2070);
and U2109 (N_2109,N_2028,N_2076);
nand U2110 (N_2110,N_2030,N_2045);
nand U2111 (N_2111,N_2093,N_2054);
nor U2112 (N_2112,N_2036,N_2064);
nor U2113 (N_2113,N_2050,N_2043);
nand U2114 (N_2114,N_2067,N_2053);
nor U2115 (N_2115,N_2042,N_2060);
or U2116 (N_2116,N_2072,N_2086);
or U2117 (N_2117,N_2098,N_2069);
nand U2118 (N_2118,N_2035,N_2052);
or U2119 (N_2119,N_2095,N_2046);
nor U2120 (N_2120,N_2074,N_2037);
or U2121 (N_2121,N_2027,N_2025);
nand U2122 (N_2122,N_2032,N_2041);
nor U2123 (N_2123,N_2082,N_2091);
nand U2124 (N_2124,N_2092,N_2065);
nor U2125 (N_2125,N_2044,N_2073);
or U2126 (N_2126,N_2081,N_2087);
nand U2127 (N_2127,N_2099,N_2059);
nand U2128 (N_2128,N_2080,N_2051);
nor U2129 (N_2129,N_2040,N_2075);
nand U2130 (N_2130,N_2057,N_2047);
and U2131 (N_2131,N_2031,N_2089);
nor U2132 (N_2132,N_2056,N_2066);
nor U2133 (N_2133,N_2049,N_2063);
and U2134 (N_2134,N_2068,N_2055);
and U2135 (N_2135,N_2034,N_2029);
nand U2136 (N_2136,N_2039,N_2062);
nor U2137 (N_2137,N_2026,N_2025);
or U2138 (N_2138,N_2035,N_2058);
and U2139 (N_2139,N_2027,N_2030);
and U2140 (N_2140,N_2044,N_2047);
nand U2141 (N_2141,N_2057,N_2050);
nor U2142 (N_2142,N_2064,N_2035);
or U2143 (N_2143,N_2065,N_2032);
nor U2144 (N_2144,N_2028,N_2060);
and U2145 (N_2145,N_2026,N_2031);
or U2146 (N_2146,N_2028,N_2049);
or U2147 (N_2147,N_2044,N_2089);
or U2148 (N_2148,N_2063,N_2055);
or U2149 (N_2149,N_2088,N_2087);
nor U2150 (N_2150,N_2058,N_2065);
or U2151 (N_2151,N_2066,N_2091);
nand U2152 (N_2152,N_2049,N_2026);
nor U2153 (N_2153,N_2026,N_2050);
or U2154 (N_2154,N_2086,N_2043);
and U2155 (N_2155,N_2029,N_2070);
nor U2156 (N_2156,N_2083,N_2080);
or U2157 (N_2157,N_2058,N_2043);
and U2158 (N_2158,N_2049,N_2094);
nor U2159 (N_2159,N_2062,N_2092);
and U2160 (N_2160,N_2094,N_2075);
and U2161 (N_2161,N_2047,N_2089);
and U2162 (N_2162,N_2093,N_2036);
and U2163 (N_2163,N_2087,N_2085);
or U2164 (N_2164,N_2068,N_2033);
or U2165 (N_2165,N_2065,N_2059);
nor U2166 (N_2166,N_2089,N_2050);
and U2167 (N_2167,N_2096,N_2060);
nor U2168 (N_2168,N_2052,N_2069);
and U2169 (N_2169,N_2039,N_2045);
nand U2170 (N_2170,N_2031,N_2095);
and U2171 (N_2171,N_2093,N_2087);
or U2172 (N_2172,N_2027,N_2064);
and U2173 (N_2173,N_2027,N_2038);
nor U2174 (N_2174,N_2074,N_2032);
nor U2175 (N_2175,N_2131,N_2133);
or U2176 (N_2176,N_2143,N_2107);
and U2177 (N_2177,N_2158,N_2164);
nor U2178 (N_2178,N_2118,N_2111);
or U2179 (N_2179,N_2152,N_2105);
or U2180 (N_2180,N_2130,N_2135);
nor U2181 (N_2181,N_2153,N_2117);
or U2182 (N_2182,N_2144,N_2171);
or U2183 (N_2183,N_2160,N_2110);
nor U2184 (N_2184,N_2157,N_2121);
and U2185 (N_2185,N_2104,N_2101);
and U2186 (N_2186,N_2162,N_2113);
nand U2187 (N_2187,N_2169,N_2165);
xor U2188 (N_2188,N_2102,N_2142);
and U2189 (N_2189,N_2108,N_2167);
and U2190 (N_2190,N_2172,N_2174);
nand U2191 (N_2191,N_2170,N_2151);
or U2192 (N_2192,N_2129,N_2137);
and U2193 (N_2193,N_2138,N_2125);
and U2194 (N_2194,N_2128,N_2140);
nand U2195 (N_2195,N_2155,N_2148);
or U2196 (N_2196,N_2159,N_2136);
nor U2197 (N_2197,N_2161,N_2163);
nor U2198 (N_2198,N_2147,N_2122);
or U2199 (N_2199,N_2132,N_2154);
nand U2200 (N_2200,N_2103,N_2106);
nand U2201 (N_2201,N_2123,N_2173);
or U2202 (N_2202,N_2109,N_2100);
and U2203 (N_2203,N_2119,N_2115);
nor U2204 (N_2204,N_2146,N_2141);
and U2205 (N_2205,N_2116,N_2139);
and U2206 (N_2206,N_2134,N_2114);
nand U2207 (N_2207,N_2120,N_2168);
nand U2208 (N_2208,N_2156,N_2150);
nand U2209 (N_2209,N_2112,N_2126);
and U2210 (N_2210,N_2124,N_2145);
and U2211 (N_2211,N_2127,N_2149);
and U2212 (N_2212,N_2166,N_2133);
or U2213 (N_2213,N_2150,N_2109);
and U2214 (N_2214,N_2164,N_2139);
nand U2215 (N_2215,N_2154,N_2146);
nand U2216 (N_2216,N_2120,N_2154);
nand U2217 (N_2217,N_2154,N_2112);
or U2218 (N_2218,N_2115,N_2107);
nand U2219 (N_2219,N_2113,N_2161);
nand U2220 (N_2220,N_2103,N_2148);
nor U2221 (N_2221,N_2136,N_2140);
nand U2222 (N_2222,N_2109,N_2115);
and U2223 (N_2223,N_2117,N_2151);
or U2224 (N_2224,N_2162,N_2167);
nor U2225 (N_2225,N_2153,N_2106);
nand U2226 (N_2226,N_2104,N_2154);
or U2227 (N_2227,N_2157,N_2126);
nand U2228 (N_2228,N_2156,N_2168);
nor U2229 (N_2229,N_2122,N_2145);
nor U2230 (N_2230,N_2105,N_2158);
nor U2231 (N_2231,N_2165,N_2153);
or U2232 (N_2232,N_2156,N_2115);
nand U2233 (N_2233,N_2143,N_2132);
or U2234 (N_2234,N_2160,N_2139);
nor U2235 (N_2235,N_2128,N_2124);
or U2236 (N_2236,N_2115,N_2111);
and U2237 (N_2237,N_2127,N_2160);
nand U2238 (N_2238,N_2109,N_2154);
nor U2239 (N_2239,N_2167,N_2107);
nand U2240 (N_2240,N_2106,N_2165);
or U2241 (N_2241,N_2128,N_2159);
nand U2242 (N_2242,N_2171,N_2136);
or U2243 (N_2243,N_2161,N_2150);
and U2244 (N_2244,N_2167,N_2165);
and U2245 (N_2245,N_2159,N_2137);
nor U2246 (N_2246,N_2145,N_2100);
and U2247 (N_2247,N_2105,N_2119);
and U2248 (N_2248,N_2156,N_2131);
nand U2249 (N_2249,N_2117,N_2128);
nand U2250 (N_2250,N_2211,N_2224);
nand U2251 (N_2251,N_2241,N_2185);
and U2252 (N_2252,N_2226,N_2231);
and U2253 (N_2253,N_2215,N_2229);
nand U2254 (N_2254,N_2225,N_2187);
or U2255 (N_2255,N_2216,N_2210);
or U2256 (N_2256,N_2236,N_2181);
nor U2257 (N_2257,N_2192,N_2218);
or U2258 (N_2258,N_2177,N_2244);
or U2259 (N_2259,N_2238,N_2197);
and U2260 (N_2260,N_2249,N_2203);
and U2261 (N_2261,N_2220,N_2184);
nor U2262 (N_2262,N_2230,N_2235);
nand U2263 (N_2263,N_2195,N_2199);
and U2264 (N_2264,N_2222,N_2182);
or U2265 (N_2265,N_2239,N_2204);
or U2266 (N_2266,N_2189,N_2196);
and U2267 (N_2267,N_2246,N_2213);
nor U2268 (N_2268,N_2221,N_2217);
and U2269 (N_2269,N_2242,N_2180);
or U2270 (N_2270,N_2179,N_2223);
nor U2271 (N_2271,N_2191,N_2219);
nand U2272 (N_2272,N_2201,N_2227);
and U2273 (N_2273,N_2186,N_2206);
nor U2274 (N_2274,N_2248,N_2243);
nand U2275 (N_2275,N_2228,N_2247);
nor U2276 (N_2276,N_2234,N_2208);
nand U2277 (N_2277,N_2176,N_2207);
nand U2278 (N_2278,N_2200,N_2205);
or U2279 (N_2279,N_2190,N_2202);
and U2280 (N_2280,N_2237,N_2188);
and U2281 (N_2281,N_2233,N_2175);
and U2282 (N_2282,N_2212,N_2240);
nor U2283 (N_2283,N_2193,N_2214);
nand U2284 (N_2284,N_2232,N_2245);
nand U2285 (N_2285,N_2183,N_2178);
nand U2286 (N_2286,N_2209,N_2198);
and U2287 (N_2287,N_2194,N_2235);
nand U2288 (N_2288,N_2213,N_2183);
nand U2289 (N_2289,N_2208,N_2219);
nor U2290 (N_2290,N_2242,N_2217);
nor U2291 (N_2291,N_2204,N_2225);
nand U2292 (N_2292,N_2181,N_2200);
nor U2293 (N_2293,N_2217,N_2200);
and U2294 (N_2294,N_2244,N_2219);
nor U2295 (N_2295,N_2189,N_2210);
and U2296 (N_2296,N_2175,N_2198);
or U2297 (N_2297,N_2205,N_2178);
nor U2298 (N_2298,N_2212,N_2207);
nand U2299 (N_2299,N_2245,N_2233);
nand U2300 (N_2300,N_2241,N_2195);
or U2301 (N_2301,N_2182,N_2200);
nor U2302 (N_2302,N_2231,N_2238);
nand U2303 (N_2303,N_2248,N_2210);
or U2304 (N_2304,N_2230,N_2222);
or U2305 (N_2305,N_2187,N_2231);
or U2306 (N_2306,N_2230,N_2204);
or U2307 (N_2307,N_2213,N_2210);
or U2308 (N_2308,N_2229,N_2223);
and U2309 (N_2309,N_2247,N_2241);
and U2310 (N_2310,N_2229,N_2205);
and U2311 (N_2311,N_2216,N_2229);
nand U2312 (N_2312,N_2187,N_2232);
nand U2313 (N_2313,N_2248,N_2249);
xnor U2314 (N_2314,N_2181,N_2194);
nand U2315 (N_2315,N_2227,N_2223);
nand U2316 (N_2316,N_2180,N_2220);
or U2317 (N_2317,N_2231,N_2189);
nand U2318 (N_2318,N_2175,N_2193);
or U2319 (N_2319,N_2198,N_2225);
or U2320 (N_2320,N_2241,N_2236);
or U2321 (N_2321,N_2180,N_2231);
nand U2322 (N_2322,N_2245,N_2214);
nand U2323 (N_2323,N_2176,N_2178);
and U2324 (N_2324,N_2240,N_2203);
or U2325 (N_2325,N_2278,N_2304);
and U2326 (N_2326,N_2277,N_2294);
nor U2327 (N_2327,N_2252,N_2300);
nand U2328 (N_2328,N_2314,N_2320);
nor U2329 (N_2329,N_2299,N_2279);
and U2330 (N_2330,N_2290,N_2310);
and U2331 (N_2331,N_2324,N_2266);
and U2332 (N_2332,N_2311,N_2303);
xnor U2333 (N_2333,N_2260,N_2276);
nand U2334 (N_2334,N_2273,N_2254);
nand U2335 (N_2335,N_2307,N_2264);
nor U2336 (N_2336,N_2272,N_2270);
nand U2337 (N_2337,N_2301,N_2262);
nand U2338 (N_2338,N_2287,N_2306);
and U2339 (N_2339,N_2297,N_2323);
nand U2340 (N_2340,N_2282,N_2263);
or U2341 (N_2341,N_2256,N_2308);
and U2342 (N_2342,N_2318,N_2313);
and U2343 (N_2343,N_2316,N_2293);
nor U2344 (N_2344,N_2305,N_2283);
nand U2345 (N_2345,N_2269,N_2261);
nor U2346 (N_2346,N_2275,N_2259);
or U2347 (N_2347,N_2288,N_2255);
nand U2348 (N_2348,N_2284,N_2265);
or U2349 (N_2349,N_2291,N_2285);
or U2350 (N_2350,N_2292,N_2251);
nand U2351 (N_2351,N_2274,N_2253);
nor U2352 (N_2352,N_2312,N_2296);
xor U2353 (N_2353,N_2317,N_2271);
and U2354 (N_2354,N_2280,N_2289);
or U2355 (N_2355,N_2321,N_2302);
nand U2356 (N_2356,N_2281,N_2257);
nor U2357 (N_2357,N_2298,N_2309);
or U2358 (N_2358,N_2268,N_2250);
nor U2359 (N_2359,N_2295,N_2286);
or U2360 (N_2360,N_2319,N_2315);
nand U2361 (N_2361,N_2267,N_2258);
and U2362 (N_2362,N_2322,N_2266);
nor U2363 (N_2363,N_2275,N_2276);
nor U2364 (N_2364,N_2296,N_2270);
or U2365 (N_2365,N_2298,N_2302);
nand U2366 (N_2366,N_2323,N_2278);
nand U2367 (N_2367,N_2272,N_2251);
or U2368 (N_2368,N_2267,N_2314);
and U2369 (N_2369,N_2265,N_2252);
xnor U2370 (N_2370,N_2293,N_2319);
and U2371 (N_2371,N_2257,N_2301);
nor U2372 (N_2372,N_2263,N_2276);
nand U2373 (N_2373,N_2277,N_2311);
and U2374 (N_2374,N_2263,N_2285);
and U2375 (N_2375,N_2274,N_2311);
nor U2376 (N_2376,N_2303,N_2319);
and U2377 (N_2377,N_2312,N_2291);
nand U2378 (N_2378,N_2273,N_2298);
and U2379 (N_2379,N_2311,N_2322);
and U2380 (N_2380,N_2297,N_2286);
nor U2381 (N_2381,N_2323,N_2315);
nor U2382 (N_2382,N_2292,N_2253);
and U2383 (N_2383,N_2266,N_2259);
and U2384 (N_2384,N_2309,N_2260);
or U2385 (N_2385,N_2318,N_2292);
nand U2386 (N_2386,N_2290,N_2315);
or U2387 (N_2387,N_2300,N_2277);
and U2388 (N_2388,N_2322,N_2306);
nor U2389 (N_2389,N_2277,N_2309);
nor U2390 (N_2390,N_2259,N_2311);
and U2391 (N_2391,N_2303,N_2272);
xnor U2392 (N_2392,N_2276,N_2289);
or U2393 (N_2393,N_2293,N_2292);
or U2394 (N_2394,N_2265,N_2288);
or U2395 (N_2395,N_2292,N_2320);
or U2396 (N_2396,N_2250,N_2311);
and U2397 (N_2397,N_2287,N_2293);
or U2398 (N_2398,N_2276,N_2269);
nand U2399 (N_2399,N_2284,N_2262);
nand U2400 (N_2400,N_2339,N_2391);
nand U2401 (N_2401,N_2377,N_2331);
nor U2402 (N_2402,N_2363,N_2342);
xnor U2403 (N_2403,N_2369,N_2373);
nor U2404 (N_2404,N_2336,N_2395);
nor U2405 (N_2405,N_2375,N_2338);
and U2406 (N_2406,N_2359,N_2365);
nand U2407 (N_2407,N_2355,N_2328);
and U2408 (N_2408,N_2352,N_2333);
xnor U2409 (N_2409,N_2362,N_2335);
nor U2410 (N_2410,N_2383,N_2329);
and U2411 (N_2411,N_2364,N_2354);
or U2412 (N_2412,N_2374,N_2337);
nor U2413 (N_2413,N_2393,N_2350);
nand U2414 (N_2414,N_2327,N_2372);
or U2415 (N_2415,N_2399,N_2357);
nor U2416 (N_2416,N_2325,N_2340);
nand U2417 (N_2417,N_2398,N_2386);
nor U2418 (N_2418,N_2351,N_2347);
or U2419 (N_2419,N_2379,N_2349);
and U2420 (N_2420,N_2326,N_2366);
xnor U2421 (N_2421,N_2387,N_2388);
and U2422 (N_2422,N_2384,N_2345);
nor U2423 (N_2423,N_2332,N_2330);
and U2424 (N_2424,N_2346,N_2367);
nand U2425 (N_2425,N_2348,N_2358);
nor U2426 (N_2426,N_2394,N_2397);
and U2427 (N_2427,N_2344,N_2361);
and U2428 (N_2428,N_2390,N_2382);
nand U2429 (N_2429,N_2343,N_2371);
nor U2430 (N_2430,N_2370,N_2380);
and U2431 (N_2431,N_2378,N_2392);
nor U2432 (N_2432,N_2353,N_2385);
nand U2433 (N_2433,N_2396,N_2356);
nor U2434 (N_2434,N_2368,N_2389);
nand U2435 (N_2435,N_2381,N_2341);
and U2436 (N_2436,N_2360,N_2376);
nand U2437 (N_2437,N_2334,N_2349);
nand U2438 (N_2438,N_2353,N_2372);
and U2439 (N_2439,N_2328,N_2383);
and U2440 (N_2440,N_2382,N_2398);
nand U2441 (N_2441,N_2378,N_2385);
nand U2442 (N_2442,N_2331,N_2371);
nand U2443 (N_2443,N_2332,N_2360);
nor U2444 (N_2444,N_2349,N_2374);
and U2445 (N_2445,N_2352,N_2337);
or U2446 (N_2446,N_2349,N_2340);
or U2447 (N_2447,N_2363,N_2360);
nor U2448 (N_2448,N_2398,N_2355);
and U2449 (N_2449,N_2341,N_2368);
xnor U2450 (N_2450,N_2328,N_2326);
nor U2451 (N_2451,N_2348,N_2386);
nor U2452 (N_2452,N_2378,N_2359);
nor U2453 (N_2453,N_2356,N_2393);
nor U2454 (N_2454,N_2370,N_2342);
and U2455 (N_2455,N_2346,N_2375);
and U2456 (N_2456,N_2368,N_2359);
and U2457 (N_2457,N_2338,N_2392);
and U2458 (N_2458,N_2330,N_2370);
or U2459 (N_2459,N_2345,N_2392);
xnor U2460 (N_2460,N_2395,N_2328);
nor U2461 (N_2461,N_2373,N_2365);
and U2462 (N_2462,N_2379,N_2376);
and U2463 (N_2463,N_2368,N_2391);
and U2464 (N_2464,N_2393,N_2380);
nand U2465 (N_2465,N_2370,N_2374);
or U2466 (N_2466,N_2368,N_2352);
nor U2467 (N_2467,N_2347,N_2383);
nand U2468 (N_2468,N_2372,N_2357);
nor U2469 (N_2469,N_2385,N_2377);
nor U2470 (N_2470,N_2376,N_2345);
and U2471 (N_2471,N_2384,N_2382);
xnor U2472 (N_2472,N_2393,N_2383);
nor U2473 (N_2473,N_2387,N_2376);
and U2474 (N_2474,N_2331,N_2380);
nor U2475 (N_2475,N_2440,N_2439);
nand U2476 (N_2476,N_2468,N_2401);
xnor U2477 (N_2477,N_2433,N_2412);
nor U2478 (N_2478,N_2416,N_2428);
nand U2479 (N_2479,N_2406,N_2462);
nand U2480 (N_2480,N_2420,N_2432);
nor U2481 (N_2481,N_2469,N_2441);
or U2482 (N_2482,N_2460,N_2407);
nand U2483 (N_2483,N_2446,N_2471);
nand U2484 (N_2484,N_2431,N_2419);
and U2485 (N_2485,N_2421,N_2413);
and U2486 (N_2486,N_2418,N_2409);
nand U2487 (N_2487,N_2467,N_2404);
and U2488 (N_2488,N_2426,N_2405);
and U2489 (N_2489,N_2455,N_2459);
or U2490 (N_2490,N_2465,N_2402);
xnor U2491 (N_2491,N_2423,N_2451);
nand U2492 (N_2492,N_2422,N_2457);
and U2493 (N_2493,N_2452,N_2415);
and U2494 (N_2494,N_2414,N_2400);
nor U2495 (N_2495,N_2408,N_2466);
nand U2496 (N_2496,N_2464,N_2458);
nor U2497 (N_2497,N_2453,N_2472);
nor U2498 (N_2498,N_2429,N_2430);
or U2499 (N_2499,N_2470,N_2417);
and U2500 (N_2500,N_2463,N_2473);
nor U2501 (N_2501,N_2456,N_2448);
nand U2502 (N_2502,N_2445,N_2403);
nor U2503 (N_2503,N_2435,N_2474);
and U2504 (N_2504,N_2425,N_2442);
nand U2505 (N_2505,N_2443,N_2424);
nor U2506 (N_2506,N_2438,N_2410);
or U2507 (N_2507,N_2434,N_2454);
nand U2508 (N_2508,N_2436,N_2450);
or U2509 (N_2509,N_2427,N_2437);
nand U2510 (N_2510,N_2411,N_2444);
or U2511 (N_2511,N_2461,N_2449);
xor U2512 (N_2512,N_2447,N_2441);
or U2513 (N_2513,N_2438,N_2403);
or U2514 (N_2514,N_2410,N_2427);
nand U2515 (N_2515,N_2458,N_2410);
nand U2516 (N_2516,N_2447,N_2472);
nor U2517 (N_2517,N_2467,N_2468);
nand U2518 (N_2518,N_2415,N_2445);
and U2519 (N_2519,N_2451,N_2409);
nand U2520 (N_2520,N_2462,N_2441);
or U2521 (N_2521,N_2457,N_2458);
and U2522 (N_2522,N_2448,N_2426);
or U2523 (N_2523,N_2466,N_2407);
nand U2524 (N_2524,N_2424,N_2433);
and U2525 (N_2525,N_2419,N_2422);
or U2526 (N_2526,N_2415,N_2473);
and U2527 (N_2527,N_2420,N_2428);
and U2528 (N_2528,N_2460,N_2469);
or U2529 (N_2529,N_2439,N_2441);
xnor U2530 (N_2530,N_2467,N_2412);
nand U2531 (N_2531,N_2432,N_2405);
or U2532 (N_2532,N_2428,N_2413);
or U2533 (N_2533,N_2469,N_2458);
or U2534 (N_2534,N_2414,N_2423);
or U2535 (N_2535,N_2453,N_2410);
nand U2536 (N_2536,N_2438,N_2413);
and U2537 (N_2537,N_2470,N_2469);
or U2538 (N_2538,N_2432,N_2401);
or U2539 (N_2539,N_2438,N_2400);
nor U2540 (N_2540,N_2409,N_2404);
and U2541 (N_2541,N_2462,N_2472);
or U2542 (N_2542,N_2405,N_2456);
nand U2543 (N_2543,N_2416,N_2448);
nor U2544 (N_2544,N_2405,N_2419);
or U2545 (N_2545,N_2451,N_2426);
nand U2546 (N_2546,N_2437,N_2435);
nand U2547 (N_2547,N_2436,N_2415);
or U2548 (N_2548,N_2473,N_2439);
nor U2549 (N_2549,N_2423,N_2427);
nand U2550 (N_2550,N_2522,N_2530);
or U2551 (N_2551,N_2524,N_2539);
nor U2552 (N_2552,N_2487,N_2549);
and U2553 (N_2553,N_2493,N_2481);
nor U2554 (N_2554,N_2529,N_2525);
nand U2555 (N_2555,N_2517,N_2528);
nand U2556 (N_2556,N_2509,N_2478);
nor U2557 (N_2557,N_2484,N_2491);
nor U2558 (N_2558,N_2510,N_2486);
nand U2559 (N_2559,N_2523,N_2512);
nand U2560 (N_2560,N_2503,N_2479);
nor U2561 (N_2561,N_2507,N_2489);
nand U2562 (N_2562,N_2496,N_2542);
or U2563 (N_2563,N_2537,N_2521);
and U2564 (N_2564,N_2514,N_2515);
and U2565 (N_2565,N_2520,N_2482);
nand U2566 (N_2566,N_2527,N_2536);
nor U2567 (N_2567,N_2492,N_2504);
and U2568 (N_2568,N_2519,N_2511);
nand U2569 (N_2569,N_2547,N_2495);
nor U2570 (N_2570,N_2480,N_2485);
nand U2571 (N_2571,N_2506,N_2502);
or U2572 (N_2572,N_2490,N_2513);
nor U2573 (N_2573,N_2535,N_2518);
nand U2574 (N_2574,N_2505,N_2488);
and U2575 (N_2575,N_2494,N_2544);
and U2576 (N_2576,N_2498,N_2540);
and U2577 (N_2577,N_2543,N_2534);
or U2578 (N_2578,N_2477,N_2541);
xor U2579 (N_2579,N_2545,N_2531);
nor U2580 (N_2580,N_2516,N_2476);
and U2581 (N_2581,N_2499,N_2501);
and U2582 (N_2582,N_2526,N_2548);
nand U2583 (N_2583,N_2532,N_2533);
nand U2584 (N_2584,N_2508,N_2500);
nand U2585 (N_2585,N_2546,N_2497);
nand U2586 (N_2586,N_2483,N_2538);
and U2587 (N_2587,N_2475,N_2521);
and U2588 (N_2588,N_2525,N_2501);
or U2589 (N_2589,N_2531,N_2528);
nand U2590 (N_2590,N_2483,N_2521);
nor U2591 (N_2591,N_2486,N_2547);
nor U2592 (N_2592,N_2520,N_2511);
nand U2593 (N_2593,N_2484,N_2532);
nand U2594 (N_2594,N_2536,N_2499);
nand U2595 (N_2595,N_2486,N_2525);
nor U2596 (N_2596,N_2499,N_2502);
or U2597 (N_2597,N_2512,N_2521);
nand U2598 (N_2598,N_2483,N_2531);
or U2599 (N_2599,N_2501,N_2507);
nor U2600 (N_2600,N_2533,N_2539);
and U2601 (N_2601,N_2531,N_2484);
nand U2602 (N_2602,N_2547,N_2483);
or U2603 (N_2603,N_2512,N_2506);
and U2604 (N_2604,N_2485,N_2521);
nand U2605 (N_2605,N_2498,N_2486);
and U2606 (N_2606,N_2502,N_2526);
nand U2607 (N_2607,N_2496,N_2523);
nor U2608 (N_2608,N_2520,N_2507);
nand U2609 (N_2609,N_2502,N_2519);
or U2610 (N_2610,N_2479,N_2514);
nor U2611 (N_2611,N_2477,N_2489);
or U2612 (N_2612,N_2475,N_2501);
or U2613 (N_2613,N_2520,N_2542);
and U2614 (N_2614,N_2498,N_2491);
and U2615 (N_2615,N_2484,N_2523);
nor U2616 (N_2616,N_2519,N_2499);
or U2617 (N_2617,N_2508,N_2491);
nand U2618 (N_2618,N_2502,N_2478);
nor U2619 (N_2619,N_2528,N_2518);
or U2620 (N_2620,N_2478,N_2491);
nand U2621 (N_2621,N_2522,N_2504);
or U2622 (N_2622,N_2546,N_2502);
or U2623 (N_2623,N_2497,N_2500);
and U2624 (N_2624,N_2534,N_2477);
nand U2625 (N_2625,N_2556,N_2588);
nand U2626 (N_2626,N_2598,N_2604);
or U2627 (N_2627,N_2596,N_2622);
xor U2628 (N_2628,N_2565,N_2583);
or U2629 (N_2629,N_2559,N_2582);
and U2630 (N_2630,N_2602,N_2555);
and U2631 (N_2631,N_2561,N_2608);
nand U2632 (N_2632,N_2550,N_2558);
or U2633 (N_2633,N_2621,N_2593);
or U2634 (N_2634,N_2616,N_2610);
nor U2635 (N_2635,N_2562,N_2568);
nand U2636 (N_2636,N_2574,N_2599);
nand U2637 (N_2637,N_2603,N_2609);
or U2638 (N_2638,N_2612,N_2611);
and U2639 (N_2639,N_2569,N_2578);
or U2640 (N_2640,N_2560,N_2551);
nor U2641 (N_2641,N_2586,N_2619);
and U2642 (N_2642,N_2600,N_2595);
and U2643 (N_2643,N_2594,N_2591);
and U2644 (N_2644,N_2575,N_2614);
nor U2645 (N_2645,N_2570,N_2607);
or U2646 (N_2646,N_2587,N_2572);
and U2647 (N_2647,N_2557,N_2564);
and U2648 (N_2648,N_2601,N_2605);
nand U2649 (N_2649,N_2590,N_2554);
and U2650 (N_2650,N_2624,N_2566);
and U2651 (N_2651,N_2597,N_2585);
or U2652 (N_2652,N_2563,N_2620);
nor U2653 (N_2653,N_2573,N_2615);
nor U2654 (N_2654,N_2553,N_2581);
nand U2655 (N_2655,N_2567,N_2577);
and U2656 (N_2656,N_2606,N_2623);
and U2657 (N_2657,N_2618,N_2617);
or U2658 (N_2658,N_2580,N_2576);
xor U2659 (N_2659,N_2592,N_2589);
xnor U2660 (N_2660,N_2571,N_2552);
nor U2661 (N_2661,N_2584,N_2579);
nand U2662 (N_2662,N_2613,N_2559);
nor U2663 (N_2663,N_2580,N_2562);
nor U2664 (N_2664,N_2620,N_2583);
nor U2665 (N_2665,N_2591,N_2580);
and U2666 (N_2666,N_2601,N_2598);
or U2667 (N_2667,N_2621,N_2552);
and U2668 (N_2668,N_2566,N_2552);
and U2669 (N_2669,N_2573,N_2568);
and U2670 (N_2670,N_2604,N_2557);
or U2671 (N_2671,N_2589,N_2571);
nand U2672 (N_2672,N_2622,N_2588);
and U2673 (N_2673,N_2578,N_2579);
nor U2674 (N_2674,N_2594,N_2550);
or U2675 (N_2675,N_2601,N_2603);
nor U2676 (N_2676,N_2616,N_2588);
nand U2677 (N_2677,N_2594,N_2621);
or U2678 (N_2678,N_2555,N_2580);
nor U2679 (N_2679,N_2563,N_2589);
or U2680 (N_2680,N_2572,N_2605);
and U2681 (N_2681,N_2603,N_2556);
xnor U2682 (N_2682,N_2615,N_2569);
and U2683 (N_2683,N_2599,N_2561);
nand U2684 (N_2684,N_2604,N_2555);
and U2685 (N_2685,N_2598,N_2619);
nand U2686 (N_2686,N_2592,N_2555);
nand U2687 (N_2687,N_2559,N_2568);
nor U2688 (N_2688,N_2581,N_2584);
or U2689 (N_2689,N_2571,N_2586);
or U2690 (N_2690,N_2588,N_2601);
and U2691 (N_2691,N_2617,N_2576);
or U2692 (N_2692,N_2601,N_2624);
nor U2693 (N_2693,N_2551,N_2603);
nand U2694 (N_2694,N_2574,N_2569);
or U2695 (N_2695,N_2562,N_2617);
nand U2696 (N_2696,N_2590,N_2583);
and U2697 (N_2697,N_2570,N_2579);
and U2698 (N_2698,N_2558,N_2570);
nor U2699 (N_2699,N_2585,N_2550);
nor U2700 (N_2700,N_2632,N_2672);
xnor U2701 (N_2701,N_2650,N_2691);
and U2702 (N_2702,N_2629,N_2639);
and U2703 (N_2703,N_2670,N_2685);
nand U2704 (N_2704,N_2643,N_2654);
and U2705 (N_2705,N_2641,N_2687);
nand U2706 (N_2706,N_2686,N_2625);
nor U2707 (N_2707,N_2692,N_2675);
xnor U2708 (N_2708,N_2626,N_2667);
nand U2709 (N_2709,N_2668,N_2659);
nor U2710 (N_2710,N_2658,N_2642);
and U2711 (N_2711,N_2634,N_2682);
nand U2712 (N_2712,N_2655,N_2663);
or U2713 (N_2713,N_2628,N_2681);
nand U2714 (N_2714,N_2673,N_2679);
and U2715 (N_2715,N_2683,N_2678);
nand U2716 (N_2716,N_2677,N_2631);
nor U2717 (N_2717,N_2669,N_2693);
nor U2718 (N_2718,N_2697,N_2660);
and U2719 (N_2719,N_2696,N_2637);
nor U2720 (N_2720,N_2690,N_2636);
nand U2721 (N_2721,N_2646,N_2651);
nor U2722 (N_2722,N_2680,N_2627);
or U2723 (N_2723,N_2666,N_2688);
nor U2724 (N_2724,N_2694,N_2676);
nor U2725 (N_2725,N_2698,N_2657);
and U2726 (N_2726,N_2664,N_2662);
nor U2727 (N_2727,N_2665,N_2638);
nand U2728 (N_2728,N_2649,N_2671);
nand U2729 (N_2729,N_2633,N_2699);
nand U2730 (N_2730,N_2674,N_2640);
nand U2731 (N_2731,N_2635,N_2684);
nor U2732 (N_2732,N_2653,N_2644);
nand U2733 (N_2733,N_2645,N_2695);
nor U2734 (N_2734,N_2656,N_2652);
nor U2735 (N_2735,N_2689,N_2647);
nand U2736 (N_2736,N_2630,N_2661);
nand U2737 (N_2737,N_2648,N_2660);
nor U2738 (N_2738,N_2675,N_2681);
and U2739 (N_2739,N_2662,N_2653);
nand U2740 (N_2740,N_2643,N_2677);
nand U2741 (N_2741,N_2646,N_2664);
nor U2742 (N_2742,N_2698,N_2677);
and U2743 (N_2743,N_2650,N_2695);
or U2744 (N_2744,N_2693,N_2625);
nor U2745 (N_2745,N_2645,N_2662);
or U2746 (N_2746,N_2633,N_2649);
or U2747 (N_2747,N_2627,N_2698);
or U2748 (N_2748,N_2687,N_2640);
and U2749 (N_2749,N_2644,N_2678);
and U2750 (N_2750,N_2691,N_2666);
and U2751 (N_2751,N_2691,N_2631);
and U2752 (N_2752,N_2632,N_2666);
and U2753 (N_2753,N_2690,N_2680);
and U2754 (N_2754,N_2682,N_2630);
or U2755 (N_2755,N_2654,N_2626);
and U2756 (N_2756,N_2629,N_2671);
or U2757 (N_2757,N_2645,N_2631);
nand U2758 (N_2758,N_2677,N_2671);
or U2759 (N_2759,N_2657,N_2638);
nor U2760 (N_2760,N_2689,N_2665);
or U2761 (N_2761,N_2668,N_2698);
and U2762 (N_2762,N_2632,N_2631);
or U2763 (N_2763,N_2681,N_2699);
or U2764 (N_2764,N_2668,N_2636);
or U2765 (N_2765,N_2660,N_2654);
and U2766 (N_2766,N_2640,N_2663);
or U2767 (N_2767,N_2650,N_2688);
nor U2768 (N_2768,N_2653,N_2691);
nor U2769 (N_2769,N_2657,N_2655);
nand U2770 (N_2770,N_2628,N_2644);
and U2771 (N_2771,N_2696,N_2629);
nand U2772 (N_2772,N_2652,N_2678);
or U2773 (N_2773,N_2687,N_2674);
nand U2774 (N_2774,N_2679,N_2699);
or U2775 (N_2775,N_2751,N_2703);
and U2776 (N_2776,N_2748,N_2735);
nand U2777 (N_2777,N_2759,N_2730);
or U2778 (N_2778,N_2734,N_2701);
nand U2779 (N_2779,N_2756,N_2757);
or U2780 (N_2780,N_2749,N_2768);
nor U2781 (N_2781,N_2740,N_2736);
and U2782 (N_2782,N_2764,N_2720);
nor U2783 (N_2783,N_2743,N_2726);
nor U2784 (N_2784,N_2754,N_2700);
nor U2785 (N_2785,N_2772,N_2760);
or U2786 (N_2786,N_2728,N_2761);
and U2787 (N_2787,N_2707,N_2729);
nand U2788 (N_2788,N_2765,N_2774);
or U2789 (N_2789,N_2706,N_2709);
and U2790 (N_2790,N_2771,N_2752);
nand U2791 (N_2791,N_2763,N_2705);
and U2792 (N_2792,N_2741,N_2731);
nand U2793 (N_2793,N_2702,N_2715);
nor U2794 (N_2794,N_2717,N_2739);
or U2795 (N_2795,N_2737,N_2744);
nand U2796 (N_2796,N_2745,N_2714);
nor U2797 (N_2797,N_2753,N_2710);
or U2798 (N_2798,N_2773,N_2723);
nand U2799 (N_2799,N_2758,N_2755);
nand U2800 (N_2800,N_2767,N_2732);
nand U2801 (N_2801,N_2769,N_2738);
nand U2802 (N_2802,N_2750,N_2722);
nand U2803 (N_2803,N_2704,N_2746);
nor U2804 (N_2804,N_2708,N_2711);
nor U2805 (N_2805,N_2718,N_2716);
nor U2806 (N_2806,N_2770,N_2733);
or U2807 (N_2807,N_2727,N_2762);
and U2808 (N_2808,N_2713,N_2719);
nor U2809 (N_2809,N_2724,N_2712);
or U2810 (N_2810,N_2725,N_2742);
nand U2811 (N_2811,N_2766,N_2747);
nor U2812 (N_2812,N_2721,N_2728);
and U2813 (N_2813,N_2711,N_2712);
nand U2814 (N_2814,N_2752,N_2743);
nor U2815 (N_2815,N_2774,N_2719);
or U2816 (N_2816,N_2755,N_2726);
nand U2817 (N_2817,N_2724,N_2750);
nor U2818 (N_2818,N_2733,N_2764);
or U2819 (N_2819,N_2736,N_2731);
and U2820 (N_2820,N_2768,N_2750);
nand U2821 (N_2821,N_2705,N_2702);
nand U2822 (N_2822,N_2711,N_2709);
nand U2823 (N_2823,N_2706,N_2714);
nor U2824 (N_2824,N_2756,N_2705);
and U2825 (N_2825,N_2718,N_2721);
nand U2826 (N_2826,N_2763,N_2749);
and U2827 (N_2827,N_2761,N_2707);
or U2828 (N_2828,N_2724,N_2755);
and U2829 (N_2829,N_2766,N_2736);
and U2830 (N_2830,N_2724,N_2762);
and U2831 (N_2831,N_2750,N_2749);
or U2832 (N_2832,N_2744,N_2764);
nor U2833 (N_2833,N_2717,N_2741);
xor U2834 (N_2834,N_2710,N_2740);
nor U2835 (N_2835,N_2756,N_2718);
or U2836 (N_2836,N_2767,N_2755);
nor U2837 (N_2837,N_2709,N_2743);
nor U2838 (N_2838,N_2774,N_2747);
nand U2839 (N_2839,N_2720,N_2767);
or U2840 (N_2840,N_2731,N_2754);
or U2841 (N_2841,N_2702,N_2706);
nor U2842 (N_2842,N_2724,N_2758);
or U2843 (N_2843,N_2711,N_2768);
and U2844 (N_2844,N_2765,N_2728);
or U2845 (N_2845,N_2756,N_2752);
nor U2846 (N_2846,N_2716,N_2742);
nor U2847 (N_2847,N_2718,N_2730);
and U2848 (N_2848,N_2746,N_2720);
and U2849 (N_2849,N_2748,N_2725);
nand U2850 (N_2850,N_2819,N_2848);
and U2851 (N_2851,N_2785,N_2792);
and U2852 (N_2852,N_2783,N_2781);
and U2853 (N_2853,N_2817,N_2839);
and U2854 (N_2854,N_2812,N_2809);
nand U2855 (N_2855,N_2811,N_2798);
nor U2856 (N_2856,N_2802,N_2824);
nand U2857 (N_2857,N_2825,N_2830);
nand U2858 (N_2858,N_2820,N_2799);
and U2859 (N_2859,N_2776,N_2804);
xor U2860 (N_2860,N_2784,N_2789);
nor U2861 (N_2861,N_2777,N_2788);
nand U2862 (N_2862,N_2801,N_2842);
and U2863 (N_2863,N_2818,N_2829);
or U2864 (N_2864,N_2833,N_2822);
nor U2865 (N_2865,N_2835,N_2797);
nand U2866 (N_2866,N_2780,N_2836);
or U2867 (N_2867,N_2816,N_2845);
or U2868 (N_2868,N_2807,N_2778);
nand U2869 (N_2869,N_2849,N_2834);
nor U2870 (N_2870,N_2794,N_2841);
or U2871 (N_2871,N_2775,N_2805);
nor U2872 (N_2872,N_2826,N_2828);
nor U2873 (N_2873,N_2844,N_2815);
nor U2874 (N_2874,N_2827,N_2786);
and U2875 (N_2875,N_2813,N_2800);
nand U2876 (N_2876,N_2790,N_2793);
or U2877 (N_2877,N_2791,N_2806);
or U2878 (N_2878,N_2787,N_2803);
nand U2879 (N_2879,N_2846,N_2832);
and U2880 (N_2880,N_2837,N_2810);
nand U2881 (N_2881,N_2814,N_2823);
nor U2882 (N_2882,N_2843,N_2838);
nor U2883 (N_2883,N_2782,N_2795);
and U2884 (N_2884,N_2840,N_2831);
and U2885 (N_2885,N_2821,N_2808);
nand U2886 (N_2886,N_2847,N_2779);
and U2887 (N_2887,N_2796,N_2790);
nor U2888 (N_2888,N_2778,N_2805);
or U2889 (N_2889,N_2777,N_2804);
or U2890 (N_2890,N_2805,N_2801);
or U2891 (N_2891,N_2799,N_2783);
nor U2892 (N_2892,N_2780,N_2809);
or U2893 (N_2893,N_2824,N_2836);
nand U2894 (N_2894,N_2810,N_2814);
and U2895 (N_2895,N_2841,N_2813);
and U2896 (N_2896,N_2783,N_2788);
nor U2897 (N_2897,N_2849,N_2792);
or U2898 (N_2898,N_2788,N_2825);
or U2899 (N_2899,N_2806,N_2829);
nor U2900 (N_2900,N_2848,N_2807);
nand U2901 (N_2901,N_2840,N_2788);
or U2902 (N_2902,N_2783,N_2787);
or U2903 (N_2903,N_2839,N_2814);
or U2904 (N_2904,N_2832,N_2786);
nor U2905 (N_2905,N_2843,N_2805);
nand U2906 (N_2906,N_2793,N_2788);
nand U2907 (N_2907,N_2837,N_2832);
nor U2908 (N_2908,N_2843,N_2777);
nor U2909 (N_2909,N_2843,N_2849);
or U2910 (N_2910,N_2802,N_2799);
or U2911 (N_2911,N_2794,N_2813);
nand U2912 (N_2912,N_2841,N_2844);
nor U2913 (N_2913,N_2812,N_2803);
and U2914 (N_2914,N_2829,N_2781);
or U2915 (N_2915,N_2776,N_2832);
and U2916 (N_2916,N_2803,N_2783);
or U2917 (N_2917,N_2830,N_2808);
or U2918 (N_2918,N_2825,N_2803);
nand U2919 (N_2919,N_2839,N_2778);
or U2920 (N_2920,N_2828,N_2815);
nor U2921 (N_2921,N_2824,N_2826);
nand U2922 (N_2922,N_2802,N_2791);
or U2923 (N_2923,N_2781,N_2809);
nand U2924 (N_2924,N_2811,N_2819);
nor U2925 (N_2925,N_2899,N_2917);
nor U2926 (N_2926,N_2858,N_2904);
and U2927 (N_2927,N_2887,N_2896);
and U2928 (N_2928,N_2876,N_2853);
or U2929 (N_2929,N_2875,N_2923);
nand U2930 (N_2930,N_2878,N_2888);
and U2931 (N_2931,N_2909,N_2901);
or U2932 (N_2932,N_2921,N_2877);
and U2933 (N_2933,N_2869,N_2920);
nor U2934 (N_2934,N_2889,N_2865);
nand U2935 (N_2935,N_2903,N_2908);
or U2936 (N_2936,N_2855,N_2859);
and U2937 (N_2937,N_2857,N_2868);
and U2938 (N_2938,N_2919,N_2883);
or U2939 (N_2939,N_2884,N_2885);
nand U2940 (N_2940,N_2879,N_2914);
nand U2941 (N_2941,N_2852,N_2922);
xnor U2942 (N_2942,N_2910,N_2861);
and U2943 (N_2943,N_2850,N_2912);
or U2944 (N_2944,N_2911,N_2892);
or U2945 (N_2945,N_2866,N_2895);
nand U2946 (N_2946,N_2874,N_2893);
nand U2947 (N_2947,N_2898,N_2906);
nor U2948 (N_2948,N_2905,N_2916);
and U2949 (N_2949,N_2900,N_2907);
nand U2950 (N_2950,N_2856,N_2851);
nand U2951 (N_2951,N_2918,N_2870);
nand U2952 (N_2952,N_2860,N_2891);
nand U2953 (N_2953,N_2881,N_2863);
or U2954 (N_2954,N_2902,N_2872);
nand U2955 (N_2955,N_2867,N_2924);
nand U2956 (N_2956,N_2871,N_2894);
and U2957 (N_2957,N_2854,N_2886);
nor U2958 (N_2958,N_2880,N_2897);
nor U2959 (N_2959,N_2862,N_2873);
or U2960 (N_2960,N_2864,N_2882);
nand U2961 (N_2961,N_2913,N_2890);
and U2962 (N_2962,N_2915,N_2900);
nand U2963 (N_2963,N_2894,N_2851);
nor U2964 (N_2964,N_2856,N_2884);
nand U2965 (N_2965,N_2900,N_2877);
nand U2966 (N_2966,N_2878,N_2889);
and U2967 (N_2967,N_2903,N_2884);
nor U2968 (N_2968,N_2868,N_2850);
nand U2969 (N_2969,N_2857,N_2917);
or U2970 (N_2970,N_2858,N_2884);
nor U2971 (N_2971,N_2857,N_2905);
or U2972 (N_2972,N_2922,N_2893);
nor U2973 (N_2973,N_2888,N_2857);
or U2974 (N_2974,N_2894,N_2896);
and U2975 (N_2975,N_2912,N_2855);
or U2976 (N_2976,N_2920,N_2864);
nand U2977 (N_2977,N_2850,N_2904);
and U2978 (N_2978,N_2858,N_2876);
nor U2979 (N_2979,N_2912,N_2885);
nand U2980 (N_2980,N_2890,N_2860);
or U2981 (N_2981,N_2900,N_2861);
or U2982 (N_2982,N_2862,N_2917);
and U2983 (N_2983,N_2906,N_2900);
nor U2984 (N_2984,N_2882,N_2883);
nand U2985 (N_2985,N_2877,N_2851);
or U2986 (N_2986,N_2870,N_2914);
and U2987 (N_2987,N_2904,N_2851);
nand U2988 (N_2988,N_2911,N_2918);
nand U2989 (N_2989,N_2901,N_2894);
or U2990 (N_2990,N_2898,N_2907);
and U2991 (N_2991,N_2850,N_2885);
nand U2992 (N_2992,N_2861,N_2860);
or U2993 (N_2993,N_2867,N_2850);
or U2994 (N_2994,N_2871,N_2857);
nor U2995 (N_2995,N_2914,N_2888);
or U2996 (N_2996,N_2903,N_2866);
nand U2997 (N_2997,N_2923,N_2913);
nor U2998 (N_2998,N_2901,N_2850);
nor U2999 (N_2999,N_2857,N_2906);
and UO_0 (O_0,N_2987,N_2961);
nor UO_1 (O_1,N_2998,N_2954);
or UO_2 (O_2,N_2973,N_2943);
nor UO_3 (O_3,N_2926,N_2934);
nor UO_4 (O_4,N_2980,N_2938);
and UO_5 (O_5,N_2992,N_2999);
nand UO_6 (O_6,N_2931,N_2988);
or UO_7 (O_7,N_2997,N_2994);
and UO_8 (O_8,N_2978,N_2964);
or UO_9 (O_9,N_2953,N_2963);
or UO_10 (O_10,N_2936,N_2945);
nor UO_11 (O_11,N_2927,N_2925);
nor UO_12 (O_12,N_2983,N_2949);
nand UO_13 (O_13,N_2944,N_2939);
nor UO_14 (O_14,N_2941,N_2962);
or UO_15 (O_15,N_2975,N_2946);
nand UO_16 (O_16,N_2929,N_2981);
nand UO_17 (O_17,N_2977,N_2976);
nor UO_18 (O_18,N_2955,N_2935);
or UO_19 (O_19,N_2948,N_2947);
and UO_20 (O_20,N_2989,N_2979);
and UO_21 (O_21,N_2942,N_2986);
nand UO_22 (O_22,N_2951,N_2937);
nor UO_23 (O_23,N_2996,N_2940);
nand UO_24 (O_24,N_2985,N_2969);
nand UO_25 (O_25,N_2991,N_2984);
or UO_26 (O_26,N_2932,N_2982);
or UO_27 (O_27,N_2968,N_2958);
or UO_28 (O_28,N_2957,N_2966);
nor UO_29 (O_29,N_2965,N_2930);
or UO_30 (O_30,N_2928,N_2933);
nand UO_31 (O_31,N_2990,N_2995);
or UO_32 (O_32,N_2971,N_2952);
nor UO_33 (O_33,N_2974,N_2993);
and UO_34 (O_34,N_2950,N_2967);
and UO_35 (O_35,N_2970,N_2972);
nor UO_36 (O_36,N_2959,N_2956);
and UO_37 (O_37,N_2960,N_2963);
and UO_38 (O_38,N_2936,N_2976);
or UO_39 (O_39,N_2930,N_2976);
and UO_40 (O_40,N_2955,N_2930);
nand UO_41 (O_41,N_2989,N_2988);
nand UO_42 (O_42,N_2940,N_2957);
nor UO_43 (O_43,N_2933,N_2992);
nor UO_44 (O_44,N_2942,N_2984);
and UO_45 (O_45,N_2969,N_2992);
nor UO_46 (O_46,N_2990,N_2931);
and UO_47 (O_47,N_2952,N_2990);
or UO_48 (O_48,N_2949,N_2937);
and UO_49 (O_49,N_2945,N_2942);
or UO_50 (O_50,N_2999,N_2983);
nor UO_51 (O_51,N_2958,N_2956);
nand UO_52 (O_52,N_2988,N_2940);
nor UO_53 (O_53,N_2997,N_2996);
or UO_54 (O_54,N_2966,N_2956);
nor UO_55 (O_55,N_2999,N_2936);
and UO_56 (O_56,N_2956,N_2955);
and UO_57 (O_57,N_2945,N_2954);
and UO_58 (O_58,N_2943,N_2980);
nor UO_59 (O_59,N_2993,N_2994);
nand UO_60 (O_60,N_2927,N_2926);
nor UO_61 (O_61,N_2961,N_2926);
and UO_62 (O_62,N_2997,N_2941);
or UO_63 (O_63,N_2943,N_2948);
or UO_64 (O_64,N_2928,N_2957);
and UO_65 (O_65,N_2933,N_2942);
and UO_66 (O_66,N_2948,N_2994);
and UO_67 (O_67,N_2958,N_2963);
and UO_68 (O_68,N_2974,N_2970);
nor UO_69 (O_69,N_2949,N_2944);
nor UO_70 (O_70,N_2974,N_2980);
and UO_71 (O_71,N_2949,N_2979);
nor UO_72 (O_72,N_2925,N_2997);
and UO_73 (O_73,N_2960,N_2957);
or UO_74 (O_74,N_2988,N_2933);
and UO_75 (O_75,N_2940,N_2986);
or UO_76 (O_76,N_2949,N_2953);
nor UO_77 (O_77,N_2994,N_2985);
or UO_78 (O_78,N_2999,N_2970);
or UO_79 (O_79,N_2963,N_2933);
and UO_80 (O_80,N_2941,N_2996);
nor UO_81 (O_81,N_2962,N_2997);
nor UO_82 (O_82,N_2952,N_2972);
and UO_83 (O_83,N_2997,N_2937);
or UO_84 (O_84,N_2979,N_2930);
nor UO_85 (O_85,N_2940,N_2946);
nor UO_86 (O_86,N_2975,N_2961);
and UO_87 (O_87,N_2951,N_2988);
nand UO_88 (O_88,N_2928,N_2993);
or UO_89 (O_89,N_2978,N_2977);
and UO_90 (O_90,N_2978,N_2935);
nand UO_91 (O_91,N_2981,N_2971);
nand UO_92 (O_92,N_2996,N_2937);
or UO_93 (O_93,N_2939,N_2949);
nand UO_94 (O_94,N_2986,N_2977);
and UO_95 (O_95,N_2946,N_2953);
and UO_96 (O_96,N_2981,N_2931);
nor UO_97 (O_97,N_2968,N_2949);
or UO_98 (O_98,N_2956,N_2960);
or UO_99 (O_99,N_2973,N_2971);
nand UO_100 (O_100,N_2962,N_2992);
nor UO_101 (O_101,N_2935,N_2971);
nand UO_102 (O_102,N_2978,N_2993);
or UO_103 (O_103,N_2928,N_2992);
or UO_104 (O_104,N_2966,N_2949);
nand UO_105 (O_105,N_2963,N_2999);
or UO_106 (O_106,N_2960,N_2971);
nor UO_107 (O_107,N_2966,N_2947);
or UO_108 (O_108,N_2961,N_2940);
nand UO_109 (O_109,N_2979,N_2993);
or UO_110 (O_110,N_2994,N_2927);
nand UO_111 (O_111,N_2958,N_2995);
nor UO_112 (O_112,N_2972,N_2926);
nand UO_113 (O_113,N_2964,N_2944);
xor UO_114 (O_114,N_2970,N_2990);
nand UO_115 (O_115,N_2997,N_2951);
or UO_116 (O_116,N_2944,N_2994);
nor UO_117 (O_117,N_2952,N_2926);
or UO_118 (O_118,N_2928,N_2972);
nand UO_119 (O_119,N_2996,N_2990);
or UO_120 (O_120,N_2958,N_2967);
nor UO_121 (O_121,N_2926,N_2962);
or UO_122 (O_122,N_2977,N_2991);
nand UO_123 (O_123,N_2963,N_2984);
and UO_124 (O_124,N_2971,N_2926);
or UO_125 (O_125,N_2979,N_2956);
nand UO_126 (O_126,N_2952,N_2950);
nor UO_127 (O_127,N_2963,N_2985);
nand UO_128 (O_128,N_2936,N_2993);
and UO_129 (O_129,N_2997,N_2982);
nand UO_130 (O_130,N_2983,N_2950);
nand UO_131 (O_131,N_2986,N_2928);
and UO_132 (O_132,N_2928,N_2969);
nor UO_133 (O_133,N_2989,N_2945);
nor UO_134 (O_134,N_2990,N_2964);
nor UO_135 (O_135,N_2934,N_2930);
and UO_136 (O_136,N_2972,N_2957);
nand UO_137 (O_137,N_2957,N_2992);
nor UO_138 (O_138,N_2950,N_2926);
nor UO_139 (O_139,N_2944,N_2935);
nand UO_140 (O_140,N_2971,N_2958);
or UO_141 (O_141,N_2950,N_2938);
nand UO_142 (O_142,N_2959,N_2997);
nor UO_143 (O_143,N_2987,N_2956);
xor UO_144 (O_144,N_2937,N_2945);
and UO_145 (O_145,N_2977,N_2964);
nand UO_146 (O_146,N_2989,N_2947);
xnor UO_147 (O_147,N_2941,N_2967);
or UO_148 (O_148,N_2993,N_2998);
or UO_149 (O_149,N_2933,N_2990);
nor UO_150 (O_150,N_2977,N_2972);
and UO_151 (O_151,N_2976,N_2978);
nor UO_152 (O_152,N_2991,N_2967);
xor UO_153 (O_153,N_2930,N_2931);
and UO_154 (O_154,N_2944,N_2958);
nand UO_155 (O_155,N_2962,N_2935);
and UO_156 (O_156,N_2946,N_2959);
nand UO_157 (O_157,N_2980,N_2935);
nor UO_158 (O_158,N_2985,N_2954);
nor UO_159 (O_159,N_2931,N_2970);
nor UO_160 (O_160,N_2988,N_2939);
nor UO_161 (O_161,N_2926,N_2979);
nor UO_162 (O_162,N_2990,N_2994);
and UO_163 (O_163,N_2936,N_2972);
nor UO_164 (O_164,N_2971,N_2942);
and UO_165 (O_165,N_2974,N_2984);
or UO_166 (O_166,N_2932,N_2945);
or UO_167 (O_167,N_2945,N_2957);
or UO_168 (O_168,N_2938,N_2968);
nand UO_169 (O_169,N_2943,N_2997);
or UO_170 (O_170,N_2992,N_2941);
or UO_171 (O_171,N_2929,N_2997);
and UO_172 (O_172,N_2956,N_2975);
xnor UO_173 (O_173,N_2953,N_2993);
nor UO_174 (O_174,N_2961,N_2930);
and UO_175 (O_175,N_2999,N_2994);
and UO_176 (O_176,N_2973,N_2960);
nor UO_177 (O_177,N_2963,N_2938);
or UO_178 (O_178,N_2974,N_2972);
nor UO_179 (O_179,N_2993,N_2934);
nand UO_180 (O_180,N_2926,N_2946);
or UO_181 (O_181,N_2984,N_2944);
or UO_182 (O_182,N_2979,N_2953);
and UO_183 (O_183,N_2989,N_2957);
and UO_184 (O_184,N_2971,N_2940);
or UO_185 (O_185,N_2976,N_2968);
nand UO_186 (O_186,N_2965,N_2991);
nor UO_187 (O_187,N_2927,N_2989);
nor UO_188 (O_188,N_2943,N_2951);
nor UO_189 (O_189,N_2946,N_2991);
or UO_190 (O_190,N_2995,N_2986);
nand UO_191 (O_191,N_2994,N_2926);
or UO_192 (O_192,N_2968,N_2979);
or UO_193 (O_193,N_2952,N_2964);
nor UO_194 (O_194,N_2951,N_2989);
or UO_195 (O_195,N_2938,N_2977);
nand UO_196 (O_196,N_2962,N_2961);
nor UO_197 (O_197,N_2989,N_2985);
and UO_198 (O_198,N_2980,N_2953);
nand UO_199 (O_199,N_2962,N_2993);
nand UO_200 (O_200,N_2960,N_2969);
or UO_201 (O_201,N_2994,N_2975);
or UO_202 (O_202,N_2946,N_2967);
and UO_203 (O_203,N_2942,N_2944);
or UO_204 (O_204,N_2978,N_2973);
nor UO_205 (O_205,N_2977,N_2927);
xor UO_206 (O_206,N_2925,N_2935);
nand UO_207 (O_207,N_2980,N_2981);
nor UO_208 (O_208,N_2956,N_2926);
or UO_209 (O_209,N_2947,N_2929);
nor UO_210 (O_210,N_2949,N_2962);
or UO_211 (O_211,N_2960,N_2977);
nand UO_212 (O_212,N_2971,N_2961);
nor UO_213 (O_213,N_2993,N_2927);
nor UO_214 (O_214,N_2931,N_2965);
or UO_215 (O_215,N_2993,N_2964);
and UO_216 (O_216,N_2956,N_2927);
or UO_217 (O_217,N_2947,N_2954);
or UO_218 (O_218,N_2950,N_2968);
nand UO_219 (O_219,N_2990,N_2992);
nand UO_220 (O_220,N_2972,N_2959);
nand UO_221 (O_221,N_2937,N_2957);
nand UO_222 (O_222,N_2938,N_2993);
nand UO_223 (O_223,N_2976,N_2984);
or UO_224 (O_224,N_2975,N_2984);
nand UO_225 (O_225,N_2974,N_2926);
or UO_226 (O_226,N_2968,N_2933);
nor UO_227 (O_227,N_2995,N_2940);
or UO_228 (O_228,N_2991,N_2930);
or UO_229 (O_229,N_2952,N_2928);
and UO_230 (O_230,N_2963,N_2989);
nor UO_231 (O_231,N_2987,N_2934);
nor UO_232 (O_232,N_2977,N_2973);
or UO_233 (O_233,N_2948,N_2980);
and UO_234 (O_234,N_2930,N_2948);
nor UO_235 (O_235,N_2953,N_2959);
nand UO_236 (O_236,N_2960,N_2925);
and UO_237 (O_237,N_2981,N_2983);
nand UO_238 (O_238,N_2968,N_2951);
or UO_239 (O_239,N_2927,N_2955);
nor UO_240 (O_240,N_2978,N_2981);
or UO_241 (O_241,N_2969,N_2935);
nand UO_242 (O_242,N_2958,N_2985);
nor UO_243 (O_243,N_2957,N_2968);
nor UO_244 (O_244,N_2939,N_2991);
or UO_245 (O_245,N_2934,N_2961);
nand UO_246 (O_246,N_2992,N_2985);
or UO_247 (O_247,N_2982,N_2938);
nand UO_248 (O_248,N_2941,N_2928);
nor UO_249 (O_249,N_2925,N_2983);
and UO_250 (O_250,N_2933,N_2960);
and UO_251 (O_251,N_2948,N_2934);
or UO_252 (O_252,N_2975,N_2932);
and UO_253 (O_253,N_2995,N_2998);
or UO_254 (O_254,N_2983,N_2973);
or UO_255 (O_255,N_2943,N_2942);
nand UO_256 (O_256,N_2934,N_2988);
or UO_257 (O_257,N_2951,N_2965);
and UO_258 (O_258,N_2943,N_2938);
or UO_259 (O_259,N_2973,N_2975);
or UO_260 (O_260,N_2996,N_2969);
and UO_261 (O_261,N_2936,N_2942);
nor UO_262 (O_262,N_2932,N_2993);
or UO_263 (O_263,N_2968,N_2990);
nand UO_264 (O_264,N_2934,N_2986);
or UO_265 (O_265,N_2958,N_2960);
and UO_266 (O_266,N_2956,N_2992);
or UO_267 (O_267,N_2962,N_2928);
nand UO_268 (O_268,N_2927,N_2982);
or UO_269 (O_269,N_2930,N_2952);
nor UO_270 (O_270,N_2958,N_2990);
and UO_271 (O_271,N_2932,N_2998);
nand UO_272 (O_272,N_2925,N_2976);
nor UO_273 (O_273,N_2959,N_2980);
nand UO_274 (O_274,N_2996,N_2931);
nor UO_275 (O_275,N_2934,N_2956);
nand UO_276 (O_276,N_2951,N_2982);
nor UO_277 (O_277,N_2932,N_2948);
and UO_278 (O_278,N_2934,N_2974);
nand UO_279 (O_279,N_2967,N_2975);
or UO_280 (O_280,N_2977,N_2959);
or UO_281 (O_281,N_2937,N_2986);
nor UO_282 (O_282,N_2987,N_2967);
nor UO_283 (O_283,N_2940,N_2931);
nand UO_284 (O_284,N_2985,N_2977);
nor UO_285 (O_285,N_2954,N_2939);
nand UO_286 (O_286,N_2927,N_2991);
and UO_287 (O_287,N_2930,N_2973);
or UO_288 (O_288,N_2994,N_2969);
and UO_289 (O_289,N_2962,N_2972);
and UO_290 (O_290,N_2999,N_2954);
nand UO_291 (O_291,N_2992,N_2942);
or UO_292 (O_292,N_2926,N_2996);
nor UO_293 (O_293,N_2974,N_2989);
nor UO_294 (O_294,N_2963,N_2942);
or UO_295 (O_295,N_2966,N_2934);
or UO_296 (O_296,N_2968,N_2978);
or UO_297 (O_297,N_2971,N_2959);
nand UO_298 (O_298,N_2962,N_2977);
and UO_299 (O_299,N_2925,N_2943);
nand UO_300 (O_300,N_2925,N_2965);
nor UO_301 (O_301,N_2960,N_2959);
nand UO_302 (O_302,N_2960,N_2935);
and UO_303 (O_303,N_2984,N_2950);
nor UO_304 (O_304,N_2970,N_2943);
or UO_305 (O_305,N_2938,N_2948);
nand UO_306 (O_306,N_2960,N_2996);
nor UO_307 (O_307,N_2985,N_2937);
and UO_308 (O_308,N_2947,N_2957);
and UO_309 (O_309,N_2969,N_2982);
nor UO_310 (O_310,N_2959,N_2943);
or UO_311 (O_311,N_2981,N_2961);
nor UO_312 (O_312,N_2959,N_2989);
and UO_313 (O_313,N_2953,N_2968);
and UO_314 (O_314,N_2976,N_2941);
and UO_315 (O_315,N_2979,N_2994);
or UO_316 (O_316,N_2975,N_2969);
nor UO_317 (O_317,N_2979,N_2959);
and UO_318 (O_318,N_2983,N_2930);
and UO_319 (O_319,N_2959,N_2958);
nor UO_320 (O_320,N_2949,N_2933);
and UO_321 (O_321,N_2953,N_2942);
nor UO_322 (O_322,N_2997,N_2950);
or UO_323 (O_323,N_2973,N_2945);
or UO_324 (O_324,N_2947,N_2931);
or UO_325 (O_325,N_2932,N_2988);
or UO_326 (O_326,N_2957,N_2958);
or UO_327 (O_327,N_2986,N_2981);
or UO_328 (O_328,N_2996,N_2978);
or UO_329 (O_329,N_2994,N_2934);
or UO_330 (O_330,N_2980,N_2937);
or UO_331 (O_331,N_2986,N_2958);
or UO_332 (O_332,N_2958,N_2929);
xnor UO_333 (O_333,N_2974,N_2963);
nand UO_334 (O_334,N_2969,N_2929);
xnor UO_335 (O_335,N_2925,N_2988);
and UO_336 (O_336,N_2930,N_2926);
nor UO_337 (O_337,N_2930,N_2978);
and UO_338 (O_338,N_2977,N_2969);
nor UO_339 (O_339,N_2944,N_2931);
and UO_340 (O_340,N_2988,N_2946);
nand UO_341 (O_341,N_2994,N_2989);
nand UO_342 (O_342,N_2999,N_2988);
nand UO_343 (O_343,N_2947,N_2979);
and UO_344 (O_344,N_2952,N_2995);
nand UO_345 (O_345,N_2941,N_2948);
or UO_346 (O_346,N_2978,N_2936);
or UO_347 (O_347,N_2942,N_2952);
nand UO_348 (O_348,N_2997,N_2939);
and UO_349 (O_349,N_2932,N_2987);
nand UO_350 (O_350,N_2932,N_2991);
nand UO_351 (O_351,N_2928,N_2989);
nor UO_352 (O_352,N_2960,N_2934);
and UO_353 (O_353,N_2947,N_2956);
nor UO_354 (O_354,N_2943,N_2933);
nor UO_355 (O_355,N_2961,N_2956);
or UO_356 (O_356,N_2993,N_2925);
nor UO_357 (O_357,N_2964,N_2945);
nand UO_358 (O_358,N_2988,N_2937);
nor UO_359 (O_359,N_2990,N_2983);
xor UO_360 (O_360,N_2999,N_2991);
nor UO_361 (O_361,N_2939,N_2959);
nor UO_362 (O_362,N_2939,N_2942);
nor UO_363 (O_363,N_2975,N_2955);
nand UO_364 (O_364,N_2965,N_2950);
nor UO_365 (O_365,N_2959,N_2988);
nand UO_366 (O_366,N_2955,N_2976);
nand UO_367 (O_367,N_2943,N_2939);
or UO_368 (O_368,N_2997,N_2989);
or UO_369 (O_369,N_2964,N_2961);
nor UO_370 (O_370,N_2933,N_2938);
nand UO_371 (O_371,N_2959,N_2974);
or UO_372 (O_372,N_2959,N_2926);
nor UO_373 (O_373,N_2948,N_2976);
nand UO_374 (O_374,N_2986,N_2948);
nand UO_375 (O_375,N_2937,N_2987);
nand UO_376 (O_376,N_2994,N_2940);
and UO_377 (O_377,N_2989,N_2934);
and UO_378 (O_378,N_2964,N_2991);
and UO_379 (O_379,N_2965,N_2946);
or UO_380 (O_380,N_2981,N_2952);
and UO_381 (O_381,N_2962,N_2954);
or UO_382 (O_382,N_2960,N_2990);
nand UO_383 (O_383,N_2982,N_2948);
and UO_384 (O_384,N_2955,N_2953);
nand UO_385 (O_385,N_2928,N_2934);
nand UO_386 (O_386,N_2954,N_2950);
nor UO_387 (O_387,N_2969,N_2981);
and UO_388 (O_388,N_2944,N_2985);
nor UO_389 (O_389,N_2939,N_2936);
nor UO_390 (O_390,N_2932,N_2949);
nor UO_391 (O_391,N_2983,N_2943);
nor UO_392 (O_392,N_2958,N_2937);
or UO_393 (O_393,N_2960,N_2994);
nor UO_394 (O_394,N_2937,N_2989);
nand UO_395 (O_395,N_2926,N_2986);
nor UO_396 (O_396,N_2957,N_2965);
nand UO_397 (O_397,N_2986,N_2982);
nand UO_398 (O_398,N_2961,N_2999);
and UO_399 (O_399,N_2947,N_2952);
or UO_400 (O_400,N_2991,N_2995);
and UO_401 (O_401,N_2985,N_2960);
nor UO_402 (O_402,N_2936,N_2935);
nand UO_403 (O_403,N_2966,N_2992);
nand UO_404 (O_404,N_2992,N_2949);
or UO_405 (O_405,N_2983,N_2932);
nor UO_406 (O_406,N_2934,N_2937);
nand UO_407 (O_407,N_2944,N_2925);
or UO_408 (O_408,N_2961,N_2966);
and UO_409 (O_409,N_2999,N_2945);
nor UO_410 (O_410,N_2939,N_2931);
nand UO_411 (O_411,N_2998,N_2963);
or UO_412 (O_412,N_2964,N_2955);
or UO_413 (O_413,N_2988,N_2979);
and UO_414 (O_414,N_2939,N_2966);
nand UO_415 (O_415,N_2969,N_2952);
nor UO_416 (O_416,N_2943,N_2978);
and UO_417 (O_417,N_2990,N_2966);
or UO_418 (O_418,N_2973,N_2933);
nand UO_419 (O_419,N_2993,N_2946);
nor UO_420 (O_420,N_2974,N_2976);
and UO_421 (O_421,N_2974,N_2941);
or UO_422 (O_422,N_2930,N_2969);
and UO_423 (O_423,N_2979,N_2986);
nor UO_424 (O_424,N_2929,N_2941);
or UO_425 (O_425,N_2980,N_2961);
or UO_426 (O_426,N_2952,N_2996);
or UO_427 (O_427,N_2944,N_2976);
nand UO_428 (O_428,N_2963,N_2988);
nor UO_429 (O_429,N_2935,N_2982);
nand UO_430 (O_430,N_2925,N_2956);
nor UO_431 (O_431,N_2932,N_2947);
and UO_432 (O_432,N_2928,N_2926);
nand UO_433 (O_433,N_2992,N_2967);
nand UO_434 (O_434,N_2997,N_2990);
or UO_435 (O_435,N_2992,N_2979);
nor UO_436 (O_436,N_2983,N_2951);
and UO_437 (O_437,N_2935,N_2976);
nand UO_438 (O_438,N_2982,N_2949);
nor UO_439 (O_439,N_2977,N_2945);
nor UO_440 (O_440,N_2963,N_2925);
and UO_441 (O_441,N_2988,N_2982);
and UO_442 (O_442,N_2968,N_2999);
nand UO_443 (O_443,N_2942,N_2996);
and UO_444 (O_444,N_2947,N_2943);
nand UO_445 (O_445,N_2983,N_2966);
or UO_446 (O_446,N_2976,N_2956);
and UO_447 (O_447,N_2958,N_2992);
nor UO_448 (O_448,N_2966,N_2998);
or UO_449 (O_449,N_2997,N_2935);
or UO_450 (O_450,N_2978,N_2940);
nor UO_451 (O_451,N_2940,N_2960);
nand UO_452 (O_452,N_2966,N_2948);
and UO_453 (O_453,N_2974,N_2927);
or UO_454 (O_454,N_2978,N_2982);
and UO_455 (O_455,N_2946,N_2952);
and UO_456 (O_456,N_2957,N_2988);
nand UO_457 (O_457,N_2961,N_2925);
xor UO_458 (O_458,N_2950,N_2990);
nand UO_459 (O_459,N_2956,N_2969);
nor UO_460 (O_460,N_2973,N_2934);
nand UO_461 (O_461,N_2979,N_2969);
nor UO_462 (O_462,N_2986,N_2989);
and UO_463 (O_463,N_2996,N_2999);
nor UO_464 (O_464,N_2991,N_2958);
and UO_465 (O_465,N_2987,N_2989);
nor UO_466 (O_466,N_2931,N_2936);
or UO_467 (O_467,N_2976,N_2942);
nor UO_468 (O_468,N_2925,N_2954);
and UO_469 (O_469,N_2934,N_2940);
nand UO_470 (O_470,N_2995,N_2968);
and UO_471 (O_471,N_2984,N_2937);
nand UO_472 (O_472,N_2994,N_2984);
and UO_473 (O_473,N_2990,N_2947);
nand UO_474 (O_474,N_2983,N_2965);
and UO_475 (O_475,N_2971,N_2970);
nor UO_476 (O_476,N_2987,N_2966);
nand UO_477 (O_477,N_2989,N_2981);
and UO_478 (O_478,N_2935,N_2951);
and UO_479 (O_479,N_2989,N_2960);
nor UO_480 (O_480,N_2944,N_2993);
or UO_481 (O_481,N_2964,N_2929);
or UO_482 (O_482,N_2982,N_2973);
nor UO_483 (O_483,N_2964,N_2975);
nor UO_484 (O_484,N_2926,N_2945);
and UO_485 (O_485,N_2931,N_2960);
or UO_486 (O_486,N_2948,N_2999);
or UO_487 (O_487,N_2992,N_2963);
or UO_488 (O_488,N_2939,N_2969);
nand UO_489 (O_489,N_2936,N_2977);
or UO_490 (O_490,N_2937,N_2925);
or UO_491 (O_491,N_2943,N_2960);
nor UO_492 (O_492,N_2960,N_2930);
nand UO_493 (O_493,N_2941,N_2990);
or UO_494 (O_494,N_2935,N_2963);
and UO_495 (O_495,N_2943,N_2944);
nor UO_496 (O_496,N_2977,N_2963);
xnor UO_497 (O_497,N_2986,N_2930);
nand UO_498 (O_498,N_2988,N_2974);
nor UO_499 (O_499,N_2954,N_2960);
endmodule