module basic_500_3000_500_30_levels_2xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_354,In_36);
or U1 (N_1,In_332,In_189);
or U2 (N_2,In_163,In_208);
nor U3 (N_3,In_307,In_203);
nor U4 (N_4,In_190,In_29);
nor U5 (N_5,In_37,In_458);
or U6 (N_6,In_169,In_402);
nand U7 (N_7,In_6,In_1);
nand U8 (N_8,In_272,In_202);
or U9 (N_9,In_434,In_339);
or U10 (N_10,In_448,In_247);
xnor U11 (N_11,In_97,In_289);
nor U12 (N_12,In_368,In_445);
and U13 (N_13,In_422,In_323);
and U14 (N_14,In_432,In_59);
nand U15 (N_15,In_39,In_285);
nor U16 (N_16,In_188,In_362);
nand U17 (N_17,In_137,In_386);
or U18 (N_18,In_266,In_216);
or U19 (N_19,In_337,In_33);
nand U20 (N_20,In_122,In_199);
nor U21 (N_21,In_172,In_485);
nor U22 (N_22,In_437,In_406);
or U23 (N_23,In_193,In_38);
and U24 (N_24,In_222,In_17);
nand U25 (N_25,In_306,In_413);
nand U26 (N_26,In_235,In_333);
nor U27 (N_27,In_239,In_185);
nor U28 (N_28,In_79,In_494);
and U29 (N_29,In_255,In_241);
or U30 (N_30,In_423,In_293);
or U31 (N_31,In_420,In_352);
nor U32 (N_32,In_135,In_336);
xor U33 (N_33,In_488,In_277);
and U34 (N_34,In_91,In_451);
nor U35 (N_35,In_150,In_35);
nor U36 (N_36,In_80,In_356);
nor U37 (N_37,In_56,In_378);
nand U38 (N_38,In_117,In_462);
nor U39 (N_39,In_81,In_447);
and U40 (N_40,In_477,In_192);
or U41 (N_41,In_391,In_63);
nand U42 (N_42,In_111,In_128);
nand U43 (N_43,In_262,In_85);
nand U44 (N_44,In_438,In_347);
or U45 (N_45,In_148,In_384);
or U46 (N_46,In_357,In_496);
and U47 (N_47,In_471,In_53);
and U48 (N_48,In_180,In_321);
nand U49 (N_49,In_344,In_3);
nand U50 (N_50,In_475,In_160);
or U51 (N_51,In_400,In_147);
nand U52 (N_52,In_416,In_8);
or U53 (N_53,In_32,In_196);
nand U54 (N_54,In_125,In_304);
nor U55 (N_55,In_72,In_0);
nor U56 (N_56,In_459,In_58);
nor U57 (N_57,In_449,In_439);
nor U58 (N_58,In_452,In_179);
or U59 (N_59,In_65,In_280);
nor U60 (N_60,In_234,In_489);
nor U61 (N_61,In_48,In_399);
nand U62 (N_62,In_456,In_22);
and U63 (N_63,In_139,In_71);
or U64 (N_64,In_98,In_134);
nand U65 (N_65,In_90,In_204);
nor U66 (N_66,In_294,In_338);
and U67 (N_67,In_40,In_110);
nand U68 (N_68,In_360,In_151);
and U69 (N_69,In_181,In_237);
nand U70 (N_70,In_232,In_211);
nand U71 (N_71,In_14,In_5);
and U72 (N_72,In_206,In_101);
nand U73 (N_73,In_153,In_442);
or U74 (N_74,In_259,In_92);
or U75 (N_75,In_453,In_220);
nand U76 (N_76,In_13,In_213);
nand U77 (N_77,In_491,In_34);
nand U78 (N_78,In_371,In_457);
or U79 (N_79,In_184,In_55);
or U80 (N_80,In_230,In_221);
or U81 (N_81,In_301,In_21);
or U82 (N_82,In_102,In_145);
nand U83 (N_83,In_446,In_300);
xor U84 (N_84,In_397,In_274);
nor U85 (N_85,In_279,In_299);
nor U86 (N_86,In_162,In_296);
and U87 (N_87,In_465,In_467);
and U88 (N_88,In_257,In_398);
or U89 (N_89,In_317,In_4);
xor U90 (N_90,In_144,In_407);
nor U91 (N_91,In_325,In_115);
nor U92 (N_92,In_320,In_395);
nand U93 (N_93,In_200,In_236);
nor U94 (N_94,In_46,In_297);
nand U95 (N_95,In_108,In_426);
nor U96 (N_96,In_404,In_441);
nor U97 (N_97,In_224,In_27);
nand U98 (N_98,In_258,In_41);
and U99 (N_99,In_478,In_312);
nand U100 (N_100,In_363,N_95);
nand U101 (N_101,N_53,N_70);
and U102 (N_102,In_149,In_86);
nand U103 (N_103,In_248,N_67);
and U104 (N_104,N_86,N_96);
nor U105 (N_105,In_177,N_54);
nor U106 (N_106,In_468,In_89);
and U107 (N_107,In_374,In_167);
and U108 (N_108,N_60,In_346);
nand U109 (N_109,In_493,In_201);
or U110 (N_110,In_340,In_264);
and U111 (N_111,In_245,In_372);
or U112 (N_112,N_77,In_12);
or U113 (N_113,In_73,In_311);
and U114 (N_114,N_4,In_136);
and U115 (N_115,In_278,In_409);
nor U116 (N_116,In_256,In_127);
nand U117 (N_117,N_61,N_6);
or U118 (N_118,In_242,In_394);
and U119 (N_119,N_33,N_32);
or U120 (N_120,N_55,In_268);
nand U121 (N_121,In_76,In_315);
nor U122 (N_122,In_411,In_252);
nand U123 (N_123,In_49,In_381);
nor U124 (N_124,N_64,In_164);
nor U125 (N_125,In_157,In_263);
and U126 (N_126,In_298,N_69);
and U127 (N_127,N_16,In_25);
or U128 (N_128,In_143,N_52);
nand U129 (N_129,N_29,N_8);
nor U130 (N_130,In_480,In_385);
nand U131 (N_131,N_2,In_95);
nor U132 (N_132,In_31,In_361);
nand U133 (N_133,In_440,In_223);
nor U134 (N_134,N_35,In_341);
or U135 (N_135,N_5,In_225);
or U136 (N_136,In_316,In_209);
and U137 (N_137,In_50,In_173);
or U138 (N_138,In_205,In_295);
or U139 (N_139,N_87,In_355);
nand U140 (N_140,In_93,N_93);
or U141 (N_141,In_42,In_82);
nand U142 (N_142,In_331,In_335);
nand U143 (N_143,N_36,In_229);
nor U144 (N_144,N_31,N_30);
or U145 (N_145,In_275,In_328);
and U146 (N_146,In_365,In_15);
nor U147 (N_147,In_116,In_84);
and U148 (N_148,In_104,In_123);
nand U149 (N_149,In_159,In_175);
and U150 (N_150,N_63,In_253);
or U151 (N_151,In_318,In_350);
or U152 (N_152,N_68,N_83);
nand U153 (N_153,In_51,In_393);
or U154 (N_154,In_133,In_497);
and U155 (N_155,In_178,N_80);
nor U156 (N_156,In_120,In_498);
nor U157 (N_157,In_26,In_313);
and U158 (N_158,In_342,In_228);
and U159 (N_159,In_246,In_182);
nor U160 (N_160,In_219,In_415);
nor U161 (N_161,In_210,In_414);
or U162 (N_162,N_37,In_10);
and U163 (N_163,In_45,N_65);
nand U164 (N_164,In_158,N_50);
or U165 (N_165,In_270,N_58);
and U166 (N_166,N_38,In_130);
or U167 (N_167,In_142,In_240);
nor U168 (N_168,In_118,In_377);
nor U169 (N_169,N_78,In_330);
and U170 (N_170,In_176,In_309);
nor U171 (N_171,In_233,In_212);
nand U172 (N_172,In_19,N_79);
nor U173 (N_173,In_484,N_14);
nand U174 (N_174,N_57,N_94);
nor U175 (N_175,In_74,In_121);
nand U176 (N_176,N_48,In_387);
nand U177 (N_177,In_100,In_288);
and U178 (N_178,In_345,N_42);
nor U179 (N_179,In_170,In_47);
xnor U180 (N_180,N_82,In_479);
or U181 (N_181,N_71,In_326);
or U182 (N_182,In_124,In_249);
nand U183 (N_183,In_291,N_98);
nor U184 (N_184,N_46,N_21);
or U185 (N_185,N_40,In_197);
or U186 (N_186,In_113,In_367);
and U187 (N_187,In_69,In_392);
or U188 (N_188,N_56,In_303);
nand U189 (N_189,N_92,In_418);
nor U190 (N_190,In_161,In_2);
nand U191 (N_191,In_433,In_88);
and U192 (N_192,N_25,In_310);
or U193 (N_193,N_0,In_66);
or U194 (N_194,In_429,In_43);
nand U195 (N_195,In_70,In_54);
nor U196 (N_196,In_327,In_155);
and U197 (N_197,N_9,In_366);
nand U198 (N_198,N_49,In_322);
or U199 (N_199,In_427,In_218);
nand U200 (N_200,N_91,In_67);
and U201 (N_201,In_382,In_75);
and U202 (N_202,N_34,N_162);
nor U203 (N_203,N_3,In_403);
and U204 (N_204,N_152,In_112);
nand U205 (N_205,N_66,N_127);
and U206 (N_206,In_482,In_383);
nand U207 (N_207,In_343,N_169);
nor U208 (N_208,N_139,N_19);
and U209 (N_209,N_85,N_108);
and U210 (N_210,N_13,In_472);
nand U211 (N_211,N_188,In_138);
or U212 (N_212,N_51,N_181);
nor U213 (N_213,In_455,In_460);
or U214 (N_214,In_454,In_349);
or U215 (N_215,N_124,In_131);
nand U216 (N_216,N_153,In_492);
or U217 (N_217,In_469,In_373);
or U218 (N_218,N_116,N_190);
nor U219 (N_219,In_412,N_185);
nand U220 (N_220,In_271,In_464);
nand U221 (N_221,N_155,In_474);
nand U222 (N_222,In_466,In_62);
or U223 (N_223,N_187,N_84);
and U224 (N_224,N_100,N_20);
and U225 (N_225,N_39,N_151);
and U226 (N_226,In_430,N_141);
nand U227 (N_227,N_115,In_292);
nand U228 (N_228,In_94,N_43);
nor U229 (N_229,N_73,In_132);
nand U230 (N_230,In_281,N_74);
or U231 (N_231,N_111,N_182);
nand U232 (N_232,In_99,In_261);
nand U233 (N_233,N_176,In_227);
and U234 (N_234,In_370,N_109);
nor U235 (N_235,N_17,N_22);
nor U236 (N_236,N_107,N_158);
and U237 (N_237,In_334,In_165);
nor U238 (N_238,N_113,N_179);
and U239 (N_239,In_435,N_163);
or U240 (N_240,In_23,N_75);
nor U241 (N_241,In_364,In_156);
nand U242 (N_242,In_30,In_96);
and U243 (N_243,In_9,In_276);
nand U244 (N_244,N_183,N_101);
nand U245 (N_245,In_408,In_486);
nor U246 (N_246,N_129,N_135);
nand U247 (N_247,In_114,N_97);
nand U248 (N_248,N_89,N_122);
or U249 (N_249,N_167,In_61);
or U250 (N_250,N_11,In_286);
and U251 (N_251,In_140,In_390);
and U252 (N_252,In_238,In_183);
nor U253 (N_253,In_166,N_119);
and U254 (N_254,N_146,N_136);
nand U255 (N_255,In_282,In_87);
and U256 (N_256,In_254,In_380);
or U257 (N_257,N_18,In_405);
nand U258 (N_258,N_166,N_159);
xor U259 (N_259,N_154,In_436);
xor U260 (N_260,N_145,In_473);
or U261 (N_261,In_251,N_149);
and U262 (N_262,In_107,In_152);
or U263 (N_263,N_7,N_157);
or U264 (N_264,N_103,N_106);
or U265 (N_265,In_119,In_444);
nor U266 (N_266,N_112,N_137);
nand U267 (N_267,N_125,N_1);
nand U268 (N_268,In_284,In_106);
nor U269 (N_269,In_187,In_267);
and U270 (N_270,In_18,In_290);
nand U271 (N_271,In_305,N_41);
and U272 (N_272,In_215,In_194);
nor U273 (N_273,N_142,In_421);
nor U274 (N_274,In_481,In_324);
nor U275 (N_275,In_483,N_134);
or U276 (N_276,In_287,N_104);
and U277 (N_277,In_129,In_7);
nand U278 (N_278,In_103,In_250);
nand U279 (N_279,N_150,In_171);
and U280 (N_280,N_102,In_191);
or U281 (N_281,In_265,N_59);
nand U282 (N_282,N_88,N_128);
nand U283 (N_283,N_133,In_353);
and U284 (N_284,In_243,In_146);
nor U285 (N_285,N_175,N_143);
nand U286 (N_286,N_105,N_138);
or U287 (N_287,In_425,In_490);
nor U288 (N_288,N_193,In_283);
or U289 (N_289,N_81,N_148);
nor U290 (N_290,In_260,N_99);
nor U291 (N_291,In_207,N_172);
or U292 (N_292,N_24,In_389);
or U293 (N_293,In_16,N_195);
nand U294 (N_294,In_154,In_375);
nand U295 (N_295,In_186,N_45);
nand U296 (N_296,In_64,In_359);
and U297 (N_297,N_178,In_77);
nand U298 (N_298,In_308,N_170);
or U299 (N_299,In_168,In_329);
nand U300 (N_300,N_267,N_207);
and U301 (N_301,N_173,In_24);
nand U302 (N_302,N_232,N_214);
and U303 (N_303,N_277,N_215);
nor U304 (N_304,N_228,In_495);
nor U305 (N_305,N_28,N_272);
and U306 (N_306,N_191,N_250);
nor U307 (N_307,In_68,N_126);
and U308 (N_308,N_171,In_476);
nand U309 (N_309,N_262,In_463);
and U310 (N_310,N_230,In_109);
and U311 (N_311,In_44,N_288);
nor U312 (N_312,N_246,In_388);
nand U313 (N_313,N_144,N_217);
or U314 (N_314,N_239,N_275);
nor U315 (N_315,In_376,N_202);
and U316 (N_316,N_118,In_52);
and U317 (N_317,In_417,In_450);
and U318 (N_318,In_20,N_210);
nor U319 (N_319,N_226,In_379);
nor U320 (N_320,In_105,N_248);
nand U321 (N_321,N_121,N_203);
or U322 (N_322,N_130,N_254);
or U323 (N_323,N_23,N_256);
or U324 (N_324,N_278,N_114);
and U325 (N_325,N_238,In_78);
nor U326 (N_326,N_297,N_299);
nand U327 (N_327,N_276,N_12);
nand U328 (N_328,N_160,In_126);
or U329 (N_329,In_273,N_235);
or U330 (N_330,N_231,N_257);
xnor U331 (N_331,In_214,N_253);
nor U332 (N_332,N_205,In_410);
and U333 (N_333,N_192,In_348);
nand U334 (N_334,N_10,N_216);
nor U335 (N_335,In_470,N_177);
and U336 (N_336,N_211,N_266);
nand U337 (N_337,N_229,N_281);
nor U338 (N_338,N_298,N_237);
nor U339 (N_339,N_280,In_424);
or U340 (N_340,N_196,N_180);
nand U341 (N_341,In_198,N_295);
and U342 (N_342,In_351,N_225);
and U343 (N_343,In_28,N_234);
or U344 (N_344,N_164,N_209);
and U345 (N_345,N_251,N_223);
nand U346 (N_346,N_44,N_165);
and U347 (N_347,In_57,In_401);
nand U348 (N_348,N_156,N_247);
nand U349 (N_349,In_244,N_282);
nand U350 (N_350,N_62,N_200);
nand U351 (N_351,N_258,N_279);
or U352 (N_352,In_269,N_199);
nand U353 (N_353,In_396,In_431);
nor U354 (N_354,N_236,N_287);
nand U355 (N_355,In_83,In_314);
nor U356 (N_356,N_168,N_290);
or U357 (N_357,N_218,N_184);
nor U358 (N_358,N_213,N_240);
or U359 (N_359,In_499,N_15);
and U360 (N_360,N_221,In_358);
and U361 (N_361,In_217,In_369);
and U362 (N_362,N_27,N_110);
or U363 (N_363,N_132,In_461);
or U364 (N_364,In_174,N_194);
and U365 (N_365,N_220,N_123);
nor U366 (N_366,N_47,In_443);
nor U367 (N_367,In_60,N_197);
nand U368 (N_368,N_90,In_195);
and U369 (N_369,N_186,N_249);
or U370 (N_370,N_189,N_72);
or U371 (N_371,N_76,N_296);
or U372 (N_372,N_269,N_233);
nand U373 (N_373,N_292,N_283);
and U374 (N_374,N_243,N_265);
or U375 (N_375,N_212,In_419);
nand U376 (N_376,N_293,N_255);
nor U377 (N_377,In_319,N_260);
or U378 (N_378,In_141,N_264);
or U379 (N_379,In_226,N_244);
and U380 (N_380,N_284,N_219);
or U381 (N_381,N_261,N_263);
nand U382 (N_382,N_274,N_294);
or U383 (N_383,N_289,N_241);
nor U384 (N_384,In_428,N_270);
nor U385 (N_385,N_245,N_147);
or U386 (N_386,N_117,N_161);
xnor U387 (N_387,In_231,N_273);
nor U388 (N_388,N_198,N_26);
nand U389 (N_389,N_286,N_201);
xnor U390 (N_390,N_208,N_206);
nand U391 (N_391,N_227,In_487);
and U392 (N_392,N_131,N_285);
and U393 (N_393,N_174,N_204);
nor U394 (N_394,N_291,N_140);
nor U395 (N_395,N_259,In_302);
nor U396 (N_396,In_11,N_268);
nor U397 (N_397,N_271,N_222);
and U398 (N_398,N_224,N_120);
nor U399 (N_399,N_242,N_252);
or U400 (N_400,N_398,N_386);
or U401 (N_401,N_343,N_371);
and U402 (N_402,N_362,N_395);
nand U403 (N_403,N_321,N_388);
nor U404 (N_404,N_363,N_380);
and U405 (N_405,N_366,N_342);
nand U406 (N_406,N_399,N_346);
or U407 (N_407,N_300,N_344);
nor U408 (N_408,N_307,N_308);
and U409 (N_409,N_365,N_327);
and U410 (N_410,N_373,N_370);
nor U411 (N_411,N_301,N_368);
or U412 (N_412,N_339,N_312);
nand U413 (N_413,N_340,N_337);
nor U414 (N_414,N_392,N_377);
nand U415 (N_415,N_330,N_379);
or U416 (N_416,N_320,N_316);
and U417 (N_417,N_352,N_317);
and U418 (N_418,N_331,N_303);
and U419 (N_419,N_335,N_310);
and U420 (N_420,N_322,N_372);
and U421 (N_421,N_378,N_354);
nor U422 (N_422,N_383,N_324);
and U423 (N_423,N_391,N_338);
and U424 (N_424,N_359,N_393);
nand U425 (N_425,N_396,N_357);
xor U426 (N_426,N_328,N_302);
nor U427 (N_427,N_315,N_348);
and U428 (N_428,N_332,N_358);
and U429 (N_429,N_345,N_385);
nor U430 (N_430,N_319,N_361);
nand U431 (N_431,N_323,N_318);
and U432 (N_432,N_341,N_376);
and U433 (N_433,N_360,N_326);
and U434 (N_434,N_333,N_390);
and U435 (N_435,N_334,N_336);
nor U436 (N_436,N_364,N_355);
and U437 (N_437,N_347,N_349);
nor U438 (N_438,N_313,N_314);
or U439 (N_439,N_382,N_305);
or U440 (N_440,N_329,N_394);
nand U441 (N_441,N_374,N_397);
and U442 (N_442,N_309,N_304);
nand U443 (N_443,N_381,N_351);
nand U444 (N_444,N_384,N_369);
or U445 (N_445,N_306,N_356);
nand U446 (N_446,N_353,N_387);
and U447 (N_447,N_389,N_367);
or U448 (N_448,N_350,N_375);
or U449 (N_449,N_325,N_311);
nand U450 (N_450,N_368,N_316);
nor U451 (N_451,N_378,N_370);
and U452 (N_452,N_356,N_313);
xor U453 (N_453,N_318,N_303);
and U454 (N_454,N_353,N_373);
and U455 (N_455,N_387,N_364);
nor U456 (N_456,N_382,N_302);
and U457 (N_457,N_385,N_360);
nand U458 (N_458,N_331,N_381);
or U459 (N_459,N_330,N_393);
nor U460 (N_460,N_375,N_342);
nor U461 (N_461,N_350,N_394);
xor U462 (N_462,N_342,N_347);
nor U463 (N_463,N_386,N_302);
and U464 (N_464,N_393,N_382);
nor U465 (N_465,N_363,N_310);
nor U466 (N_466,N_345,N_356);
or U467 (N_467,N_300,N_375);
nor U468 (N_468,N_393,N_348);
xor U469 (N_469,N_334,N_379);
nand U470 (N_470,N_363,N_334);
xnor U471 (N_471,N_357,N_351);
xor U472 (N_472,N_368,N_382);
and U473 (N_473,N_326,N_346);
and U474 (N_474,N_368,N_363);
and U475 (N_475,N_335,N_320);
and U476 (N_476,N_372,N_391);
or U477 (N_477,N_380,N_381);
nand U478 (N_478,N_331,N_364);
or U479 (N_479,N_351,N_372);
nand U480 (N_480,N_308,N_328);
nand U481 (N_481,N_330,N_339);
or U482 (N_482,N_361,N_375);
or U483 (N_483,N_354,N_375);
or U484 (N_484,N_337,N_350);
nor U485 (N_485,N_363,N_348);
xnor U486 (N_486,N_399,N_385);
nor U487 (N_487,N_314,N_320);
nand U488 (N_488,N_369,N_358);
nand U489 (N_489,N_315,N_337);
nor U490 (N_490,N_374,N_363);
nand U491 (N_491,N_302,N_329);
or U492 (N_492,N_390,N_349);
nor U493 (N_493,N_396,N_361);
nand U494 (N_494,N_354,N_381);
nand U495 (N_495,N_349,N_309);
and U496 (N_496,N_310,N_307);
or U497 (N_497,N_364,N_322);
nor U498 (N_498,N_301,N_394);
nor U499 (N_499,N_305,N_339);
nand U500 (N_500,N_467,N_417);
or U501 (N_501,N_435,N_414);
nor U502 (N_502,N_453,N_405);
or U503 (N_503,N_494,N_424);
nand U504 (N_504,N_448,N_442);
and U505 (N_505,N_427,N_416);
and U506 (N_506,N_400,N_466);
or U507 (N_507,N_479,N_464);
or U508 (N_508,N_406,N_452);
or U509 (N_509,N_401,N_458);
and U510 (N_510,N_477,N_402);
and U511 (N_511,N_476,N_480);
nand U512 (N_512,N_440,N_426);
or U513 (N_513,N_407,N_498);
nand U514 (N_514,N_475,N_481);
or U515 (N_515,N_432,N_403);
and U516 (N_516,N_444,N_418);
or U517 (N_517,N_422,N_486);
nand U518 (N_518,N_437,N_430);
or U519 (N_519,N_445,N_492);
and U520 (N_520,N_409,N_443);
or U521 (N_521,N_439,N_462);
nor U522 (N_522,N_471,N_413);
or U523 (N_523,N_461,N_491);
nand U524 (N_524,N_499,N_436);
nand U525 (N_525,N_421,N_433);
nor U526 (N_526,N_425,N_497);
and U527 (N_527,N_455,N_482);
nor U528 (N_528,N_454,N_408);
and U529 (N_529,N_457,N_485);
nor U530 (N_530,N_419,N_493);
or U531 (N_531,N_465,N_447);
nor U532 (N_532,N_496,N_484);
nor U533 (N_533,N_410,N_434);
nor U534 (N_534,N_428,N_429);
nor U535 (N_535,N_472,N_474);
or U536 (N_536,N_463,N_423);
and U537 (N_537,N_473,N_459);
and U538 (N_538,N_488,N_446);
nand U539 (N_539,N_412,N_415);
or U540 (N_540,N_456,N_431);
nor U541 (N_541,N_490,N_489);
nor U542 (N_542,N_478,N_470);
or U543 (N_543,N_441,N_487);
nor U544 (N_544,N_460,N_420);
and U545 (N_545,N_449,N_451);
or U546 (N_546,N_468,N_483);
nor U547 (N_547,N_438,N_469);
and U548 (N_548,N_495,N_411);
nor U549 (N_549,N_450,N_404);
or U550 (N_550,N_455,N_470);
nand U551 (N_551,N_459,N_482);
or U552 (N_552,N_479,N_407);
nand U553 (N_553,N_495,N_484);
or U554 (N_554,N_449,N_459);
nand U555 (N_555,N_481,N_421);
nand U556 (N_556,N_414,N_433);
nor U557 (N_557,N_497,N_433);
and U558 (N_558,N_430,N_424);
nand U559 (N_559,N_457,N_404);
or U560 (N_560,N_410,N_457);
nor U561 (N_561,N_485,N_468);
nand U562 (N_562,N_463,N_419);
and U563 (N_563,N_471,N_410);
or U564 (N_564,N_433,N_408);
nor U565 (N_565,N_406,N_458);
and U566 (N_566,N_454,N_418);
nor U567 (N_567,N_438,N_463);
or U568 (N_568,N_415,N_465);
and U569 (N_569,N_475,N_449);
nand U570 (N_570,N_424,N_434);
and U571 (N_571,N_479,N_409);
nor U572 (N_572,N_433,N_411);
or U573 (N_573,N_414,N_446);
nor U574 (N_574,N_407,N_416);
nand U575 (N_575,N_428,N_456);
or U576 (N_576,N_403,N_407);
nand U577 (N_577,N_413,N_485);
or U578 (N_578,N_495,N_475);
nand U579 (N_579,N_443,N_415);
nor U580 (N_580,N_403,N_428);
nor U581 (N_581,N_413,N_497);
nand U582 (N_582,N_433,N_442);
nand U583 (N_583,N_406,N_429);
nand U584 (N_584,N_492,N_441);
nor U585 (N_585,N_421,N_459);
nor U586 (N_586,N_470,N_493);
nor U587 (N_587,N_415,N_470);
nand U588 (N_588,N_471,N_474);
or U589 (N_589,N_471,N_480);
nor U590 (N_590,N_418,N_435);
and U591 (N_591,N_480,N_415);
nor U592 (N_592,N_483,N_422);
and U593 (N_593,N_494,N_468);
xnor U594 (N_594,N_460,N_433);
and U595 (N_595,N_496,N_448);
or U596 (N_596,N_470,N_438);
nor U597 (N_597,N_458,N_439);
and U598 (N_598,N_467,N_488);
or U599 (N_599,N_473,N_406);
and U600 (N_600,N_562,N_517);
nand U601 (N_601,N_544,N_588);
xor U602 (N_602,N_583,N_599);
and U603 (N_603,N_530,N_592);
nand U604 (N_604,N_569,N_561);
nor U605 (N_605,N_507,N_548);
nor U606 (N_606,N_524,N_591);
or U607 (N_607,N_582,N_556);
nor U608 (N_608,N_564,N_539);
nor U609 (N_609,N_595,N_543);
nor U610 (N_610,N_594,N_545);
nand U611 (N_611,N_542,N_538);
and U612 (N_612,N_554,N_553);
or U613 (N_613,N_541,N_527);
or U614 (N_614,N_509,N_515);
or U615 (N_615,N_523,N_516);
nand U616 (N_616,N_536,N_597);
nor U617 (N_617,N_547,N_549);
or U618 (N_618,N_508,N_528);
or U619 (N_619,N_537,N_511);
nor U620 (N_620,N_574,N_560);
nor U621 (N_621,N_503,N_550);
and U622 (N_622,N_525,N_581);
or U623 (N_623,N_533,N_532);
nor U624 (N_624,N_555,N_577);
nor U625 (N_625,N_589,N_552);
nand U626 (N_626,N_534,N_519);
and U627 (N_627,N_522,N_535);
or U628 (N_628,N_518,N_573);
and U629 (N_629,N_558,N_586);
and U630 (N_630,N_578,N_563);
nor U631 (N_631,N_585,N_514);
and U632 (N_632,N_566,N_506);
nand U633 (N_633,N_593,N_584);
nor U634 (N_634,N_504,N_575);
nand U635 (N_635,N_513,N_526);
or U636 (N_636,N_598,N_531);
or U637 (N_637,N_502,N_510);
and U638 (N_638,N_546,N_557);
and U639 (N_639,N_540,N_551);
nand U640 (N_640,N_590,N_580);
and U641 (N_641,N_521,N_579);
nand U642 (N_642,N_587,N_520);
nor U643 (N_643,N_559,N_565);
and U644 (N_644,N_512,N_567);
or U645 (N_645,N_596,N_570);
nand U646 (N_646,N_505,N_568);
or U647 (N_647,N_529,N_501);
nor U648 (N_648,N_500,N_576);
nor U649 (N_649,N_572,N_571);
and U650 (N_650,N_580,N_506);
nor U651 (N_651,N_567,N_582);
and U652 (N_652,N_503,N_588);
or U653 (N_653,N_582,N_558);
nor U654 (N_654,N_555,N_512);
nand U655 (N_655,N_557,N_552);
or U656 (N_656,N_503,N_559);
or U657 (N_657,N_542,N_580);
nand U658 (N_658,N_533,N_510);
nor U659 (N_659,N_541,N_540);
nand U660 (N_660,N_518,N_531);
and U661 (N_661,N_575,N_583);
nor U662 (N_662,N_564,N_506);
nor U663 (N_663,N_573,N_581);
nor U664 (N_664,N_535,N_586);
nand U665 (N_665,N_509,N_528);
or U666 (N_666,N_506,N_548);
nor U667 (N_667,N_529,N_569);
nor U668 (N_668,N_562,N_540);
nand U669 (N_669,N_502,N_584);
nand U670 (N_670,N_598,N_589);
nand U671 (N_671,N_589,N_526);
nor U672 (N_672,N_503,N_509);
nand U673 (N_673,N_528,N_561);
and U674 (N_674,N_521,N_530);
and U675 (N_675,N_580,N_531);
nor U676 (N_676,N_521,N_558);
nand U677 (N_677,N_554,N_593);
nor U678 (N_678,N_532,N_587);
and U679 (N_679,N_504,N_592);
or U680 (N_680,N_518,N_538);
and U681 (N_681,N_542,N_514);
nor U682 (N_682,N_520,N_525);
nor U683 (N_683,N_527,N_519);
xor U684 (N_684,N_595,N_541);
and U685 (N_685,N_514,N_523);
nor U686 (N_686,N_562,N_594);
nand U687 (N_687,N_593,N_571);
or U688 (N_688,N_557,N_599);
nand U689 (N_689,N_501,N_558);
nand U690 (N_690,N_525,N_551);
and U691 (N_691,N_502,N_580);
nand U692 (N_692,N_551,N_591);
nor U693 (N_693,N_562,N_597);
nor U694 (N_694,N_509,N_507);
nand U695 (N_695,N_536,N_576);
and U696 (N_696,N_552,N_597);
nand U697 (N_697,N_523,N_542);
or U698 (N_698,N_529,N_568);
nand U699 (N_699,N_531,N_561);
and U700 (N_700,N_607,N_631);
nand U701 (N_701,N_686,N_619);
or U702 (N_702,N_637,N_674);
nand U703 (N_703,N_673,N_676);
nand U704 (N_704,N_697,N_687);
nand U705 (N_705,N_698,N_652);
or U706 (N_706,N_616,N_650);
nand U707 (N_707,N_618,N_634);
or U708 (N_708,N_683,N_656);
and U709 (N_709,N_608,N_612);
nor U710 (N_710,N_659,N_661);
nand U711 (N_711,N_672,N_633);
or U712 (N_712,N_691,N_694);
nor U713 (N_713,N_638,N_651);
or U714 (N_714,N_693,N_664);
or U715 (N_715,N_685,N_681);
or U716 (N_716,N_602,N_635);
and U717 (N_717,N_632,N_643);
nand U718 (N_718,N_665,N_626);
and U719 (N_719,N_614,N_645);
and U720 (N_720,N_613,N_670);
xor U721 (N_721,N_625,N_623);
and U722 (N_722,N_679,N_649);
and U723 (N_723,N_621,N_646);
nand U724 (N_724,N_636,N_688);
or U725 (N_725,N_699,N_690);
and U726 (N_726,N_678,N_641);
nand U727 (N_727,N_689,N_684);
nand U728 (N_728,N_629,N_604);
nor U729 (N_729,N_657,N_640);
nand U730 (N_730,N_671,N_677);
nand U731 (N_731,N_620,N_617);
nand U732 (N_732,N_695,N_644);
or U733 (N_733,N_655,N_639);
nor U734 (N_734,N_603,N_653);
nand U735 (N_735,N_611,N_669);
nor U736 (N_736,N_647,N_696);
or U737 (N_737,N_609,N_660);
or U738 (N_738,N_628,N_658);
and U739 (N_739,N_622,N_610);
and U740 (N_740,N_627,N_682);
nor U741 (N_741,N_630,N_675);
or U742 (N_742,N_667,N_624);
nand U743 (N_743,N_680,N_692);
nand U744 (N_744,N_615,N_666);
and U745 (N_745,N_601,N_668);
or U746 (N_746,N_648,N_600);
nand U747 (N_747,N_606,N_662);
nand U748 (N_748,N_663,N_654);
nor U749 (N_749,N_605,N_642);
and U750 (N_750,N_695,N_651);
nand U751 (N_751,N_642,N_606);
nand U752 (N_752,N_645,N_628);
or U753 (N_753,N_607,N_676);
xnor U754 (N_754,N_670,N_648);
or U755 (N_755,N_695,N_679);
and U756 (N_756,N_657,N_655);
nor U757 (N_757,N_676,N_654);
and U758 (N_758,N_616,N_622);
or U759 (N_759,N_630,N_649);
and U760 (N_760,N_680,N_613);
and U761 (N_761,N_647,N_691);
and U762 (N_762,N_627,N_694);
and U763 (N_763,N_611,N_622);
nor U764 (N_764,N_693,N_690);
nand U765 (N_765,N_683,N_615);
and U766 (N_766,N_646,N_663);
nand U767 (N_767,N_679,N_618);
xor U768 (N_768,N_600,N_641);
nand U769 (N_769,N_665,N_674);
nand U770 (N_770,N_638,N_673);
nor U771 (N_771,N_666,N_665);
nor U772 (N_772,N_633,N_621);
nand U773 (N_773,N_623,N_634);
or U774 (N_774,N_609,N_692);
and U775 (N_775,N_666,N_678);
and U776 (N_776,N_629,N_680);
nand U777 (N_777,N_696,N_607);
and U778 (N_778,N_652,N_604);
nor U779 (N_779,N_699,N_665);
nand U780 (N_780,N_673,N_608);
and U781 (N_781,N_651,N_614);
nor U782 (N_782,N_683,N_667);
nor U783 (N_783,N_638,N_672);
nor U784 (N_784,N_627,N_642);
or U785 (N_785,N_609,N_675);
and U786 (N_786,N_640,N_605);
and U787 (N_787,N_641,N_610);
nor U788 (N_788,N_666,N_663);
nand U789 (N_789,N_673,N_637);
xor U790 (N_790,N_639,N_644);
or U791 (N_791,N_699,N_630);
and U792 (N_792,N_683,N_687);
nor U793 (N_793,N_627,N_634);
or U794 (N_794,N_615,N_665);
and U795 (N_795,N_644,N_628);
nor U796 (N_796,N_626,N_696);
nand U797 (N_797,N_670,N_617);
or U798 (N_798,N_622,N_663);
nor U799 (N_799,N_657,N_613);
nand U800 (N_800,N_793,N_708);
nand U801 (N_801,N_755,N_736);
nor U802 (N_802,N_782,N_789);
xor U803 (N_803,N_728,N_723);
or U804 (N_804,N_750,N_764);
nand U805 (N_805,N_705,N_735);
and U806 (N_806,N_798,N_781);
and U807 (N_807,N_751,N_703);
and U808 (N_808,N_761,N_718);
or U809 (N_809,N_763,N_756);
nand U810 (N_810,N_715,N_720);
or U811 (N_811,N_706,N_709);
and U812 (N_812,N_775,N_722);
and U813 (N_813,N_730,N_743);
and U814 (N_814,N_727,N_719);
and U815 (N_815,N_776,N_739);
nor U816 (N_816,N_767,N_765);
nor U817 (N_817,N_740,N_790);
xor U818 (N_818,N_721,N_791);
nor U819 (N_819,N_794,N_734);
or U820 (N_820,N_712,N_766);
or U821 (N_821,N_757,N_738);
xor U822 (N_822,N_747,N_724);
or U823 (N_823,N_759,N_714);
xor U824 (N_824,N_783,N_742);
nor U825 (N_825,N_771,N_778);
nand U826 (N_826,N_774,N_741);
nand U827 (N_827,N_716,N_754);
nor U828 (N_828,N_758,N_770);
xnor U829 (N_829,N_786,N_762);
or U830 (N_830,N_784,N_737);
or U831 (N_831,N_769,N_745);
nand U832 (N_832,N_787,N_772);
or U833 (N_833,N_768,N_704);
nor U834 (N_834,N_701,N_773);
nand U835 (N_835,N_777,N_779);
xnor U836 (N_836,N_726,N_753);
and U837 (N_837,N_796,N_707);
and U838 (N_838,N_785,N_780);
or U839 (N_839,N_700,N_713);
nor U840 (N_840,N_799,N_788);
nor U841 (N_841,N_792,N_717);
and U842 (N_842,N_744,N_797);
nor U843 (N_843,N_711,N_752);
nor U844 (N_844,N_702,N_749);
or U845 (N_845,N_760,N_748);
and U846 (N_846,N_710,N_732);
nand U847 (N_847,N_746,N_729);
or U848 (N_848,N_795,N_731);
or U849 (N_849,N_725,N_733);
and U850 (N_850,N_779,N_798);
and U851 (N_851,N_719,N_782);
nor U852 (N_852,N_710,N_708);
or U853 (N_853,N_775,N_789);
and U854 (N_854,N_710,N_766);
or U855 (N_855,N_787,N_731);
nand U856 (N_856,N_796,N_772);
or U857 (N_857,N_786,N_744);
or U858 (N_858,N_722,N_768);
nand U859 (N_859,N_793,N_705);
and U860 (N_860,N_792,N_767);
and U861 (N_861,N_782,N_729);
nand U862 (N_862,N_742,N_751);
and U863 (N_863,N_759,N_744);
and U864 (N_864,N_744,N_795);
and U865 (N_865,N_762,N_787);
nor U866 (N_866,N_730,N_719);
and U867 (N_867,N_795,N_735);
or U868 (N_868,N_771,N_798);
nand U869 (N_869,N_753,N_712);
nor U870 (N_870,N_734,N_799);
xor U871 (N_871,N_767,N_743);
xnor U872 (N_872,N_776,N_771);
or U873 (N_873,N_768,N_721);
or U874 (N_874,N_775,N_794);
nand U875 (N_875,N_711,N_748);
and U876 (N_876,N_729,N_794);
or U877 (N_877,N_777,N_780);
and U878 (N_878,N_788,N_768);
nor U879 (N_879,N_754,N_729);
or U880 (N_880,N_716,N_731);
nand U881 (N_881,N_740,N_752);
nor U882 (N_882,N_791,N_719);
nand U883 (N_883,N_737,N_789);
nor U884 (N_884,N_782,N_772);
nand U885 (N_885,N_707,N_749);
or U886 (N_886,N_772,N_771);
nor U887 (N_887,N_747,N_774);
nor U888 (N_888,N_746,N_706);
nand U889 (N_889,N_727,N_799);
and U890 (N_890,N_779,N_706);
nor U891 (N_891,N_780,N_773);
nor U892 (N_892,N_769,N_792);
or U893 (N_893,N_728,N_715);
nand U894 (N_894,N_783,N_763);
and U895 (N_895,N_776,N_782);
nor U896 (N_896,N_724,N_752);
nor U897 (N_897,N_760,N_753);
nor U898 (N_898,N_780,N_751);
nor U899 (N_899,N_774,N_772);
nor U900 (N_900,N_841,N_877);
or U901 (N_901,N_813,N_819);
or U902 (N_902,N_894,N_859);
or U903 (N_903,N_838,N_829);
and U904 (N_904,N_863,N_897);
or U905 (N_905,N_816,N_846);
nand U906 (N_906,N_873,N_839);
and U907 (N_907,N_888,N_832);
nand U908 (N_908,N_810,N_896);
nand U909 (N_909,N_817,N_870);
and U910 (N_910,N_895,N_802);
or U911 (N_911,N_872,N_854);
nand U912 (N_912,N_828,N_861);
nor U913 (N_913,N_853,N_801);
nor U914 (N_914,N_822,N_883);
nor U915 (N_915,N_833,N_857);
nor U916 (N_916,N_837,N_890);
nor U917 (N_917,N_821,N_809);
nand U918 (N_918,N_805,N_834);
nand U919 (N_919,N_862,N_899);
nor U920 (N_920,N_858,N_885);
nand U921 (N_921,N_893,N_812);
nand U922 (N_922,N_827,N_820);
nand U923 (N_923,N_845,N_851);
nand U924 (N_924,N_880,N_878);
nor U925 (N_925,N_825,N_835);
xor U926 (N_926,N_867,N_865);
and U927 (N_927,N_881,N_823);
xor U928 (N_928,N_855,N_876);
and U929 (N_929,N_842,N_814);
nor U930 (N_930,N_844,N_874);
nor U931 (N_931,N_850,N_889);
nor U932 (N_932,N_892,N_868);
and U933 (N_933,N_800,N_818);
nor U934 (N_934,N_887,N_840);
and U935 (N_935,N_831,N_898);
and U936 (N_936,N_856,N_866);
or U937 (N_937,N_879,N_826);
nor U938 (N_938,N_824,N_852);
nor U939 (N_939,N_811,N_804);
or U940 (N_940,N_836,N_808);
or U941 (N_941,N_843,N_807);
nand U942 (N_942,N_860,N_849);
nand U943 (N_943,N_847,N_830);
nor U944 (N_944,N_864,N_803);
or U945 (N_945,N_882,N_806);
or U946 (N_946,N_871,N_815);
or U947 (N_947,N_886,N_869);
and U948 (N_948,N_848,N_875);
or U949 (N_949,N_891,N_884);
nor U950 (N_950,N_809,N_857);
or U951 (N_951,N_805,N_886);
and U952 (N_952,N_872,N_865);
nor U953 (N_953,N_890,N_832);
nand U954 (N_954,N_831,N_872);
and U955 (N_955,N_856,N_813);
and U956 (N_956,N_835,N_809);
xor U957 (N_957,N_810,N_806);
or U958 (N_958,N_825,N_870);
nor U959 (N_959,N_840,N_802);
nand U960 (N_960,N_874,N_885);
nor U961 (N_961,N_832,N_889);
and U962 (N_962,N_825,N_848);
and U963 (N_963,N_855,N_856);
nand U964 (N_964,N_802,N_827);
nand U965 (N_965,N_811,N_814);
nand U966 (N_966,N_819,N_816);
nand U967 (N_967,N_898,N_825);
xnor U968 (N_968,N_898,N_848);
or U969 (N_969,N_834,N_877);
nand U970 (N_970,N_842,N_804);
nor U971 (N_971,N_819,N_824);
or U972 (N_972,N_878,N_809);
and U973 (N_973,N_840,N_829);
nand U974 (N_974,N_845,N_816);
and U975 (N_975,N_844,N_892);
and U976 (N_976,N_838,N_832);
nor U977 (N_977,N_877,N_859);
and U978 (N_978,N_849,N_816);
nor U979 (N_979,N_846,N_847);
nor U980 (N_980,N_897,N_810);
nor U981 (N_981,N_886,N_883);
and U982 (N_982,N_871,N_897);
nand U983 (N_983,N_844,N_899);
or U984 (N_984,N_834,N_803);
nor U985 (N_985,N_820,N_872);
nor U986 (N_986,N_839,N_875);
or U987 (N_987,N_820,N_839);
nor U988 (N_988,N_847,N_837);
or U989 (N_989,N_827,N_891);
nand U990 (N_990,N_861,N_848);
nand U991 (N_991,N_890,N_889);
nand U992 (N_992,N_829,N_817);
nor U993 (N_993,N_837,N_844);
and U994 (N_994,N_810,N_817);
nor U995 (N_995,N_889,N_873);
nor U996 (N_996,N_838,N_828);
and U997 (N_997,N_840,N_807);
nand U998 (N_998,N_882,N_864);
or U999 (N_999,N_820,N_891);
or U1000 (N_1000,N_914,N_971);
nand U1001 (N_1001,N_919,N_922);
nor U1002 (N_1002,N_954,N_900);
or U1003 (N_1003,N_952,N_959);
or U1004 (N_1004,N_988,N_964);
and U1005 (N_1005,N_985,N_918);
nor U1006 (N_1006,N_925,N_906);
nand U1007 (N_1007,N_960,N_938);
nand U1008 (N_1008,N_904,N_937);
or U1009 (N_1009,N_981,N_902);
nor U1010 (N_1010,N_977,N_956);
nor U1011 (N_1011,N_991,N_982);
or U1012 (N_1012,N_984,N_989);
xnor U1013 (N_1013,N_951,N_963);
nand U1014 (N_1014,N_903,N_908);
and U1015 (N_1015,N_910,N_943);
and U1016 (N_1016,N_934,N_999);
nor U1017 (N_1017,N_940,N_912);
and U1018 (N_1018,N_987,N_969);
or U1019 (N_1019,N_945,N_929);
nor U1020 (N_1020,N_920,N_993);
nor U1021 (N_1021,N_973,N_974);
or U1022 (N_1022,N_979,N_970);
or U1023 (N_1023,N_961,N_953);
nand U1024 (N_1024,N_928,N_965);
and U1025 (N_1025,N_976,N_916);
xor U1026 (N_1026,N_930,N_966);
and U1027 (N_1027,N_913,N_932);
and U1028 (N_1028,N_923,N_915);
nor U1029 (N_1029,N_983,N_975);
and U1030 (N_1030,N_911,N_990);
and U1031 (N_1031,N_997,N_962);
or U1032 (N_1032,N_927,N_967);
nor U1033 (N_1033,N_907,N_931);
nor U1034 (N_1034,N_992,N_972);
nand U1035 (N_1035,N_950,N_958);
or U1036 (N_1036,N_968,N_994);
nand U1037 (N_1037,N_998,N_955);
or U1038 (N_1038,N_978,N_924);
and U1039 (N_1039,N_980,N_926);
nor U1040 (N_1040,N_995,N_996);
nand U1041 (N_1041,N_949,N_942);
or U1042 (N_1042,N_939,N_947);
nand U1043 (N_1043,N_905,N_944);
and U1044 (N_1044,N_941,N_957);
and U1045 (N_1045,N_933,N_909);
or U1046 (N_1046,N_935,N_917);
and U1047 (N_1047,N_948,N_921);
or U1048 (N_1048,N_936,N_901);
nand U1049 (N_1049,N_986,N_946);
and U1050 (N_1050,N_973,N_903);
nor U1051 (N_1051,N_900,N_920);
or U1052 (N_1052,N_939,N_938);
nor U1053 (N_1053,N_966,N_968);
xor U1054 (N_1054,N_972,N_924);
nor U1055 (N_1055,N_964,N_962);
or U1056 (N_1056,N_933,N_934);
or U1057 (N_1057,N_951,N_985);
and U1058 (N_1058,N_906,N_996);
nor U1059 (N_1059,N_913,N_942);
nor U1060 (N_1060,N_967,N_929);
nand U1061 (N_1061,N_999,N_928);
nand U1062 (N_1062,N_915,N_929);
nor U1063 (N_1063,N_978,N_918);
nand U1064 (N_1064,N_979,N_902);
nor U1065 (N_1065,N_953,N_994);
and U1066 (N_1066,N_954,N_901);
nand U1067 (N_1067,N_909,N_981);
and U1068 (N_1068,N_950,N_978);
nand U1069 (N_1069,N_987,N_955);
nand U1070 (N_1070,N_935,N_951);
or U1071 (N_1071,N_974,N_927);
or U1072 (N_1072,N_966,N_919);
and U1073 (N_1073,N_974,N_941);
nor U1074 (N_1074,N_999,N_954);
nor U1075 (N_1075,N_977,N_940);
or U1076 (N_1076,N_965,N_903);
or U1077 (N_1077,N_918,N_912);
or U1078 (N_1078,N_927,N_952);
or U1079 (N_1079,N_971,N_957);
nor U1080 (N_1080,N_955,N_937);
or U1081 (N_1081,N_930,N_927);
nor U1082 (N_1082,N_956,N_924);
nor U1083 (N_1083,N_994,N_942);
nand U1084 (N_1084,N_974,N_995);
nand U1085 (N_1085,N_927,N_909);
or U1086 (N_1086,N_901,N_942);
nand U1087 (N_1087,N_917,N_910);
or U1088 (N_1088,N_984,N_993);
or U1089 (N_1089,N_990,N_901);
nand U1090 (N_1090,N_991,N_970);
or U1091 (N_1091,N_971,N_966);
or U1092 (N_1092,N_928,N_903);
and U1093 (N_1093,N_929,N_913);
nor U1094 (N_1094,N_912,N_964);
nand U1095 (N_1095,N_930,N_929);
nor U1096 (N_1096,N_987,N_918);
nor U1097 (N_1097,N_917,N_959);
and U1098 (N_1098,N_913,N_916);
and U1099 (N_1099,N_925,N_958);
and U1100 (N_1100,N_1036,N_1071);
nor U1101 (N_1101,N_1058,N_1009);
or U1102 (N_1102,N_1012,N_1039);
and U1103 (N_1103,N_1018,N_1049);
or U1104 (N_1104,N_1003,N_1042);
nand U1105 (N_1105,N_1079,N_1059);
nand U1106 (N_1106,N_1043,N_1019);
or U1107 (N_1107,N_1061,N_1027);
and U1108 (N_1108,N_1002,N_1052);
nor U1109 (N_1109,N_1090,N_1053);
or U1110 (N_1110,N_1044,N_1066);
or U1111 (N_1111,N_1099,N_1074);
and U1112 (N_1112,N_1089,N_1023);
nand U1113 (N_1113,N_1087,N_1032);
or U1114 (N_1114,N_1047,N_1054);
and U1115 (N_1115,N_1062,N_1063);
nor U1116 (N_1116,N_1038,N_1091);
nand U1117 (N_1117,N_1035,N_1085);
nor U1118 (N_1118,N_1057,N_1028);
nand U1119 (N_1119,N_1065,N_1072);
nor U1120 (N_1120,N_1026,N_1021);
and U1121 (N_1121,N_1006,N_1051);
nand U1122 (N_1122,N_1075,N_1076);
nand U1123 (N_1123,N_1025,N_1082);
and U1124 (N_1124,N_1073,N_1095);
or U1125 (N_1125,N_1093,N_1060);
and U1126 (N_1126,N_1098,N_1040);
or U1127 (N_1127,N_1050,N_1094);
nand U1128 (N_1128,N_1068,N_1022);
nand U1129 (N_1129,N_1092,N_1004);
nand U1130 (N_1130,N_1015,N_1014);
or U1131 (N_1131,N_1010,N_1046);
nor U1132 (N_1132,N_1077,N_1048);
nor U1133 (N_1133,N_1080,N_1037);
or U1134 (N_1134,N_1017,N_1086);
and U1135 (N_1135,N_1083,N_1078);
nor U1136 (N_1136,N_1041,N_1056);
xnor U1137 (N_1137,N_1005,N_1001);
and U1138 (N_1138,N_1029,N_1088);
nand U1139 (N_1139,N_1097,N_1011);
nand U1140 (N_1140,N_1034,N_1084);
and U1141 (N_1141,N_1070,N_1033);
or U1142 (N_1142,N_1024,N_1096);
and U1143 (N_1143,N_1031,N_1069);
and U1144 (N_1144,N_1030,N_1020);
or U1145 (N_1145,N_1007,N_1064);
or U1146 (N_1146,N_1045,N_1008);
or U1147 (N_1147,N_1067,N_1013);
and U1148 (N_1148,N_1016,N_1055);
nand U1149 (N_1149,N_1000,N_1081);
or U1150 (N_1150,N_1098,N_1069);
or U1151 (N_1151,N_1074,N_1014);
or U1152 (N_1152,N_1064,N_1079);
nor U1153 (N_1153,N_1054,N_1033);
and U1154 (N_1154,N_1005,N_1061);
and U1155 (N_1155,N_1081,N_1091);
or U1156 (N_1156,N_1033,N_1098);
and U1157 (N_1157,N_1009,N_1028);
nor U1158 (N_1158,N_1014,N_1063);
nand U1159 (N_1159,N_1002,N_1042);
nand U1160 (N_1160,N_1042,N_1050);
and U1161 (N_1161,N_1081,N_1006);
nand U1162 (N_1162,N_1037,N_1075);
or U1163 (N_1163,N_1067,N_1036);
nor U1164 (N_1164,N_1077,N_1039);
nor U1165 (N_1165,N_1093,N_1037);
and U1166 (N_1166,N_1094,N_1064);
or U1167 (N_1167,N_1024,N_1003);
nand U1168 (N_1168,N_1095,N_1056);
or U1169 (N_1169,N_1049,N_1024);
and U1170 (N_1170,N_1080,N_1079);
nor U1171 (N_1171,N_1030,N_1060);
or U1172 (N_1172,N_1021,N_1046);
nor U1173 (N_1173,N_1085,N_1060);
and U1174 (N_1174,N_1086,N_1030);
nand U1175 (N_1175,N_1090,N_1020);
or U1176 (N_1176,N_1084,N_1050);
and U1177 (N_1177,N_1033,N_1088);
or U1178 (N_1178,N_1033,N_1028);
nand U1179 (N_1179,N_1050,N_1048);
nand U1180 (N_1180,N_1048,N_1091);
nor U1181 (N_1181,N_1080,N_1066);
and U1182 (N_1182,N_1075,N_1094);
nand U1183 (N_1183,N_1027,N_1080);
and U1184 (N_1184,N_1016,N_1039);
or U1185 (N_1185,N_1005,N_1097);
nor U1186 (N_1186,N_1022,N_1039);
and U1187 (N_1187,N_1025,N_1013);
or U1188 (N_1188,N_1075,N_1062);
nor U1189 (N_1189,N_1038,N_1033);
nor U1190 (N_1190,N_1088,N_1080);
nor U1191 (N_1191,N_1054,N_1080);
nor U1192 (N_1192,N_1054,N_1072);
and U1193 (N_1193,N_1018,N_1098);
nor U1194 (N_1194,N_1022,N_1036);
or U1195 (N_1195,N_1001,N_1030);
nor U1196 (N_1196,N_1026,N_1071);
nor U1197 (N_1197,N_1034,N_1047);
nor U1198 (N_1198,N_1051,N_1046);
nor U1199 (N_1199,N_1047,N_1072);
nand U1200 (N_1200,N_1163,N_1177);
xor U1201 (N_1201,N_1199,N_1176);
nor U1202 (N_1202,N_1148,N_1184);
and U1203 (N_1203,N_1182,N_1164);
or U1204 (N_1204,N_1193,N_1105);
nor U1205 (N_1205,N_1112,N_1131);
or U1206 (N_1206,N_1165,N_1135);
and U1207 (N_1207,N_1140,N_1126);
nor U1208 (N_1208,N_1189,N_1120);
and U1209 (N_1209,N_1158,N_1139);
or U1210 (N_1210,N_1116,N_1117);
nor U1211 (N_1211,N_1128,N_1124);
nor U1212 (N_1212,N_1153,N_1188);
and U1213 (N_1213,N_1143,N_1191);
nand U1214 (N_1214,N_1181,N_1194);
or U1215 (N_1215,N_1113,N_1161);
nor U1216 (N_1216,N_1154,N_1168);
and U1217 (N_1217,N_1170,N_1162);
and U1218 (N_1218,N_1137,N_1108);
nand U1219 (N_1219,N_1109,N_1149);
and U1220 (N_1220,N_1174,N_1145);
nand U1221 (N_1221,N_1147,N_1185);
nand U1222 (N_1222,N_1133,N_1198);
or U1223 (N_1223,N_1125,N_1169);
nor U1224 (N_1224,N_1192,N_1102);
or U1225 (N_1225,N_1142,N_1138);
or U1226 (N_1226,N_1160,N_1107);
nor U1227 (N_1227,N_1106,N_1151);
or U1228 (N_1228,N_1118,N_1127);
nor U1229 (N_1229,N_1103,N_1197);
or U1230 (N_1230,N_1155,N_1175);
or U1231 (N_1231,N_1119,N_1171);
or U1232 (N_1232,N_1183,N_1178);
nor U1233 (N_1233,N_1132,N_1152);
nor U1234 (N_1234,N_1123,N_1150);
nor U1235 (N_1235,N_1144,N_1195);
or U1236 (N_1236,N_1159,N_1179);
nand U1237 (N_1237,N_1129,N_1141);
or U1238 (N_1238,N_1101,N_1122);
nand U1239 (N_1239,N_1190,N_1115);
nor U1240 (N_1240,N_1104,N_1130);
and U1241 (N_1241,N_1136,N_1173);
and U1242 (N_1242,N_1196,N_1187);
nor U1243 (N_1243,N_1172,N_1121);
nand U1244 (N_1244,N_1167,N_1110);
xor U1245 (N_1245,N_1157,N_1186);
or U1246 (N_1246,N_1156,N_1114);
nand U1247 (N_1247,N_1180,N_1134);
nor U1248 (N_1248,N_1146,N_1166);
or U1249 (N_1249,N_1100,N_1111);
or U1250 (N_1250,N_1112,N_1198);
xor U1251 (N_1251,N_1154,N_1142);
nand U1252 (N_1252,N_1198,N_1127);
and U1253 (N_1253,N_1111,N_1150);
and U1254 (N_1254,N_1126,N_1188);
and U1255 (N_1255,N_1145,N_1177);
or U1256 (N_1256,N_1167,N_1135);
nor U1257 (N_1257,N_1141,N_1114);
nor U1258 (N_1258,N_1194,N_1165);
or U1259 (N_1259,N_1109,N_1148);
and U1260 (N_1260,N_1131,N_1192);
or U1261 (N_1261,N_1112,N_1101);
or U1262 (N_1262,N_1184,N_1185);
or U1263 (N_1263,N_1165,N_1143);
nand U1264 (N_1264,N_1139,N_1103);
or U1265 (N_1265,N_1110,N_1140);
nand U1266 (N_1266,N_1173,N_1130);
nand U1267 (N_1267,N_1169,N_1132);
and U1268 (N_1268,N_1153,N_1116);
nand U1269 (N_1269,N_1168,N_1102);
or U1270 (N_1270,N_1194,N_1186);
nand U1271 (N_1271,N_1188,N_1194);
and U1272 (N_1272,N_1171,N_1160);
nor U1273 (N_1273,N_1147,N_1103);
and U1274 (N_1274,N_1171,N_1193);
or U1275 (N_1275,N_1164,N_1120);
or U1276 (N_1276,N_1114,N_1116);
nand U1277 (N_1277,N_1113,N_1159);
nand U1278 (N_1278,N_1161,N_1189);
and U1279 (N_1279,N_1169,N_1117);
nor U1280 (N_1280,N_1191,N_1182);
or U1281 (N_1281,N_1142,N_1197);
nand U1282 (N_1282,N_1102,N_1133);
nor U1283 (N_1283,N_1111,N_1127);
and U1284 (N_1284,N_1150,N_1107);
and U1285 (N_1285,N_1194,N_1124);
and U1286 (N_1286,N_1138,N_1139);
or U1287 (N_1287,N_1131,N_1193);
nor U1288 (N_1288,N_1132,N_1108);
nor U1289 (N_1289,N_1189,N_1187);
or U1290 (N_1290,N_1127,N_1190);
and U1291 (N_1291,N_1142,N_1124);
nand U1292 (N_1292,N_1186,N_1120);
nand U1293 (N_1293,N_1193,N_1117);
nor U1294 (N_1294,N_1190,N_1104);
and U1295 (N_1295,N_1131,N_1194);
and U1296 (N_1296,N_1139,N_1118);
nand U1297 (N_1297,N_1119,N_1128);
and U1298 (N_1298,N_1175,N_1108);
and U1299 (N_1299,N_1151,N_1104);
or U1300 (N_1300,N_1298,N_1220);
and U1301 (N_1301,N_1242,N_1213);
or U1302 (N_1302,N_1279,N_1227);
or U1303 (N_1303,N_1225,N_1273);
or U1304 (N_1304,N_1212,N_1297);
nand U1305 (N_1305,N_1202,N_1214);
and U1306 (N_1306,N_1271,N_1266);
and U1307 (N_1307,N_1296,N_1267);
nand U1308 (N_1308,N_1243,N_1253);
and U1309 (N_1309,N_1265,N_1247);
or U1310 (N_1310,N_1275,N_1291);
nor U1311 (N_1311,N_1250,N_1223);
nor U1312 (N_1312,N_1260,N_1224);
xnor U1313 (N_1313,N_1238,N_1240);
and U1314 (N_1314,N_1234,N_1210);
or U1315 (N_1315,N_1219,N_1264);
and U1316 (N_1316,N_1285,N_1204);
nand U1317 (N_1317,N_1235,N_1241);
nand U1318 (N_1318,N_1277,N_1228);
nor U1319 (N_1319,N_1274,N_1278);
and U1320 (N_1320,N_1248,N_1269);
or U1321 (N_1321,N_1268,N_1226);
or U1322 (N_1322,N_1231,N_1292);
and U1323 (N_1323,N_1254,N_1258);
and U1324 (N_1324,N_1205,N_1282);
or U1325 (N_1325,N_1259,N_1262);
or U1326 (N_1326,N_1209,N_1289);
or U1327 (N_1327,N_1290,N_1272);
or U1328 (N_1328,N_1263,N_1201);
xnor U1329 (N_1329,N_1221,N_1233);
and U1330 (N_1330,N_1257,N_1270);
nor U1331 (N_1331,N_1200,N_1208);
or U1332 (N_1332,N_1288,N_1244);
nor U1333 (N_1333,N_1256,N_1239);
or U1334 (N_1334,N_1249,N_1237);
nor U1335 (N_1335,N_1218,N_1207);
nor U1336 (N_1336,N_1280,N_1217);
nor U1337 (N_1337,N_1211,N_1229);
nand U1338 (N_1338,N_1276,N_1255);
or U1339 (N_1339,N_1245,N_1252);
or U1340 (N_1340,N_1203,N_1230);
and U1341 (N_1341,N_1215,N_1251);
nand U1342 (N_1342,N_1283,N_1281);
and U1343 (N_1343,N_1286,N_1287);
nor U1344 (N_1344,N_1294,N_1299);
and U1345 (N_1345,N_1216,N_1295);
nand U1346 (N_1346,N_1236,N_1232);
xor U1347 (N_1347,N_1261,N_1284);
xor U1348 (N_1348,N_1246,N_1206);
and U1349 (N_1349,N_1293,N_1222);
nor U1350 (N_1350,N_1214,N_1247);
xnor U1351 (N_1351,N_1243,N_1203);
nor U1352 (N_1352,N_1268,N_1235);
nor U1353 (N_1353,N_1225,N_1260);
or U1354 (N_1354,N_1280,N_1290);
nand U1355 (N_1355,N_1292,N_1202);
and U1356 (N_1356,N_1275,N_1235);
nand U1357 (N_1357,N_1227,N_1283);
nor U1358 (N_1358,N_1212,N_1226);
or U1359 (N_1359,N_1245,N_1237);
and U1360 (N_1360,N_1220,N_1211);
and U1361 (N_1361,N_1220,N_1226);
and U1362 (N_1362,N_1268,N_1237);
or U1363 (N_1363,N_1263,N_1271);
or U1364 (N_1364,N_1232,N_1216);
or U1365 (N_1365,N_1231,N_1264);
nand U1366 (N_1366,N_1291,N_1210);
nand U1367 (N_1367,N_1292,N_1297);
nand U1368 (N_1368,N_1207,N_1282);
or U1369 (N_1369,N_1279,N_1208);
or U1370 (N_1370,N_1230,N_1210);
nand U1371 (N_1371,N_1212,N_1251);
and U1372 (N_1372,N_1267,N_1206);
or U1373 (N_1373,N_1266,N_1219);
nor U1374 (N_1374,N_1259,N_1226);
nand U1375 (N_1375,N_1201,N_1245);
or U1376 (N_1376,N_1266,N_1250);
nor U1377 (N_1377,N_1295,N_1298);
nand U1378 (N_1378,N_1289,N_1201);
nor U1379 (N_1379,N_1209,N_1275);
or U1380 (N_1380,N_1272,N_1252);
and U1381 (N_1381,N_1289,N_1224);
or U1382 (N_1382,N_1273,N_1218);
or U1383 (N_1383,N_1200,N_1262);
nand U1384 (N_1384,N_1248,N_1284);
and U1385 (N_1385,N_1278,N_1212);
and U1386 (N_1386,N_1236,N_1237);
nor U1387 (N_1387,N_1232,N_1257);
nand U1388 (N_1388,N_1280,N_1238);
nor U1389 (N_1389,N_1212,N_1236);
or U1390 (N_1390,N_1255,N_1266);
or U1391 (N_1391,N_1285,N_1279);
nand U1392 (N_1392,N_1284,N_1281);
nor U1393 (N_1393,N_1298,N_1297);
nand U1394 (N_1394,N_1238,N_1290);
nor U1395 (N_1395,N_1243,N_1216);
nand U1396 (N_1396,N_1211,N_1287);
and U1397 (N_1397,N_1267,N_1234);
or U1398 (N_1398,N_1208,N_1265);
nor U1399 (N_1399,N_1204,N_1289);
or U1400 (N_1400,N_1325,N_1314);
nand U1401 (N_1401,N_1359,N_1357);
nor U1402 (N_1402,N_1385,N_1381);
nor U1403 (N_1403,N_1316,N_1305);
nand U1404 (N_1404,N_1354,N_1344);
nand U1405 (N_1405,N_1343,N_1345);
and U1406 (N_1406,N_1347,N_1317);
nor U1407 (N_1407,N_1307,N_1389);
nand U1408 (N_1408,N_1304,N_1320);
nor U1409 (N_1409,N_1391,N_1348);
and U1410 (N_1410,N_1332,N_1378);
and U1411 (N_1411,N_1399,N_1319);
xnor U1412 (N_1412,N_1318,N_1342);
and U1413 (N_1413,N_1383,N_1312);
nand U1414 (N_1414,N_1392,N_1313);
and U1415 (N_1415,N_1361,N_1376);
and U1416 (N_1416,N_1300,N_1339);
nand U1417 (N_1417,N_1355,N_1368);
nand U1418 (N_1418,N_1302,N_1323);
nand U1419 (N_1419,N_1337,N_1321);
nand U1420 (N_1420,N_1340,N_1334);
nor U1421 (N_1421,N_1366,N_1328);
and U1422 (N_1422,N_1309,N_1322);
and U1423 (N_1423,N_1333,N_1379);
and U1424 (N_1424,N_1353,N_1352);
or U1425 (N_1425,N_1371,N_1356);
nor U1426 (N_1426,N_1370,N_1303);
nor U1427 (N_1427,N_1324,N_1384);
xor U1428 (N_1428,N_1349,N_1346);
and U1429 (N_1429,N_1335,N_1393);
nor U1430 (N_1430,N_1308,N_1397);
and U1431 (N_1431,N_1375,N_1358);
nand U1432 (N_1432,N_1377,N_1311);
or U1433 (N_1433,N_1380,N_1398);
and U1434 (N_1434,N_1327,N_1351);
nand U1435 (N_1435,N_1326,N_1374);
and U1436 (N_1436,N_1310,N_1336);
or U1437 (N_1437,N_1395,N_1341);
or U1438 (N_1438,N_1363,N_1372);
nor U1439 (N_1439,N_1331,N_1364);
and U1440 (N_1440,N_1338,N_1301);
or U1441 (N_1441,N_1350,N_1365);
nand U1442 (N_1442,N_1369,N_1390);
and U1443 (N_1443,N_1387,N_1373);
nor U1444 (N_1444,N_1306,N_1382);
nand U1445 (N_1445,N_1362,N_1386);
and U1446 (N_1446,N_1330,N_1388);
nand U1447 (N_1447,N_1396,N_1360);
and U1448 (N_1448,N_1329,N_1367);
and U1449 (N_1449,N_1394,N_1315);
and U1450 (N_1450,N_1382,N_1319);
nor U1451 (N_1451,N_1393,N_1319);
nor U1452 (N_1452,N_1371,N_1308);
nand U1453 (N_1453,N_1307,N_1342);
nor U1454 (N_1454,N_1365,N_1328);
nand U1455 (N_1455,N_1373,N_1344);
xor U1456 (N_1456,N_1394,N_1317);
xnor U1457 (N_1457,N_1302,N_1393);
nand U1458 (N_1458,N_1325,N_1316);
and U1459 (N_1459,N_1355,N_1345);
or U1460 (N_1460,N_1381,N_1375);
nand U1461 (N_1461,N_1322,N_1396);
or U1462 (N_1462,N_1393,N_1382);
and U1463 (N_1463,N_1346,N_1318);
xor U1464 (N_1464,N_1323,N_1318);
or U1465 (N_1465,N_1349,N_1372);
and U1466 (N_1466,N_1393,N_1380);
xor U1467 (N_1467,N_1373,N_1330);
nand U1468 (N_1468,N_1365,N_1390);
or U1469 (N_1469,N_1320,N_1360);
or U1470 (N_1470,N_1389,N_1314);
nor U1471 (N_1471,N_1338,N_1307);
nand U1472 (N_1472,N_1300,N_1399);
nor U1473 (N_1473,N_1378,N_1368);
nor U1474 (N_1474,N_1324,N_1382);
nand U1475 (N_1475,N_1378,N_1349);
nand U1476 (N_1476,N_1393,N_1369);
nor U1477 (N_1477,N_1335,N_1361);
or U1478 (N_1478,N_1329,N_1391);
or U1479 (N_1479,N_1310,N_1369);
nand U1480 (N_1480,N_1357,N_1354);
and U1481 (N_1481,N_1316,N_1306);
nand U1482 (N_1482,N_1335,N_1369);
or U1483 (N_1483,N_1392,N_1382);
and U1484 (N_1484,N_1356,N_1397);
nand U1485 (N_1485,N_1387,N_1349);
nand U1486 (N_1486,N_1387,N_1319);
nor U1487 (N_1487,N_1348,N_1356);
nand U1488 (N_1488,N_1372,N_1344);
and U1489 (N_1489,N_1348,N_1305);
and U1490 (N_1490,N_1330,N_1348);
nand U1491 (N_1491,N_1316,N_1382);
nor U1492 (N_1492,N_1338,N_1319);
and U1493 (N_1493,N_1372,N_1314);
nand U1494 (N_1494,N_1377,N_1367);
and U1495 (N_1495,N_1350,N_1382);
and U1496 (N_1496,N_1357,N_1317);
nand U1497 (N_1497,N_1376,N_1355);
nand U1498 (N_1498,N_1330,N_1334);
or U1499 (N_1499,N_1327,N_1334);
or U1500 (N_1500,N_1455,N_1459);
nand U1501 (N_1501,N_1418,N_1400);
xnor U1502 (N_1502,N_1488,N_1443);
or U1503 (N_1503,N_1444,N_1402);
and U1504 (N_1504,N_1433,N_1463);
nand U1505 (N_1505,N_1496,N_1493);
or U1506 (N_1506,N_1422,N_1431);
or U1507 (N_1507,N_1419,N_1439);
or U1508 (N_1508,N_1435,N_1489);
nand U1509 (N_1509,N_1448,N_1407);
or U1510 (N_1510,N_1420,N_1413);
nor U1511 (N_1511,N_1470,N_1414);
nand U1512 (N_1512,N_1412,N_1456);
and U1513 (N_1513,N_1475,N_1458);
and U1514 (N_1514,N_1410,N_1424);
nand U1515 (N_1515,N_1405,N_1490);
nand U1516 (N_1516,N_1482,N_1478);
and U1517 (N_1517,N_1468,N_1401);
nand U1518 (N_1518,N_1461,N_1462);
nor U1519 (N_1519,N_1440,N_1421);
and U1520 (N_1520,N_1471,N_1426);
and U1521 (N_1521,N_1434,N_1449);
and U1522 (N_1522,N_1497,N_1445);
nor U1523 (N_1523,N_1408,N_1432);
or U1524 (N_1524,N_1442,N_1466);
and U1525 (N_1525,N_1423,N_1452);
and U1526 (N_1526,N_1465,N_1403);
and U1527 (N_1527,N_1483,N_1450);
and U1528 (N_1528,N_1474,N_1467);
and U1529 (N_1529,N_1409,N_1469);
and U1530 (N_1530,N_1486,N_1484);
or U1531 (N_1531,N_1457,N_1441);
or U1532 (N_1532,N_1411,N_1480);
nand U1533 (N_1533,N_1430,N_1417);
and U1534 (N_1534,N_1476,N_1473);
nor U1535 (N_1535,N_1472,N_1487);
nand U1536 (N_1536,N_1429,N_1436);
nor U1537 (N_1537,N_1477,N_1427);
and U1538 (N_1538,N_1479,N_1499);
or U1539 (N_1539,N_1454,N_1437);
nor U1540 (N_1540,N_1428,N_1447);
nand U1541 (N_1541,N_1481,N_1495);
nand U1542 (N_1542,N_1453,N_1498);
or U1543 (N_1543,N_1415,N_1494);
nor U1544 (N_1544,N_1460,N_1491);
nand U1545 (N_1545,N_1446,N_1485);
nand U1546 (N_1546,N_1451,N_1492);
or U1547 (N_1547,N_1425,N_1404);
nand U1548 (N_1548,N_1464,N_1406);
nand U1549 (N_1549,N_1438,N_1416);
nor U1550 (N_1550,N_1413,N_1446);
and U1551 (N_1551,N_1463,N_1489);
nand U1552 (N_1552,N_1467,N_1407);
and U1553 (N_1553,N_1430,N_1403);
nand U1554 (N_1554,N_1432,N_1436);
or U1555 (N_1555,N_1461,N_1487);
nand U1556 (N_1556,N_1467,N_1494);
nor U1557 (N_1557,N_1483,N_1422);
nor U1558 (N_1558,N_1499,N_1414);
nand U1559 (N_1559,N_1404,N_1496);
nand U1560 (N_1560,N_1486,N_1414);
nor U1561 (N_1561,N_1483,N_1421);
nand U1562 (N_1562,N_1407,N_1468);
nand U1563 (N_1563,N_1453,N_1422);
nand U1564 (N_1564,N_1454,N_1476);
and U1565 (N_1565,N_1491,N_1485);
nand U1566 (N_1566,N_1456,N_1455);
or U1567 (N_1567,N_1499,N_1470);
or U1568 (N_1568,N_1488,N_1430);
or U1569 (N_1569,N_1495,N_1409);
and U1570 (N_1570,N_1470,N_1477);
nand U1571 (N_1571,N_1403,N_1468);
nor U1572 (N_1572,N_1432,N_1456);
and U1573 (N_1573,N_1471,N_1407);
or U1574 (N_1574,N_1472,N_1432);
or U1575 (N_1575,N_1424,N_1417);
nor U1576 (N_1576,N_1439,N_1475);
or U1577 (N_1577,N_1439,N_1446);
nand U1578 (N_1578,N_1466,N_1407);
or U1579 (N_1579,N_1420,N_1417);
nand U1580 (N_1580,N_1476,N_1495);
nor U1581 (N_1581,N_1422,N_1427);
nand U1582 (N_1582,N_1470,N_1443);
nand U1583 (N_1583,N_1460,N_1494);
or U1584 (N_1584,N_1415,N_1466);
or U1585 (N_1585,N_1464,N_1423);
or U1586 (N_1586,N_1446,N_1480);
nand U1587 (N_1587,N_1443,N_1453);
or U1588 (N_1588,N_1459,N_1410);
or U1589 (N_1589,N_1481,N_1479);
nor U1590 (N_1590,N_1450,N_1467);
or U1591 (N_1591,N_1456,N_1496);
nand U1592 (N_1592,N_1429,N_1454);
or U1593 (N_1593,N_1413,N_1466);
or U1594 (N_1594,N_1477,N_1448);
xor U1595 (N_1595,N_1443,N_1414);
nor U1596 (N_1596,N_1413,N_1421);
nand U1597 (N_1597,N_1407,N_1425);
or U1598 (N_1598,N_1459,N_1426);
or U1599 (N_1599,N_1447,N_1463);
or U1600 (N_1600,N_1541,N_1530);
nor U1601 (N_1601,N_1503,N_1584);
nand U1602 (N_1602,N_1583,N_1517);
and U1603 (N_1603,N_1590,N_1593);
or U1604 (N_1604,N_1597,N_1527);
nand U1605 (N_1605,N_1522,N_1552);
and U1606 (N_1606,N_1510,N_1540);
nand U1607 (N_1607,N_1576,N_1551);
nand U1608 (N_1608,N_1521,N_1505);
nor U1609 (N_1609,N_1561,N_1514);
nand U1610 (N_1610,N_1586,N_1566);
nor U1611 (N_1611,N_1578,N_1538);
or U1612 (N_1612,N_1526,N_1594);
or U1613 (N_1613,N_1547,N_1544);
nand U1614 (N_1614,N_1553,N_1592);
nor U1615 (N_1615,N_1548,N_1542);
or U1616 (N_1616,N_1562,N_1588);
or U1617 (N_1617,N_1589,N_1533);
nand U1618 (N_1618,N_1509,N_1571);
nor U1619 (N_1619,N_1504,N_1502);
nor U1620 (N_1620,N_1535,N_1567);
or U1621 (N_1621,N_1557,N_1536);
nor U1622 (N_1622,N_1574,N_1528);
or U1623 (N_1623,N_1556,N_1596);
and U1624 (N_1624,N_1559,N_1520);
or U1625 (N_1625,N_1579,N_1555);
nand U1626 (N_1626,N_1532,N_1585);
nand U1627 (N_1627,N_1572,N_1543);
or U1628 (N_1628,N_1519,N_1513);
nor U1629 (N_1629,N_1569,N_1549);
or U1630 (N_1630,N_1587,N_1577);
nand U1631 (N_1631,N_1564,N_1515);
or U1632 (N_1632,N_1550,N_1531);
nor U1633 (N_1633,N_1570,N_1563);
or U1634 (N_1634,N_1534,N_1529);
or U1635 (N_1635,N_1523,N_1518);
nand U1636 (N_1636,N_1537,N_1580);
or U1637 (N_1637,N_1595,N_1591);
nor U1638 (N_1638,N_1545,N_1501);
and U1639 (N_1639,N_1582,N_1560);
or U1640 (N_1640,N_1512,N_1516);
nor U1641 (N_1641,N_1558,N_1581);
or U1642 (N_1642,N_1524,N_1599);
and U1643 (N_1643,N_1500,N_1507);
nor U1644 (N_1644,N_1565,N_1539);
or U1645 (N_1645,N_1546,N_1573);
and U1646 (N_1646,N_1525,N_1554);
xnor U1647 (N_1647,N_1508,N_1506);
xnor U1648 (N_1648,N_1568,N_1511);
nor U1649 (N_1649,N_1598,N_1575);
and U1650 (N_1650,N_1575,N_1518);
or U1651 (N_1651,N_1537,N_1515);
or U1652 (N_1652,N_1574,N_1522);
nor U1653 (N_1653,N_1550,N_1561);
xor U1654 (N_1654,N_1588,N_1572);
and U1655 (N_1655,N_1558,N_1587);
or U1656 (N_1656,N_1571,N_1510);
and U1657 (N_1657,N_1588,N_1509);
and U1658 (N_1658,N_1592,N_1504);
and U1659 (N_1659,N_1502,N_1584);
xnor U1660 (N_1660,N_1532,N_1525);
nand U1661 (N_1661,N_1503,N_1598);
and U1662 (N_1662,N_1545,N_1593);
or U1663 (N_1663,N_1537,N_1543);
nor U1664 (N_1664,N_1509,N_1521);
and U1665 (N_1665,N_1500,N_1593);
and U1666 (N_1666,N_1514,N_1544);
nor U1667 (N_1667,N_1512,N_1557);
or U1668 (N_1668,N_1512,N_1513);
and U1669 (N_1669,N_1518,N_1553);
nor U1670 (N_1670,N_1596,N_1579);
and U1671 (N_1671,N_1522,N_1581);
or U1672 (N_1672,N_1506,N_1538);
nand U1673 (N_1673,N_1564,N_1514);
and U1674 (N_1674,N_1509,N_1564);
or U1675 (N_1675,N_1536,N_1556);
or U1676 (N_1676,N_1589,N_1501);
or U1677 (N_1677,N_1536,N_1563);
nand U1678 (N_1678,N_1514,N_1507);
or U1679 (N_1679,N_1530,N_1500);
xor U1680 (N_1680,N_1538,N_1541);
nor U1681 (N_1681,N_1579,N_1591);
or U1682 (N_1682,N_1500,N_1579);
nand U1683 (N_1683,N_1587,N_1580);
or U1684 (N_1684,N_1550,N_1513);
and U1685 (N_1685,N_1522,N_1507);
nand U1686 (N_1686,N_1511,N_1569);
nor U1687 (N_1687,N_1505,N_1557);
or U1688 (N_1688,N_1513,N_1500);
nand U1689 (N_1689,N_1577,N_1571);
and U1690 (N_1690,N_1504,N_1507);
or U1691 (N_1691,N_1551,N_1514);
and U1692 (N_1692,N_1547,N_1540);
nand U1693 (N_1693,N_1502,N_1543);
and U1694 (N_1694,N_1505,N_1540);
or U1695 (N_1695,N_1584,N_1526);
nor U1696 (N_1696,N_1578,N_1556);
nand U1697 (N_1697,N_1573,N_1519);
nor U1698 (N_1698,N_1540,N_1560);
and U1699 (N_1699,N_1556,N_1575);
nor U1700 (N_1700,N_1638,N_1651);
or U1701 (N_1701,N_1697,N_1663);
xnor U1702 (N_1702,N_1614,N_1681);
and U1703 (N_1703,N_1600,N_1680);
nor U1704 (N_1704,N_1628,N_1645);
and U1705 (N_1705,N_1679,N_1676);
nor U1706 (N_1706,N_1612,N_1684);
nor U1707 (N_1707,N_1683,N_1664);
xnor U1708 (N_1708,N_1662,N_1627);
nor U1709 (N_1709,N_1678,N_1691);
or U1710 (N_1710,N_1670,N_1690);
and U1711 (N_1711,N_1687,N_1647);
or U1712 (N_1712,N_1633,N_1617);
nor U1713 (N_1713,N_1696,N_1686);
and U1714 (N_1714,N_1650,N_1671);
or U1715 (N_1715,N_1619,N_1674);
nand U1716 (N_1716,N_1640,N_1605);
or U1717 (N_1717,N_1603,N_1656);
nand U1718 (N_1718,N_1622,N_1698);
and U1719 (N_1719,N_1616,N_1639);
nor U1720 (N_1720,N_1611,N_1637);
and U1721 (N_1721,N_1675,N_1644);
and U1722 (N_1722,N_1694,N_1667);
and U1723 (N_1723,N_1655,N_1669);
nor U1724 (N_1724,N_1653,N_1643);
nor U1725 (N_1725,N_1642,N_1661);
or U1726 (N_1726,N_1615,N_1607);
nor U1727 (N_1727,N_1609,N_1648);
or U1728 (N_1728,N_1641,N_1626);
and U1729 (N_1729,N_1672,N_1652);
and U1730 (N_1730,N_1695,N_1625);
nor U1731 (N_1731,N_1613,N_1693);
nand U1732 (N_1732,N_1606,N_1677);
nand U1733 (N_1733,N_1632,N_1620);
nor U1734 (N_1734,N_1602,N_1646);
nor U1735 (N_1735,N_1631,N_1699);
nor U1736 (N_1736,N_1657,N_1659);
nand U1737 (N_1737,N_1601,N_1665);
nand U1738 (N_1738,N_1660,N_1629);
and U1739 (N_1739,N_1608,N_1634);
nand U1740 (N_1740,N_1630,N_1635);
and U1741 (N_1741,N_1623,N_1610);
nand U1742 (N_1742,N_1604,N_1689);
or U1743 (N_1743,N_1654,N_1673);
nor U1744 (N_1744,N_1688,N_1618);
nor U1745 (N_1745,N_1649,N_1658);
nand U1746 (N_1746,N_1624,N_1636);
or U1747 (N_1747,N_1621,N_1666);
nand U1748 (N_1748,N_1692,N_1668);
nand U1749 (N_1749,N_1685,N_1682);
nor U1750 (N_1750,N_1699,N_1672);
and U1751 (N_1751,N_1637,N_1647);
and U1752 (N_1752,N_1604,N_1629);
nand U1753 (N_1753,N_1631,N_1635);
nor U1754 (N_1754,N_1610,N_1679);
and U1755 (N_1755,N_1630,N_1658);
nor U1756 (N_1756,N_1619,N_1673);
nor U1757 (N_1757,N_1633,N_1641);
or U1758 (N_1758,N_1650,N_1651);
and U1759 (N_1759,N_1653,N_1646);
or U1760 (N_1760,N_1666,N_1642);
or U1761 (N_1761,N_1675,N_1672);
nand U1762 (N_1762,N_1660,N_1655);
or U1763 (N_1763,N_1638,N_1611);
nand U1764 (N_1764,N_1620,N_1693);
nand U1765 (N_1765,N_1676,N_1687);
nand U1766 (N_1766,N_1681,N_1655);
and U1767 (N_1767,N_1630,N_1626);
or U1768 (N_1768,N_1630,N_1603);
and U1769 (N_1769,N_1640,N_1691);
nor U1770 (N_1770,N_1658,N_1629);
and U1771 (N_1771,N_1650,N_1664);
and U1772 (N_1772,N_1645,N_1642);
or U1773 (N_1773,N_1655,N_1622);
nor U1774 (N_1774,N_1639,N_1659);
nor U1775 (N_1775,N_1639,N_1655);
and U1776 (N_1776,N_1683,N_1679);
nand U1777 (N_1777,N_1669,N_1690);
nor U1778 (N_1778,N_1642,N_1698);
or U1779 (N_1779,N_1603,N_1620);
and U1780 (N_1780,N_1611,N_1621);
nand U1781 (N_1781,N_1620,N_1610);
nor U1782 (N_1782,N_1635,N_1625);
nor U1783 (N_1783,N_1642,N_1670);
and U1784 (N_1784,N_1690,N_1662);
or U1785 (N_1785,N_1693,N_1636);
nand U1786 (N_1786,N_1695,N_1649);
and U1787 (N_1787,N_1607,N_1668);
xor U1788 (N_1788,N_1655,N_1645);
and U1789 (N_1789,N_1623,N_1650);
or U1790 (N_1790,N_1667,N_1645);
and U1791 (N_1791,N_1637,N_1655);
nor U1792 (N_1792,N_1616,N_1651);
nor U1793 (N_1793,N_1636,N_1685);
and U1794 (N_1794,N_1618,N_1608);
or U1795 (N_1795,N_1661,N_1689);
nand U1796 (N_1796,N_1683,N_1637);
nand U1797 (N_1797,N_1609,N_1623);
or U1798 (N_1798,N_1646,N_1607);
nand U1799 (N_1799,N_1626,N_1675);
or U1800 (N_1800,N_1786,N_1788);
or U1801 (N_1801,N_1771,N_1753);
and U1802 (N_1802,N_1750,N_1798);
nand U1803 (N_1803,N_1792,N_1730);
and U1804 (N_1804,N_1704,N_1711);
nor U1805 (N_1805,N_1791,N_1759);
nand U1806 (N_1806,N_1713,N_1790);
and U1807 (N_1807,N_1762,N_1712);
or U1808 (N_1808,N_1744,N_1718);
and U1809 (N_1809,N_1701,N_1787);
and U1810 (N_1810,N_1706,N_1741);
nand U1811 (N_1811,N_1761,N_1794);
or U1812 (N_1812,N_1746,N_1723);
nand U1813 (N_1813,N_1767,N_1766);
and U1814 (N_1814,N_1782,N_1708);
nand U1815 (N_1815,N_1780,N_1755);
nor U1816 (N_1816,N_1726,N_1764);
nand U1817 (N_1817,N_1740,N_1789);
nand U1818 (N_1818,N_1720,N_1745);
and U1819 (N_1819,N_1770,N_1700);
or U1820 (N_1820,N_1751,N_1727);
or U1821 (N_1821,N_1775,N_1776);
and U1822 (N_1822,N_1724,N_1736);
nor U1823 (N_1823,N_1747,N_1722);
or U1824 (N_1824,N_1783,N_1779);
nor U1825 (N_1825,N_1749,N_1763);
nor U1826 (N_1826,N_1717,N_1777);
nand U1827 (N_1827,N_1796,N_1793);
nand U1828 (N_1828,N_1799,N_1731);
or U1829 (N_1829,N_1739,N_1773);
nor U1830 (N_1830,N_1702,N_1754);
or U1831 (N_1831,N_1728,N_1715);
and U1832 (N_1832,N_1714,N_1719);
nand U1833 (N_1833,N_1705,N_1752);
nand U1834 (N_1834,N_1743,N_1769);
or U1835 (N_1835,N_1760,N_1758);
and U1836 (N_1836,N_1772,N_1756);
or U1837 (N_1837,N_1765,N_1768);
nand U1838 (N_1838,N_1709,N_1703);
and U1839 (N_1839,N_1784,N_1732);
or U1840 (N_1840,N_1737,N_1757);
nand U1841 (N_1841,N_1742,N_1729);
nor U1842 (N_1842,N_1721,N_1778);
nand U1843 (N_1843,N_1733,N_1738);
and U1844 (N_1844,N_1725,N_1797);
nand U1845 (N_1845,N_1735,N_1710);
or U1846 (N_1846,N_1707,N_1795);
and U1847 (N_1847,N_1748,N_1781);
nor U1848 (N_1848,N_1734,N_1785);
or U1849 (N_1849,N_1716,N_1774);
and U1850 (N_1850,N_1721,N_1763);
or U1851 (N_1851,N_1711,N_1777);
or U1852 (N_1852,N_1733,N_1796);
or U1853 (N_1853,N_1704,N_1795);
or U1854 (N_1854,N_1779,N_1715);
and U1855 (N_1855,N_1784,N_1792);
nor U1856 (N_1856,N_1745,N_1791);
nor U1857 (N_1857,N_1749,N_1743);
nor U1858 (N_1858,N_1767,N_1716);
nor U1859 (N_1859,N_1799,N_1752);
nand U1860 (N_1860,N_1700,N_1726);
or U1861 (N_1861,N_1798,N_1762);
nand U1862 (N_1862,N_1724,N_1765);
nor U1863 (N_1863,N_1789,N_1777);
nand U1864 (N_1864,N_1704,N_1777);
nand U1865 (N_1865,N_1726,N_1757);
nor U1866 (N_1866,N_1739,N_1715);
or U1867 (N_1867,N_1707,N_1755);
or U1868 (N_1868,N_1768,N_1759);
and U1869 (N_1869,N_1723,N_1772);
nand U1870 (N_1870,N_1718,N_1793);
nor U1871 (N_1871,N_1791,N_1744);
and U1872 (N_1872,N_1782,N_1757);
nor U1873 (N_1873,N_1796,N_1795);
nand U1874 (N_1874,N_1740,N_1735);
nor U1875 (N_1875,N_1758,N_1764);
or U1876 (N_1876,N_1764,N_1736);
or U1877 (N_1877,N_1789,N_1731);
and U1878 (N_1878,N_1757,N_1791);
or U1879 (N_1879,N_1725,N_1763);
and U1880 (N_1880,N_1721,N_1720);
nand U1881 (N_1881,N_1727,N_1787);
nand U1882 (N_1882,N_1740,N_1705);
and U1883 (N_1883,N_1716,N_1765);
nand U1884 (N_1884,N_1750,N_1733);
xnor U1885 (N_1885,N_1711,N_1721);
or U1886 (N_1886,N_1745,N_1710);
nand U1887 (N_1887,N_1743,N_1766);
or U1888 (N_1888,N_1720,N_1718);
or U1889 (N_1889,N_1779,N_1755);
nand U1890 (N_1890,N_1768,N_1774);
nor U1891 (N_1891,N_1711,N_1738);
nor U1892 (N_1892,N_1777,N_1743);
nand U1893 (N_1893,N_1730,N_1799);
or U1894 (N_1894,N_1752,N_1716);
nand U1895 (N_1895,N_1790,N_1754);
nand U1896 (N_1896,N_1730,N_1760);
nand U1897 (N_1897,N_1724,N_1713);
and U1898 (N_1898,N_1771,N_1716);
or U1899 (N_1899,N_1798,N_1776);
nor U1900 (N_1900,N_1878,N_1883);
and U1901 (N_1901,N_1825,N_1801);
nand U1902 (N_1902,N_1882,N_1800);
and U1903 (N_1903,N_1829,N_1876);
nand U1904 (N_1904,N_1897,N_1852);
and U1905 (N_1905,N_1816,N_1884);
nor U1906 (N_1906,N_1822,N_1824);
nand U1907 (N_1907,N_1867,N_1812);
or U1908 (N_1908,N_1870,N_1838);
or U1909 (N_1909,N_1844,N_1891);
nor U1910 (N_1910,N_1862,N_1809);
nand U1911 (N_1911,N_1858,N_1803);
nor U1912 (N_1912,N_1811,N_1814);
nor U1913 (N_1913,N_1842,N_1863);
nand U1914 (N_1914,N_1874,N_1806);
or U1915 (N_1915,N_1872,N_1894);
and U1916 (N_1916,N_1854,N_1828);
and U1917 (N_1917,N_1850,N_1837);
or U1918 (N_1918,N_1818,N_1804);
nand U1919 (N_1919,N_1830,N_1857);
nor U1920 (N_1920,N_1865,N_1864);
xnor U1921 (N_1921,N_1895,N_1855);
or U1922 (N_1922,N_1845,N_1898);
nand U1923 (N_1923,N_1885,N_1846);
or U1924 (N_1924,N_1817,N_1831);
or U1925 (N_1925,N_1851,N_1869);
nand U1926 (N_1926,N_1813,N_1890);
nand U1927 (N_1927,N_1880,N_1821);
nand U1928 (N_1928,N_1834,N_1886);
or U1929 (N_1929,N_1839,N_1808);
and U1930 (N_1930,N_1881,N_1848);
or U1931 (N_1931,N_1823,N_1879);
nor U1932 (N_1932,N_1827,N_1859);
nor U1933 (N_1933,N_1819,N_1815);
or U1934 (N_1934,N_1853,N_1840);
xor U1935 (N_1935,N_1866,N_1802);
or U1936 (N_1936,N_1875,N_1860);
nand U1937 (N_1937,N_1868,N_1826);
nor U1938 (N_1938,N_1871,N_1899);
or U1939 (N_1939,N_1861,N_1841);
nor U1940 (N_1940,N_1896,N_1820);
and U1941 (N_1941,N_1893,N_1873);
nand U1942 (N_1942,N_1877,N_1833);
or U1943 (N_1943,N_1836,N_1805);
nand U1944 (N_1944,N_1856,N_1847);
nor U1945 (N_1945,N_1843,N_1889);
nor U1946 (N_1946,N_1849,N_1888);
and U1947 (N_1947,N_1832,N_1807);
xnor U1948 (N_1948,N_1887,N_1810);
and U1949 (N_1949,N_1835,N_1892);
and U1950 (N_1950,N_1810,N_1809);
nor U1951 (N_1951,N_1806,N_1861);
nor U1952 (N_1952,N_1871,N_1811);
nand U1953 (N_1953,N_1810,N_1868);
nand U1954 (N_1954,N_1875,N_1894);
or U1955 (N_1955,N_1810,N_1804);
nor U1956 (N_1956,N_1838,N_1850);
or U1957 (N_1957,N_1863,N_1892);
and U1958 (N_1958,N_1810,N_1853);
nor U1959 (N_1959,N_1872,N_1810);
nand U1960 (N_1960,N_1811,N_1889);
xor U1961 (N_1961,N_1810,N_1819);
nor U1962 (N_1962,N_1815,N_1842);
and U1963 (N_1963,N_1883,N_1861);
nand U1964 (N_1964,N_1845,N_1828);
nor U1965 (N_1965,N_1850,N_1874);
nand U1966 (N_1966,N_1852,N_1836);
or U1967 (N_1967,N_1895,N_1874);
nor U1968 (N_1968,N_1893,N_1839);
nand U1969 (N_1969,N_1866,N_1818);
nand U1970 (N_1970,N_1840,N_1888);
and U1971 (N_1971,N_1852,N_1867);
nand U1972 (N_1972,N_1819,N_1889);
nand U1973 (N_1973,N_1815,N_1856);
or U1974 (N_1974,N_1820,N_1819);
and U1975 (N_1975,N_1853,N_1805);
and U1976 (N_1976,N_1844,N_1816);
nand U1977 (N_1977,N_1896,N_1842);
nand U1978 (N_1978,N_1800,N_1883);
nor U1979 (N_1979,N_1804,N_1829);
and U1980 (N_1980,N_1843,N_1825);
nor U1981 (N_1981,N_1824,N_1848);
or U1982 (N_1982,N_1803,N_1849);
or U1983 (N_1983,N_1840,N_1808);
and U1984 (N_1984,N_1880,N_1842);
and U1985 (N_1985,N_1812,N_1878);
or U1986 (N_1986,N_1881,N_1849);
and U1987 (N_1987,N_1899,N_1861);
and U1988 (N_1988,N_1827,N_1826);
or U1989 (N_1989,N_1877,N_1814);
nor U1990 (N_1990,N_1850,N_1813);
nand U1991 (N_1991,N_1824,N_1857);
nor U1992 (N_1992,N_1865,N_1852);
and U1993 (N_1993,N_1836,N_1840);
nor U1994 (N_1994,N_1808,N_1849);
xnor U1995 (N_1995,N_1829,N_1849);
nor U1996 (N_1996,N_1889,N_1872);
or U1997 (N_1997,N_1838,N_1804);
and U1998 (N_1998,N_1847,N_1858);
and U1999 (N_1999,N_1808,N_1817);
nand U2000 (N_2000,N_1951,N_1960);
or U2001 (N_2001,N_1906,N_1907);
nand U2002 (N_2002,N_1950,N_1957);
and U2003 (N_2003,N_1970,N_1979);
and U2004 (N_2004,N_1943,N_1937);
nor U2005 (N_2005,N_1972,N_1940);
and U2006 (N_2006,N_1963,N_1985);
nand U2007 (N_2007,N_1915,N_1909);
or U2008 (N_2008,N_1930,N_1922);
nor U2009 (N_2009,N_1928,N_1965);
nor U2010 (N_2010,N_1923,N_1980);
or U2011 (N_2011,N_1953,N_1990);
or U2012 (N_2012,N_1992,N_1955);
or U2013 (N_2013,N_1925,N_1976);
or U2014 (N_2014,N_1968,N_1958);
nor U2015 (N_2015,N_1993,N_1926);
or U2016 (N_2016,N_1971,N_1933);
nand U2017 (N_2017,N_1978,N_1936);
nand U2018 (N_2018,N_1910,N_1938);
and U2019 (N_2019,N_1920,N_1918);
nor U2020 (N_2020,N_1945,N_1994);
nand U2021 (N_2021,N_1961,N_1959);
nor U2022 (N_2022,N_1946,N_1973);
and U2023 (N_2023,N_1902,N_1916);
and U2024 (N_2024,N_1989,N_1988);
or U2025 (N_2025,N_1941,N_1975);
nand U2026 (N_2026,N_1952,N_1991);
or U2027 (N_2027,N_1939,N_1969);
nand U2028 (N_2028,N_1964,N_1948);
or U2029 (N_2029,N_1904,N_1944);
nor U2030 (N_2030,N_1934,N_1967);
or U2031 (N_2031,N_1900,N_1942);
nor U2032 (N_2032,N_1929,N_1903);
and U2033 (N_2033,N_1914,N_1901);
nand U2034 (N_2034,N_1935,N_1995);
nand U2035 (N_2035,N_1996,N_1912);
nor U2036 (N_2036,N_1947,N_1962);
or U2037 (N_2037,N_1987,N_1927);
or U2038 (N_2038,N_1954,N_1924);
nand U2039 (N_2039,N_1983,N_1977);
nor U2040 (N_2040,N_1966,N_1986);
and U2041 (N_2041,N_1999,N_1932);
nand U2042 (N_2042,N_1931,N_1905);
nor U2043 (N_2043,N_1913,N_1997);
and U2044 (N_2044,N_1921,N_1917);
nor U2045 (N_2045,N_1984,N_1908);
or U2046 (N_2046,N_1974,N_1919);
or U2047 (N_2047,N_1911,N_1956);
nor U2048 (N_2048,N_1981,N_1982);
and U2049 (N_2049,N_1949,N_1998);
nor U2050 (N_2050,N_1989,N_1966);
nor U2051 (N_2051,N_1997,N_1984);
nand U2052 (N_2052,N_1936,N_1900);
nand U2053 (N_2053,N_1950,N_1995);
and U2054 (N_2054,N_1925,N_1933);
or U2055 (N_2055,N_1990,N_1905);
or U2056 (N_2056,N_1923,N_1913);
nor U2057 (N_2057,N_1966,N_1925);
nand U2058 (N_2058,N_1975,N_1968);
or U2059 (N_2059,N_1901,N_1906);
and U2060 (N_2060,N_1914,N_1928);
nand U2061 (N_2061,N_1909,N_1939);
and U2062 (N_2062,N_1922,N_1906);
nand U2063 (N_2063,N_1988,N_1906);
xor U2064 (N_2064,N_1925,N_1916);
or U2065 (N_2065,N_1944,N_1963);
nand U2066 (N_2066,N_1965,N_1910);
nor U2067 (N_2067,N_1976,N_1900);
nor U2068 (N_2068,N_1919,N_1995);
or U2069 (N_2069,N_1911,N_1958);
nor U2070 (N_2070,N_1982,N_1997);
nand U2071 (N_2071,N_1973,N_1970);
nor U2072 (N_2072,N_1930,N_1933);
nor U2073 (N_2073,N_1992,N_1905);
and U2074 (N_2074,N_1988,N_1997);
or U2075 (N_2075,N_1974,N_1980);
nor U2076 (N_2076,N_1974,N_1983);
nor U2077 (N_2077,N_1945,N_1944);
nand U2078 (N_2078,N_1929,N_1933);
nand U2079 (N_2079,N_1990,N_1901);
or U2080 (N_2080,N_1970,N_1942);
nand U2081 (N_2081,N_1997,N_1953);
and U2082 (N_2082,N_1961,N_1941);
nand U2083 (N_2083,N_1995,N_1906);
and U2084 (N_2084,N_1922,N_1958);
and U2085 (N_2085,N_1920,N_1950);
nand U2086 (N_2086,N_1914,N_1911);
nor U2087 (N_2087,N_1930,N_1907);
or U2088 (N_2088,N_1949,N_1986);
nand U2089 (N_2089,N_1990,N_1910);
xor U2090 (N_2090,N_1982,N_1998);
and U2091 (N_2091,N_1952,N_1962);
or U2092 (N_2092,N_1962,N_1925);
and U2093 (N_2093,N_1963,N_1943);
nor U2094 (N_2094,N_1940,N_1929);
nor U2095 (N_2095,N_1945,N_1987);
or U2096 (N_2096,N_1950,N_1969);
nand U2097 (N_2097,N_1990,N_1909);
nor U2098 (N_2098,N_1940,N_1998);
nor U2099 (N_2099,N_1981,N_1915);
nand U2100 (N_2100,N_2090,N_2050);
nor U2101 (N_2101,N_2023,N_2034);
nor U2102 (N_2102,N_2084,N_2081);
nor U2103 (N_2103,N_2055,N_2086);
nor U2104 (N_2104,N_2027,N_2096);
nand U2105 (N_2105,N_2028,N_2058);
and U2106 (N_2106,N_2012,N_2040);
or U2107 (N_2107,N_2005,N_2016);
or U2108 (N_2108,N_2066,N_2026);
and U2109 (N_2109,N_2010,N_2018);
and U2110 (N_2110,N_2036,N_2059);
nor U2111 (N_2111,N_2099,N_2035);
nand U2112 (N_2112,N_2075,N_2015);
and U2113 (N_2113,N_2051,N_2047);
or U2114 (N_2114,N_2093,N_2007);
or U2115 (N_2115,N_2082,N_2098);
or U2116 (N_2116,N_2030,N_2078);
or U2117 (N_2117,N_2006,N_2073);
nor U2118 (N_2118,N_2003,N_2032);
nor U2119 (N_2119,N_2038,N_2048);
and U2120 (N_2120,N_2046,N_2063);
or U2121 (N_2121,N_2087,N_2002);
or U2122 (N_2122,N_2029,N_2061);
and U2123 (N_2123,N_2019,N_2094);
nand U2124 (N_2124,N_2085,N_2014);
nand U2125 (N_2125,N_2049,N_2072);
nor U2126 (N_2126,N_2000,N_2079);
and U2127 (N_2127,N_2062,N_2069);
nor U2128 (N_2128,N_2031,N_2053);
and U2129 (N_2129,N_2043,N_2025);
or U2130 (N_2130,N_2020,N_2071);
and U2131 (N_2131,N_2057,N_2088);
and U2132 (N_2132,N_2091,N_2065);
and U2133 (N_2133,N_2037,N_2008);
xor U2134 (N_2134,N_2022,N_2076);
nor U2135 (N_2135,N_2044,N_2033);
and U2136 (N_2136,N_2054,N_2064);
nor U2137 (N_2137,N_2097,N_2067);
or U2138 (N_2138,N_2089,N_2017);
and U2139 (N_2139,N_2070,N_2092);
and U2140 (N_2140,N_2001,N_2080);
nand U2141 (N_2141,N_2009,N_2042);
nor U2142 (N_2142,N_2013,N_2039);
nand U2143 (N_2143,N_2021,N_2004);
nand U2144 (N_2144,N_2052,N_2068);
nand U2145 (N_2145,N_2095,N_2045);
and U2146 (N_2146,N_2024,N_2041);
and U2147 (N_2147,N_2083,N_2011);
nand U2148 (N_2148,N_2056,N_2060);
nand U2149 (N_2149,N_2074,N_2077);
nor U2150 (N_2150,N_2015,N_2083);
nand U2151 (N_2151,N_2001,N_2079);
nand U2152 (N_2152,N_2062,N_2040);
nor U2153 (N_2153,N_2087,N_2018);
nand U2154 (N_2154,N_2074,N_2002);
or U2155 (N_2155,N_2037,N_2018);
nand U2156 (N_2156,N_2090,N_2005);
nor U2157 (N_2157,N_2098,N_2008);
or U2158 (N_2158,N_2085,N_2000);
or U2159 (N_2159,N_2084,N_2046);
or U2160 (N_2160,N_2024,N_2080);
nand U2161 (N_2161,N_2008,N_2022);
and U2162 (N_2162,N_2095,N_2000);
or U2163 (N_2163,N_2045,N_2077);
and U2164 (N_2164,N_2074,N_2022);
or U2165 (N_2165,N_2041,N_2076);
nand U2166 (N_2166,N_2008,N_2039);
and U2167 (N_2167,N_2083,N_2010);
nand U2168 (N_2168,N_2061,N_2026);
nor U2169 (N_2169,N_2061,N_2073);
or U2170 (N_2170,N_2032,N_2063);
and U2171 (N_2171,N_2000,N_2015);
or U2172 (N_2172,N_2003,N_2057);
xnor U2173 (N_2173,N_2008,N_2083);
nand U2174 (N_2174,N_2091,N_2023);
nor U2175 (N_2175,N_2037,N_2055);
nand U2176 (N_2176,N_2077,N_2019);
nor U2177 (N_2177,N_2089,N_2025);
or U2178 (N_2178,N_2087,N_2072);
and U2179 (N_2179,N_2062,N_2098);
nand U2180 (N_2180,N_2044,N_2049);
and U2181 (N_2181,N_2037,N_2026);
nand U2182 (N_2182,N_2059,N_2016);
and U2183 (N_2183,N_2031,N_2043);
or U2184 (N_2184,N_2034,N_2047);
and U2185 (N_2185,N_2095,N_2053);
nand U2186 (N_2186,N_2051,N_2092);
xor U2187 (N_2187,N_2099,N_2074);
and U2188 (N_2188,N_2083,N_2037);
xor U2189 (N_2189,N_2027,N_2059);
nand U2190 (N_2190,N_2005,N_2099);
and U2191 (N_2191,N_2094,N_2010);
nor U2192 (N_2192,N_2095,N_2071);
xor U2193 (N_2193,N_2009,N_2036);
nand U2194 (N_2194,N_2098,N_2051);
nand U2195 (N_2195,N_2088,N_2064);
nand U2196 (N_2196,N_2009,N_2012);
nand U2197 (N_2197,N_2001,N_2091);
xor U2198 (N_2198,N_2022,N_2086);
nand U2199 (N_2199,N_2039,N_2048);
and U2200 (N_2200,N_2196,N_2136);
nor U2201 (N_2201,N_2113,N_2182);
nor U2202 (N_2202,N_2118,N_2131);
nor U2203 (N_2203,N_2175,N_2110);
nor U2204 (N_2204,N_2111,N_2160);
nor U2205 (N_2205,N_2163,N_2193);
and U2206 (N_2206,N_2103,N_2186);
nor U2207 (N_2207,N_2106,N_2185);
or U2208 (N_2208,N_2161,N_2166);
nand U2209 (N_2209,N_2101,N_2127);
nor U2210 (N_2210,N_2192,N_2194);
nand U2211 (N_2211,N_2138,N_2139);
nand U2212 (N_2212,N_2158,N_2148);
or U2213 (N_2213,N_2123,N_2120);
and U2214 (N_2214,N_2143,N_2117);
and U2215 (N_2215,N_2112,N_2109);
and U2216 (N_2216,N_2119,N_2184);
nor U2217 (N_2217,N_2159,N_2199);
nand U2218 (N_2218,N_2122,N_2133);
and U2219 (N_2219,N_2132,N_2169);
and U2220 (N_2220,N_2188,N_2107);
or U2221 (N_2221,N_2147,N_2198);
or U2222 (N_2222,N_2181,N_2171);
nand U2223 (N_2223,N_2174,N_2170);
or U2224 (N_2224,N_2183,N_2145);
or U2225 (N_2225,N_2130,N_2167);
or U2226 (N_2226,N_2153,N_2154);
or U2227 (N_2227,N_2126,N_2105);
nor U2228 (N_2228,N_2157,N_2142);
nor U2229 (N_2229,N_2173,N_2197);
nor U2230 (N_2230,N_2108,N_2125);
nor U2231 (N_2231,N_2168,N_2189);
and U2232 (N_2232,N_2178,N_2137);
or U2233 (N_2233,N_2165,N_2129);
or U2234 (N_2234,N_2114,N_2187);
or U2235 (N_2235,N_2152,N_2164);
nand U2236 (N_2236,N_2179,N_2116);
and U2237 (N_2237,N_2134,N_2180);
or U2238 (N_2238,N_2151,N_2104);
xor U2239 (N_2239,N_2195,N_2149);
or U2240 (N_2240,N_2190,N_2124);
nand U2241 (N_2241,N_2102,N_2176);
or U2242 (N_2242,N_2100,N_2155);
nor U2243 (N_2243,N_2128,N_2140);
nand U2244 (N_2244,N_2162,N_2121);
nor U2245 (N_2245,N_2115,N_2156);
or U2246 (N_2246,N_2172,N_2191);
or U2247 (N_2247,N_2150,N_2135);
nor U2248 (N_2248,N_2146,N_2177);
nor U2249 (N_2249,N_2141,N_2144);
or U2250 (N_2250,N_2171,N_2102);
nand U2251 (N_2251,N_2189,N_2192);
nor U2252 (N_2252,N_2160,N_2197);
nor U2253 (N_2253,N_2157,N_2191);
nor U2254 (N_2254,N_2124,N_2106);
or U2255 (N_2255,N_2152,N_2173);
or U2256 (N_2256,N_2194,N_2133);
and U2257 (N_2257,N_2159,N_2117);
or U2258 (N_2258,N_2152,N_2125);
nor U2259 (N_2259,N_2166,N_2108);
and U2260 (N_2260,N_2138,N_2129);
xor U2261 (N_2261,N_2191,N_2187);
and U2262 (N_2262,N_2174,N_2155);
and U2263 (N_2263,N_2197,N_2195);
nor U2264 (N_2264,N_2166,N_2175);
xor U2265 (N_2265,N_2166,N_2126);
nand U2266 (N_2266,N_2165,N_2124);
or U2267 (N_2267,N_2119,N_2146);
and U2268 (N_2268,N_2161,N_2164);
nor U2269 (N_2269,N_2155,N_2140);
nor U2270 (N_2270,N_2168,N_2143);
and U2271 (N_2271,N_2158,N_2141);
and U2272 (N_2272,N_2132,N_2198);
nand U2273 (N_2273,N_2192,N_2107);
xnor U2274 (N_2274,N_2183,N_2160);
nor U2275 (N_2275,N_2167,N_2151);
and U2276 (N_2276,N_2165,N_2121);
or U2277 (N_2277,N_2127,N_2157);
or U2278 (N_2278,N_2191,N_2131);
nand U2279 (N_2279,N_2126,N_2154);
nor U2280 (N_2280,N_2175,N_2179);
or U2281 (N_2281,N_2111,N_2179);
nand U2282 (N_2282,N_2149,N_2111);
nand U2283 (N_2283,N_2190,N_2151);
nor U2284 (N_2284,N_2108,N_2175);
nand U2285 (N_2285,N_2102,N_2186);
or U2286 (N_2286,N_2104,N_2192);
or U2287 (N_2287,N_2115,N_2151);
or U2288 (N_2288,N_2187,N_2182);
nand U2289 (N_2289,N_2162,N_2194);
nor U2290 (N_2290,N_2145,N_2190);
or U2291 (N_2291,N_2188,N_2128);
or U2292 (N_2292,N_2156,N_2193);
nand U2293 (N_2293,N_2171,N_2150);
nand U2294 (N_2294,N_2163,N_2104);
nor U2295 (N_2295,N_2193,N_2132);
nor U2296 (N_2296,N_2183,N_2123);
nand U2297 (N_2297,N_2129,N_2189);
nor U2298 (N_2298,N_2113,N_2129);
nand U2299 (N_2299,N_2152,N_2145);
nand U2300 (N_2300,N_2227,N_2211);
nand U2301 (N_2301,N_2216,N_2210);
or U2302 (N_2302,N_2239,N_2203);
or U2303 (N_2303,N_2281,N_2296);
and U2304 (N_2304,N_2254,N_2285);
and U2305 (N_2305,N_2206,N_2232);
or U2306 (N_2306,N_2267,N_2247);
and U2307 (N_2307,N_2255,N_2208);
nand U2308 (N_2308,N_2229,N_2260);
nand U2309 (N_2309,N_2237,N_2269);
xnor U2310 (N_2310,N_2231,N_2212);
or U2311 (N_2311,N_2228,N_2209);
or U2312 (N_2312,N_2282,N_2249);
and U2313 (N_2313,N_2276,N_2256);
or U2314 (N_2314,N_2295,N_2214);
and U2315 (N_2315,N_2258,N_2207);
nor U2316 (N_2316,N_2291,N_2221);
and U2317 (N_2317,N_2200,N_2243);
nand U2318 (N_2318,N_2244,N_2293);
nand U2319 (N_2319,N_2220,N_2248);
nor U2320 (N_2320,N_2297,N_2218);
and U2321 (N_2321,N_2292,N_2251);
nor U2322 (N_2322,N_2274,N_2266);
and U2323 (N_2323,N_2259,N_2271);
and U2324 (N_2324,N_2280,N_2235);
nor U2325 (N_2325,N_2287,N_2230);
nand U2326 (N_2326,N_2253,N_2277);
nand U2327 (N_2327,N_2261,N_2290);
nor U2328 (N_2328,N_2246,N_2275);
and U2329 (N_2329,N_2264,N_2205);
nor U2330 (N_2330,N_2283,N_2257);
or U2331 (N_2331,N_2202,N_2299);
nor U2332 (N_2332,N_2201,N_2224);
nor U2333 (N_2333,N_2272,N_2289);
nand U2334 (N_2334,N_2222,N_2252);
nand U2335 (N_2335,N_2263,N_2223);
nand U2336 (N_2336,N_2204,N_2286);
nor U2337 (N_2337,N_2233,N_2241);
nor U2338 (N_2338,N_2238,N_2219);
nand U2339 (N_2339,N_2245,N_2236);
nor U2340 (N_2340,N_2273,N_2234);
nand U2341 (N_2341,N_2215,N_2279);
nor U2342 (N_2342,N_2240,N_2262);
or U2343 (N_2343,N_2270,N_2284);
xnor U2344 (N_2344,N_2225,N_2278);
nor U2345 (N_2345,N_2226,N_2288);
nor U2346 (N_2346,N_2265,N_2294);
nand U2347 (N_2347,N_2250,N_2298);
or U2348 (N_2348,N_2268,N_2242);
nand U2349 (N_2349,N_2213,N_2217);
nand U2350 (N_2350,N_2236,N_2296);
nand U2351 (N_2351,N_2224,N_2222);
or U2352 (N_2352,N_2250,N_2293);
nand U2353 (N_2353,N_2275,N_2255);
nand U2354 (N_2354,N_2241,N_2248);
nand U2355 (N_2355,N_2279,N_2293);
nor U2356 (N_2356,N_2203,N_2281);
xnor U2357 (N_2357,N_2223,N_2280);
nor U2358 (N_2358,N_2260,N_2247);
nand U2359 (N_2359,N_2232,N_2201);
nand U2360 (N_2360,N_2289,N_2223);
nor U2361 (N_2361,N_2239,N_2259);
nand U2362 (N_2362,N_2262,N_2245);
nand U2363 (N_2363,N_2217,N_2211);
and U2364 (N_2364,N_2288,N_2224);
nand U2365 (N_2365,N_2272,N_2224);
nor U2366 (N_2366,N_2235,N_2283);
or U2367 (N_2367,N_2233,N_2216);
nor U2368 (N_2368,N_2219,N_2201);
or U2369 (N_2369,N_2297,N_2264);
and U2370 (N_2370,N_2265,N_2268);
xnor U2371 (N_2371,N_2277,N_2234);
or U2372 (N_2372,N_2200,N_2238);
nand U2373 (N_2373,N_2240,N_2288);
or U2374 (N_2374,N_2296,N_2222);
and U2375 (N_2375,N_2275,N_2200);
or U2376 (N_2376,N_2252,N_2263);
or U2377 (N_2377,N_2287,N_2245);
and U2378 (N_2378,N_2232,N_2222);
nor U2379 (N_2379,N_2224,N_2267);
and U2380 (N_2380,N_2244,N_2212);
or U2381 (N_2381,N_2210,N_2291);
or U2382 (N_2382,N_2233,N_2240);
nand U2383 (N_2383,N_2231,N_2223);
or U2384 (N_2384,N_2248,N_2214);
nor U2385 (N_2385,N_2258,N_2223);
nor U2386 (N_2386,N_2298,N_2221);
and U2387 (N_2387,N_2294,N_2256);
xor U2388 (N_2388,N_2206,N_2228);
and U2389 (N_2389,N_2253,N_2264);
nand U2390 (N_2390,N_2220,N_2283);
xor U2391 (N_2391,N_2266,N_2293);
or U2392 (N_2392,N_2298,N_2253);
or U2393 (N_2393,N_2201,N_2247);
nand U2394 (N_2394,N_2261,N_2276);
or U2395 (N_2395,N_2296,N_2218);
or U2396 (N_2396,N_2215,N_2211);
nand U2397 (N_2397,N_2223,N_2264);
nor U2398 (N_2398,N_2284,N_2213);
nand U2399 (N_2399,N_2224,N_2261);
nor U2400 (N_2400,N_2326,N_2363);
or U2401 (N_2401,N_2309,N_2386);
nor U2402 (N_2402,N_2350,N_2397);
or U2403 (N_2403,N_2346,N_2337);
nor U2404 (N_2404,N_2303,N_2329);
or U2405 (N_2405,N_2387,N_2321);
nor U2406 (N_2406,N_2314,N_2370);
or U2407 (N_2407,N_2368,N_2365);
and U2408 (N_2408,N_2349,N_2327);
nand U2409 (N_2409,N_2367,N_2347);
nand U2410 (N_2410,N_2374,N_2355);
nand U2411 (N_2411,N_2335,N_2330);
xor U2412 (N_2412,N_2394,N_2356);
nand U2413 (N_2413,N_2308,N_2392);
or U2414 (N_2414,N_2305,N_2302);
and U2415 (N_2415,N_2377,N_2336);
or U2416 (N_2416,N_2301,N_2340);
or U2417 (N_2417,N_2385,N_2364);
nand U2418 (N_2418,N_2338,N_2310);
nor U2419 (N_2419,N_2396,N_2324);
xor U2420 (N_2420,N_2322,N_2333);
nand U2421 (N_2421,N_2360,N_2379);
or U2422 (N_2422,N_2378,N_2345);
nor U2423 (N_2423,N_2313,N_2357);
or U2424 (N_2424,N_2341,N_2316);
nor U2425 (N_2425,N_2371,N_2351);
and U2426 (N_2426,N_2300,N_2306);
nand U2427 (N_2427,N_2307,N_2376);
nand U2428 (N_2428,N_2398,N_2372);
and U2429 (N_2429,N_2331,N_2384);
or U2430 (N_2430,N_2315,N_2382);
and U2431 (N_2431,N_2366,N_2348);
or U2432 (N_2432,N_2328,N_2334);
nand U2433 (N_2433,N_2380,N_2361);
or U2434 (N_2434,N_2375,N_2332);
nand U2435 (N_2435,N_2359,N_2318);
or U2436 (N_2436,N_2395,N_2399);
nand U2437 (N_2437,N_2352,N_2354);
nor U2438 (N_2438,N_2342,N_2383);
and U2439 (N_2439,N_2344,N_2311);
or U2440 (N_2440,N_2343,N_2390);
and U2441 (N_2441,N_2369,N_2373);
and U2442 (N_2442,N_2381,N_2323);
nor U2443 (N_2443,N_2362,N_2312);
and U2444 (N_2444,N_2319,N_2353);
nor U2445 (N_2445,N_2339,N_2320);
or U2446 (N_2446,N_2391,N_2325);
nand U2447 (N_2447,N_2304,N_2358);
nor U2448 (N_2448,N_2317,N_2389);
nor U2449 (N_2449,N_2388,N_2393);
and U2450 (N_2450,N_2308,N_2367);
and U2451 (N_2451,N_2363,N_2340);
nor U2452 (N_2452,N_2381,N_2375);
nand U2453 (N_2453,N_2380,N_2347);
nand U2454 (N_2454,N_2345,N_2390);
and U2455 (N_2455,N_2324,N_2359);
and U2456 (N_2456,N_2324,N_2337);
xnor U2457 (N_2457,N_2338,N_2332);
nand U2458 (N_2458,N_2327,N_2385);
nor U2459 (N_2459,N_2343,N_2385);
or U2460 (N_2460,N_2316,N_2366);
or U2461 (N_2461,N_2319,N_2379);
xor U2462 (N_2462,N_2311,N_2376);
and U2463 (N_2463,N_2328,N_2375);
or U2464 (N_2464,N_2307,N_2301);
nand U2465 (N_2465,N_2356,N_2348);
nand U2466 (N_2466,N_2362,N_2375);
nor U2467 (N_2467,N_2351,N_2379);
nor U2468 (N_2468,N_2389,N_2388);
and U2469 (N_2469,N_2312,N_2350);
nor U2470 (N_2470,N_2365,N_2362);
nor U2471 (N_2471,N_2354,N_2310);
nor U2472 (N_2472,N_2393,N_2336);
and U2473 (N_2473,N_2316,N_2373);
or U2474 (N_2474,N_2376,N_2366);
nand U2475 (N_2475,N_2338,N_2321);
or U2476 (N_2476,N_2393,N_2349);
nand U2477 (N_2477,N_2384,N_2398);
nand U2478 (N_2478,N_2316,N_2372);
or U2479 (N_2479,N_2388,N_2396);
and U2480 (N_2480,N_2370,N_2359);
or U2481 (N_2481,N_2308,N_2371);
nand U2482 (N_2482,N_2345,N_2319);
nor U2483 (N_2483,N_2384,N_2346);
nor U2484 (N_2484,N_2338,N_2393);
nand U2485 (N_2485,N_2320,N_2334);
nor U2486 (N_2486,N_2379,N_2332);
or U2487 (N_2487,N_2329,N_2388);
nor U2488 (N_2488,N_2362,N_2355);
or U2489 (N_2489,N_2365,N_2359);
nor U2490 (N_2490,N_2390,N_2384);
and U2491 (N_2491,N_2330,N_2370);
and U2492 (N_2492,N_2351,N_2370);
or U2493 (N_2493,N_2329,N_2339);
nand U2494 (N_2494,N_2393,N_2351);
nand U2495 (N_2495,N_2332,N_2342);
and U2496 (N_2496,N_2389,N_2338);
nand U2497 (N_2497,N_2325,N_2390);
nor U2498 (N_2498,N_2370,N_2317);
nand U2499 (N_2499,N_2364,N_2396);
or U2500 (N_2500,N_2404,N_2488);
and U2501 (N_2501,N_2465,N_2456);
nand U2502 (N_2502,N_2425,N_2418);
nand U2503 (N_2503,N_2431,N_2498);
and U2504 (N_2504,N_2476,N_2473);
nor U2505 (N_2505,N_2437,N_2478);
or U2506 (N_2506,N_2484,N_2499);
nor U2507 (N_2507,N_2426,N_2494);
nand U2508 (N_2508,N_2485,N_2451);
and U2509 (N_2509,N_2452,N_2496);
or U2510 (N_2510,N_2470,N_2443);
nand U2511 (N_2511,N_2413,N_2407);
or U2512 (N_2512,N_2475,N_2435);
or U2513 (N_2513,N_2439,N_2497);
and U2514 (N_2514,N_2448,N_2412);
nand U2515 (N_2515,N_2422,N_2408);
or U2516 (N_2516,N_2424,N_2416);
nor U2517 (N_2517,N_2491,N_2495);
nor U2518 (N_2518,N_2441,N_2467);
and U2519 (N_2519,N_2474,N_2483);
nor U2520 (N_2520,N_2487,N_2444);
nand U2521 (N_2521,N_2414,N_2460);
or U2522 (N_2522,N_2405,N_2489);
nand U2523 (N_2523,N_2410,N_2486);
nor U2524 (N_2524,N_2477,N_2461);
or U2525 (N_2525,N_2403,N_2417);
nand U2526 (N_2526,N_2490,N_2445);
or U2527 (N_2527,N_2419,N_2442);
or U2528 (N_2528,N_2415,N_2454);
and U2529 (N_2529,N_2469,N_2421);
and U2530 (N_2530,N_2453,N_2458);
and U2531 (N_2531,N_2446,N_2447);
and U2532 (N_2532,N_2429,N_2432);
nor U2533 (N_2533,N_2406,N_2423);
nor U2534 (N_2534,N_2400,N_2401);
or U2535 (N_2535,N_2472,N_2466);
nand U2536 (N_2536,N_2482,N_2433);
nor U2537 (N_2537,N_2464,N_2420);
xor U2538 (N_2538,N_2440,N_2457);
and U2539 (N_2539,N_2428,N_2479);
nand U2540 (N_2540,N_2430,N_2481);
nor U2541 (N_2541,N_2492,N_2436);
and U2542 (N_2542,N_2409,N_2462);
nand U2543 (N_2543,N_2434,N_2411);
nor U2544 (N_2544,N_2455,N_2459);
nand U2545 (N_2545,N_2463,N_2402);
and U2546 (N_2546,N_2471,N_2480);
nand U2547 (N_2547,N_2493,N_2468);
xor U2548 (N_2548,N_2449,N_2450);
or U2549 (N_2549,N_2438,N_2427);
and U2550 (N_2550,N_2439,N_2451);
nor U2551 (N_2551,N_2442,N_2420);
or U2552 (N_2552,N_2481,N_2494);
or U2553 (N_2553,N_2482,N_2472);
nor U2554 (N_2554,N_2422,N_2433);
nand U2555 (N_2555,N_2485,N_2407);
nor U2556 (N_2556,N_2423,N_2432);
nor U2557 (N_2557,N_2464,N_2435);
nand U2558 (N_2558,N_2481,N_2478);
nor U2559 (N_2559,N_2472,N_2408);
or U2560 (N_2560,N_2441,N_2472);
xor U2561 (N_2561,N_2457,N_2400);
nor U2562 (N_2562,N_2434,N_2450);
and U2563 (N_2563,N_2448,N_2481);
nand U2564 (N_2564,N_2477,N_2443);
and U2565 (N_2565,N_2404,N_2435);
or U2566 (N_2566,N_2496,N_2420);
or U2567 (N_2567,N_2443,N_2485);
nand U2568 (N_2568,N_2486,N_2408);
and U2569 (N_2569,N_2445,N_2464);
nand U2570 (N_2570,N_2409,N_2422);
nor U2571 (N_2571,N_2415,N_2433);
and U2572 (N_2572,N_2478,N_2444);
and U2573 (N_2573,N_2437,N_2471);
and U2574 (N_2574,N_2487,N_2489);
nand U2575 (N_2575,N_2437,N_2440);
nor U2576 (N_2576,N_2415,N_2416);
or U2577 (N_2577,N_2404,N_2406);
nor U2578 (N_2578,N_2421,N_2417);
nor U2579 (N_2579,N_2401,N_2445);
nor U2580 (N_2580,N_2475,N_2451);
nand U2581 (N_2581,N_2454,N_2436);
nand U2582 (N_2582,N_2419,N_2410);
and U2583 (N_2583,N_2482,N_2403);
and U2584 (N_2584,N_2472,N_2445);
nor U2585 (N_2585,N_2441,N_2449);
and U2586 (N_2586,N_2432,N_2458);
or U2587 (N_2587,N_2479,N_2482);
nand U2588 (N_2588,N_2453,N_2418);
nand U2589 (N_2589,N_2427,N_2421);
xor U2590 (N_2590,N_2448,N_2495);
nor U2591 (N_2591,N_2491,N_2446);
nand U2592 (N_2592,N_2457,N_2451);
nor U2593 (N_2593,N_2492,N_2401);
nor U2594 (N_2594,N_2427,N_2434);
nor U2595 (N_2595,N_2426,N_2465);
or U2596 (N_2596,N_2481,N_2400);
nor U2597 (N_2597,N_2448,N_2403);
nor U2598 (N_2598,N_2422,N_2496);
nor U2599 (N_2599,N_2458,N_2493);
nor U2600 (N_2600,N_2586,N_2508);
nand U2601 (N_2601,N_2550,N_2530);
or U2602 (N_2602,N_2592,N_2512);
nor U2603 (N_2603,N_2598,N_2504);
nor U2604 (N_2604,N_2558,N_2522);
nor U2605 (N_2605,N_2511,N_2525);
nor U2606 (N_2606,N_2572,N_2545);
nand U2607 (N_2607,N_2516,N_2531);
nor U2608 (N_2608,N_2595,N_2551);
nor U2609 (N_2609,N_2515,N_2500);
and U2610 (N_2610,N_2538,N_2555);
nand U2611 (N_2611,N_2503,N_2571);
or U2612 (N_2612,N_2528,N_2544);
and U2613 (N_2613,N_2510,N_2566);
nor U2614 (N_2614,N_2539,N_2573);
or U2615 (N_2615,N_2589,N_2523);
or U2616 (N_2616,N_2599,N_2518);
nor U2617 (N_2617,N_2554,N_2574);
and U2618 (N_2618,N_2564,N_2557);
or U2619 (N_2619,N_2524,N_2583);
nand U2620 (N_2620,N_2570,N_2556);
nor U2621 (N_2621,N_2547,N_2502);
or U2622 (N_2622,N_2563,N_2553);
and U2623 (N_2623,N_2535,N_2552);
or U2624 (N_2624,N_2529,N_2519);
or U2625 (N_2625,N_2596,N_2505);
nand U2626 (N_2626,N_2548,N_2517);
and U2627 (N_2627,N_2584,N_2579);
nand U2628 (N_2628,N_2533,N_2565);
nand U2629 (N_2629,N_2514,N_2567);
or U2630 (N_2630,N_2536,N_2540);
or U2631 (N_2631,N_2534,N_2526);
xnor U2632 (N_2632,N_2585,N_2587);
nor U2633 (N_2633,N_2521,N_2513);
or U2634 (N_2634,N_2590,N_2542);
and U2635 (N_2635,N_2506,N_2575);
nand U2636 (N_2636,N_2507,N_2569);
or U2637 (N_2637,N_2581,N_2561);
or U2638 (N_2638,N_2568,N_2520);
and U2639 (N_2639,N_2578,N_2560);
nand U2640 (N_2640,N_2591,N_2509);
nand U2641 (N_2641,N_2537,N_2582);
nand U2642 (N_2642,N_2577,N_2588);
or U2643 (N_2643,N_2546,N_2580);
nor U2644 (N_2644,N_2594,N_2501);
nor U2645 (N_2645,N_2562,N_2527);
and U2646 (N_2646,N_2541,N_2576);
nor U2647 (N_2647,N_2549,N_2593);
nand U2648 (N_2648,N_2543,N_2559);
nor U2649 (N_2649,N_2532,N_2597);
or U2650 (N_2650,N_2572,N_2590);
nor U2651 (N_2651,N_2590,N_2557);
nand U2652 (N_2652,N_2548,N_2562);
nor U2653 (N_2653,N_2543,N_2532);
and U2654 (N_2654,N_2573,N_2507);
nor U2655 (N_2655,N_2584,N_2537);
or U2656 (N_2656,N_2589,N_2569);
and U2657 (N_2657,N_2511,N_2581);
xor U2658 (N_2658,N_2550,N_2507);
nor U2659 (N_2659,N_2597,N_2580);
nand U2660 (N_2660,N_2532,N_2529);
nor U2661 (N_2661,N_2534,N_2545);
and U2662 (N_2662,N_2566,N_2563);
or U2663 (N_2663,N_2515,N_2510);
and U2664 (N_2664,N_2526,N_2517);
nor U2665 (N_2665,N_2595,N_2530);
nor U2666 (N_2666,N_2585,N_2512);
and U2667 (N_2667,N_2568,N_2565);
nand U2668 (N_2668,N_2503,N_2551);
and U2669 (N_2669,N_2524,N_2561);
nand U2670 (N_2670,N_2599,N_2511);
or U2671 (N_2671,N_2549,N_2585);
nor U2672 (N_2672,N_2501,N_2522);
or U2673 (N_2673,N_2580,N_2505);
nand U2674 (N_2674,N_2572,N_2512);
nor U2675 (N_2675,N_2516,N_2506);
nor U2676 (N_2676,N_2518,N_2574);
or U2677 (N_2677,N_2506,N_2546);
nand U2678 (N_2678,N_2558,N_2571);
and U2679 (N_2679,N_2506,N_2595);
nand U2680 (N_2680,N_2507,N_2590);
nor U2681 (N_2681,N_2577,N_2532);
and U2682 (N_2682,N_2591,N_2558);
nor U2683 (N_2683,N_2571,N_2590);
or U2684 (N_2684,N_2525,N_2514);
or U2685 (N_2685,N_2570,N_2583);
nor U2686 (N_2686,N_2573,N_2581);
or U2687 (N_2687,N_2549,N_2569);
nor U2688 (N_2688,N_2556,N_2526);
nor U2689 (N_2689,N_2595,N_2574);
nand U2690 (N_2690,N_2550,N_2515);
and U2691 (N_2691,N_2540,N_2587);
nand U2692 (N_2692,N_2544,N_2581);
or U2693 (N_2693,N_2560,N_2528);
or U2694 (N_2694,N_2596,N_2509);
nor U2695 (N_2695,N_2510,N_2567);
or U2696 (N_2696,N_2500,N_2595);
nand U2697 (N_2697,N_2559,N_2589);
nor U2698 (N_2698,N_2576,N_2565);
nand U2699 (N_2699,N_2599,N_2534);
or U2700 (N_2700,N_2639,N_2675);
and U2701 (N_2701,N_2661,N_2627);
nor U2702 (N_2702,N_2643,N_2679);
and U2703 (N_2703,N_2640,N_2688);
and U2704 (N_2704,N_2648,N_2670);
and U2705 (N_2705,N_2676,N_2609);
nand U2706 (N_2706,N_2645,N_2642);
nand U2707 (N_2707,N_2697,N_2604);
nand U2708 (N_2708,N_2618,N_2600);
and U2709 (N_2709,N_2625,N_2685);
nor U2710 (N_2710,N_2692,N_2665);
xnor U2711 (N_2711,N_2674,N_2690);
and U2712 (N_2712,N_2686,N_2696);
nor U2713 (N_2713,N_2647,N_2663);
and U2714 (N_2714,N_2624,N_2681);
or U2715 (N_2715,N_2636,N_2629);
nand U2716 (N_2716,N_2602,N_2694);
nor U2717 (N_2717,N_2605,N_2668);
nand U2718 (N_2718,N_2666,N_2684);
nand U2719 (N_2719,N_2673,N_2650);
nand U2720 (N_2720,N_2606,N_2626);
or U2721 (N_2721,N_2659,N_2635);
and U2722 (N_2722,N_2691,N_2695);
nand U2723 (N_2723,N_2613,N_2693);
nand U2724 (N_2724,N_2680,N_2628);
nand U2725 (N_2725,N_2644,N_2633);
or U2726 (N_2726,N_2699,N_2608);
nor U2727 (N_2727,N_2652,N_2638);
and U2728 (N_2728,N_2667,N_2614);
or U2729 (N_2729,N_2641,N_2630);
and U2730 (N_2730,N_2617,N_2672);
and U2731 (N_2731,N_2664,N_2634);
and U2732 (N_2732,N_2610,N_2607);
or U2733 (N_2733,N_2616,N_2603);
and U2734 (N_2734,N_2615,N_2669);
nor U2735 (N_2735,N_2649,N_2646);
and U2736 (N_2736,N_2623,N_2620);
and U2737 (N_2737,N_2671,N_2689);
nor U2738 (N_2738,N_2632,N_2682);
or U2739 (N_2739,N_2612,N_2678);
or U2740 (N_2740,N_2654,N_2622);
nor U2741 (N_2741,N_2677,N_2657);
or U2742 (N_2742,N_2653,N_2687);
or U2743 (N_2743,N_2698,N_2656);
nor U2744 (N_2744,N_2651,N_2619);
and U2745 (N_2745,N_2658,N_2683);
nand U2746 (N_2746,N_2621,N_2662);
or U2747 (N_2747,N_2637,N_2601);
and U2748 (N_2748,N_2655,N_2611);
and U2749 (N_2749,N_2631,N_2660);
nor U2750 (N_2750,N_2652,N_2688);
nor U2751 (N_2751,N_2667,N_2604);
or U2752 (N_2752,N_2640,N_2691);
or U2753 (N_2753,N_2609,N_2602);
and U2754 (N_2754,N_2625,N_2695);
nor U2755 (N_2755,N_2609,N_2679);
nand U2756 (N_2756,N_2663,N_2640);
nand U2757 (N_2757,N_2661,N_2619);
nor U2758 (N_2758,N_2685,N_2653);
and U2759 (N_2759,N_2613,N_2628);
or U2760 (N_2760,N_2676,N_2605);
nor U2761 (N_2761,N_2672,N_2634);
and U2762 (N_2762,N_2656,N_2687);
nor U2763 (N_2763,N_2664,N_2691);
nor U2764 (N_2764,N_2605,N_2634);
xor U2765 (N_2765,N_2623,N_2601);
and U2766 (N_2766,N_2661,N_2650);
nor U2767 (N_2767,N_2656,N_2699);
or U2768 (N_2768,N_2653,N_2609);
and U2769 (N_2769,N_2677,N_2663);
or U2770 (N_2770,N_2688,N_2606);
nand U2771 (N_2771,N_2661,N_2665);
nand U2772 (N_2772,N_2628,N_2610);
or U2773 (N_2773,N_2600,N_2699);
nand U2774 (N_2774,N_2604,N_2603);
nand U2775 (N_2775,N_2651,N_2697);
and U2776 (N_2776,N_2648,N_2626);
and U2777 (N_2777,N_2601,N_2628);
xnor U2778 (N_2778,N_2608,N_2668);
and U2779 (N_2779,N_2632,N_2645);
and U2780 (N_2780,N_2630,N_2615);
nand U2781 (N_2781,N_2655,N_2688);
and U2782 (N_2782,N_2672,N_2676);
and U2783 (N_2783,N_2637,N_2602);
xor U2784 (N_2784,N_2668,N_2671);
and U2785 (N_2785,N_2691,N_2699);
nand U2786 (N_2786,N_2628,N_2626);
nand U2787 (N_2787,N_2628,N_2627);
nor U2788 (N_2788,N_2670,N_2630);
or U2789 (N_2789,N_2628,N_2600);
nand U2790 (N_2790,N_2683,N_2688);
and U2791 (N_2791,N_2613,N_2664);
nor U2792 (N_2792,N_2600,N_2637);
nand U2793 (N_2793,N_2627,N_2678);
nor U2794 (N_2794,N_2618,N_2623);
or U2795 (N_2795,N_2644,N_2666);
nand U2796 (N_2796,N_2635,N_2617);
nor U2797 (N_2797,N_2676,N_2643);
nand U2798 (N_2798,N_2653,N_2661);
or U2799 (N_2799,N_2697,N_2688);
nand U2800 (N_2800,N_2783,N_2730);
or U2801 (N_2801,N_2748,N_2727);
nand U2802 (N_2802,N_2705,N_2763);
and U2803 (N_2803,N_2747,N_2788);
nor U2804 (N_2804,N_2790,N_2741);
or U2805 (N_2805,N_2767,N_2765);
nand U2806 (N_2806,N_2782,N_2724);
nand U2807 (N_2807,N_2738,N_2701);
and U2808 (N_2808,N_2789,N_2770);
or U2809 (N_2809,N_2754,N_2710);
nand U2810 (N_2810,N_2713,N_2784);
nor U2811 (N_2811,N_2703,N_2775);
and U2812 (N_2812,N_2781,N_2744);
nor U2813 (N_2813,N_2752,N_2751);
or U2814 (N_2814,N_2786,N_2702);
nand U2815 (N_2815,N_2750,N_2795);
nor U2816 (N_2816,N_2712,N_2773);
and U2817 (N_2817,N_2761,N_2745);
nand U2818 (N_2818,N_2711,N_2715);
nor U2819 (N_2819,N_2785,N_2728);
or U2820 (N_2820,N_2708,N_2725);
or U2821 (N_2821,N_2778,N_2777);
nor U2822 (N_2822,N_2739,N_2706);
and U2823 (N_2823,N_2719,N_2764);
nand U2824 (N_2824,N_2792,N_2735);
nor U2825 (N_2825,N_2793,N_2717);
and U2826 (N_2826,N_2740,N_2716);
and U2827 (N_2827,N_2759,N_2731);
nor U2828 (N_2828,N_2758,N_2753);
or U2829 (N_2829,N_2772,N_2714);
nor U2830 (N_2830,N_2776,N_2771);
nor U2831 (N_2831,N_2762,N_2755);
nor U2832 (N_2832,N_2760,N_2707);
or U2833 (N_2833,N_2720,N_2796);
or U2834 (N_2834,N_2718,N_2791);
nor U2835 (N_2835,N_2787,N_2766);
xnor U2836 (N_2836,N_2726,N_2722);
and U2837 (N_2837,N_2729,N_2700);
nor U2838 (N_2838,N_2734,N_2799);
xor U2839 (N_2839,N_2743,N_2749);
nand U2840 (N_2840,N_2737,N_2746);
or U2841 (N_2841,N_2798,N_2797);
nor U2842 (N_2842,N_2721,N_2757);
or U2843 (N_2843,N_2732,N_2780);
or U2844 (N_2844,N_2709,N_2794);
or U2845 (N_2845,N_2768,N_2704);
nand U2846 (N_2846,N_2736,N_2733);
nor U2847 (N_2847,N_2756,N_2774);
nor U2848 (N_2848,N_2723,N_2769);
nor U2849 (N_2849,N_2742,N_2779);
nand U2850 (N_2850,N_2749,N_2716);
and U2851 (N_2851,N_2768,N_2788);
nand U2852 (N_2852,N_2700,N_2737);
or U2853 (N_2853,N_2795,N_2797);
nor U2854 (N_2854,N_2762,N_2702);
nor U2855 (N_2855,N_2727,N_2768);
nand U2856 (N_2856,N_2709,N_2718);
or U2857 (N_2857,N_2743,N_2791);
nor U2858 (N_2858,N_2712,N_2748);
and U2859 (N_2859,N_2715,N_2771);
and U2860 (N_2860,N_2795,N_2759);
nor U2861 (N_2861,N_2714,N_2749);
nand U2862 (N_2862,N_2742,N_2717);
or U2863 (N_2863,N_2783,N_2737);
nand U2864 (N_2864,N_2729,N_2716);
or U2865 (N_2865,N_2704,N_2744);
or U2866 (N_2866,N_2716,N_2717);
xnor U2867 (N_2867,N_2767,N_2787);
nand U2868 (N_2868,N_2765,N_2776);
and U2869 (N_2869,N_2716,N_2786);
and U2870 (N_2870,N_2767,N_2737);
nor U2871 (N_2871,N_2760,N_2706);
and U2872 (N_2872,N_2759,N_2758);
and U2873 (N_2873,N_2700,N_2768);
and U2874 (N_2874,N_2783,N_2777);
nand U2875 (N_2875,N_2700,N_2799);
and U2876 (N_2876,N_2724,N_2735);
nor U2877 (N_2877,N_2731,N_2717);
or U2878 (N_2878,N_2796,N_2725);
nor U2879 (N_2879,N_2752,N_2757);
nand U2880 (N_2880,N_2728,N_2709);
and U2881 (N_2881,N_2769,N_2743);
nor U2882 (N_2882,N_2715,N_2774);
nand U2883 (N_2883,N_2778,N_2711);
and U2884 (N_2884,N_2767,N_2795);
nand U2885 (N_2885,N_2744,N_2726);
nand U2886 (N_2886,N_2745,N_2719);
and U2887 (N_2887,N_2764,N_2737);
nand U2888 (N_2888,N_2746,N_2781);
nor U2889 (N_2889,N_2721,N_2795);
or U2890 (N_2890,N_2794,N_2780);
or U2891 (N_2891,N_2769,N_2762);
nand U2892 (N_2892,N_2728,N_2764);
or U2893 (N_2893,N_2727,N_2795);
xnor U2894 (N_2894,N_2702,N_2794);
or U2895 (N_2895,N_2764,N_2708);
and U2896 (N_2896,N_2710,N_2775);
and U2897 (N_2897,N_2798,N_2727);
nand U2898 (N_2898,N_2718,N_2734);
or U2899 (N_2899,N_2702,N_2759);
or U2900 (N_2900,N_2892,N_2876);
nor U2901 (N_2901,N_2853,N_2834);
xnor U2902 (N_2902,N_2840,N_2804);
and U2903 (N_2903,N_2822,N_2809);
or U2904 (N_2904,N_2819,N_2894);
or U2905 (N_2905,N_2813,N_2868);
nand U2906 (N_2906,N_2856,N_2878);
nand U2907 (N_2907,N_2869,N_2865);
or U2908 (N_2908,N_2898,N_2891);
or U2909 (N_2909,N_2827,N_2854);
and U2910 (N_2910,N_2860,N_2800);
or U2911 (N_2911,N_2855,N_2887);
nand U2912 (N_2912,N_2806,N_2862);
and U2913 (N_2913,N_2875,N_2835);
and U2914 (N_2914,N_2814,N_2803);
or U2915 (N_2915,N_2881,N_2861);
and U2916 (N_2916,N_2820,N_2808);
nor U2917 (N_2917,N_2851,N_2897);
or U2918 (N_2918,N_2818,N_2866);
or U2919 (N_2919,N_2810,N_2848);
and U2920 (N_2920,N_2849,N_2859);
nand U2921 (N_2921,N_2807,N_2880);
nand U2922 (N_2922,N_2852,N_2872);
nand U2923 (N_2923,N_2850,N_2847);
and U2924 (N_2924,N_2864,N_2817);
nand U2925 (N_2925,N_2885,N_2844);
nor U2926 (N_2926,N_2842,N_2833);
nand U2927 (N_2927,N_2899,N_2893);
and U2928 (N_2928,N_2873,N_2883);
nor U2929 (N_2929,N_2829,N_2838);
and U2930 (N_2930,N_2871,N_2890);
nand U2931 (N_2931,N_2828,N_2889);
or U2932 (N_2932,N_2879,N_2858);
or U2933 (N_2933,N_2884,N_2826);
nor U2934 (N_2934,N_2812,N_2867);
and U2935 (N_2935,N_2801,N_2863);
or U2936 (N_2936,N_2836,N_2839);
nor U2937 (N_2937,N_2805,N_2888);
nor U2938 (N_2938,N_2825,N_2832);
and U2939 (N_2939,N_2857,N_2824);
nand U2940 (N_2940,N_2823,N_2886);
nand U2941 (N_2941,N_2895,N_2837);
nor U2942 (N_2942,N_2846,N_2816);
or U2943 (N_2943,N_2882,N_2811);
and U2944 (N_2944,N_2815,N_2896);
nand U2945 (N_2945,N_2845,N_2874);
and U2946 (N_2946,N_2831,N_2841);
and U2947 (N_2947,N_2870,N_2802);
and U2948 (N_2948,N_2843,N_2830);
xnor U2949 (N_2949,N_2877,N_2821);
or U2950 (N_2950,N_2861,N_2806);
or U2951 (N_2951,N_2858,N_2850);
or U2952 (N_2952,N_2816,N_2872);
and U2953 (N_2953,N_2832,N_2883);
and U2954 (N_2954,N_2826,N_2852);
or U2955 (N_2955,N_2854,N_2816);
nand U2956 (N_2956,N_2829,N_2867);
and U2957 (N_2957,N_2849,N_2810);
nor U2958 (N_2958,N_2856,N_2830);
nand U2959 (N_2959,N_2850,N_2869);
nor U2960 (N_2960,N_2804,N_2803);
nand U2961 (N_2961,N_2895,N_2873);
nor U2962 (N_2962,N_2849,N_2845);
nand U2963 (N_2963,N_2843,N_2859);
and U2964 (N_2964,N_2860,N_2892);
nand U2965 (N_2965,N_2811,N_2898);
and U2966 (N_2966,N_2805,N_2898);
nand U2967 (N_2967,N_2838,N_2821);
and U2968 (N_2968,N_2866,N_2869);
nand U2969 (N_2969,N_2860,N_2845);
nor U2970 (N_2970,N_2887,N_2850);
nand U2971 (N_2971,N_2807,N_2862);
nand U2972 (N_2972,N_2805,N_2867);
nand U2973 (N_2973,N_2819,N_2868);
and U2974 (N_2974,N_2807,N_2866);
or U2975 (N_2975,N_2837,N_2884);
nand U2976 (N_2976,N_2886,N_2876);
or U2977 (N_2977,N_2887,N_2852);
or U2978 (N_2978,N_2869,N_2842);
nand U2979 (N_2979,N_2818,N_2803);
and U2980 (N_2980,N_2885,N_2890);
xnor U2981 (N_2981,N_2861,N_2845);
nor U2982 (N_2982,N_2879,N_2842);
and U2983 (N_2983,N_2849,N_2802);
nor U2984 (N_2984,N_2883,N_2863);
nor U2985 (N_2985,N_2863,N_2884);
nand U2986 (N_2986,N_2894,N_2841);
nor U2987 (N_2987,N_2848,N_2819);
nand U2988 (N_2988,N_2851,N_2811);
and U2989 (N_2989,N_2843,N_2888);
nand U2990 (N_2990,N_2867,N_2824);
and U2991 (N_2991,N_2862,N_2872);
and U2992 (N_2992,N_2819,N_2849);
nor U2993 (N_2993,N_2861,N_2814);
or U2994 (N_2994,N_2819,N_2885);
nor U2995 (N_2995,N_2806,N_2856);
nor U2996 (N_2996,N_2851,N_2849);
nor U2997 (N_2997,N_2885,N_2894);
or U2998 (N_2998,N_2808,N_2872);
nand U2999 (N_2999,N_2891,N_2873);
and UO_0 (O_0,N_2903,N_2931);
nand UO_1 (O_1,N_2946,N_2963);
nand UO_2 (O_2,N_2913,N_2923);
or UO_3 (O_3,N_2935,N_2916);
xor UO_4 (O_4,N_2978,N_2995);
or UO_5 (O_5,N_2981,N_2970);
nor UO_6 (O_6,N_2974,N_2956);
nand UO_7 (O_7,N_2993,N_2934);
or UO_8 (O_8,N_2914,N_2959);
and UO_9 (O_9,N_2911,N_2945);
nor UO_10 (O_10,N_2984,N_2969);
nor UO_11 (O_11,N_2907,N_2972);
nand UO_12 (O_12,N_2988,N_2926);
and UO_13 (O_13,N_2941,N_2998);
nand UO_14 (O_14,N_2976,N_2932);
or UO_15 (O_15,N_2922,N_2975);
and UO_16 (O_16,N_2902,N_2912);
and UO_17 (O_17,N_2989,N_2985);
nand UO_18 (O_18,N_2944,N_2929);
and UO_19 (O_19,N_2971,N_2937);
or UO_20 (O_20,N_2953,N_2982);
or UO_21 (O_21,N_2938,N_2983);
nand UO_22 (O_22,N_2901,N_2994);
nand UO_23 (O_23,N_2909,N_2980);
nand UO_24 (O_24,N_2967,N_2962);
nor UO_25 (O_25,N_2952,N_2947);
nand UO_26 (O_26,N_2979,N_2992);
or UO_27 (O_27,N_2930,N_2900);
nor UO_28 (O_28,N_2951,N_2990);
and UO_29 (O_29,N_2957,N_2966);
or UO_30 (O_30,N_2997,N_2936);
and UO_31 (O_31,N_2977,N_2910);
and UO_32 (O_32,N_2955,N_2954);
nand UO_33 (O_33,N_2986,N_2961);
and UO_34 (O_34,N_2968,N_2924);
or UO_35 (O_35,N_2904,N_2921);
or UO_36 (O_36,N_2958,N_2987);
or UO_37 (O_37,N_2948,N_2996);
or UO_38 (O_38,N_2973,N_2918);
nand UO_39 (O_39,N_2915,N_2991);
nand UO_40 (O_40,N_2927,N_2965);
xor UO_41 (O_41,N_2919,N_2960);
or UO_42 (O_42,N_2933,N_2906);
and UO_43 (O_43,N_2940,N_2943);
or UO_44 (O_44,N_2942,N_2939);
or UO_45 (O_45,N_2925,N_2950);
nor UO_46 (O_46,N_2928,N_2999);
and UO_47 (O_47,N_2905,N_2917);
nand UO_48 (O_48,N_2908,N_2920);
nand UO_49 (O_49,N_2949,N_2964);
nor UO_50 (O_50,N_2934,N_2907);
nor UO_51 (O_51,N_2950,N_2936);
nand UO_52 (O_52,N_2930,N_2974);
and UO_53 (O_53,N_2902,N_2995);
nand UO_54 (O_54,N_2952,N_2965);
or UO_55 (O_55,N_2925,N_2952);
nand UO_56 (O_56,N_2971,N_2951);
or UO_57 (O_57,N_2968,N_2983);
or UO_58 (O_58,N_2974,N_2987);
nand UO_59 (O_59,N_2986,N_2969);
nor UO_60 (O_60,N_2988,N_2930);
and UO_61 (O_61,N_2922,N_2971);
nand UO_62 (O_62,N_2912,N_2959);
nor UO_63 (O_63,N_2922,N_2936);
nor UO_64 (O_64,N_2959,N_2947);
and UO_65 (O_65,N_2927,N_2992);
nor UO_66 (O_66,N_2917,N_2932);
or UO_67 (O_67,N_2911,N_2929);
and UO_68 (O_68,N_2952,N_2988);
or UO_69 (O_69,N_2947,N_2992);
nand UO_70 (O_70,N_2997,N_2947);
nor UO_71 (O_71,N_2928,N_2923);
xnor UO_72 (O_72,N_2990,N_2904);
and UO_73 (O_73,N_2966,N_2903);
nor UO_74 (O_74,N_2992,N_2980);
or UO_75 (O_75,N_2995,N_2990);
nor UO_76 (O_76,N_2984,N_2974);
or UO_77 (O_77,N_2925,N_2996);
nand UO_78 (O_78,N_2905,N_2912);
and UO_79 (O_79,N_2975,N_2946);
nor UO_80 (O_80,N_2944,N_2911);
nor UO_81 (O_81,N_2949,N_2938);
and UO_82 (O_82,N_2904,N_2909);
and UO_83 (O_83,N_2985,N_2964);
or UO_84 (O_84,N_2969,N_2937);
nor UO_85 (O_85,N_2935,N_2985);
or UO_86 (O_86,N_2962,N_2919);
nor UO_87 (O_87,N_2974,N_2964);
or UO_88 (O_88,N_2952,N_2995);
nor UO_89 (O_89,N_2962,N_2925);
or UO_90 (O_90,N_2997,N_2991);
nand UO_91 (O_91,N_2903,N_2963);
nand UO_92 (O_92,N_2921,N_2981);
or UO_93 (O_93,N_2908,N_2911);
xor UO_94 (O_94,N_2955,N_2928);
or UO_95 (O_95,N_2916,N_2952);
nor UO_96 (O_96,N_2984,N_2915);
and UO_97 (O_97,N_2954,N_2900);
xnor UO_98 (O_98,N_2971,N_2923);
nand UO_99 (O_99,N_2985,N_2979);
nor UO_100 (O_100,N_2984,N_2962);
xor UO_101 (O_101,N_2904,N_2919);
nand UO_102 (O_102,N_2961,N_2915);
and UO_103 (O_103,N_2934,N_2955);
nor UO_104 (O_104,N_2973,N_2917);
and UO_105 (O_105,N_2905,N_2993);
nand UO_106 (O_106,N_2959,N_2901);
nor UO_107 (O_107,N_2929,N_2919);
nand UO_108 (O_108,N_2948,N_2960);
and UO_109 (O_109,N_2919,N_2990);
or UO_110 (O_110,N_2957,N_2982);
nor UO_111 (O_111,N_2946,N_2943);
and UO_112 (O_112,N_2904,N_2971);
nand UO_113 (O_113,N_2911,N_2931);
nor UO_114 (O_114,N_2990,N_2942);
nor UO_115 (O_115,N_2943,N_2948);
and UO_116 (O_116,N_2914,N_2930);
or UO_117 (O_117,N_2928,N_2968);
and UO_118 (O_118,N_2922,N_2996);
or UO_119 (O_119,N_2973,N_2998);
xor UO_120 (O_120,N_2972,N_2939);
nor UO_121 (O_121,N_2963,N_2910);
nor UO_122 (O_122,N_2920,N_2968);
nor UO_123 (O_123,N_2984,N_2911);
or UO_124 (O_124,N_2948,N_2917);
nor UO_125 (O_125,N_2947,N_2977);
or UO_126 (O_126,N_2917,N_2946);
nand UO_127 (O_127,N_2915,N_2979);
nor UO_128 (O_128,N_2948,N_2912);
nand UO_129 (O_129,N_2931,N_2991);
nand UO_130 (O_130,N_2980,N_2935);
nand UO_131 (O_131,N_2945,N_2997);
or UO_132 (O_132,N_2908,N_2988);
and UO_133 (O_133,N_2939,N_2901);
nand UO_134 (O_134,N_2923,N_2944);
nand UO_135 (O_135,N_2916,N_2999);
xor UO_136 (O_136,N_2969,N_2926);
or UO_137 (O_137,N_2948,N_2967);
or UO_138 (O_138,N_2914,N_2951);
nand UO_139 (O_139,N_2956,N_2921);
and UO_140 (O_140,N_2943,N_2952);
nand UO_141 (O_141,N_2944,N_2966);
and UO_142 (O_142,N_2906,N_2939);
and UO_143 (O_143,N_2997,N_2987);
or UO_144 (O_144,N_2944,N_2948);
or UO_145 (O_145,N_2988,N_2956);
and UO_146 (O_146,N_2926,N_2975);
or UO_147 (O_147,N_2944,N_2922);
and UO_148 (O_148,N_2923,N_2982);
nand UO_149 (O_149,N_2906,N_2947);
or UO_150 (O_150,N_2985,N_2950);
and UO_151 (O_151,N_2914,N_2981);
or UO_152 (O_152,N_2923,N_2947);
and UO_153 (O_153,N_2964,N_2900);
nand UO_154 (O_154,N_2961,N_2960);
or UO_155 (O_155,N_2976,N_2921);
nand UO_156 (O_156,N_2971,N_2987);
nor UO_157 (O_157,N_2906,N_2903);
nand UO_158 (O_158,N_2970,N_2919);
and UO_159 (O_159,N_2974,N_2953);
nor UO_160 (O_160,N_2951,N_2984);
and UO_161 (O_161,N_2997,N_2914);
and UO_162 (O_162,N_2976,N_2963);
nand UO_163 (O_163,N_2905,N_2903);
or UO_164 (O_164,N_2993,N_2945);
or UO_165 (O_165,N_2932,N_2909);
or UO_166 (O_166,N_2983,N_2913);
and UO_167 (O_167,N_2989,N_2921);
nand UO_168 (O_168,N_2986,N_2906);
or UO_169 (O_169,N_2923,N_2958);
xor UO_170 (O_170,N_2918,N_2974);
nor UO_171 (O_171,N_2948,N_2921);
nand UO_172 (O_172,N_2980,N_2928);
nand UO_173 (O_173,N_2985,N_2988);
or UO_174 (O_174,N_2987,N_2966);
nand UO_175 (O_175,N_2966,N_2946);
nor UO_176 (O_176,N_2935,N_2943);
or UO_177 (O_177,N_2957,N_2946);
and UO_178 (O_178,N_2958,N_2922);
and UO_179 (O_179,N_2975,N_2968);
nor UO_180 (O_180,N_2914,N_2940);
and UO_181 (O_181,N_2923,N_2945);
and UO_182 (O_182,N_2988,N_2922);
and UO_183 (O_183,N_2907,N_2923);
nor UO_184 (O_184,N_2957,N_2914);
xnor UO_185 (O_185,N_2906,N_2950);
nor UO_186 (O_186,N_2958,N_2949);
nor UO_187 (O_187,N_2927,N_2991);
or UO_188 (O_188,N_2914,N_2938);
nand UO_189 (O_189,N_2974,N_2959);
nand UO_190 (O_190,N_2964,N_2970);
or UO_191 (O_191,N_2941,N_2983);
or UO_192 (O_192,N_2979,N_2922);
or UO_193 (O_193,N_2932,N_2979);
nand UO_194 (O_194,N_2950,N_2979);
or UO_195 (O_195,N_2938,N_2990);
and UO_196 (O_196,N_2906,N_2957);
or UO_197 (O_197,N_2957,N_2907);
and UO_198 (O_198,N_2992,N_2985);
or UO_199 (O_199,N_2907,N_2994);
nand UO_200 (O_200,N_2978,N_2957);
and UO_201 (O_201,N_2952,N_2997);
nand UO_202 (O_202,N_2975,N_2969);
nor UO_203 (O_203,N_2928,N_2916);
and UO_204 (O_204,N_2946,N_2936);
or UO_205 (O_205,N_2971,N_2967);
and UO_206 (O_206,N_2922,N_2950);
nor UO_207 (O_207,N_2993,N_2920);
and UO_208 (O_208,N_2914,N_2946);
nand UO_209 (O_209,N_2909,N_2933);
nor UO_210 (O_210,N_2954,N_2991);
nand UO_211 (O_211,N_2930,N_2916);
nand UO_212 (O_212,N_2906,N_2980);
nor UO_213 (O_213,N_2967,N_2922);
and UO_214 (O_214,N_2954,N_2909);
or UO_215 (O_215,N_2995,N_2904);
or UO_216 (O_216,N_2927,N_2969);
nand UO_217 (O_217,N_2946,N_2999);
or UO_218 (O_218,N_2948,N_2904);
nor UO_219 (O_219,N_2980,N_2924);
or UO_220 (O_220,N_2935,N_2987);
or UO_221 (O_221,N_2901,N_2991);
nand UO_222 (O_222,N_2961,N_2903);
nand UO_223 (O_223,N_2916,N_2956);
and UO_224 (O_224,N_2935,N_2982);
or UO_225 (O_225,N_2966,N_2965);
nor UO_226 (O_226,N_2972,N_2976);
nand UO_227 (O_227,N_2992,N_2955);
or UO_228 (O_228,N_2985,N_2975);
nand UO_229 (O_229,N_2988,N_2948);
nand UO_230 (O_230,N_2900,N_2984);
nand UO_231 (O_231,N_2940,N_2967);
and UO_232 (O_232,N_2991,N_2994);
nand UO_233 (O_233,N_2973,N_2987);
and UO_234 (O_234,N_2984,N_2920);
and UO_235 (O_235,N_2917,N_2943);
and UO_236 (O_236,N_2936,N_2913);
and UO_237 (O_237,N_2965,N_2907);
nor UO_238 (O_238,N_2903,N_2922);
nand UO_239 (O_239,N_2946,N_2976);
or UO_240 (O_240,N_2924,N_2974);
and UO_241 (O_241,N_2944,N_2997);
nor UO_242 (O_242,N_2966,N_2999);
nor UO_243 (O_243,N_2986,N_2947);
nor UO_244 (O_244,N_2980,N_2968);
nor UO_245 (O_245,N_2979,N_2946);
nor UO_246 (O_246,N_2943,N_2958);
nand UO_247 (O_247,N_2914,N_2954);
or UO_248 (O_248,N_2990,N_2963);
or UO_249 (O_249,N_2939,N_2964);
nand UO_250 (O_250,N_2960,N_2940);
or UO_251 (O_251,N_2962,N_2907);
nand UO_252 (O_252,N_2995,N_2949);
or UO_253 (O_253,N_2915,N_2977);
nor UO_254 (O_254,N_2902,N_2907);
xnor UO_255 (O_255,N_2910,N_2961);
nand UO_256 (O_256,N_2945,N_2964);
nor UO_257 (O_257,N_2981,N_2922);
nand UO_258 (O_258,N_2952,N_2900);
or UO_259 (O_259,N_2952,N_2986);
and UO_260 (O_260,N_2976,N_2900);
nand UO_261 (O_261,N_2908,N_2952);
nand UO_262 (O_262,N_2994,N_2909);
and UO_263 (O_263,N_2938,N_2916);
or UO_264 (O_264,N_2988,N_2992);
nor UO_265 (O_265,N_2943,N_2939);
and UO_266 (O_266,N_2996,N_2992);
nor UO_267 (O_267,N_2947,N_2901);
and UO_268 (O_268,N_2939,N_2933);
nor UO_269 (O_269,N_2967,N_2908);
or UO_270 (O_270,N_2951,N_2915);
nand UO_271 (O_271,N_2976,N_2948);
xor UO_272 (O_272,N_2974,N_2990);
or UO_273 (O_273,N_2980,N_2937);
or UO_274 (O_274,N_2956,N_2914);
and UO_275 (O_275,N_2913,N_2987);
nand UO_276 (O_276,N_2977,N_2963);
and UO_277 (O_277,N_2991,N_2929);
nor UO_278 (O_278,N_2962,N_2910);
and UO_279 (O_279,N_2939,N_2998);
or UO_280 (O_280,N_2999,N_2961);
or UO_281 (O_281,N_2987,N_2929);
or UO_282 (O_282,N_2973,N_2964);
nand UO_283 (O_283,N_2966,N_2967);
nor UO_284 (O_284,N_2944,N_2986);
nor UO_285 (O_285,N_2948,N_2937);
nor UO_286 (O_286,N_2948,N_2991);
and UO_287 (O_287,N_2929,N_2993);
or UO_288 (O_288,N_2960,N_2979);
nor UO_289 (O_289,N_2996,N_2938);
xnor UO_290 (O_290,N_2973,N_2938);
nand UO_291 (O_291,N_2922,N_2985);
xnor UO_292 (O_292,N_2924,N_2972);
and UO_293 (O_293,N_2968,N_2958);
or UO_294 (O_294,N_2952,N_2940);
nor UO_295 (O_295,N_2941,N_2920);
or UO_296 (O_296,N_2922,N_2948);
nor UO_297 (O_297,N_2967,N_2904);
and UO_298 (O_298,N_2956,N_2966);
and UO_299 (O_299,N_2919,N_2900);
nand UO_300 (O_300,N_2910,N_2957);
nand UO_301 (O_301,N_2961,N_2938);
and UO_302 (O_302,N_2900,N_2916);
nand UO_303 (O_303,N_2938,N_2998);
nor UO_304 (O_304,N_2950,N_2920);
nor UO_305 (O_305,N_2945,N_2950);
nor UO_306 (O_306,N_2984,N_2954);
nor UO_307 (O_307,N_2915,N_2960);
or UO_308 (O_308,N_2902,N_2926);
or UO_309 (O_309,N_2905,N_2945);
nor UO_310 (O_310,N_2953,N_2971);
nand UO_311 (O_311,N_2983,N_2963);
nand UO_312 (O_312,N_2933,N_2931);
or UO_313 (O_313,N_2995,N_2996);
or UO_314 (O_314,N_2986,N_2916);
nand UO_315 (O_315,N_2961,N_2981);
or UO_316 (O_316,N_2975,N_2915);
and UO_317 (O_317,N_2923,N_2956);
and UO_318 (O_318,N_2910,N_2980);
nand UO_319 (O_319,N_2935,N_2962);
nand UO_320 (O_320,N_2924,N_2925);
xnor UO_321 (O_321,N_2975,N_2992);
nor UO_322 (O_322,N_2997,N_2998);
or UO_323 (O_323,N_2960,N_2936);
nand UO_324 (O_324,N_2910,N_2966);
and UO_325 (O_325,N_2973,N_2977);
nor UO_326 (O_326,N_2950,N_2935);
nor UO_327 (O_327,N_2961,N_2942);
and UO_328 (O_328,N_2903,N_2938);
nor UO_329 (O_329,N_2945,N_2932);
nand UO_330 (O_330,N_2907,N_2953);
nand UO_331 (O_331,N_2947,N_2995);
and UO_332 (O_332,N_2901,N_2926);
nand UO_333 (O_333,N_2936,N_2903);
and UO_334 (O_334,N_2974,N_2923);
or UO_335 (O_335,N_2959,N_2918);
or UO_336 (O_336,N_2963,N_2952);
or UO_337 (O_337,N_2981,N_2942);
nand UO_338 (O_338,N_2960,N_2942);
nand UO_339 (O_339,N_2939,N_2930);
nand UO_340 (O_340,N_2978,N_2981);
nand UO_341 (O_341,N_2990,N_2914);
nand UO_342 (O_342,N_2907,N_2943);
nor UO_343 (O_343,N_2921,N_2986);
nor UO_344 (O_344,N_2938,N_2940);
and UO_345 (O_345,N_2946,N_2995);
and UO_346 (O_346,N_2925,N_2943);
nand UO_347 (O_347,N_2937,N_2911);
nand UO_348 (O_348,N_2972,N_2978);
nor UO_349 (O_349,N_2995,N_2987);
nand UO_350 (O_350,N_2976,N_2962);
nand UO_351 (O_351,N_2966,N_2923);
nor UO_352 (O_352,N_2950,N_2978);
nor UO_353 (O_353,N_2954,N_2931);
nand UO_354 (O_354,N_2941,N_2939);
or UO_355 (O_355,N_2916,N_2991);
or UO_356 (O_356,N_2901,N_2912);
and UO_357 (O_357,N_2948,N_2930);
nand UO_358 (O_358,N_2956,N_2969);
xnor UO_359 (O_359,N_2950,N_2923);
nor UO_360 (O_360,N_2902,N_2915);
nand UO_361 (O_361,N_2997,N_2984);
nand UO_362 (O_362,N_2990,N_2979);
or UO_363 (O_363,N_2967,N_2960);
nor UO_364 (O_364,N_2987,N_2970);
xor UO_365 (O_365,N_2975,N_2917);
nor UO_366 (O_366,N_2935,N_2902);
nor UO_367 (O_367,N_2907,N_2906);
and UO_368 (O_368,N_2961,N_2991);
nor UO_369 (O_369,N_2965,N_2934);
and UO_370 (O_370,N_2984,N_2985);
nor UO_371 (O_371,N_2992,N_2990);
nand UO_372 (O_372,N_2904,N_2992);
nor UO_373 (O_373,N_2964,N_2987);
and UO_374 (O_374,N_2962,N_2957);
nor UO_375 (O_375,N_2970,N_2934);
nor UO_376 (O_376,N_2936,N_2991);
or UO_377 (O_377,N_2954,N_2973);
xnor UO_378 (O_378,N_2962,N_2980);
or UO_379 (O_379,N_2937,N_2975);
nor UO_380 (O_380,N_2912,N_2985);
or UO_381 (O_381,N_2941,N_2984);
and UO_382 (O_382,N_2946,N_2916);
or UO_383 (O_383,N_2941,N_2949);
nand UO_384 (O_384,N_2955,N_2924);
nor UO_385 (O_385,N_2926,N_2973);
and UO_386 (O_386,N_2964,N_2994);
nand UO_387 (O_387,N_2921,N_2950);
or UO_388 (O_388,N_2991,N_2990);
or UO_389 (O_389,N_2980,N_2965);
nor UO_390 (O_390,N_2993,N_2906);
nor UO_391 (O_391,N_2981,N_2963);
nand UO_392 (O_392,N_2948,N_2974);
nor UO_393 (O_393,N_2977,N_2961);
nor UO_394 (O_394,N_2919,N_2947);
nand UO_395 (O_395,N_2963,N_2930);
nor UO_396 (O_396,N_2968,N_2935);
nand UO_397 (O_397,N_2974,N_2968);
and UO_398 (O_398,N_2978,N_2953);
nand UO_399 (O_399,N_2947,N_2915);
nand UO_400 (O_400,N_2996,N_2969);
nor UO_401 (O_401,N_2925,N_2933);
nand UO_402 (O_402,N_2936,N_2947);
or UO_403 (O_403,N_2986,N_2979);
nor UO_404 (O_404,N_2919,N_2986);
and UO_405 (O_405,N_2958,N_2982);
or UO_406 (O_406,N_2974,N_2997);
and UO_407 (O_407,N_2976,N_2981);
nor UO_408 (O_408,N_2954,N_2998);
and UO_409 (O_409,N_2905,N_2942);
or UO_410 (O_410,N_2900,N_2965);
and UO_411 (O_411,N_2934,N_2938);
or UO_412 (O_412,N_2992,N_2911);
and UO_413 (O_413,N_2902,N_2932);
and UO_414 (O_414,N_2971,N_2909);
nor UO_415 (O_415,N_2941,N_2989);
and UO_416 (O_416,N_2937,N_2959);
and UO_417 (O_417,N_2962,N_2954);
and UO_418 (O_418,N_2992,N_2956);
and UO_419 (O_419,N_2950,N_2952);
or UO_420 (O_420,N_2961,N_2907);
or UO_421 (O_421,N_2907,N_2964);
nand UO_422 (O_422,N_2922,N_2938);
nand UO_423 (O_423,N_2966,N_2916);
nor UO_424 (O_424,N_2912,N_2907);
nor UO_425 (O_425,N_2935,N_2986);
nand UO_426 (O_426,N_2994,N_2969);
or UO_427 (O_427,N_2991,N_2943);
nand UO_428 (O_428,N_2903,N_2994);
nand UO_429 (O_429,N_2953,N_2944);
or UO_430 (O_430,N_2901,N_2958);
and UO_431 (O_431,N_2978,N_2900);
nand UO_432 (O_432,N_2901,N_2981);
or UO_433 (O_433,N_2992,N_2922);
and UO_434 (O_434,N_2977,N_2981);
nor UO_435 (O_435,N_2916,N_2933);
nor UO_436 (O_436,N_2978,N_2903);
and UO_437 (O_437,N_2997,N_2968);
nor UO_438 (O_438,N_2943,N_2909);
nor UO_439 (O_439,N_2921,N_2915);
or UO_440 (O_440,N_2900,N_2915);
and UO_441 (O_441,N_2988,N_2954);
nand UO_442 (O_442,N_2947,N_2975);
and UO_443 (O_443,N_2954,N_2938);
nor UO_444 (O_444,N_2980,N_2973);
nor UO_445 (O_445,N_2999,N_2907);
and UO_446 (O_446,N_2909,N_2979);
and UO_447 (O_447,N_2972,N_2917);
xor UO_448 (O_448,N_2969,N_2955);
and UO_449 (O_449,N_2948,N_2986);
or UO_450 (O_450,N_2967,N_2956);
or UO_451 (O_451,N_2913,N_2976);
nand UO_452 (O_452,N_2994,N_2941);
or UO_453 (O_453,N_2960,N_2912);
or UO_454 (O_454,N_2962,N_2901);
or UO_455 (O_455,N_2993,N_2950);
or UO_456 (O_456,N_2964,N_2926);
nand UO_457 (O_457,N_2945,N_2980);
xnor UO_458 (O_458,N_2941,N_2921);
and UO_459 (O_459,N_2990,N_2952);
or UO_460 (O_460,N_2977,N_2911);
nand UO_461 (O_461,N_2907,N_2905);
or UO_462 (O_462,N_2929,N_2928);
and UO_463 (O_463,N_2954,N_2966);
nand UO_464 (O_464,N_2971,N_2945);
and UO_465 (O_465,N_2902,N_2992);
nand UO_466 (O_466,N_2990,N_2968);
nand UO_467 (O_467,N_2993,N_2978);
or UO_468 (O_468,N_2994,N_2935);
nand UO_469 (O_469,N_2990,N_2935);
nand UO_470 (O_470,N_2970,N_2942);
and UO_471 (O_471,N_2965,N_2983);
or UO_472 (O_472,N_2901,N_2922);
nand UO_473 (O_473,N_2992,N_2969);
and UO_474 (O_474,N_2905,N_2977);
nand UO_475 (O_475,N_2901,N_2907);
nor UO_476 (O_476,N_2963,N_2964);
nand UO_477 (O_477,N_2911,N_2922);
nor UO_478 (O_478,N_2980,N_2936);
and UO_479 (O_479,N_2939,N_2949);
nor UO_480 (O_480,N_2920,N_2921);
or UO_481 (O_481,N_2969,N_2922);
and UO_482 (O_482,N_2974,N_2995);
nand UO_483 (O_483,N_2980,N_2955);
nand UO_484 (O_484,N_2920,N_2905);
nor UO_485 (O_485,N_2948,N_2965);
or UO_486 (O_486,N_2924,N_2984);
nor UO_487 (O_487,N_2950,N_2946);
or UO_488 (O_488,N_2949,N_2986);
nor UO_489 (O_489,N_2996,N_2985);
nand UO_490 (O_490,N_2909,N_2923);
or UO_491 (O_491,N_2993,N_2901);
or UO_492 (O_492,N_2909,N_2914);
nand UO_493 (O_493,N_2979,N_2920);
or UO_494 (O_494,N_2994,N_2927);
or UO_495 (O_495,N_2995,N_2956);
and UO_496 (O_496,N_2905,N_2999);
or UO_497 (O_497,N_2918,N_2948);
or UO_498 (O_498,N_2943,N_2901);
nor UO_499 (O_499,N_2977,N_2946);
endmodule