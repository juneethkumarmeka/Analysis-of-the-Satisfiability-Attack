module basic_750_5000_1000_2_levels_1xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2501,N_2502,N_2507,N_2509,N_2510,N_2511,N_2512,N_2513,N_2515,N_2516,N_2517,N_2518,N_2521,N_2522,N_2524,N_2525,N_2526,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2540,N_2541,N_2542,N_2543,N_2545,N_2546,N_2547,N_2548,N_2549,N_2551,N_2552,N_2553,N_2554,N_2555,N_2557,N_2558,N_2559,N_2560,N_2561,N_2563,N_2565,N_2567,N_2568,N_2569,N_2570,N_2573,N_2574,N_2575,N_2576,N_2577,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2615,N_2617,N_2618,N_2620,N_2621,N_2622,N_2624,N_2625,N_2627,N_2628,N_2629,N_2631,N_2632,N_2634,N_2636,N_2637,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2655,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2670,N_2673,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2692,N_2694,N_2695,N_2696,N_2697,N_2698,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2782,N_2784,N_2785,N_2786,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2820,N_2822,N_2824,N_2825,N_2827,N_2828,N_2829,N_2830,N_2832,N_2833,N_2834,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2852,N_2853,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2867,N_2868,N_2869,N_2870,N_2872,N_2874,N_2876,N_2877,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2899,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2910,N_2911,N_2912,N_2914,N_2915,N_2916,N_2917,N_2919,N_2920,N_2921,N_2922,N_2923,N_2925,N_2926,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2936,N_2937,N_2938,N_2939,N_2940,N_2942,N_2943,N_2944,N_2946,N_2948,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2964,N_2966,N_2968,N_2969,N_2970,N_2971,N_2972,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2982,N_2983,N_2986,N_2988,N_2990,N_2991,N_2992,N_2993,N_2994,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3022,N_3023,N_3024,N_3025,N_3026,N_3028,N_3029,N_3030,N_3031,N_3032,N_3034,N_3035,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3044,N_3045,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3075,N_3076,N_3077,N_3078,N_3080,N_3081,N_3082,N_3083,N_3084,N_3086,N_3087,N_3088,N_3089,N_3091,N_3092,N_3093,N_3095,N_3096,N_3097,N_3098,N_3099,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3113,N_3114,N_3115,N_3116,N_3117,N_3119,N_3125,N_3127,N_3128,N_3129,N_3130,N_3132,N_3133,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3144,N_3145,N_3147,N_3148,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3159,N_3160,N_3162,N_3164,N_3165,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3184,N_3185,N_3186,N_3188,N_3189,N_3191,N_3192,N_3193,N_3194,N_3195,N_3197,N_3198,N_3199,N_3201,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3235,N_3236,N_3237,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3274,N_3276,N_3277,N_3278,N_3279,N_3280,N_3282,N_3284,N_3287,N_3288,N_3290,N_3292,N_3293,N_3294,N_3295,N_3297,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3309,N_3310,N_3311,N_3312,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3350,N_3351,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3391,N_3392,N_3393,N_3394,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3410,N_3411,N_3412,N_3413,N_3415,N_3416,N_3417,N_3418,N_3420,N_3422,N_3423,N_3424,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3438,N_3439,N_3440,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3450,N_3451,N_3453,N_3454,N_3455,N_3457,N_3458,N_3459,N_3460,N_3462,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3477,N_3479,N_3480,N_3481,N_3482,N_3483,N_3485,N_3486,N_3487,N_3488,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3504,N_3505,N_3506,N_3508,N_3509,N_3510,N_3511,N_3512,N_3514,N_3517,N_3518,N_3520,N_3522,N_3523,N_3525,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3548,N_3550,N_3551,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3577,N_3578,N_3579,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3592,N_3593,N_3594,N_3595,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3607,N_3608,N_3609,N_3611,N_3614,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3628,N_3629,N_3630,N_3631,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3653,N_3654,N_3655,N_3656,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3680,N_3681,N_3683,N_3685,N_3686,N_3687,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3721,N_3724,N_3725,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3737,N_3739,N_3740,N_3743,N_3744,N_3746,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3763,N_3764,N_3765,N_3768,N_3769,N_3770,N_3771,N_3772,N_3774,N_3776,N_3777,N_3778,N_3779,N_3780,N_3782,N_3783,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3792,N_3793,N_3796,N_3797,N_3798,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3810,N_3812,N_3813,N_3814,N_3817,N_3818,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3829,N_3830,N_3831,N_3832,N_3833,N_3836,N_3838,N_3839,N_3840,N_3841,N_3843,N_3844,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3859,N_3860,N_3861,N_3862,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3885,N_3886,N_3888,N_3889,N_3890,N_3891,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3900,N_3901,N_3902,N_3903,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3925,N_3926,N_3927,N_3928,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3942,N_3943,N_3945,N_3946,N_3947,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3961,N_3962,N_3965,N_3967,N_3968,N_3969,N_3970,N_3972,N_3973,N_3974,N_3976,N_3977,N_3979,N_3980,N_3981,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3997,N_3998,N_4000,N_4003,N_4004,N_4005,N_4007,N_4008,N_4010,N_4011,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4023,N_4024,N_4025,N_4026,N_4028,N_4030,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4058,N_4059,N_4060,N_4061,N_4062,N_4065,N_4066,N_4067,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4087,N_4088,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4129,N_4131,N_4133,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4148,N_4149,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4161,N_4162,N_4163,N_4164,N_4166,N_4167,N_4170,N_4171,N_4173,N_4174,N_4175,N_4177,N_4180,N_4181,N_4183,N_4184,N_4187,N_4188,N_4189,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4208,N_4209,N_4210,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4255,N_4256,N_4257,N_4259,N_4260,N_4261,N_4263,N_4265,N_4266,N_4268,N_4270,N_4271,N_4273,N_4276,N_4277,N_4278,N_4280,N_4281,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4303,N_4305,N_4306,N_4307,N_4308,N_4309,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4318,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4345,N_4346,N_4347,N_4348,N_4350,N_4351,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4360,N_4361,N_4362,N_4363,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4375,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4396,N_4398,N_4399,N_4400,N_4401,N_4402,N_4404,N_4405,N_4406,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4425,N_4426,N_4427,N_4428,N_4429,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4441,N_4442,N_4443,N_4444,N_4445,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4455,N_4457,N_4458,N_4463,N_4464,N_4466,N_4467,N_4468,N_4469,N_4472,N_4473,N_4474,N_4475,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4490,N_4491,N_4492,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4509,N_4510,N_4511,N_4512,N_4514,N_4515,N_4516,N_4517,N_4518,N_4521,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4572,N_4573,N_4574,N_4575,N_4576,N_4579,N_4580,N_4583,N_4584,N_4585,N_4586,N_4588,N_4589,N_4590,N_4592,N_4593,N_4594,N_4595,N_4598,N_4599,N_4600,N_4601,N_4602,N_4604,N_4605,N_4606,N_4607,N_4608,N_4610,N_4611,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4641,N_4643,N_4644,N_4645,N_4646,N_4648,N_4649,N_4650,N_4651,N_4652,N_4654,N_4656,N_4657,N_4658,N_4660,N_4661,N_4663,N_4664,N_4666,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4676,N_4677,N_4678,N_4679,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4701,N_4703,N_4704,N_4705,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4719,N_4721,N_4722,N_4723,N_4724,N_4725,N_4727,N_4728,N_4729,N_4730,N_4732,N_4733,N_4734,N_4736,N_4737,N_4738,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4752,N_4754,N_4755,N_4757,N_4759,N_4761,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4783,N_4784,N_4787,N_4788,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4822,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4834,N_4835,N_4836,N_4838,N_4840,N_4842,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4856,N_4859,N_4860,N_4861,N_4863,N_4864,N_4866,N_4867,N_4869,N_4870,N_4872,N_4873,N_4874,N_4875,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4907,N_4908,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4918,N_4919,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4933,N_4935,N_4936,N_4937,N_4938,N_4940,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4993,N_4994,N_4996,N_4997,N_4998,N_4999;
or U0 (N_0,In_220,In_195);
or U1 (N_1,In_495,In_62);
or U2 (N_2,In_446,In_688);
or U3 (N_3,In_118,In_645);
nor U4 (N_4,In_655,In_735);
or U5 (N_5,In_368,In_472);
nor U6 (N_6,In_620,In_516);
or U7 (N_7,In_573,In_320);
nand U8 (N_8,In_25,In_461);
nand U9 (N_9,In_672,In_494);
nor U10 (N_10,In_304,In_242);
nor U11 (N_11,In_355,In_568);
and U12 (N_12,In_718,In_422);
and U13 (N_13,In_239,In_389);
nor U14 (N_14,In_679,In_59);
or U15 (N_15,In_405,In_84);
and U16 (N_16,In_361,In_262);
or U17 (N_17,In_120,In_581);
or U18 (N_18,In_580,In_247);
or U19 (N_19,In_159,In_678);
or U20 (N_20,In_636,In_417);
nor U21 (N_21,In_456,In_458);
xnor U22 (N_22,In_504,In_332);
nand U23 (N_23,In_130,In_505);
nor U24 (N_24,In_670,In_272);
and U25 (N_25,In_275,In_696);
nor U26 (N_26,In_148,In_280);
nand U27 (N_27,In_96,In_309);
nand U28 (N_28,In_101,In_509);
and U29 (N_29,In_337,In_265);
nor U30 (N_30,In_499,In_685);
nand U31 (N_31,In_734,In_575);
nor U32 (N_32,In_481,In_419);
or U33 (N_33,In_281,In_73);
and U34 (N_34,In_233,In_119);
nand U35 (N_35,In_199,In_576);
and U36 (N_36,In_661,In_204);
nor U37 (N_37,In_168,In_567);
and U38 (N_38,In_630,In_677);
nand U39 (N_39,In_742,In_595);
nand U40 (N_40,In_531,In_364);
nand U41 (N_41,In_705,In_79);
nor U42 (N_42,In_122,In_253);
nand U43 (N_43,In_135,In_534);
nor U44 (N_44,In_442,In_229);
and U45 (N_45,In_26,In_517);
or U46 (N_46,In_428,In_268);
nor U47 (N_47,In_542,In_522);
nor U48 (N_48,In_338,In_411);
and U49 (N_49,In_3,In_91);
nand U50 (N_50,In_453,In_160);
or U51 (N_51,In_746,In_290);
nand U52 (N_52,In_185,In_241);
and U53 (N_53,In_19,In_56);
nor U54 (N_54,In_165,In_455);
or U55 (N_55,In_487,In_612);
and U56 (N_56,In_631,In_106);
and U57 (N_57,In_139,In_403);
or U58 (N_58,In_98,In_225);
nor U59 (N_59,In_182,In_342);
or U60 (N_60,In_484,In_408);
or U61 (N_61,In_215,In_552);
nor U62 (N_62,In_97,In_550);
or U63 (N_63,In_180,In_614);
xor U64 (N_64,In_64,In_643);
nand U65 (N_65,In_189,In_291);
and U66 (N_66,In_113,In_109);
nand U67 (N_67,In_114,In_434);
nand U68 (N_68,In_223,In_142);
or U69 (N_69,In_704,In_549);
nor U70 (N_70,In_156,In_8);
xor U71 (N_71,In_424,In_398);
and U72 (N_72,In_302,In_43);
nor U73 (N_73,In_232,In_33);
or U74 (N_74,In_99,In_406);
nand U75 (N_75,In_506,In_384);
nand U76 (N_76,In_492,In_731);
nand U77 (N_77,In_635,In_6);
or U78 (N_78,In_149,In_154);
and U79 (N_79,In_22,In_42);
and U80 (N_80,In_543,In_21);
or U81 (N_81,In_333,In_465);
nor U82 (N_82,In_521,In_31);
and U83 (N_83,In_212,In_387);
or U84 (N_84,In_664,In_489);
or U85 (N_85,In_603,In_48);
and U86 (N_86,In_681,In_571);
or U87 (N_87,In_736,In_277);
nand U88 (N_88,In_605,In_482);
nor U89 (N_89,In_133,In_538);
nor U90 (N_90,In_607,In_452);
and U91 (N_91,In_315,In_564);
and U92 (N_92,In_536,In_283);
nand U93 (N_93,In_723,In_151);
and U94 (N_94,In_222,In_602);
nor U95 (N_95,In_341,In_9);
nand U96 (N_96,In_47,In_488);
and U97 (N_97,In_193,In_732);
nor U98 (N_98,In_418,In_323);
nand U99 (N_99,In_625,In_11);
nor U100 (N_100,In_658,In_54);
nor U101 (N_101,In_574,In_646);
nor U102 (N_102,In_739,In_624);
and U103 (N_103,In_695,In_29);
xor U104 (N_104,In_445,In_640);
nand U105 (N_105,In_279,In_432);
nand U106 (N_106,In_708,In_713);
nand U107 (N_107,In_250,In_533);
or U108 (N_108,In_390,In_157);
or U109 (N_109,In_294,In_256);
nand U110 (N_110,In_125,In_164);
nor U111 (N_111,In_553,In_15);
nor U112 (N_112,In_409,In_621);
nand U113 (N_113,In_414,In_116);
nand U114 (N_114,In_490,In_558);
nand U115 (N_115,In_184,In_244);
and U116 (N_116,In_377,In_298);
nor U117 (N_117,In_90,In_747);
and U118 (N_118,In_447,In_429);
or U119 (N_119,In_383,In_236);
nor U120 (N_120,In_629,In_599);
or U121 (N_121,In_200,In_136);
nand U122 (N_122,In_86,In_107);
nor U123 (N_123,In_243,In_28);
nand U124 (N_124,In_311,In_444);
or U125 (N_125,In_124,In_528);
and U126 (N_126,In_588,In_210);
or U127 (N_127,In_176,In_617);
or U128 (N_128,In_61,In_394);
and U129 (N_129,In_637,In_660);
or U130 (N_130,In_402,In_146);
or U131 (N_131,In_95,In_515);
nor U132 (N_132,In_716,In_360);
and U133 (N_133,In_194,In_134);
and U134 (N_134,In_70,In_308);
or U135 (N_135,In_448,In_724);
nand U136 (N_136,In_652,In_17);
or U137 (N_137,In_108,In_684);
nor U138 (N_138,In_667,In_305);
nor U139 (N_139,In_740,In_545);
or U140 (N_140,In_464,In_58);
or U141 (N_141,In_657,In_715);
nor U142 (N_142,In_435,In_717);
and U143 (N_143,In_354,In_166);
nand U144 (N_144,In_642,In_327);
and U145 (N_145,In_16,In_299);
and U146 (N_146,In_57,In_51);
nor U147 (N_147,In_325,In_619);
nand U148 (N_148,In_85,In_501);
nand U149 (N_149,In_334,In_479);
and U150 (N_150,In_219,In_745);
nor U151 (N_151,In_20,In_317);
or U152 (N_152,In_510,In_45);
and U153 (N_153,In_474,In_246);
nand U154 (N_154,In_153,In_507);
nor U155 (N_155,In_560,In_513);
and U156 (N_156,In_727,In_82);
or U157 (N_157,In_140,In_608);
nor U158 (N_158,In_141,In_30);
nor U159 (N_159,In_729,In_412);
nor U160 (N_160,In_248,In_80);
nor U161 (N_161,In_350,In_654);
and U162 (N_162,In_663,In_44);
nand U163 (N_163,In_421,In_511);
nand U164 (N_164,In_473,In_584);
and U165 (N_165,In_703,In_36);
nor U166 (N_166,In_459,In_152);
or U167 (N_167,In_137,In_451);
or U168 (N_168,In_230,In_207);
nor U169 (N_169,In_145,In_376);
nor U170 (N_170,In_121,In_351);
and U171 (N_171,In_470,In_183);
nor U172 (N_172,In_129,In_525);
nand U173 (N_173,In_535,In_301);
nor U174 (N_174,In_362,In_514);
and U175 (N_175,In_710,In_601);
nand U176 (N_176,In_375,In_240);
nor U177 (N_177,In_478,In_425);
nor U178 (N_178,In_622,In_413);
or U179 (N_179,In_616,In_187);
nor U180 (N_180,In_726,In_190);
nor U181 (N_181,In_65,In_117);
nor U182 (N_182,In_345,In_530);
and U183 (N_183,In_391,In_300);
nand U184 (N_184,In_237,In_615);
nand U185 (N_185,In_379,In_673);
or U186 (N_186,In_730,In_55);
or U187 (N_187,In_569,In_683);
nor U188 (N_188,In_328,In_198);
or U189 (N_189,In_523,In_208);
and U190 (N_190,In_466,In_597);
nand U191 (N_191,In_344,In_486);
nor U192 (N_192,In_177,In_496);
and U193 (N_193,In_380,In_527);
nand U194 (N_194,In_356,In_261);
nor U195 (N_195,In_537,In_372);
or U196 (N_196,In_467,In_722);
nor U197 (N_197,In_306,In_254);
nand U198 (N_198,In_609,In_500);
nand U199 (N_199,In_647,In_4);
or U200 (N_200,In_547,In_469);
nand U201 (N_201,In_659,In_638);
nor U202 (N_202,In_450,In_206);
nor U203 (N_203,In_5,In_278);
or U204 (N_204,In_143,In_102);
or U205 (N_205,In_287,In_626);
nand U206 (N_206,In_353,In_382);
or U207 (N_207,In_395,In_540);
nor U208 (N_208,In_14,In_503);
and U209 (N_209,In_357,In_214);
nand U210 (N_210,In_594,In_709);
nand U211 (N_211,In_628,In_266);
nand U212 (N_212,In_743,In_669);
or U213 (N_213,In_675,In_393);
nor U214 (N_214,In_544,In_52);
nand U215 (N_215,In_426,In_63);
and U216 (N_216,In_593,In_158);
nor U217 (N_217,In_163,In_430);
nor U218 (N_218,In_346,In_582);
nor U219 (N_219,In_252,In_221);
and U220 (N_220,In_416,In_369);
nor U221 (N_221,In_680,In_512);
and U222 (N_222,In_712,In_738);
and U223 (N_223,In_518,In_115);
or U224 (N_224,In_559,In_570);
nand U225 (N_225,In_373,In_555);
or U226 (N_226,In_94,In_284);
or U227 (N_227,In_330,In_358);
or U228 (N_228,In_653,In_319);
and U229 (N_229,In_363,In_589);
and U230 (N_230,In_267,In_460);
nand U231 (N_231,In_554,In_491);
nand U232 (N_232,In_24,In_697);
or U233 (N_233,In_707,In_572);
nor U234 (N_234,In_485,In_437);
nor U235 (N_235,In_181,In_126);
and U236 (N_236,In_60,In_420);
nand U237 (N_237,In_50,In_441);
and U238 (N_238,In_269,In_132);
nor U239 (N_239,In_35,In_71);
nor U240 (N_240,In_359,In_583);
and U241 (N_241,In_577,In_228);
and U242 (N_242,In_270,In_226);
nand U243 (N_243,In_668,In_175);
or U244 (N_244,In_604,In_191);
nand U245 (N_245,In_67,In_596);
nand U246 (N_246,In_127,In_725);
and U247 (N_247,In_144,In_179);
or U248 (N_248,In_415,In_75);
nand U249 (N_249,In_37,In_557);
nand U250 (N_250,In_310,In_463);
nand U251 (N_251,In_378,In_285);
and U252 (N_252,In_519,In_561);
nand U253 (N_253,In_255,In_88);
nor U254 (N_254,In_314,In_706);
nand U255 (N_255,In_7,In_392);
or U256 (N_256,In_468,In_296);
or U257 (N_257,In_340,In_186);
and U258 (N_258,In_161,In_273);
or U259 (N_259,In_123,In_105);
nor U260 (N_260,In_634,In_641);
and U261 (N_261,In_566,In_662);
and U262 (N_262,In_699,In_686);
or U263 (N_263,In_648,In_565);
or U264 (N_264,In_656,In_39);
nor U265 (N_265,In_258,In_639);
nor U266 (N_266,In_714,In_245);
nor U267 (N_267,In_307,In_150);
and U268 (N_268,In_76,In_100);
nor U269 (N_269,In_623,In_613);
and U270 (N_270,In_335,In_196);
nor U271 (N_271,In_173,In_322);
or U272 (N_272,In_744,In_440);
and U273 (N_273,In_532,In_627);
nand U274 (N_274,In_676,In_192);
or U275 (N_275,In_556,In_457);
nand U276 (N_276,In_234,In_665);
or U277 (N_277,In_78,In_77);
or U278 (N_278,In_366,In_477);
and U279 (N_279,In_702,In_349);
nand U280 (N_280,In_397,In_502);
nand U281 (N_281,In_651,In_400);
and U282 (N_282,In_721,In_49);
and U283 (N_283,In_27,In_689);
or U284 (N_284,In_271,In_203);
nand U285 (N_285,In_374,In_381);
or U286 (N_286,In_282,In_40);
nand U287 (N_287,In_227,In_288);
and U288 (N_288,In_748,In_548);
nand U289 (N_289,In_449,In_737);
xnor U290 (N_290,In_520,In_498);
nor U291 (N_291,In_316,In_471);
or U292 (N_292,In_10,In_541);
or U293 (N_293,In_687,In_224);
nor U294 (N_294,In_401,In_443);
nor U295 (N_295,In_693,In_66);
and U296 (N_296,In_286,In_274);
nor U297 (N_297,In_303,In_352);
nor U298 (N_298,In_103,In_719);
or U299 (N_299,In_590,In_201);
or U300 (N_300,In_147,In_347);
nor U301 (N_301,In_694,In_649);
or U302 (N_302,In_329,In_2);
nand U303 (N_303,In_563,In_217);
nor U304 (N_304,In_41,In_483);
nand U305 (N_305,In_546,In_318);
and U306 (N_306,In_92,In_436);
nor U307 (N_307,In_343,In_438);
or U308 (N_308,In_167,In_529);
nor U309 (N_309,In_698,In_480);
nand U310 (N_310,In_87,In_728);
nor U311 (N_311,In_749,In_578);
nor U312 (N_312,In_386,In_68);
or U313 (N_313,In_202,In_231);
or U314 (N_314,In_293,In_586);
or U315 (N_315,In_598,In_399);
or U316 (N_316,In_292,In_89);
nand U317 (N_317,In_439,In_493);
nor U318 (N_318,In_348,In_111);
nor U319 (N_319,In_23,In_587);
nand U320 (N_320,In_331,In_295);
and U321 (N_321,In_433,In_38);
nor U322 (N_322,In_410,In_666);
or U323 (N_323,In_611,In_12);
nand U324 (N_324,In_213,In_72);
nor U325 (N_325,In_74,In_610);
and U326 (N_326,In_682,In_526);
xnor U327 (N_327,In_188,In_591);
or U328 (N_328,In_249,In_579);
or U329 (N_329,In_524,In_83);
nor U330 (N_330,In_312,In_497);
nand U331 (N_331,In_427,In_289);
nand U332 (N_332,In_128,In_632);
nor U333 (N_333,In_155,In_34);
nor U334 (N_334,In_131,In_385);
and U335 (N_335,In_592,In_110);
and U336 (N_336,In_197,In_0);
nand U337 (N_337,In_321,In_326);
or U338 (N_338,In_454,In_169);
nand U339 (N_339,In_171,In_260);
or U340 (N_340,In_733,In_585);
and U341 (N_341,In_690,In_69);
nor U342 (N_342,In_431,In_257);
or U343 (N_343,In_606,In_701);
and U344 (N_344,In_93,In_13);
or U345 (N_345,In_562,In_462);
nand U346 (N_346,In_170,In_423);
nor U347 (N_347,In_371,In_81);
nand U348 (N_348,In_367,In_370);
nor U349 (N_349,In_264,In_138);
nand U350 (N_350,In_174,In_276);
or U351 (N_351,In_600,In_388);
and U352 (N_352,In_1,In_238);
nand U353 (N_353,In_53,In_700);
nor U354 (N_354,In_46,In_551);
or U355 (N_355,In_32,In_205);
nand U356 (N_356,In_396,In_178);
nor U357 (N_357,In_218,In_324);
and U358 (N_358,In_720,In_235);
nor U359 (N_359,In_211,In_209);
nand U360 (N_360,In_475,In_404);
nand U361 (N_361,In_741,In_671);
or U362 (N_362,In_644,In_259);
nor U363 (N_363,In_297,In_339);
or U364 (N_364,In_112,In_674);
and U365 (N_365,In_365,In_216);
and U366 (N_366,In_172,In_251);
nor U367 (N_367,In_407,In_711);
and U368 (N_368,In_476,In_633);
nor U369 (N_369,In_539,In_18);
nand U370 (N_370,In_104,In_650);
nor U371 (N_371,In_313,In_618);
or U372 (N_372,In_508,In_336);
nor U373 (N_373,In_691,In_263);
or U374 (N_374,In_692,In_162);
and U375 (N_375,In_27,In_208);
nor U376 (N_376,In_337,In_683);
and U377 (N_377,In_694,In_27);
nand U378 (N_378,In_698,In_557);
nor U379 (N_379,In_748,In_158);
or U380 (N_380,In_324,In_416);
or U381 (N_381,In_600,In_456);
nand U382 (N_382,In_318,In_75);
nand U383 (N_383,In_583,In_300);
or U384 (N_384,In_666,In_644);
or U385 (N_385,In_175,In_64);
nand U386 (N_386,In_254,In_284);
nand U387 (N_387,In_191,In_321);
or U388 (N_388,In_318,In_746);
nor U389 (N_389,In_498,In_630);
nand U390 (N_390,In_435,In_103);
nand U391 (N_391,In_611,In_312);
and U392 (N_392,In_227,In_214);
nand U393 (N_393,In_7,In_628);
and U394 (N_394,In_552,In_369);
nor U395 (N_395,In_457,In_487);
nor U396 (N_396,In_33,In_744);
or U397 (N_397,In_119,In_296);
xor U398 (N_398,In_23,In_742);
nor U399 (N_399,In_271,In_702);
or U400 (N_400,In_122,In_339);
nand U401 (N_401,In_199,In_651);
nand U402 (N_402,In_637,In_327);
or U403 (N_403,In_285,In_27);
nor U404 (N_404,In_700,In_69);
or U405 (N_405,In_676,In_738);
or U406 (N_406,In_560,In_484);
nand U407 (N_407,In_354,In_44);
nand U408 (N_408,In_745,In_541);
or U409 (N_409,In_675,In_481);
nor U410 (N_410,In_625,In_298);
nand U411 (N_411,In_227,In_675);
nand U412 (N_412,In_452,In_508);
nand U413 (N_413,In_482,In_224);
nor U414 (N_414,In_406,In_399);
nor U415 (N_415,In_12,In_532);
nor U416 (N_416,In_215,In_514);
nor U417 (N_417,In_549,In_271);
or U418 (N_418,In_360,In_646);
nor U419 (N_419,In_101,In_575);
and U420 (N_420,In_171,In_553);
and U421 (N_421,In_549,In_722);
and U422 (N_422,In_70,In_553);
nor U423 (N_423,In_408,In_334);
and U424 (N_424,In_283,In_230);
nor U425 (N_425,In_141,In_739);
nand U426 (N_426,In_103,In_175);
or U427 (N_427,In_286,In_638);
or U428 (N_428,In_364,In_460);
nand U429 (N_429,In_421,In_371);
nor U430 (N_430,In_82,In_480);
nand U431 (N_431,In_582,In_29);
and U432 (N_432,In_334,In_424);
or U433 (N_433,In_390,In_234);
and U434 (N_434,In_691,In_185);
nor U435 (N_435,In_172,In_335);
nor U436 (N_436,In_409,In_471);
nand U437 (N_437,In_242,In_33);
and U438 (N_438,In_489,In_666);
or U439 (N_439,In_188,In_25);
nor U440 (N_440,In_140,In_423);
and U441 (N_441,In_703,In_421);
nor U442 (N_442,In_152,In_566);
or U443 (N_443,In_321,In_552);
and U444 (N_444,In_671,In_519);
or U445 (N_445,In_665,In_252);
or U446 (N_446,In_564,In_478);
or U447 (N_447,In_35,In_580);
and U448 (N_448,In_424,In_623);
nor U449 (N_449,In_726,In_171);
nand U450 (N_450,In_143,In_148);
nand U451 (N_451,In_120,In_179);
and U452 (N_452,In_419,In_581);
nand U453 (N_453,In_632,In_539);
nor U454 (N_454,In_246,In_442);
or U455 (N_455,In_285,In_65);
and U456 (N_456,In_383,In_714);
or U457 (N_457,In_367,In_577);
or U458 (N_458,In_176,In_92);
or U459 (N_459,In_212,In_567);
and U460 (N_460,In_229,In_366);
or U461 (N_461,In_250,In_107);
nand U462 (N_462,In_140,In_644);
or U463 (N_463,In_237,In_108);
nand U464 (N_464,In_474,In_238);
nor U465 (N_465,In_511,In_656);
and U466 (N_466,In_129,In_473);
nand U467 (N_467,In_254,In_503);
or U468 (N_468,In_734,In_145);
nand U469 (N_469,In_417,In_61);
nand U470 (N_470,In_272,In_164);
nand U471 (N_471,In_690,In_110);
or U472 (N_472,In_435,In_689);
and U473 (N_473,In_654,In_44);
or U474 (N_474,In_653,In_195);
nand U475 (N_475,In_716,In_452);
nand U476 (N_476,In_162,In_347);
nor U477 (N_477,In_101,In_201);
nor U478 (N_478,In_194,In_273);
or U479 (N_479,In_395,In_628);
and U480 (N_480,In_519,In_473);
or U481 (N_481,In_523,In_312);
nand U482 (N_482,In_381,In_276);
nand U483 (N_483,In_284,In_541);
or U484 (N_484,In_199,In_139);
nand U485 (N_485,In_277,In_92);
and U486 (N_486,In_636,In_529);
nand U487 (N_487,In_317,In_12);
xor U488 (N_488,In_55,In_707);
nand U489 (N_489,In_33,In_730);
nor U490 (N_490,In_677,In_609);
and U491 (N_491,In_675,In_272);
nor U492 (N_492,In_735,In_525);
xor U493 (N_493,In_169,In_521);
nand U494 (N_494,In_611,In_695);
nor U495 (N_495,In_361,In_142);
or U496 (N_496,In_152,In_131);
nor U497 (N_497,In_646,In_81);
and U498 (N_498,In_401,In_289);
and U499 (N_499,In_716,In_381);
and U500 (N_500,In_41,In_528);
nand U501 (N_501,In_294,In_721);
nor U502 (N_502,In_245,In_715);
nor U503 (N_503,In_657,In_194);
and U504 (N_504,In_309,In_362);
and U505 (N_505,In_354,In_21);
nand U506 (N_506,In_318,In_98);
or U507 (N_507,In_455,In_273);
and U508 (N_508,In_76,In_582);
nand U509 (N_509,In_424,In_721);
and U510 (N_510,In_261,In_249);
nand U511 (N_511,In_306,In_674);
nand U512 (N_512,In_378,In_146);
and U513 (N_513,In_258,In_665);
nand U514 (N_514,In_13,In_48);
nand U515 (N_515,In_144,In_568);
or U516 (N_516,In_673,In_190);
and U517 (N_517,In_517,In_178);
and U518 (N_518,In_600,In_538);
and U519 (N_519,In_160,In_364);
or U520 (N_520,In_116,In_680);
nand U521 (N_521,In_66,In_92);
and U522 (N_522,In_206,In_251);
and U523 (N_523,In_199,In_345);
and U524 (N_524,In_88,In_460);
and U525 (N_525,In_470,In_258);
nor U526 (N_526,In_144,In_265);
and U527 (N_527,In_716,In_408);
nand U528 (N_528,In_186,In_616);
or U529 (N_529,In_278,In_442);
nor U530 (N_530,In_126,In_271);
nor U531 (N_531,In_203,In_302);
nand U532 (N_532,In_212,In_22);
or U533 (N_533,In_483,In_515);
nand U534 (N_534,In_158,In_675);
nor U535 (N_535,In_167,In_663);
nand U536 (N_536,In_303,In_86);
or U537 (N_537,In_36,In_598);
or U538 (N_538,In_328,In_732);
and U539 (N_539,In_9,In_218);
nand U540 (N_540,In_174,In_529);
nor U541 (N_541,In_307,In_152);
nand U542 (N_542,In_673,In_22);
nand U543 (N_543,In_600,In_589);
or U544 (N_544,In_239,In_18);
nand U545 (N_545,In_537,In_587);
nor U546 (N_546,In_553,In_414);
nand U547 (N_547,In_194,In_685);
nor U548 (N_548,In_574,In_221);
nor U549 (N_549,In_682,In_418);
nor U550 (N_550,In_467,In_626);
or U551 (N_551,In_449,In_182);
nand U552 (N_552,In_305,In_664);
nor U553 (N_553,In_723,In_663);
and U554 (N_554,In_183,In_492);
or U555 (N_555,In_614,In_485);
nand U556 (N_556,In_636,In_215);
or U557 (N_557,In_68,In_539);
and U558 (N_558,In_318,In_386);
or U559 (N_559,In_571,In_516);
or U560 (N_560,In_649,In_512);
or U561 (N_561,In_337,In_6);
or U562 (N_562,In_745,In_299);
and U563 (N_563,In_603,In_568);
and U564 (N_564,In_287,In_49);
and U565 (N_565,In_571,In_680);
or U566 (N_566,In_304,In_154);
or U567 (N_567,In_679,In_306);
nor U568 (N_568,In_84,In_559);
nor U569 (N_569,In_184,In_103);
or U570 (N_570,In_8,In_439);
and U571 (N_571,In_211,In_350);
or U572 (N_572,In_195,In_184);
and U573 (N_573,In_461,In_702);
and U574 (N_574,In_656,In_336);
nand U575 (N_575,In_580,In_515);
and U576 (N_576,In_576,In_200);
and U577 (N_577,In_508,In_11);
nand U578 (N_578,In_439,In_365);
and U579 (N_579,In_574,In_51);
nor U580 (N_580,In_589,In_583);
nor U581 (N_581,In_602,In_547);
nor U582 (N_582,In_542,In_129);
and U583 (N_583,In_344,In_504);
or U584 (N_584,In_311,In_374);
or U585 (N_585,In_721,In_22);
or U586 (N_586,In_9,In_412);
nand U587 (N_587,In_614,In_293);
nand U588 (N_588,In_749,In_53);
nand U589 (N_589,In_515,In_664);
nand U590 (N_590,In_717,In_180);
nor U591 (N_591,In_333,In_50);
nand U592 (N_592,In_531,In_297);
and U593 (N_593,In_404,In_591);
and U594 (N_594,In_445,In_141);
nand U595 (N_595,In_60,In_4);
nand U596 (N_596,In_697,In_198);
or U597 (N_597,In_665,In_94);
nand U598 (N_598,In_80,In_544);
nand U599 (N_599,In_186,In_562);
nand U600 (N_600,In_172,In_424);
nor U601 (N_601,In_524,In_477);
nor U602 (N_602,In_252,In_514);
and U603 (N_603,In_405,In_1);
and U604 (N_604,In_396,In_181);
and U605 (N_605,In_297,In_384);
or U606 (N_606,In_195,In_123);
nand U607 (N_607,In_438,In_371);
nor U608 (N_608,In_307,In_585);
and U609 (N_609,In_56,In_670);
nand U610 (N_610,In_314,In_365);
nor U611 (N_611,In_392,In_43);
nand U612 (N_612,In_247,In_38);
and U613 (N_613,In_481,In_361);
and U614 (N_614,In_256,In_13);
nand U615 (N_615,In_576,In_112);
nor U616 (N_616,In_660,In_351);
or U617 (N_617,In_450,In_367);
and U618 (N_618,In_697,In_57);
or U619 (N_619,In_97,In_597);
or U620 (N_620,In_649,In_598);
and U621 (N_621,In_229,In_252);
nor U622 (N_622,In_683,In_373);
nand U623 (N_623,In_604,In_114);
nor U624 (N_624,In_123,In_403);
and U625 (N_625,In_652,In_47);
nand U626 (N_626,In_99,In_423);
nand U627 (N_627,In_56,In_240);
nor U628 (N_628,In_667,In_609);
nor U629 (N_629,In_11,In_474);
nor U630 (N_630,In_227,In_417);
or U631 (N_631,In_498,In_421);
nand U632 (N_632,In_619,In_630);
nand U633 (N_633,In_622,In_383);
nor U634 (N_634,In_381,In_119);
nand U635 (N_635,In_603,In_631);
nand U636 (N_636,In_272,In_662);
nand U637 (N_637,In_313,In_270);
nor U638 (N_638,In_107,In_225);
or U639 (N_639,In_575,In_396);
and U640 (N_640,In_622,In_675);
nor U641 (N_641,In_508,In_362);
or U642 (N_642,In_145,In_402);
and U643 (N_643,In_363,In_46);
nor U644 (N_644,In_125,In_22);
and U645 (N_645,In_405,In_82);
nand U646 (N_646,In_295,In_271);
nand U647 (N_647,In_277,In_162);
nor U648 (N_648,In_4,In_687);
or U649 (N_649,In_59,In_412);
or U650 (N_650,In_719,In_692);
nor U651 (N_651,In_375,In_393);
and U652 (N_652,In_419,In_46);
and U653 (N_653,In_405,In_331);
nand U654 (N_654,In_2,In_87);
nor U655 (N_655,In_99,In_215);
nor U656 (N_656,In_94,In_714);
nand U657 (N_657,In_148,In_308);
or U658 (N_658,In_377,In_279);
or U659 (N_659,In_30,In_455);
or U660 (N_660,In_453,In_377);
nand U661 (N_661,In_324,In_514);
and U662 (N_662,In_185,In_657);
nor U663 (N_663,In_160,In_218);
nor U664 (N_664,In_248,In_421);
and U665 (N_665,In_551,In_412);
nor U666 (N_666,In_214,In_647);
nand U667 (N_667,In_507,In_65);
and U668 (N_668,In_395,In_43);
and U669 (N_669,In_353,In_532);
nand U670 (N_670,In_492,In_263);
and U671 (N_671,In_209,In_450);
and U672 (N_672,In_89,In_738);
nand U673 (N_673,In_543,In_140);
nor U674 (N_674,In_31,In_739);
or U675 (N_675,In_126,In_250);
nand U676 (N_676,In_394,In_310);
and U677 (N_677,In_648,In_698);
nor U678 (N_678,In_454,In_227);
nor U679 (N_679,In_484,In_5);
and U680 (N_680,In_303,In_549);
nand U681 (N_681,In_417,In_715);
nand U682 (N_682,In_4,In_43);
nand U683 (N_683,In_63,In_353);
and U684 (N_684,In_228,In_282);
nor U685 (N_685,In_136,In_377);
and U686 (N_686,In_704,In_583);
and U687 (N_687,In_523,In_128);
nand U688 (N_688,In_240,In_650);
and U689 (N_689,In_311,In_435);
nand U690 (N_690,In_700,In_158);
or U691 (N_691,In_641,In_671);
or U692 (N_692,In_121,In_562);
or U693 (N_693,In_501,In_82);
and U694 (N_694,In_519,In_304);
or U695 (N_695,In_109,In_98);
nand U696 (N_696,In_687,In_688);
and U697 (N_697,In_355,In_419);
nor U698 (N_698,In_611,In_390);
nand U699 (N_699,In_714,In_146);
and U700 (N_700,In_179,In_552);
and U701 (N_701,In_110,In_719);
and U702 (N_702,In_680,In_38);
nor U703 (N_703,In_73,In_58);
nor U704 (N_704,In_173,In_479);
nor U705 (N_705,In_3,In_724);
nand U706 (N_706,In_39,In_18);
and U707 (N_707,In_105,In_535);
nand U708 (N_708,In_305,In_237);
or U709 (N_709,In_401,In_364);
nor U710 (N_710,In_742,In_712);
nor U711 (N_711,In_528,In_358);
or U712 (N_712,In_692,In_190);
nand U713 (N_713,In_635,In_484);
nand U714 (N_714,In_408,In_698);
and U715 (N_715,In_19,In_363);
or U716 (N_716,In_663,In_332);
nor U717 (N_717,In_477,In_588);
and U718 (N_718,In_599,In_292);
and U719 (N_719,In_469,In_187);
nand U720 (N_720,In_491,In_6);
and U721 (N_721,In_195,In_438);
and U722 (N_722,In_741,In_258);
or U723 (N_723,In_399,In_487);
nand U724 (N_724,In_289,In_95);
and U725 (N_725,In_1,In_263);
or U726 (N_726,In_712,In_650);
or U727 (N_727,In_584,In_472);
nor U728 (N_728,In_741,In_424);
nor U729 (N_729,In_726,In_592);
and U730 (N_730,In_27,In_479);
nand U731 (N_731,In_158,In_598);
or U732 (N_732,In_658,In_236);
and U733 (N_733,In_499,In_235);
and U734 (N_734,In_487,In_174);
xor U735 (N_735,In_184,In_504);
nor U736 (N_736,In_623,In_332);
and U737 (N_737,In_581,In_644);
nor U738 (N_738,In_302,In_326);
nand U739 (N_739,In_275,In_214);
nor U740 (N_740,In_236,In_543);
and U741 (N_741,In_619,In_175);
xor U742 (N_742,In_472,In_572);
nand U743 (N_743,In_1,In_350);
or U744 (N_744,In_194,In_700);
nor U745 (N_745,In_114,In_213);
nand U746 (N_746,In_406,In_613);
and U747 (N_747,In_307,In_120);
and U748 (N_748,In_190,In_238);
nor U749 (N_749,In_565,In_58);
nand U750 (N_750,In_375,In_323);
and U751 (N_751,In_184,In_444);
and U752 (N_752,In_719,In_462);
nand U753 (N_753,In_35,In_390);
nor U754 (N_754,In_577,In_256);
and U755 (N_755,In_270,In_326);
nand U756 (N_756,In_68,In_521);
and U757 (N_757,In_201,In_397);
nand U758 (N_758,In_459,In_60);
and U759 (N_759,In_73,In_704);
nand U760 (N_760,In_22,In_449);
nand U761 (N_761,In_459,In_107);
nor U762 (N_762,In_717,In_732);
xor U763 (N_763,In_566,In_448);
nor U764 (N_764,In_738,In_621);
nor U765 (N_765,In_584,In_325);
nor U766 (N_766,In_154,In_555);
and U767 (N_767,In_506,In_533);
or U768 (N_768,In_709,In_470);
xnor U769 (N_769,In_656,In_510);
nor U770 (N_770,In_664,In_5);
nor U771 (N_771,In_647,In_167);
and U772 (N_772,In_420,In_480);
or U773 (N_773,In_699,In_157);
and U774 (N_774,In_186,In_142);
or U775 (N_775,In_107,In_41);
nand U776 (N_776,In_728,In_556);
or U777 (N_777,In_748,In_65);
nand U778 (N_778,In_103,In_682);
and U779 (N_779,In_510,In_215);
nor U780 (N_780,In_63,In_113);
and U781 (N_781,In_619,In_84);
and U782 (N_782,In_251,In_730);
nand U783 (N_783,In_333,In_630);
or U784 (N_784,In_200,In_570);
or U785 (N_785,In_45,In_315);
and U786 (N_786,In_354,In_337);
or U787 (N_787,In_341,In_647);
nand U788 (N_788,In_456,In_155);
nand U789 (N_789,In_542,In_240);
and U790 (N_790,In_132,In_144);
nand U791 (N_791,In_603,In_461);
or U792 (N_792,In_82,In_649);
nand U793 (N_793,In_380,In_651);
and U794 (N_794,In_144,In_519);
and U795 (N_795,In_430,In_476);
and U796 (N_796,In_614,In_567);
or U797 (N_797,In_429,In_57);
or U798 (N_798,In_345,In_367);
nor U799 (N_799,In_64,In_624);
nor U800 (N_800,In_392,In_511);
nand U801 (N_801,In_542,In_361);
or U802 (N_802,In_721,In_60);
or U803 (N_803,In_712,In_179);
or U804 (N_804,In_662,In_626);
and U805 (N_805,In_97,In_438);
or U806 (N_806,In_220,In_113);
nor U807 (N_807,In_321,In_206);
nand U808 (N_808,In_159,In_390);
and U809 (N_809,In_232,In_690);
nand U810 (N_810,In_100,In_116);
nor U811 (N_811,In_54,In_82);
or U812 (N_812,In_604,In_631);
nand U813 (N_813,In_516,In_1);
or U814 (N_814,In_96,In_91);
nand U815 (N_815,In_150,In_249);
nand U816 (N_816,In_278,In_270);
nand U817 (N_817,In_41,In_266);
nand U818 (N_818,In_569,In_496);
and U819 (N_819,In_118,In_726);
nand U820 (N_820,In_384,In_88);
and U821 (N_821,In_6,In_155);
or U822 (N_822,In_160,In_599);
nor U823 (N_823,In_13,In_328);
nand U824 (N_824,In_465,In_540);
or U825 (N_825,In_4,In_404);
nand U826 (N_826,In_339,In_482);
nand U827 (N_827,In_224,In_144);
nand U828 (N_828,In_320,In_229);
nor U829 (N_829,In_614,In_202);
nand U830 (N_830,In_250,In_381);
or U831 (N_831,In_18,In_144);
nand U832 (N_832,In_478,In_553);
and U833 (N_833,In_371,In_635);
nand U834 (N_834,In_246,In_670);
or U835 (N_835,In_442,In_425);
nand U836 (N_836,In_146,In_696);
nor U837 (N_837,In_734,In_396);
and U838 (N_838,In_696,In_241);
nor U839 (N_839,In_643,In_48);
nor U840 (N_840,In_396,In_398);
and U841 (N_841,In_444,In_450);
or U842 (N_842,In_432,In_347);
or U843 (N_843,In_481,In_436);
and U844 (N_844,In_159,In_327);
or U845 (N_845,In_544,In_516);
and U846 (N_846,In_289,In_390);
nand U847 (N_847,In_241,In_99);
and U848 (N_848,In_87,In_139);
and U849 (N_849,In_328,In_100);
and U850 (N_850,In_285,In_504);
nor U851 (N_851,In_76,In_503);
nor U852 (N_852,In_556,In_8);
or U853 (N_853,In_321,In_699);
nor U854 (N_854,In_280,In_186);
nand U855 (N_855,In_500,In_93);
nor U856 (N_856,In_622,In_315);
nor U857 (N_857,In_741,In_492);
and U858 (N_858,In_462,In_670);
and U859 (N_859,In_413,In_1);
or U860 (N_860,In_488,In_38);
nand U861 (N_861,In_343,In_22);
or U862 (N_862,In_251,In_571);
nor U863 (N_863,In_637,In_514);
or U864 (N_864,In_726,In_148);
nand U865 (N_865,In_604,In_309);
nor U866 (N_866,In_434,In_436);
nor U867 (N_867,In_146,In_549);
or U868 (N_868,In_356,In_16);
nor U869 (N_869,In_222,In_346);
nor U870 (N_870,In_111,In_39);
nor U871 (N_871,In_419,In_638);
and U872 (N_872,In_42,In_132);
nand U873 (N_873,In_565,In_115);
or U874 (N_874,In_702,In_2);
or U875 (N_875,In_149,In_541);
nor U876 (N_876,In_393,In_561);
nand U877 (N_877,In_202,In_1);
or U878 (N_878,In_395,In_487);
nand U879 (N_879,In_720,In_229);
nor U880 (N_880,In_268,In_511);
nor U881 (N_881,In_252,In_136);
nor U882 (N_882,In_112,In_104);
and U883 (N_883,In_587,In_6);
nand U884 (N_884,In_203,In_696);
and U885 (N_885,In_86,In_453);
nor U886 (N_886,In_74,In_427);
and U887 (N_887,In_543,In_279);
or U888 (N_888,In_424,In_647);
or U889 (N_889,In_46,In_635);
nand U890 (N_890,In_243,In_479);
or U891 (N_891,In_403,In_57);
nor U892 (N_892,In_166,In_50);
nor U893 (N_893,In_391,In_665);
nand U894 (N_894,In_355,In_42);
and U895 (N_895,In_148,In_336);
and U896 (N_896,In_212,In_264);
nor U897 (N_897,In_660,In_184);
nand U898 (N_898,In_44,In_264);
nor U899 (N_899,In_230,In_554);
or U900 (N_900,In_468,In_148);
or U901 (N_901,In_233,In_726);
or U902 (N_902,In_119,In_382);
nor U903 (N_903,In_571,In_64);
and U904 (N_904,In_558,In_181);
or U905 (N_905,In_703,In_371);
and U906 (N_906,In_595,In_671);
nand U907 (N_907,In_636,In_8);
nand U908 (N_908,In_422,In_687);
or U909 (N_909,In_543,In_392);
and U910 (N_910,In_437,In_527);
or U911 (N_911,In_506,In_680);
nor U912 (N_912,In_417,In_12);
nand U913 (N_913,In_176,In_128);
nand U914 (N_914,In_657,In_101);
nor U915 (N_915,In_225,In_489);
or U916 (N_916,In_671,In_356);
xnor U917 (N_917,In_313,In_389);
nand U918 (N_918,In_445,In_540);
nor U919 (N_919,In_84,In_121);
nand U920 (N_920,In_424,In_422);
and U921 (N_921,In_41,In_695);
nor U922 (N_922,In_624,In_610);
and U923 (N_923,In_746,In_436);
nor U924 (N_924,In_216,In_471);
and U925 (N_925,In_353,In_545);
or U926 (N_926,In_176,In_520);
and U927 (N_927,In_431,In_218);
or U928 (N_928,In_286,In_205);
and U929 (N_929,In_398,In_659);
and U930 (N_930,In_381,In_151);
and U931 (N_931,In_83,In_262);
or U932 (N_932,In_69,In_526);
and U933 (N_933,In_430,In_523);
and U934 (N_934,In_357,In_369);
or U935 (N_935,In_343,In_428);
and U936 (N_936,In_308,In_379);
nand U937 (N_937,In_640,In_212);
nand U938 (N_938,In_400,In_83);
or U939 (N_939,In_142,In_484);
nand U940 (N_940,In_207,In_691);
nand U941 (N_941,In_588,In_202);
and U942 (N_942,In_377,In_525);
and U943 (N_943,In_124,In_312);
or U944 (N_944,In_550,In_497);
nand U945 (N_945,In_697,In_360);
and U946 (N_946,In_123,In_581);
or U947 (N_947,In_140,In_86);
nand U948 (N_948,In_506,In_435);
and U949 (N_949,In_515,In_475);
nand U950 (N_950,In_290,In_118);
and U951 (N_951,In_314,In_252);
nand U952 (N_952,In_53,In_31);
nor U953 (N_953,In_213,In_604);
nor U954 (N_954,In_714,In_440);
nor U955 (N_955,In_237,In_228);
and U956 (N_956,In_733,In_439);
nor U957 (N_957,In_118,In_584);
nor U958 (N_958,In_360,In_444);
nand U959 (N_959,In_570,In_466);
nand U960 (N_960,In_274,In_557);
nor U961 (N_961,In_413,In_486);
and U962 (N_962,In_682,In_496);
nand U963 (N_963,In_620,In_722);
and U964 (N_964,In_82,In_493);
nor U965 (N_965,In_509,In_670);
and U966 (N_966,In_652,In_143);
nor U967 (N_967,In_285,In_331);
or U968 (N_968,In_392,In_618);
nor U969 (N_969,In_491,In_318);
nor U970 (N_970,In_351,In_66);
nand U971 (N_971,In_702,In_21);
nor U972 (N_972,In_652,In_540);
nor U973 (N_973,In_540,In_282);
nor U974 (N_974,In_714,In_731);
nand U975 (N_975,In_632,In_316);
nand U976 (N_976,In_328,In_177);
nand U977 (N_977,In_401,In_259);
nor U978 (N_978,In_467,In_399);
nor U979 (N_979,In_211,In_457);
nor U980 (N_980,In_624,In_239);
nor U981 (N_981,In_136,In_212);
nor U982 (N_982,In_359,In_13);
or U983 (N_983,In_296,In_315);
nand U984 (N_984,In_75,In_451);
and U985 (N_985,In_538,In_58);
and U986 (N_986,In_45,In_161);
nand U987 (N_987,In_452,In_100);
nand U988 (N_988,In_518,In_494);
nor U989 (N_989,In_174,In_75);
nand U990 (N_990,In_436,In_232);
or U991 (N_991,In_497,In_482);
nor U992 (N_992,In_226,In_197);
or U993 (N_993,In_395,In_624);
or U994 (N_994,In_724,In_739);
or U995 (N_995,In_626,In_131);
and U996 (N_996,In_746,In_58);
nand U997 (N_997,In_511,In_547);
nor U998 (N_998,In_279,In_547);
nand U999 (N_999,In_558,In_57);
nor U1000 (N_1000,In_119,In_348);
nor U1001 (N_1001,In_308,In_375);
nand U1002 (N_1002,In_424,In_293);
and U1003 (N_1003,In_445,In_300);
nand U1004 (N_1004,In_266,In_13);
or U1005 (N_1005,In_521,In_359);
and U1006 (N_1006,In_117,In_719);
or U1007 (N_1007,In_512,In_198);
or U1008 (N_1008,In_355,In_311);
nor U1009 (N_1009,In_731,In_522);
nor U1010 (N_1010,In_148,In_37);
nand U1011 (N_1011,In_310,In_429);
and U1012 (N_1012,In_317,In_233);
and U1013 (N_1013,In_174,In_63);
and U1014 (N_1014,In_193,In_312);
and U1015 (N_1015,In_279,In_527);
nand U1016 (N_1016,In_132,In_73);
and U1017 (N_1017,In_746,In_166);
nor U1018 (N_1018,In_284,In_224);
nor U1019 (N_1019,In_48,In_713);
and U1020 (N_1020,In_398,In_506);
and U1021 (N_1021,In_696,In_132);
nor U1022 (N_1022,In_89,In_385);
nand U1023 (N_1023,In_62,In_521);
nor U1024 (N_1024,In_446,In_253);
or U1025 (N_1025,In_115,In_255);
nor U1026 (N_1026,In_560,In_148);
nor U1027 (N_1027,In_387,In_711);
and U1028 (N_1028,In_585,In_91);
nand U1029 (N_1029,In_724,In_329);
or U1030 (N_1030,In_512,In_73);
nand U1031 (N_1031,In_553,In_503);
and U1032 (N_1032,In_469,In_363);
and U1033 (N_1033,In_730,In_403);
nand U1034 (N_1034,In_694,In_393);
or U1035 (N_1035,In_214,In_272);
nor U1036 (N_1036,In_332,In_38);
nand U1037 (N_1037,In_193,In_106);
nor U1038 (N_1038,In_616,In_528);
and U1039 (N_1039,In_466,In_98);
or U1040 (N_1040,In_79,In_446);
nand U1041 (N_1041,In_589,In_636);
or U1042 (N_1042,In_149,In_163);
xor U1043 (N_1043,In_327,In_593);
and U1044 (N_1044,In_445,In_293);
and U1045 (N_1045,In_264,In_626);
nand U1046 (N_1046,In_274,In_589);
nor U1047 (N_1047,In_219,In_578);
nand U1048 (N_1048,In_169,In_554);
nand U1049 (N_1049,In_387,In_708);
and U1050 (N_1050,In_248,In_361);
nor U1051 (N_1051,In_685,In_91);
nand U1052 (N_1052,In_307,In_448);
and U1053 (N_1053,In_726,In_123);
and U1054 (N_1054,In_126,In_156);
and U1055 (N_1055,In_524,In_288);
or U1056 (N_1056,In_215,In_211);
nor U1057 (N_1057,In_549,In_82);
or U1058 (N_1058,In_143,In_553);
and U1059 (N_1059,In_182,In_38);
and U1060 (N_1060,In_158,In_156);
or U1061 (N_1061,In_116,In_384);
or U1062 (N_1062,In_251,In_578);
nand U1063 (N_1063,In_33,In_696);
nor U1064 (N_1064,In_594,In_344);
or U1065 (N_1065,In_282,In_405);
and U1066 (N_1066,In_701,In_46);
or U1067 (N_1067,In_607,In_692);
nor U1068 (N_1068,In_679,In_158);
nor U1069 (N_1069,In_665,In_667);
and U1070 (N_1070,In_295,In_560);
nand U1071 (N_1071,In_417,In_650);
nor U1072 (N_1072,In_404,In_437);
nand U1073 (N_1073,In_394,In_248);
nand U1074 (N_1074,In_434,In_40);
nor U1075 (N_1075,In_245,In_397);
or U1076 (N_1076,In_134,In_570);
nor U1077 (N_1077,In_745,In_253);
nor U1078 (N_1078,In_381,In_516);
nand U1079 (N_1079,In_269,In_685);
nand U1080 (N_1080,In_719,In_238);
and U1081 (N_1081,In_287,In_289);
or U1082 (N_1082,In_383,In_725);
or U1083 (N_1083,In_421,In_57);
xnor U1084 (N_1084,In_502,In_556);
nand U1085 (N_1085,In_718,In_9);
nand U1086 (N_1086,In_167,In_282);
nor U1087 (N_1087,In_181,In_74);
and U1088 (N_1088,In_715,In_377);
or U1089 (N_1089,In_154,In_87);
or U1090 (N_1090,In_421,In_669);
and U1091 (N_1091,In_555,In_631);
nand U1092 (N_1092,In_311,In_510);
xor U1093 (N_1093,In_288,In_637);
nand U1094 (N_1094,In_239,In_369);
and U1095 (N_1095,In_79,In_304);
nand U1096 (N_1096,In_350,In_102);
nand U1097 (N_1097,In_569,In_466);
xor U1098 (N_1098,In_665,In_87);
or U1099 (N_1099,In_213,In_84);
nand U1100 (N_1100,In_317,In_231);
and U1101 (N_1101,In_731,In_506);
or U1102 (N_1102,In_219,In_661);
nor U1103 (N_1103,In_162,In_78);
nand U1104 (N_1104,In_729,In_69);
or U1105 (N_1105,In_674,In_34);
or U1106 (N_1106,In_337,In_718);
and U1107 (N_1107,In_95,In_135);
nor U1108 (N_1108,In_580,In_279);
and U1109 (N_1109,In_502,In_34);
nor U1110 (N_1110,In_0,In_495);
nand U1111 (N_1111,In_407,In_423);
and U1112 (N_1112,In_634,In_36);
and U1113 (N_1113,In_327,In_517);
nor U1114 (N_1114,In_99,In_284);
or U1115 (N_1115,In_453,In_23);
nor U1116 (N_1116,In_687,In_543);
nand U1117 (N_1117,In_557,In_664);
nand U1118 (N_1118,In_697,In_150);
nor U1119 (N_1119,In_480,In_452);
and U1120 (N_1120,In_356,In_478);
or U1121 (N_1121,In_672,In_115);
nand U1122 (N_1122,In_411,In_741);
nand U1123 (N_1123,In_641,In_406);
nand U1124 (N_1124,In_665,In_118);
nand U1125 (N_1125,In_4,In_466);
nand U1126 (N_1126,In_392,In_238);
and U1127 (N_1127,In_409,In_615);
nor U1128 (N_1128,In_99,In_125);
nand U1129 (N_1129,In_214,In_391);
nor U1130 (N_1130,In_400,In_686);
or U1131 (N_1131,In_654,In_119);
and U1132 (N_1132,In_407,In_90);
and U1133 (N_1133,In_12,In_709);
nand U1134 (N_1134,In_322,In_438);
or U1135 (N_1135,In_101,In_317);
xor U1136 (N_1136,In_474,In_542);
and U1137 (N_1137,In_490,In_171);
and U1138 (N_1138,In_139,In_501);
and U1139 (N_1139,In_353,In_233);
or U1140 (N_1140,In_193,In_272);
nor U1141 (N_1141,In_694,In_733);
nand U1142 (N_1142,In_461,In_674);
and U1143 (N_1143,In_577,In_134);
or U1144 (N_1144,In_549,In_607);
nor U1145 (N_1145,In_688,In_73);
nor U1146 (N_1146,In_354,In_686);
nor U1147 (N_1147,In_534,In_20);
nand U1148 (N_1148,In_728,In_463);
and U1149 (N_1149,In_510,In_70);
and U1150 (N_1150,In_410,In_540);
or U1151 (N_1151,In_691,In_579);
and U1152 (N_1152,In_50,In_275);
or U1153 (N_1153,In_101,In_630);
nand U1154 (N_1154,In_736,In_470);
nor U1155 (N_1155,In_597,In_484);
nor U1156 (N_1156,In_150,In_8);
and U1157 (N_1157,In_414,In_240);
nor U1158 (N_1158,In_168,In_741);
or U1159 (N_1159,In_159,In_639);
and U1160 (N_1160,In_218,In_535);
nor U1161 (N_1161,In_175,In_684);
xnor U1162 (N_1162,In_512,In_618);
and U1163 (N_1163,In_266,In_39);
or U1164 (N_1164,In_352,In_141);
and U1165 (N_1165,In_174,In_407);
nand U1166 (N_1166,In_611,In_590);
nor U1167 (N_1167,In_700,In_663);
or U1168 (N_1168,In_279,In_494);
and U1169 (N_1169,In_562,In_733);
or U1170 (N_1170,In_104,In_80);
or U1171 (N_1171,In_268,In_603);
xor U1172 (N_1172,In_606,In_53);
nand U1173 (N_1173,In_692,In_315);
or U1174 (N_1174,In_63,In_99);
nor U1175 (N_1175,In_141,In_493);
nor U1176 (N_1176,In_64,In_653);
or U1177 (N_1177,In_536,In_577);
nor U1178 (N_1178,In_78,In_520);
nor U1179 (N_1179,In_181,In_23);
nand U1180 (N_1180,In_424,In_34);
nor U1181 (N_1181,In_315,In_291);
and U1182 (N_1182,In_76,In_75);
and U1183 (N_1183,In_19,In_390);
or U1184 (N_1184,In_708,In_608);
and U1185 (N_1185,In_718,In_685);
or U1186 (N_1186,In_283,In_200);
nor U1187 (N_1187,In_725,In_341);
nand U1188 (N_1188,In_70,In_194);
nor U1189 (N_1189,In_667,In_695);
and U1190 (N_1190,In_169,In_330);
nand U1191 (N_1191,In_92,In_342);
nor U1192 (N_1192,In_194,In_66);
and U1193 (N_1193,In_197,In_127);
xor U1194 (N_1194,In_449,In_418);
and U1195 (N_1195,In_318,In_659);
and U1196 (N_1196,In_35,In_301);
nand U1197 (N_1197,In_309,In_671);
nand U1198 (N_1198,In_699,In_559);
and U1199 (N_1199,In_305,In_688);
nor U1200 (N_1200,In_104,In_565);
and U1201 (N_1201,In_330,In_63);
or U1202 (N_1202,In_10,In_481);
nand U1203 (N_1203,In_356,In_643);
and U1204 (N_1204,In_430,In_291);
nand U1205 (N_1205,In_160,In_534);
or U1206 (N_1206,In_128,In_391);
nand U1207 (N_1207,In_242,In_709);
nand U1208 (N_1208,In_151,In_581);
nor U1209 (N_1209,In_166,In_121);
nand U1210 (N_1210,In_4,In_112);
and U1211 (N_1211,In_10,In_352);
and U1212 (N_1212,In_481,In_623);
or U1213 (N_1213,In_159,In_662);
and U1214 (N_1214,In_345,In_138);
and U1215 (N_1215,In_333,In_212);
and U1216 (N_1216,In_202,In_595);
and U1217 (N_1217,In_457,In_445);
and U1218 (N_1218,In_678,In_160);
nand U1219 (N_1219,In_543,In_198);
nand U1220 (N_1220,In_589,In_466);
or U1221 (N_1221,In_326,In_274);
or U1222 (N_1222,In_326,In_9);
nor U1223 (N_1223,In_622,In_533);
and U1224 (N_1224,In_647,In_24);
nor U1225 (N_1225,In_125,In_483);
nor U1226 (N_1226,In_18,In_365);
nor U1227 (N_1227,In_451,In_465);
or U1228 (N_1228,In_74,In_421);
nand U1229 (N_1229,In_334,In_744);
nor U1230 (N_1230,In_225,In_724);
and U1231 (N_1231,In_487,In_591);
nor U1232 (N_1232,In_177,In_385);
and U1233 (N_1233,In_553,In_24);
and U1234 (N_1234,In_58,In_583);
or U1235 (N_1235,In_545,In_604);
or U1236 (N_1236,In_515,In_531);
and U1237 (N_1237,In_150,In_144);
and U1238 (N_1238,In_587,In_514);
nor U1239 (N_1239,In_153,In_319);
or U1240 (N_1240,In_701,In_207);
or U1241 (N_1241,In_586,In_344);
and U1242 (N_1242,In_619,In_736);
and U1243 (N_1243,In_193,In_567);
nor U1244 (N_1244,In_380,In_17);
or U1245 (N_1245,In_437,In_357);
xnor U1246 (N_1246,In_670,In_146);
and U1247 (N_1247,In_704,In_180);
or U1248 (N_1248,In_722,In_396);
or U1249 (N_1249,In_141,In_578);
or U1250 (N_1250,In_100,In_208);
or U1251 (N_1251,In_670,In_480);
and U1252 (N_1252,In_91,In_488);
or U1253 (N_1253,In_472,In_596);
and U1254 (N_1254,In_75,In_573);
nand U1255 (N_1255,In_233,In_554);
or U1256 (N_1256,In_649,In_412);
and U1257 (N_1257,In_295,In_619);
or U1258 (N_1258,In_416,In_558);
or U1259 (N_1259,In_175,In_211);
or U1260 (N_1260,In_370,In_610);
or U1261 (N_1261,In_290,In_109);
and U1262 (N_1262,In_510,In_439);
and U1263 (N_1263,In_588,In_279);
nand U1264 (N_1264,In_673,In_571);
nand U1265 (N_1265,In_489,In_68);
nand U1266 (N_1266,In_37,In_283);
nor U1267 (N_1267,In_15,In_126);
nor U1268 (N_1268,In_571,In_235);
and U1269 (N_1269,In_291,In_8);
and U1270 (N_1270,In_582,In_187);
or U1271 (N_1271,In_184,In_568);
nand U1272 (N_1272,In_141,In_85);
and U1273 (N_1273,In_469,In_444);
or U1274 (N_1274,In_581,In_538);
nand U1275 (N_1275,In_662,In_458);
and U1276 (N_1276,In_478,In_296);
nand U1277 (N_1277,In_3,In_509);
nand U1278 (N_1278,In_464,In_655);
and U1279 (N_1279,In_729,In_302);
and U1280 (N_1280,In_160,In_558);
nand U1281 (N_1281,In_38,In_725);
and U1282 (N_1282,In_357,In_255);
nor U1283 (N_1283,In_254,In_331);
and U1284 (N_1284,In_360,In_300);
and U1285 (N_1285,In_221,In_519);
and U1286 (N_1286,In_462,In_308);
or U1287 (N_1287,In_125,In_16);
nor U1288 (N_1288,In_307,In_415);
or U1289 (N_1289,In_704,In_260);
and U1290 (N_1290,In_710,In_718);
and U1291 (N_1291,In_123,In_700);
nor U1292 (N_1292,In_711,In_160);
nor U1293 (N_1293,In_657,In_621);
nor U1294 (N_1294,In_459,In_249);
xor U1295 (N_1295,In_128,In_531);
nand U1296 (N_1296,In_512,In_382);
nor U1297 (N_1297,In_396,In_747);
and U1298 (N_1298,In_572,In_387);
nor U1299 (N_1299,In_442,In_236);
nor U1300 (N_1300,In_599,In_206);
nand U1301 (N_1301,In_275,In_600);
nor U1302 (N_1302,In_406,In_394);
nor U1303 (N_1303,In_542,In_644);
nand U1304 (N_1304,In_346,In_102);
or U1305 (N_1305,In_719,In_172);
nand U1306 (N_1306,In_171,In_40);
nor U1307 (N_1307,In_579,In_314);
nor U1308 (N_1308,In_603,In_409);
nor U1309 (N_1309,In_169,In_605);
or U1310 (N_1310,In_576,In_684);
nand U1311 (N_1311,In_47,In_302);
nor U1312 (N_1312,In_395,In_80);
nor U1313 (N_1313,In_631,In_628);
or U1314 (N_1314,In_219,In_363);
nand U1315 (N_1315,In_584,In_613);
nand U1316 (N_1316,In_284,In_617);
nand U1317 (N_1317,In_74,In_354);
and U1318 (N_1318,In_644,In_246);
or U1319 (N_1319,In_122,In_47);
or U1320 (N_1320,In_487,In_25);
nor U1321 (N_1321,In_203,In_353);
nand U1322 (N_1322,In_603,In_626);
nand U1323 (N_1323,In_112,In_555);
and U1324 (N_1324,In_744,In_521);
or U1325 (N_1325,In_587,In_166);
or U1326 (N_1326,In_561,In_485);
nand U1327 (N_1327,In_263,In_103);
nand U1328 (N_1328,In_321,In_251);
and U1329 (N_1329,In_317,In_134);
or U1330 (N_1330,In_224,In_98);
nand U1331 (N_1331,In_400,In_390);
or U1332 (N_1332,In_229,In_158);
or U1333 (N_1333,In_686,In_747);
nand U1334 (N_1334,In_258,In_298);
nand U1335 (N_1335,In_612,In_61);
or U1336 (N_1336,In_719,In_737);
or U1337 (N_1337,In_564,In_32);
nor U1338 (N_1338,In_433,In_418);
and U1339 (N_1339,In_216,In_288);
nor U1340 (N_1340,In_81,In_74);
or U1341 (N_1341,In_726,In_259);
or U1342 (N_1342,In_409,In_13);
or U1343 (N_1343,In_133,In_706);
nand U1344 (N_1344,In_36,In_347);
and U1345 (N_1345,In_303,In_623);
or U1346 (N_1346,In_513,In_248);
or U1347 (N_1347,In_318,In_193);
or U1348 (N_1348,In_233,In_51);
nand U1349 (N_1349,In_701,In_469);
nand U1350 (N_1350,In_573,In_703);
nand U1351 (N_1351,In_524,In_535);
nor U1352 (N_1352,In_368,In_59);
nand U1353 (N_1353,In_741,In_441);
and U1354 (N_1354,In_231,In_568);
and U1355 (N_1355,In_475,In_52);
nor U1356 (N_1356,In_435,In_710);
nor U1357 (N_1357,In_452,In_312);
nand U1358 (N_1358,In_499,In_202);
or U1359 (N_1359,In_64,In_159);
nand U1360 (N_1360,In_103,In_510);
or U1361 (N_1361,In_173,In_460);
and U1362 (N_1362,In_493,In_193);
nor U1363 (N_1363,In_651,In_270);
nor U1364 (N_1364,In_422,In_130);
or U1365 (N_1365,In_424,In_385);
nor U1366 (N_1366,In_740,In_445);
nor U1367 (N_1367,In_538,In_313);
nor U1368 (N_1368,In_332,In_693);
and U1369 (N_1369,In_625,In_465);
nand U1370 (N_1370,In_160,In_273);
or U1371 (N_1371,In_394,In_714);
nor U1372 (N_1372,In_93,In_240);
nor U1373 (N_1373,In_63,In_195);
nand U1374 (N_1374,In_237,In_137);
or U1375 (N_1375,In_595,In_76);
nand U1376 (N_1376,In_550,In_54);
nand U1377 (N_1377,In_620,In_107);
nand U1378 (N_1378,In_300,In_214);
and U1379 (N_1379,In_433,In_703);
and U1380 (N_1380,In_500,In_485);
nor U1381 (N_1381,In_160,In_491);
or U1382 (N_1382,In_332,In_383);
nand U1383 (N_1383,In_243,In_117);
and U1384 (N_1384,In_696,In_735);
or U1385 (N_1385,In_615,In_484);
or U1386 (N_1386,In_436,In_250);
and U1387 (N_1387,In_359,In_569);
or U1388 (N_1388,In_436,In_46);
nand U1389 (N_1389,In_749,In_569);
and U1390 (N_1390,In_487,In_185);
nor U1391 (N_1391,In_333,In_502);
or U1392 (N_1392,In_227,In_528);
nor U1393 (N_1393,In_648,In_725);
or U1394 (N_1394,In_226,In_557);
and U1395 (N_1395,In_216,In_314);
nand U1396 (N_1396,In_159,In_407);
and U1397 (N_1397,In_320,In_306);
nand U1398 (N_1398,In_724,In_224);
or U1399 (N_1399,In_670,In_735);
or U1400 (N_1400,In_511,In_34);
nor U1401 (N_1401,In_573,In_587);
nand U1402 (N_1402,In_60,In_574);
nor U1403 (N_1403,In_229,In_240);
or U1404 (N_1404,In_646,In_27);
nor U1405 (N_1405,In_93,In_386);
and U1406 (N_1406,In_355,In_305);
nor U1407 (N_1407,In_220,In_329);
or U1408 (N_1408,In_725,In_177);
xnor U1409 (N_1409,In_660,In_129);
nor U1410 (N_1410,In_422,In_216);
nand U1411 (N_1411,In_668,In_2);
and U1412 (N_1412,In_656,In_159);
or U1413 (N_1413,In_433,In_526);
nand U1414 (N_1414,In_656,In_739);
nor U1415 (N_1415,In_247,In_12);
nor U1416 (N_1416,In_313,In_547);
or U1417 (N_1417,In_686,In_38);
and U1418 (N_1418,In_449,In_212);
xnor U1419 (N_1419,In_589,In_432);
or U1420 (N_1420,In_672,In_675);
and U1421 (N_1421,In_247,In_395);
or U1422 (N_1422,In_31,In_19);
and U1423 (N_1423,In_735,In_593);
or U1424 (N_1424,In_669,In_668);
or U1425 (N_1425,In_749,In_561);
and U1426 (N_1426,In_94,In_258);
nand U1427 (N_1427,In_319,In_205);
or U1428 (N_1428,In_644,In_187);
and U1429 (N_1429,In_278,In_153);
nand U1430 (N_1430,In_611,In_424);
nor U1431 (N_1431,In_21,In_392);
and U1432 (N_1432,In_336,In_519);
and U1433 (N_1433,In_487,In_71);
xor U1434 (N_1434,In_381,In_535);
and U1435 (N_1435,In_687,In_546);
nand U1436 (N_1436,In_159,In_0);
nor U1437 (N_1437,In_378,In_387);
nor U1438 (N_1438,In_232,In_6);
and U1439 (N_1439,In_482,In_49);
and U1440 (N_1440,In_466,In_438);
nor U1441 (N_1441,In_669,In_717);
nor U1442 (N_1442,In_658,In_598);
or U1443 (N_1443,In_335,In_555);
xnor U1444 (N_1444,In_293,In_171);
nor U1445 (N_1445,In_347,In_56);
and U1446 (N_1446,In_485,In_748);
or U1447 (N_1447,In_482,In_347);
and U1448 (N_1448,In_221,In_689);
and U1449 (N_1449,In_339,In_435);
or U1450 (N_1450,In_345,In_621);
nor U1451 (N_1451,In_219,In_237);
or U1452 (N_1452,In_381,In_218);
and U1453 (N_1453,In_678,In_358);
nand U1454 (N_1454,In_394,In_723);
nor U1455 (N_1455,In_76,In_340);
xnor U1456 (N_1456,In_407,In_85);
and U1457 (N_1457,In_587,In_389);
and U1458 (N_1458,In_281,In_627);
nor U1459 (N_1459,In_401,In_170);
nand U1460 (N_1460,In_238,In_292);
and U1461 (N_1461,In_275,In_585);
nor U1462 (N_1462,In_325,In_615);
nand U1463 (N_1463,In_57,In_24);
and U1464 (N_1464,In_118,In_181);
nor U1465 (N_1465,In_550,In_452);
nor U1466 (N_1466,In_213,In_283);
nor U1467 (N_1467,In_146,In_641);
nand U1468 (N_1468,In_364,In_376);
or U1469 (N_1469,In_239,In_434);
nor U1470 (N_1470,In_77,In_600);
and U1471 (N_1471,In_312,In_65);
and U1472 (N_1472,In_741,In_504);
nor U1473 (N_1473,In_589,In_229);
nor U1474 (N_1474,In_574,In_269);
or U1475 (N_1475,In_629,In_167);
or U1476 (N_1476,In_552,In_749);
nand U1477 (N_1477,In_120,In_358);
nor U1478 (N_1478,In_386,In_295);
or U1479 (N_1479,In_463,In_733);
nand U1480 (N_1480,In_296,In_0);
and U1481 (N_1481,In_325,In_146);
nor U1482 (N_1482,In_202,In_389);
nand U1483 (N_1483,In_508,In_335);
and U1484 (N_1484,In_345,In_268);
nor U1485 (N_1485,In_648,In_537);
nand U1486 (N_1486,In_370,In_112);
nand U1487 (N_1487,In_588,In_700);
nand U1488 (N_1488,In_748,In_665);
and U1489 (N_1489,In_199,In_542);
and U1490 (N_1490,In_106,In_139);
or U1491 (N_1491,In_60,In_63);
nand U1492 (N_1492,In_159,In_247);
nand U1493 (N_1493,In_195,In_282);
nand U1494 (N_1494,In_444,In_537);
or U1495 (N_1495,In_65,In_361);
nand U1496 (N_1496,In_690,In_97);
nand U1497 (N_1497,In_526,In_234);
and U1498 (N_1498,In_174,In_11);
nor U1499 (N_1499,In_349,In_447);
and U1500 (N_1500,In_654,In_545);
and U1501 (N_1501,In_103,In_310);
nand U1502 (N_1502,In_464,In_419);
nor U1503 (N_1503,In_549,In_78);
nand U1504 (N_1504,In_168,In_157);
nor U1505 (N_1505,In_436,In_125);
or U1506 (N_1506,In_503,In_429);
and U1507 (N_1507,In_238,In_597);
or U1508 (N_1508,In_550,In_283);
nand U1509 (N_1509,In_130,In_451);
nor U1510 (N_1510,In_667,In_686);
or U1511 (N_1511,In_88,In_43);
nor U1512 (N_1512,In_36,In_516);
nor U1513 (N_1513,In_556,In_222);
or U1514 (N_1514,In_346,In_572);
and U1515 (N_1515,In_268,In_157);
or U1516 (N_1516,In_337,In_608);
or U1517 (N_1517,In_310,In_511);
nand U1518 (N_1518,In_1,In_30);
nor U1519 (N_1519,In_344,In_266);
nand U1520 (N_1520,In_377,In_163);
or U1521 (N_1521,In_588,In_349);
nor U1522 (N_1522,In_376,In_573);
nand U1523 (N_1523,In_18,In_10);
or U1524 (N_1524,In_487,In_91);
nand U1525 (N_1525,In_703,In_231);
nand U1526 (N_1526,In_69,In_57);
and U1527 (N_1527,In_154,In_582);
or U1528 (N_1528,In_710,In_733);
xnor U1529 (N_1529,In_242,In_208);
nand U1530 (N_1530,In_411,In_571);
nor U1531 (N_1531,In_380,In_656);
xor U1532 (N_1532,In_352,In_186);
and U1533 (N_1533,In_393,In_265);
and U1534 (N_1534,In_234,In_583);
or U1535 (N_1535,In_702,In_258);
nand U1536 (N_1536,In_678,In_31);
nor U1537 (N_1537,In_363,In_105);
and U1538 (N_1538,In_4,In_125);
nor U1539 (N_1539,In_249,In_95);
and U1540 (N_1540,In_320,In_551);
and U1541 (N_1541,In_319,In_389);
or U1542 (N_1542,In_20,In_225);
or U1543 (N_1543,In_619,In_588);
or U1544 (N_1544,In_670,In_76);
and U1545 (N_1545,In_166,In_602);
nand U1546 (N_1546,In_165,In_732);
nand U1547 (N_1547,In_314,In_482);
and U1548 (N_1548,In_14,In_739);
or U1549 (N_1549,In_652,In_89);
and U1550 (N_1550,In_408,In_371);
nand U1551 (N_1551,In_621,In_269);
nand U1552 (N_1552,In_46,In_518);
or U1553 (N_1553,In_476,In_623);
nor U1554 (N_1554,In_226,In_692);
or U1555 (N_1555,In_103,In_467);
nor U1556 (N_1556,In_136,In_209);
and U1557 (N_1557,In_233,In_121);
or U1558 (N_1558,In_164,In_534);
or U1559 (N_1559,In_317,In_406);
xor U1560 (N_1560,In_563,In_450);
or U1561 (N_1561,In_584,In_652);
nand U1562 (N_1562,In_76,In_259);
and U1563 (N_1563,In_150,In_389);
and U1564 (N_1564,In_353,In_148);
nand U1565 (N_1565,In_180,In_705);
nor U1566 (N_1566,In_626,In_207);
or U1567 (N_1567,In_608,In_603);
nand U1568 (N_1568,In_148,In_346);
nor U1569 (N_1569,In_479,In_203);
or U1570 (N_1570,In_638,In_402);
and U1571 (N_1571,In_103,In_666);
nand U1572 (N_1572,In_120,In_403);
or U1573 (N_1573,In_479,In_56);
or U1574 (N_1574,In_502,In_39);
or U1575 (N_1575,In_604,In_65);
nor U1576 (N_1576,In_309,In_724);
or U1577 (N_1577,In_467,In_514);
nor U1578 (N_1578,In_741,In_129);
nor U1579 (N_1579,In_638,In_278);
nand U1580 (N_1580,In_303,In_15);
nand U1581 (N_1581,In_186,In_251);
nor U1582 (N_1582,In_308,In_438);
or U1583 (N_1583,In_514,In_591);
or U1584 (N_1584,In_67,In_405);
nor U1585 (N_1585,In_130,In_294);
and U1586 (N_1586,In_507,In_207);
or U1587 (N_1587,In_388,In_446);
and U1588 (N_1588,In_21,In_532);
nor U1589 (N_1589,In_543,In_138);
nor U1590 (N_1590,In_433,In_212);
and U1591 (N_1591,In_511,In_308);
nor U1592 (N_1592,In_722,In_497);
nor U1593 (N_1593,In_197,In_27);
nand U1594 (N_1594,In_583,In_615);
or U1595 (N_1595,In_321,In_118);
and U1596 (N_1596,In_395,In_235);
or U1597 (N_1597,In_741,In_450);
or U1598 (N_1598,In_642,In_109);
nand U1599 (N_1599,In_726,In_427);
or U1600 (N_1600,In_425,In_620);
or U1601 (N_1601,In_34,In_256);
or U1602 (N_1602,In_192,In_471);
or U1603 (N_1603,In_112,In_661);
and U1604 (N_1604,In_346,In_219);
nand U1605 (N_1605,In_20,In_578);
nand U1606 (N_1606,In_172,In_291);
nor U1607 (N_1607,In_510,In_397);
nand U1608 (N_1608,In_620,In_482);
nand U1609 (N_1609,In_682,In_25);
and U1610 (N_1610,In_507,In_217);
nor U1611 (N_1611,In_135,In_301);
nor U1612 (N_1612,In_378,In_403);
nor U1613 (N_1613,In_745,In_10);
nor U1614 (N_1614,In_136,In_18);
or U1615 (N_1615,In_152,In_85);
and U1616 (N_1616,In_101,In_0);
nand U1617 (N_1617,In_576,In_340);
or U1618 (N_1618,In_170,In_557);
nand U1619 (N_1619,In_609,In_578);
and U1620 (N_1620,In_470,In_191);
or U1621 (N_1621,In_664,In_19);
and U1622 (N_1622,In_397,In_445);
and U1623 (N_1623,In_328,In_88);
nand U1624 (N_1624,In_450,In_733);
nand U1625 (N_1625,In_499,In_164);
nor U1626 (N_1626,In_31,In_469);
nand U1627 (N_1627,In_365,In_590);
and U1628 (N_1628,In_559,In_120);
and U1629 (N_1629,In_55,In_184);
nor U1630 (N_1630,In_18,In_522);
nand U1631 (N_1631,In_212,In_34);
nor U1632 (N_1632,In_316,In_339);
and U1633 (N_1633,In_603,In_289);
nand U1634 (N_1634,In_647,In_330);
nor U1635 (N_1635,In_409,In_57);
and U1636 (N_1636,In_366,In_565);
nand U1637 (N_1637,In_654,In_25);
nor U1638 (N_1638,In_680,In_391);
nand U1639 (N_1639,In_317,In_491);
and U1640 (N_1640,In_26,In_66);
nand U1641 (N_1641,In_329,In_19);
nand U1642 (N_1642,In_166,In_291);
and U1643 (N_1643,In_97,In_567);
or U1644 (N_1644,In_67,In_392);
nand U1645 (N_1645,In_218,In_202);
nand U1646 (N_1646,In_38,In_96);
nand U1647 (N_1647,In_68,In_421);
nand U1648 (N_1648,In_303,In_422);
nor U1649 (N_1649,In_138,In_173);
nand U1650 (N_1650,In_605,In_696);
nor U1651 (N_1651,In_333,In_350);
and U1652 (N_1652,In_745,In_230);
nand U1653 (N_1653,In_473,In_301);
or U1654 (N_1654,In_219,In_125);
and U1655 (N_1655,In_488,In_507);
or U1656 (N_1656,In_208,In_651);
nor U1657 (N_1657,In_9,In_319);
and U1658 (N_1658,In_379,In_380);
nand U1659 (N_1659,In_141,In_496);
and U1660 (N_1660,In_551,In_316);
nand U1661 (N_1661,In_403,In_641);
nor U1662 (N_1662,In_674,In_579);
nand U1663 (N_1663,In_193,In_302);
or U1664 (N_1664,In_213,In_74);
or U1665 (N_1665,In_230,In_222);
and U1666 (N_1666,In_537,In_315);
or U1667 (N_1667,In_464,In_713);
nor U1668 (N_1668,In_382,In_19);
nand U1669 (N_1669,In_46,In_614);
and U1670 (N_1670,In_648,In_188);
nand U1671 (N_1671,In_401,In_699);
nand U1672 (N_1672,In_249,In_556);
nor U1673 (N_1673,In_480,In_26);
and U1674 (N_1674,In_608,In_718);
and U1675 (N_1675,In_251,In_156);
nand U1676 (N_1676,In_227,In_232);
and U1677 (N_1677,In_456,In_78);
or U1678 (N_1678,In_422,In_648);
or U1679 (N_1679,In_481,In_202);
and U1680 (N_1680,In_52,In_258);
and U1681 (N_1681,In_50,In_723);
nor U1682 (N_1682,In_162,In_58);
nor U1683 (N_1683,In_582,In_580);
and U1684 (N_1684,In_212,In_402);
nand U1685 (N_1685,In_346,In_336);
nor U1686 (N_1686,In_11,In_505);
or U1687 (N_1687,In_328,In_381);
nor U1688 (N_1688,In_703,In_406);
nor U1689 (N_1689,In_644,In_407);
and U1690 (N_1690,In_333,In_362);
or U1691 (N_1691,In_371,In_405);
and U1692 (N_1692,In_535,In_172);
and U1693 (N_1693,In_353,In_218);
and U1694 (N_1694,In_49,In_470);
or U1695 (N_1695,In_327,In_300);
nor U1696 (N_1696,In_210,In_600);
or U1697 (N_1697,In_524,In_608);
nor U1698 (N_1698,In_701,In_172);
nor U1699 (N_1699,In_540,In_702);
nand U1700 (N_1700,In_124,In_10);
nand U1701 (N_1701,In_724,In_273);
and U1702 (N_1702,In_625,In_482);
and U1703 (N_1703,In_672,In_325);
and U1704 (N_1704,In_401,In_674);
or U1705 (N_1705,In_466,In_553);
nand U1706 (N_1706,In_76,In_458);
and U1707 (N_1707,In_468,In_414);
nor U1708 (N_1708,In_505,In_334);
nand U1709 (N_1709,In_555,In_651);
and U1710 (N_1710,In_285,In_7);
or U1711 (N_1711,In_627,In_623);
and U1712 (N_1712,In_166,In_675);
nor U1713 (N_1713,In_248,In_605);
nor U1714 (N_1714,In_420,In_523);
or U1715 (N_1715,In_151,In_272);
and U1716 (N_1716,In_94,In_236);
nand U1717 (N_1717,In_692,In_560);
nand U1718 (N_1718,In_222,In_683);
and U1719 (N_1719,In_67,In_731);
and U1720 (N_1720,In_130,In_559);
or U1721 (N_1721,In_173,In_622);
nand U1722 (N_1722,In_572,In_527);
nor U1723 (N_1723,In_644,In_237);
nor U1724 (N_1724,In_58,In_622);
nand U1725 (N_1725,In_16,In_187);
and U1726 (N_1726,In_46,In_739);
nand U1727 (N_1727,In_250,In_256);
or U1728 (N_1728,In_31,In_236);
or U1729 (N_1729,In_364,In_61);
nor U1730 (N_1730,In_112,In_289);
and U1731 (N_1731,In_501,In_477);
nor U1732 (N_1732,In_140,In_714);
and U1733 (N_1733,In_508,In_17);
or U1734 (N_1734,In_373,In_353);
or U1735 (N_1735,In_376,In_304);
or U1736 (N_1736,In_172,In_80);
nor U1737 (N_1737,In_301,In_27);
and U1738 (N_1738,In_170,In_165);
nand U1739 (N_1739,In_72,In_315);
nand U1740 (N_1740,In_611,In_632);
and U1741 (N_1741,In_728,In_611);
nand U1742 (N_1742,In_551,In_120);
nor U1743 (N_1743,In_422,In_547);
and U1744 (N_1744,In_225,In_418);
nand U1745 (N_1745,In_344,In_90);
or U1746 (N_1746,In_65,In_283);
nor U1747 (N_1747,In_324,In_197);
or U1748 (N_1748,In_731,In_159);
or U1749 (N_1749,In_126,In_176);
or U1750 (N_1750,In_192,In_455);
or U1751 (N_1751,In_199,In_35);
and U1752 (N_1752,In_64,In_132);
and U1753 (N_1753,In_3,In_425);
nor U1754 (N_1754,In_367,In_359);
or U1755 (N_1755,In_313,In_391);
nor U1756 (N_1756,In_327,In_653);
nor U1757 (N_1757,In_319,In_542);
or U1758 (N_1758,In_335,In_606);
or U1759 (N_1759,In_517,In_120);
xor U1760 (N_1760,In_311,In_505);
and U1761 (N_1761,In_129,In_396);
or U1762 (N_1762,In_573,In_64);
and U1763 (N_1763,In_583,In_635);
nor U1764 (N_1764,In_328,In_185);
and U1765 (N_1765,In_468,In_129);
nor U1766 (N_1766,In_719,In_45);
or U1767 (N_1767,In_573,In_339);
nand U1768 (N_1768,In_201,In_273);
nor U1769 (N_1769,In_458,In_531);
and U1770 (N_1770,In_59,In_406);
and U1771 (N_1771,In_76,In_344);
or U1772 (N_1772,In_243,In_335);
nand U1773 (N_1773,In_453,In_188);
nand U1774 (N_1774,In_307,In_108);
nand U1775 (N_1775,In_96,In_443);
nand U1776 (N_1776,In_111,In_749);
and U1777 (N_1777,In_726,In_481);
and U1778 (N_1778,In_172,In_224);
nor U1779 (N_1779,In_282,In_183);
or U1780 (N_1780,In_478,In_143);
nand U1781 (N_1781,In_676,In_191);
and U1782 (N_1782,In_695,In_522);
nand U1783 (N_1783,In_745,In_631);
nor U1784 (N_1784,In_236,In_517);
nand U1785 (N_1785,In_290,In_460);
nand U1786 (N_1786,In_375,In_444);
and U1787 (N_1787,In_612,In_532);
and U1788 (N_1788,In_705,In_625);
nand U1789 (N_1789,In_244,In_200);
nor U1790 (N_1790,In_113,In_270);
nor U1791 (N_1791,In_404,In_745);
or U1792 (N_1792,In_631,In_521);
and U1793 (N_1793,In_492,In_74);
or U1794 (N_1794,In_585,In_584);
nand U1795 (N_1795,In_705,In_452);
and U1796 (N_1796,In_586,In_248);
nor U1797 (N_1797,In_320,In_371);
nand U1798 (N_1798,In_207,In_322);
or U1799 (N_1799,In_402,In_323);
and U1800 (N_1800,In_502,In_169);
or U1801 (N_1801,In_165,In_700);
or U1802 (N_1802,In_6,In_105);
nor U1803 (N_1803,In_206,In_655);
and U1804 (N_1804,In_721,In_487);
nor U1805 (N_1805,In_275,In_675);
or U1806 (N_1806,In_302,In_252);
and U1807 (N_1807,In_63,In_662);
nor U1808 (N_1808,In_374,In_574);
nor U1809 (N_1809,In_741,In_135);
or U1810 (N_1810,In_721,In_192);
nor U1811 (N_1811,In_243,In_722);
and U1812 (N_1812,In_49,In_339);
nor U1813 (N_1813,In_404,In_555);
or U1814 (N_1814,In_497,In_397);
nand U1815 (N_1815,In_727,In_645);
xnor U1816 (N_1816,In_309,In_5);
nand U1817 (N_1817,In_65,In_709);
and U1818 (N_1818,In_366,In_412);
nor U1819 (N_1819,In_228,In_400);
or U1820 (N_1820,In_325,In_391);
nand U1821 (N_1821,In_59,In_701);
and U1822 (N_1822,In_600,In_375);
nor U1823 (N_1823,In_79,In_578);
nor U1824 (N_1824,In_314,In_529);
nor U1825 (N_1825,In_304,In_187);
or U1826 (N_1826,In_326,In_170);
nand U1827 (N_1827,In_440,In_445);
nor U1828 (N_1828,In_126,In_297);
or U1829 (N_1829,In_517,In_125);
nand U1830 (N_1830,In_322,In_159);
or U1831 (N_1831,In_609,In_535);
xnor U1832 (N_1832,In_703,In_222);
and U1833 (N_1833,In_602,In_389);
nand U1834 (N_1834,In_321,In_451);
and U1835 (N_1835,In_188,In_248);
and U1836 (N_1836,In_323,In_483);
nand U1837 (N_1837,In_269,In_503);
or U1838 (N_1838,In_190,In_194);
nand U1839 (N_1839,In_260,In_379);
nand U1840 (N_1840,In_151,In_719);
or U1841 (N_1841,In_531,In_339);
nor U1842 (N_1842,In_622,In_268);
nor U1843 (N_1843,In_465,In_537);
or U1844 (N_1844,In_517,In_131);
nor U1845 (N_1845,In_100,In_31);
nand U1846 (N_1846,In_166,In_214);
nand U1847 (N_1847,In_254,In_452);
nand U1848 (N_1848,In_447,In_639);
nor U1849 (N_1849,In_685,In_36);
xnor U1850 (N_1850,In_117,In_75);
and U1851 (N_1851,In_305,In_590);
nor U1852 (N_1852,In_346,In_720);
nand U1853 (N_1853,In_194,In_50);
or U1854 (N_1854,In_3,In_18);
nand U1855 (N_1855,In_381,In_126);
or U1856 (N_1856,In_525,In_403);
nor U1857 (N_1857,In_538,In_78);
nor U1858 (N_1858,In_317,In_220);
nand U1859 (N_1859,In_177,In_257);
and U1860 (N_1860,In_373,In_617);
and U1861 (N_1861,In_525,In_197);
and U1862 (N_1862,In_674,In_519);
and U1863 (N_1863,In_131,In_583);
nand U1864 (N_1864,In_130,In_551);
nor U1865 (N_1865,In_462,In_704);
nor U1866 (N_1866,In_388,In_216);
or U1867 (N_1867,In_218,In_390);
nor U1868 (N_1868,In_632,In_447);
nand U1869 (N_1869,In_43,In_521);
nand U1870 (N_1870,In_516,In_427);
nor U1871 (N_1871,In_212,In_191);
and U1872 (N_1872,In_254,In_31);
nand U1873 (N_1873,In_133,In_111);
or U1874 (N_1874,In_502,In_691);
and U1875 (N_1875,In_302,In_329);
and U1876 (N_1876,In_682,In_217);
nand U1877 (N_1877,In_275,In_201);
nor U1878 (N_1878,In_87,In_243);
nor U1879 (N_1879,In_422,In_234);
nor U1880 (N_1880,In_609,In_308);
nand U1881 (N_1881,In_36,In_125);
nand U1882 (N_1882,In_704,In_339);
or U1883 (N_1883,In_247,In_328);
and U1884 (N_1884,In_18,In_351);
or U1885 (N_1885,In_667,In_353);
nor U1886 (N_1886,In_40,In_623);
or U1887 (N_1887,In_537,In_139);
and U1888 (N_1888,In_34,In_459);
and U1889 (N_1889,In_671,In_329);
and U1890 (N_1890,In_454,In_175);
nand U1891 (N_1891,In_396,In_691);
nor U1892 (N_1892,In_550,In_708);
nand U1893 (N_1893,In_35,In_720);
and U1894 (N_1894,In_595,In_179);
and U1895 (N_1895,In_292,In_654);
or U1896 (N_1896,In_671,In_467);
and U1897 (N_1897,In_463,In_164);
nand U1898 (N_1898,In_31,In_307);
nand U1899 (N_1899,In_500,In_375);
and U1900 (N_1900,In_63,In_112);
and U1901 (N_1901,In_543,In_102);
xor U1902 (N_1902,In_97,In_186);
or U1903 (N_1903,In_315,In_421);
or U1904 (N_1904,In_613,In_389);
and U1905 (N_1905,In_613,In_660);
nand U1906 (N_1906,In_426,In_99);
and U1907 (N_1907,In_134,In_550);
nor U1908 (N_1908,In_127,In_20);
xor U1909 (N_1909,In_93,In_90);
and U1910 (N_1910,In_696,In_559);
nor U1911 (N_1911,In_187,In_62);
and U1912 (N_1912,In_656,In_112);
nand U1913 (N_1913,In_610,In_183);
or U1914 (N_1914,In_714,In_348);
or U1915 (N_1915,In_113,In_698);
or U1916 (N_1916,In_220,In_43);
nor U1917 (N_1917,In_594,In_179);
nor U1918 (N_1918,In_682,In_354);
nand U1919 (N_1919,In_454,In_119);
and U1920 (N_1920,In_455,In_23);
nor U1921 (N_1921,In_608,In_702);
and U1922 (N_1922,In_449,In_596);
nand U1923 (N_1923,In_405,In_733);
or U1924 (N_1924,In_193,In_546);
and U1925 (N_1925,In_108,In_320);
and U1926 (N_1926,In_452,In_728);
and U1927 (N_1927,In_14,In_688);
nand U1928 (N_1928,In_190,In_699);
and U1929 (N_1929,In_748,In_711);
and U1930 (N_1930,In_746,In_601);
nand U1931 (N_1931,In_457,In_632);
nor U1932 (N_1932,In_694,In_142);
and U1933 (N_1933,In_539,In_126);
nand U1934 (N_1934,In_63,In_405);
nor U1935 (N_1935,In_7,In_325);
nand U1936 (N_1936,In_401,In_244);
nor U1937 (N_1937,In_465,In_153);
nor U1938 (N_1938,In_294,In_264);
nor U1939 (N_1939,In_535,In_564);
nor U1940 (N_1940,In_208,In_108);
nand U1941 (N_1941,In_188,In_422);
nand U1942 (N_1942,In_205,In_518);
or U1943 (N_1943,In_505,In_101);
and U1944 (N_1944,In_255,In_323);
nor U1945 (N_1945,In_464,In_288);
nand U1946 (N_1946,In_73,In_210);
nand U1947 (N_1947,In_40,In_241);
nor U1948 (N_1948,In_391,In_122);
or U1949 (N_1949,In_303,In_46);
or U1950 (N_1950,In_325,In_525);
or U1951 (N_1951,In_618,In_236);
or U1952 (N_1952,In_531,In_713);
nand U1953 (N_1953,In_572,In_268);
xnor U1954 (N_1954,In_197,In_89);
nor U1955 (N_1955,In_695,In_563);
nor U1956 (N_1956,In_160,In_428);
or U1957 (N_1957,In_295,In_345);
nand U1958 (N_1958,In_323,In_626);
or U1959 (N_1959,In_479,In_505);
and U1960 (N_1960,In_304,In_575);
xor U1961 (N_1961,In_688,In_58);
or U1962 (N_1962,In_278,In_287);
or U1963 (N_1963,In_59,In_172);
and U1964 (N_1964,In_71,In_302);
nand U1965 (N_1965,In_168,In_668);
or U1966 (N_1966,In_470,In_102);
or U1967 (N_1967,In_518,In_130);
nor U1968 (N_1968,In_576,In_353);
and U1969 (N_1969,In_129,In_552);
nand U1970 (N_1970,In_567,In_24);
and U1971 (N_1971,In_475,In_705);
or U1972 (N_1972,In_718,In_293);
nor U1973 (N_1973,In_459,In_175);
nand U1974 (N_1974,In_375,In_573);
and U1975 (N_1975,In_728,In_602);
nor U1976 (N_1976,In_551,In_285);
or U1977 (N_1977,In_731,In_106);
nand U1978 (N_1978,In_247,In_669);
nor U1979 (N_1979,In_615,In_491);
nand U1980 (N_1980,In_646,In_720);
nand U1981 (N_1981,In_78,In_562);
and U1982 (N_1982,In_271,In_679);
and U1983 (N_1983,In_191,In_639);
nor U1984 (N_1984,In_513,In_292);
or U1985 (N_1985,In_471,In_699);
nor U1986 (N_1986,In_669,In_546);
nor U1987 (N_1987,In_480,In_22);
or U1988 (N_1988,In_211,In_557);
or U1989 (N_1989,In_160,In_223);
nand U1990 (N_1990,In_221,In_676);
or U1991 (N_1991,In_191,In_736);
and U1992 (N_1992,In_99,In_688);
or U1993 (N_1993,In_230,In_645);
and U1994 (N_1994,In_310,In_222);
and U1995 (N_1995,In_60,In_126);
or U1996 (N_1996,In_21,In_585);
nor U1997 (N_1997,In_679,In_123);
nand U1998 (N_1998,In_209,In_162);
and U1999 (N_1999,In_66,In_110);
or U2000 (N_2000,In_280,In_730);
nor U2001 (N_2001,In_102,In_59);
and U2002 (N_2002,In_667,In_621);
nor U2003 (N_2003,In_133,In_230);
or U2004 (N_2004,In_678,In_427);
nor U2005 (N_2005,In_298,In_21);
or U2006 (N_2006,In_582,In_747);
nor U2007 (N_2007,In_552,In_347);
nand U2008 (N_2008,In_370,In_29);
nand U2009 (N_2009,In_683,In_745);
or U2010 (N_2010,In_697,In_464);
and U2011 (N_2011,In_443,In_514);
nor U2012 (N_2012,In_209,In_706);
and U2013 (N_2013,In_167,In_212);
nor U2014 (N_2014,In_141,In_183);
and U2015 (N_2015,In_423,In_710);
nor U2016 (N_2016,In_41,In_359);
nand U2017 (N_2017,In_745,In_153);
nor U2018 (N_2018,In_120,In_499);
or U2019 (N_2019,In_478,In_223);
and U2020 (N_2020,In_146,In_615);
or U2021 (N_2021,In_43,In_140);
nor U2022 (N_2022,In_508,In_61);
or U2023 (N_2023,In_199,In_363);
nand U2024 (N_2024,In_360,In_459);
nand U2025 (N_2025,In_176,In_277);
nor U2026 (N_2026,In_698,In_476);
or U2027 (N_2027,In_587,In_605);
and U2028 (N_2028,In_101,In_251);
and U2029 (N_2029,In_571,In_735);
xnor U2030 (N_2030,In_586,In_520);
nor U2031 (N_2031,In_555,In_482);
and U2032 (N_2032,In_609,In_687);
or U2033 (N_2033,In_113,In_575);
or U2034 (N_2034,In_636,In_482);
nor U2035 (N_2035,In_58,In_611);
nor U2036 (N_2036,In_599,In_528);
and U2037 (N_2037,In_434,In_619);
nand U2038 (N_2038,In_673,In_357);
or U2039 (N_2039,In_692,In_375);
and U2040 (N_2040,In_149,In_103);
or U2041 (N_2041,In_390,In_542);
nor U2042 (N_2042,In_188,In_384);
and U2043 (N_2043,In_214,In_95);
nand U2044 (N_2044,In_386,In_144);
nor U2045 (N_2045,In_591,In_454);
and U2046 (N_2046,In_622,In_216);
or U2047 (N_2047,In_544,In_417);
nand U2048 (N_2048,In_55,In_415);
nand U2049 (N_2049,In_687,In_512);
or U2050 (N_2050,In_688,In_545);
nand U2051 (N_2051,In_203,In_731);
nor U2052 (N_2052,In_275,In_117);
nor U2053 (N_2053,In_682,In_598);
nor U2054 (N_2054,In_628,In_619);
and U2055 (N_2055,In_311,In_502);
or U2056 (N_2056,In_244,In_442);
and U2057 (N_2057,In_115,In_712);
or U2058 (N_2058,In_649,In_201);
nand U2059 (N_2059,In_37,In_143);
or U2060 (N_2060,In_65,In_741);
nand U2061 (N_2061,In_81,In_653);
nand U2062 (N_2062,In_121,In_640);
nand U2063 (N_2063,In_465,In_712);
and U2064 (N_2064,In_564,In_692);
and U2065 (N_2065,In_700,In_76);
nor U2066 (N_2066,In_599,In_272);
or U2067 (N_2067,In_305,In_172);
or U2068 (N_2068,In_414,In_120);
xor U2069 (N_2069,In_578,In_481);
nand U2070 (N_2070,In_152,In_352);
or U2071 (N_2071,In_543,In_596);
or U2072 (N_2072,In_182,In_503);
or U2073 (N_2073,In_707,In_7);
and U2074 (N_2074,In_97,In_328);
or U2075 (N_2075,In_702,In_316);
and U2076 (N_2076,In_90,In_647);
nor U2077 (N_2077,In_2,In_510);
nor U2078 (N_2078,In_530,In_247);
and U2079 (N_2079,In_52,In_242);
nor U2080 (N_2080,In_604,In_139);
and U2081 (N_2081,In_319,In_126);
nor U2082 (N_2082,In_296,In_612);
nor U2083 (N_2083,In_206,In_613);
nor U2084 (N_2084,In_193,In_8);
or U2085 (N_2085,In_582,In_428);
nor U2086 (N_2086,In_590,In_238);
nor U2087 (N_2087,In_17,In_182);
nor U2088 (N_2088,In_275,In_640);
and U2089 (N_2089,In_685,In_533);
nor U2090 (N_2090,In_741,In_425);
nor U2091 (N_2091,In_46,In_10);
nand U2092 (N_2092,In_184,In_506);
and U2093 (N_2093,In_666,In_523);
or U2094 (N_2094,In_639,In_676);
and U2095 (N_2095,In_256,In_409);
nand U2096 (N_2096,In_76,In_709);
and U2097 (N_2097,In_392,In_239);
nor U2098 (N_2098,In_164,In_747);
nor U2099 (N_2099,In_142,In_629);
and U2100 (N_2100,In_581,In_444);
nand U2101 (N_2101,In_478,In_199);
nor U2102 (N_2102,In_607,In_601);
nor U2103 (N_2103,In_327,In_608);
nor U2104 (N_2104,In_454,In_316);
nor U2105 (N_2105,In_74,In_524);
or U2106 (N_2106,In_457,In_0);
nand U2107 (N_2107,In_703,In_102);
and U2108 (N_2108,In_349,In_46);
and U2109 (N_2109,In_16,In_579);
nor U2110 (N_2110,In_75,In_288);
and U2111 (N_2111,In_191,In_666);
xor U2112 (N_2112,In_565,In_574);
nand U2113 (N_2113,In_745,In_75);
and U2114 (N_2114,In_31,In_445);
and U2115 (N_2115,In_734,In_518);
nor U2116 (N_2116,In_237,In_10);
nor U2117 (N_2117,In_416,In_450);
or U2118 (N_2118,In_620,In_64);
or U2119 (N_2119,In_144,In_8);
nor U2120 (N_2120,In_247,In_197);
or U2121 (N_2121,In_390,In_30);
and U2122 (N_2122,In_341,In_248);
or U2123 (N_2123,In_282,In_71);
and U2124 (N_2124,In_466,In_236);
and U2125 (N_2125,In_76,In_216);
nand U2126 (N_2126,In_202,In_268);
nor U2127 (N_2127,In_325,In_663);
nor U2128 (N_2128,In_675,In_280);
nand U2129 (N_2129,In_147,In_534);
nor U2130 (N_2130,In_399,In_110);
nor U2131 (N_2131,In_169,In_1);
and U2132 (N_2132,In_68,In_57);
nand U2133 (N_2133,In_711,In_113);
or U2134 (N_2134,In_617,In_124);
or U2135 (N_2135,In_43,In_691);
or U2136 (N_2136,In_84,In_191);
nand U2137 (N_2137,In_21,In_725);
or U2138 (N_2138,In_570,In_84);
or U2139 (N_2139,In_717,In_683);
or U2140 (N_2140,In_535,In_693);
nand U2141 (N_2141,In_645,In_671);
nor U2142 (N_2142,In_481,In_593);
nor U2143 (N_2143,In_408,In_670);
nor U2144 (N_2144,In_91,In_386);
and U2145 (N_2145,In_12,In_575);
xor U2146 (N_2146,In_125,In_463);
nor U2147 (N_2147,In_155,In_255);
nor U2148 (N_2148,In_176,In_197);
and U2149 (N_2149,In_701,In_119);
nor U2150 (N_2150,In_499,In_690);
nor U2151 (N_2151,In_445,In_27);
or U2152 (N_2152,In_729,In_199);
or U2153 (N_2153,In_458,In_25);
and U2154 (N_2154,In_717,In_256);
and U2155 (N_2155,In_722,In_682);
xor U2156 (N_2156,In_51,In_128);
nand U2157 (N_2157,In_375,In_140);
or U2158 (N_2158,In_181,In_114);
nor U2159 (N_2159,In_603,In_120);
or U2160 (N_2160,In_729,In_675);
or U2161 (N_2161,In_66,In_331);
or U2162 (N_2162,In_308,In_517);
and U2163 (N_2163,In_221,In_88);
nor U2164 (N_2164,In_155,In_545);
and U2165 (N_2165,In_488,In_565);
nor U2166 (N_2166,In_2,In_485);
nand U2167 (N_2167,In_256,In_331);
or U2168 (N_2168,In_638,In_617);
nand U2169 (N_2169,In_424,In_287);
and U2170 (N_2170,In_408,In_611);
nor U2171 (N_2171,In_327,In_420);
and U2172 (N_2172,In_260,In_637);
nor U2173 (N_2173,In_190,In_346);
nand U2174 (N_2174,In_749,In_143);
nor U2175 (N_2175,In_590,In_483);
nand U2176 (N_2176,In_548,In_422);
and U2177 (N_2177,In_729,In_305);
nor U2178 (N_2178,In_388,In_471);
or U2179 (N_2179,In_485,In_555);
or U2180 (N_2180,In_480,In_688);
nor U2181 (N_2181,In_503,In_341);
or U2182 (N_2182,In_264,In_538);
and U2183 (N_2183,In_166,In_193);
nand U2184 (N_2184,In_516,In_80);
nor U2185 (N_2185,In_532,In_685);
xor U2186 (N_2186,In_32,In_184);
nor U2187 (N_2187,In_699,In_688);
xnor U2188 (N_2188,In_428,In_140);
nand U2189 (N_2189,In_745,In_213);
nor U2190 (N_2190,In_607,In_516);
or U2191 (N_2191,In_612,In_672);
nand U2192 (N_2192,In_342,In_38);
nand U2193 (N_2193,In_335,In_129);
nor U2194 (N_2194,In_508,In_723);
and U2195 (N_2195,In_195,In_145);
nor U2196 (N_2196,In_76,In_554);
nand U2197 (N_2197,In_262,In_733);
nand U2198 (N_2198,In_159,In_6);
nand U2199 (N_2199,In_399,In_59);
nand U2200 (N_2200,In_495,In_49);
or U2201 (N_2201,In_515,In_133);
nor U2202 (N_2202,In_687,In_190);
nand U2203 (N_2203,In_60,In_389);
xor U2204 (N_2204,In_237,In_554);
nand U2205 (N_2205,In_551,In_167);
or U2206 (N_2206,In_218,In_54);
or U2207 (N_2207,In_63,In_182);
and U2208 (N_2208,In_637,In_230);
nor U2209 (N_2209,In_60,In_202);
nor U2210 (N_2210,In_612,In_221);
xnor U2211 (N_2211,In_734,In_87);
nor U2212 (N_2212,In_309,In_677);
and U2213 (N_2213,In_547,In_207);
nand U2214 (N_2214,In_746,In_482);
and U2215 (N_2215,In_485,In_226);
nand U2216 (N_2216,In_431,In_628);
and U2217 (N_2217,In_511,In_644);
nand U2218 (N_2218,In_200,In_195);
and U2219 (N_2219,In_739,In_113);
nor U2220 (N_2220,In_187,In_208);
nand U2221 (N_2221,In_264,In_463);
nor U2222 (N_2222,In_337,In_102);
or U2223 (N_2223,In_455,In_216);
and U2224 (N_2224,In_127,In_506);
nand U2225 (N_2225,In_694,In_544);
or U2226 (N_2226,In_219,In_160);
nor U2227 (N_2227,In_411,In_38);
xnor U2228 (N_2228,In_225,In_524);
or U2229 (N_2229,In_39,In_491);
and U2230 (N_2230,In_116,In_107);
nor U2231 (N_2231,In_280,In_54);
nand U2232 (N_2232,In_531,In_93);
or U2233 (N_2233,In_707,In_297);
or U2234 (N_2234,In_286,In_152);
nor U2235 (N_2235,In_269,In_124);
or U2236 (N_2236,In_668,In_42);
nand U2237 (N_2237,In_280,In_191);
nand U2238 (N_2238,In_446,In_739);
xnor U2239 (N_2239,In_524,In_707);
or U2240 (N_2240,In_334,In_96);
or U2241 (N_2241,In_445,In_568);
nand U2242 (N_2242,In_267,In_220);
nand U2243 (N_2243,In_328,In_441);
nor U2244 (N_2244,In_368,In_223);
nor U2245 (N_2245,In_443,In_128);
nand U2246 (N_2246,In_315,In_48);
and U2247 (N_2247,In_578,In_409);
or U2248 (N_2248,In_117,In_720);
and U2249 (N_2249,In_461,In_606);
nor U2250 (N_2250,In_314,In_238);
nand U2251 (N_2251,In_169,In_196);
or U2252 (N_2252,In_133,In_716);
and U2253 (N_2253,In_698,In_699);
nor U2254 (N_2254,In_419,In_301);
and U2255 (N_2255,In_40,In_109);
nor U2256 (N_2256,In_528,In_718);
or U2257 (N_2257,In_533,In_341);
and U2258 (N_2258,In_746,In_121);
or U2259 (N_2259,In_749,In_265);
or U2260 (N_2260,In_187,In_527);
or U2261 (N_2261,In_222,In_434);
nand U2262 (N_2262,In_62,In_254);
nor U2263 (N_2263,In_158,In_53);
and U2264 (N_2264,In_727,In_88);
nand U2265 (N_2265,In_661,In_12);
nor U2266 (N_2266,In_740,In_234);
nand U2267 (N_2267,In_540,In_166);
nor U2268 (N_2268,In_242,In_412);
and U2269 (N_2269,In_188,In_351);
nand U2270 (N_2270,In_733,In_643);
nand U2271 (N_2271,In_180,In_571);
nor U2272 (N_2272,In_636,In_232);
and U2273 (N_2273,In_376,In_680);
nor U2274 (N_2274,In_470,In_435);
xnor U2275 (N_2275,In_422,In_400);
xor U2276 (N_2276,In_382,In_477);
or U2277 (N_2277,In_485,In_639);
and U2278 (N_2278,In_29,In_654);
nand U2279 (N_2279,In_637,In_138);
nor U2280 (N_2280,In_668,In_515);
or U2281 (N_2281,In_4,In_301);
and U2282 (N_2282,In_281,In_102);
nand U2283 (N_2283,In_670,In_463);
or U2284 (N_2284,In_177,In_573);
nor U2285 (N_2285,In_681,In_146);
and U2286 (N_2286,In_595,In_578);
and U2287 (N_2287,In_714,In_224);
or U2288 (N_2288,In_37,In_39);
or U2289 (N_2289,In_502,In_511);
nand U2290 (N_2290,In_522,In_628);
nand U2291 (N_2291,In_443,In_102);
nor U2292 (N_2292,In_588,In_438);
and U2293 (N_2293,In_90,In_406);
nor U2294 (N_2294,In_73,In_374);
or U2295 (N_2295,In_291,In_422);
or U2296 (N_2296,In_57,In_445);
nor U2297 (N_2297,In_18,In_73);
nand U2298 (N_2298,In_304,In_414);
and U2299 (N_2299,In_593,In_701);
nor U2300 (N_2300,In_664,In_394);
nand U2301 (N_2301,In_629,In_92);
or U2302 (N_2302,In_414,In_552);
nor U2303 (N_2303,In_711,In_242);
nor U2304 (N_2304,In_216,In_113);
and U2305 (N_2305,In_635,In_677);
and U2306 (N_2306,In_77,In_337);
or U2307 (N_2307,In_620,In_24);
nand U2308 (N_2308,In_468,In_383);
and U2309 (N_2309,In_549,In_394);
nor U2310 (N_2310,In_121,In_585);
or U2311 (N_2311,In_103,In_258);
nor U2312 (N_2312,In_713,In_534);
or U2313 (N_2313,In_331,In_238);
nor U2314 (N_2314,In_440,In_433);
nor U2315 (N_2315,In_460,In_481);
or U2316 (N_2316,In_639,In_710);
nor U2317 (N_2317,In_111,In_76);
nand U2318 (N_2318,In_572,In_653);
nand U2319 (N_2319,In_109,In_680);
nand U2320 (N_2320,In_389,In_735);
and U2321 (N_2321,In_485,In_667);
nor U2322 (N_2322,In_587,In_646);
and U2323 (N_2323,In_715,In_566);
nand U2324 (N_2324,In_402,In_338);
nor U2325 (N_2325,In_588,In_445);
and U2326 (N_2326,In_143,In_679);
nand U2327 (N_2327,In_91,In_631);
xor U2328 (N_2328,In_730,In_131);
nand U2329 (N_2329,In_16,In_644);
and U2330 (N_2330,In_27,In_535);
or U2331 (N_2331,In_344,In_411);
nand U2332 (N_2332,In_369,In_63);
and U2333 (N_2333,In_239,In_333);
or U2334 (N_2334,In_706,In_558);
nand U2335 (N_2335,In_715,In_748);
nor U2336 (N_2336,In_744,In_342);
nor U2337 (N_2337,In_277,In_61);
nor U2338 (N_2338,In_57,In_334);
and U2339 (N_2339,In_593,In_46);
and U2340 (N_2340,In_670,In_481);
nor U2341 (N_2341,In_668,In_537);
or U2342 (N_2342,In_273,In_472);
or U2343 (N_2343,In_23,In_557);
nand U2344 (N_2344,In_710,In_465);
xor U2345 (N_2345,In_309,In_0);
or U2346 (N_2346,In_387,In_559);
nor U2347 (N_2347,In_459,In_628);
or U2348 (N_2348,In_530,In_537);
or U2349 (N_2349,In_528,In_368);
or U2350 (N_2350,In_336,In_621);
and U2351 (N_2351,In_312,In_36);
nor U2352 (N_2352,In_207,In_522);
nor U2353 (N_2353,In_213,In_689);
and U2354 (N_2354,In_352,In_308);
and U2355 (N_2355,In_591,In_464);
or U2356 (N_2356,In_202,In_287);
nand U2357 (N_2357,In_643,In_9);
nor U2358 (N_2358,In_433,In_321);
nor U2359 (N_2359,In_38,In_348);
or U2360 (N_2360,In_482,In_269);
nor U2361 (N_2361,In_358,In_426);
and U2362 (N_2362,In_705,In_234);
nand U2363 (N_2363,In_407,In_739);
and U2364 (N_2364,In_374,In_259);
nand U2365 (N_2365,In_549,In_128);
or U2366 (N_2366,In_258,In_23);
or U2367 (N_2367,In_560,In_543);
nand U2368 (N_2368,In_519,In_408);
nor U2369 (N_2369,In_136,In_234);
and U2370 (N_2370,In_541,In_67);
and U2371 (N_2371,In_402,In_273);
or U2372 (N_2372,In_269,In_697);
nand U2373 (N_2373,In_410,In_558);
or U2374 (N_2374,In_576,In_593);
nand U2375 (N_2375,In_561,In_408);
nor U2376 (N_2376,In_246,In_343);
nand U2377 (N_2377,In_61,In_689);
nand U2378 (N_2378,In_38,In_519);
nand U2379 (N_2379,In_556,In_56);
nand U2380 (N_2380,In_385,In_349);
and U2381 (N_2381,In_609,In_379);
and U2382 (N_2382,In_162,In_128);
nand U2383 (N_2383,In_631,In_36);
nand U2384 (N_2384,In_533,In_671);
and U2385 (N_2385,In_251,In_139);
or U2386 (N_2386,In_419,In_415);
and U2387 (N_2387,In_356,In_650);
nor U2388 (N_2388,In_343,In_624);
or U2389 (N_2389,In_729,In_703);
nor U2390 (N_2390,In_566,In_173);
nor U2391 (N_2391,In_716,In_417);
or U2392 (N_2392,In_292,In_613);
nand U2393 (N_2393,In_396,In_127);
or U2394 (N_2394,In_599,In_397);
nor U2395 (N_2395,In_19,In_369);
and U2396 (N_2396,In_719,In_324);
and U2397 (N_2397,In_78,In_294);
nand U2398 (N_2398,In_427,In_152);
or U2399 (N_2399,In_744,In_84);
nor U2400 (N_2400,In_364,In_398);
and U2401 (N_2401,In_424,In_290);
and U2402 (N_2402,In_631,In_7);
or U2403 (N_2403,In_244,In_514);
nor U2404 (N_2404,In_579,In_195);
or U2405 (N_2405,In_518,In_726);
or U2406 (N_2406,In_130,In_211);
or U2407 (N_2407,In_542,In_88);
nand U2408 (N_2408,In_7,In_460);
nand U2409 (N_2409,In_164,In_507);
or U2410 (N_2410,In_148,In_465);
and U2411 (N_2411,In_276,In_596);
xnor U2412 (N_2412,In_10,In_470);
or U2413 (N_2413,In_706,In_493);
nand U2414 (N_2414,In_731,In_649);
nor U2415 (N_2415,In_436,In_280);
or U2416 (N_2416,In_622,In_653);
or U2417 (N_2417,In_74,In_447);
nor U2418 (N_2418,In_324,In_178);
nor U2419 (N_2419,In_275,In_370);
or U2420 (N_2420,In_262,In_189);
nor U2421 (N_2421,In_722,In_314);
xor U2422 (N_2422,In_411,In_590);
xnor U2423 (N_2423,In_723,In_680);
or U2424 (N_2424,In_129,In_364);
and U2425 (N_2425,In_675,In_130);
and U2426 (N_2426,In_711,In_103);
nor U2427 (N_2427,In_663,In_297);
and U2428 (N_2428,In_562,In_270);
or U2429 (N_2429,In_373,In_206);
nor U2430 (N_2430,In_310,In_677);
or U2431 (N_2431,In_367,In_59);
nand U2432 (N_2432,In_633,In_76);
and U2433 (N_2433,In_35,In_317);
nand U2434 (N_2434,In_172,In_348);
nor U2435 (N_2435,In_644,In_394);
nor U2436 (N_2436,In_261,In_173);
or U2437 (N_2437,In_583,In_79);
nor U2438 (N_2438,In_42,In_479);
nor U2439 (N_2439,In_480,In_726);
nor U2440 (N_2440,In_708,In_547);
or U2441 (N_2441,In_18,In_679);
nand U2442 (N_2442,In_253,In_495);
or U2443 (N_2443,In_40,In_320);
nor U2444 (N_2444,In_743,In_119);
or U2445 (N_2445,In_194,In_401);
nand U2446 (N_2446,In_652,In_322);
nor U2447 (N_2447,In_302,In_352);
and U2448 (N_2448,In_301,In_56);
nor U2449 (N_2449,In_686,In_730);
nand U2450 (N_2450,In_646,In_363);
nand U2451 (N_2451,In_178,In_625);
nor U2452 (N_2452,In_650,In_450);
or U2453 (N_2453,In_548,In_303);
or U2454 (N_2454,In_689,In_43);
nor U2455 (N_2455,In_522,In_209);
and U2456 (N_2456,In_741,In_499);
nor U2457 (N_2457,In_87,In_105);
nor U2458 (N_2458,In_298,In_409);
nor U2459 (N_2459,In_29,In_545);
or U2460 (N_2460,In_243,In_711);
nand U2461 (N_2461,In_396,In_742);
nor U2462 (N_2462,In_280,In_668);
and U2463 (N_2463,In_576,In_117);
xor U2464 (N_2464,In_717,In_504);
nor U2465 (N_2465,In_328,In_261);
or U2466 (N_2466,In_683,In_368);
or U2467 (N_2467,In_203,In_176);
or U2468 (N_2468,In_474,In_250);
or U2469 (N_2469,In_633,In_52);
nand U2470 (N_2470,In_395,In_663);
and U2471 (N_2471,In_384,In_376);
and U2472 (N_2472,In_377,In_415);
or U2473 (N_2473,In_673,In_728);
and U2474 (N_2474,In_663,In_377);
nand U2475 (N_2475,In_380,In_371);
or U2476 (N_2476,In_105,In_648);
or U2477 (N_2477,In_592,In_395);
or U2478 (N_2478,In_601,In_550);
or U2479 (N_2479,In_628,In_164);
or U2480 (N_2480,In_730,In_521);
or U2481 (N_2481,In_446,In_392);
nor U2482 (N_2482,In_381,In_539);
or U2483 (N_2483,In_183,In_357);
nand U2484 (N_2484,In_304,In_196);
nand U2485 (N_2485,In_511,In_708);
nor U2486 (N_2486,In_566,In_160);
nand U2487 (N_2487,In_721,In_188);
nor U2488 (N_2488,In_280,In_212);
or U2489 (N_2489,In_195,In_27);
nor U2490 (N_2490,In_264,In_23);
nand U2491 (N_2491,In_654,In_127);
nor U2492 (N_2492,In_183,In_616);
nand U2493 (N_2493,In_360,In_689);
or U2494 (N_2494,In_418,In_322);
and U2495 (N_2495,In_675,In_418);
nor U2496 (N_2496,In_339,In_638);
and U2497 (N_2497,In_458,In_150);
or U2498 (N_2498,In_647,In_295);
nor U2499 (N_2499,In_344,In_508);
or U2500 (N_2500,N_1808,N_2490);
nand U2501 (N_2501,N_1390,N_112);
nand U2502 (N_2502,N_898,N_1813);
nor U2503 (N_2503,N_1603,N_1129);
nand U2504 (N_2504,N_1733,N_1880);
nor U2505 (N_2505,N_251,N_1252);
nand U2506 (N_2506,N_2299,N_2326);
nand U2507 (N_2507,N_1137,N_178);
or U2508 (N_2508,N_1376,N_1158);
nand U2509 (N_2509,N_844,N_2209);
or U2510 (N_2510,N_1184,N_951);
and U2511 (N_2511,N_1094,N_1499);
nand U2512 (N_2512,N_1117,N_1998);
and U2513 (N_2513,N_297,N_1598);
nand U2514 (N_2514,N_2342,N_1367);
nand U2515 (N_2515,N_2460,N_1550);
nor U2516 (N_2516,N_2290,N_1220);
nor U2517 (N_2517,N_1820,N_509);
or U2518 (N_2518,N_516,N_293);
nor U2519 (N_2519,N_455,N_1156);
or U2520 (N_2520,N_893,N_481);
or U2521 (N_2521,N_1883,N_1860);
or U2522 (N_2522,N_860,N_2391);
nand U2523 (N_2523,N_244,N_1115);
nand U2524 (N_2524,N_687,N_171);
nor U2525 (N_2525,N_148,N_1047);
or U2526 (N_2526,N_1189,N_435);
nand U2527 (N_2527,N_595,N_1249);
or U2528 (N_2528,N_2124,N_2106);
and U2529 (N_2529,N_2385,N_2278);
nor U2530 (N_2530,N_1073,N_1964);
or U2531 (N_2531,N_1203,N_374);
nor U2532 (N_2532,N_2184,N_1728);
nand U2533 (N_2533,N_2113,N_1482);
or U2534 (N_2534,N_1887,N_1072);
or U2535 (N_2535,N_413,N_2314);
nor U2536 (N_2536,N_2218,N_1606);
or U2537 (N_2537,N_2330,N_1230);
and U2538 (N_2538,N_2028,N_895);
and U2539 (N_2539,N_240,N_544);
or U2540 (N_2540,N_700,N_1471);
nand U2541 (N_2541,N_1140,N_2424);
nand U2542 (N_2542,N_1186,N_404);
or U2543 (N_2543,N_51,N_1676);
and U2544 (N_2544,N_1922,N_1750);
and U2545 (N_2545,N_426,N_1875);
or U2546 (N_2546,N_368,N_1934);
nand U2547 (N_2547,N_241,N_470);
nor U2548 (N_2548,N_645,N_1768);
and U2549 (N_2549,N_680,N_1504);
nand U2550 (N_2550,N_1635,N_474);
nor U2551 (N_2551,N_2320,N_1191);
or U2552 (N_2552,N_2008,N_493);
or U2553 (N_2553,N_661,N_472);
nand U2554 (N_2554,N_1544,N_1175);
nor U2555 (N_2555,N_130,N_2307);
nand U2556 (N_2556,N_85,N_543);
or U2557 (N_2557,N_1508,N_2012);
nand U2558 (N_2558,N_405,N_217);
nor U2559 (N_2559,N_330,N_823);
or U2560 (N_2560,N_1561,N_408);
and U2561 (N_2561,N_2036,N_59);
and U2562 (N_2562,N_1283,N_2011);
or U2563 (N_2563,N_226,N_1358);
and U2564 (N_2564,N_1991,N_2402);
or U2565 (N_2565,N_335,N_1659);
or U2566 (N_2566,N_2009,N_2386);
nor U2567 (N_2567,N_1334,N_642);
nand U2568 (N_2568,N_2434,N_416);
nand U2569 (N_2569,N_2403,N_2436);
or U2570 (N_2570,N_400,N_826);
and U2571 (N_2571,N_41,N_228);
nand U2572 (N_2572,N_1004,N_314);
or U2573 (N_2573,N_104,N_1793);
nor U2574 (N_2574,N_1753,N_1003);
nand U2575 (N_2575,N_1285,N_526);
or U2576 (N_2576,N_1086,N_152);
or U2577 (N_2577,N_1802,N_1155);
and U2578 (N_2578,N_1861,N_98);
nor U2579 (N_2579,N_1268,N_1233);
and U2580 (N_2580,N_2020,N_879);
or U2581 (N_2581,N_1143,N_954);
xnor U2582 (N_2582,N_2381,N_74);
nand U2583 (N_2583,N_2498,N_2491);
or U2584 (N_2584,N_1,N_2241);
nor U2585 (N_2585,N_26,N_2423);
nor U2586 (N_2586,N_1325,N_1655);
and U2587 (N_2587,N_185,N_1902);
nand U2588 (N_2588,N_2282,N_1412);
and U2589 (N_2589,N_884,N_385);
or U2590 (N_2590,N_1899,N_2492);
nor U2591 (N_2591,N_1149,N_210);
nor U2592 (N_2592,N_2428,N_1159);
nand U2593 (N_2593,N_1862,N_1209);
nor U2594 (N_2594,N_1244,N_1965);
nand U2595 (N_2595,N_934,N_92);
nand U2596 (N_2596,N_2013,N_2056);
nor U2597 (N_2597,N_2194,N_2488);
or U2598 (N_2598,N_453,N_1890);
nor U2599 (N_2599,N_1792,N_615);
and U2600 (N_2600,N_2213,N_1667);
nor U2601 (N_2601,N_342,N_533);
nor U2602 (N_2602,N_624,N_1199);
nor U2603 (N_2603,N_960,N_237);
and U2604 (N_2604,N_1262,N_588);
nand U2605 (N_2605,N_425,N_1301);
or U2606 (N_2606,N_181,N_2067);
nor U2607 (N_2607,N_1596,N_935);
and U2608 (N_2608,N_1122,N_1788);
nor U2609 (N_2609,N_696,N_1421);
or U2610 (N_2610,N_360,N_729);
and U2611 (N_2611,N_1510,N_2172);
or U2612 (N_2612,N_773,N_1697);
nor U2613 (N_2613,N_465,N_636);
and U2614 (N_2614,N_1552,N_850);
or U2615 (N_2615,N_2211,N_1652);
nand U2616 (N_2616,N_880,N_1927);
or U2617 (N_2617,N_2446,N_311);
and U2618 (N_2618,N_1031,N_401);
or U2619 (N_2619,N_1312,N_2359);
nand U2620 (N_2620,N_1384,N_1282);
nand U2621 (N_2621,N_2471,N_587);
nand U2622 (N_2622,N_3,N_1270);
nor U2623 (N_2623,N_1258,N_2397);
and U2624 (N_2624,N_2458,N_565);
nor U2625 (N_2625,N_977,N_1123);
nor U2626 (N_2626,N_1810,N_1196);
nand U2627 (N_2627,N_1082,N_1898);
nor U2628 (N_2628,N_673,N_1629);
nand U2629 (N_2629,N_2162,N_2137);
nor U2630 (N_2630,N_136,N_859);
nand U2631 (N_2631,N_825,N_497);
or U2632 (N_2632,N_1636,N_2132);
nor U2633 (N_2633,N_398,N_1027);
and U2634 (N_2634,N_1352,N_1957);
and U2635 (N_2635,N_1326,N_1008);
and U2636 (N_2636,N_904,N_2064);
and U2637 (N_2637,N_103,N_788);
or U2638 (N_2638,N_2233,N_44);
nand U2639 (N_2639,N_306,N_2409);
and U2640 (N_2640,N_1055,N_123);
nand U2641 (N_2641,N_1167,N_1035);
nor U2642 (N_2642,N_1833,N_436);
or U2643 (N_2643,N_169,N_2293);
or U2644 (N_2644,N_348,N_2117);
nand U2645 (N_2645,N_276,N_1610);
and U2646 (N_2646,N_2268,N_35);
nor U2647 (N_2647,N_2096,N_215);
or U2648 (N_2648,N_1313,N_1058);
nand U2649 (N_2649,N_150,N_1618);
and U2650 (N_2650,N_1751,N_55);
nand U2651 (N_2651,N_381,N_781);
nor U2652 (N_2652,N_604,N_467);
and U2653 (N_2653,N_78,N_1328);
nand U2654 (N_2654,N_1870,N_1053);
nand U2655 (N_2655,N_2238,N_177);
and U2656 (N_2656,N_2379,N_2199);
or U2657 (N_2657,N_412,N_327);
nand U2658 (N_2658,N_849,N_957);
nand U2659 (N_2659,N_1542,N_1604);
and U2660 (N_2660,N_706,N_2392);
and U2661 (N_2661,N_568,N_1425);
nor U2662 (N_2662,N_2226,N_864);
or U2663 (N_2663,N_1400,N_203);
nor U2664 (N_2664,N_1147,N_2158);
and U2665 (N_2665,N_2154,N_1903);
or U2666 (N_2666,N_641,N_2485);
or U2667 (N_2667,N_1966,N_1744);
nor U2668 (N_2668,N_958,N_2244);
and U2669 (N_2669,N_429,N_2255);
nor U2670 (N_2670,N_175,N_1056);
nand U2671 (N_2671,N_596,N_569);
nor U2672 (N_2672,N_1840,N_767);
or U2673 (N_2673,N_170,N_2463);
and U2674 (N_2674,N_1713,N_2134);
or U2675 (N_2675,N_2388,N_144);
nand U2676 (N_2676,N_608,N_1615);
or U2677 (N_2677,N_1319,N_1578);
nand U2678 (N_2678,N_548,N_252);
nor U2679 (N_2679,N_963,N_40);
nand U2680 (N_2680,N_2181,N_1928);
xnor U2681 (N_2681,N_1772,N_189);
nand U2682 (N_2682,N_444,N_1799);
and U2683 (N_2683,N_1944,N_1557);
nand U2684 (N_2684,N_329,N_1483);
and U2685 (N_2685,N_683,N_1626);
nand U2686 (N_2686,N_558,N_86);
nor U2687 (N_2687,N_2075,N_1148);
and U2688 (N_2688,N_1969,N_776);
or U2689 (N_2689,N_2177,N_198);
and U2690 (N_2690,N_1917,N_892);
or U2691 (N_2691,N_733,N_281);
nor U2692 (N_2692,N_503,N_2489);
or U2693 (N_2693,N_1476,N_100);
or U2694 (N_2694,N_1242,N_1719);
nand U2695 (N_2695,N_920,N_2029);
nand U2696 (N_2696,N_2195,N_1625);
or U2697 (N_2697,N_452,N_654);
or U2698 (N_2698,N_1670,N_67);
nand U2699 (N_2699,N_585,N_220);
and U2700 (N_2700,N_1439,N_578);
and U2701 (N_2701,N_1468,N_667);
and U2702 (N_2702,N_1278,N_1386);
or U2703 (N_2703,N_1422,N_1487);
nor U2704 (N_2704,N_261,N_876);
or U2705 (N_2705,N_1079,N_1113);
nand U2706 (N_2706,N_862,N_291);
nor U2707 (N_2707,N_1748,N_1878);
nor U2708 (N_2708,N_1216,N_31);
and U2709 (N_2709,N_1593,N_354);
nor U2710 (N_2710,N_1681,N_295);
and U2711 (N_2711,N_1896,N_1017);
nor U2712 (N_2712,N_468,N_2322);
nand U2713 (N_2713,N_469,N_1206);
nand U2714 (N_2714,N_2419,N_1423);
nand U2715 (N_2715,N_2149,N_1275);
or U2716 (N_2716,N_106,N_117);
and U2717 (N_2717,N_1682,N_1491);
and U2718 (N_2718,N_2193,N_1018);
and U2719 (N_2719,N_82,N_54);
and U2720 (N_2720,N_1740,N_511);
nand U2721 (N_2721,N_151,N_820);
and U2722 (N_2722,N_1030,N_411);
or U2723 (N_2723,N_437,N_1663);
nand U2724 (N_2724,N_2478,N_1540);
or U2725 (N_2725,N_1770,N_1782);
and U2726 (N_2726,N_1284,N_1228);
or U2727 (N_2727,N_1281,N_222);
nor U2728 (N_2728,N_658,N_1107);
and U2729 (N_2729,N_1801,N_504);
nand U2730 (N_2730,N_2310,N_2201);
and U2731 (N_2731,N_406,N_141);
and U2732 (N_2732,N_1163,N_1752);
and U2733 (N_2733,N_1503,N_403);
and U2734 (N_2734,N_1872,N_1842);
xor U2735 (N_2735,N_1293,N_1646);
nand U2736 (N_2736,N_529,N_1064);
or U2737 (N_2737,N_1683,N_2237);
or U2738 (N_2738,N_1885,N_1198);
or U2739 (N_2739,N_813,N_268);
and U2740 (N_2740,N_882,N_1469);
xnor U2741 (N_2741,N_1797,N_1498);
nand U2742 (N_2742,N_671,N_379);
nand U2743 (N_2743,N_1513,N_1102);
nand U2744 (N_2744,N_1823,N_208);
or U2745 (N_2745,N_1597,N_583);
nor U2746 (N_2746,N_2225,N_1316);
or U2747 (N_2747,N_1536,N_2119);
or U2748 (N_2748,N_640,N_1357);
and U2749 (N_2749,N_1583,N_2470);
nor U2750 (N_2750,N_372,N_149);
nor U2751 (N_2751,N_168,N_1600);
or U2752 (N_2752,N_1723,N_118);
nand U2753 (N_2753,N_264,N_1088);
and U2754 (N_2754,N_32,N_931);
and U2755 (N_2755,N_37,N_541);
or U2756 (N_2756,N_1116,N_2331);
nand U2757 (N_2757,N_1466,N_1034);
nor U2758 (N_2758,N_1224,N_902);
nor U2759 (N_2759,N_2465,N_1179);
nand U2760 (N_2760,N_745,N_2219);
nand U2761 (N_2761,N_2484,N_1131);
and U2762 (N_2762,N_775,N_2239);
or U2763 (N_2763,N_557,N_430);
or U2764 (N_2764,N_2450,N_146);
xor U2765 (N_2765,N_1006,N_322);
nor U2766 (N_2766,N_972,N_1895);
nand U2767 (N_2767,N_774,N_24);
and U2768 (N_2768,N_1634,N_964);
nand U2769 (N_2769,N_1338,N_1307);
nor U2770 (N_2770,N_839,N_111);
nor U2771 (N_2771,N_952,N_351);
nor U2772 (N_2772,N_637,N_1559);
and U2773 (N_2773,N_1257,N_1581);
and U2774 (N_2774,N_2001,N_1255);
nand U2775 (N_2775,N_2155,N_1647);
nor U2776 (N_2776,N_1311,N_1584);
nand U2777 (N_2777,N_871,N_2315);
or U2778 (N_2778,N_319,N_2110);
nand U2779 (N_2779,N_552,N_1401);
nand U2780 (N_2780,N_532,N_1521);
and U2781 (N_2781,N_2130,N_1190);
or U2782 (N_2782,N_865,N_1771);
and U2783 (N_2783,N_2196,N_2205);
or U2784 (N_2784,N_60,N_807);
or U2785 (N_2785,N_1945,N_866);
or U2786 (N_2786,N_912,N_1248);
nor U2787 (N_2787,N_2269,N_681);
nand U2788 (N_2788,N_205,N_1722);
and U2789 (N_2789,N_1675,N_383);
nor U2790 (N_2790,N_182,N_1574);
nand U2791 (N_2791,N_2325,N_1101);
or U2792 (N_2792,N_517,N_101);
and U2793 (N_2793,N_1570,N_2439);
nor U2794 (N_2794,N_685,N_1791);
nand U2795 (N_2795,N_914,N_2412);
and U2796 (N_2796,N_108,N_975);
nor U2797 (N_2797,N_2191,N_423);
and U2798 (N_2798,N_1280,N_1543);
xnor U2799 (N_2799,N_1648,N_861);
nor U2800 (N_2800,N_2174,N_919);
nor U2801 (N_2801,N_2369,N_2311);
or U2802 (N_2802,N_2267,N_1114);
nor U2803 (N_2803,N_200,N_2222);
nand U2804 (N_2804,N_736,N_1843);
xor U2805 (N_2805,N_2298,N_2408);
nor U2806 (N_2806,N_1141,N_1051);
and U2807 (N_2807,N_1560,N_138);
nand U2808 (N_2808,N_2058,N_921);
or U2809 (N_2809,N_1958,N_2127);
and U2810 (N_2810,N_784,N_1548);
or U2811 (N_2811,N_1208,N_764);
or U2812 (N_2812,N_1726,N_1711);
nor U2813 (N_2813,N_1746,N_2279);
nor U2814 (N_2814,N_326,N_345);
and U2815 (N_2815,N_325,N_2277);
or U2816 (N_2816,N_932,N_1492);
and U2817 (N_2817,N_827,N_1452);
nand U2818 (N_2818,N_973,N_1707);
or U2819 (N_2819,N_1500,N_900);
and U2820 (N_2820,N_2276,N_1721);
and U2821 (N_2821,N_1020,N_821);
and U2822 (N_2822,N_87,N_277);
or U2823 (N_2823,N_1085,N_757);
or U2824 (N_2824,N_1142,N_2050);
nor U2825 (N_2825,N_959,N_576);
nor U2826 (N_2826,N_1005,N_1622);
and U2827 (N_2827,N_431,N_1680);
nor U2828 (N_2828,N_1028,N_2285);
xnor U2829 (N_2829,N_2236,N_1865);
or U2830 (N_2830,N_531,N_1049);
or U2831 (N_2831,N_2247,N_589);
and U2832 (N_2832,N_1549,N_1154);
nand U2833 (N_2833,N_908,N_1343);
nor U2834 (N_2834,N_289,N_1590);
nor U2835 (N_2835,N_323,N_1764);
nand U2836 (N_2836,N_950,N_2281);
nor U2837 (N_2837,N_581,N_1481);
xnor U2838 (N_2838,N_2227,N_2494);
nand U2839 (N_2839,N_365,N_16);
and U2840 (N_2840,N_2171,N_2179);
or U2841 (N_2841,N_2347,N_2387);
or U2842 (N_2842,N_600,N_1730);
or U2843 (N_2843,N_896,N_993);
nand U2844 (N_2844,N_214,N_2121);
nand U2845 (N_2845,N_1591,N_689);
or U2846 (N_2846,N_835,N_193);
or U2847 (N_2847,N_843,N_650);
and U2848 (N_2848,N_507,N_1857);
or U2849 (N_2849,N_1377,N_1294);
nor U2850 (N_2850,N_1514,N_1260);
nor U2851 (N_2851,N_447,N_129);
nand U2852 (N_2852,N_157,N_211);
and U2853 (N_2853,N_1767,N_131);
nor U2854 (N_2854,N_1745,N_2057);
and U2855 (N_2855,N_2414,N_513);
or U2856 (N_2856,N_786,N_282);
and U2857 (N_2857,N_936,N_611);
and U2858 (N_2858,N_2431,N_1331);
or U2859 (N_2859,N_2437,N_153);
and U2860 (N_2860,N_925,N_724);
nand U2861 (N_2861,N_1525,N_274);
or U2862 (N_2862,N_1608,N_1786);
and U2863 (N_2863,N_1558,N_2461);
nand U2864 (N_2864,N_755,N_2467);
nand U2865 (N_2865,N_2382,N_1332);
and U2866 (N_2866,N_328,N_612);
nor U2867 (N_2867,N_852,N_313);
and U2868 (N_2868,N_2457,N_1506);
or U2869 (N_2869,N_2187,N_2002);
or U2870 (N_2870,N_1656,N_1990);
nor U2871 (N_2871,N_347,N_2445);
nor U2872 (N_2872,N_2348,N_2416);
nor U2873 (N_2873,N_2144,N_1187);
nor U2874 (N_2874,N_1348,N_249);
nand U2875 (N_2875,N_2356,N_1994);
nor U2876 (N_2876,N_2432,N_2280);
and U2877 (N_2877,N_2480,N_842);
and U2878 (N_2878,N_207,N_1973);
nor U2879 (N_2879,N_2366,N_1716);
nor U2880 (N_2880,N_28,N_1126);
nor U2881 (N_2881,N_2077,N_1534);
or U2882 (N_2882,N_454,N_397);
nand U2883 (N_2883,N_180,N_165);
nand U2884 (N_2884,N_1518,N_593);
or U2885 (N_2885,N_858,N_362);
or U2886 (N_2886,N_1961,N_473);
nand U2887 (N_2887,N_2059,N_2295);
or U2888 (N_2888,N_2455,N_2232);
or U2889 (N_2889,N_1404,N_723);
nor U2890 (N_2890,N_549,N_783);
and U2891 (N_2891,N_1546,N_29);
and U2892 (N_2892,N_2027,N_1065);
or U2893 (N_2893,N_1405,N_392);
and U2894 (N_2894,N_1237,N_1761);
nand U2895 (N_2895,N_2313,N_1967);
nor U2896 (N_2896,N_2350,N_948);
nand U2897 (N_2897,N_540,N_2486);
nand U2898 (N_2898,N_747,N_794);
nand U2899 (N_2899,N_955,N_2005);
nor U2900 (N_2900,N_1677,N_370);
and U2901 (N_2901,N_885,N_731);
and U2902 (N_2902,N_1435,N_1850);
nand U2903 (N_2903,N_324,N_1916);
or U2904 (N_2904,N_805,N_1355);
nor U2905 (N_2905,N_653,N_1327);
or U2906 (N_2906,N_57,N_1956);
and U2907 (N_2907,N_45,N_1061);
nor U2908 (N_2908,N_907,N_2100);
or U2909 (N_2909,N_1599,N_646);
or U2910 (N_2910,N_535,N_889);
or U2911 (N_2911,N_793,N_828);
and U2912 (N_2912,N_66,N_366);
or U2913 (N_2913,N_2087,N_1605);
or U2914 (N_2914,N_2118,N_1133);
nand U2915 (N_2915,N_357,N_1099);
nor U2916 (N_2916,N_1951,N_2259);
nand U2917 (N_2917,N_769,N_915);
nor U2918 (N_2918,N_937,N_377);
nor U2919 (N_2919,N_1125,N_1866);
xor U2920 (N_2920,N_1620,N_1756);
nor U2921 (N_2921,N_2234,N_1617);
or U2922 (N_2922,N_2321,N_2139);
and U2923 (N_2923,N_2010,N_2499);
nor U2924 (N_2924,N_1059,N_1938);
nor U2925 (N_2925,N_1960,N_812);
or U2926 (N_2926,N_1690,N_488);
or U2927 (N_2927,N_2192,N_720);
nor U2928 (N_2928,N_979,N_1876);
nand U2929 (N_2929,N_305,N_1953);
or U2930 (N_2930,N_1774,N_176);
nand U2931 (N_2931,N_187,N_1795);
nor U2932 (N_2932,N_554,N_448);
and U2933 (N_2933,N_737,N_1024);
and U2934 (N_2934,N_1264,N_881);
or U2935 (N_2935,N_1735,N_142);
nand U2936 (N_2936,N_143,N_2405);
or U2937 (N_2937,N_2039,N_2204);
nor U2938 (N_2938,N_1614,N_1362);
nor U2939 (N_2939,N_1434,N_1124);
nor U2940 (N_2940,N_966,N_2327);
nor U2941 (N_2941,N_1385,N_262);
and U2942 (N_2942,N_2301,N_128);
nor U2943 (N_2943,N_1022,N_590);
nand U2944 (N_2944,N_2346,N_47);
or U2945 (N_2945,N_1339,N_566);
nand U2946 (N_2946,N_20,N_579);
and U2947 (N_2947,N_216,N_838);
xnor U2948 (N_2948,N_1829,N_816);
or U2949 (N_2949,N_1909,N_651);
nand U2950 (N_2950,N_953,N_1528);
and U2951 (N_2951,N_1105,N_353);
or U2952 (N_2952,N_1170,N_2074);
nand U2953 (N_2953,N_1830,N_1729);
or U2954 (N_2954,N_1908,N_1449);
or U2955 (N_2955,N_371,N_522);
nand U2956 (N_2956,N_1408,N_439);
nor U2957 (N_2957,N_2245,N_1463);
or U2958 (N_2958,N_728,N_363);
or U2959 (N_2959,N_1344,N_308);
nand U2960 (N_2960,N_1251,N_1212);
and U2961 (N_2961,N_1804,N_1461);
nor U2962 (N_2962,N_2426,N_2150);
or U2963 (N_2963,N_2340,N_854);
nor U2964 (N_2964,N_797,N_2368);
nand U2965 (N_2965,N_2069,N_771);
and U2966 (N_2966,N_2034,N_484);
nor U2967 (N_2967,N_1462,N_1845);
or U2968 (N_2968,N_1023,N_334);
xnor U2969 (N_2969,N_722,N_1999);
or U2970 (N_2970,N_1373,N_1040);
nand U2971 (N_2971,N_1522,N_584);
or U2972 (N_2972,N_2168,N_1305);
nor U2973 (N_2973,N_461,N_1446);
or U2974 (N_2974,N_88,N_545);
and U2975 (N_2975,N_1480,N_1662);
or U2976 (N_2976,N_1076,N_318);
nor U2977 (N_2977,N_2185,N_2324);
or U2978 (N_2978,N_1341,N_2060);
or U2979 (N_2979,N_894,N_657);
or U2980 (N_2980,N_1259,N_1858);
nor U2981 (N_2981,N_1638,N_2125);
and U2982 (N_2982,N_1145,N_462);
nor U2983 (N_2983,N_1985,N_833);
nor U2984 (N_2984,N_647,N_458);
nor U2985 (N_2985,N_1692,N_1315);
or U2986 (N_2986,N_450,N_2042);
and U2987 (N_2987,N_1200,N_753);
nand U2988 (N_2988,N_1688,N_1743);
nand U2989 (N_2989,N_930,N_2082);
or U2990 (N_2990,N_2252,N_494);
or U2991 (N_2991,N_750,N_996);
or U2992 (N_2992,N_1241,N_2076);
nor U2993 (N_2993,N_34,N_903);
nor U2994 (N_2994,N_536,N_410);
and U2995 (N_2995,N_1180,N_1393);
nor U2996 (N_2996,N_631,N_1340);
or U2997 (N_2997,N_2109,N_2);
nor U2998 (N_2998,N_460,N_2377);
or U2999 (N_2999,N_350,N_223);
and U3000 (N_3000,N_284,N_2122);
or U3001 (N_3001,N_830,N_1151);
or U3002 (N_3002,N_25,N_804);
or U3003 (N_3003,N_2248,N_2120);
nand U3004 (N_3004,N_1366,N_2270);
nor U3005 (N_3005,N_445,N_2367);
nor U3006 (N_3006,N_974,N_2230);
nor U3007 (N_3007,N_154,N_906);
and U3008 (N_3008,N_1042,N_675);
and U3009 (N_3009,N_1486,N_570);
or U3010 (N_3010,N_46,N_758);
and U3011 (N_3011,N_1738,N_1855);
nand U3012 (N_3012,N_1849,N_2371);
or U3013 (N_3013,N_1083,N_275);
nor U3014 (N_3014,N_1353,N_2095);
and U3015 (N_3015,N_341,N_1387);
nor U3016 (N_3016,N_2145,N_1112);
or U3017 (N_3017,N_1821,N_1399);
nor U3018 (N_3018,N_1074,N_709);
nor U3019 (N_3019,N_2294,N_2173);
or U3020 (N_3020,N_2357,N_1856);
and U3021 (N_3021,N_1223,N_2464);
and U3022 (N_3022,N_891,N_346);
xnor U3023 (N_3023,N_2440,N_1637);
and U3024 (N_3024,N_1213,N_1271);
or U3025 (N_3025,N_814,N_785);
or U3026 (N_3026,N_1426,N_2286);
nor U3027 (N_3027,N_521,N_2469);
nor U3028 (N_3028,N_1739,N_1523);
xor U3029 (N_3029,N_527,N_1696);
and U3030 (N_3030,N_2396,N_195);
and U3031 (N_3031,N_1437,N_482);
and U3032 (N_3032,N_2355,N_1930);
and U3033 (N_3033,N_440,N_1070);
nor U3034 (N_3034,N_33,N_1886);
or U3035 (N_3035,N_79,N_1417);
and U3036 (N_3036,N_997,N_2098);
and U3037 (N_3037,N_1464,N_0);
nor U3038 (N_3038,N_267,N_2215);
nor U3039 (N_3039,N_1096,N_989);
nand U3040 (N_3040,N_1502,N_1243);
and U3041 (N_3041,N_1227,N_751);
or U3042 (N_3042,N_2115,N_421);
nand U3043 (N_3043,N_1274,N_2182);
and U3044 (N_3044,N_2049,N_2415);
and U3045 (N_3045,N_1925,N_212);
and U3046 (N_3046,N_1624,N_1779);
nand U3047 (N_3047,N_2062,N_114);
or U3048 (N_3048,N_1451,N_1572);
or U3049 (N_3049,N_1568,N_1816);
or U3050 (N_3050,N_2136,N_2107);
nand U3051 (N_3051,N_422,N_1672);
nand U3052 (N_3052,N_434,N_1477);
nor U3053 (N_3053,N_299,N_616);
nand U3054 (N_3054,N_69,N_1937);
and U3055 (N_3055,N_1882,N_2148);
or U3056 (N_3056,N_715,N_1585);
nand U3057 (N_3057,N_983,N_1374);
and U3058 (N_3058,N_6,N_22);
nor U3059 (N_3059,N_1941,N_1848);
nor U3060 (N_3060,N_1645,N_1569);
and U3061 (N_3061,N_23,N_464);
nand U3062 (N_3062,N_245,N_840);
and U3063 (N_3063,N_1780,N_234);
and U3064 (N_3064,N_2335,N_480);
or U3065 (N_3065,N_302,N_1695);
and U3066 (N_3066,N_1447,N_1397);
and U3067 (N_3067,N_1798,N_1381);
xor U3068 (N_3068,N_2103,N_878);
or U3069 (N_3069,N_2143,N_2170);
nand U3070 (N_3070,N_847,N_1277);
or U3071 (N_3071,N_601,N_2417);
and U3072 (N_3072,N_132,N_155);
nor U3073 (N_3073,N_1438,N_286);
or U3074 (N_3074,N_1587,N_725);
or U3075 (N_3075,N_1710,N_1512);
nor U3076 (N_3076,N_831,N_515);
and U3077 (N_3077,N_162,N_1673);
nor U3078 (N_3078,N_1913,N_1556);
nor U3079 (N_3079,N_1914,N_1108);
nand U3080 (N_3080,N_792,N_486);
nor U3081 (N_3081,N_2114,N_992);
and U3082 (N_3082,N_373,N_1098);
and U3083 (N_3083,N_2015,N_1347);
nand U3084 (N_3084,N_1715,N_272);
nor U3085 (N_3085,N_417,N_610);
and U3086 (N_3086,N_2214,N_752);
and U3087 (N_3087,N_1734,N_2479);
nor U3088 (N_3088,N_853,N_339);
and U3089 (N_3089,N_320,N_1225);
nor U3090 (N_3090,N_2061,N_1160);
nor U3091 (N_3091,N_1253,N_2105);
and U3092 (N_3092,N_1100,N_599);
or U3093 (N_3093,N_2456,N_125);
and U3094 (N_3094,N_710,N_2296);
nand U3095 (N_3095,N_12,N_2048);
nor U3096 (N_3096,N_1554,N_1863);
and U3097 (N_3097,N_1787,N_121);
nor U3098 (N_3098,N_534,N_1853);
nor U3099 (N_3099,N_1702,N_508);
nor U3100 (N_3100,N_183,N_968);
nor U3101 (N_3101,N_1837,N_1000);
nand U3102 (N_3102,N_2070,N_2216);
or U3103 (N_3103,N_2260,N_2261);
and U3104 (N_3104,N_1193,N_564);
nand U3105 (N_3105,N_218,N_609);
nand U3106 (N_3106,N_161,N_846);
and U3107 (N_3107,N_2338,N_2256);
and U3108 (N_3108,N_2086,N_2474);
and U3109 (N_3109,N_1644,N_707);
nand U3110 (N_3110,N_1963,N_1416);
nor U3111 (N_3111,N_1666,N_1911);
or U3112 (N_3112,N_711,N_1947);
nor U3113 (N_3113,N_815,N_1807);
or U3114 (N_3114,N_1317,N_759);
or U3115 (N_3115,N_873,N_206);
nand U3116 (N_3116,N_61,N_2341);
nand U3117 (N_3117,N_1380,N_537);
nand U3118 (N_3118,N_841,N_338);
nor U3119 (N_3119,N_304,N_998);
or U3120 (N_3120,N_1057,N_1345);
or U3121 (N_3121,N_102,N_15);
and U3122 (N_3122,N_575,N_1246);
and U3123 (N_3123,N_1877,N_1081);
nand U3124 (N_3124,N_1276,N_1411);
nor U3125 (N_3125,N_867,N_1302);
or U3126 (N_3126,N_1250,N_666);
nand U3127 (N_3127,N_1714,N_238);
nor U3128 (N_3128,N_1939,N_2041);
and U3129 (N_3129,N_648,N_1157);
or U3130 (N_3130,N_2309,N_1153);
and U3131 (N_3131,N_1701,N_1161);
and U3132 (N_3132,N_686,N_2482);
and U3133 (N_3133,N_2175,N_1515);
nor U3134 (N_3134,N_2206,N_1952);
or U3135 (N_3135,N_2370,N_1631);
nor U3136 (N_3136,N_883,N_99);
and U3137 (N_3137,N_1643,N_1395);
nor U3138 (N_3138,N_2000,N_1651);
and U3139 (N_3139,N_414,N_697);
and U3140 (N_3140,N_787,N_1201);
nor U3141 (N_3141,N_1704,N_2344);
nor U3142 (N_3142,N_188,N_2052);
nor U3143 (N_3143,N_1488,N_1448);
nand U3144 (N_3144,N_2242,N_56);
nor U3145 (N_3145,N_1781,N_940);
and U3146 (N_3146,N_1440,N_1363);
nand U3147 (N_3147,N_2129,N_186);
and U3148 (N_3148,N_8,N_510);
nor U3149 (N_3149,N_2487,N_122);
or U3150 (N_3150,N_762,N_574);
nor U3151 (N_3151,N_1940,N_560);
nor U3152 (N_3152,N_1444,N_789);
nand U3153 (N_3153,N_75,N_137);
nand U3154 (N_3154,N_1467,N_2349);
nand U3155 (N_3155,N_1359,N_296);
or U3156 (N_3156,N_765,N_1509);
nor U3157 (N_3157,N_1612,N_2262);
and U3158 (N_3158,N_1299,N_1234);
and U3159 (N_3159,N_115,N_2065);
nand U3160 (N_3160,N_1906,N_1864);
nand U3161 (N_3161,N_984,N_2004);
nor U3162 (N_3162,N_2334,N_2413);
and U3163 (N_3163,N_818,N_888);
or U3164 (N_3164,N_2221,N_778);
nor U3165 (N_3165,N_1517,N_27);
nor U3166 (N_3166,N_676,N_479);
and U3167 (N_3167,N_1755,N_1674);
nor U3168 (N_3168,N_1531,N_1516);
nand U3169 (N_3169,N_1778,N_2452);
nor U3170 (N_3170,N_1306,N_438);
nand U3171 (N_3171,N_982,N_824);
or U3172 (N_3172,N_2164,N_1240);
and U3173 (N_3173,N_1904,N_1485);
and U3174 (N_3174,N_2147,N_2046);
and U3175 (N_3175,N_1535,N_1595);
nor U3176 (N_3176,N_1982,N_2240);
nand U3177 (N_3177,N_1263,N_1080);
nand U3178 (N_3178,N_556,N_1144);
nor U3179 (N_3179,N_396,N_364);
nand U3180 (N_3180,N_242,N_639);
nand U3181 (N_3181,N_991,N_1641);
and U3182 (N_3182,N_1974,N_1171);
nor U3183 (N_3183,N_2085,N_1060);
nand U3184 (N_3184,N_2207,N_1127);
and U3185 (N_3185,N_1538,N_550);
and U3186 (N_3186,N_1458,N_717);
and U3187 (N_3187,N_1784,N_985);
or U3188 (N_3188,N_1297,N_2273);
nand U3189 (N_3189,N_555,N_395);
nor U3190 (N_3190,N_2291,N_714);
nor U3191 (N_3191,N_1992,N_970);
or U3192 (N_3192,N_2343,N_690);
nor U3193 (N_3193,N_1501,N_2017);
and U3194 (N_3194,N_1633,N_2319);
or U3195 (N_3195,N_1091,N_419);
nand U3196 (N_3196,N_2312,N_1507);
nor U3197 (N_3197,N_2102,N_1565);
nand U3198 (N_3198,N_2229,N_2475);
nor U3199 (N_3199,N_1943,N_1759);
nor U3200 (N_3200,N_1011,N_1836);
nand U3201 (N_3201,N_127,N_1640);
or U3202 (N_3202,N_2123,N_68);
nor U3203 (N_3203,N_664,N_1443);
or U3204 (N_3204,N_1290,N_1727);
and U3205 (N_3205,N_1825,N_1827);
and U3206 (N_3206,N_1287,N_18);
and U3207 (N_3207,N_2352,N_1616);
and U3208 (N_3208,N_2258,N_163);
and U3209 (N_3209,N_1970,N_336);
nand U3210 (N_3210,N_754,N_204);
nand U3211 (N_3211,N_1869,N_120);
and U3212 (N_3212,N_113,N_743);
nand U3213 (N_3213,N_1314,N_278);
and U3214 (N_3214,N_1669,N_246);
or U3215 (N_3215,N_1146,N_42);
nand U3216 (N_3216,N_909,N_271);
or U3217 (N_3217,N_303,N_2272);
nor U3218 (N_3218,N_1236,N_1188);
and U3219 (N_3219,N_1564,N_1218);
and U3220 (N_3220,N_2031,N_1001);
or U3221 (N_3221,N_525,N_808);
and U3222 (N_3222,N_1229,N_505);
nor U3223 (N_3223,N_459,N_580);
nor U3224 (N_3224,N_1136,N_803);
or U3225 (N_3225,N_744,N_1490);
or U3226 (N_3226,N_947,N_1594);
nand U3227 (N_3227,N_1354,N_1176);
nor U3228 (N_3228,N_806,N_868);
nand U3229 (N_3229,N_1817,N_1497);
nand U3230 (N_3230,N_698,N_309);
or U3231 (N_3231,N_1984,N_1718);
nand U3232 (N_3232,N_1068,N_2176);
or U3233 (N_3233,N_1298,N_810);
nand U3234 (N_3234,N_2235,N_1361);
and U3235 (N_3235,N_708,N_1699);
and U3236 (N_3236,N_1474,N_905);
nor U3237 (N_3237,N_1602,N_2200);
nand U3238 (N_3238,N_1232,N_1613);
or U3239 (N_3239,N_1424,N_746);
or U3240 (N_3240,N_2003,N_1292);
nand U3241 (N_3241,N_2043,N_735);
nor U3242 (N_3242,N_748,N_2166);
nand U3243 (N_3243,N_2410,N_1494);
nor U3244 (N_3244,N_1418,N_2339);
or U3245 (N_3245,N_1420,N_2038);
or U3246 (N_3246,N_443,N_2165);
nor U3247 (N_3247,N_1981,N_1368);
and U3248 (N_3248,N_1879,N_1962);
nand U3249 (N_3249,N_1472,N_1762);
and U3250 (N_3250,N_1320,N_1433);
and U3251 (N_3251,N_196,N_1679);
or U3252 (N_3252,N_298,N_1664);
and U3253 (N_3253,N_923,N_799);
nor U3254 (N_3254,N_2406,N_1336);
and U3255 (N_3255,N_321,N_2019);
or U3256 (N_3256,N_192,N_2302);
or U3257 (N_3257,N_1077,N_2398);
nor U3258 (N_3258,N_1709,N_260);
and U3259 (N_3259,N_1095,N_1295);
and U3260 (N_3260,N_1231,N_614);
nor U3261 (N_3261,N_201,N_739);
or U3262 (N_3262,N_756,N_1582);
nand U3263 (N_3263,N_19,N_2351);
or U3264 (N_3264,N_1470,N_1431);
or U3265 (N_3265,N_768,N_378);
nor U3266 (N_3266,N_1834,N_1211);
and U3267 (N_3267,N_1010,N_1846);
nand U3268 (N_3268,N_918,N_2284);
and U3269 (N_3269,N_795,N_1609);
or U3270 (N_3270,N_80,N_2444);
nand U3271 (N_3271,N_1724,N_64);
nand U3272 (N_3272,N_1712,N_1084);
nor U3273 (N_3273,N_688,N_1689);
and U3274 (N_3274,N_1693,N_811);
nor U3275 (N_3275,N_2047,N_1364);
or U3276 (N_3276,N_602,N_1265);
and U3277 (N_3277,N_367,N_2153);
and U3278 (N_3278,N_2097,N_184);
or U3279 (N_3279,N_834,N_1279);
and U3280 (N_3280,N_310,N_1529);
and U3281 (N_3281,N_1226,N_1021);
and U3282 (N_3282,N_36,N_231);
nand U3283 (N_3283,N_391,N_279);
nand U3284 (N_3284,N_420,N_1104);
or U3285 (N_3285,N_1217,N_967);
and U3286 (N_3286,N_1983,N_916);
nand U3287 (N_3287,N_2289,N_941);
or U3288 (N_3288,N_386,N_933);
nand U3289 (N_3289,N_1950,N_1811);
nand U3290 (N_3290,N_927,N_179);
and U3291 (N_3291,N_1409,N_135);
nand U3292 (N_3292,N_1794,N_1071);
nor U3293 (N_3293,N_2390,N_1731);
and U3294 (N_3294,N_1378,N_1684);
nand U3295 (N_3295,N_2429,N_1777);
nand U3296 (N_3296,N_1575,N_2014);
nor U3297 (N_3297,N_1168,N_2303);
and U3298 (N_3298,N_53,N_4);
and U3299 (N_3299,N_1221,N_1454);
or U3300 (N_3300,N_1009,N_2271);
or U3301 (N_3301,N_292,N_1205);
and U3302 (N_3302,N_1867,N_1658);
nand U3303 (N_3303,N_1757,N_618);
and U3304 (N_3304,N_332,N_1592);
or U3305 (N_3305,N_1029,N_48);
and U3306 (N_3306,N_1563,N_1106);
or U3307 (N_3307,N_1933,N_2411);
or U3308 (N_3308,N_2140,N_331);
and U3309 (N_3309,N_358,N_692);
nand U3310 (N_3310,N_490,N_2198);
or U3311 (N_3311,N_2323,N_1455);
and U3312 (N_3312,N_2212,N_1815);
or U3313 (N_3313,N_1720,N_1222);
nand U3314 (N_3314,N_911,N_2138);
and U3315 (N_3315,N_598,N_1033);
nor U3316 (N_3316,N_1166,N_230);
nand U3317 (N_3317,N_2283,N_1014);
and U3318 (N_3318,N_1379,N_2045);
or U3319 (N_3319,N_1993,N_999);
nand U3320 (N_3320,N_542,N_961);
or U3321 (N_3321,N_2180,N_1526);
nor U3322 (N_3322,N_1356,N_670);
nor U3323 (N_3323,N_1632,N_2449);
nor U3324 (N_3324,N_1407,N_90);
nor U3325 (N_3325,N_855,N_1954);
and U3326 (N_3326,N_553,N_2468);
or U3327 (N_3327,N_2068,N_1267);
and U3328 (N_3328,N_2151,N_1800);
nor U3329 (N_3329,N_1121,N_628);
nand U3330 (N_3330,N_2090,N_1016);
nor U3331 (N_3331,N_1323,N_1370);
and U3332 (N_3332,N_2133,N_2089);
nand U3333 (N_3333,N_1032,N_1892);
or U3334 (N_3334,N_1959,N_2372);
nor U3335 (N_3335,N_730,N_2223);
nor U3336 (N_3336,N_390,N_2266);
or U3337 (N_3337,N_1457,N_2418);
nand U3338 (N_3338,N_1551,N_716);
or U3339 (N_3339,N_1747,N_50);
nand U3340 (N_3340,N_477,N_343);
or U3341 (N_3341,N_194,N_14);
or U3342 (N_3342,N_976,N_623);
nand U3343 (N_3343,N_2399,N_938);
nor U3344 (N_3344,N_38,N_1576);
or U3345 (N_3345,N_990,N_1553);
and U3346 (N_3346,N_83,N_1182);
nand U3347 (N_3347,N_344,N_1803);
and U3348 (N_3348,N_1375,N_283);
or U3349 (N_3349,N_1002,N_2496);
or U3350 (N_3350,N_2477,N_402);
nand U3351 (N_3351,N_761,N_1588);
nor U3352 (N_3352,N_1247,N_969);
nor U3353 (N_3353,N_1132,N_432);
or U3354 (N_3354,N_2257,N_2016);
nor U3355 (N_3355,N_1383,N_2454);
and U3356 (N_3356,N_704,N_1537);
or U3357 (N_3357,N_2425,N_1912);
nor U3358 (N_3358,N_1988,N_669);
and U3359 (N_3359,N_290,N_1173);
nor U3360 (N_3360,N_2353,N_1854);
or U3361 (N_3361,N_1918,N_1841);
and U3362 (N_3362,N_2030,N_446);
and U3363 (N_3363,N_2092,N_73);
and U3364 (N_3364,N_1177,N_1495);
nand U3365 (N_3365,N_790,N_1350);
or U3366 (N_3366,N_269,N_1814);
and U3367 (N_3367,N_134,N_2394);
nor U3368 (N_3368,N_980,N_617);
nor U3369 (N_3369,N_52,N_682);
or U3370 (N_3370,N_1219,N_1705);
nand U3371 (N_3371,N_502,N_2251);
nand U3372 (N_3372,N_956,N_1150);
and U3373 (N_3373,N_506,N_2430);
nand U3374 (N_3374,N_1195,N_546);
or U3375 (N_3375,N_219,N_1272);
nor U3376 (N_3376,N_2023,N_9);
nand U3377 (N_3377,N_2112,N_457);
nor U3378 (N_3378,N_1562,N_2407);
nand U3379 (N_3379,N_2384,N_1183);
or U3380 (N_3380,N_819,N_1844);
nand U3381 (N_3381,N_1162,N_1948);
or U3382 (N_3382,N_1742,N_780);
nand U3383 (N_3383,N_1202,N_699);
nand U3384 (N_3384,N_524,N_1619);
or U3385 (N_3385,N_2263,N_1093);
nor U3386 (N_3386,N_2389,N_1050);
nor U3387 (N_3387,N_1092,N_300);
or U3388 (N_3388,N_562,N_1296);
nor U3389 (N_3389,N_1831,N_2099);
nor U3390 (N_3390,N_591,N_2264);
nor U3391 (N_3391,N_857,N_738);
nor U3392 (N_3392,N_140,N_1324);
nand U3393 (N_3393,N_656,N_2421);
nor U3394 (N_3394,N_632,N_5);
nor U3395 (N_3395,N_663,N_167);
nand U3396 (N_3396,N_1322,N_2345);
nand U3397 (N_3397,N_1478,N_199);
nand U3398 (N_3398,N_856,N_1089);
and U3399 (N_3399,N_213,N_13);
nor U3400 (N_3400,N_929,N_483);
nand U3401 (N_3401,N_2497,N_1822);
nor U3402 (N_3402,N_713,N_2094);
nand U3403 (N_3403,N_1979,N_428);
nand U3404 (N_3404,N_2156,N_1181);
or U3405 (N_3405,N_1884,N_1445);
or U3406 (N_3406,N_2072,N_285);
nor U3407 (N_3407,N_433,N_870);
nand U3408 (N_3408,N_1300,N_2274);
nand U3409 (N_3409,N_1429,N_2078);
and U3410 (N_3410,N_124,N_848);
or U3411 (N_3411,N_1754,N_1138);
nor U3412 (N_3412,N_586,N_1577);
nor U3413 (N_3413,N_1796,N_897);
nor U3414 (N_3414,N_2108,N_1996);
and U3415 (N_3415,N_312,N_1627);
nor U3416 (N_3416,N_110,N_81);
nand U3417 (N_3417,N_126,N_561);
nor U3418 (N_3418,N_874,N_678);
and U3419 (N_3419,N_1062,N_2231);
nor U3420 (N_3420,N_197,N_1660);
or U3421 (N_3421,N_97,N_913);
nand U3422 (N_3422,N_1571,N_1410);
or U3423 (N_3423,N_2018,N_559);
or U3424 (N_3424,N_2364,N_1891);
or U3425 (N_3425,N_2063,N_2079);
and U3426 (N_3426,N_978,N_2401);
and U3427 (N_3427,N_145,N_1046);
or U3428 (N_3428,N_2373,N_802);
nor U3429 (N_3429,N_1955,N_1308);
nand U3430 (N_3430,N_399,N_2126);
nand U3431 (N_3431,N_1977,N_962);
nand U3432 (N_3432,N_1043,N_1269);
nor U3433 (N_3433,N_107,N_2336);
or U3434 (N_3434,N_1763,N_2022);
or U3435 (N_3435,N_2188,N_1976);
and U3436 (N_3436,N_471,N_236);
and U3437 (N_3437,N_2202,N_1567);
and U3438 (N_3438,N_84,N_2427);
nand U3439 (N_3439,N_1520,N_718);
and U3440 (N_3440,N_1036,N_1194);
nor U3441 (N_3441,N_2318,N_2161);
nor U3442 (N_3442,N_734,N_890);
nor U3443 (N_3443,N_2035,N_1266);
nor U3444 (N_3444,N_1414,N_1694);
nor U3445 (N_3445,N_1809,N_2083);
nor U3446 (N_3446,N_732,N_1760);
nor U3447 (N_3447,N_1769,N_315);
nor U3448 (N_3448,N_721,N_94);
nor U3449 (N_3449,N_530,N_89);
nand U3450 (N_3450,N_1790,N_741);
nand U3451 (N_3451,N_1178,N_160);
and U3452 (N_3452,N_605,N_777);
or U3453 (N_3453,N_1832,N_1919);
and U3454 (N_3454,N_265,N_622);
nand U3455 (N_3455,N_626,N_705);
and U3456 (N_3456,N_2328,N_945);
or U3457 (N_3457,N_491,N_375);
and U3458 (N_3458,N_1090,N_1881);
or U3459 (N_3459,N_2084,N_1496);
nand U3460 (N_3460,N_1717,N_1621);
and U3461 (N_3461,N_1475,N_356);
nand U3462 (N_3462,N_971,N_1893);
nor U3463 (N_3463,N_2378,N_1453);
nand U3464 (N_3464,N_2250,N_944);
and U3465 (N_3465,N_551,N_1128);
or U3466 (N_3466,N_1396,N_2395);
nor U3467 (N_3467,N_424,N_567);
or U3468 (N_3468,N_1130,N_779);
xnor U3469 (N_3469,N_164,N_409);
nor U3470 (N_3470,N_1054,N_2217);
nand U3471 (N_3471,N_924,N_1894);
nand U3472 (N_3472,N_703,N_760);
or U3473 (N_3473,N_1725,N_2111);
or U3474 (N_3474,N_202,N_1533);
nor U3475 (N_3475,N_2249,N_832);
and U3476 (N_3476,N_1351,N_597);
nor U3477 (N_3477,N_1812,N_58);
nor U3478 (N_3478,N_2288,N_243);
nor U3479 (N_3479,N_662,N_1589);
or U3480 (N_3480,N_2466,N_1256);
nand U3481 (N_3481,N_994,N_1924);
and U3482 (N_3482,N_369,N_1649);
or U3483 (N_3483,N_498,N_1045);
and U3484 (N_3484,N_1736,N_1566);
nor U3485 (N_3485,N_2160,N_229);
nor U3486 (N_3486,N_2131,N_2186);
and U3487 (N_3487,N_2448,N_1749);
nor U3488 (N_3488,N_2443,N_875);
nand U3489 (N_3489,N_1766,N_672);
nand U3490 (N_3490,N_2157,N_2383);
and U3491 (N_3491,N_394,N_1484);
nand U3492 (N_3492,N_147,N_1936);
and U3493 (N_3493,N_2462,N_701);
nor U3494 (N_3494,N_2007,N_809);
or U3495 (N_3495,N_2093,N_1532);
and U3496 (N_3496,N_987,N_910);
nand U3497 (N_3497,N_1687,N_2375);
or U3498 (N_3498,N_280,N_288);
nor U3499 (N_3499,N_489,N_2040);
nand U3500 (N_3500,N_1685,N_63);
or U3501 (N_3501,N_442,N_1403);
and U3502 (N_3502,N_1839,N_539);
and U3503 (N_3503,N_2146,N_2178);
and U3504 (N_3504,N_287,N_1369);
xnor U3505 (N_3505,N_2024,N_49);
nor U3506 (N_3506,N_1360,N_2292);
and U3507 (N_3507,N_1286,N_1773);
nand U3508 (N_3508,N_119,N_939);
or U3509 (N_3509,N_478,N_643);
and U3510 (N_3510,N_965,N_1910);
nand U3511 (N_3511,N_1479,N_1432);
nand U3512 (N_3512,N_523,N_2365);
and U3513 (N_3513,N_1980,N_1665);
or U3514 (N_3514,N_301,N_317);
or U3515 (N_3515,N_886,N_512);
nand U3516 (N_3516,N_235,N_684);
nor U3517 (N_3517,N_800,N_869);
nand U3518 (N_3518,N_2053,N_1968);
nand U3519 (N_3519,N_926,N_415);
or U3520 (N_3520,N_1776,N_1921);
nor U3521 (N_3521,N_1402,N_829);
nand U3522 (N_3522,N_1489,N_1580);
nand U3523 (N_3523,N_547,N_2404);
or U3524 (N_3524,N_1835,N_652);
nand U3525 (N_3525,N_492,N_1078);
nand U3526 (N_3526,N_1737,N_665);
and U3527 (N_3527,N_1111,N_1579);
xor U3528 (N_3528,N_2329,N_1819);
nand U3529 (N_3529,N_340,N_2476);
and U3530 (N_3530,N_772,N_239);
nand U3531 (N_3531,N_726,N_133);
and U3532 (N_3532,N_2208,N_257);
nand U3533 (N_3533,N_1932,N_352);
and U3534 (N_3534,N_899,N_2101);
nand U3535 (N_3535,N_1349,N_763);
nand U3536 (N_3536,N_1365,N_1019);
nor U3537 (N_3537,N_943,N_2453);
nand U3538 (N_3538,N_1436,N_791);
or U3539 (N_3539,N_1037,N_782);
nor U3540 (N_3540,N_2438,N_456);
nor U3541 (N_3541,N_11,N_487);
nand U3542 (N_3542,N_1110,N_1775);
and U3543 (N_3543,N_2073,N_227);
and U3544 (N_3544,N_427,N_2442);
nand U3545 (N_3545,N_1995,N_837);
nand U3546 (N_3546,N_1852,N_466);
and U3547 (N_3547,N_2493,N_1859);
and U3548 (N_3548,N_248,N_538);
nand U3549 (N_3549,N_270,N_712);
nor U3550 (N_3550,N_693,N_191);
and U3551 (N_3551,N_1291,N_2362);
nand U3552 (N_3552,N_649,N_1907);
and U3553 (N_3553,N_2159,N_2305);
nor U3554 (N_3554,N_259,N_355);
nand U3555 (N_3555,N_1828,N_1428);
and U3556 (N_3556,N_1245,N_817);
nand U3557 (N_3557,N_96,N_501);
nand U3558 (N_3558,N_1686,N_917);
nor U3559 (N_3559,N_1118,N_70);
and U3560 (N_3560,N_1653,N_1935);
and U3561 (N_3561,N_1505,N_1639);
nand U3562 (N_3562,N_451,N_2287);
nor U3563 (N_3563,N_1989,N_1038);
and U3564 (N_3564,N_1668,N_2358);
or U3565 (N_3565,N_1459,N_294);
or U3566 (N_3566,N_316,N_232);
xnor U3567 (N_3567,N_1333,N_380);
nor U3568 (N_3568,N_1971,N_2435);
nand U3569 (N_3569,N_224,N_1289);
and U3570 (N_3570,N_1765,N_1923);
nand U3571 (N_3571,N_93,N_1703);
nand U3572 (N_3572,N_1321,N_1586);
nand U3573 (N_3573,N_2091,N_607);
xnor U3574 (N_3574,N_2055,N_1330);
nor U3575 (N_3575,N_1210,N_1103);
nor U3576 (N_3576,N_1547,N_1607);
nor U3577 (N_3577,N_1337,N_1235);
and U3578 (N_3578,N_877,N_109);
nand U3579 (N_3579,N_1450,N_500);
or U3580 (N_3580,N_2374,N_159);
and U3581 (N_3581,N_1041,N_1657);
nand U3582 (N_3582,N_1273,N_863);
and U3583 (N_3583,N_2363,N_887);
and U3584 (N_3584,N_72,N_2275);
or U3585 (N_3585,N_1398,N_627);
or U3586 (N_3586,N_1389,N_679);
and U3587 (N_3587,N_1700,N_2297);
and U3588 (N_3588,N_2224,N_225);
nor U3589 (N_3589,N_266,N_2243);
nand U3590 (N_3590,N_1382,N_2006);
or U3591 (N_3591,N_603,N_1698);
nor U3592 (N_3592,N_384,N_621);
or U3593 (N_3593,N_77,N_476);
or U3594 (N_3594,N_2081,N_1539);
and U3595 (N_3595,N_17,N_1897);
nor U3596 (N_3596,N_633,N_2308);
or U3597 (N_3597,N_2400,N_221);
nor U3598 (N_3598,N_349,N_1007);
and U3599 (N_3599,N_988,N_946);
xor U3600 (N_3600,N_2183,N_2152);
and U3601 (N_3601,N_796,N_2354);
or U3602 (N_3602,N_393,N_2253);
and U3603 (N_3603,N_1406,N_337);
nand U3604 (N_3604,N_634,N_2473);
and U3605 (N_3605,N_1915,N_1427);
or U3606 (N_3606,N_1025,N_1623);
nand U3607 (N_3607,N_2337,N_845);
xor U3608 (N_3608,N_39,N_635);
and U3609 (N_3609,N_1678,N_475);
nand U3610 (N_3610,N_1650,N_1473);
or U3611 (N_3611,N_2265,N_2246);
and U3612 (N_3612,N_2447,N_1039);
nor U3613 (N_3613,N_677,N_2361);
and U3614 (N_3614,N_2197,N_1671);
nand U3615 (N_3615,N_1601,N_981);
nand U3616 (N_3616,N_668,N_1871);
and U3617 (N_3617,N_1239,N_674);
nand U3618 (N_3618,N_1630,N_1204);
or U3619 (N_3619,N_21,N_256);
nor U3620 (N_3620,N_1192,N_255);
nand U3621 (N_3621,N_172,N_2422);
and U3622 (N_3622,N_1888,N_2433);
nor U3623 (N_3623,N_2104,N_1134);
nor U3624 (N_3624,N_1785,N_62);
nor U3625 (N_3625,N_441,N_1942);
nor U3626 (N_3626,N_1874,N_2306);
and U3627 (N_3627,N_836,N_2167);
and U3628 (N_3628,N_166,N_659);
nor U3629 (N_3629,N_333,N_2254);
nor U3630 (N_3630,N_2332,N_1119);
nand U3631 (N_3631,N_95,N_1708);
nor U3632 (N_3632,N_1152,N_495);
and U3633 (N_3633,N_1905,N_520);
nor U3634 (N_3634,N_1066,N_1493);
nand U3635 (N_3635,N_1304,N_1826);
nor U3636 (N_3636,N_901,N_749);
and U3637 (N_3637,N_2472,N_2054);
nor U3638 (N_3638,N_1847,N_2483);
and U3639 (N_3639,N_801,N_2203);
nor U3640 (N_3640,N_770,N_1628);
nand U3641 (N_3641,N_209,N_190);
nor U3642 (N_3642,N_2021,N_2441);
nor U3643 (N_3643,N_2189,N_1335);
nor U3644 (N_3644,N_1303,N_250);
nor U3645 (N_3645,N_2495,N_644);
nand U3646 (N_3646,N_872,N_2300);
nand U3647 (N_3647,N_116,N_105);
nand U3648 (N_3648,N_2190,N_1026);
nor U3649 (N_3649,N_449,N_1164);
and U3650 (N_3650,N_518,N_1456);
or U3651 (N_3651,N_2304,N_254);
or U3652 (N_3652,N_30,N_1013);
nand U3653 (N_3653,N_359,N_407);
nor U3654 (N_3654,N_1430,N_2459);
or U3655 (N_3655,N_1931,N_1783);
nand U3656 (N_3656,N_1371,N_1067);
and U3657 (N_3657,N_2169,N_2317);
nand U3658 (N_3658,N_1207,N_1465);
nor U3659 (N_3659,N_1511,N_1261);
nand U3660 (N_3660,N_156,N_1214);
or U3661 (N_3661,N_1109,N_1169);
or U3662 (N_3662,N_630,N_519);
nor U3663 (N_3663,N_233,N_928);
or U3664 (N_3664,N_1135,N_1611);
and U3665 (N_3665,N_10,N_1758);
nand U3666 (N_3666,N_577,N_2163);
and U3667 (N_3667,N_1015,N_2026);
nor U3668 (N_3668,N_620,N_2066);
or U3669 (N_3669,N_1838,N_694);
and U3670 (N_3670,N_2051,N_91);
nor U3671 (N_3671,N_71,N_43);
or U3672 (N_3672,N_1441,N_1318);
and U3673 (N_3673,N_1732,N_258);
nand U3674 (N_3674,N_619,N_1949);
and U3675 (N_3675,N_1063,N_1069);
or U3676 (N_3676,N_1997,N_740);
xnor U3677 (N_3677,N_387,N_139);
and U3678 (N_3678,N_563,N_2032);
or U3679 (N_3679,N_1873,N_1920);
xnor U3680 (N_3680,N_1139,N_307);
nor U3681 (N_3681,N_1097,N_1372);
or U3682 (N_3682,N_2080,N_1900);
or U3683 (N_3683,N_1197,N_2025);
and U3684 (N_3684,N_2376,N_174);
or U3685 (N_3685,N_1254,N_1288);
xor U3686 (N_3686,N_1824,N_1818);
or U3687 (N_3687,N_606,N_1987);
nand U3688 (N_3688,N_65,N_2116);
nor U3689 (N_3689,N_2380,N_695);
nand U3690 (N_3690,N_1889,N_1545);
and U3691 (N_3691,N_613,N_625);
and U3692 (N_3692,N_1165,N_2451);
and U3693 (N_3693,N_1442,N_1975);
and U3694 (N_3694,N_727,N_2393);
nand U3695 (N_3695,N_1215,N_361);
nand U3696 (N_3696,N_1413,N_1391);
nand U3697 (N_3697,N_1419,N_418);
nor U3698 (N_3698,N_382,N_273);
or U3699 (N_3699,N_1901,N_1048);
and U3700 (N_3700,N_592,N_496);
nor U3701 (N_3701,N_2044,N_1120);
and U3702 (N_3702,N_719,N_1741);
or U3703 (N_3703,N_76,N_949);
nor U3704 (N_3704,N_263,N_1868);
xor U3705 (N_3705,N_1805,N_822);
or U3706 (N_3706,N_1946,N_986);
and U3707 (N_3707,N_2316,N_1174);
or U3708 (N_3708,N_376,N_1415);
or U3709 (N_3709,N_691,N_485);
nor U3710 (N_3710,N_1530,N_388);
or U3711 (N_3711,N_1394,N_1654);
nor U3712 (N_3712,N_573,N_1642);
or U3713 (N_3713,N_2210,N_1392);
nand U3714 (N_3714,N_1044,N_1806);
and U3715 (N_3715,N_1789,N_1460);
nor U3716 (N_3716,N_1310,N_655);
nand U3717 (N_3717,N_942,N_629);
nand U3718 (N_3718,N_1986,N_514);
and U3719 (N_3719,N_247,N_1075);
nor U3720 (N_3720,N_1978,N_1388);
and U3721 (N_3721,N_1926,N_1519);
and U3722 (N_3722,N_2360,N_1052);
nand U3723 (N_3723,N_1329,N_2033);
and U3724 (N_3724,N_742,N_2220);
nor U3725 (N_3725,N_2071,N_7);
or U3726 (N_3726,N_528,N_571);
or U3727 (N_3727,N_1238,N_1691);
nand U3728 (N_3728,N_1555,N_1573);
nand U3729 (N_3729,N_1309,N_253);
nand U3730 (N_3730,N_2088,N_463);
nand U3731 (N_3731,N_1342,N_389);
nor U3732 (N_3732,N_851,N_594);
nor U3733 (N_3733,N_2037,N_922);
xor U3734 (N_3734,N_582,N_2228);
nor U3735 (N_3735,N_1706,N_660);
nor U3736 (N_3736,N_2481,N_2135);
nand U3737 (N_3737,N_1087,N_572);
and U3738 (N_3738,N_2142,N_2141);
or U3739 (N_3739,N_1524,N_158);
and U3740 (N_3740,N_1541,N_702);
or U3741 (N_3741,N_173,N_499);
nor U3742 (N_3742,N_995,N_766);
or U3743 (N_3743,N_1185,N_2333);
and U3744 (N_3744,N_1972,N_798);
and U3745 (N_3745,N_1929,N_2128);
nand U3746 (N_3746,N_638,N_1527);
or U3747 (N_3747,N_1851,N_1346);
nand U3748 (N_3748,N_1012,N_2420);
and U3749 (N_3749,N_1661,N_1172);
and U3750 (N_3750,N_679,N_114);
nand U3751 (N_3751,N_2234,N_2173);
nand U3752 (N_3752,N_624,N_1225);
nand U3753 (N_3753,N_1579,N_448);
or U3754 (N_3754,N_1702,N_1534);
nor U3755 (N_3755,N_1982,N_2277);
nor U3756 (N_3756,N_2381,N_1651);
nand U3757 (N_3757,N_2115,N_1454);
nor U3758 (N_3758,N_1005,N_662);
nand U3759 (N_3759,N_2113,N_1469);
nor U3760 (N_3760,N_992,N_368);
or U3761 (N_3761,N_1256,N_1720);
nand U3762 (N_3762,N_919,N_123);
and U3763 (N_3763,N_1745,N_1270);
and U3764 (N_3764,N_228,N_2268);
and U3765 (N_3765,N_1773,N_1203);
and U3766 (N_3766,N_1210,N_2314);
and U3767 (N_3767,N_670,N_2296);
or U3768 (N_3768,N_39,N_828);
and U3769 (N_3769,N_429,N_1982);
nor U3770 (N_3770,N_18,N_2443);
or U3771 (N_3771,N_191,N_305);
nor U3772 (N_3772,N_2076,N_1123);
or U3773 (N_3773,N_1132,N_2220);
and U3774 (N_3774,N_1822,N_1007);
or U3775 (N_3775,N_670,N_1936);
and U3776 (N_3776,N_970,N_210);
and U3777 (N_3777,N_360,N_1333);
nor U3778 (N_3778,N_2376,N_1740);
nor U3779 (N_3779,N_2018,N_1286);
or U3780 (N_3780,N_1495,N_2038);
or U3781 (N_3781,N_1014,N_1124);
and U3782 (N_3782,N_2498,N_1063);
or U3783 (N_3783,N_756,N_1298);
and U3784 (N_3784,N_2096,N_2460);
nand U3785 (N_3785,N_19,N_1661);
or U3786 (N_3786,N_1118,N_304);
nand U3787 (N_3787,N_1374,N_681);
and U3788 (N_3788,N_732,N_482);
nand U3789 (N_3789,N_347,N_41);
nand U3790 (N_3790,N_596,N_645);
or U3791 (N_3791,N_2309,N_548);
nand U3792 (N_3792,N_1450,N_29);
nor U3793 (N_3793,N_1443,N_1051);
or U3794 (N_3794,N_694,N_1910);
and U3795 (N_3795,N_1816,N_1144);
or U3796 (N_3796,N_1501,N_177);
nand U3797 (N_3797,N_2088,N_1842);
and U3798 (N_3798,N_2186,N_1620);
nand U3799 (N_3799,N_0,N_1740);
nor U3800 (N_3800,N_990,N_834);
or U3801 (N_3801,N_1426,N_206);
and U3802 (N_3802,N_2429,N_1802);
nand U3803 (N_3803,N_1419,N_465);
and U3804 (N_3804,N_1605,N_831);
and U3805 (N_3805,N_1823,N_982);
nand U3806 (N_3806,N_985,N_1950);
nor U3807 (N_3807,N_1797,N_46);
or U3808 (N_3808,N_297,N_2372);
and U3809 (N_3809,N_1471,N_736);
nor U3810 (N_3810,N_837,N_864);
and U3811 (N_3811,N_232,N_1638);
nor U3812 (N_3812,N_396,N_1449);
nand U3813 (N_3813,N_393,N_780);
or U3814 (N_3814,N_1348,N_110);
nor U3815 (N_3815,N_2207,N_2229);
nor U3816 (N_3816,N_1512,N_1209);
nand U3817 (N_3817,N_1916,N_2470);
nor U3818 (N_3818,N_1143,N_1295);
nand U3819 (N_3819,N_174,N_2347);
or U3820 (N_3820,N_2001,N_89);
nor U3821 (N_3821,N_522,N_383);
or U3822 (N_3822,N_1168,N_1638);
nand U3823 (N_3823,N_2058,N_2126);
or U3824 (N_3824,N_711,N_263);
or U3825 (N_3825,N_728,N_523);
and U3826 (N_3826,N_701,N_1581);
nand U3827 (N_3827,N_2312,N_1008);
nor U3828 (N_3828,N_416,N_1735);
or U3829 (N_3829,N_318,N_347);
or U3830 (N_3830,N_2101,N_530);
or U3831 (N_3831,N_1116,N_1632);
or U3832 (N_3832,N_849,N_1721);
and U3833 (N_3833,N_2474,N_495);
nor U3834 (N_3834,N_521,N_1068);
nand U3835 (N_3835,N_1601,N_2248);
and U3836 (N_3836,N_1763,N_1698);
nand U3837 (N_3837,N_1057,N_1245);
nand U3838 (N_3838,N_983,N_2300);
and U3839 (N_3839,N_1409,N_63);
and U3840 (N_3840,N_649,N_792);
nand U3841 (N_3841,N_1773,N_2040);
or U3842 (N_3842,N_1201,N_346);
nand U3843 (N_3843,N_600,N_2007);
or U3844 (N_3844,N_1655,N_508);
or U3845 (N_3845,N_2258,N_1907);
and U3846 (N_3846,N_1763,N_490);
nor U3847 (N_3847,N_20,N_352);
and U3848 (N_3848,N_1185,N_862);
and U3849 (N_3849,N_1001,N_1830);
and U3850 (N_3850,N_401,N_1019);
nor U3851 (N_3851,N_36,N_1442);
and U3852 (N_3852,N_1581,N_1154);
nand U3853 (N_3853,N_2423,N_2031);
nor U3854 (N_3854,N_179,N_1300);
nor U3855 (N_3855,N_1185,N_1423);
nand U3856 (N_3856,N_979,N_1470);
or U3857 (N_3857,N_1547,N_554);
and U3858 (N_3858,N_344,N_1048);
nand U3859 (N_3859,N_460,N_377);
nand U3860 (N_3860,N_346,N_800);
and U3861 (N_3861,N_2279,N_1343);
or U3862 (N_3862,N_747,N_2285);
or U3863 (N_3863,N_50,N_1077);
and U3864 (N_3864,N_1410,N_1467);
nand U3865 (N_3865,N_1449,N_549);
nand U3866 (N_3866,N_1361,N_1264);
or U3867 (N_3867,N_1326,N_1991);
nand U3868 (N_3868,N_1743,N_788);
and U3869 (N_3869,N_944,N_2188);
nor U3870 (N_3870,N_317,N_891);
nand U3871 (N_3871,N_882,N_2485);
or U3872 (N_3872,N_964,N_1595);
or U3873 (N_3873,N_1143,N_2383);
nand U3874 (N_3874,N_2227,N_927);
nor U3875 (N_3875,N_1501,N_847);
or U3876 (N_3876,N_1354,N_315);
or U3877 (N_3877,N_474,N_677);
nand U3878 (N_3878,N_503,N_1524);
xnor U3879 (N_3879,N_6,N_2147);
and U3880 (N_3880,N_379,N_949);
nor U3881 (N_3881,N_1816,N_888);
nand U3882 (N_3882,N_963,N_80);
or U3883 (N_3883,N_1773,N_2402);
nand U3884 (N_3884,N_406,N_2142);
nor U3885 (N_3885,N_569,N_892);
nand U3886 (N_3886,N_1771,N_1644);
nand U3887 (N_3887,N_585,N_558);
nand U3888 (N_3888,N_1768,N_1832);
nor U3889 (N_3889,N_1472,N_2471);
or U3890 (N_3890,N_1128,N_168);
nand U3891 (N_3891,N_1099,N_2116);
and U3892 (N_3892,N_1336,N_1960);
and U3893 (N_3893,N_785,N_224);
nand U3894 (N_3894,N_1388,N_1062);
and U3895 (N_3895,N_879,N_1921);
or U3896 (N_3896,N_1564,N_50);
nand U3897 (N_3897,N_112,N_2361);
nor U3898 (N_3898,N_465,N_961);
and U3899 (N_3899,N_1673,N_1178);
and U3900 (N_3900,N_1252,N_1661);
and U3901 (N_3901,N_680,N_1705);
or U3902 (N_3902,N_1918,N_1166);
nand U3903 (N_3903,N_480,N_1502);
nor U3904 (N_3904,N_2038,N_601);
and U3905 (N_3905,N_2289,N_1035);
or U3906 (N_3906,N_940,N_31);
and U3907 (N_3907,N_1999,N_68);
and U3908 (N_3908,N_2348,N_1278);
nor U3909 (N_3909,N_298,N_2042);
nor U3910 (N_3910,N_232,N_101);
nand U3911 (N_3911,N_1211,N_483);
and U3912 (N_3912,N_444,N_1338);
or U3913 (N_3913,N_2208,N_459);
and U3914 (N_3914,N_471,N_758);
nor U3915 (N_3915,N_1205,N_1957);
nand U3916 (N_3916,N_620,N_919);
nand U3917 (N_3917,N_1335,N_1310);
or U3918 (N_3918,N_2023,N_1146);
or U3919 (N_3919,N_2333,N_1746);
nor U3920 (N_3920,N_1826,N_1364);
and U3921 (N_3921,N_2331,N_1514);
and U3922 (N_3922,N_1738,N_1349);
or U3923 (N_3923,N_1236,N_1057);
nand U3924 (N_3924,N_538,N_950);
and U3925 (N_3925,N_1744,N_461);
or U3926 (N_3926,N_2447,N_303);
nor U3927 (N_3927,N_2427,N_1515);
nor U3928 (N_3928,N_2155,N_2175);
nor U3929 (N_3929,N_881,N_928);
and U3930 (N_3930,N_905,N_1124);
or U3931 (N_3931,N_2320,N_1247);
nor U3932 (N_3932,N_112,N_1675);
and U3933 (N_3933,N_2402,N_817);
nand U3934 (N_3934,N_1690,N_1346);
nand U3935 (N_3935,N_349,N_1888);
nand U3936 (N_3936,N_1994,N_1716);
nor U3937 (N_3937,N_735,N_2238);
nor U3938 (N_3938,N_29,N_1714);
or U3939 (N_3939,N_2114,N_289);
nor U3940 (N_3940,N_870,N_2347);
and U3941 (N_3941,N_2138,N_1852);
nor U3942 (N_3942,N_621,N_1398);
or U3943 (N_3943,N_1202,N_2017);
or U3944 (N_3944,N_1433,N_1498);
nor U3945 (N_3945,N_796,N_2249);
and U3946 (N_3946,N_579,N_1326);
or U3947 (N_3947,N_615,N_2259);
nand U3948 (N_3948,N_1563,N_91);
nor U3949 (N_3949,N_938,N_1123);
nand U3950 (N_3950,N_1732,N_156);
nand U3951 (N_3951,N_1804,N_1955);
or U3952 (N_3952,N_239,N_285);
nor U3953 (N_3953,N_2302,N_1463);
or U3954 (N_3954,N_814,N_2496);
nor U3955 (N_3955,N_1550,N_351);
nor U3956 (N_3956,N_1573,N_1596);
or U3957 (N_3957,N_1002,N_2247);
or U3958 (N_3958,N_59,N_2452);
or U3959 (N_3959,N_1215,N_171);
and U3960 (N_3960,N_1694,N_527);
nand U3961 (N_3961,N_2310,N_1637);
and U3962 (N_3962,N_856,N_2159);
and U3963 (N_3963,N_146,N_1712);
nor U3964 (N_3964,N_736,N_1968);
and U3965 (N_3965,N_1408,N_447);
and U3966 (N_3966,N_1380,N_2436);
or U3967 (N_3967,N_2310,N_1686);
or U3968 (N_3968,N_2162,N_680);
nor U3969 (N_3969,N_1073,N_1239);
nor U3970 (N_3970,N_2029,N_732);
or U3971 (N_3971,N_2141,N_785);
nand U3972 (N_3972,N_56,N_370);
nand U3973 (N_3973,N_720,N_631);
and U3974 (N_3974,N_1214,N_1358);
or U3975 (N_3975,N_403,N_2462);
and U3976 (N_3976,N_2197,N_159);
nand U3977 (N_3977,N_1419,N_376);
and U3978 (N_3978,N_1635,N_898);
nand U3979 (N_3979,N_1961,N_677);
and U3980 (N_3980,N_2241,N_2358);
and U3981 (N_3981,N_274,N_1924);
or U3982 (N_3982,N_1710,N_2183);
and U3983 (N_3983,N_1093,N_151);
and U3984 (N_3984,N_1021,N_1530);
or U3985 (N_3985,N_1384,N_442);
or U3986 (N_3986,N_1989,N_2354);
nand U3987 (N_3987,N_1186,N_929);
nand U3988 (N_3988,N_1536,N_1086);
or U3989 (N_3989,N_119,N_47);
nand U3990 (N_3990,N_1862,N_624);
or U3991 (N_3991,N_585,N_1852);
nand U3992 (N_3992,N_1785,N_312);
or U3993 (N_3993,N_1032,N_616);
nand U3994 (N_3994,N_2408,N_1386);
nor U3995 (N_3995,N_34,N_2194);
and U3996 (N_3996,N_986,N_1955);
and U3997 (N_3997,N_270,N_1031);
nor U3998 (N_3998,N_376,N_1919);
or U3999 (N_3999,N_2156,N_1330);
and U4000 (N_4000,N_1184,N_870);
nand U4001 (N_4001,N_373,N_37);
or U4002 (N_4002,N_1486,N_58);
or U4003 (N_4003,N_768,N_2081);
nand U4004 (N_4004,N_1624,N_2411);
nor U4005 (N_4005,N_1101,N_2321);
and U4006 (N_4006,N_2310,N_1889);
and U4007 (N_4007,N_854,N_69);
nand U4008 (N_4008,N_528,N_1961);
xor U4009 (N_4009,N_922,N_393);
nand U4010 (N_4010,N_475,N_674);
and U4011 (N_4011,N_1211,N_2249);
nand U4012 (N_4012,N_241,N_1684);
nor U4013 (N_4013,N_2091,N_266);
or U4014 (N_4014,N_1988,N_109);
and U4015 (N_4015,N_672,N_201);
and U4016 (N_4016,N_395,N_1748);
or U4017 (N_4017,N_2312,N_186);
nand U4018 (N_4018,N_994,N_1928);
nor U4019 (N_4019,N_1087,N_2179);
nand U4020 (N_4020,N_867,N_175);
and U4021 (N_4021,N_1324,N_1687);
nand U4022 (N_4022,N_2210,N_1756);
nand U4023 (N_4023,N_1933,N_820);
nor U4024 (N_4024,N_126,N_179);
nand U4025 (N_4025,N_799,N_110);
nand U4026 (N_4026,N_1633,N_1040);
or U4027 (N_4027,N_1932,N_1487);
and U4028 (N_4028,N_394,N_1117);
and U4029 (N_4029,N_575,N_1227);
or U4030 (N_4030,N_2160,N_318);
nand U4031 (N_4031,N_237,N_1518);
or U4032 (N_4032,N_2426,N_756);
and U4033 (N_4033,N_1496,N_715);
and U4034 (N_4034,N_2312,N_979);
and U4035 (N_4035,N_1186,N_1782);
nand U4036 (N_4036,N_858,N_651);
nand U4037 (N_4037,N_1011,N_464);
and U4038 (N_4038,N_799,N_325);
and U4039 (N_4039,N_1429,N_1657);
nand U4040 (N_4040,N_2168,N_50);
nand U4041 (N_4041,N_485,N_2006);
nand U4042 (N_4042,N_1041,N_1825);
and U4043 (N_4043,N_220,N_656);
nor U4044 (N_4044,N_1583,N_957);
nand U4045 (N_4045,N_1027,N_171);
nand U4046 (N_4046,N_879,N_1937);
or U4047 (N_4047,N_825,N_1097);
nand U4048 (N_4048,N_1855,N_361);
nand U4049 (N_4049,N_1103,N_963);
and U4050 (N_4050,N_2226,N_1475);
nand U4051 (N_4051,N_1824,N_887);
nand U4052 (N_4052,N_1025,N_2489);
nor U4053 (N_4053,N_957,N_1575);
and U4054 (N_4054,N_2341,N_105);
nand U4055 (N_4055,N_1523,N_456);
xnor U4056 (N_4056,N_82,N_1092);
and U4057 (N_4057,N_1241,N_1761);
nor U4058 (N_4058,N_2358,N_1759);
nand U4059 (N_4059,N_1220,N_1524);
and U4060 (N_4060,N_1757,N_1455);
or U4061 (N_4061,N_1970,N_765);
nor U4062 (N_4062,N_2415,N_1774);
nand U4063 (N_4063,N_2043,N_1227);
and U4064 (N_4064,N_466,N_363);
xnor U4065 (N_4065,N_402,N_958);
nand U4066 (N_4066,N_139,N_429);
nor U4067 (N_4067,N_2285,N_1830);
or U4068 (N_4068,N_370,N_1764);
nand U4069 (N_4069,N_125,N_1552);
nand U4070 (N_4070,N_121,N_476);
or U4071 (N_4071,N_2112,N_2029);
nand U4072 (N_4072,N_561,N_2008);
nand U4073 (N_4073,N_348,N_2235);
and U4074 (N_4074,N_2400,N_465);
nand U4075 (N_4075,N_412,N_1227);
and U4076 (N_4076,N_1614,N_2497);
and U4077 (N_4077,N_1473,N_2226);
or U4078 (N_4078,N_883,N_1425);
or U4079 (N_4079,N_2427,N_2036);
and U4080 (N_4080,N_1787,N_2068);
xnor U4081 (N_4081,N_1445,N_2249);
nor U4082 (N_4082,N_431,N_1928);
and U4083 (N_4083,N_1467,N_1708);
xor U4084 (N_4084,N_230,N_1169);
and U4085 (N_4085,N_841,N_906);
or U4086 (N_4086,N_1441,N_1404);
or U4087 (N_4087,N_1859,N_2020);
and U4088 (N_4088,N_2044,N_657);
nor U4089 (N_4089,N_2416,N_2135);
or U4090 (N_4090,N_1378,N_2374);
and U4091 (N_4091,N_892,N_1114);
or U4092 (N_4092,N_712,N_947);
nor U4093 (N_4093,N_1087,N_2418);
nand U4094 (N_4094,N_502,N_1301);
and U4095 (N_4095,N_1406,N_182);
or U4096 (N_4096,N_823,N_883);
nand U4097 (N_4097,N_1222,N_112);
nor U4098 (N_4098,N_1111,N_380);
nor U4099 (N_4099,N_1777,N_247);
nor U4100 (N_4100,N_1962,N_1995);
and U4101 (N_4101,N_2079,N_158);
nand U4102 (N_4102,N_33,N_2261);
nand U4103 (N_4103,N_1784,N_2198);
nor U4104 (N_4104,N_493,N_1066);
nor U4105 (N_4105,N_628,N_1666);
nand U4106 (N_4106,N_1761,N_1139);
or U4107 (N_4107,N_1665,N_2399);
or U4108 (N_4108,N_2254,N_226);
and U4109 (N_4109,N_452,N_1869);
and U4110 (N_4110,N_2095,N_1777);
nor U4111 (N_4111,N_1126,N_218);
nor U4112 (N_4112,N_2310,N_826);
nand U4113 (N_4113,N_2251,N_1730);
nor U4114 (N_4114,N_409,N_1712);
xor U4115 (N_4115,N_670,N_270);
and U4116 (N_4116,N_1337,N_1872);
or U4117 (N_4117,N_1283,N_787);
or U4118 (N_4118,N_502,N_2471);
nand U4119 (N_4119,N_2343,N_1049);
and U4120 (N_4120,N_1365,N_1565);
nor U4121 (N_4121,N_962,N_1393);
or U4122 (N_4122,N_1858,N_1645);
nor U4123 (N_4123,N_339,N_1355);
and U4124 (N_4124,N_1745,N_1350);
nor U4125 (N_4125,N_630,N_927);
nand U4126 (N_4126,N_165,N_2401);
nor U4127 (N_4127,N_966,N_865);
and U4128 (N_4128,N_901,N_1600);
nor U4129 (N_4129,N_1954,N_257);
and U4130 (N_4130,N_876,N_431);
nor U4131 (N_4131,N_550,N_507);
or U4132 (N_4132,N_1052,N_1607);
or U4133 (N_4133,N_2197,N_861);
or U4134 (N_4134,N_1202,N_2241);
nor U4135 (N_4135,N_87,N_2124);
nand U4136 (N_4136,N_875,N_354);
nor U4137 (N_4137,N_1276,N_2302);
nor U4138 (N_4138,N_2312,N_1847);
or U4139 (N_4139,N_1587,N_226);
or U4140 (N_4140,N_638,N_1535);
nand U4141 (N_4141,N_1068,N_1140);
and U4142 (N_4142,N_1437,N_704);
nand U4143 (N_4143,N_2449,N_1333);
or U4144 (N_4144,N_1082,N_1495);
nand U4145 (N_4145,N_1839,N_107);
and U4146 (N_4146,N_616,N_331);
or U4147 (N_4147,N_108,N_1385);
nor U4148 (N_4148,N_1056,N_1766);
nor U4149 (N_4149,N_1816,N_1683);
nor U4150 (N_4150,N_1253,N_245);
nor U4151 (N_4151,N_1955,N_189);
or U4152 (N_4152,N_1741,N_620);
nand U4153 (N_4153,N_481,N_718);
and U4154 (N_4154,N_2438,N_2297);
nor U4155 (N_4155,N_133,N_2028);
nand U4156 (N_4156,N_1396,N_833);
and U4157 (N_4157,N_635,N_1536);
and U4158 (N_4158,N_1387,N_291);
and U4159 (N_4159,N_244,N_1912);
nor U4160 (N_4160,N_1326,N_1504);
nor U4161 (N_4161,N_778,N_751);
and U4162 (N_4162,N_2295,N_1441);
nand U4163 (N_4163,N_982,N_1697);
or U4164 (N_4164,N_1047,N_399);
nor U4165 (N_4165,N_1292,N_1108);
and U4166 (N_4166,N_988,N_2382);
and U4167 (N_4167,N_1742,N_385);
nor U4168 (N_4168,N_1346,N_2326);
nand U4169 (N_4169,N_844,N_2370);
nor U4170 (N_4170,N_2353,N_640);
and U4171 (N_4171,N_1396,N_1610);
nor U4172 (N_4172,N_1975,N_924);
and U4173 (N_4173,N_806,N_798);
nor U4174 (N_4174,N_2005,N_923);
or U4175 (N_4175,N_1286,N_1342);
and U4176 (N_4176,N_212,N_939);
and U4177 (N_4177,N_2232,N_802);
nor U4178 (N_4178,N_2220,N_605);
and U4179 (N_4179,N_2250,N_1768);
xor U4180 (N_4180,N_1890,N_2360);
and U4181 (N_4181,N_970,N_2125);
and U4182 (N_4182,N_522,N_2499);
and U4183 (N_4183,N_880,N_99);
and U4184 (N_4184,N_1307,N_1831);
nand U4185 (N_4185,N_2002,N_739);
nor U4186 (N_4186,N_1280,N_858);
nand U4187 (N_4187,N_299,N_2437);
nor U4188 (N_4188,N_309,N_194);
and U4189 (N_4189,N_1114,N_254);
or U4190 (N_4190,N_1426,N_1665);
nor U4191 (N_4191,N_117,N_601);
or U4192 (N_4192,N_764,N_971);
nor U4193 (N_4193,N_591,N_2241);
nand U4194 (N_4194,N_424,N_1551);
nor U4195 (N_4195,N_417,N_210);
nand U4196 (N_4196,N_2031,N_1874);
nor U4197 (N_4197,N_428,N_1643);
or U4198 (N_4198,N_178,N_2129);
and U4199 (N_4199,N_1507,N_1632);
or U4200 (N_4200,N_2126,N_485);
and U4201 (N_4201,N_863,N_1598);
nand U4202 (N_4202,N_1813,N_1101);
or U4203 (N_4203,N_219,N_652);
nand U4204 (N_4204,N_1335,N_660);
nor U4205 (N_4205,N_1776,N_661);
xor U4206 (N_4206,N_1651,N_1863);
or U4207 (N_4207,N_1367,N_2340);
or U4208 (N_4208,N_72,N_2064);
nor U4209 (N_4209,N_115,N_1477);
nor U4210 (N_4210,N_1410,N_2443);
and U4211 (N_4211,N_955,N_1477);
nor U4212 (N_4212,N_235,N_2197);
nor U4213 (N_4213,N_1141,N_1090);
nor U4214 (N_4214,N_1704,N_333);
nand U4215 (N_4215,N_1769,N_250);
or U4216 (N_4216,N_533,N_1385);
nor U4217 (N_4217,N_1370,N_1075);
nor U4218 (N_4218,N_1248,N_968);
and U4219 (N_4219,N_253,N_1773);
nand U4220 (N_4220,N_597,N_1378);
nor U4221 (N_4221,N_330,N_963);
or U4222 (N_4222,N_0,N_1881);
or U4223 (N_4223,N_965,N_1800);
nor U4224 (N_4224,N_2463,N_855);
nor U4225 (N_4225,N_962,N_134);
nor U4226 (N_4226,N_1574,N_1298);
or U4227 (N_4227,N_1229,N_917);
or U4228 (N_4228,N_2134,N_103);
and U4229 (N_4229,N_2232,N_1230);
nor U4230 (N_4230,N_509,N_1031);
nand U4231 (N_4231,N_1672,N_1287);
and U4232 (N_4232,N_352,N_424);
nand U4233 (N_4233,N_1972,N_2070);
nor U4234 (N_4234,N_1507,N_550);
nor U4235 (N_4235,N_2151,N_448);
or U4236 (N_4236,N_122,N_1407);
or U4237 (N_4237,N_522,N_2327);
nor U4238 (N_4238,N_1607,N_1769);
and U4239 (N_4239,N_243,N_1922);
nor U4240 (N_4240,N_1897,N_718);
nand U4241 (N_4241,N_358,N_2433);
nor U4242 (N_4242,N_1608,N_681);
nor U4243 (N_4243,N_1310,N_658);
nor U4244 (N_4244,N_705,N_2358);
or U4245 (N_4245,N_886,N_2341);
nor U4246 (N_4246,N_2348,N_141);
xnor U4247 (N_4247,N_1472,N_1873);
nor U4248 (N_4248,N_1011,N_400);
nand U4249 (N_4249,N_2340,N_696);
and U4250 (N_4250,N_404,N_1282);
or U4251 (N_4251,N_1182,N_1391);
and U4252 (N_4252,N_1370,N_2000);
nand U4253 (N_4253,N_1070,N_2237);
xor U4254 (N_4254,N_1288,N_303);
nor U4255 (N_4255,N_643,N_116);
or U4256 (N_4256,N_1299,N_1529);
or U4257 (N_4257,N_656,N_1032);
nand U4258 (N_4258,N_463,N_1224);
nand U4259 (N_4259,N_1939,N_2302);
nor U4260 (N_4260,N_1916,N_407);
nor U4261 (N_4261,N_1505,N_1357);
or U4262 (N_4262,N_564,N_2279);
or U4263 (N_4263,N_1353,N_562);
nor U4264 (N_4264,N_1784,N_1695);
and U4265 (N_4265,N_2326,N_1813);
and U4266 (N_4266,N_1523,N_1732);
or U4267 (N_4267,N_808,N_2478);
nand U4268 (N_4268,N_1557,N_2104);
or U4269 (N_4269,N_8,N_543);
and U4270 (N_4270,N_974,N_667);
nand U4271 (N_4271,N_490,N_1043);
and U4272 (N_4272,N_94,N_366);
nor U4273 (N_4273,N_244,N_2053);
and U4274 (N_4274,N_2272,N_925);
nand U4275 (N_4275,N_1053,N_1849);
and U4276 (N_4276,N_2381,N_1164);
and U4277 (N_4277,N_123,N_2011);
nor U4278 (N_4278,N_2185,N_221);
nand U4279 (N_4279,N_1462,N_2457);
and U4280 (N_4280,N_1836,N_539);
nor U4281 (N_4281,N_2227,N_1661);
nor U4282 (N_4282,N_1976,N_2108);
nand U4283 (N_4283,N_1800,N_626);
nand U4284 (N_4284,N_568,N_1030);
nor U4285 (N_4285,N_2402,N_2092);
and U4286 (N_4286,N_871,N_2497);
and U4287 (N_4287,N_419,N_905);
or U4288 (N_4288,N_179,N_543);
and U4289 (N_4289,N_2469,N_949);
or U4290 (N_4290,N_1174,N_2462);
and U4291 (N_4291,N_1294,N_2330);
nand U4292 (N_4292,N_1716,N_2075);
nand U4293 (N_4293,N_577,N_1870);
or U4294 (N_4294,N_1641,N_773);
and U4295 (N_4295,N_161,N_1690);
nor U4296 (N_4296,N_87,N_934);
nor U4297 (N_4297,N_867,N_1753);
and U4298 (N_4298,N_2390,N_701);
or U4299 (N_4299,N_1355,N_315);
and U4300 (N_4300,N_211,N_1689);
or U4301 (N_4301,N_1415,N_1904);
or U4302 (N_4302,N_1168,N_1752);
nor U4303 (N_4303,N_1328,N_218);
nor U4304 (N_4304,N_728,N_1089);
nor U4305 (N_4305,N_862,N_2098);
and U4306 (N_4306,N_2147,N_979);
nand U4307 (N_4307,N_1147,N_829);
nor U4308 (N_4308,N_973,N_2158);
and U4309 (N_4309,N_1905,N_880);
or U4310 (N_4310,N_1173,N_737);
nor U4311 (N_4311,N_312,N_2285);
nand U4312 (N_4312,N_347,N_1695);
and U4313 (N_4313,N_1578,N_207);
or U4314 (N_4314,N_22,N_1835);
nor U4315 (N_4315,N_1502,N_2395);
and U4316 (N_4316,N_139,N_2375);
or U4317 (N_4317,N_1969,N_2270);
and U4318 (N_4318,N_2474,N_865);
and U4319 (N_4319,N_1003,N_147);
or U4320 (N_4320,N_938,N_631);
nand U4321 (N_4321,N_499,N_791);
nand U4322 (N_4322,N_1858,N_1616);
or U4323 (N_4323,N_2246,N_373);
nand U4324 (N_4324,N_1226,N_361);
nand U4325 (N_4325,N_245,N_1678);
or U4326 (N_4326,N_1451,N_740);
nand U4327 (N_4327,N_801,N_1462);
nor U4328 (N_4328,N_642,N_2121);
nand U4329 (N_4329,N_1725,N_197);
and U4330 (N_4330,N_440,N_570);
and U4331 (N_4331,N_2106,N_2445);
or U4332 (N_4332,N_436,N_1619);
nor U4333 (N_4333,N_24,N_2036);
nor U4334 (N_4334,N_127,N_662);
and U4335 (N_4335,N_849,N_1005);
nor U4336 (N_4336,N_2109,N_2301);
and U4337 (N_4337,N_958,N_2078);
nand U4338 (N_4338,N_881,N_650);
nand U4339 (N_4339,N_1953,N_1117);
and U4340 (N_4340,N_2081,N_566);
and U4341 (N_4341,N_614,N_1029);
nor U4342 (N_4342,N_135,N_571);
nor U4343 (N_4343,N_842,N_1997);
nor U4344 (N_4344,N_180,N_2238);
nand U4345 (N_4345,N_1704,N_664);
nor U4346 (N_4346,N_1169,N_1583);
nor U4347 (N_4347,N_138,N_2252);
or U4348 (N_4348,N_1109,N_1591);
nor U4349 (N_4349,N_1478,N_2184);
and U4350 (N_4350,N_414,N_2098);
nor U4351 (N_4351,N_1959,N_355);
nor U4352 (N_4352,N_2314,N_2236);
nor U4353 (N_4353,N_2283,N_514);
or U4354 (N_4354,N_1680,N_1270);
or U4355 (N_4355,N_794,N_1974);
or U4356 (N_4356,N_1883,N_71);
or U4357 (N_4357,N_1884,N_2201);
and U4358 (N_4358,N_485,N_1107);
and U4359 (N_4359,N_174,N_383);
nor U4360 (N_4360,N_1132,N_414);
or U4361 (N_4361,N_827,N_2165);
nor U4362 (N_4362,N_1978,N_1299);
nor U4363 (N_4363,N_1166,N_2185);
or U4364 (N_4364,N_1724,N_2040);
nand U4365 (N_4365,N_911,N_1412);
nor U4366 (N_4366,N_1334,N_2352);
nand U4367 (N_4367,N_252,N_746);
nand U4368 (N_4368,N_1539,N_2047);
and U4369 (N_4369,N_1788,N_62);
and U4370 (N_4370,N_2470,N_44);
and U4371 (N_4371,N_1468,N_609);
and U4372 (N_4372,N_1751,N_1473);
and U4373 (N_4373,N_525,N_1916);
or U4374 (N_4374,N_171,N_1988);
nor U4375 (N_4375,N_1718,N_936);
and U4376 (N_4376,N_1844,N_2100);
and U4377 (N_4377,N_243,N_1786);
and U4378 (N_4378,N_1815,N_1295);
or U4379 (N_4379,N_671,N_871);
and U4380 (N_4380,N_485,N_420);
nand U4381 (N_4381,N_2389,N_706);
and U4382 (N_4382,N_1089,N_37);
nand U4383 (N_4383,N_666,N_2343);
or U4384 (N_4384,N_2100,N_642);
xor U4385 (N_4385,N_1460,N_998);
and U4386 (N_4386,N_2490,N_254);
nor U4387 (N_4387,N_1651,N_9);
nor U4388 (N_4388,N_1160,N_1740);
nor U4389 (N_4389,N_2476,N_1875);
and U4390 (N_4390,N_1298,N_591);
and U4391 (N_4391,N_45,N_1701);
or U4392 (N_4392,N_1505,N_420);
nor U4393 (N_4393,N_42,N_200);
nor U4394 (N_4394,N_952,N_988);
or U4395 (N_4395,N_1295,N_337);
nand U4396 (N_4396,N_311,N_1403);
and U4397 (N_4397,N_1506,N_757);
nor U4398 (N_4398,N_140,N_1463);
nor U4399 (N_4399,N_338,N_1795);
nor U4400 (N_4400,N_1230,N_101);
nand U4401 (N_4401,N_400,N_2008);
and U4402 (N_4402,N_422,N_352);
or U4403 (N_4403,N_1840,N_653);
nor U4404 (N_4404,N_515,N_1238);
nor U4405 (N_4405,N_597,N_1306);
nand U4406 (N_4406,N_1197,N_1050);
nor U4407 (N_4407,N_1351,N_1086);
nand U4408 (N_4408,N_1864,N_256);
xnor U4409 (N_4409,N_2126,N_2494);
and U4410 (N_4410,N_1902,N_437);
or U4411 (N_4411,N_2487,N_1429);
nor U4412 (N_4412,N_1510,N_488);
nor U4413 (N_4413,N_1010,N_1534);
or U4414 (N_4414,N_1902,N_2148);
nand U4415 (N_4415,N_2243,N_245);
or U4416 (N_4416,N_69,N_833);
or U4417 (N_4417,N_1706,N_1882);
or U4418 (N_4418,N_1444,N_318);
and U4419 (N_4419,N_1437,N_283);
nor U4420 (N_4420,N_226,N_253);
and U4421 (N_4421,N_1941,N_0);
or U4422 (N_4422,N_491,N_88);
and U4423 (N_4423,N_1543,N_1935);
nor U4424 (N_4424,N_2074,N_187);
and U4425 (N_4425,N_1987,N_448);
or U4426 (N_4426,N_1468,N_196);
or U4427 (N_4427,N_1269,N_465);
nor U4428 (N_4428,N_805,N_1366);
nand U4429 (N_4429,N_116,N_865);
or U4430 (N_4430,N_684,N_2006);
or U4431 (N_4431,N_576,N_2056);
nand U4432 (N_4432,N_1107,N_1654);
nor U4433 (N_4433,N_901,N_1910);
nor U4434 (N_4434,N_2130,N_905);
or U4435 (N_4435,N_1232,N_1900);
or U4436 (N_4436,N_1238,N_1653);
and U4437 (N_4437,N_2194,N_1112);
nand U4438 (N_4438,N_1832,N_1776);
nand U4439 (N_4439,N_1547,N_1630);
and U4440 (N_4440,N_2099,N_2339);
and U4441 (N_4441,N_948,N_145);
nand U4442 (N_4442,N_813,N_1605);
nor U4443 (N_4443,N_211,N_1615);
nor U4444 (N_4444,N_796,N_1831);
or U4445 (N_4445,N_1500,N_1868);
nand U4446 (N_4446,N_784,N_2450);
and U4447 (N_4447,N_58,N_2240);
or U4448 (N_4448,N_1081,N_1992);
nor U4449 (N_4449,N_2360,N_1239);
or U4450 (N_4450,N_304,N_2000);
nand U4451 (N_4451,N_2396,N_826);
nor U4452 (N_4452,N_34,N_1907);
nand U4453 (N_4453,N_1545,N_2302);
and U4454 (N_4454,N_661,N_1819);
nor U4455 (N_4455,N_1124,N_252);
and U4456 (N_4456,N_1928,N_1116);
and U4457 (N_4457,N_570,N_538);
or U4458 (N_4458,N_1932,N_373);
nor U4459 (N_4459,N_962,N_2112);
nand U4460 (N_4460,N_562,N_2122);
or U4461 (N_4461,N_1245,N_437);
nor U4462 (N_4462,N_437,N_587);
and U4463 (N_4463,N_2092,N_1947);
nor U4464 (N_4464,N_474,N_2017);
or U4465 (N_4465,N_978,N_1472);
nand U4466 (N_4466,N_1010,N_1783);
nor U4467 (N_4467,N_610,N_2055);
nor U4468 (N_4468,N_1592,N_686);
and U4469 (N_4469,N_1689,N_656);
nand U4470 (N_4470,N_363,N_1798);
nand U4471 (N_4471,N_196,N_2278);
and U4472 (N_4472,N_405,N_465);
and U4473 (N_4473,N_2013,N_579);
nor U4474 (N_4474,N_392,N_706);
and U4475 (N_4475,N_499,N_1497);
and U4476 (N_4476,N_1979,N_467);
or U4477 (N_4477,N_1684,N_1127);
and U4478 (N_4478,N_1156,N_1107);
nor U4479 (N_4479,N_1558,N_98);
nand U4480 (N_4480,N_584,N_1459);
nor U4481 (N_4481,N_268,N_806);
and U4482 (N_4482,N_2089,N_1154);
nand U4483 (N_4483,N_797,N_1405);
and U4484 (N_4484,N_932,N_2193);
or U4485 (N_4485,N_1424,N_442);
and U4486 (N_4486,N_2007,N_405);
nand U4487 (N_4487,N_1851,N_992);
nand U4488 (N_4488,N_1832,N_1815);
nand U4489 (N_4489,N_796,N_1680);
and U4490 (N_4490,N_1930,N_2228);
or U4491 (N_4491,N_1550,N_195);
or U4492 (N_4492,N_2335,N_707);
or U4493 (N_4493,N_436,N_1239);
nor U4494 (N_4494,N_1059,N_2070);
or U4495 (N_4495,N_571,N_1453);
and U4496 (N_4496,N_1138,N_813);
nand U4497 (N_4497,N_523,N_2037);
and U4498 (N_4498,N_884,N_2189);
nand U4499 (N_4499,N_2210,N_640);
nor U4500 (N_4500,N_1346,N_1451);
nor U4501 (N_4501,N_1215,N_494);
or U4502 (N_4502,N_1823,N_388);
or U4503 (N_4503,N_598,N_681);
or U4504 (N_4504,N_195,N_1231);
nor U4505 (N_4505,N_415,N_974);
and U4506 (N_4506,N_457,N_899);
or U4507 (N_4507,N_1260,N_203);
nand U4508 (N_4508,N_1452,N_2265);
nor U4509 (N_4509,N_2364,N_1881);
and U4510 (N_4510,N_1199,N_1587);
nor U4511 (N_4511,N_33,N_330);
nor U4512 (N_4512,N_572,N_2373);
and U4513 (N_4513,N_979,N_871);
or U4514 (N_4514,N_1675,N_415);
and U4515 (N_4515,N_75,N_1196);
or U4516 (N_4516,N_2021,N_2120);
or U4517 (N_4517,N_1704,N_2200);
or U4518 (N_4518,N_2148,N_645);
and U4519 (N_4519,N_1481,N_2102);
nand U4520 (N_4520,N_1159,N_1025);
nand U4521 (N_4521,N_452,N_893);
nor U4522 (N_4522,N_1599,N_630);
nand U4523 (N_4523,N_1354,N_2240);
and U4524 (N_4524,N_1306,N_1537);
nand U4525 (N_4525,N_1521,N_260);
nand U4526 (N_4526,N_1247,N_477);
nor U4527 (N_4527,N_506,N_394);
nor U4528 (N_4528,N_1123,N_1249);
or U4529 (N_4529,N_1114,N_1856);
nand U4530 (N_4530,N_2397,N_1690);
nand U4531 (N_4531,N_1952,N_1831);
nand U4532 (N_4532,N_2034,N_2354);
nand U4533 (N_4533,N_799,N_10);
and U4534 (N_4534,N_1493,N_309);
and U4535 (N_4535,N_2481,N_230);
nor U4536 (N_4536,N_2262,N_1415);
or U4537 (N_4537,N_116,N_576);
and U4538 (N_4538,N_1199,N_2043);
or U4539 (N_4539,N_1965,N_1072);
nand U4540 (N_4540,N_1658,N_1252);
nand U4541 (N_4541,N_200,N_1779);
or U4542 (N_4542,N_950,N_207);
or U4543 (N_4543,N_2125,N_2331);
nor U4544 (N_4544,N_1963,N_935);
nand U4545 (N_4545,N_1500,N_363);
and U4546 (N_4546,N_2029,N_1620);
or U4547 (N_4547,N_586,N_1546);
or U4548 (N_4548,N_322,N_446);
nand U4549 (N_4549,N_1195,N_2082);
nand U4550 (N_4550,N_1336,N_1346);
and U4551 (N_4551,N_2090,N_253);
nor U4552 (N_4552,N_1050,N_1593);
and U4553 (N_4553,N_2169,N_164);
and U4554 (N_4554,N_1262,N_1376);
and U4555 (N_4555,N_407,N_1980);
or U4556 (N_4556,N_2376,N_2005);
nor U4557 (N_4557,N_1164,N_1179);
nor U4558 (N_4558,N_2477,N_2316);
or U4559 (N_4559,N_1376,N_337);
nor U4560 (N_4560,N_629,N_1077);
nor U4561 (N_4561,N_150,N_1135);
or U4562 (N_4562,N_1973,N_1775);
and U4563 (N_4563,N_2005,N_1751);
and U4564 (N_4564,N_54,N_921);
nor U4565 (N_4565,N_1740,N_1558);
or U4566 (N_4566,N_2098,N_513);
nand U4567 (N_4567,N_1661,N_1193);
nand U4568 (N_4568,N_1203,N_1913);
and U4569 (N_4569,N_510,N_1476);
or U4570 (N_4570,N_60,N_1776);
nor U4571 (N_4571,N_1725,N_295);
nand U4572 (N_4572,N_890,N_1706);
nand U4573 (N_4573,N_1962,N_2129);
nor U4574 (N_4574,N_721,N_1406);
nand U4575 (N_4575,N_2180,N_1797);
or U4576 (N_4576,N_2494,N_1182);
nor U4577 (N_4577,N_1720,N_588);
nand U4578 (N_4578,N_1488,N_2119);
nand U4579 (N_4579,N_786,N_1301);
and U4580 (N_4580,N_1941,N_1664);
and U4581 (N_4581,N_2027,N_2357);
nor U4582 (N_4582,N_1434,N_725);
or U4583 (N_4583,N_493,N_419);
and U4584 (N_4584,N_58,N_291);
and U4585 (N_4585,N_2278,N_2424);
and U4586 (N_4586,N_1311,N_623);
or U4587 (N_4587,N_806,N_1769);
nand U4588 (N_4588,N_1291,N_1854);
and U4589 (N_4589,N_402,N_803);
nor U4590 (N_4590,N_753,N_1635);
xor U4591 (N_4591,N_735,N_2392);
and U4592 (N_4592,N_731,N_834);
nand U4593 (N_4593,N_16,N_1396);
and U4594 (N_4594,N_1386,N_552);
nor U4595 (N_4595,N_465,N_1376);
or U4596 (N_4596,N_1158,N_2009);
nor U4597 (N_4597,N_2132,N_2021);
nor U4598 (N_4598,N_349,N_440);
or U4599 (N_4599,N_1076,N_1320);
nand U4600 (N_4600,N_1729,N_1741);
nand U4601 (N_4601,N_1495,N_193);
nor U4602 (N_4602,N_823,N_392);
and U4603 (N_4603,N_1379,N_914);
or U4604 (N_4604,N_770,N_2381);
and U4605 (N_4605,N_143,N_2361);
and U4606 (N_4606,N_603,N_1057);
or U4607 (N_4607,N_1264,N_1371);
nor U4608 (N_4608,N_1949,N_288);
nand U4609 (N_4609,N_1046,N_322);
nand U4610 (N_4610,N_648,N_2212);
or U4611 (N_4611,N_803,N_712);
and U4612 (N_4612,N_1041,N_2438);
or U4613 (N_4613,N_2076,N_2168);
and U4614 (N_4614,N_2449,N_2353);
or U4615 (N_4615,N_2187,N_1310);
nor U4616 (N_4616,N_1759,N_1411);
and U4617 (N_4617,N_192,N_2233);
nand U4618 (N_4618,N_62,N_389);
or U4619 (N_4619,N_550,N_1882);
nand U4620 (N_4620,N_1664,N_1401);
or U4621 (N_4621,N_749,N_785);
and U4622 (N_4622,N_886,N_2178);
or U4623 (N_4623,N_119,N_613);
or U4624 (N_4624,N_1656,N_852);
nor U4625 (N_4625,N_321,N_79);
nand U4626 (N_4626,N_928,N_374);
or U4627 (N_4627,N_954,N_1572);
and U4628 (N_4628,N_2037,N_1750);
nor U4629 (N_4629,N_2492,N_805);
nand U4630 (N_4630,N_359,N_473);
or U4631 (N_4631,N_244,N_146);
and U4632 (N_4632,N_2002,N_1759);
and U4633 (N_4633,N_2023,N_1447);
or U4634 (N_4634,N_2081,N_913);
nand U4635 (N_4635,N_692,N_427);
nor U4636 (N_4636,N_610,N_1023);
and U4637 (N_4637,N_136,N_340);
and U4638 (N_4638,N_756,N_1639);
or U4639 (N_4639,N_167,N_1722);
or U4640 (N_4640,N_1277,N_1466);
nand U4641 (N_4641,N_1494,N_1082);
nor U4642 (N_4642,N_2093,N_1973);
nor U4643 (N_4643,N_1133,N_2191);
nor U4644 (N_4644,N_581,N_565);
xnor U4645 (N_4645,N_1354,N_1618);
or U4646 (N_4646,N_1025,N_1030);
nor U4647 (N_4647,N_915,N_1672);
and U4648 (N_4648,N_603,N_497);
nand U4649 (N_4649,N_2327,N_761);
xnor U4650 (N_4650,N_1048,N_2342);
or U4651 (N_4651,N_2486,N_1938);
or U4652 (N_4652,N_544,N_2391);
and U4653 (N_4653,N_977,N_1068);
nor U4654 (N_4654,N_1714,N_1517);
nand U4655 (N_4655,N_1182,N_1082);
nor U4656 (N_4656,N_854,N_2266);
nor U4657 (N_4657,N_780,N_371);
and U4658 (N_4658,N_1790,N_2148);
nor U4659 (N_4659,N_365,N_2479);
or U4660 (N_4660,N_551,N_1461);
nor U4661 (N_4661,N_388,N_1331);
or U4662 (N_4662,N_485,N_2212);
nand U4663 (N_4663,N_2237,N_1556);
nand U4664 (N_4664,N_2234,N_1995);
nor U4665 (N_4665,N_957,N_1319);
nand U4666 (N_4666,N_1620,N_642);
nand U4667 (N_4667,N_2128,N_1405);
or U4668 (N_4668,N_117,N_34);
and U4669 (N_4669,N_1185,N_413);
nand U4670 (N_4670,N_208,N_1447);
or U4671 (N_4671,N_695,N_1551);
nor U4672 (N_4672,N_934,N_1976);
and U4673 (N_4673,N_2165,N_507);
or U4674 (N_4674,N_308,N_402);
nor U4675 (N_4675,N_39,N_1688);
nand U4676 (N_4676,N_870,N_456);
xor U4677 (N_4677,N_529,N_975);
nor U4678 (N_4678,N_2057,N_151);
and U4679 (N_4679,N_1688,N_1400);
and U4680 (N_4680,N_778,N_1743);
nor U4681 (N_4681,N_961,N_2050);
and U4682 (N_4682,N_2493,N_913);
nand U4683 (N_4683,N_1162,N_1721);
and U4684 (N_4684,N_1881,N_937);
and U4685 (N_4685,N_205,N_683);
or U4686 (N_4686,N_2374,N_1476);
or U4687 (N_4687,N_1646,N_446);
nand U4688 (N_4688,N_2465,N_2453);
nand U4689 (N_4689,N_13,N_2118);
nand U4690 (N_4690,N_2377,N_1437);
and U4691 (N_4691,N_1908,N_21);
and U4692 (N_4692,N_2343,N_639);
xnor U4693 (N_4693,N_750,N_7);
or U4694 (N_4694,N_2325,N_1328);
nor U4695 (N_4695,N_340,N_1288);
nor U4696 (N_4696,N_481,N_1758);
and U4697 (N_4697,N_1705,N_1291);
nand U4698 (N_4698,N_1414,N_329);
or U4699 (N_4699,N_713,N_2174);
and U4700 (N_4700,N_797,N_431);
nor U4701 (N_4701,N_1036,N_2092);
and U4702 (N_4702,N_561,N_282);
or U4703 (N_4703,N_529,N_2162);
or U4704 (N_4704,N_2286,N_444);
or U4705 (N_4705,N_1946,N_1058);
or U4706 (N_4706,N_185,N_1365);
nor U4707 (N_4707,N_611,N_2379);
nor U4708 (N_4708,N_264,N_1959);
nor U4709 (N_4709,N_1434,N_1105);
and U4710 (N_4710,N_2244,N_1598);
or U4711 (N_4711,N_1209,N_1237);
nand U4712 (N_4712,N_1701,N_1139);
or U4713 (N_4713,N_2139,N_85);
nand U4714 (N_4714,N_1779,N_290);
xor U4715 (N_4715,N_2240,N_680);
nand U4716 (N_4716,N_1461,N_2296);
and U4717 (N_4717,N_140,N_1615);
and U4718 (N_4718,N_2221,N_329);
and U4719 (N_4719,N_51,N_1996);
nor U4720 (N_4720,N_1474,N_221);
or U4721 (N_4721,N_2211,N_1478);
nand U4722 (N_4722,N_1022,N_1299);
and U4723 (N_4723,N_626,N_2457);
xnor U4724 (N_4724,N_1893,N_1073);
or U4725 (N_4725,N_2429,N_2016);
or U4726 (N_4726,N_2057,N_1603);
nand U4727 (N_4727,N_1669,N_2142);
nor U4728 (N_4728,N_16,N_2056);
and U4729 (N_4729,N_98,N_128);
nand U4730 (N_4730,N_2208,N_1250);
and U4731 (N_4731,N_1414,N_901);
or U4732 (N_4732,N_375,N_11);
or U4733 (N_4733,N_627,N_2454);
and U4734 (N_4734,N_1448,N_261);
nor U4735 (N_4735,N_2482,N_389);
nand U4736 (N_4736,N_2465,N_2334);
or U4737 (N_4737,N_59,N_2131);
or U4738 (N_4738,N_496,N_2449);
and U4739 (N_4739,N_728,N_2475);
or U4740 (N_4740,N_1844,N_104);
and U4741 (N_4741,N_1737,N_945);
nor U4742 (N_4742,N_1285,N_2278);
or U4743 (N_4743,N_520,N_847);
nor U4744 (N_4744,N_1375,N_785);
and U4745 (N_4745,N_481,N_1451);
and U4746 (N_4746,N_2029,N_2237);
and U4747 (N_4747,N_686,N_34);
nor U4748 (N_4748,N_1604,N_1562);
or U4749 (N_4749,N_1845,N_1681);
nand U4750 (N_4750,N_2289,N_2107);
nor U4751 (N_4751,N_1955,N_2185);
nor U4752 (N_4752,N_1696,N_1819);
nor U4753 (N_4753,N_642,N_993);
nand U4754 (N_4754,N_1028,N_695);
nor U4755 (N_4755,N_816,N_2330);
nand U4756 (N_4756,N_917,N_1684);
and U4757 (N_4757,N_1542,N_1950);
nor U4758 (N_4758,N_803,N_1009);
nand U4759 (N_4759,N_1542,N_632);
nand U4760 (N_4760,N_637,N_361);
nand U4761 (N_4761,N_1311,N_17);
and U4762 (N_4762,N_1758,N_1687);
nand U4763 (N_4763,N_280,N_1140);
nand U4764 (N_4764,N_1618,N_1356);
nor U4765 (N_4765,N_1097,N_618);
or U4766 (N_4766,N_1345,N_1238);
or U4767 (N_4767,N_1299,N_1873);
and U4768 (N_4768,N_1014,N_2357);
nand U4769 (N_4769,N_1500,N_631);
nand U4770 (N_4770,N_53,N_935);
nor U4771 (N_4771,N_1625,N_2083);
and U4772 (N_4772,N_1718,N_131);
nor U4773 (N_4773,N_142,N_1143);
nor U4774 (N_4774,N_1678,N_625);
nand U4775 (N_4775,N_1439,N_210);
nand U4776 (N_4776,N_581,N_159);
and U4777 (N_4777,N_1730,N_1795);
nand U4778 (N_4778,N_1255,N_1347);
nand U4779 (N_4779,N_1587,N_1486);
xor U4780 (N_4780,N_887,N_1434);
nor U4781 (N_4781,N_2162,N_872);
nand U4782 (N_4782,N_1147,N_1176);
nand U4783 (N_4783,N_2190,N_404);
or U4784 (N_4784,N_1570,N_428);
nor U4785 (N_4785,N_29,N_1819);
nand U4786 (N_4786,N_2458,N_1794);
and U4787 (N_4787,N_2455,N_1286);
nor U4788 (N_4788,N_1877,N_1046);
and U4789 (N_4789,N_358,N_2206);
nand U4790 (N_4790,N_937,N_18);
nand U4791 (N_4791,N_2396,N_1482);
or U4792 (N_4792,N_1052,N_2048);
nor U4793 (N_4793,N_659,N_2026);
nand U4794 (N_4794,N_769,N_1493);
and U4795 (N_4795,N_1689,N_631);
nor U4796 (N_4796,N_493,N_2051);
or U4797 (N_4797,N_2364,N_972);
nor U4798 (N_4798,N_1298,N_1714);
and U4799 (N_4799,N_1404,N_1403);
or U4800 (N_4800,N_2016,N_58);
nor U4801 (N_4801,N_390,N_1990);
nor U4802 (N_4802,N_345,N_241);
or U4803 (N_4803,N_612,N_1876);
and U4804 (N_4804,N_201,N_1475);
or U4805 (N_4805,N_1130,N_1593);
and U4806 (N_4806,N_1835,N_1375);
nand U4807 (N_4807,N_822,N_1496);
or U4808 (N_4808,N_2266,N_583);
and U4809 (N_4809,N_487,N_66);
and U4810 (N_4810,N_1357,N_242);
or U4811 (N_4811,N_395,N_979);
nand U4812 (N_4812,N_1620,N_293);
nor U4813 (N_4813,N_1808,N_1213);
xnor U4814 (N_4814,N_628,N_734);
nand U4815 (N_4815,N_147,N_268);
and U4816 (N_4816,N_1427,N_554);
and U4817 (N_4817,N_2332,N_650);
and U4818 (N_4818,N_1704,N_2381);
and U4819 (N_4819,N_42,N_575);
nor U4820 (N_4820,N_175,N_455);
and U4821 (N_4821,N_2415,N_1661);
or U4822 (N_4822,N_13,N_733);
and U4823 (N_4823,N_1869,N_709);
nor U4824 (N_4824,N_268,N_585);
xnor U4825 (N_4825,N_2184,N_2341);
and U4826 (N_4826,N_1358,N_1841);
nand U4827 (N_4827,N_609,N_2176);
nand U4828 (N_4828,N_2188,N_748);
nor U4829 (N_4829,N_2461,N_2085);
and U4830 (N_4830,N_214,N_2186);
nand U4831 (N_4831,N_403,N_1311);
nor U4832 (N_4832,N_1785,N_714);
and U4833 (N_4833,N_2492,N_1303);
nor U4834 (N_4834,N_1224,N_1820);
nor U4835 (N_4835,N_1442,N_283);
nor U4836 (N_4836,N_273,N_1420);
or U4837 (N_4837,N_2230,N_1840);
or U4838 (N_4838,N_859,N_2481);
nand U4839 (N_4839,N_1247,N_2124);
and U4840 (N_4840,N_1452,N_1007);
or U4841 (N_4841,N_1457,N_2378);
nand U4842 (N_4842,N_1754,N_1573);
and U4843 (N_4843,N_2441,N_284);
nor U4844 (N_4844,N_882,N_1521);
nor U4845 (N_4845,N_470,N_1676);
or U4846 (N_4846,N_739,N_2296);
or U4847 (N_4847,N_810,N_1828);
xnor U4848 (N_4848,N_2295,N_1622);
or U4849 (N_4849,N_2240,N_1642);
or U4850 (N_4850,N_2400,N_251);
and U4851 (N_4851,N_27,N_1522);
nand U4852 (N_4852,N_95,N_566);
or U4853 (N_4853,N_2228,N_2085);
nand U4854 (N_4854,N_973,N_1120);
nand U4855 (N_4855,N_735,N_160);
nand U4856 (N_4856,N_5,N_1547);
or U4857 (N_4857,N_1167,N_2073);
nand U4858 (N_4858,N_1079,N_1792);
nor U4859 (N_4859,N_750,N_1765);
nor U4860 (N_4860,N_1225,N_2351);
nor U4861 (N_4861,N_410,N_295);
nor U4862 (N_4862,N_2317,N_698);
or U4863 (N_4863,N_170,N_1031);
and U4864 (N_4864,N_2260,N_1908);
nand U4865 (N_4865,N_661,N_1453);
or U4866 (N_4866,N_2458,N_901);
or U4867 (N_4867,N_666,N_2074);
or U4868 (N_4868,N_661,N_505);
and U4869 (N_4869,N_1896,N_2125);
nand U4870 (N_4870,N_120,N_103);
nor U4871 (N_4871,N_349,N_2095);
nand U4872 (N_4872,N_1124,N_256);
and U4873 (N_4873,N_2321,N_829);
and U4874 (N_4874,N_370,N_1726);
nor U4875 (N_4875,N_774,N_1491);
nor U4876 (N_4876,N_1214,N_2136);
nor U4877 (N_4877,N_205,N_545);
nor U4878 (N_4878,N_486,N_2443);
or U4879 (N_4879,N_2237,N_751);
and U4880 (N_4880,N_2397,N_1409);
or U4881 (N_4881,N_1253,N_1040);
and U4882 (N_4882,N_1270,N_1249);
or U4883 (N_4883,N_2298,N_1773);
nor U4884 (N_4884,N_307,N_1843);
or U4885 (N_4885,N_511,N_607);
nand U4886 (N_4886,N_17,N_679);
or U4887 (N_4887,N_384,N_2206);
nor U4888 (N_4888,N_784,N_533);
and U4889 (N_4889,N_787,N_826);
nand U4890 (N_4890,N_68,N_1045);
or U4891 (N_4891,N_1333,N_174);
and U4892 (N_4892,N_2403,N_526);
nor U4893 (N_4893,N_914,N_611);
and U4894 (N_4894,N_960,N_2264);
and U4895 (N_4895,N_363,N_543);
or U4896 (N_4896,N_1132,N_200);
nor U4897 (N_4897,N_1642,N_511);
or U4898 (N_4898,N_1548,N_957);
nand U4899 (N_4899,N_134,N_750);
and U4900 (N_4900,N_91,N_2114);
or U4901 (N_4901,N_1867,N_17);
or U4902 (N_4902,N_1230,N_763);
and U4903 (N_4903,N_1068,N_215);
nor U4904 (N_4904,N_1522,N_1545);
nand U4905 (N_4905,N_793,N_2166);
nand U4906 (N_4906,N_1150,N_630);
and U4907 (N_4907,N_1409,N_1846);
nand U4908 (N_4908,N_1194,N_23);
and U4909 (N_4909,N_88,N_880);
nand U4910 (N_4910,N_1265,N_1962);
and U4911 (N_4911,N_837,N_669);
nand U4912 (N_4912,N_789,N_84);
nor U4913 (N_4913,N_1098,N_2250);
or U4914 (N_4914,N_766,N_2184);
and U4915 (N_4915,N_1487,N_312);
and U4916 (N_4916,N_1550,N_1480);
nand U4917 (N_4917,N_1716,N_164);
nor U4918 (N_4918,N_1234,N_2441);
nor U4919 (N_4919,N_1741,N_1009);
nand U4920 (N_4920,N_1420,N_1367);
or U4921 (N_4921,N_5,N_1877);
or U4922 (N_4922,N_976,N_2210);
and U4923 (N_4923,N_437,N_210);
nor U4924 (N_4924,N_1628,N_1512);
and U4925 (N_4925,N_1922,N_762);
and U4926 (N_4926,N_752,N_913);
and U4927 (N_4927,N_2429,N_1296);
and U4928 (N_4928,N_61,N_677);
nand U4929 (N_4929,N_2235,N_2033);
nand U4930 (N_4930,N_1819,N_1888);
nor U4931 (N_4931,N_213,N_140);
nor U4932 (N_4932,N_1108,N_1546);
nand U4933 (N_4933,N_526,N_798);
nand U4934 (N_4934,N_1198,N_104);
or U4935 (N_4935,N_1421,N_1637);
nor U4936 (N_4936,N_2282,N_1655);
and U4937 (N_4937,N_515,N_2188);
nand U4938 (N_4938,N_1098,N_660);
and U4939 (N_4939,N_375,N_2111);
nand U4940 (N_4940,N_1885,N_536);
nor U4941 (N_4941,N_1199,N_303);
and U4942 (N_4942,N_2047,N_2289);
and U4943 (N_4943,N_835,N_722);
nand U4944 (N_4944,N_2147,N_349);
nand U4945 (N_4945,N_1704,N_1878);
or U4946 (N_4946,N_1172,N_685);
nor U4947 (N_4947,N_2398,N_1189);
or U4948 (N_4948,N_343,N_1060);
nor U4949 (N_4949,N_726,N_1874);
xnor U4950 (N_4950,N_224,N_17);
or U4951 (N_4951,N_1649,N_834);
nor U4952 (N_4952,N_1367,N_95);
nand U4953 (N_4953,N_321,N_1842);
and U4954 (N_4954,N_1646,N_1810);
and U4955 (N_4955,N_1237,N_142);
and U4956 (N_4956,N_490,N_1207);
and U4957 (N_4957,N_1761,N_683);
nand U4958 (N_4958,N_1612,N_205);
nand U4959 (N_4959,N_2339,N_771);
or U4960 (N_4960,N_1549,N_2327);
and U4961 (N_4961,N_928,N_1943);
nor U4962 (N_4962,N_594,N_1030);
nor U4963 (N_4963,N_1991,N_690);
nor U4964 (N_4964,N_1369,N_2328);
and U4965 (N_4965,N_2251,N_597);
and U4966 (N_4966,N_1822,N_577);
and U4967 (N_4967,N_2128,N_1374);
or U4968 (N_4968,N_205,N_1917);
or U4969 (N_4969,N_1253,N_1022);
or U4970 (N_4970,N_660,N_2401);
or U4971 (N_4971,N_390,N_1733);
and U4972 (N_4972,N_1098,N_451);
nand U4973 (N_4973,N_2004,N_1859);
and U4974 (N_4974,N_2374,N_1296);
and U4975 (N_4975,N_62,N_414);
nand U4976 (N_4976,N_86,N_1221);
and U4977 (N_4977,N_1674,N_924);
or U4978 (N_4978,N_1093,N_288);
and U4979 (N_4979,N_2390,N_605);
nor U4980 (N_4980,N_181,N_1423);
nor U4981 (N_4981,N_226,N_578);
or U4982 (N_4982,N_49,N_148);
or U4983 (N_4983,N_1570,N_1569);
or U4984 (N_4984,N_326,N_1068);
or U4985 (N_4985,N_2100,N_1377);
nor U4986 (N_4986,N_2024,N_2401);
or U4987 (N_4987,N_607,N_1995);
or U4988 (N_4988,N_1434,N_2145);
and U4989 (N_4989,N_219,N_2392);
or U4990 (N_4990,N_533,N_226);
nand U4991 (N_4991,N_2392,N_2166);
and U4992 (N_4992,N_1524,N_806);
nand U4993 (N_4993,N_454,N_1390);
or U4994 (N_4994,N_2256,N_1561);
nand U4995 (N_4995,N_35,N_1893);
nand U4996 (N_4996,N_410,N_1150);
and U4997 (N_4997,N_392,N_813);
or U4998 (N_4998,N_122,N_1124);
or U4999 (N_4999,N_521,N_192);
nor UO_0 (O_0,N_4834,N_3533);
or UO_1 (O_1,N_4678,N_3629);
and UO_2 (O_2,N_4145,N_2501);
or UO_3 (O_3,N_3025,N_4195);
nand UO_4 (O_4,N_4887,N_4572);
and UO_5 (O_5,N_4861,N_3468);
or UO_6 (O_6,N_4634,N_2732);
nor UO_7 (O_7,N_2749,N_2822);
or UO_8 (O_8,N_2776,N_4260);
nand UO_9 (O_9,N_4730,N_2726);
or UO_10 (O_10,N_2773,N_2711);
nand UO_11 (O_11,N_3740,N_3159);
nor UO_12 (O_12,N_4284,N_3434);
nor UO_13 (O_13,N_4690,N_3443);
nand UO_14 (O_14,N_3510,N_3771);
and UO_15 (O_15,N_3950,N_3382);
nor UO_16 (O_16,N_3422,N_3268);
or UO_17 (O_17,N_4362,N_2622);
and UO_18 (O_18,N_3602,N_3305);
nor UO_19 (O_19,N_4103,N_3912);
and UO_20 (O_20,N_3776,N_4123);
nor UO_21 (O_21,N_4386,N_4297);
and UO_22 (O_22,N_2793,N_3779);
and UO_23 (O_23,N_4261,N_2670);
nand UO_24 (O_24,N_4240,N_3562);
nor UO_25 (O_25,N_4280,N_4767);
nand UO_26 (O_26,N_3398,N_2795);
nand UO_27 (O_27,N_4543,N_4869);
and UO_28 (O_28,N_4442,N_3316);
or UO_29 (O_29,N_4712,N_3707);
or UO_30 (O_30,N_2993,N_4890);
and UO_31 (O_31,N_4631,N_2754);
nor UO_32 (O_32,N_2937,N_3481);
nand UO_33 (O_33,N_4518,N_4676);
nor UO_34 (O_34,N_3990,N_4278);
or UO_35 (O_35,N_2923,N_4725);
and UO_36 (O_36,N_3934,N_3508);
and UO_37 (O_37,N_2808,N_3983);
or UO_38 (O_38,N_2646,N_4115);
or UO_39 (O_39,N_4241,N_3081);
nand UO_40 (O_40,N_4455,N_3825);
or UO_41 (O_41,N_4481,N_3631);
nor UO_42 (O_42,N_4614,N_4065);
nand UO_43 (O_43,N_4342,N_4387);
or UO_44 (O_44,N_2511,N_3675);
and UO_45 (O_45,N_2772,N_3910);
or UO_46 (O_46,N_4794,N_2794);
and UO_47 (O_47,N_2908,N_3194);
or UO_48 (O_48,N_4658,N_2882);
and UO_49 (O_49,N_3109,N_2917);
and UO_50 (O_50,N_4050,N_4265);
nor UO_51 (O_51,N_3251,N_2959);
or UO_52 (O_52,N_4618,N_3748);
and UO_53 (O_53,N_4480,N_4648);
nor UO_54 (O_54,N_4713,N_4469);
and UO_55 (O_55,N_4812,N_3969);
and UO_56 (O_56,N_4149,N_4765);
or UO_57 (O_57,N_4445,N_4701);
nor UO_58 (O_58,N_3522,N_4853);
nand UO_59 (O_59,N_2892,N_3186);
nand UO_60 (O_60,N_2720,N_4569);
and UO_61 (O_61,N_3125,N_3790);
nand UO_62 (O_62,N_4894,N_3977);
nor UO_63 (O_63,N_4356,N_2978);
nor UO_64 (O_64,N_2943,N_3826);
nand UO_65 (O_65,N_4844,N_2747);
or UO_66 (O_66,N_3551,N_4972);
nand UO_67 (O_67,N_2944,N_4256);
nor UO_68 (O_68,N_3304,N_2583);
or UO_69 (O_69,N_4860,N_3603);
nand UO_70 (O_70,N_4392,N_4757);
or UO_71 (O_71,N_3648,N_2832);
and UO_72 (O_72,N_3700,N_2939);
nand UO_73 (O_73,N_4580,N_2748);
and UO_74 (O_74,N_2687,N_2784);
or UO_75 (O_75,N_2607,N_3015);
nand UO_76 (O_76,N_4929,N_3764);
nor UO_77 (O_77,N_2759,N_3732);
or UO_78 (O_78,N_3894,N_3737);
nor UO_79 (O_79,N_4277,N_4693);
or UO_80 (O_80,N_4177,N_3957);
and UO_81 (O_81,N_3860,N_3730);
or UO_82 (O_82,N_4340,N_3307);
and UO_83 (O_83,N_3247,N_3936);
or UO_84 (O_84,N_4209,N_2842);
nor UO_85 (O_85,N_2510,N_3663);
and UO_86 (O_86,N_4804,N_3710);
and UO_87 (O_87,N_2914,N_4573);
nand UO_88 (O_88,N_2904,N_4083);
nor UO_89 (O_89,N_3375,N_2922);
or UO_90 (O_90,N_3529,N_3590);
and UO_91 (O_91,N_2810,N_3412);
and UO_92 (O_92,N_3691,N_2535);
nor UO_93 (O_93,N_3350,N_4621);
or UO_94 (O_94,N_3497,N_2552);
and UO_95 (O_95,N_3038,N_3727);
nor UO_96 (O_96,N_3788,N_3199);
and UO_97 (O_97,N_3649,N_3587);
or UO_98 (O_98,N_4399,N_2990);
or UO_99 (O_99,N_2651,N_4506);
or UO_100 (O_100,N_3334,N_3113);
and UO_101 (O_101,N_3645,N_2644);
nor UO_102 (O_102,N_4396,N_3023);
nand UO_103 (O_103,N_4944,N_3890);
nand UO_104 (O_104,N_4069,N_4743);
nand UO_105 (O_105,N_3408,N_3426);
or UO_106 (O_106,N_2568,N_3415);
xnor UO_107 (O_107,N_4248,N_3839);
nor UO_108 (O_108,N_4684,N_3827);
nand UO_109 (O_109,N_3488,N_4276);
nor UO_110 (O_110,N_4092,N_4322);
and UO_111 (O_111,N_4670,N_4601);
nor UO_112 (O_112,N_3107,N_4541);
nor UO_113 (O_113,N_3406,N_3692);
or UO_114 (O_114,N_3173,N_2717);
and UO_115 (O_115,N_3665,N_3420);
nand UO_116 (O_116,N_4892,N_2742);
or UO_117 (O_117,N_4779,N_2879);
and UO_118 (O_118,N_2980,N_3428);
or UO_119 (O_119,N_4872,N_4237);
nor UO_120 (O_120,N_2721,N_3227);
nor UO_121 (O_121,N_4933,N_2603);
nand UO_122 (O_122,N_2734,N_2513);
nand UO_123 (O_123,N_4525,N_4491);
nor UO_124 (O_124,N_4023,N_3623);
and UO_125 (O_125,N_3136,N_4918);
nand UO_126 (O_126,N_3859,N_2750);
nor UO_127 (O_127,N_3365,N_2530);
nand UO_128 (O_128,N_4903,N_4110);
nand UO_129 (O_129,N_4514,N_4413);
nor UO_130 (O_130,N_4497,N_3117);
nand UO_131 (O_131,N_3254,N_4797);
and UO_132 (O_132,N_3168,N_4321);
nand UO_133 (O_133,N_2637,N_3698);
and UO_134 (O_134,N_4020,N_4215);
nor UO_135 (O_135,N_4363,N_3457);
nand UO_136 (O_136,N_4568,N_4874);
and UO_137 (O_137,N_4666,N_4250);
and UO_138 (O_138,N_4963,N_4347);
nand UO_139 (O_139,N_4435,N_4727);
or UO_140 (O_140,N_4979,N_4964);
nor UO_141 (O_141,N_4637,N_2640);
or UO_142 (O_142,N_3638,N_4734);
or UO_143 (O_143,N_2969,N_3592);
nor UO_144 (O_144,N_2692,N_3051);
or UO_145 (O_145,N_3848,N_4883);
and UO_146 (O_146,N_3861,N_3042);
nand UO_147 (O_147,N_4345,N_4711);
nand UO_148 (O_148,N_3058,N_4859);
nand UO_149 (O_149,N_3405,N_3364);
nand UO_150 (O_150,N_4432,N_4117);
and UO_151 (O_151,N_4788,N_3271);
nand UO_152 (O_152,N_4315,N_3011);
nor UO_153 (O_153,N_4243,N_3699);
nor UO_154 (O_154,N_3110,N_2785);
or UO_155 (O_155,N_3013,N_4875);
and UO_156 (O_156,N_4778,N_4041);
nor UO_157 (O_157,N_2960,N_3755);
nand UO_158 (O_158,N_4820,N_4594);
or UO_159 (O_159,N_4077,N_3913);
nand UO_160 (O_160,N_4755,N_3244);
or UO_161 (O_161,N_4370,N_3981);
or UO_162 (O_162,N_3132,N_4738);
and UO_163 (O_163,N_4681,N_2824);
and UO_164 (O_164,N_3725,N_3817);
nand UO_165 (O_165,N_4987,N_3879);
nor UO_166 (O_166,N_4792,N_4045);
nand UO_167 (O_167,N_3763,N_3616);
nand UO_168 (O_168,N_4367,N_2590);
nand UO_169 (O_169,N_2517,N_4512);
or UO_170 (O_170,N_4203,N_3226);
nand UO_171 (O_171,N_3252,N_4624);
or UO_172 (O_172,N_3272,N_4784);
nand UO_173 (O_173,N_3267,N_4805);
nor UO_174 (O_174,N_3031,N_3193);
and UO_175 (O_175,N_2727,N_4246);
and UO_176 (O_176,N_2952,N_2587);
nor UO_177 (O_177,N_3442,N_3701);
or UO_178 (O_178,N_2696,N_3141);
nor UO_179 (O_179,N_4638,N_4070);
and UO_180 (O_180,N_2838,N_4511);
nor UO_181 (O_181,N_3309,N_4978);
and UO_182 (O_182,N_3397,N_4592);
nor UO_183 (O_183,N_3404,N_4208);
and UO_184 (O_184,N_3782,N_3487);
or UO_185 (O_185,N_3403,N_3430);
or UO_186 (O_186,N_4324,N_3362);
nand UO_187 (O_187,N_4305,N_3739);
and UO_188 (O_188,N_2573,N_3972);
nand UO_189 (O_189,N_4080,N_4732);
nand UO_190 (O_190,N_3312,N_3248);
nor UO_191 (O_191,N_4244,N_3906);
nor UO_192 (O_192,N_4575,N_2859);
nor UO_193 (O_193,N_4206,N_3997);
or UO_194 (O_194,N_2841,N_4338);
nand UO_195 (O_195,N_3232,N_4059);
nor UO_196 (O_196,N_4312,N_2507);
and UO_197 (O_197,N_4960,N_4218);
nor UO_198 (O_198,N_4896,N_4949);
nor UO_199 (O_199,N_3045,N_2712);
xor UO_200 (O_200,N_4194,N_2611);
nand UO_201 (O_201,N_4611,N_3466);
nor UO_202 (O_202,N_4966,N_3564);
and UO_203 (O_203,N_3575,N_4990);
nor UO_204 (O_204,N_2694,N_4422);
and UO_205 (O_205,N_3578,N_3810);
or UO_206 (O_206,N_4482,N_3891);
and UO_207 (O_207,N_3261,N_4040);
nor UO_208 (O_208,N_3995,N_4102);
nor UO_209 (O_209,N_4810,N_3467);
and UO_210 (O_210,N_2845,N_4968);
nand UO_211 (O_211,N_3588,N_4210);
or UO_212 (O_212,N_4505,N_4709);
or UO_213 (O_213,N_4122,N_2666);
nor UO_214 (O_214,N_4426,N_4078);
nand UO_215 (O_215,N_3235,N_4807);
or UO_216 (O_216,N_3625,N_3841);
and UO_217 (O_217,N_4971,N_4938);
and UO_218 (O_218,N_4381,N_3477);
or UO_219 (O_219,N_4851,N_3148);
or UO_220 (O_220,N_3265,N_4551);
or UO_221 (O_221,N_3020,N_4831);
or UO_222 (O_222,N_3077,N_4689);
nor UO_223 (O_223,N_4908,N_3862);
and UO_224 (O_224,N_4329,N_4477);
nor UO_225 (O_225,N_4721,N_4119);
and UO_226 (O_226,N_4073,N_2868);
nor UO_227 (O_227,N_3293,N_3274);
and UO_228 (O_228,N_3565,N_3703);
nand UO_229 (O_229,N_2782,N_3231);
and UO_230 (O_230,N_3242,N_3536);
or UO_231 (O_231,N_3035,N_2738);
nor UO_232 (O_232,N_3968,N_2804);
nor UO_233 (O_233,N_2522,N_4028);
nor UO_234 (O_234,N_4052,N_4888);
nor UO_235 (O_235,N_4744,N_3353);
nor UO_236 (O_236,N_3804,N_3808);
nor UO_237 (O_237,N_2902,N_2958);
and UO_238 (O_238,N_3402,N_4054);
or UO_239 (O_239,N_3577,N_3925);
and UO_240 (O_240,N_3853,N_2988);
nor UO_241 (O_241,N_4382,N_2893);
nand UO_242 (O_242,N_2817,N_4610);
nor UO_243 (O_243,N_3517,N_4925);
and UO_244 (O_244,N_4954,N_3880);
and UO_245 (O_245,N_4704,N_4848);
nor UO_246 (O_246,N_3160,N_2688);
nor UO_247 (O_247,N_3881,N_2968);
nand UO_248 (O_248,N_3731,N_3607);
nor UO_249 (O_249,N_3935,N_4801);
nor UO_250 (O_250,N_3133,N_3651);
or UO_251 (O_251,N_4120,N_3153);
or UO_252 (O_252,N_3769,N_4891);
nand UO_253 (O_253,N_4969,N_4644);
or UO_254 (O_254,N_3294,N_2894);
and UO_255 (O_255,N_4427,N_4733);
and UO_256 (O_256,N_3180,N_4942);
nand UO_257 (O_257,N_4595,N_4556);
or UO_258 (O_258,N_4316,N_3531);
and UO_259 (O_259,N_4475,N_4563);
nand UO_260 (O_260,N_2570,N_3974);
or UO_261 (O_261,N_3473,N_4991);
or UO_262 (O_262,N_4548,N_3303);
or UO_263 (O_263,N_4341,N_2864);
nand UO_264 (O_264,N_2581,N_3067);
nor UO_265 (O_265,N_3851,N_3844);
nor UO_266 (O_266,N_2661,N_4444);
and UO_267 (O_267,N_3451,N_2675);
nand UO_268 (O_268,N_4574,N_3854);
and UO_269 (O_269,N_4053,N_2627);
nor UO_270 (O_270,N_2563,N_4346);
and UO_271 (O_271,N_2950,N_4313);
nor UO_272 (O_272,N_4048,N_3465);
and UO_273 (O_273,N_2986,N_3483);
and UO_274 (O_274,N_3181,N_3905);
nand UO_275 (O_275,N_3095,N_2617);
and UO_276 (O_276,N_4953,N_2531);
and UO_277 (O_277,N_3920,N_4291);
or UO_278 (O_278,N_2874,N_3805);
or UO_279 (O_279,N_3144,N_4682);
and UO_280 (O_280,N_4554,N_4759);
or UO_281 (O_281,N_3016,N_4795);
nand UO_282 (O_282,N_3973,N_3681);
nor UO_283 (O_283,N_3801,N_4602);
nor UO_284 (O_284,N_2946,N_4479);
nand UO_285 (O_285,N_3438,N_3347);
and UO_286 (O_286,N_3351,N_4714);
or UO_287 (O_287,N_3253,N_4635);
and UO_288 (O_288,N_3018,N_3407);
nor UO_289 (O_289,N_3676,N_4438);
nand UO_290 (O_290,N_2545,N_4143);
nor UO_291 (O_291,N_2788,N_4327);
and UO_292 (O_292,N_4959,N_4472);
or UO_293 (O_293,N_2885,N_4636);
and UO_294 (O_294,N_3360,N_3535);
and UO_295 (O_295,N_4656,N_4688);
and UO_296 (O_296,N_2610,N_4881);
or UO_297 (O_297,N_3878,N_2709);
or UO_298 (O_298,N_3734,N_2777);
nor UO_299 (O_299,N_2848,N_3902);
and UO_300 (O_300,N_2998,N_4290);
nor UO_301 (O_301,N_3646,N_3705);
and UO_302 (O_302,N_2502,N_3876);
nor UO_303 (O_303,N_2537,N_3236);
and UO_304 (O_304,N_3993,N_3680);
nand UO_305 (O_305,N_3204,N_2828);
nor UO_306 (O_306,N_2903,N_4016);
nand UO_307 (O_307,N_3938,N_3918);
xnor UO_308 (O_308,N_3059,N_3728);
nor UO_309 (O_309,N_3091,N_3778);
nor UO_310 (O_310,N_3520,N_4623);
nor UO_311 (O_311,N_4526,N_3257);
or UO_312 (O_312,N_3342,N_3435);
and UO_313 (O_313,N_3514,N_4478);
nor UO_314 (O_314,N_2628,N_4952);
and UO_315 (O_315,N_4036,N_4532);
and UO_316 (O_316,N_3084,N_3384);
and UO_317 (O_317,N_4660,N_3399);
or UO_318 (O_318,N_4947,N_4153);
nand UO_319 (O_319,N_3014,N_4588);
nand UO_320 (O_320,N_3752,N_4373);
nor UO_321 (O_321,N_4997,N_4409);
nor UO_322 (O_322,N_3119,N_4184);
and UO_323 (O_323,N_2999,N_2798);
and UO_324 (O_324,N_4451,N_4965);
nor UO_325 (O_325,N_4895,N_3439);
nor UO_326 (O_326,N_4406,N_4371);
nor UO_327 (O_327,N_2542,N_3992);
nor UO_328 (O_328,N_4547,N_2555);
or UO_329 (O_329,N_2602,N_3389);
or UO_330 (O_330,N_3945,N_4458);
and UO_331 (O_331,N_4946,N_2786);
or UO_332 (O_332,N_4360,N_4450);
nor UO_333 (O_333,N_3916,N_4741);
nor UO_334 (O_334,N_4641,N_4893);
or UO_335 (O_335,N_4950,N_3417);
and UO_336 (O_336,N_3583,N_3987);
nor UO_337 (O_337,N_4369,N_2559);
nor UO_338 (O_338,N_3197,N_4948);
and UO_339 (O_339,N_2899,N_4198);
nor UO_340 (O_340,N_3370,N_2609);
and UO_341 (O_341,N_4590,N_4131);
and UO_342 (O_342,N_3846,N_4380);
nor UO_343 (O_343,N_4441,N_4084);
and UO_344 (O_344,N_2733,N_2895);
nor UO_345 (O_345,N_4420,N_3156);
nor UO_346 (O_346,N_4228,N_4695);
and UO_347 (O_347,N_4286,N_2789);
nor UO_348 (O_348,N_4783,N_3696);
nor UO_349 (O_349,N_3873,N_4263);
and UO_350 (O_350,N_4005,N_2612);
nor UO_351 (O_351,N_4484,N_2929);
or UO_352 (O_352,N_4106,N_4113);
or UO_353 (O_353,N_4565,N_3953);
nand UO_354 (O_354,N_2920,N_3462);
or UO_355 (O_355,N_3746,N_4545);
and UO_356 (O_356,N_3470,N_4232);
nor UO_357 (O_357,N_4060,N_3431);
nor UO_358 (O_358,N_4379,N_4091);
nand UO_359 (O_359,N_3621,N_4809);
and UO_360 (O_360,N_2553,N_2839);
and UO_361 (O_361,N_2608,N_3620);
and UO_362 (O_362,N_3581,N_4354);
or UO_363 (O_363,N_4366,N_3856);
nor UO_364 (O_364,N_4298,N_3246);
and UO_365 (O_365,N_4747,N_4417);
nand UO_366 (O_366,N_3030,N_3530);
nand UO_367 (O_367,N_4283,N_3440);
or UO_368 (O_368,N_3758,N_2807);
and UO_369 (O_369,N_4372,N_3955);
and UO_370 (O_370,N_3541,N_3026);
nand UO_371 (O_371,N_4819,N_3669);
or UO_372 (O_372,N_3151,N_3986);
and UO_373 (O_373,N_4473,N_4527);
nand UO_374 (O_374,N_4633,N_3793);
nor UO_375 (O_375,N_4943,N_2774);
or UO_376 (O_376,N_4748,N_2702);
nor UO_377 (O_377,N_3172,N_3206);
nand UO_378 (O_378,N_3777,N_3374);
and UO_379 (O_379,N_3177,N_4133);
or UO_380 (O_380,N_2953,N_2569);
nand UO_381 (O_381,N_2560,N_3062);
nand UO_382 (O_382,N_3065,N_4761);
and UO_383 (O_383,N_3256,N_3459);
and UO_384 (O_384,N_4351,N_3114);
nor UO_385 (O_385,N_3500,N_3589);
and UO_386 (O_386,N_4095,N_4410);
and UO_387 (O_387,N_2698,N_2906);
and UO_388 (O_388,N_3927,N_4032);
and UO_389 (O_389,N_3509,N_4097);
nand UO_390 (O_390,N_4447,N_4937);
nand UO_391 (O_391,N_4815,N_3070);
and UO_392 (O_392,N_3970,N_3798);
and UO_393 (O_393,N_2757,N_3917);
or UO_394 (O_394,N_4668,N_2714);
or UO_395 (O_395,N_2858,N_3321);
or UO_396 (O_396,N_4607,N_4308);
and UO_397 (O_397,N_2974,N_4156);
or UO_398 (O_398,N_3893,N_4552);
and UO_399 (O_399,N_3836,N_2585);
and UO_400 (O_400,N_4287,N_4296);
nor UO_401 (O_401,N_3167,N_3689);
or UO_402 (O_402,N_4255,N_4567);
nand UO_403 (O_403,N_3505,N_3032);
nand UO_404 (O_404,N_3243,N_3750);
or UO_405 (O_405,N_3495,N_4295);
or UO_406 (O_406,N_3259,N_3909);
or UO_407 (O_407,N_3693,N_4501);
nand UO_408 (O_408,N_4980,N_3108);
nand UO_409 (O_409,N_4817,N_3840);
or UO_410 (O_410,N_2663,N_2532);
nand UO_411 (O_411,N_2775,N_3656);
or UO_412 (O_412,N_2557,N_4796);
and UO_413 (O_413,N_2991,N_2586);
nand UO_414 (O_414,N_2592,N_3868);
or UO_415 (O_415,N_4742,N_3219);
nor UO_416 (O_416,N_4021,N_2865);
and UO_417 (O_417,N_4856,N_4047);
nor UO_418 (O_418,N_3496,N_3498);
nor UO_419 (O_419,N_4583,N_4847);
nand UO_420 (O_420,N_3928,N_3223);
and UO_421 (O_421,N_4079,N_3301);
and UO_422 (O_422,N_3571,N_3474);
and UO_423 (O_423,N_3083,N_4221);
nand UO_424 (O_424,N_4174,N_2673);
or UO_425 (O_425,N_4886,N_4495);
and UO_426 (O_426,N_3743,N_4806);
and UO_427 (O_427,N_3331,N_4018);
nor UO_428 (O_428,N_4829,N_4104);
nand UO_429 (O_429,N_4616,N_2996);
or UO_430 (O_430,N_3056,N_3744);
nor UO_431 (O_431,N_2928,N_2870);
nand UO_432 (O_432,N_2708,N_3661);
nor UO_433 (O_433,N_3677,N_3096);
nand UO_434 (O_434,N_3295,N_2689);
nand UO_435 (O_435,N_3239,N_3019);
and UO_436 (O_436,N_2728,N_3877);
nand UO_437 (O_437,N_2915,N_3076);
nor UO_438 (O_438,N_2938,N_2704);
nand UO_439 (O_439,N_4919,N_4772);
or UO_440 (O_440,N_2731,N_4273);
nor UO_441 (O_441,N_4775,N_3548);
nand UO_442 (O_442,N_3636,N_4694);
or UO_443 (O_443,N_3525,N_3341);
nand UO_444 (O_444,N_4125,N_4605);
or UO_445 (O_445,N_3952,N_2942);
and UO_446 (O_446,N_4416,N_3574);
nor UO_447 (O_447,N_2825,N_3277);
nor UO_448 (O_448,N_2884,N_4500);
nor UO_449 (O_449,N_3174,N_2554);
nor UO_450 (O_450,N_3637,N_3947);
nand UO_451 (O_451,N_3073,N_3523);
xor UO_452 (O_452,N_4650,N_4314);
or UO_453 (O_453,N_3780,N_3086);
nand UO_454 (O_454,N_3066,N_4604);
nand UO_455 (O_455,N_3998,N_3209);
and UO_456 (O_456,N_4109,N_3685);
or UO_457 (O_457,N_2664,N_3075);
xor UO_458 (O_458,N_4723,N_2931);
or UO_459 (O_459,N_3895,N_2621);
nand UO_460 (O_460,N_4173,N_2964);
nand UO_461 (O_461,N_2769,N_4803);
nand UO_462 (O_462,N_2796,N_4646);
nor UO_463 (O_463,N_2719,N_4663);
and UO_464 (O_464,N_3245,N_3175);
or UO_465 (O_465,N_4285,N_4385);
nor UO_466 (O_466,N_4171,N_4503);
and UO_467 (O_467,N_2681,N_3584);
nand UO_468 (O_468,N_3325,N_4516);
and UO_469 (O_469,N_3544,N_4266);
xor UO_470 (O_470,N_4087,N_4499);
or UO_471 (O_471,N_2768,N_2618);
and UO_472 (O_472,N_2600,N_3356);
or UO_473 (O_473,N_3189,N_3711);
or UO_474 (O_474,N_3889,N_4696);
or UO_475 (O_475,N_3619,N_3105);
nor UO_476 (O_476,N_2652,N_4201);
and UO_477 (O_477,N_2659,N_4967);
and UO_478 (O_478,N_3214,N_2843);
and UO_479 (O_479,N_2705,N_2629);
or UO_480 (O_480,N_4686,N_4566);
or UO_481 (O_481,N_3432,N_3504);
or UO_482 (O_482,N_4930,N_4973);
and UO_483 (O_483,N_4745,N_3543);
and UO_484 (O_484,N_2597,N_3088);
or UO_485 (O_485,N_2576,N_2926);
and UO_486 (O_486,N_2655,N_4231);
or UO_487 (O_487,N_4075,N_4530);
nand UO_488 (O_488,N_4632,N_3220);
or UO_489 (O_489,N_4722,N_4425);
nand UO_490 (O_490,N_2525,N_4835);
nor UO_491 (O_491,N_4076,N_3785);
nand UO_492 (O_492,N_3831,N_4271);
nand UO_493 (O_493,N_3756,N_3511);
nand UO_494 (O_494,N_2976,N_3400);
nand UO_495 (O_495,N_3326,N_4724);
or UO_496 (O_496,N_3445,N_3958);
or UO_497 (O_497,N_4220,N_2911);
or UO_498 (O_498,N_4845,N_3116);
nand UO_499 (O_499,N_4880,N_3857);
or UO_500 (O_500,N_4222,N_4300);
or UO_501 (O_501,N_3716,N_4651);
and UO_502 (O_502,N_2872,N_4234);
or UO_503 (O_503,N_3709,N_4365);
or UO_504 (O_504,N_3410,N_3729);
nand UO_505 (O_505,N_3796,N_2827);
nor UO_506 (O_506,N_2580,N_4498);
or UO_507 (O_507,N_4043,N_3639);
nor UO_508 (O_508,N_2620,N_3287);
or UO_509 (O_509,N_4657,N_4825);
nand UO_510 (O_510,N_3628,N_4957);
or UO_511 (O_511,N_3102,N_3482);
or UO_512 (O_512,N_4598,N_4649);
or UO_513 (O_513,N_2818,N_2746);
and UO_514 (O_514,N_3299,N_4798);
and UO_515 (O_515,N_4331,N_4816);
nor UO_516 (O_516,N_3413,N_4769);
and UO_517 (O_517,N_4911,N_4328);
or UO_518 (O_518,N_3464,N_4443);
nor UO_519 (O_519,N_2765,N_4787);
and UO_520 (O_520,N_2605,N_3212);
and UO_521 (O_521,N_2589,N_2933);
nand UO_522 (O_522,N_4175,N_3372);
or UO_523 (O_523,N_3753,N_3178);
nor UO_524 (O_524,N_3322,N_3492);
and UO_525 (O_525,N_3939,N_2575);
or UO_526 (O_526,N_4517,N_4985);
or UO_527 (O_527,N_4528,N_3850);
nor UO_528 (O_528,N_2797,N_4096);
nor UO_529 (O_529,N_3593,N_4901);
or UO_530 (O_530,N_4061,N_3617);
nand UO_531 (O_531,N_3933,N_3339);
or UO_532 (O_532,N_3213,N_2853);
xor UO_533 (O_533,N_4873,N_3956);
nor UO_534 (O_534,N_3211,N_4910);
and UO_535 (O_535,N_4672,N_2534);
nor UO_536 (O_536,N_4008,N_2812);
or UO_537 (O_537,N_2584,N_3323);
and UO_538 (O_538,N_2840,N_4166);
or UO_539 (O_539,N_2814,N_4151);
and UO_540 (O_540,N_3207,N_4193);
or UO_541 (O_541,N_3931,N_4114);
nand UO_542 (O_542,N_4414,N_4229);
or UO_543 (O_543,N_2697,N_4852);
and UO_544 (O_544,N_3647,N_2561);
and UO_545 (O_545,N_3866,N_4025);
or UO_546 (O_546,N_4746,N_2703);
xnor UO_547 (O_547,N_4453,N_4214);
nor UO_548 (O_548,N_3005,N_2515);
nor UO_549 (O_549,N_4669,N_4192);
and UO_550 (O_550,N_3269,N_3152);
nor UO_551 (O_551,N_3635,N_3262);
and UO_552 (O_552,N_4034,N_3140);
or UO_553 (O_553,N_4703,N_4301);
and UO_554 (O_554,N_3237,N_4389);
nand UO_555 (O_555,N_2809,N_4715);
or UO_556 (O_556,N_2737,N_4487);
or UO_557 (O_557,N_3715,N_3683);
and UO_558 (O_558,N_2548,N_4507);
and UO_559 (O_559,N_3567,N_3937);
nor UO_560 (O_560,N_4586,N_3988);
and UO_561 (O_561,N_4773,N_3418);
nor UO_562 (O_562,N_3068,N_2710);
or UO_563 (O_563,N_4200,N_4584);
or UO_564 (O_564,N_4926,N_3358);
or UO_565 (O_565,N_4223,N_4405);
or UO_566 (O_566,N_3039,N_3800);
and UO_567 (O_567,N_3518,N_4233);
nor UO_568 (O_568,N_3870,N_2685);
and UO_569 (O_569,N_4905,N_3554);
and UO_570 (O_570,N_2521,N_4159);
nor UO_571 (O_571,N_3130,N_3634);
nor UO_572 (O_572,N_4553,N_4729);
or UO_573 (O_573,N_4306,N_3849);
nor UO_574 (O_574,N_2863,N_3369);
nand UO_575 (O_575,N_3555,N_4249);
or UO_576 (O_576,N_3923,N_2925);
or UO_577 (O_577,N_2723,N_4502);
and UO_578 (O_578,N_3192,N_4155);
and UO_579 (O_579,N_2970,N_3599);
or UO_580 (O_580,N_3965,N_4400);
and UO_581 (O_581,N_4840,N_2979);
or UO_582 (O_582,N_3191,N_4253);
and UO_583 (O_583,N_4270,N_4419);
or UO_584 (O_584,N_4375,N_4026);
nand UO_585 (O_585,N_3004,N_2615);
nor UO_586 (O_586,N_4627,N_4509);
and UO_587 (O_587,N_2551,N_2634);
nand UO_588 (O_588,N_2955,N_4421);
and UO_589 (O_589,N_3922,N_3319);
and UO_590 (O_590,N_4494,N_2833);
or UO_591 (O_591,N_3914,N_2668);
or UO_592 (O_592,N_2791,N_4202);
nor UO_593 (O_593,N_4088,N_3225);
or UO_594 (O_594,N_2546,N_3915);
nor UO_595 (O_595,N_2803,N_4108);
or UO_596 (O_596,N_3361,N_4466);
nand UO_597 (O_597,N_2558,N_2657);
or UO_598 (O_598,N_4105,N_3783);
xnor UO_599 (O_599,N_3882,N_4533);
or UO_600 (O_600,N_3537,N_4067);
and UO_601 (O_601,N_3611,N_4619);
or UO_602 (O_602,N_4754,N_4538);
nand UO_603 (O_603,N_4062,N_3770);
or UO_604 (O_604,N_4140,N_4428);
nand UO_605 (O_605,N_4353,N_4599);
or UO_606 (O_606,N_3486,N_4247);
nand UO_607 (O_607,N_4643,N_4864);
or UO_608 (O_608,N_2891,N_3673);
nand UO_609 (O_609,N_2636,N_2861);
and UO_610 (O_610,N_4698,N_3494);
nand UO_611 (O_611,N_3092,N_3932);
nor UO_612 (O_612,N_4557,N_2678);
or UO_613 (O_613,N_2852,N_4654);
nor UO_614 (O_614,N_3886,N_3155);
and UO_615 (O_615,N_2745,N_3142);
and UO_616 (O_616,N_3813,N_2730);
nand UO_617 (O_617,N_4936,N_2860);
nor UO_618 (O_618,N_3164,N_3097);
nand UO_619 (O_619,N_4549,N_3888);
nand UO_620 (O_620,N_4368,N_2982);
or UO_621 (O_621,N_2799,N_4982);
nand UO_622 (O_622,N_3962,N_3802);
nor UO_623 (O_623,N_4677,N_4626);
xnor UO_624 (O_624,N_3184,N_4093);
and UO_625 (O_625,N_4989,N_2954);
or UO_626 (O_626,N_3786,N_3311);
nand UO_627 (O_627,N_2625,N_4617);
or UO_628 (O_628,N_4913,N_2846);
or UO_629 (O_629,N_4928,N_4309);
nor UO_630 (O_630,N_2718,N_4531);
and UO_631 (O_631,N_3208,N_3823);
nand UO_632 (O_632,N_4042,N_4924);
nor UO_633 (O_633,N_3821,N_4988);
and UO_634 (O_634,N_4161,N_2880);
and UO_635 (O_635,N_2665,N_3867);
or UO_636 (O_636,N_3749,N_4673);
nand UO_637 (O_637,N_4010,N_4188);
nor UO_638 (O_638,N_4534,N_2516);
or UO_639 (O_639,N_4292,N_3491);
nor UO_640 (O_640,N_3614,N_3328);
or UO_641 (O_641,N_3344,N_3640);
and UO_642 (O_642,N_4555,N_4986);
or UO_643 (O_643,N_2813,N_2601);
nor UO_644 (O_644,N_2977,N_4536);
nand UO_645 (O_645,N_4390,N_3718);
nor UO_646 (O_646,N_3241,N_4003);
nand UO_647 (O_647,N_3885,N_3061);
nand UO_648 (O_648,N_3052,N_3022);
nand UO_649 (O_649,N_4158,N_4217);
and UO_650 (O_650,N_3157,N_4303);
or UO_651 (O_651,N_4415,N_3774);
nand UO_652 (O_652,N_3205,N_3908);
nor UO_653 (O_653,N_3573,N_4033);
and UO_654 (O_654,N_3566,N_2764);
nand UO_655 (O_655,N_4813,N_4049);
nor UO_656 (O_656,N_3216,N_3453);
or UO_657 (O_657,N_3686,N_3006);
nand UO_658 (O_658,N_2577,N_3812);
nor UO_659 (O_659,N_2806,N_3697);
nand UO_660 (O_660,N_3528,N_3195);
or UO_661 (O_661,N_4776,N_4763);
nand UO_662 (O_662,N_3754,N_3332);
or UO_663 (O_663,N_2690,N_3290);
or UO_664 (O_664,N_2512,N_3318);
or UO_665 (O_665,N_4996,N_4705);
or UO_666 (O_666,N_3424,N_4474);
and UO_667 (O_667,N_3919,N_3447);
nor UO_668 (O_668,N_2743,N_4251);
nor UO_669 (O_669,N_4814,N_3991);
and UO_670 (O_670,N_3871,N_2643);
or UO_671 (O_671,N_2951,N_3792);
or UO_672 (O_672,N_3594,N_4935);
nand UO_673 (O_673,N_3896,N_2631);
nand UO_674 (O_674,N_3306,N_4863);
or UO_675 (O_675,N_4608,N_4542);
or UO_676 (O_676,N_3655,N_4708);
or UO_677 (O_677,N_3448,N_3721);
and UO_678 (O_678,N_3506,N_2679);
and UO_679 (O_679,N_4781,N_4094);
nand UO_680 (O_680,N_3276,N_4766);
nor UO_681 (O_681,N_3653,N_3690);
nor UO_682 (O_682,N_4827,N_4204);
nor UO_683 (O_683,N_3672,N_3662);
nor UO_684 (O_684,N_3660,N_3024);
and UO_685 (O_685,N_4398,N_3559);
or UO_686 (O_686,N_4391,N_2889);
nor UO_687 (O_687,N_2888,N_3280);
or UO_688 (O_688,N_3082,N_4189);
or UO_689 (O_689,N_3540,N_3377);
and UO_690 (O_690,N_4383,N_4927);
nor UO_691 (O_691,N_4822,N_2756);
nand UO_692 (O_692,N_3847,N_4307);
nand UO_693 (O_693,N_4163,N_4606);
and UO_694 (O_694,N_4697,N_3501);
or UO_695 (O_695,N_4661,N_4793);
nand UO_696 (O_696,N_4157,N_3093);
nor UO_697 (O_697,N_3485,N_4970);
nand UO_698 (O_698,N_4540,N_3940);
and UO_699 (O_699,N_4357,N_3446);
nor UO_700 (O_700,N_4152,N_4652);
nor UO_701 (O_701,N_2829,N_3230);
and UO_702 (O_702,N_2820,N_4378);
nand UO_703 (O_703,N_3806,N_3532);
nor UO_704 (O_704,N_4437,N_3179);
and UO_705 (O_705,N_2881,N_2966);
nand UO_706 (O_706,N_3714,N_2624);
and UO_707 (O_707,N_3210,N_3822);
and UO_708 (O_708,N_4850,N_2910);
or UO_709 (O_709,N_4339,N_3218);
nor UO_710 (O_710,N_3668,N_3391);
and UO_711 (O_711,N_3137,N_2751);
or UO_712 (O_712,N_2680,N_4854);
nor UO_713 (O_713,N_3475,N_3297);
nand UO_714 (O_714,N_3641,N_4216);
or UO_715 (O_715,N_3162,N_2700);
nor UO_716 (O_716,N_3708,N_3818);
or UO_717 (O_717,N_3250,N_4900);
or UO_718 (O_718,N_3138,N_4912);
and UO_719 (O_719,N_3429,N_4183);
or UO_720 (O_720,N_3512,N_3176);
nand UO_721 (O_721,N_2574,N_4139);
nor UO_722 (O_722,N_4771,N_4752);
and UO_723 (O_723,N_3388,N_3980);
and UO_724 (O_724,N_2596,N_4402);
nand UO_725 (O_725,N_4015,N_3171);
or UO_726 (O_726,N_3336,N_4112);
nand UO_727 (O_727,N_2760,N_2536);
nor UO_728 (O_728,N_4355,N_2957);
nand UO_729 (O_729,N_4167,N_3436);
nand UO_730 (O_730,N_4866,N_4024);
nand UO_731 (O_731,N_4333,N_3003);
and UO_732 (O_732,N_4332,N_3898);
or UO_733 (O_733,N_3907,N_3630);
and UO_734 (O_734,N_4035,N_4750);
nand UO_735 (O_735,N_4164,N_3874);
nor UO_736 (O_736,N_4710,N_4579);
and UO_737 (O_737,N_3057,N_3601);
or UO_738 (O_738,N_2758,N_3865);
or UO_739 (O_739,N_4081,N_3128);
nor UO_740 (O_740,N_4141,N_4504);
or UO_741 (O_741,N_4600,N_2932);
or UO_742 (O_742,N_2936,N_2752);
and UO_743 (O_743,N_2647,N_2862);
and UO_744 (O_744,N_4560,N_4558);
nor UO_745 (O_745,N_3667,N_3926);
nand UO_746 (O_746,N_3666,N_3455);
nand UO_747 (O_747,N_2667,N_3371);
or UO_748 (O_748,N_2816,N_3472);
nand UO_749 (O_749,N_4828,N_4838);
nor UO_750 (O_750,N_4335,N_2736);
nand UO_751 (O_751,N_4836,N_2847);
nand UO_752 (O_752,N_4492,N_2919);
nor UO_753 (O_753,N_3624,N_3376);
and UO_754 (O_754,N_4774,N_2632);
nand UO_755 (O_755,N_3961,N_3279);
and UO_756 (O_756,N_3330,N_2921);
or UO_757 (O_757,N_4199,N_3534);
nand UO_758 (O_758,N_3354,N_4664);
nor UO_759 (O_759,N_2724,N_3444);
and UO_760 (O_760,N_4259,N_3034);
nand UO_761 (O_761,N_2658,N_3787);
and UO_762 (O_762,N_2849,N_3949);
and UO_763 (O_763,N_3579,N_4213);
and UO_764 (O_764,N_2767,N_4897);
and UO_765 (O_765,N_3010,N_3201);
or UO_766 (O_766,N_3345,N_4326);
and UO_767 (O_767,N_3855,N_2650);
and UO_768 (O_768,N_3597,N_3314);
or UO_769 (O_769,N_4388,N_3363);
xnor UO_770 (O_770,N_4072,N_3600);
nand UO_771 (O_771,N_2606,N_4121);
nand UO_772 (O_772,N_3049,N_2565);
and UO_773 (O_773,N_4683,N_2844);
nor UO_774 (O_774,N_4434,N_3320);
and UO_775 (O_775,N_4137,N_4468);
and UO_776 (O_776,N_2518,N_2887);
and UO_777 (O_777,N_3994,N_3654);
or UO_778 (O_778,N_3270,N_3585);
nor UO_779 (O_779,N_3659,N_4529);
nor UO_780 (O_780,N_3582,N_2582);
nand UO_781 (O_781,N_4975,N_2579);
and UO_782 (O_782,N_2547,N_3921);
or UO_783 (O_783,N_4824,N_3458);
nand UO_784 (O_784,N_3979,N_3258);
and UO_785 (O_785,N_3278,N_3550);
and UO_786 (O_786,N_4154,N_3976);
nand UO_787 (O_787,N_3942,N_3622);
and UO_788 (O_788,N_4849,N_3240);
and UO_789 (O_789,N_4561,N_4082);
and UO_790 (O_790,N_4884,N_4768);
nor UO_791 (O_791,N_3381,N_3869);
nand UO_792 (O_792,N_4719,N_2940);
and UO_793 (O_793,N_4994,N_3000);
or UO_794 (O_794,N_3129,N_4984);
nand UO_795 (O_795,N_4483,N_4842);
nor UO_796 (O_796,N_4830,N_3609);
nor UO_797 (O_797,N_3644,N_4236);
or UO_798 (O_798,N_3954,N_4961);
nor UO_799 (O_799,N_3797,N_4889);
xor UO_800 (O_800,N_2856,N_4993);
nand UO_801 (O_801,N_4281,N_4974);
and UO_802 (O_802,N_4485,N_3028);
nand UO_803 (O_803,N_4800,N_4448);
nand UO_804 (O_804,N_3724,N_3104);
nor UO_805 (O_805,N_4085,N_2695);
nand UO_806 (O_806,N_3337,N_4977);
and UO_807 (O_807,N_4433,N_3292);
nor UO_808 (O_808,N_4224,N_3224);
nor UO_809 (O_809,N_3229,N_2543);
or UO_810 (O_810,N_4037,N_4000);
nor UO_811 (O_811,N_2541,N_3127);
or UO_812 (O_812,N_3903,N_4685);
and UO_813 (O_813,N_3423,N_4124);
and UO_814 (O_814,N_4515,N_2744);
or UO_815 (O_815,N_2778,N_4429);
or UO_816 (O_816,N_4162,N_4239);
nor UO_817 (O_817,N_3338,N_4907);
and UO_818 (O_818,N_4962,N_3735);
nor UO_819 (O_819,N_3608,N_4449);
nor UO_820 (O_820,N_4323,N_3984);
nand UO_821 (O_821,N_4242,N_4692);
xor UO_822 (O_822,N_2905,N_4107);
or UO_823 (O_823,N_3985,N_3327);
nor UO_824 (O_824,N_2595,N_3386);
nor UO_825 (O_825,N_4645,N_4521);
nand UO_826 (O_826,N_2763,N_3315);
or UO_827 (O_827,N_3664,N_4334);
or UO_828 (O_828,N_4496,N_2591);
nor UO_829 (O_829,N_4983,N_3288);
nand UO_830 (O_830,N_4764,N_3249);
or UO_831 (O_831,N_4411,N_4404);
or UO_832 (O_832,N_2684,N_3145);
nor UO_833 (O_833,N_3355,N_3557);
and UO_834 (O_834,N_3832,N_3618);
or UO_835 (O_835,N_4299,N_4998);
nand UO_836 (O_836,N_4620,N_4951);
and UO_837 (O_837,N_3480,N_4802);
and UO_838 (O_838,N_3765,N_3704);
or UO_839 (O_839,N_3379,N_3041);
and UO_840 (O_840,N_2912,N_3215);
nand UO_841 (O_841,N_4257,N_2802);
nor UO_842 (O_842,N_4030,N_4544);
and UO_843 (O_843,N_3427,N_2594);
xor UO_844 (O_844,N_3335,N_4613);
and UO_845 (O_845,N_4885,N_4004);
and UO_846 (O_846,N_4187,N_3348);
or UO_847 (O_847,N_2706,N_4914);
and UO_848 (O_848,N_2524,N_2567);
or UO_849 (O_849,N_2604,N_4348);
and UO_850 (O_850,N_4629,N_3872);
nor UO_851 (O_851,N_2509,N_4205);
nand UO_852 (O_852,N_2588,N_3479);
and UO_853 (O_853,N_4293,N_4615);
and UO_854 (O_854,N_4452,N_3340);
or UO_855 (O_855,N_2779,N_4142);
or UO_856 (O_856,N_4230,N_2837);
and UO_857 (O_857,N_2642,N_2755);
nor UO_858 (O_858,N_4737,N_4490);
or UO_859 (O_859,N_4808,N_3037);
nor UO_860 (O_860,N_3687,N_3165);
and UO_861 (O_861,N_2916,N_3586);
nor UO_862 (O_862,N_3393,N_2800);
and UO_863 (O_863,N_3115,N_2770);
nand UO_864 (O_864,N_2701,N_4728);
and UO_865 (O_865,N_4051,N_3054);
or UO_866 (O_866,N_3642,N_4870);
and UO_867 (O_867,N_3838,N_4846);
nor UO_868 (O_868,N_4019,N_2676);
nand UO_869 (O_869,N_3460,N_4570);
nand UO_870 (O_870,N_2792,N_4101);
nand UO_871 (O_871,N_3717,N_4463);
and UO_872 (O_872,N_4350,N_3814);
nor UO_873 (O_873,N_3263,N_3558);
nor UO_874 (O_874,N_3545,N_4780);
nand UO_875 (O_875,N_4749,N_3373);
or UO_876 (O_876,N_3284,N_2877);
or UO_877 (O_877,N_3064,N_3198);
nand UO_878 (O_878,N_4288,N_3807);
nand UO_879 (O_879,N_3188,N_2857);
and UO_880 (O_880,N_4252,N_3329);
or UO_881 (O_881,N_2686,N_4691);
nand UO_882 (O_882,N_4628,N_4510);
nor UO_883 (O_883,N_3454,N_4915);
or UO_884 (O_884,N_2735,N_3433);
and UO_885 (O_885,N_2713,N_2975);
nor UO_886 (O_886,N_3471,N_3598);
or UO_887 (O_887,N_4958,N_2593);
or UO_888 (O_888,N_4882,N_2729);
or UO_889 (O_889,N_4170,N_3829);
or UO_890 (O_890,N_4439,N_3733);
or UO_891 (O_891,N_3411,N_3103);
nand UO_892 (O_892,N_4336,N_2805);
nor UO_893 (O_893,N_3833,N_4017);
nand UO_894 (O_894,N_3048,N_2526);
or UO_895 (O_895,N_2948,N_3069);
nand UO_896 (O_896,N_4238,N_4111);
or UO_897 (O_897,N_4191,N_3561);
and UO_898 (O_898,N_2540,N_4401);
or UO_899 (O_899,N_2962,N_2876);
nor UO_900 (O_900,N_4671,N_3385);
nor UO_901 (O_901,N_3343,N_3357);
nand UO_902 (O_902,N_3897,N_4011);
nand UO_903 (O_903,N_4826,N_3050);
and UO_904 (O_904,N_2983,N_2801);
nand UO_905 (O_905,N_2599,N_4358);
nor UO_906 (O_906,N_2707,N_3650);
and UO_907 (O_907,N_4007,N_3001);
or UO_908 (O_908,N_3012,N_4235);
nand UO_909 (O_909,N_4679,N_3900);
or UO_910 (O_910,N_4325,N_3392);
nor UO_911 (O_911,N_2890,N_2715);
and UO_912 (O_912,N_2662,N_4777);
or UO_913 (O_913,N_3595,N_4116);
or UO_914 (O_914,N_3378,N_4100);
or UO_915 (O_915,N_3719,N_2722);
nand UO_916 (O_916,N_3150,N_3310);
nor UO_917 (O_917,N_2869,N_2790);
nand UO_918 (O_918,N_3416,N_2815);
and UO_919 (O_919,N_3099,N_2683);
nor UO_920 (O_920,N_3080,N_3380);
nand UO_921 (O_921,N_4129,N_3147);
nand UO_922 (O_922,N_3493,N_3569);
nand UO_923 (O_923,N_3078,N_3563);
and UO_924 (O_924,N_2997,N_2529);
nor UO_925 (O_925,N_3266,N_4564);
nor UO_926 (O_926,N_4337,N_4418);
and UO_927 (O_927,N_4044,N_4546);
and UO_928 (O_928,N_3556,N_4539);
or UO_929 (O_929,N_4940,N_4408);
nor UO_930 (O_930,N_3469,N_4576);
or UO_931 (O_931,N_4535,N_4562);
and UO_932 (O_932,N_2883,N_4071);
and UO_933 (O_933,N_3282,N_2830);
and UO_934 (O_934,N_3255,N_3943);
or UO_935 (O_935,N_4945,N_4225);
nor UO_936 (O_936,N_3053,N_4289);
nand UO_937 (O_937,N_3072,N_3989);
nand UO_938 (O_938,N_3098,N_4144);
nand UO_939 (O_939,N_2930,N_3368);
nand UO_940 (O_940,N_4867,N_3911);
nand UO_941 (O_941,N_3757,N_3396);
nand UO_942 (O_942,N_2867,N_2649);
nor UO_943 (O_943,N_3060,N_3570);
nand UO_944 (O_944,N_4138,N_3499);
nand UO_945 (O_945,N_4294,N_4981);
and UO_946 (O_946,N_4879,N_3959);
nand UO_947 (O_947,N_3946,N_2766);
nand UO_948 (O_948,N_3401,N_4180);
nor UO_949 (O_949,N_4486,N_3017);
and UO_950 (O_950,N_3539,N_4904);
and UO_951 (O_951,N_4736,N_3706);
nand UO_952 (O_952,N_3087,N_3228);
and UO_953 (O_953,N_4311,N_3044);
or UO_954 (O_954,N_4148,N_4268);
nand UO_955 (O_955,N_4090,N_3170);
or UO_956 (O_956,N_3300,N_3824);
nand UO_957 (O_957,N_3203,N_3875);
nor UO_958 (O_958,N_4622,N_2613);
nand UO_959 (O_959,N_4074,N_4589);
and UO_960 (O_960,N_4818,N_3695);
or UO_961 (O_961,N_2771,N_3803);
or UO_962 (O_962,N_3154,N_2992);
or UO_963 (O_963,N_4318,N_3029);
or UO_964 (O_964,N_3901,N_3772);
and UO_965 (O_965,N_3951,N_3071);
nor UO_966 (O_966,N_3450,N_3538);
nand UO_967 (O_967,N_4361,N_4039);
and UO_968 (O_968,N_2677,N_3553);
and UO_969 (O_969,N_4196,N_3674);
or UO_970 (O_970,N_3217,N_3089);
nor UO_971 (O_971,N_3002,N_4630);
nor UO_972 (O_972,N_3843,N_3394);
nor UO_973 (O_973,N_2549,N_3040);
nand UO_974 (O_974,N_4146,N_4181);
nor UO_975 (O_975,N_3387,N_4585);
nor UO_976 (O_976,N_3852,N_4118);
and UO_977 (O_977,N_4464,N_3317);
nand UO_978 (O_978,N_3789,N_4467);
nand UO_979 (O_979,N_3346,N_4436);
or UO_980 (O_980,N_3768,N_2653);
and UO_981 (O_981,N_2641,N_3106);
nor UO_982 (O_982,N_3139,N_3333);
or UO_983 (O_983,N_3324,N_3185);
nand UO_984 (O_984,N_3694,N_3751);
nor UO_985 (O_985,N_4058,N_3572);
nand UO_986 (O_986,N_2533,N_2660);
nor UO_987 (O_987,N_2648,N_3633);
or UO_988 (O_988,N_2886,N_2834);
nor UO_989 (O_989,N_3063,N_2961);
nand UO_990 (O_990,N_2645,N_4066);
nand UO_991 (O_991,N_3169,N_3047);
xor UO_992 (O_992,N_3542,N_4412);
nand UO_993 (O_993,N_3302,N_3967);
nor UO_994 (O_994,N_3626,N_4923);
or UO_995 (O_995,N_2972,N_3264);
nor UO_996 (O_996,N_2907,N_2971);
nor UO_997 (O_997,N_2994,N_4902);
nand UO_998 (O_998,N_4457,N_3830);
nor UO_999 (O_999,N_4999,N_4593);
endmodule