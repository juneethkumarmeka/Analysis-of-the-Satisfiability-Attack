module basic_500_3000_500_60_levels_5xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_203,In_419);
and U1 (N_1,In_49,In_57);
nor U2 (N_2,In_476,In_348);
nand U3 (N_3,In_421,In_273);
nor U4 (N_4,In_136,In_343);
nor U5 (N_5,In_339,In_63);
and U6 (N_6,In_303,In_312);
nand U7 (N_7,In_7,In_200);
nor U8 (N_8,In_179,In_239);
nor U9 (N_9,In_141,In_69);
or U10 (N_10,In_415,In_199);
or U11 (N_11,In_389,In_361);
nor U12 (N_12,In_456,In_107);
nand U13 (N_13,In_326,In_87);
and U14 (N_14,In_497,In_324);
xnor U15 (N_15,In_446,In_182);
nand U16 (N_16,In_146,In_349);
and U17 (N_17,In_311,In_400);
nor U18 (N_18,In_298,In_469);
nor U19 (N_19,In_11,In_213);
and U20 (N_20,In_499,In_404);
or U21 (N_21,In_208,In_166);
nor U22 (N_22,In_186,In_309);
nor U23 (N_23,In_245,In_76);
xnor U24 (N_24,In_442,In_33);
xnor U25 (N_25,In_485,In_431);
nor U26 (N_26,In_280,In_54);
and U27 (N_27,In_1,In_114);
nand U28 (N_28,In_91,In_342);
nand U29 (N_29,In_140,In_29);
and U30 (N_30,In_392,In_51);
and U31 (N_31,In_101,In_160);
and U32 (N_32,In_109,In_444);
nand U33 (N_33,In_331,In_391);
and U34 (N_34,In_460,In_180);
nor U35 (N_35,In_484,In_15);
and U36 (N_36,In_170,In_367);
xnor U37 (N_37,In_297,In_46);
nor U38 (N_38,In_206,In_218);
nor U39 (N_39,In_489,In_375);
and U40 (N_40,In_128,In_338);
or U41 (N_41,In_435,In_441);
xor U42 (N_42,In_59,In_424);
nor U43 (N_43,In_267,In_439);
nand U44 (N_44,In_156,In_27);
xor U45 (N_45,In_426,In_32);
nor U46 (N_46,In_238,In_145);
nand U47 (N_47,In_110,In_173);
nand U48 (N_48,In_299,In_372);
nor U49 (N_49,In_482,In_0);
and U50 (N_50,N_23,In_65);
nand U51 (N_51,In_294,In_353);
nand U52 (N_52,In_39,In_6);
or U53 (N_53,In_257,In_41);
and U54 (N_54,N_37,In_20);
nand U55 (N_55,In_467,In_158);
nor U56 (N_56,N_26,In_67);
or U57 (N_57,In_210,In_346);
nor U58 (N_58,N_18,In_288);
nand U59 (N_59,In_452,In_410);
or U60 (N_60,In_261,In_73);
nor U61 (N_61,In_80,In_266);
or U62 (N_62,In_85,In_232);
or U63 (N_63,In_418,In_42);
and U64 (N_64,In_422,In_378);
nor U65 (N_65,In_117,In_58);
nand U66 (N_66,In_387,In_249);
and U67 (N_67,In_480,In_108);
nand U68 (N_68,In_293,In_328);
nand U69 (N_69,In_162,In_115);
or U70 (N_70,N_6,In_472);
nand U71 (N_71,In_366,In_398);
nand U72 (N_72,In_19,In_92);
nand U73 (N_73,In_285,In_88);
xnor U74 (N_74,In_132,In_106);
nand U75 (N_75,In_474,In_263);
nand U76 (N_76,N_12,In_171);
or U77 (N_77,In_495,In_282);
nor U78 (N_78,In_9,In_190);
nor U79 (N_79,In_151,In_194);
or U80 (N_80,In_177,In_479);
nand U81 (N_81,In_433,N_30);
or U82 (N_82,N_44,In_152);
nor U83 (N_83,In_408,In_251);
nand U84 (N_84,In_370,In_153);
and U85 (N_85,In_413,In_229);
nor U86 (N_86,In_248,In_374);
and U87 (N_87,In_430,In_350);
nand U88 (N_88,In_473,In_79);
or U89 (N_89,In_345,In_385);
or U90 (N_90,In_130,In_258);
xor U91 (N_91,In_211,In_16);
or U92 (N_92,In_149,N_39);
xnor U93 (N_93,In_191,In_207);
nand U94 (N_94,In_230,In_143);
nor U95 (N_95,In_195,In_397);
or U96 (N_96,In_97,In_71);
and U97 (N_97,In_93,In_396);
and U98 (N_98,In_302,In_490);
xnor U99 (N_99,In_260,In_368);
and U100 (N_100,In_333,In_355);
or U101 (N_101,In_187,In_75);
and U102 (N_102,In_226,In_196);
nor U103 (N_103,In_23,In_21);
nand U104 (N_104,In_70,In_221);
nor U105 (N_105,In_255,In_197);
and U106 (N_106,In_82,In_376);
nor U107 (N_107,In_77,N_1);
or U108 (N_108,In_487,N_67);
or U109 (N_109,In_364,In_465);
or U110 (N_110,In_118,N_43);
and U111 (N_111,N_53,N_33);
or U112 (N_112,In_235,In_250);
xor U113 (N_113,In_244,In_236);
and U114 (N_114,In_332,In_185);
nand U115 (N_115,In_443,In_329);
nand U116 (N_116,In_55,In_278);
or U117 (N_117,In_135,N_10);
nand U118 (N_118,In_60,In_379);
nand U119 (N_119,In_386,In_181);
or U120 (N_120,In_215,N_49);
and U121 (N_121,In_129,In_306);
nor U122 (N_122,In_31,In_287);
and U123 (N_123,In_100,In_466);
or U124 (N_124,In_253,In_411);
nor U125 (N_125,N_50,N_93);
nand U126 (N_126,In_102,N_66);
or U127 (N_127,In_256,In_459);
nand U128 (N_128,N_14,In_72);
nand U129 (N_129,N_82,In_274);
and U130 (N_130,In_395,N_62);
or U131 (N_131,In_453,In_390);
nand U132 (N_132,In_341,In_14);
and U133 (N_133,In_159,N_96);
nand U134 (N_134,N_32,In_279);
and U135 (N_135,N_40,In_481);
or U136 (N_136,In_323,In_315);
nand U137 (N_137,N_13,In_157);
or U138 (N_138,In_24,In_74);
or U139 (N_139,In_313,N_64);
nand U140 (N_140,In_103,In_125);
or U141 (N_141,In_436,In_425);
nand U142 (N_142,In_448,In_254);
xnor U143 (N_143,In_420,In_275);
and U144 (N_144,N_92,In_493);
nand U145 (N_145,In_336,In_131);
nand U146 (N_146,In_454,In_407);
and U147 (N_147,In_35,In_308);
and U148 (N_148,N_15,N_20);
xor U149 (N_149,In_119,In_150);
and U150 (N_150,In_458,N_88);
xnor U151 (N_151,In_50,In_432);
nor U152 (N_152,In_296,In_330);
or U153 (N_153,In_95,N_59);
nor U154 (N_154,In_5,N_76);
nand U155 (N_155,N_89,N_7);
nor U156 (N_156,N_83,N_123);
nand U157 (N_157,N_90,N_127);
nand U158 (N_158,N_35,In_219);
or U159 (N_159,In_335,In_96);
nand U160 (N_160,N_54,In_234);
xor U161 (N_161,In_227,N_46);
or U162 (N_162,In_305,In_295);
nor U163 (N_163,In_222,N_100);
nor U164 (N_164,In_310,N_58);
and U165 (N_165,In_449,N_138);
nand U166 (N_166,N_122,N_126);
nor U167 (N_167,In_137,N_8);
xor U168 (N_168,In_98,In_445);
nor U169 (N_169,In_317,N_129);
and U170 (N_170,N_85,In_401);
nor U171 (N_171,In_17,N_69);
nand U172 (N_172,N_140,In_428);
nor U173 (N_173,In_47,In_344);
nor U174 (N_174,N_98,In_112);
and U175 (N_175,N_145,In_365);
and U176 (N_176,In_247,N_80);
xor U177 (N_177,In_45,In_123);
or U178 (N_178,N_41,In_417);
nand U179 (N_179,In_381,In_167);
nand U180 (N_180,N_125,N_81);
nor U181 (N_181,N_143,In_252);
nand U182 (N_182,In_168,In_455);
or U183 (N_183,N_113,In_8);
and U184 (N_184,In_43,In_155);
or U185 (N_185,In_44,N_139);
and U186 (N_186,In_10,N_136);
or U187 (N_187,N_146,In_62);
nand U188 (N_188,In_204,In_144);
or U189 (N_189,In_380,N_134);
xor U190 (N_190,In_37,In_268);
or U191 (N_191,In_165,In_3);
nand U192 (N_192,N_60,In_53);
and U193 (N_193,In_447,N_61);
nand U194 (N_194,N_107,In_347);
nor U195 (N_195,In_192,In_154);
nand U196 (N_196,In_105,In_269);
nor U197 (N_197,In_371,In_318);
nor U198 (N_198,N_135,In_496);
nand U199 (N_199,N_4,In_405);
and U200 (N_200,In_147,N_45);
and U201 (N_201,N_0,In_22);
nor U202 (N_202,In_99,In_120);
or U203 (N_203,In_450,In_325);
nor U204 (N_204,In_412,N_133);
nor U205 (N_205,In_286,In_126);
and U206 (N_206,N_29,In_40);
and U207 (N_207,N_108,In_242);
and U208 (N_208,In_356,N_180);
and U209 (N_209,In_139,N_179);
nor U210 (N_210,In_277,In_104);
or U211 (N_211,In_178,In_90);
nand U212 (N_212,In_265,In_81);
nand U213 (N_213,N_103,In_363);
or U214 (N_214,N_16,N_21);
xor U215 (N_215,N_84,In_264);
or U216 (N_216,N_112,In_61);
or U217 (N_217,In_18,In_13);
nand U218 (N_218,In_327,In_461);
and U219 (N_219,In_468,In_176);
or U220 (N_220,In_172,N_141);
or U221 (N_221,N_102,In_133);
nand U222 (N_222,In_111,N_194);
and U223 (N_223,N_91,In_188);
xor U224 (N_224,N_147,In_307);
nand U225 (N_225,In_233,N_74);
xor U226 (N_226,N_144,In_66);
or U227 (N_227,In_351,In_369);
and U228 (N_228,In_457,In_217);
or U229 (N_229,In_406,In_321);
nand U230 (N_230,In_174,In_113);
nand U231 (N_231,N_158,N_106);
nand U232 (N_232,In_36,In_440);
and U233 (N_233,In_228,N_110);
or U234 (N_234,In_394,N_199);
and U235 (N_235,N_181,In_201);
or U236 (N_236,In_427,N_68);
and U237 (N_237,In_270,In_464);
nand U238 (N_238,In_290,N_155);
nand U239 (N_239,N_118,N_27);
or U240 (N_240,N_131,N_99);
nand U241 (N_241,N_153,N_128);
xnor U242 (N_242,In_12,N_5);
nand U243 (N_243,In_246,N_191);
and U244 (N_244,In_383,In_451);
or U245 (N_245,In_360,N_114);
and U246 (N_246,N_195,N_132);
nand U247 (N_247,N_188,N_48);
nand U248 (N_248,N_111,In_475);
xor U249 (N_249,N_154,In_189);
nor U250 (N_250,N_206,In_216);
nand U251 (N_251,In_354,In_30);
and U252 (N_252,In_434,In_300);
and U253 (N_253,N_75,In_134);
nor U254 (N_254,N_215,In_423);
nor U255 (N_255,In_488,N_198);
xnor U256 (N_256,N_234,In_220);
nand U257 (N_257,N_177,N_17);
nor U258 (N_258,N_163,In_402);
xnor U259 (N_259,N_42,N_216);
nand U260 (N_260,N_238,N_200);
nor U261 (N_261,N_51,N_34);
xor U262 (N_262,In_163,N_63);
nand U263 (N_263,N_189,N_52);
and U264 (N_264,N_220,In_198);
or U265 (N_265,N_36,In_78);
and U266 (N_266,In_292,N_165);
and U267 (N_267,N_94,N_65);
and U268 (N_268,In_304,In_301);
or U269 (N_269,In_340,N_222);
and U270 (N_270,In_283,In_86);
or U271 (N_271,In_470,In_281);
or U272 (N_272,In_409,N_116);
xor U273 (N_273,In_34,In_477);
nor U274 (N_274,In_382,N_170);
nor U275 (N_275,In_212,In_384);
nand U276 (N_276,N_225,In_357);
nor U277 (N_277,In_403,In_52);
nand U278 (N_278,In_142,In_463);
and U279 (N_279,In_316,In_291);
and U280 (N_280,In_122,N_237);
nor U281 (N_281,N_185,N_9);
or U282 (N_282,In_56,N_167);
nand U283 (N_283,N_242,N_47);
xnor U284 (N_284,N_79,N_183);
nor U285 (N_285,N_164,N_160);
nand U286 (N_286,N_224,N_223);
nand U287 (N_287,In_214,N_78);
or U288 (N_288,N_117,N_187);
nand U289 (N_289,N_207,N_232);
xor U290 (N_290,In_438,N_202);
xnor U291 (N_291,In_486,N_56);
xnor U292 (N_292,N_156,In_388);
nor U293 (N_293,N_70,In_225);
nor U294 (N_294,In_184,N_24);
nor U295 (N_295,N_105,N_115);
nor U296 (N_296,In_183,N_229);
xor U297 (N_297,N_159,In_314);
or U298 (N_298,N_205,N_176);
xor U299 (N_299,N_28,In_416);
and U300 (N_300,In_161,In_223);
nor U301 (N_301,In_373,N_269);
xnor U302 (N_302,N_19,N_152);
or U303 (N_303,N_22,N_231);
nand U304 (N_304,N_11,N_250);
nand U305 (N_305,N_137,In_124);
nand U306 (N_306,N_246,N_260);
and U307 (N_307,N_284,N_287);
or U308 (N_308,N_213,In_337);
and U309 (N_309,In_202,N_262);
nor U310 (N_310,N_203,N_55);
nand U311 (N_311,N_173,N_174);
xor U312 (N_312,In_276,N_193);
nand U313 (N_313,N_278,N_275);
nand U314 (N_314,N_263,In_414);
or U315 (N_315,N_124,In_492);
nor U316 (N_316,N_291,In_38);
xnor U317 (N_317,In_193,N_182);
or U318 (N_318,N_204,In_498);
nand U319 (N_319,N_212,N_130);
and U320 (N_320,In_272,N_192);
and U321 (N_321,N_119,In_399);
nand U322 (N_322,N_253,N_261);
or U323 (N_323,N_101,In_28);
nand U324 (N_324,N_217,In_84);
and U325 (N_325,N_244,N_211);
and U326 (N_326,N_273,N_218);
nand U327 (N_327,N_190,N_274);
and U328 (N_328,N_264,N_162);
nand U329 (N_329,N_248,In_89);
nor U330 (N_330,In_334,In_175);
or U331 (N_331,N_57,N_295);
and U332 (N_332,In_2,N_25);
xor U333 (N_333,N_172,In_462);
nand U334 (N_334,N_161,In_359);
or U335 (N_335,N_97,In_358);
nand U336 (N_336,In_352,N_209);
nand U337 (N_337,N_236,N_281);
nand U338 (N_338,In_320,In_478);
or U339 (N_339,N_270,In_271);
and U340 (N_340,N_184,N_233);
or U341 (N_341,N_265,In_241);
and U342 (N_342,N_230,N_228);
nor U343 (N_343,N_294,N_31);
and U344 (N_344,N_95,N_277);
nor U345 (N_345,N_226,In_289);
and U346 (N_346,N_247,N_235);
nand U347 (N_347,N_297,In_121);
or U348 (N_348,N_121,In_362);
nor U349 (N_349,N_149,In_64);
or U350 (N_350,N_290,N_349);
nand U351 (N_351,N_221,N_339);
or U352 (N_352,In_483,N_298);
xnor U353 (N_353,N_293,In_94);
nand U354 (N_354,N_309,In_116);
or U355 (N_355,N_296,N_307);
and U356 (N_356,In_471,In_127);
and U357 (N_357,N_344,In_148);
and U358 (N_358,N_322,N_208);
xor U359 (N_359,In_164,N_186);
and U360 (N_360,N_157,N_227);
nand U361 (N_361,N_109,N_201);
and U362 (N_362,In_240,N_314);
nor U363 (N_363,In_224,In_205);
nand U364 (N_364,In_491,N_310);
or U365 (N_365,N_169,N_299);
or U366 (N_366,N_303,N_286);
nor U367 (N_367,N_2,N_245);
or U368 (N_368,N_257,In_393);
or U369 (N_369,N_3,N_289);
or U370 (N_370,N_325,N_341);
and U371 (N_371,N_142,In_68);
or U372 (N_372,N_288,N_306);
and U373 (N_373,N_327,In_243);
or U374 (N_374,N_87,N_268);
or U375 (N_375,N_318,N_171);
nor U376 (N_376,N_319,N_340);
xnor U377 (N_377,In_284,In_259);
nand U378 (N_378,N_283,N_324);
or U379 (N_379,In_83,N_346);
or U380 (N_380,N_239,In_377);
and U381 (N_381,N_241,N_120);
or U382 (N_382,N_334,N_321);
or U383 (N_383,N_285,N_266);
nor U384 (N_384,N_343,N_342);
nand U385 (N_385,N_271,N_258);
or U386 (N_386,N_151,N_243);
nand U387 (N_387,N_254,N_276);
and U388 (N_388,N_312,N_335);
or U389 (N_389,In_138,In_169);
nor U390 (N_390,N_302,N_175);
nand U391 (N_391,N_168,N_256);
and U392 (N_392,N_104,N_308);
nand U393 (N_393,N_336,N_300);
nor U394 (N_394,In_319,N_348);
nor U395 (N_395,In_262,N_347);
nand U396 (N_396,In_26,N_280);
nor U397 (N_397,In_231,N_73);
or U398 (N_398,N_214,N_148);
and U399 (N_399,N_328,N_219);
or U400 (N_400,N_361,N_392);
and U401 (N_401,N_345,N_369);
nor U402 (N_402,N_393,N_384);
nand U403 (N_403,N_368,N_380);
or U404 (N_404,N_375,N_399);
nand U405 (N_405,N_330,N_353);
or U406 (N_406,N_355,N_150);
xnor U407 (N_407,In_48,N_255);
or U408 (N_408,In_437,N_357);
or U409 (N_409,N_383,N_367);
xnor U410 (N_410,N_364,N_398);
or U411 (N_411,N_259,N_166);
xnor U412 (N_412,In_25,N_323);
nor U413 (N_413,N_350,N_292);
and U414 (N_414,N_210,N_352);
or U415 (N_415,N_365,N_372);
nor U416 (N_416,N_390,N_272);
nand U417 (N_417,N_337,N_360);
nand U418 (N_418,N_366,N_391);
and U419 (N_419,N_326,N_316);
and U420 (N_420,N_386,N_377);
and U421 (N_421,N_362,N_267);
nand U422 (N_422,N_351,N_240);
or U423 (N_423,N_354,N_329);
and U424 (N_424,In_322,N_389);
or U425 (N_425,N_77,N_396);
or U426 (N_426,N_313,N_197);
or U427 (N_427,N_395,N_356);
and U428 (N_428,N_397,In_209);
and U429 (N_429,N_394,N_38);
or U430 (N_430,In_4,N_381);
and U431 (N_431,N_379,N_252);
or U432 (N_432,N_333,N_178);
nor U433 (N_433,N_385,N_376);
and U434 (N_434,N_387,N_388);
or U435 (N_435,N_370,N_373);
nand U436 (N_436,N_301,N_282);
nor U437 (N_437,N_382,N_304);
nor U438 (N_438,N_371,In_429);
or U439 (N_439,N_359,N_249);
and U440 (N_440,N_251,In_237);
or U441 (N_441,N_311,N_331);
or U442 (N_442,N_72,N_358);
xor U443 (N_443,N_71,N_338);
xor U444 (N_444,N_279,In_494);
nor U445 (N_445,N_363,N_317);
or U446 (N_446,N_196,N_86);
and U447 (N_447,N_332,N_315);
nand U448 (N_448,N_305,N_320);
nor U449 (N_449,N_378,N_374);
or U450 (N_450,N_404,N_407);
nand U451 (N_451,N_412,N_425);
nor U452 (N_452,N_441,N_430);
nand U453 (N_453,N_431,N_447);
nand U454 (N_454,N_413,N_448);
xor U455 (N_455,N_439,N_408);
or U456 (N_456,N_438,N_409);
or U457 (N_457,N_415,N_401);
and U458 (N_458,N_428,N_406);
nor U459 (N_459,N_427,N_426);
or U460 (N_460,N_435,N_443);
and U461 (N_461,N_422,N_423);
nor U462 (N_462,N_416,N_440);
and U463 (N_463,N_429,N_419);
xnor U464 (N_464,N_442,N_411);
nand U465 (N_465,N_418,N_432);
nor U466 (N_466,N_400,N_421);
nand U467 (N_467,N_437,N_420);
nand U468 (N_468,N_433,N_449);
nor U469 (N_469,N_444,N_403);
nor U470 (N_470,N_410,N_414);
nand U471 (N_471,N_417,N_405);
or U472 (N_472,N_402,N_436);
nor U473 (N_473,N_424,N_446);
nand U474 (N_474,N_445,N_434);
nor U475 (N_475,N_440,N_435);
or U476 (N_476,N_413,N_409);
xor U477 (N_477,N_426,N_448);
and U478 (N_478,N_408,N_443);
nor U479 (N_479,N_420,N_414);
or U480 (N_480,N_442,N_400);
and U481 (N_481,N_420,N_422);
xnor U482 (N_482,N_447,N_419);
or U483 (N_483,N_427,N_401);
nand U484 (N_484,N_438,N_440);
nor U485 (N_485,N_444,N_442);
nor U486 (N_486,N_407,N_436);
xor U487 (N_487,N_401,N_421);
xor U488 (N_488,N_419,N_402);
nand U489 (N_489,N_411,N_403);
nor U490 (N_490,N_400,N_420);
nand U491 (N_491,N_423,N_421);
or U492 (N_492,N_444,N_409);
nor U493 (N_493,N_427,N_423);
xor U494 (N_494,N_401,N_448);
and U495 (N_495,N_448,N_436);
nand U496 (N_496,N_430,N_407);
xor U497 (N_497,N_439,N_449);
nor U498 (N_498,N_437,N_412);
and U499 (N_499,N_444,N_424);
nor U500 (N_500,N_453,N_466);
xnor U501 (N_501,N_486,N_450);
nand U502 (N_502,N_482,N_460);
xor U503 (N_503,N_476,N_494);
nor U504 (N_504,N_457,N_477);
nor U505 (N_505,N_461,N_479);
and U506 (N_506,N_459,N_464);
xnor U507 (N_507,N_483,N_451);
and U508 (N_508,N_465,N_480);
nor U509 (N_509,N_487,N_462);
nor U510 (N_510,N_467,N_485);
nand U511 (N_511,N_495,N_468);
and U512 (N_512,N_499,N_496);
nor U513 (N_513,N_478,N_481);
or U514 (N_514,N_458,N_469);
nor U515 (N_515,N_454,N_463);
nand U516 (N_516,N_490,N_489);
xor U517 (N_517,N_473,N_491);
nor U518 (N_518,N_452,N_455);
and U519 (N_519,N_456,N_471);
nor U520 (N_520,N_497,N_470);
nor U521 (N_521,N_474,N_493);
and U522 (N_522,N_492,N_472);
xnor U523 (N_523,N_498,N_488);
and U524 (N_524,N_475,N_484);
and U525 (N_525,N_475,N_457);
and U526 (N_526,N_494,N_460);
and U527 (N_527,N_489,N_475);
or U528 (N_528,N_466,N_450);
nand U529 (N_529,N_480,N_481);
and U530 (N_530,N_469,N_475);
nor U531 (N_531,N_486,N_496);
or U532 (N_532,N_483,N_484);
or U533 (N_533,N_456,N_460);
nor U534 (N_534,N_487,N_481);
nor U535 (N_535,N_489,N_476);
or U536 (N_536,N_478,N_452);
and U537 (N_537,N_453,N_485);
nor U538 (N_538,N_497,N_479);
and U539 (N_539,N_490,N_459);
xor U540 (N_540,N_469,N_465);
and U541 (N_541,N_455,N_463);
nand U542 (N_542,N_493,N_456);
nor U543 (N_543,N_487,N_465);
or U544 (N_544,N_491,N_454);
and U545 (N_545,N_478,N_455);
and U546 (N_546,N_470,N_462);
and U547 (N_547,N_467,N_499);
nor U548 (N_548,N_477,N_470);
or U549 (N_549,N_473,N_476);
xor U550 (N_550,N_520,N_543);
nor U551 (N_551,N_516,N_505);
nor U552 (N_552,N_518,N_529);
nor U553 (N_553,N_524,N_510);
or U554 (N_554,N_509,N_508);
nor U555 (N_555,N_503,N_500);
or U556 (N_556,N_546,N_539);
and U557 (N_557,N_526,N_547);
nor U558 (N_558,N_541,N_548);
nor U559 (N_559,N_502,N_519);
and U560 (N_560,N_528,N_512);
or U561 (N_561,N_527,N_536);
and U562 (N_562,N_533,N_506);
and U563 (N_563,N_549,N_525);
or U564 (N_564,N_522,N_514);
nor U565 (N_565,N_545,N_534);
nand U566 (N_566,N_542,N_517);
xor U567 (N_567,N_531,N_523);
and U568 (N_568,N_504,N_507);
nand U569 (N_569,N_537,N_532);
and U570 (N_570,N_511,N_540);
or U571 (N_571,N_521,N_501);
nand U572 (N_572,N_544,N_535);
nor U573 (N_573,N_538,N_515);
nand U574 (N_574,N_513,N_530);
nand U575 (N_575,N_539,N_541);
nand U576 (N_576,N_510,N_533);
or U577 (N_577,N_525,N_506);
and U578 (N_578,N_511,N_549);
nor U579 (N_579,N_529,N_500);
and U580 (N_580,N_521,N_509);
nand U581 (N_581,N_516,N_535);
xnor U582 (N_582,N_524,N_513);
xnor U583 (N_583,N_507,N_541);
xor U584 (N_584,N_516,N_527);
xnor U585 (N_585,N_518,N_528);
nor U586 (N_586,N_537,N_523);
or U587 (N_587,N_536,N_531);
and U588 (N_588,N_537,N_516);
or U589 (N_589,N_515,N_548);
nor U590 (N_590,N_536,N_521);
nand U591 (N_591,N_517,N_512);
nor U592 (N_592,N_517,N_538);
or U593 (N_593,N_543,N_525);
nand U594 (N_594,N_518,N_500);
and U595 (N_595,N_502,N_518);
and U596 (N_596,N_524,N_503);
xor U597 (N_597,N_546,N_511);
or U598 (N_598,N_519,N_536);
or U599 (N_599,N_544,N_514);
nor U600 (N_600,N_560,N_579);
nor U601 (N_601,N_597,N_570);
nor U602 (N_602,N_588,N_556);
and U603 (N_603,N_594,N_554);
nand U604 (N_604,N_595,N_567);
or U605 (N_605,N_555,N_584);
xor U606 (N_606,N_577,N_550);
nand U607 (N_607,N_551,N_598);
xor U608 (N_608,N_580,N_592);
and U609 (N_609,N_557,N_578);
or U610 (N_610,N_562,N_574);
nor U611 (N_611,N_552,N_568);
and U612 (N_612,N_582,N_569);
and U613 (N_613,N_553,N_559);
nand U614 (N_614,N_576,N_589);
and U615 (N_615,N_587,N_591);
and U616 (N_616,N_575,N_571);
nor U617 (N_617,N_566,N_585);
or U618 (N_618,N_581,N_564);
xor U619 (N_619,N_599,N_593);
or U620 (N_620,N_586,N_573);
and U621 (N_621,N_583,N_572);
and U622 (N_622,N_565,N_561);
nor U623 (N_623,N_563,N_590);
nand U624 (N_624,N_558,N_596);
nand U625 (N_625,N_595,N_599);
xor U626 (N_626,N_553,N_594);
or U627 (N_627,N_582,N_571);
or U628 (N_628,N_594,N_570);
and U629 (N_629,N_577,N_573);
and U630 (N_630,N_569,N_598);
xnor U631 (N_631,N_575,N_581);
or U632 (N_632,N_557,N_553);
or U633 (N_633,N_566,N_595);
and U634 (N_634,N_570,N_589);
and U635 (N_635,N_589,N_599);
nand U636 (N_636,N_593,N_583);
nor U637 (N_637,N_582,N_562);
xnor U638 (N_638,N_559,N_550);
and U639 (N_639,N_567,N_575);
nand U640 (N_640,N_589,N_567);
or U641 (N_641,N_584,N_568);
nor U642 (N_642,N_551,N_587);
or U643 (N_643,N_590,N_570);
nor U644 (N_644,N_573,N_579);
and U645 (N_645,N_552,N_584);
or U646 (N_646,N_597,N_588);
or U647 (N_647,N_571,N_557);
and U648 (N_648,N_589,N_551);
nor U649 (N_649,N_597,N_564);
xnor U650 (N_650,N_608,N_639);
nor U651 (N_651,N_624,N_610);
or U652 (N_652,N_606,N_614);
xnor U653 (N_653,N_617,N_629);
nor U654 (N_654,N_605,N_625);
nor U655 (N_655,N_634,N_603);
nor U656 (N_656,N_633,N_601);
and U657 (N_657,N_649,N_641);
xnor U658 (N_658,N_602,N_609);
and U659 (N_659,N_635,N_636);
nand U660 (N_660,N_646,N_607);
xor U661 (N_661,N_615,N_628);
nand U662 (N_662,N_643,N_621);
nand U663 (N_663,N_630,N_640);
nand U664 (N_664,N_648,N_604);
and U665 (N_665,N_600,N_642);
or U666 (N_666,N_631,N_618);
and U667 (N_667,N_616,N_638);
or U668 (N_668,N_632,N_623);
nor U669 (N_669,N_622,N_647);
or U670 (N_670,N_620,N_612);
nand U671 (N_671,N_613,N_637);
or U672 (N_672,N_619,N_626);
xor U673 (N_673,N_627,N_645);
and U674 (N_674,N_611,N_644);
or U675 (N_675,N_614,N_603);
xor U676 (N_676,N_638,N_645);
and U677 (N_677,N_639,N_632);
nand U678 (N_678,N_638,N_617);
nand U679 (N_679,N_608,N_646);
or U680 (N_680,N_619,N_601);
or U681 (N_681,N_604,N_633);
and U682 (N_682,N_602,N_617);
and U683 (N_683,N_633,N_606);
nor U684 (N_684,N_641,N_620);
or U685 (N_685,N_609,N_636);
or U686 (N_686,N_636,N_618);
xor U687 (N_687,N_606,N_605);
or U688 (N_688,N_600,N_638);
nor U689 (N_689,N_636,N_610);
xnor U690 (N_690,N_637,N_628);
nor U691 (N_691,N_646,N_636);
and U692 (N_692,N_613,N_624);
and U693 (N_693,N_601,N_612);
xnor U694 (N_694,N_623,N_638);
and U695 (N_695,N_630,N_638);
or U696 (N_696,N_614,N_624);
and U697 (N_697,N_624,N_638);
and U698 (N_698,N_629,N_643);
and U699 (N_699,N_619,N_636);
xor U700 (N_700,N_694,N_693);
nor U701 (N_701,N_681,N_690);
or U702 (N_702,N_656,N_657);
nand U703 (N_703,N_670,N_689);
nand U704 (N_704,N_673,N_668);
xor U705 (N_705,N_651,N_652);
nand U706 (N_706,N_675,N_660);
nor U707 (N_707,N_671,N_659);
and U708 (N_708,N_682,N_695);
xnor U709 (N_709,N_697,N_672);
nor U710 (N_710,N_685,N_687);
or U711 (N_711,N_662,N_663);
nand U712 (N_712,N_684,N_679);
or U713 (N_713,N_686,N_664);
nand U714 (N_714,N_661,N_676);
nand U715 (N_715,N_653,N_680);
nand U716 (N_716,N_677,N_667);
or U717 (N_717,N_655,N_650);
nor U718 (N_718,N_692,N_666);
nand U719 (N_719,N_699,N_654);
nor U720 (N_720,N_688,N_691);
and U721 (N_721,N_674,N_658);
and U722 (N_722,N_698,N_669);
and U723 (N_723,N_678,N_665);
nor U724 (N_724,N_683,N_696);
nor U725 (N_725,N_697,N_661);
and U726 (N_726,N_696,N_675);
xor U727 (N_727,N_657,N_675);
nand U728 (N_728,N_655,N_675);
nor U729 (N_729,N_656,N_658);
nor U730 (N_730,N_667,N_669);
or U731 (N_731,N_659,N_653);
nand U732 (N_732,N_672,N_690);
nor U733 (N_733,N_653,N_666);
or U734 (N_734,N_664,N_691);
nor U735 (N_735,N_682,N_660);
nand U736 (N_736,N_674,N_691);
and U737 (N_737,N_664,N_650);
nor U738 (N_738,N_689,N_694);
and U739 (N_739,N_670,N_655);
nor U740 (N_740,N_676,N_666);
nand U741 (N_741,N_697,N_687);
nor U742 (N_742,N_656,N_673);
or U743 (N_743,N_659,N_696);
or U744 (N_744,N_654,N_681);
nand U745 (N_745,N_659,N_676);
or U746 (N_746,N_678,N_655);
nor U747 (N_747,N_695,N_668);
nor U748 (N_748,N_683,N_693);
nand U749 (N_749,N_691,N_672);
or U750 (N_750,N_736,N_716);
or U751 (N_751,N_734,N_749);
or U752 (N_752,N_710,N_722);
and U753 (N_753,N_747,N_735);
xnor U754 (N_754,N_719,N_709);
nor U755 (N_755,N_744,N_739);
nor U756 (N_756,N_702,N_725);
and U757 (N_757,N_721,N_714);
or U758 (N_758,N_733,N_738);
nand U759 (N_759,N_746,N_742);
and U760 (N_760,N_730,N_707);
or U761 (N_761,N_727,N_718);
nor U762 (N_762,N_706,N_720);
nor U763 (N_763,N_740,N_711);
and U764 (N_764,N_701,N_712);
or U765 (N_765,N_708,N_748);
and U766 (N_766,N_713,N_728);
nand U767 (N_767,N_723,N_726);
and U768 (N_768,N_704,N_745);
nor U769 (N_769,N_715,N_700);
or U770 (N_770,N_731,N_724);
and U771 (N_771,N_703,N_732);
xor U772 (N_772,N_737,N_743);
nor U773 (N_773,N_717,N_741);
and U774 (N_774,N_705,N_729);
nand U775 (N_775,N_718,N_704);
nand U776 (N_776,N_745,N_744);
or U777 (N_777,N_742,N_707);
nand U778 (N_778,N_720,N_702);
nand U779 (N_779,N_734,N_703);
and U780 (N_780,N_721,N_731);
nor U781 (N_781,N_710,N_715);
or U782 (N_782,N_714,N_707);
nand U783 (N_783,N_704,N_722);
nor U784 (N_784,N_730,N_706);
nor U785 (N_785,N_743,N_713);
nand U786 (N_786,N_708,N_728);
nand U787 (N_787,N_732,N_729);
nand U788 (N_788,N_713,N_739);
nor U789 (N_789,N_736,N_731);
and U790 (N_790,N_726,N_739);
nand U791 (N_791,N_713,N_747);
nor U792 (N_792,N_735,N_711);
and U793 (N_793,N_744,N_746);
xnor U794 (N_794,N_746,N_743);
nand U795 (N_795,N_723,N_725);
and U796 (N_796,N_714,N_700);
nor U797 (N_797,N_713,N_725);
nor U798 (N_798,N_742,N_715);
nor U799 (N_799,N_719,N_713);
and U800 (N_800,N_786,N_753);
or U801 (N_801,N_765,N_759);
nand U802 (N_802,N_789,N_787);
and U803 (N_803,N_782,N_758);
or U804 (N_804,N_764,N_785);
or U805 (N_805,N_756,N_781);
xor U806 (N_806,N_796,N_768);
nor U807 (N_807,N_751,N_761);
or U808 (N_808,N_755,N_788);
nand U809 (N_809,N_763,N_773);
or U810 (N_810,N_780,N_792);
or U811 (N_811,N_775,N_799);
nor U812 (N_812,N_771,N_798);
and U813 (N_813,N_770,N_769);
nand U814 (N_814,N_757,N_762);
or U815 (N_815,N_766,N_774);
nand U816 (N_816,N_776,N_794);
nor U817 (N_817,N_767,N_783);
or U818 (N_818,N_784,N_778);
nand U819 (N_819,N_760,N_754);
or U820 (N_820,N_795,N_772);
nand U821 (N_821,N_790,N_777);
nor U822 (N_822,N_797,N_750);
nand U823 (N_823,N_793,N_752);
xnor U824 (N_824,N_791,N_779);
nand U825 (N_825,N_753,N_756);
and U826 (N_826,N_763,N_774);
or U827 (N_827,N_767,N_764);
and U828 (N_828,N_781,N_785);
nor U829 (N_829,N_783,N_792);
and U830 (N_830,N_751,N_780);
nand U831 (N_831,N_793,N_756);
nand U832 (N_832,N_791,N_792);
nand U833 (N_833,N_754,N_796);
nor U834 (N_834,N_772,N_798);
xor U835 (N_835,N_798,N_775);
nor U836 (N_836,N_793,N_775);
and U837 (N_837,N_774,N_754);
nand U838 (N_838,N_772,N_779);
and U839 (N_839,N_772,N_771);
xnor U840 (N_840,N_796,N_771);
nor U841 (N_841,N_761,N_775);
and U842 (N_842,N_775,N_764);
nor U843 (N_843,N_776,N_754);
nor U844 (N_844,N_795,N_755);
nand U845 (N_845,N_755,N_778);
nand U846 (N_846,N_760,N_752);
nor U847 (N_847,N_782,N_764);
or U848 (N_848,N_794,N_753);
nor U849 (N_849,N_783,N_780);
nand U850 (N_850,N_846,N_836);
or U851 (N_851,N_839,N_842);
or U852 (N_852,N_805,N_834);
or U853 (N_853,N_826,N_820);
nor U854 (N_854,N_832,N_838);
or U855 (N_855,N_843,N_808);
xor U856 (N_856,N_827,N_831);
nor U857 (N_857,N_803,N_822);
and U858 (N_858,N_801,N_810);
and U859 (N_859,N_804,N_811);
nand U860 (N_860,N_819,N_848);
and U861 (N_861,N_828,N_802);
xor U862 (N_862,N_833,N_835);
or U863 (N_863,N_818,N_837);
or U864 (N_864,N_809,N_847);
nor U865 (N_865,N_829,N_800);
or U866 (N_866,N_813,N_807);
and U867 (N_867,N_845,N_815);
nor U868 (N_868,N_821,N_840);
and U869 (N_869,N_841,N_817);
nand U870 (N_870,N_812,N_830);
nand U871 (N_871,N_849,N_816);
nand U872 (N_872,N_844,N_824);
nand U873 (N_873,N_814,N_823);
xnor U874 (N_874,N_806,N_825);
nand U875 (N_875,N_841,N_820);
or U876 (N_876,N_846,N_801);
nor U877 (N_877,N_809,N_810);
and U878 (N_878,N_821,N_800);
nand U879 (N_879,N_822,N_820);
xor U880 (N_880,N_801,N_800);
nor U881 (N_881,N_841,N_838);
nand U882 (N_882,N_808,N_845);
and U883 (N_883,N_830,N_845);
or U884 (N_884,N_823,N_825);
or U885 (N_885,N_848,N_831);
and U886 (N_886,N_844,N_830);
and U887 (N_887,N_829,N_826);
or U888 (N_888,N_833,N_803);
nand U889 (N_889,N_811,N_809);
or U890 (N_890,N_812,N_800);
nor U891 (N_891,N_823,N_836);
or U892 (N_892,N_831,N_837);
or U893 (N_893,N_801,N_842);
nor U894 (N_894,N_842,N_831);
and U895 (N_895,N_839,N_829);
nor U896 (N_896,N_846,N_818);
or U897 (N_897,N_812,N_804);
xor U898 (N_898,N_823,N_803);
and U899 (N_899,N_840,N_817);
nand U900 (N_900,N_865,N_890);
nand U901 (N_901,N_897,N_853);
nand U902 (N_902,N_895,N_893);
or U903 (N_903,N_858,N_862);
nor U904 (N_904,N_892,N_857);
or U905 (N_905,N_866,N_898);
or U906 (N_906,N_870,N_874);
nor U907 (N_907,N_888,N_859);
or U908 (N_908,N_887,N_861);
or U909 (N_909,N_869,N_882);
or U910 (N_910,N_876,N_871);
or U911 (N_911,N_889,N_881);
nand U912 (N_912,N_875,N_899);
and U913 (N_913,N_872,N_864);
nand U914 (N_914,N_851,N_880);
nor U915 (N_915,N_877,N_860);
nand U916 (N_916,N_854,N_883);
nor U917 (N_917,N_873,N_868);
and U918 (N_918,N_886,N_885);
nor U919 (N_919,N_863,N_884);
nor U920 (N_920,N_896,N_878);
nor U921 (N_921,N_891,N_894);
and U922 (N_922,N_850,N_855);
nor U923 (N_923,N_879,N_867);
and U924 (N_924,N_856,N_852);
and U925 (N_925,N_854,N_851);
nor U926 (N_926,N_866,N_874);
or U927 (N_927,N_857,N_860);
or U928 (N_928,N_853,N_870);
and U929 (N_929,N_887,N_863);
xnor U930 (N_930,N_881,N_892);
or U931 (N_931,N_866,N_865);
and U932 (N_932,N_886,N_898);
and U933 (N_933,N_883,N_869);
or U934 (N_934,N_895,N_882);
or U935 (N_935,N_864,N_852);
or U936 (N_936,N_854,N_852);
and U937 (N_937,N_851,N_876);
and U938 (N_938,N_882,N_871);
xor U939 (N_939,N_864,N_890);
and U940 (N_940,N_851,N_896);
nand U941 (N_941,N_885,N_869);
and U942 (N_942,N_851,N_886);
nor U943 (N_943,N_866,N_891);
nor U944 (N_944,N_864,N_857);
nand U945 (N_945,N_885,N_884);
and U946 (N_946,N_887,N_853);
xnor U947 (N_947,N_874,N_856);
or U948 (N_948,N_856,N_897);
nand U949 (N_949,N_892,N_876);
nor U950 (N_950,N_913,N_911);
or U951 (N_951,N_915,N_917);
nor U952 (N_952,N_949,N_907);
and U953 (N_953,N_905,N_928);
or U954 (N_954,N_947,N_902);
nand U955 (N_955,N_936,N_943);
nor U956 (N_956,N_916,N_935);
xor U957 (N_957,N_904,N_909);
nand U958 (N_958,N_941,N_940);
and U959 (N_959,N_944,N_914);
nand U960 (N_960,N_920,N_929);
or U961 (N_961,N_925,N_906);
or U962 (N_962,N_927,N_918);
and U963 (N_963,N_939,N_930);
or U964 (N_964,N_923,N_933);
nor U965 (N_965,N_924,N_919);
nand U966 (N_966,N_945,N_903);
nor U967 (N_967,N_900,N_932);
and U968 (N_968,N_942,N_901);
nand U969 (N_969,N_948,N_912);
xor U970 (N_970,N_926,N_934);
xor U971 (N_971,N_910,N_921);
nand U972 (N_972,N_922,N_908);
nand U973 (N_973,N_946,N_937);
and U974 (N_974,N_938,N_931);
nor U975 (N_975,N_914,N_909);
xor U976 (N_976,N_949,N_933);
and U977 (N_977,N_918,N_945);
nor U978 (N_978,N_911,N_920);
nor U979 (N_979,N_915,N_918);
or U980 (N_980,N_904,N_912);
and U981 (N_981,N_914,N_919);
nand U982 (N_982,N_915,N_906);
and U983 (N_983,N_944,N_933);
or U984 (N_984,N_920,N_927);
nand U985 (N_985,N_903,N_915);
xnor U986 (N_986,N_917,N_900);
and U987 (N_987,N_913,N_909);
and U988 (N_988,N_913,N_928);
nand U989 (N_989,N_909,N_900);
nor U990 (N_990,N_917,N_902);
and U991 (N_991,N_903,N_947);
and U992 (N_992,N_913,N_907);
xnor U993 (N_993,N_933,N_914);
nand U994 (N_994,N_924,N_942);
and U995 (N_995,N_945,N_932);
or U996 (N_996,N_909,N_922);
xnor U997 (N_997,N_942,N_915);
and U998 (N_998,N_933,N_941);
nor U999 (N_999,N_914,N_949);
and U1000 (N_1000,N_959,N_977);
xnor U1001 (N_1001,N_962,N_955);
or U1002 (N_1002,N_963,N_991);
or U1003 (N_1003,N_999,N_972);
or U1004 (N_1004,N_951,N_979);
nor U1005 (N_1005,N_970,N_974);
nor U1006 (N_1006,N_950,N_984);
nand U1007 (N_1007,N_964,N_957);
or U1008 (N_1008,N_996,N_987);
or U1009 (N_1009,N_986,N_988);
nor U1010 (N_1010,N_966,N_980);
or U1011 (N_1011,N_995,N_975);
nor U1012 (N_1012,N_990,N_971);
or U1013 (N_1013,N_956,N_989);
nand U1014 (N_1014,N_973,N_983);
or U1015 (N_1015,N_961,N_981);
nor U1016 (N_1016,N_998,N_992);
nor U1017 (N_1017,N_954,N_969);
nand U1018 (N_1018,N_968,N_952);
and U1019 (N_1019,N_978,N_967);
nor U1020 (N_1020,N_993,N_960);
and U1021 (N_1021,N_976,N_997);
xor U1022 (N_1022,N_958,N_982);
nand U1023 (N_1023,N_994,N_965);
nor U1024 (N_1024,N_985,N_953);
nor U1025 (N_1025,N_995,N_986);
xnor U1026 (N_1026,N_966,N_985);
nor U1027 (N_1027,N_981,N_965);
and U1028 (N_1028,N_997,N_967);
nand U1029 (N_1029,N_983,N_959);
or U1030 (N_1030,N_972,N_981);
nand U1031 (N_1031,N_985,N_978);
and U1032 (N_1032,N_996,N_997);
xnor U1033 (N_1033,N_954,N_979);
nand U1034 (N_1034,N_982,N_991);
xnor U1035 (N_1035,N_978,N_962);
nor U1036 (N_1036,N_979,N_994);
and U1037 (N_1037,N_973,N_964);
nand U1038 (N_1038,N_956,N_978);
nand U1039 (N_1039,N_956,N_983);
or U1040 (N_1040,N_969,N_983);
nor U1041 (N_1041,N_962,N_966);
nor U1042 (N_1042,N_982,N_998);
and U1043 (N_1043,N_990,N_957);
nand U1044 (N_1044,N_965,N_989);
or U1045 (N_1045,N_959,N_957);
and U1046 (N_1046,N_982,N_965);
or U1047 (N_1047,N_995,N_991);
and U1048 (N_1048,N_967,N_984);
and U1049 (N_1049,N_993,N_974);
nand U1050 (N_1050,N_1049,N_1017);
and U1051 (N_1051,N_1047,N_1002);
nand U1052 (N_1052,N_1026,N_1037);
nand U1053 (N_1053,N_1030,N_1000);
xor U1054 (N_1054,N_1019,N_1048);
nor U1055 (N_1055,N_1009,N_1029);
or U1056 (N_1056,N_1040,N_1023);
and U1057 (N_1057,N_1007,N_1033);
nand U1058 (N_1058,N_1018,N_1043);
nand U1059 (N_1059,N_1012,N_1025);
nand U1060 (N_1060,N_1015,N_1013);
and U1061 (N_1061,N_1008,N_1011);
and U1062 (N_1062,N_1020,N_1045);
nor U1063 (N_1063,N_1016,N_1039);
and U1064 (N_1064,N_1010,N_1036);
nor U1065 (N_1065,N_1044,N_1014);
and U1066 (N_1066,N_1001,N_1032);
and U1067 (N_1067,N_1035,N_1028);
nand U1068 (N_1068,N_1004,N_1024);
xor U1069 (N_1069,N_1022,N_1005);
or U1070 (N_1070,N_1031,N_1034);
and U1071 (N_1071,N_1041,N_1046);
xnor U1072 (N_1072,N_1021,N_1038);
nand U1073 (N_1073,N_1006,N_1027);
nand U1074 (N_1074,N_1003,N_1042);
nand U1075 (N_1075,N_1045,N_1032);
or U1076 (N_1076,N_1046,N_1017);
and U1077 (N_1077,N_1008,N_1033);
and U1078 (N_1078,N_1031,N_1017);
nand U1079 (N_1079,N_1016,N_1030);
and U1080 (N_1080,N_1010,N_1014);
or U1081 (N_1081,N_1045,N_1029);
and U1082 (N_1082,N_1030,N_1034);
xor U1083 (N_1083,N_1040,N_1013);
nor U1084 (N_1084,N_1028,N_1005);
nor U1085 (N_1085,N_1010,N_1006);
or U1086 (N_1086,N_1027,N_1023);
or U1087 (N_1087,N_1003,N_1033);
nor U1088 (N_1088,N_1049,N_1001);
nor U1089 (N_1089,N_1018,N_1015);
nand U1090 (N_1090,N_1023,N_1021);
and U1091 (N_1091,N_1012,N_1032);
or U1092 (N_1092,N_1010,N_1023);
or U1093 (N_1093,N_1028,N_1010);
or U1094 (N_1094,N_1031,N_1026);
nand U1095 (N_1095,N_1016,N_1047);
xnor U1096 (N_1096,N_1010,N_1039);
nor U1097 (N_1097,N_1029,N_1039);
nor U1098 (N_1098,N_1002,N_1043);
or U1099 (N_1099,N_1041,N_1032);
and U1100 (N_1100,N_1057,N_1064);
or U1101 (N_1101,N_1070,N_1088);
xor U1102 (N_1102,N_1083,N_1071);
or U1103 (N_1103,N_1074,N_1072);
or U1104 (N_1104,N_1065,N_1096);
nand U1105 (N_1105,N_1087,N_1086);
or U1106 (N_1106,N_1077,N_1060);
xnor U1107 (N_1107,N_1051,N_1095);
or U1108 (N_1108,N_1056,N_1066);
xor U1109 (N_1109,N_1078,N_1058);
nor U1110 (N_1110,N_1093,N_1090);
xor U1111 (N_1111,N_1097,N_1053);
or U1112 (N_1112,N_1085,N_1063);
nor U1113 (N_1113,N_1059,N_1094);
and U1114 (N_1114,N_1080,N_1098);
nor U1115 (N_1115,N_1069,N_1075);
xor U1116 (N_1116,N_1067,N_1089);
or U1117 (N_1117,N_1054,N_1068);
nand U1118 (N_1118,N_1055,N_1081);
or U1119 (N_1119,N_1076,N_1099);
xnor U1120 (N_1120,N_1082,N_1091);
and U1121 (N_1121,N_1073,N_1084);
and U1122 (N_1122,N_1050,N_1092);
and U1123 (N_1123,N_1052,N_1061);
nor U1124 (N_1124,N_1079,N_1062);
or U1125 (N_1125,N_1054,N_1077);
nor U1126 (N_1126,N_1062,N_1082);
nand U1127 (N_1127,N_1095,N_1071);
nor U1128 (N_1128,N_1064,N_1098);
nor U1129 (N_1129,N_1078,N_1053);
and U1130 (N_1130,N_1056,N_1075);
or U1131 (N_1131,N_1077,N_1096);
nand U1132 (N_1132,N_1073,N_1074);
and U1133 (N_1133,N_1087,N_1090);
or U1134 (N_1134,N_1085,N_1058);
or U1135 (N_1135,N_1060,N_1061);
nor U1136 (N_1136,N_1064,N_1083);
nor U1137 (N_1137,N_1095,N_1093);
or U1138 (N_1138,N_1098,N_1095);
and U1139 (N_1139,N_1083,N_1053);
and U1140 (N_1140,N_1070,N_1062);
or U1141 (N_1141,N_1071,N_1081);
nor U1142 (N_1142,N_1088,N_1058);
or U1143 (N_1143,N_1063,N_1057);
or U1144 (N_1144,N_1068,N_1093);
xnor U1145 (N_1145,N_1078,N_1068);
and U1146 (N_1146,N_1057,N_1069);
nor U1147 (N_1147,N_1093,N_1096);
nand U1148 (N_1148,N_1084,N_1078);
or U1149 (N_1149,N_1081,N_1099);
nor U1150 (N_1150,N_1114,N_1138);
nor U1151 (N_1151,N_1103,N_1110);
nand U1152 (N_1152,N_1140,N_1111);
or U1153 (N_1153,N_1116,N_1130);
or U1154 (N_1154,N_1137,N_1134);
nor U1155 (N_1155,N_1104,N_1136);
or U1156 (N_1156,N_1117,N_1126);
and U1157 (N_1157,N_1112,N_1147);
xnor U1158 (N_1158,N_1143,N_1113);
nand U1159 (N_1159,N_1124,N_1142);
nand U1160 (N_1160,N_1135,N_1146);
nand U1161 (N_1161,N_1122,N_1123);
nand U1162 (N_1162,N_1101,N_1131);
nand U1163 (N_1163,N_1121,N_1139);
or U1164 (N_1164,N_1141,N_1127);
or U1165 (N_1165,N_1148,N_1125);
xnor U1166 (N_1166,N_1120,N_1144);
or U1167 (N_1167,N_1129,N_1105);
nand U1168 (N_1168,N_1132,N_1128);
nand U1169 (N_1169,N_1119,N_1118);
or U1170 (N_1170,N_1145,N_1149);
or U1171 (N_1171,N_1108,N_1109);
xor U1172 (N_1172,N_1107,N_1102);
nor U1173 (N_1173,N_1133,N_1106);
xor U1174 (N_1174,N_1115,N_1100);
nand U1175 (N_1175,N_1106,N_1107);
and U1176 (N_1176,N_1114,N_1140);
nand U1177 (N_1177,N_1134,N_1143);
nand U1178 (N_1178,N_1114,N_1133);
nand U1179 (N_1179,N_1104,N_1143);
or U1180 (N_1180,N_1136,N_1112);
nor U1181 (N_1181,N_1101,N_1132);
nand U1182 (N_1182,N_1122,N_1133);
nand U1183 (N_1183,N_1108,N_1127);
nand U1184 (N_1184,N_1122,N_1149);
nor U1185 (N_1185,N_1116,N_1138);
or U1186 (N_1186,N_1118,N_1103);
or U1187 (N_1187,N_1139,N_1108);
xor U1188 (N_1188,N_1143,N_1107);
xnor U1189 (N_1189,N_1134,N_1138);
or U1190 (N_1190,N_1137,N_1109);
or U1191 (N_1191,N_1146,N_1128);
nand U1192 (N_1192,N_1136,N_1111);
and U1193 (N_1193,N_1137,N_1111);
nand U1194 (N_1194,N_1137,N_1102);
xnor U1195 (N_1195,N_1146,N_1100);
or U1196 (N_1196,N_1129,N_1145);
nor U1197 (N_1197,N_1115,N_1106);
or U1198 (N_1198,N_1114,N_1141);
xnor U1199 (N_1199,N_1116,N_1145);
nand U1200 (N_1200,N_1172,N_1189);
nand U1201 (N_1201,N_1194,N_1185);
and U1202 (N_1202,N_1152,N_1174);
and U1203 (N_1203,N_1159,N_1171);
or U1204 (N_1204,N_1170,N_1175);
xor U1205 (N_1205,N_1162,N_1163);
and U1206 (N_1206,N_1184,N_1176);
or U1207 (N_1207,N_1173,N_1197);
or U1208 (N_1208,N_1180,N_1154);
and U1209 (N_1209,N_1198,N_1160);
nor U1210 (N_1210,N_1181,N_1192);
xor U1211 (N_1211,N_1179,N_1195);
and U1212 (N_1212,N_1183,N_1153);
nand U1213 (N_1213,N_1165,N_1168);
nor U1214 (N_1214,N_1188,N_1164);
and U1215 (N_1215,N_1186,N_1177);
nand U1216 (N_1216,N_1182,N_1190);
or U1217 (N_1217,N_1187,N_1196);
nor U1218 (N_1218,N_1161,N_1167);
nand U1219 (N_1219,N_1191,N_1166);
xor U1220 (N_1220,N_1178,N_1158);
or U1221 (N_1221,N_1199,N_1157);
nor U1222 (N_1222,N_1193,N_1156);
and U1223 (N_1223,N_1169,N_1150);
or U1224 (N_1224,N_1155,N_1151);
nor U1225 (N_1225,N_1181,N_1150);
or U1226 (N_1226,N_1183,N_1193);
xnor U1227 (N_1227,N_1166,N_1176);
and U1228 (N_1228,N_1187,N_1192);
and U1229 (N_1229,N_1190,N_1187);
and U1230 (N_1230,N_1155,N_1179);
or U1231 (N_1231,N_1192,N_1193);
nor U1232 (N_1232,N_1171,N_1182);
and U1233 (N_1233,N_1168,N_1172);
nor U1234 (N_1234,N_1172,N_1194);
and U1235 (N_1235,N_1153,N_1182);
nand U1236 (N_1236,N_1179,N_1164);
nand U1237 (N_1237,N_1191,N_1158);
nor U1238 (N_1238,N_1197,N_1157);
xnor U1239 (N_1239,N_1152,N_1183);
and U1240 (N_1240,N_1155,N_1165);
and U1241 (N_1241,N_1176,N_1199);
nand U1242 (N_1242,N_1166,N_1195);
nor U1243 (N_1243,N_1172,N_1154);
and U1244 (N_1244,N_1198,N_1197);
nor U1245 (N_1245,N_1169,N_1155);
nor U1246 (N_1246,N_1187,N_1156);
nand U1247 (N_1247,N_1157,N_1165);
or U1248 (N_1248,N_1189,N_1198);
nand U1249 (N_1249,N_1186,N_1152);
or U1250 (N_1250,N_1241,N_1244);
and U1251 (N_1251,N_1237,N_1212);
and U1252 (N_1252,N_1233,N_1203);
nand U1253 (N_1253,N_1248,N_1235);
nand U1254 (N_1254,N_1206,N_1204);
nor U1255 (N_1255,N_1238,N_1240);
nand U1256 (N_1256,N_1239,N_1207);
nand U1257 (N_1257,N_1224,N_1215);
and U1258 (N_1258,N_1220,N_1231);
and U1259 (N_1259,N_1201,N_1227);
xnor U1260 (N_1260,N_1242,N_1243);
or U1261 (N_1261,N_1223,N_1226);
xor U1262 (N_1262,N_1247,N_1229);
and U1263 (N_1263,N_1200,N_1225);
nand U1264 (N_1264,N_1214,N_1232);
xnor U1265 (N_1265,N_1245,N_1230);
nor U1266 (N_1266,N_1218,N_1249);
or U1267 (N_1267,N_1202,N_1216);
nor U1268 (N_1268,N_1236,N_1213);
and U1269 (N_1269,N_1210,N_1208);
or U1270 (N_1270,N_1228,N_1246);
nand U1271 (N_1271,N_1234,N_1221);
and U1272 (N_1272,N_1209,N_1205);
xor U1273 (N_1273,N_1211,N_1222);
xnor U1274 (N_1274,N_1219,N_1217);
or U1275 (N_1275,N_1240,N_1239);
and U1276 (N_1276,N_1233,N_1212);
nor U1277 (N_1277,N_1204,N_1245);
or U1278 (N_1278,N_1217,N_1232);
or U1279 (N_1279,N_1208,N_1232);
nand U1280 (N_1280,N_1228,N_1203);
and U1281 (N_1281,N_1202,N_1227);
nand U1282 (N_1282,N_1200,N_1234);
nor U1283 (N_1283,N_1214,N_1207);
and U1284 (N_1284,N_1212,N_1204);
nor U1285 (N_1285,N_1246,N_1244);
nor U1286 (N_1286,N_1219,N_1221);
nand U1287 (N_1287,N_1201,N_1218);
xnor U1288 (N_1288,N_1213,N_1246);
nor U1289 (N_1289,N_1214,N_1218);
nor U1290 (N_1290,N_1242,N_1224);
nand U1291 (N_1291,N_1234,N_1231);
and U1292 (N_1292,N_1241,N_1233);
nand U1293 (N_1293,N_1209,N_1222);
or U1294 (N_1294,N_1219,N_1228);
nor U1295 (N_1295,N_1248,N_1225);
nor U1296 (N_1296,N_1211,N_1228);
and U1297 (N_1297,N_1207,N_1242);
nand U1298 (N_1298,N_1226,N_1206);
and U1299 (N_1299,N_1206,N_1209);
or U1300 (N_1300,N_1283,N_1263);
nand U1301 (N_1301,N_1278,N_1276);
nand U1302 (N_1302,N_1280,N_1260);
or U1303 (N_1303,N_1250,N_1294);
nand U1304 (N_1304,N_1271,N_1266);
or U1305 (N_1305,N_1255,N_1256);
and U1306 (N_1306,N_1270,N_1274);
nor U1307 (N_1307,N_1269,N_1284);
nor U1308 (N_1308,N_1287,N_1275);
nand U1309 (N_1309,N_1279,N_1257);
nor U1310 (N_1310,N_1262,N_1251);
or U1311 (N_1311,N_1277,N_1286);
nand U1312 (N_1312,N_1288,N_1299);
nand U1313 (N_1313,N_1282,N_1297);
or U1314 (N_1314,N_1291,N_1268);
nor U1315 (N_1315,N_1261,N_1292);
nor U1316 (N_1316,N_1265,N_1273);
nand U1317 (N_1317,N_1289,N_1290);
nand U1318 (N_1318,N_1252,N_1267);
nand U1319 (N_1319,N_1258,N_1272);
and U1320 (N_1320,N_1295,N_1298);
xnor U1321 (N_1321,N_1293,N_1281);
and U1322 (N_1322,N_1285,N_1259);
nor U1323 (N_1323,N_1254,N_1264);
nor U1324 (N_1324,N_1296,N_1253);
and U1325 (N_1325,N_1273,N_1251);
nor U1326 (N_1326,N_1281,N_1251);
nand U1327 (N_1327,N_1280,N_1297);
and U1328 (N_1328,N_1292,N_1273);
or U1329 (N_1329,N_1267,N_1253);
or U1330 (N_1330,N_1279,N_1273);
nand U1331 (N_1331,N_1265,N_1287);
or U1332 (N_1332,N_1255,N_1266);
nor U1333 (N_1333,N_1262,N_1284);
nand U1334 (N_1334,N_1268,N_1278);
or U1335 (N_1335,N_1275,N_1274);
or U1336 (N_1336,N_1286,N_1253);
nor U1337 (N_1337,N_1250,N_1262);
or U1338 (N_1338,N_1284,N_1251);
nor U1339 (N_1339,N_1284,N_1273);
nor U1340 (N_1340,N_1285,N_1269);
nor U1341 (N_1341,N_1279,N_1296);
and U1342 (N_1342,N_1265,N_1292);
nand U1343 (N_1343,N_1294,N_1278);
nor U1344 (N_1344,N_1258,N_1268);
or U1345 (N_1345,N_1268,N_1276);
nand U1346 (N_1346,N_1289,N_1296);
nor U1347 (N_1347,N_1271,N_1288);
or U1348 (N_1348,N_1254,N_1258);
nor U1349 (N_1349,N_1295,N_1262);
and U1350 (N_1350,N_1330,N_1304);
nor U1351 (N_1351,N_1333,N_1316);
or U1352 (N_1352,N_1341,N_1342);
or U1353 (N_1353,N_1347,N_1339);
or U1354 (N_1354,N_1307,N_1300);
nand U1355 (N_1355,N_1315,N_1346);
nand U1356 (N_1356,N_1326,N_1349);
xor U1357 (N_1357,N_1317,N_1343);
nor U1358 (N_1358,N_1320,N_1336);
and U1359 (N_1359,N_1348,N_1345);
or U1360 (N_1360,N_1344,N_1302);
nand U1361 (N_1361,N_1335,N_1308);
nand U1362 (N_1362,N_1321,N_1306);
or U1363 (N_1363,N_1324,N_1332);
and U1364 (N_1364,N_1322,N_1331);
and U1365 (N_1365,N_1319,N_1303);
nor U1366 (N_1366,N_1314,N_1318);
nor U1367 (N_1367,N_1338,N_1305);
nor U1368 (N_1368,N_1310,N_1325);
nand U1369 (N_1369,N_1312,N_1313);
and U1370 (N_1370,N_1334,N_1340);
or U1371 (N_1371,N_1337,N_1329);
xor U1372 (N_1372,N_1328,N_1309);
nand U1373 (N_1373,N_1311,N_1327);
and U1374 (N_1374,N_1323,N_1301);
or U1375 (N_1375,N_1341,N_1308);
nand U1376 (N_1376,N_1316,N_1349);
nor U1377 (N_1377,N_1330,N_1318);
and U1378 (N_1378,N_1302,N_1313);
or U1379 (N_1379,N_1338,N_1301);
and U1380 (N_1380,N_1342,N_1321);
or U1381 (N_1381,N_1310,N_1302);
or U1382 (N_1382,N_1330,N_1335);
or U1383 (N_1383,N_1315,N_1316);
xor U1384 (N_1384,N_1318,N_1309);
nor U1385 (N_1385,N_1343,N_1348);
or U1386 (N_1386,N_1326,N_1347);
nor U1387 (N_1387,N_1342,N_1330);
nand U1388 (N_1388,N_1335,N_1341);
and U1389 (N_1389,N_1333,N_1320);
and U1390 (N_1390,N_1306,N_1315);
nand U1391 (N_1391,N_1338,N_1336);
xor U1392 (N_1392,N_1323,N_1313);
or U1393 (N_1393,N_1308,N_1302);
and U1394 (N_1394,N_1303,N_1318);
and U1395 (N_1395,N_1303,N_1317);
and U1396 (N_1396,N_1333,N_1310);
nor U1397 (N_1397,N_1349,N_1343);
nand U1398 (N_1398,N_1329,N_1338);
or U1399 (N_1399,N_1308,N_1349);
nand U1400 (N_1400,N_1396,N_1370);
nand U1401 (N_1401,N_1362,N_1391);
or U1402 (N_1402,N_1380,N_1395);
and U1403 (N_1403,N_1392,N_1363);
and U1404 (N_1404,N_1382,N_1367);
and U1405 (N_1405,N_1384,N_1372);
nor U1406 (N_1406,N_1365,N_1386);
nand U1407 (N_1407,N_1366,N_1399);
and U1408 (N_1408,N_1383,N_1393);
or U1409 (N_1409,N_1354,N_1378);
nor U1410 (N_1410,N_1360,N_1356);
xnor U1411 (N_1411,N_1353,N_1387);
xnor U1412 (N_1412,N_1358,N_1361);
nand U1413 (N_1413,N_1374,N_1388);
nor U1414 (N_1414,N_1377,N_1379);
nor U1415 (N_1415,N_1368,N_1375);
and U1416 (N_1416,N_1397,N_1369);
and U1417 (N_1417,N_1390,N_1385);
and U1418 (N_1418,N_1357,N_1350);
or U1419 (N_1419,N_1376,N_1364);
nor U1420 (N_1420,N_1371,N_1381);
or U1421 (N_1421,N_1355,N_1359);
nor U1422 (N_1422,N_1351,N_1389);
nor U1423 (N_1423,N_1398,N_1394);
and U1424 (N_1424,N_1373,N_1352);
nor U1425 (N_1425,N_1398,N_1362);
nor U1426 (N_1426,N_1372,N_1381);
or U1427 (N_1427,N_1388,N_1387);
nand U1428 (N_1428,N_1386,N_1395);
and U1429 (N_1429,N_1385,N_1395);
or U1430 (N_1430,N_1397,N_1365);
or U1431 (N_1431,N_1359,N_1366);
or U1432 (N_1432,N_1387,N_1372);
or U1433 (N_1433,N_1362,N_1376);
nand U1434 (N_1434,N_1352,N_1350);
and U1435 (N_1435,N_1389,N_1372);
or U1436 (N_1436,N_1364,N_1383);
nor U1437 (N_1437,N_1371,N_1394);
or U1438 (N_1438,N_1391,N_1387);
nor U1439 (N_1439,N_1398,N_1369);
xnor U1440 (N_1440,N_1381,N_1367);
nor U1441 (N_1441,N_1362,N_1364);
nand U1442 (N_1442,N_1390,N_1396);
or U1443 (N_1443,N_1388,N_1362);
or U1444 (N_1444,N_1385,N_1366);
and U1445 (N_1445,N_1351,N_1359);
nor U1446 (N_1446,N_1355,N_1354);
nor U1447 (N_1447,N_1361,N_1389);
nand U1448 (N_1448,N_1371,N_1388);
xnor U1449 (N_1449,N_1390,N_1367);
nor U1450 (N_1450,N_1409,N_1445);
nand U1451 (N_1451,N_1427,N_1424);
xnor U1452 (N_1452,N_1447,N_1400);
or U1453 (N_1453,N_1405,N_1432);
or U1454 (N_1454,N_1414,N_1429);
nand U1455 (N_1455,N_1428,N_1412);
nor U1456 (N_1456,N_1415,N_1446);
nand U1457 (N_1457,N_1416,N_1421);
and U1458 (N_1458,N_1449,N_1418);
or U1459 (N_1459,N_1442,N_1441);
nand U1460 (N_1460,N_1439,N_1433);
nand U1461 (N_1461,N_1420,N_1411);
and U1462 (N_1462,N_1408,N_1438);
nand U1463 (N_1463,N_1435,N_1413);
or U1464 (N_1464,N_1434,N_1430);
and U1465 (N_1465,N_1403,N_1417);
nand U1466 (N_1466,N_1404,N_1448);
nand U1467 (N_1467,N_1406,N_1431);
nor U1468 (N_1468,N_1419,N_1410);
and U1469 (N_1469,N_1436,N_1437);
or U1470 (N_1470,N_1402,N_1440);
or U1471 (N_1471,N_1407,N_1426);
nor U1472 (N_1472,N_1443,N_1444);
and U1473 (N_1473,N_1425,N_1423);
nor U1474 (N_1474,N_1422,N_1401);
and U1475 (N_1475,N_1446,N_1404);
nor U1476 (N_1476,N_1403,N_1413);
nand U1477 (N_1477,N_1445,N_1405);
and U1478 (N_1478,N_1413,N_1420);
nor U1479 (N_1479,N_1419,N_1428);
and U1480 (N_1480,N_1414,N_1423);
nand U1481 (N_1481,N_1400,N_1402);
nor U1482 (N_1482,N_1427,N_1426);
or U1483 (N_1483,N_1438,N_1423);
nor U1484 (N_1484,N_1415,N_1426);
and U1485 (N_1485,N_1421,N_1427);
xor U1486 (N_1486,N_1411,N_1428);
nor U1487 (N_1487,N_1444,N_1414);
and U1488 (N_1488,N_1416,N_1427);
and U1489 (N_1489,N_1448,N_1409);
and U1490 (N_1490,N_1406,N_1421);
and U1491 (N_1491,N_1402,N_1445);
nand U1492 (N_1492,N_1412,N_1444);
nor U1493 (N_1493,N_1407,N_1413);
or U1494 (N_1494,N_1426,N_1423);
nor U1495 (N_1495,N_1438,N_1407);
and U1496 (N_1496,N_1407,N_1412);
or U1497 (N_1497,N_1442,N_1408);
nand U1498 (N_1498,N_1401,N_1403);
nor U1499 (N_1499,N_1426,N_1419);
nand U1500 (N_1500,N_1489,N_1457);
nand U1501 (N_1501,N_1497,N_1473);
nor U1502 (N_1502,N_1494,N_1471);
or U1503 (N_1503,N_1490,N_1493);
nand U1504 (N_1504,N_1480,N_1452);
xor U1505 (N_1505,N_1492,N_1466);
nor U1506 (N_1506,N_1469,N_1479);
or U1507 (N_1507,N_1476,N_1450);
nor U1508 (N_1508,N_1472,N_1496);
and U1509 (N_1509,N_1456,N_1458);
and U1510 (N_1510,N_1463,N_1478);
nor U1511 (N_1511,N_1475,N_1470);
nor U1512 (N_1512,N_1488,N_1484);
and U1513 (N_1513,N_1468,N_1495);
xnor U1514 (N_1514,N_1499,N_1454);
and U1515 (N_1515,N_1487,N_1481);
nor U1516 (N_1516,N_1462,N_1451);
and U1517 (N_1517,N_1491,N_1483);
nand U1518 (N_1518,N_1485,N_1482);
and U1519 (N_1519,N_1498,N_1465);
nand U1520 (N_1520,N_1455,N_1459);
xor U1521 (N_1521,N_1464,N_1453);
xor U1522 (N_1522,N_1460,N_1461);
nor U1523 (N_1523,N_1477,N_1467);
and U1524 (N_1524,N_1486,N_1474);
or U1525 (N_1525,N_1491,N_1498);
nand U1526 (N_1526,N_1481,N_1484);
nand U1527 (N_1527,N_1485,N_1478);
and U1528 (N_1528,N_1470,N_1473);
and U1529 (N_1529,N_1461,N_1489);
and U1530 (N_1530,N_1460,N_1451);
xor U1531 (N_1531,N_1462,N_1483);
or U1532 (N_1532,N_1472,N_1481);
nor U1533 (N_1533,N_1450,N_1451);
and U1534 (N_1534,N_1481,N_1485);
nor U1535 (N_1535,N_1472,N_1458);
or U1536 (N_1536,N_1495,N_1452);
nor U1537 (N_1537,N_1481,N_1497);
and U1538 (N_1538,N_1496,N_1480);
nor U1539 (N_1539,N_1463,N_1484);
or U1540 (N_1540,N_1467,N_1469);
nand U1541 (N_1541,N_1461,N_1452);
nor U1542 (N_1542,N_1480,N_1499);
and U1543 (N_1543,N_1491,N_1450);
nand U1544 (N_1544,N_1456,N_1454);
nor U1545 (N_1545,N_1479,N_1497);
xor U1546 (N_1546,N_1462,N_1477);
or U1547 (N_1547,N_1469,N_1466);
nor U1548 (N_1548,N_1464,N_1481);
nor U1549 (N_1549,N_1497,N_1477);
nor U1550 (N_1550,N_1548,N_1519);
or U1551 (N_1551,N_1534,N_1504);
or U1552 (N_1552,N_1516,N_1531);
nor U1553 (N_1553,N_1512,N_1541);
nor U1554 (N_1554,N_1542,N_1540);
nand U1555 (N_1555,N_1536,N_1509);
xor U1556 (N_1556,N_1535,N_1505);
nor U1557 (N_1557,N_1507,N_1511);
nor U1558 (N_1558,N_1502,N_1526);
nor U1559 (N_1559,N_1518,N_1501);
nor U1560 (N_1560,N_1515,N_1522);
or U1561 (N_1561,N_1545,N_1527);
nor U1562 (N_1562,N_1529,N_1547);
and U1563 (N_1563,N_1544,N_1539);
or U1564 (N_1564,N_1537,N_1524);
and U1565 (N_1565,N_1546,N_1508);
or U1566 (N_1566,N_1530,N_1520);
and U1567 (N_1567,N_1543,N_1503);
nor U1568 (N_1568,N_1514,N_1500);
and U1569 (N_1569,N_1538,N_1523);
or U1570 (N_1570,N_1525,N_1513);
nand U1571 (N_1571,N_1517,N_1549);
or U1572 (N_1572,N_1528,N_1510);
nor U1573 (N_1573,N_1532,N_1521);
or U1574 (N_1574,N_1506,N_1533);
xor U1575 (N_1575,N_1547,N_1527);
xor U1576 (N_1576,N_1507,N_1500);
nor U1577 (N_1577,N_1546,N_1513);
xnor U1578 (N_1578,N_1502,N_1529);
or U1579 (N_1579,N_1514,N_1520);
nand U1580 (N_1580,N_1517,N_1510);
xnor U1581 (N_1581,N_1521,N_1542);
nand U1582 (N_1582,N_1505,N_1549);
nand U1583 (N_1583,N_1523,N_1508);
xnor U1584 (N_1584,N_1517,N_1526);
xnor U1585 (N_1585,N_1535,N_1526);
nor U1586 (N_1586,N_1549,N_1545);
and U1587 (N_1587,N_1534,N_1531);
and U1588 (N_1588,N_1504,N_1508);
or U1589 (N_1589,N_1500,N_1511);
and U1590 (N_1590,N_1531,N_1524);
nor U1591 (N_1591,N_1521,N_1540);
and U1592 (N_1592,N_1503,N_1502);
or U1593 (N_1593,N_1516,N_1530);
nor U1594 (N_1594,N_1506,N_1527);
and U1595 (N_1595,N_1532,N_1511);
or U1596 (N_1596,N_1519,N_1535);
nand U1597 (N_1597,N_1529,N_1540);
or U1598 (N_1598,N_1523,N_1535);
or U1599 (N_1599,N_1509,N_1529);
nor U1600 (N_1600,N_1553,N_1566);
nand U1601 (N_1601,N_1593,N_1595);
nor U1602 (N_1602,N_1584,N_1552);
and U1603 (N_1603,N_1570,N_1581);
and U1604 (N_1604,N_1563,N_1554);
nor U1605 (N_1605,N_1556,N_1560);
nor U1606 (N_1606,N_1589,N_1591);
and U1607 (N_1607,N_1550,N_1557);
xor U1608 (N_1608,N_1599,N_1592);
nand U1609 (N_1609,N_1558,N_1583);
nor U1610 (N_1610,N_1567,N_1565);
xnor U1611 (N_1611,N_1576,N_1578);
or U1612 (N_1612,N_1568,N_1577);
or U1613 (N_1613,N_1572,N_1594);
and U1614 (N_1614,N_1596,N_1590);
nand U1615 (N_1615,N_1571,N_1573);
xor U1616 (N_1616,N_1555,N_1551);
nand U1617 (N_1617,N_1559,N_1562);
nand U1618 (N_1618,N_1569,N_1564);
nand U1619 (N_1619,N_1585,N_1580);
nor U1620 (N_1620,N_1561,N_1598);
nand U1621 (N_1621,N_1587,N_1579);
nand U1622 (N_1622,N_1597,N_1575);
or U1623 (N_1623,N_1574,N_1582);
xor U1624 (N_1624,N_1588,N_1586);
xnor U1625 (N_1625,N_1554,N_1588);
nand U1626 (N_1626,N_1555,N_1562);
or U1627 (N_1627,N_1578,N_1553);
or U1628 (N_1628,N_1578,N_1593);
xor U1629 (N_1629,N_1586,N_1558);
or U1630 (N_1630,N_1581,N_1594);
nand U1631 (N_1631,N_1560,N_1563);
nand U1632 (N_1632,N_1573,N_1576);
nand U1633 (N_1633,N_1576,N_1561);
and U1634 (N_1634,N_1591,N_1572);
or U1635 (N_1635,N_1596,N_1560);
or U1636 (N_1636,N_1578,N_1566);
and U1637 (N_1637,N_1553,N_1558);
nand U1638 (N_1638,N_1580,N_1554);
nand U1639 (N_1639,N_1596,N_1561);
nor U1640 (N_1640,N_1596,N_1550);
or U1641 (N_1641,N_1566,N_1587);
or U1642 (N_1642,N_1591,N_1599);
and U1643 (N_1643,N_1595,N_1570);
nand U1644 (N_1644,N_1592,N_1582);
xor U1645 (N_1645,N_1561,N_1582);
or U1646 (N_1646,N_1553,N_1573);
nand U1647 (N_1647,N_1550,N_1595);
or U1648 (N_1648,N_1593,N_1564);
and U1649 (N_1649,N_1553,N_1561);
and U1650 (N_1650,N_1606,N_1640);
and U1651 (N_1651,N_1627,N_1601);
nand U1652 (N_1652,N_1629,N_1602);
nand U1653 (N_1653,N_1644,N_1643);
nor U1654 (N_1654,N_1634,N_1648);
and U1655 (N_1655,N_1633,N_1647);
nand U1656 (N_1656,N_1624,N_1631);
nand U1657 (N_1657,N_1637,N_1609);
and U1658 (N_1658,N_1613,N_1617);
xor U1659 (N_1659,N_1618,N_1628);
xor U1660 (N_1660,N_1636,N_1616);
and U1661 (N_1661,N_1612,N_1623);
nor U1662 (N_1662,N_1619,N_1610);
or U1663 (N_1663,N_1611,N_1605);
or U1664 (N_1664,N_1638,N_1649);
or U1665 (N_1665,N_1646,N_1632);
nand U1666 (N_1666,N_1641,N_1608);
nand U1667 (N_1667,N_1630,N_1639);
or U1668 (N_1668,N_1642,N_1603);
xnor U1669 (N_1669,N_1622,N_1604);
nor U1670 (N_1670,N_1635,N_1645);
xnor U1671 (N_1671,N_1620,N_1600);
or U1672 (N_1672,N_1607,N_1614);
xor U1673 (N_1673,N_1626,N_1621);
nor U1674 (N_1674,N_1625,N_1615);
nor U1675 (N_1675,N_1623,N_1609);
xnor U1676 (N_1676,N_1638,N_1646);
nand U1677 (N_1677,N_1605,N_1620);
nor U1678 (N_1678,N_1635,N_1618);
and U1679 (N_1679,N_1643,N_1645);
or U1680 (N_1680,N_1621,N_1614);
or U1681 (N_1681,N_1614,N_1629);
nor U1682 (N_1682,N_1612,N_1644);
nand U1683 (N_1683,N_1628,N_1616);
nand U1684 (N_1684,N_1636,N_1603);
or U1685 (N_1685,N_1603,N_1615);
or U1686 (N_1686,N_1644,N_1641);
or U1687 (N_1687,N_1613,N_1608);
xor U1688 (N_1688,N_1635,N_1627);
and U1689 (N_1689,N_1609,N_1608);
nor U1690 (N_1690,N_1607,N_1605);
nor U1691 (N_1691,N_1600,N_1625);
and U1692 (N_1692,N_1621,N_1638);
and U1693 (N_1693,N_1642,N_1602);
nor U1694 (N_1694,N_1622,N_1632);
xnor U1695 (N_1695,N_1644,N_1613);
or U1696 (N_1696,N_1602,N_1605);
nand U1697 (N_1697,N_1616,N_1649);
nor U1698 (N_1698,N_1621,N_1630);
nand U1699 (N_1699,N_1636,N_1628);
nor U1700 (N_1700,N_1683,N_1668);
or U1701 (N_1701,N_1690,N_1678);
nand U1702 (N_1702,N_1667,N_1694);
and U1703 (N_1703,N_1681,N_1687);
nor U1704 (N_1704,N_1696,N_1672);
and U1705 (N_1705,N_1691,N_1666);
and U1706 (N_1706,N_1671,N_1673);
nor U1707 (N_1707,N_1662,N_1660);
nor U1708 (N_1708,N_1664,N_1677);
or U1709 (N_1709,N_1684,N_1679);
and U1710 (N_1710,N_1656,N_1657);
nand U1711 (N_1711,N_1692,N_1685);
nor U1712 (N_1712,N_1676,N_1686);
xor U1713 (N_1713,N_1654,N_1670);
nor U1714 (N_1714,N_1675,N_1655);
nand U1715 (N_1715,N_1697,N_1650);
xnor U1716 (N_1716,N_1665,N_1693);
and U1717 (N_1717,N_1695,N_1698);
nand U1718 (N_1718,N_1661,N_1652);
nand U1719 (N_1719,N_1699,N_1689);
nand U1720 (N_1720,N_1663,N_1669);
or U1721 (N_1721,N_1682,N_1651);
or U1722 (N_1722,N_1659,N_1653);
nand U1723 (N_1723,N_1680,N_1674);
nand U1724 (N_1724,N_1658,N_1688);
nand U1725 (N_1725,N_1681,N_1653);
or U1726 (N_1726,N_1675,N_1666);
nor U1727 (N_1727,N_1696,N_1684);
xnor U1728 (N_1728,N_1654,N_1651);
nor U1729 (N_1729,N_1667,N_1657);
or U1730 (N_1730,N_1688,N_1673);
or U1731 (N_1731,N_1676,N_1684);
xnor U1732 (N_1732,N_1675,N_1693);
nor U1733 (N_1733,N_1669,N_1659);
nand U1734 (N_1734,N_1675,N_1652);
xnor U1735 (N_1735,N_1689,N_1667);
or U1736 (N_1736,N_1696,N_1662);
and U1737 (N_1737,N_1658,N_1695);
nor U1738 (N_1738,N_1682,N_1663);
nand U1739 (N_1739,N_1678,N_1671);
and U1740 (N_1740,N_1678,N_1665);
xnor U1741 (N_1741,N_1673,N_1653);
or U1742 (N_1742,N_1676,N_1679);
nor U1743 (N_1743,N_1695,N_1678);
and U1744 (N_1744,N_1691,N_1671);
and U1745 (N_1745,N_1661,N_1688);
nor U1746 (N_1746,N_1658,N_1666);
nor U1747 (N_1747,N_1696,N_1653);
nand U1748 (N_1748,N_1670,N_1669);
and U1749 (N_1749,N_1665,N_1659);
nand U1750 (N_1750,N_1738,N_1735);
xor U1751 (N_1751,N_1722,N_1702);
nand U1752 (N_1752,N_1724,N_1726);
nand U1753 (N_1753,N_1746,N_1716);
xor U1754 (N_1754,N_1705,N_1736);
xor U1755 (N_1755,N_1741,N_1719);
and U1756 (N_1756,N_1749,N_1717);
nor U1757 (N_1757,N_1729,N_1710);
nand U1758 (N_1758,N_1707,N_1727);
nand U1759 (N_1759,N_1732,N_1714);
or U1760 (N_1760,N_1706,N_1720);
nand U1761 (N_1761,N_1737,N_1718);
nor U1762 (N_1762,N_1725,N_1740);
or U1763 (N_1763,N_1723,N_1715);
and U1764 (N_1764,N_1708,N_1742);
and U1765 (N_1765,N_1704,N_1701);
nand U1766 (N_1766,N_1709,N_1745);
and U1767 (N_1767,N_1713,N_1712);
nand U1768 (N_1768,N_1739,N_1743);
nor U1769 (N_1769,N_1747,N_1730);
nand U1770 (N_1770,N_1711,N_1733);
and U1771 (N_1771,N_1748,N_1728);
nand U1772 (N_1772,N_1700,N_1721);
nand U1773 (N_1773,N_1731,N_1734);
and U1774 (N_1774,N_1703,N_1744);
xor U1775 (N_1775,N_1742,N_1732);
and U1776 (N_1776,N_1701,N_1749);
nand U1777 (N_1777,N_1721,N_1712);
and U1778 (N_1778,N_1731,N_1724);
nand U1779 (N_1779,N_1739,N_1726);
and U1780 (N_1780,N_1737,N_1734);
nor U1781 (N_1781,N_1741,N_1700);
or U1782 (N_1782,N_1747,N_1748);
nor U1783 (N_1783,N_1726,N_1747);
nand U1784 (N_1784,N_1734,N_1711);
or U1785 (N_1785,N_1739,N_1730);
and U1786 (N_1786,N_1719,N_1733);
nand U1787 (N_1787,N_1712,N_1720);
nand U1788 (N_1788,N_1722,N_1730);
nor U1789 (N_1789,N_1720,N_1738);
and U1790 (N_1790,N_1700,N_1738);
nand U1791 (N_1791,N_1717,N_1706);
xnor U1792 (N_1792,N_1734,N_1742);
and U1793 (N_1793,N_1744,N_1731);
xor U1794 (N_1794,N_1707,N_1737);
and U1795 (N_1795,N_1704,N_1723);
nor U1796 (N_1796,N_1742,N_1701);
nand U1797 (N_1797,N_1746,N_1715);
or U1798 (N_1798,N_1700,N_1731);
and U1799 (N_1799,N_1749,N_1704);
or U1800 (N_1800,N_1793,N_1791);
nand U1801 (N_1801,N_1760,N_1770);
nand U1802 (N_1802,N_1796,N_1774);
nand U1803 (N_1803,N_1783,N_1799);
and U1804 (N_1804,N_1768,N_1781);
nand U1805 (N_1805,N_1780,N_1790);
xor U1806 (N_1806,N_1753,N_1752);
nand U1807 (N_1807,N_1764,N_1789);
and U1808 (N_1808,N_1775,N_1792);
nor U1809 (N_1809,N_1761,N_1765);
and U1810 (N_1810,N_1759,N_1762);
nor U1811 (N_1811,N_1772,N_1773);
nand U1812 (N_1812,N_1778,N_1751);
nand U1813 (N_1813,N_1757,N_1787);
nor U1814 (N_1814,N_1782,N_1766);
nor U1815 (N_1815,N_1754,N_1756);
nand U1816 (N_1816,N_1785,N_1755);
nor U1817 (N_1817,N_1779,N_1798);
or U1818 (N_1818,N_1777,N_1769);
nor U1819 (N_1819,N_1776,N_1758);
and U1820 (N_1820,N_1795,N_1750);
and U1821 (N_1821,N_1786,N_1767);
nand U1822 (N_1822,N_1794,N_1788);
nand U1823 (N_1823,N_1763,N_1771);
nor U1824 (N_1824,N_1784,N_1797);
or U1825 (N_1825,N_1755,N_1791);
and U1826 (N_1826,N_1778,N_1761);
nand U1827 (N_1827,N_1783,N_1781);
nand U1828 (N_1828,N_1775,N_1786);
nor U1829 (N_1829,N_1778,N_1756);
nor U1830 (N_1830,N_1770,N_1771);
or U1831 (N_1831,N_1775,N_1794);
or U1832 (N_1832,N_1799,N_1752);
nor U1833 (N_1833,N_1772,N_1766);
or U1834 (N_1834,N_1755,N_1756);
and U1835 (N_1835,N_1787,N_1768);
and U1836 (N_1836,N_1772,N_1797);
nand U1837 (N_1837,N_1758,N_1794);
and U1838 (N_1838,N_1772,N_1750);
nor U1839 (N_1839,N_1786,N_1764);
nand U1840 (N_1840,N_1762,N_1789);
nand U1841 (N_1841,N_1760,N_1773);
xor U1842 (N_1842,N_1783,N_1777);
and U1843 (N_1843,N_1781,N_1753);
nor U1844 (N_1844,N_1755,N_1790);
and U1845 (N_1845,N_1763,N_1775);
and U1846 (N_1846,N_1765,N_1755);
nand U1847 (N_1847,N_1754,N_1795);
nor U1848 (N_1848,N_1779,N_1752);
nor U1849 (N_1849,N_1761,N_1757);
xnor U1850 (N_1850,N_1822,N_1849);
nor U1851 (N_1851,N_1848,N_1837);
nor U1852 (N_1852,N_1832,N_1802);
nand U1853 (N_1853,N_1824,N_1814);
nand U1854 (N_1854,N_1811,N_1842);
and U1855 (N_1855,N_1805,N_1841);
nand U1856 (N_1856,N_1839,N_1846);
nand U1857 (N_1857,N_1819,N_1847);
nand U1858 (N_1858,N_1816,N_1834);
or U1859 (N_1859,N_1813,N_1817);
nor U1860 (N_1860,N_1818,N_1831);
or U1861 (N_1861,N_1815,N_1833);
or U1862 (N_1862,N_1806,N_1826);
nor U1863 (N_1863,N_1809,N_1845);
xor U1864 (N_1864,N_1830,N_1844);
or U1865 (N_1865,N_1825,N_1836);
nand U1866 (N_1866,N_1807,N_1803);
nand U1867 (N_1867,N_1829,N_1820);
nor U1868 (N_1868,N_1843,N_1835);
or U1869 (N_1869,N_1810,N_1812);
or U1870 (N_1870,N_1838,N_1808);
xor U1871 (N_1871,N_1827,N_1828);
or U1872 (N_1872,N_1804,N_1801);
nand U1873 (N_1873,N_1821,N_1840);
or U1874 (N_1874,N_1800,N_1823);
or U1875 (N_1875,N_1803,N_1843);
nor U1876 (N_1876,N_1840,N_1814);
nor U1877 (N_1877,N_1836,N_1833);
or U1878 (N_1878,N_1834,N_1818);
or U1879 (N_1879,N_1841,N_1836);
and U1880 (N_1880,N_1839,N_1818);
or U1881 (N_1881,N_1824,N_1817);
nor U1882 (N_1882,N_1828,N_1810);
nand U1883 (N_1883,N_1848,N_1800);
xor U1884 (N_1884,N_1814,N_1845);
nand U1885 (N_1885,N_1815,N_1847);
nand U1886 (N_1886,N_1832,N_1806);
nor U1887 (N_1887,N_1839,N_1826);
nand U1888 (N_1888,N_1835,N_1836);
or U1889 (N_1889,N_1845,N_1843);
or U1890 (N_1890,N_1809,N_1846);
nand U1891 (N_1891,N_1801,N_1848);
nand U1892 (N_1892,N_1838,N_1840);
nand U1893 (N_1893,N_1831,N_1802);
xor U1894 (N_1894,N_1817,N_1830);
nor U1895 (N_1895,N_1819,N_1830);
or U1896 (N_1896,N_1841,N_1815);
xor U1897 (N_1897,N_1825,N_1829);
xor U1898 (N_1898,N_1804,N_1837);
nand U1899 (N_1899,N_1822,N_1848);
and U1900 (N_1900,N_1890,N_1897);
nor U1901 (N_1901,N_1872,N_1887);
or U1902 (N_1902,N_1893,N_1861);
or U1903 (N_1903,N_1855,N_1894);
xnor U1904 (N_1904,N_1896,N_1867);
nor U1905 (N_1905,N_1865,N_1866);
and U1906 (N_1906,N_1868,N_1885);
nor U1907 (N_1907,N_1882,N_1862);
and U1908 (N_1908,N_1886,N_1891);
nor U1909 (N_1909,N_1856,N_1870);
nand U1910 (N_1910,N_1875,N_1858);
or U1911 (N_1911,N_1873,N_1878);
nor U1912 (N_1912,N_1857,N_1877);
or U1913 (N_1913,N_1853,N_1860);
nand U1914 (N_1914,N_1863,N_1898);
nand U1915 (N_1915,N_1899,N_1854);
and U1916 (N_1916,N_1888,N_1852);
xnor U1917 (N_1917,N_1869,N_1864);
or U1918 (N_1918,N_1851,N_1876);
and U1919 (N_1919,N_1895,N_1880);
or U1920 (N_1920,N_1879,N_1850);
xor U1921 (N_1921,N_1883,N_1884);
or U1922 (N_1922,N_1859,N_1881);
nor U1923 (N_1923,N_1892,N_1889);
or U1924 (N_1924,N_1871,N_1874);
nand U1925 (N_1925,N_1877,N_1860);
nor U1926 (N_1926,N_1854,N_1882);
and U1927 (N_1927,N_1871,N_1898);
nand U1928 (N_1928,N_1850,N_1889);
and U1929 (N_1929,N_1899,N_1877);
nand U1930 (N_1930,N_1876,N_1896);
and U1931 (N_1931,N_1863,N_1897);
and U1932 (N_1932,N_1890,N_1862);
and U1933 (N_1933,N_1860,N_1889);
or U1934 (N_1934,N_1883,N_1880);
nand U1935 (N_1935,N_1880,N_1859);
nand U1936 (N_1936,N_1872,N_1866);
and U1937 (N_1937,N_1861,N_1873);
nor U1938 (N_1938,N_1874,N_1853);
nor U1939 (N_1939,N_1888,N_1880);
and U1940 (N_1940,N_1853,N_1882);
xor U1941 (N_1941,N_1887,N_1877);
and U1942 (N_1942,N_1877,N_1861);
nor U1943 (N_1943,N_1866,N_1895);
nand U1944 (N_1944,N_1853,N_1850);
or U1945 (N_1945,N_1879,N_1890);
nor U1946 (N_1946,N_1864,N_1851);
or U1947 (N_1947,N_1871,N_1867);
and U1948 (N_1948,N_1863,N_1874);
and U1949 (N_1949,N_1851,N_1880);
or U1950 (N_1950,N_1909,N_1932);
and U1951 (N_1951,N_1912,N_1907);
or U1952 (N_1952,N_1929,N_1947);
and U1953 (N_1953,N_1944,N_1906);
or U1954 (N_1954,N_1915,N_1939);
nor U1955 (N_1955,N_1900,N_1946);
xor U1956 (N_1956,N_1924,N_1922);
nand U1957 (N_1957,N_1945,N_1903);
nand U1958 (N_1958,N_1926,N_1928);
or U1959 (N_1959,N_1923,N_1933);
and U1960 (N_1960,N_1943,N_1940);
nor U1961 (N_1961,N_1941,N_1921);
and U1962 (N_1962,N_1948,N_1905);
and U1963 (N_1963,N_1937,N_1925);
and U1964 (N_1964,N_1930,N_1914);
or U1965 (N_1965,N_1949,N_1942);
xnor U1966 (N_1966,N_1938,N_1911);
nor U1967 (N_1967,N_1936,N_1913);
or U1968 (N_1968,N_1931,N_1901);
or U1969 (N_1969,N_1904,N_1910);
and U1970 (N_1970,N_1916,N_1918);
and U1971 (N_1971,N_1935,N_1934);
nand U1972 (N_1972,N_1927,N_1908);
or U1973 (N_1973,N_1902,N_1920);
xnor U1974 (N_1974,N_1919,N_1917);
or U1975 (N_1975,N_1916,N_1926);
nand U1976 (N_1976,N_1949,N_1925);
nand U1977 (N_1977,N_1927,N_1935);
nor U1978 (N_1978,N_1903,N_1926);
xnor U1979 (N_1979,N_1930,N_1917);
nand U1980 (N_1980,N_1941,N_1906);
or U1981 (N_1981,N_1943,N_1922);
nor U1982 (N_1982,N_1911,N_1924);
xor U1983 (N_1983,N_1920,N_1924);
nand U1984 (N_1984,N_1902,N_1916);
or U1985 (N_1985,N_1944,N_1904);
or U1986 (N_1986,N_1949,N_1941);
and U1987 (N_1987,N_1908,N_1906);
nand U1988 (N_1988,N_1911,N_1919);
nor U1989 (N_1989,N_1912,N_1914);
and U1990 (N_1990,N_1928,N_1932);
or U1991 (N_1991,N_1903,N_1929);
nor U1992 (N_1992,N_1908,N_1936);
and U1993 (N_1993,N_1913,N_1911);
nor U1994 (N_1994,N_1928,N_1930);
nor U1995 (N_1995,N_1905,N_1909);
nor U1996 (N_1996,N_1940,N_1928);
and U1997 (N_1997,N_1903,N_1932);
nand U1998 (N_1998,N_1905,N_1919);
xor U1999 (N_1999,N_1910,N_1948);
nand U2000 (N_2000,N_1962,N_1986);
or U2001 (N_2001,N_1971,N_1998);
nor U2002 (N_2002,N_1969,N_1982);
nand U2003 (N_2003,N_1959,N_1993);
nor U2004 (N_2004,N_1960,N_1951);
and U2005 (N_2005,N_1968,N_1983);
nor U2006 (N_2006,N_1957,N_1992);
nand U2007 (N_2007,N_1994,N_1961);
nand U2008 (N_2008,N_1978,N_1975);
nor U2009 (N_2009,N_1953,N_1979);
nand U2010 (N_2010,N_1963,N_1999);
or U2011 (N_2011,N_1995,N_1952);
nor U2012 (N_2012,N_1997,N_1956);
and U2013 (N_2013,N_1950,N_1988);
nand U2014 (N_2014,N_1973,N_1974);
nand U2015 (N_2015,N_1958,N_1970);
nor U2016 (N_2016,N_1966,N_1996);
or U2017 (N_2017,N_1954,N_1972);
xor U2018 (N_2018,N_1955,N_1967);
or U2019 (N_2019,N_1984,N_1989);
nor U2020 (N_2020,N_1977,N_1981);
and U2021 (N_2021,N_1964,N_1965);
xor U2022 (N_2022,N_1985,N_1987);
or U2023 (N_2023,N_1976,N_1980);
or U2024 (N_2024,N_1990,N_1991);
nand U2025 (N_2025,N_1979,N_1973);
or U2026 (N_2026,N_1993,N_1998);
or U2027 (N_2027,N_1961,N_1962);
and U2028 (N_2028,N_1963,N_1982);
nor U2029 (N_2029,N_1966,N_1970);
nand U2030 (N_2030,N_1991,N_1973);
and U2031 (N_2031,N_1956,N_1972);
and U2032 (N_2032,N_1979,N_1958);
nand U2033 (N_2033,N_1960,N_1962);
or U2034 (N_2034,N_1969,N_1995);
and U2035 (N_2035,N_1950,N_1970);
nand U2036 (N_2036,N_1996,N_1961);
nor U2037 (N_2037,N_1975,N_1959);
nor U2038 (N_2038,N_1962,N_1965);
and U2039 (N_2039,N_1978,N_1998);
and U2040 (N_2040,N_1973,N_1963);
or U2041 (N_2041,N_1954,N_1971);
and U2042 (N_2042,N_1970,N_1969);
xnor U2043 (N_2043,N_1980,N_1991);
and U2044 (N_2044,N_1980,N_1972);
or U2045 (N_2045,N_1958,N_1959);
nand U2046 (N_2046,N_1965,N_1969);
nand U2047 (N_2047,N_1957,N_1954);
nand U2048 (N_2048,N_1962,N_1980);
nor U2049 (N_2049,N_1976,N_1972);
nand U2050 (N_2050,N_2034,N_2016);
nor U2051 (N_2051,N_2003,N_2032);
or U2052 (N_2052,N_2000,N_2004);
nand U2053 (N_2053,N_2002,N_2024);
xnor U2054 (N_2054,N_2007,N_2029);
and U2055 (N_2055,N_2036,N_2039);
nand U2056 (N_2056,N_2037,N_2045);
or U2057 (N_2057,N_2043,N_2030);
and U2058 (N_2058,N_2035,N_2010);
nand U2059 (N_2059,N_2049,N_2046);
and U2060 (N_2060,N_2013,N_2026);
nor U2061 (N_2061,N_2015,N_2025);
and U2062 (N_2062,N_2031,N_2042);
or U2063 (N_2063,N_2018,N_2008);
or U2064 (N_2064,N_2012,N_2014);
nand U2065 (N_2065,N_2009,N_2028);
nand U2066 (N_2066,N_2040,N_2021);
and U2067 (N_2067,N_2006,N_2001);
nor U2068 (N_2068,N_2041,N_2027);
or U2069 (N_2069,N_2047,N_2005);
xor U2070 (N_2070,N_2038,N_2017);
nand U2071 (N_2071,N_2020,N_2048);
nor U2072 (N_2072,N_2023,N_2022);
nor U2073 (N_2073,N_2044,N_2033);
and U2074 (N_2074,N_2011,N_2019);
nand U2075 (N_2075,N_2008,N_2036);
xor U2076 (N_2076,N_2046,N_2045);
nand U2077 (N_2077,N_2043,N_2032);
nor U2078 (N_2078,N_2014,N_2024);
xnor U2079 (N_2079,N_2001,N_2044);
and U2080 (N_2080,N_2049,N_2041);
nand U2081 (N_2081,N_2022,N_2025);
nor U2082 (N_2082,N_2013,N_2028);
and U2083 (N_2083,N_2008,N_2000);
xor U2084 (N_2084,N_2021,N_2025);
nor U2085 (N_2085,N_2021,N_2039);
or U2086 (N_2086,N_2039,N_2010);
or U2087 (N_2087,N_2034,N_2029);
and U2088 (N_2088,N_2003,N_2020);
and U2089 (N_2089,N_2044,N_2039);
xnor U2090 (N_2090,N_2035,N_2039);
or U2091 (N_2091,N_2022,N_2037);
nor U2092 (N_2092,N_2040,N_2048);
nor U2093 (N_2093,N_2038,N_2021);
nand U2094 (N_2094,N_2011,N_2002);
or U2095 (N_2095,N_2031,N_2020);
and U2096 (N_2096,N_2034,N_2019);
and U2097 (N_2097,N_2042,N_2026);
and U2098 (N_2098,N_2017,N_2046);
nand U2099 (N_2099,N_2031,N_2019);
and U2100 (N_2100,N_2078,N_2085);
and U2101 (N_2101,N_2098,N_2052);
or U2102 (N_2102,N_2055,N_2089);
nand U2103 (N_2103,N_2082,N_2080);
nor U2104 (N_2104,N_2077,N_2096);
or U2105 (N_2105,N_2050,N_2065);
nor U2106 (N_2106,N_2092,N_2069);
nor U2107 (N_2107,N_2088,N_2070);
and U2108 (N_2108,N_2075,N_2063);
nor U2109 (N_2109,N_2060,N_2058);
and U2110 (N_2110,N_2062,N_2054);
nor U2111 (N_2111,N_2067,N_2095);
xnor U2112 (N_2112,N_2087,N_2064);
and U2113 (N_2113,N_2061,N_2093);
and U2114 (N_2114,N_2074,N_2091);
or U2115 (N_2115,N_2059,N_2073);
and U2116 (N_2116,N_2094,N_2056);
nand U2117 (N_2117,N_2099,N_2086);
nand U2118 (N_2118,N_2066,N_2053);
xor U2119 (N_2119,N_2081,N_2068);
nor U2120 (N_2120,N_2057,N_2097);
nand U2121 (N_2121,N_2051,N_2079);
nand U2122 (N_2122,N_2084,N_2071);
nand U2123 (N_2123,N_2072,N_2076);
and U2124 (N_2124,N_2090,N_2083);
or U2125 (N_2125,N_2090,N_2092);
and U2126 (N_2126,N_2070,N_2051);
nand U2127 (N_2127,N_2089,N_2087);
or U2128 (N_2128,N_2066,N_2057);
or U2129 (N_2129,N_2072,N_2096);
nor U2130 (N_2130,N_2096,N_2082);
and U2131 (N_2131,N_2053,N_2091);
nand U2132 (N_2132,N_2051,N_2058);
nand U2133 (N_2133,N_2084,N_2096);
nand U2134 (N_2134,N_2093,N_2068);
and U2135 (N_2135,N_2059,N_2095);
and U2136 (N_2136,N_2054,N_2055);
or U2137 (N_2137,N_2096,N_2071);
or U2138 (N_2138,N_2099,N_2078);
nand U2139 (N_2139,N_2087,N_2081);
xor U2140 (N_2140,N_2080,N_2064);
and U2141 (N_2141,N_2053,N_2084);
nor U2142 (N_2142,N_2099,N_2064);
nor U2143 (N_2143,N_2070,N_2089);
or U2144 (N_2144,N_2072,N_2059);
or U2145 (N_2145,N_2064,N_2061);
xnor U2146 (N_2146,N_2082,N_2077);
and U2147 (N_2147,N_2057,N_2051);
nand U2148 (N_2148,N_2095,N_2074);
and U2149 (N_2149,N_2095,N_2068);
and U2150 (N_2150,N_2138,N_2126);
and U2151 (N_2151,N_2103,N_2121);
and U2152 (N_2152,N_2133,N_2107);
nand U2153 (N_2153,N_2147,N_2125);
nand U2154 (N_2154,N_2129,N_2106);
nor U2155 (N_2155,N_2122,N_2119);
or U2156 (N_2156,N_2141,N_2104);
or U2157 (N_2157,N_2117,N_2118);
and U2158 (N_2158,N_2149,N_2105);
xor U2159 (N_2159,N_2130,N_2110);
xor U2160 (N_2160,N_2144,N_2128);
and U2161 (N_2161,N_2115,N_2124);
or U2162 (N_2162,N_2100,N_2113);
or U2163 (N_2163,N_2146,N_2136);
xor U2164 (N_2164,N_2111,N_2131);
and U2165 (N_2165,N_2139,N_2134);
xor U2166 (N_2166,N_2140,N_2137);
or U2167 (N_2167,N_2109,N_2116);
nand U2168 (N_2168,N_2132,N_2135);
and U2169 (N_2169,N_2114,N_2108);
and U2170 (N_2170,N_2120,N_2148);
and U2171 (N_2171,N_2142,N_2101);
and U2172 (N_2172,N_2123,N_2145);
nor U2173 (N_2173,N_2127,N_2102);
nand U2174 (N_2174,N_2143,N_2112);
nor U2175 (N_2175,N_2147,N_2126);
or U2176 (N_2176,N_2111,N_2103);
nand U2177 (N_2177,N_2125,N_2110);
and U2178 (N_2178,N_2125,N_2141);
nor U2179 (N_2179,N_2105,N_2110);
and U2180 (N_2180,N_2103,N_2123);
and U2181 (N_2181,N_2114,N_2119);
xor U2182 (N_2182,N_2120,N_2107);
and U2183 (N_2183,N_2125,N_2103);
nor U2184 (N_2184,N_2148,N_2125);
nor U2185 (N_2185,N_2142,N_2126);
nand U2186 (N_2186,N_2142,N_2133);
nor U2187 (N_2187,N_2129,N_2126);
nor U2188 (N_2188,N_2100,N_2107);
nand U2189 (N_2189,N_2126,N_2108);
or U2190 (N_2190,N_2110,N_2148);
or U2191 (N_2191,N_2134,N_2148);
and U2192 (N_2192,N_2134,N_2123);
nor U2193 (N_2193,N_2113,N_2112);
or U2194 (N_2194,N_2118,N_2140);
nand U2195 (N_2195,N_2124,N_2129);
or U2196 (N_2196,N_2117,N_2133);
xor U2197 (N_2197,N_2118,N_2107);
nor U2198 (N_2198,N_2146,N_2113);
and U2199 (N_2199,N_2135,N_2110);
nand U2200 (N_2200,N_2171,N_2165);
nor U2201 (N_2201,N_2167,N_2194);
nand U2202 (N_2202,N_2195,N_2180);
and U2203 (N_2203,N_2160,N_2177);
and U2204 (N_2204,N_2153,N_2196);
and U2205 (N_2205,N_2162,N_2174);
nor U2206 (N_2206,N_2182,N_2166);
or U2207 (N_2207,N_2155,N_2154);
nor U2208 (N_2208,N_2184,N_2169);
nor U2209 (N_2209,N_2173,N_2158);
and U2210 (N_2210,N_2189,N_2197);
or U2211 (N_2211,N_2151,N_2152);
and U2212 (N_2212,N_2193,N_2164);
and U2213 (N_2213,N_2187,N_2163);
nor U2214 (N_2214,N_2159,N_2175);
or U2215 (N_2215,N_2181,N_2186);
xor U2216 (N_2216,N_2198,N_2179);
nand U2217 (N_2217,N_2176,N_2161);
nor U2218 (N_2218,N_2157,N_2191);
nor U2219 (N_2219,N_2156,N_2192);
nor U2220 (N_2220,N_2150,N_2199);
or U2221 (N_2221,N_2168,N_2183);
nor U2222 (N_2222,N_2172,N_2190);
and U2223 (N_2223,N_2170,N_2188);
or U2224 (N_2224,N_2185,N_2178);
nor U2225 (N_2225,N_2165,N_2189);
nor U2226 (N_2226,N_2191,N_2178);
and U2227 (N_2227,N_2188,N_2181);
and U2228 (N_2228,N_2168,N_2184);
or U2229 (N_2229,N_2185,N_2173);
and U2230 (N_2230,N_2170,N_2194);
and U2231 (N_2231,N_2178,N_2163);
nor U2232 (N_2232,N_2189,N_2158);
or U2233 (N_2233,N_2158,N_2196);
nand U2234 (N_2234,N_2167,N_2198);
and U2235 (N_2235,N_2157,N_2183);
or U2236 (N_2236,N_2193,N_2182);
and U2237 (N_2237,N_2189,N_2152);
or U2238 (N_2238,N_2182,N_2196);
nand U2239 (N_2239,N_2190,N_2171);
nand U2240 (N_2240,N_2176,N_2154);
or U2241 (N_2241,N_2151,N_2183);
nor U2242 (N_2242,N_2175,N_2155);
nor U2243 (N_2243,N_2197,N_2184);
nor U2244 (N_2244,N_2198,N_2159);
or U2245 (N_2245,N_2153,N_2183);
or U2246 (N_2246,N_2174,N_2192);
xnor U2247 (N_2247,N_2198,N_2154);
or U2248 (N_2248,N_2155,N_2198);
or U2249 (N_2249,N_2186,N_2198);
xnor U2250 (N_2250,N_2211,N_2231);
nand U2251 (N_2251,N_2219,N_2248);
and U2252 (N_2252,N_2237,N_2249);
nor U2253 (N_2253,N_2208,N_2246);
nor U2254 (N_2254,N_2210,N_2247);
or U2255 (N_2255,N_2242,N_2238);
nor U2256 (N_2256,N_2228,N_2244);
or U2257 (N_2257,N_2200,N_2240);
nand U2258 (N_2258,N_2217,N_2243);
or U2259 (N_2259,N_2204,N_2224);
nor U2260 (N_2260,N_2226,N_2239);
and U2261 (N_2261,N_2230,N_2232);
nor U2262 (N_2262,N_2236,N_2229);
nor U2263 (N_2263,N_2235,N_2212);
nand U2264 (N_2264,N_2223,N_2218);
or U2265 (N_2265,N_2209,N_2234);
or U2266 (N_2266,N_2205,N_2215);
and U2267 (N_2267,N_2233,N_2207);
or U2268 (N_2268,N_2202,N_2227);
nand U2269 (N_2269,N_2221,N_2216);
or U2270 (N_2270,N_2225,N_2214);
or U2271 (N_2271,N_2222,N_2220);
nor U2272 (N_2272,N_2245,N_2241);
or U2273 (N_2273,N_2206,N_2213);
and U2274 (N_2274,N_2201,N_2203);
xnor U2275 (N_2275,N_2205,N_2246);
and U2276 (N_2276,N_2216,N_2230);
nand U2277 (N_2277,N_2211,N_2242);
and U2278 (N_2278,N_2220,N_2240);
or U2279 (N_2279,N_2240,N_2245);
xor U2280 (N_2280,N_2211,N_2217);
or U2281 (N_2281,N_2238,N_2203);
nor U2282 (N_2282,N_2225,N_2248);
nor U2283 (N_2283,N_2218,N_2246);
nand U2284 (N_2284,N_2233,N_2208);
nand U2285 (N_2285,N_2224,N_2205);
or U2286 (N_2286,N_2225,N_2234);
or U2287 (N_2287,N_2217,N_2207);
nor U2288 (N_2288,N_2202,N_2213);
nor U2289 (N_2289,N_2219,N_2200);
nand U2290 (N_2290,N_2229,N_2249);
nor U2291 (N_2291,N_2215,N_2211);
or U2292 (N_2292,N_2215,N_2212);
and U2293 (N_2293,N_2212,N_2207);
and U2294 (N_2294,N_2244,N_2219);
or U2295 (N_2295,N_2217,N_2230);
and U2296 (N_2296,N_2201,N_2210);
and U2297 (N_2297,N_2249,N_2214);
or U2298 (N_2298,N_2241,N_2205);
nor U2299 (N_2299,N_2204,N_2245);
and U2300 (N_2300,N_2270,N_2295);
or U2301 (N_2301,N_2282,N_2251);
nor U2302 (N_2302,N_2258,N_2289);
nand U2303 (N_2303,N_2272,N_2261);
or U2304 (N_2304,N_2252,N_2250);
or U2305 (N_2305,N_2253,N_2273);
and U2306 (N_2306,N_2286,N_2263);
xnor U2307 (N_2307,N_2255,N_2294);
nor U2308 (N_2308,N_2254,N_2299);
or U2309 (N_2309,N_2268,N_2262);
or U2310 (N_2310,N_2283,N_2285);
nand U2311 (N_2311,N_2260,N_2293);
or U2312 (N_2312,N_2288,N_2265);
nand U2313 (N_2313,N_2276,N_2287);
nor U2314 (N_2314,N_2291,N_2284);
or U2315 (N_2315,N_2256,N_2267);
xnor U2316 (N_2316,N_2264,N_2274);
and U2317 (N_2317,N_2292,N_2257);
or U2318 (N_2318,N_2277,N_2271);
nor U2319 (N_2319,N_2281,N_2266);
xor U2320 (N_2320,N_2296,N_2269);
or U2321 (N_2321,N_2290,N_2280);
xnor U2322 (N_2322,N_2279,N_2298);
and U2323 (N_2323,N_2259,N_2278);
nor U2324 (N_2324,N_2297,N_2275);
nor U2325 (N_2325,N_2271,N_2260);
and U2326 (N_2326,N_2251,N_2276);
xor U2327 (N_2327,N_2261,N_2250);
xor U2328 (N_2328,N_2279,N_2274);
and U2329 (N_2329,N_2252,N_2276);
and U2330 (N_2330,N_2270,N_2275);
nor U2331 (N_2331,N_2287,N_2296);
and U2332 (N_2332,N_2299,N_2287);
xnor U2333 (N_2333,N_2284,N_2288);
or U2334 (N_2334,N_2269,N_2276);
or U2335 (N_2335,N_2257,N_2254);
nor U2336 (N_2336,N_2284,N_2251);
or U2337 (N_2337,N_2264,N_2295);
nand U2338 (N_2338,N_2292,N_2263);
nor U2339 (N_2339,N_2282,N_2279);
nand U2340 (N_2340,N_2286,N_2297);
and U2341 (N_2341,N_2257,N_2290);
xnor U2342 (N_2342,N_2267,N_2266);
nor U2343 (N_2343,N_2271,N_2289);
nand U2344 (N_2344,N_2259,N_2285);
xor U2345 (N_2345,N_2288,N_2266);
nor U2346 (N_2346,N_2284,N_2266);
and U2347 (N_2347,N_2280,N_2258);
nand U2348 (N_2348,N_2265,N_2290);
nor U2349 (N_2349,N_2289,N_2283);
or U2350 (N_2350,N_2340,N_2301);
or U2351 (N_2351,N_2342,N_2339);
and U2352 (N_2352,N_2320,N_2316);
and U2353 (N_2353,N_2338,N_2337);
or U2354 (N_2354,N_2304,N_2312);
and U2355 (N_2355,N_2319,N_2331);
and U2356 (N_2356,N_2332,N_2303);
nor U2357 (N_2357,N_2344,N_2335);
xor U2358 (N_2358,N_2322,N_2323);
or U2359 (N_2359,N_2305,N_2326);
and U2360 (N_2360,N_2309,N_2308);
nor U2361 (N_2361,N_2327,N_2347);
nand U2362 (N_2362,N_2349,N_2314);
and U2363 (N_2363,N_2302,N_2315);
nand U2364 (N_2364,N_2345,N_2329);
and U2365 (N_2365,N_2313,N_2324);
nor U2366 (N_2366,N_2348,N_2311);
xor U2367 (N_2367,N_2325,N_2336);
and U2368 (N_2368,N_2334,N_2346);
and U2369 (N_2369,N_2343,N_2328);
nor U2370 (N_2370,N_2333,N_2310);
or U2371 (N_2371,N_2307,N_2318);
and U2372 (N_2372,N_2321,N_2306);
xor U2373 (N_2373,N_2341,N_2330);
xnor U2374 (N_2374,N_2300,N_2317);
or U2375 (N_2375,N_2343,N_2310);
xnor U2376 (N_2376,N_2316,N_2317);
or U2377 (N_2377,N_2312,N_2321);
nor U2378 (N_2378,N_2310,N_2315);
nor U2379 (N_2379,N_2320,N_2342);
nor U2380 (N_2380,N_2339,N_2331);
nor U2381 (N_2381,N_2306,N_2337);
and U2382 (N_2382,N_2318,N_2336);
nor U2383 (N_2383,N_2338,N_2313);
xor U2384 (N_2384,N_2308,N_2315);
xor U2385 (N_2385,N_2321,N_2317);
and U2386 (N_2386,N_2326,N_2304);
nor U2387 (N_2387,N_2333,N_2349);
and U2388 (N_2388,N_2328,N_2321);
and U2389 (N_2389,N_2322,N_2331);
nand U2390 (N_2390,N_2344,N_2306);
and U2391 (N_2391,N_2314,N_2309);
nand U2392 (N_2392,N_2308,N_2305);
nand U2393 (N_2393,N_2333,N_2315);
or U2394 (N_2394,N_2326,N_2337);
and U2395 (N_2395,N_2335,N_2321);
nor U2396 (N_2396,N_2349,N_2343);
nand U2397 (N_2397,N_2333,N_2345);
nor U2398 (N_2398,N_2317,N_2348);
and U2399 (N_2399,N_2310,N_2330);
nand U2400 (N_2400,N_2390,N_2371);
and U2401 (N_2401,N_2363,N_2364);
or U2402 (N_2402,N_2368,N_2370);
xor U2403 (N_2403,N_2377,N_2395);
xor U2404 (N_2404,N_2385,N_2379);
nand U2405 (N_2405,N_2375,N_2356);
xor U2406 (N_2406,N_2391,N_2352);
and U2407 (N_2407,N_2369,N_2398);
nor U2408 (N_2408,N_2383,N_2365);
nand U2409 (N_2409,N_2372,N_2378);
and U2410 (N_2410,N_2399,N_2382);
xor U2411 (N_2411,N_2350,N_2393);
and U2412 (N_2412,N_2387,N_2386);
or U2413 (N_2413,N_2366,N_2380);
xnor U2414 (N_2414,N_2389,N_2384);
and U2415 (N_2415,N_2381,N_2388);
nand U2416 (N_2416,N_2353,N_2357);
or U2417 (N_2417,N_2361,N_2392);
or U2418 (N_2418,N_2394,N_2396);
nand U2419 (N_2419,N_2374,N_2354);
nor U2420 (N_2420,N_2373,N_2367);
nor U2421 (N_2421,N_2358,N_2397);
nor U2422 (N_2422,N_2359,N_2362);
nor U2423 (N_2423,N_2360,N_2351);
or U2424 (N_2424,N_2355,N_2376);
nor U2425 (N_2425,N_2353,N_2382);
or U2426 (N_2426,N_2367,N_2361);
nand U2427 (N_2427,N_2354,N_2380);
nor U2428 (N_2428,N_2390,N_2354);
and U2429 (N_2429,N_2356,N_2365);
and U2430 (N_2430,N_2368,N_2386);
xnor U2431 (N_2431,N_2374,N_2356);
nor U2432 (N_2432,N_2397,N_2366);
xor U2433 (N_2433,N_2377,N_2364);
nor U2434 (N_2434,N_2350,N_2357);
nand U2435 (N_2435,N_2375,N_2390);
nand U2436 (N_2436,N_2362,N_2389);
and U2437 (N_2437,N_2351,N_2367);
nand U2438 (N_2438,N_2359,N_2391);
or U2439 (N_2439,N_2350,N_2376);
nor U2440 (N_2440,N_2352,N_2353);
or U2441 (N_2441,N_2367,N_2362);
nor U2442 (N_2442,N_2379,N_2378);
xor U2443 (N_2443,N_2356,N_2362);
nand U2444 (N_2444,N_2351,N_2361);
or U2445 (N_2445,N_2390,N_2383);
nand U2446 (N_2446,N_2387,N_2369);
and U2447 (N_2447,N_2397,N_2398);
or U2448 (N_2448,N_2377,N_2383);
or U2449 (N_2449,N_2367,N_2370);
or U2450 (N_2450,N_2448,N_2434);
nand U2451 (N_2451,N_2421,N_2426);
or U2452 (N_2452,N_2440,N_2415);
xor U2453 (N_2453,N_2429,N_2407);
xnor U2454 (N_2454,N_2436,N_2444);
xnor U2455 (N_2455,N_2408,N_2441);
nand U2456 (N_2456,N_2420,N_2423);
nor U2457 (N_2457,N_2424,N_2437);
and U2458 (N_2458,N_2404,N_2403);
nand U2459 (N_2459,N_2438,N_2400);
xnor U2460 (N_2460,N_2442,N_2425);
nand U2461 (N_2461,N_2449,N_2418);
or U2462 (N_2462,N_2446,N_2428);
and U2463 (N_2463,N_2412,N_2422);
nand U2464 (N_2464,N_2431,N_2406);
and U2465 (N_2465,N_2405,N_2413);
nand U2466 (N_2466,N_2427,N_2443);
and U2467 (N_2467,N_2430,N_2416);
and U2468 (N_2468,N_2410,N_2401);
xnor U2469 (N_2469,N_2419,N_2414);
and U2470 (N_2470,N_2411,N_2433);
xnor U2471 (N_2471,N_2432,N_2447);
nor U2472 (N_2472,N_2402,N_2417);
and U2473 (N_2473,N_2409,N_2439);
and U2474 (N_2474,N_2435,N_2445);
nand U2475 (N_2475,N_2420,N_2447);
and U2476 (N_2476,N_2432,N_2449);
nor U2477 (N_2477,N_2430,N_2400);
and U2478 (N_2478,N_2427,N_2401);
or U2479 (N_2479,N_2430,N_2406);
and U2480 (N_2480,N_2444,N_2431);
nand U2481 (N_2481,N_2443,N_2419);
nor U2482 (N_2482,N_2436,N_2438);
and U2483 (N_2483,N_2406,N_2405);
and U2484 (N_2484,N_2419,N_2412);
or U2485 (N_2485,N_2426,N_2427);
nand U2486 (N_2486,N_2402,N_2441);
or U2487 (N_2487,N_2439,N_2402);
or U2488 (N_2488,N_2417,N_2407);
xnor U2489 (N_2489,N_2418,N_2410);
or U2490 (N_2490,N_2432,N_2420);
and U2491 (N_2491,N_2432,N_2440);
xnor U2492 (N_2492,N_2415,N_2446);
and U2493 (N_2493,N_2437,N_2421);
xor U2494 (N_2494,N_2441,N_2401);
nand U2495 (N_2495,N_2400,N_2446);
or U2496 (N_2496,N_2423,N_2407);
nand U2497 (N_2497,N_2446,N_2449);
and U2498 (N_2498,N_2421,N_2433);
or U2499 (N_2499,N_2405,N_2402);
nor U2500 (N_2500,N_2466,N_2494);
nand U2501 (N_2501,N_2451,N_2453);
and U2502 (N_2502,N_2487,N_2483);
and U2503 (N_2503,N_2455,N_2473);
xor U2504 (N_2504,N_2468,N_2452);
or U2505 (N_2505,N_2490,N_2462);
nor U2506 (N_2506,N_2459,N_2492);
and U2507 (N_2507,N_2481,N_2464);
nor U2508 (N_2508,N_2478,N_2465);
or U2509 (N_2509,N_2499,N_2456);
nor U2510 (N_2510,N_2482,N_2488);
nor U2511 (N_2511,N_2463,N_2454);
or U2512 (N_2512,N_2458,N_2484);
or U2513 (N_2513,N_2470,N_2491);
and U2514 (N_2514,N_2475,N_2480);
nor U2515 (N_2515,N_2493,N_2471);
and U2516 (N_2516,N_2460,N_2469);
or U2517 (N_2517,N_2457,N_2496);
xor U2518 (N_2518,N_2461,N_2472);
or U2519 (N_2519,N_2474,N_2486);
nand U2520 (N_2520,N_2495,N_2467);
and U2521 (N_2521,N_2489,N_2497);
and U2522 (N_2522,N_2476,N_2479);
and U2523 (N_2523,N_2477,N_2450);
and U2524 (N_2524,N_2498,N_2485);
or U2525 (N_2525,N_2482,N_2489);
nor U2526 (N_2526,N_2471,N_2467);
and U2527 (N_2527,N_2474,N_2463);
xor U2528 (N_2528,N_2454,N_2487);
nor U2529 (N_2529,N_2466,N_2481);
or U2530 (N_2530,N_2488,N_2476);
and U2531 (N_2531,N_2496,N_2472);
nor U2532 (N_2532,N_2491,N_2474);
nand U2533 (N_2533,N_2472,N_2458);
nor U2534 (N_2534,N_2481,N_2495);
or U2535 (N_2535,N_2455,N_2486);
nor U2536 (N_2536,N_2479,N_2464);
and U2537 (N_2537,N_2468,N_2495);
or U2538 (N_2538,N_2450,N_2467);
nor U2539 (N_2539,N_2461,N_2459);
nand U2540 (N_2540,N_2497,N_2491);
xor U2541 (N_2541,N_2459,N_2466);
nor U2542 (N_2542,N_2469,N_2483);
nor U2543 (N_2543,N_2487,N_2484);
nor U2544 (N_2544,N_2491,N_2465);
xor U2545 (N_2545,N_2465,N_2455);
or U2546 (N_2546,N_2487,N_2476);
and U2547 (N_2547,N_2477,N_2462);
or U2548 (N_2548,N_2465,N_2493);
nor U2549 (N_2549,N_2455,N_2479);
and U2550 (N_2550,N_2512,N_2515);
and U2551 (N_2551,N_2521,N_2531);
and U2552 (N_2552,N_2544,N_2530);
and U2553 (N_2553,N_2541,N_2523);
nand U2554 (N_2554,N_2528,N_2532);
and U2555 (N_2555,N_2534,N_2509);
nand U2556 (N_2556,N_2547,N_2539);
or U2557 (N_2557,N_2548,N_2510);
nor U2558 (N_2558,N_2517,N_2507);
or U2559 (N_2559,N_2519,N_2529);
and U2560 (N_2560,N_2536,N_2502);
or U2561 (N_2561,N_2520,N_2511);
or U2562 (N_2562,N_2545,N_2535);
or U2563 (N_2563,N_2527,N_2516);
nand U2564 (N_2564,N_2506,N_2543);
or U2565 (N_2565,N_2505,N_2501);
and U2566 (N_2566,N_2522,N_2537);
or U2567 (N_2567,N_2525,N_2504);
xnor U2568 (N_2568,N_2526,N_2538);
nor U2569 (N_2569,N_2503,N_2508);
and U2570 (N_2570,N_2514,N_2524);
nor U2571 (N_2571,N_2542,N_2518);
or U2572 (N_2572,N_2513,N_2546);
or U2573 (N_2573,N_2540,N_2533);
nor U2574 (N_2574,N_2549,N_2500);
or U2575 (N_2575,N_2548,N_2530);
nor U2576 (N_2576,N_2542,N_2509);
or U2577 (N_2577,N_2516,N_2504);
and U2578 (N_2578,N_2540,N_2515);
or U2579 (N_2579,N_2517,N_2502);
and U2580 (N_2580,N_2515,N_2509);
and U2581 (N_2581,N_2539,N_2525);
xnor U2582 (N_2582,N_2538,N_2510);
or U2583 (N_2583,N_2543,N_2541);
nand U2584 (N_2584,N_2511,N_2504);
and U2585 (N_2585,N_2549,N_2519);
xnor U2586 (N_2586,N_2527,N_2513);
xor U2587 (N_2587,N_2544,N_2547);
or U2588 (N_2588,N_2500,N_2525);
nand U2589 (N_2589,N_2542,N_2521);
and U2590 (N_2590,N_2543,N_2505);
nand U2591 (N_2591,N_2507,N_2545);
nor U2592 (N_2592,N_2540,N_2542);
nand U2593 (N_2593,N_2504,N_2534);
xor U2594 (N_2594,N_2516,N_2522);
nand U2595 (N_2595,N_2511,N_2519);
xnor U2596 (N_2596,N_2501,N_2521);
or U2597 (N_2597,N_2523,N_2502);
or U2598 (N_2598,N_2519,N_2532);
or U2599 (N_2599,N_2512,N_2534);
nand U2600 (N_2600,N_2594,N_2590);
xor U2601 (N_2601,N_2587,N_2564);
xnor U2602 (N_2602,N_2553,N_2550);
xnor U2603 (N_2603,N_2579,N_2578);
nand U2604 (N_2604,N_2561,N_2567);
or U2605 (N_2605,N_2568,N_2556);
xor U2606 (N_2606,N_2562,N_2554);
nand U2607 (N_2607,N_2584,N_2597);
and U2608 (N_2608,N_2570,N_2558);
and U2609 (N_2609,N_2566,N_2582);
nand U2610 (N_2610,N_2595,N_2551);
nor U2611 (N_2611,N_2565,N_2571);
and U2612 (N_2612,N_2588,N_2585);
nor U2613 (N_2613,N_2576,N_2569);
nand U2614 (N_2614,N_2592,N_2573);
nor U2615 (N_2615,N_2591,N_2574);
and U2616 (N_2616,N_2560,N_2555);
xor U2617 (N_2617,N_2598,N_2581);
and U2618 (N_2618,N_2577,N_2552);
or U2619 (N_2619,N_2589,N_2575);
and U2620 (N_2620,N_2596,N_2557);
and U2621 (N_2621,N_2593,N_2586);
nand U2622 (N_2622,N_2559,N_2563);
xor U2623 (N_2623,N_2583,N_2572);
nand U2624 (N_2624,N_2580,N_2599);
xor U2625 (N_2625,N_2561,N_2571);
nor U2626 (N_2626,N_2562,N_2584);
nand U2627 (N_2627,N_2579,N_2550);
nand U2628 (N_2628,N_2580,N_2577);
nand U2629 (N_2629,N_2592,N_2597);
nor U2630 (N_2630,N_2553,N_2590);
and U2631 (N_2631,N_2588,N_2567);
nor U2632 (N_2632,N_2569,N_2564);
nor U2633 (N_2633,N_2587,N_2559);
nand U2634 (N_2634,N_2589,N_2572);
xnor U2635 (N_2635,N_2563,N_2588);
and U2636 (N_2636,N_2583,N_2557);
and U2637 (N_2637,N_2593,N_2581);
nand U2638 (N_2638,N_2579,N_2595);
and U2639 (N_2639,N_2556,N_2580);
or U2640 (N_2640,N_2559,N_2588);
and U2641 (N_2641,N_2566,N_2553);
or U2642 (N_2642,N_2565,N_2570);
xor U2643 (N_2643,N_2572,N_2553);
xor U2644 (N_2644,N_2570,N_2584);
nand U2645 (N_2645,N_2598,N_2577);
nand U2646 (N_2646,N_2576,N_2556);
and U2647 (N_2647,N_2596,N_2598);
and U2648 (N_2648,N_2569,N_2554);
xnor U2649 (N_2649,N_2572,N_2570);
and U2650 (N_2650,N_2622,N_2609);
and U2651 (N_2651,N_2623,N_2641);
nor U2652 (N_2652,N_2616,N_2645);
xor U2653 (N_2653,N_2606,N_2614);
and U2654 (N_2654,N_2608,N_2602);
or U2655 (N_2655,N_2628,N_2644);
or U2656 (N_2656,N_2620,N_2640);
or U2657 (N_2657,N_2600,N_2617);
and U2658 (N_2658,N_2630,N_2607);
nand U2659 (N_2659,N_2603,N_2629);
or U2660 (N_2660,N_2634,N_2631);
nand U2661 (N_2661,N_2646,N_2613);
or U2662 (N_2662,N_2612,N_2636);
nor U2663 (N_2663,N_2615,N_2649);
and U2664 (N_2664,N_2632,N_2611);
nor U2665 (N_2665,N_2626,N_2601);
nor U2666 (N_2666,N_2635,N_2621);
or U2667 (N_2667,N_2638,N_2605);
nand U2668 (N_2668,N_2604,N_2624);
nand U2669 (N_2669,N_2647,N_2642);
nand U2670 (N_2670,N_2619,N_2637);
xnor U2671 (N_2671,N_2633,N_2610);
or U2672 (N_2672,N_2648,N_2627);
and U2673 (N_2673,N_2625,N_2639);
nand U2674 (N_2674,N_2643,N_2618);
xor U2675 (N_2675,N_2616,N_2612);
or U2676 (N_2676,N_2612,N_2615);
or U2677 (N_2677,N_2623,N_2636);
nor U2678 (N_2678,N_2619,N_2625);
and U2679 (N_2679,N_2640,N_2607);
and U2680 (N_2680,N_2629,N_2605);
and U2681 (N_2681,N_2616,N_2606);
and U2682 (N_2682,N_2618,N_2609);
and U2683 (N_2683,N_2615,N_2603);
or U2684 (N_2684,N_2605,N_2642);
or U2685 (N_2685,N_2602,N_2627);
nor U2686 (N_2686,N_2605,N_2604);
nand U2687 (N_2687,N_2609,N_2644);
nor U2688 (N_2688,N_2636,N_2606);
nor U2689 (N_2689,N_2608,N_2617);
nor U2690 (N_2690,N_2635,N_2614);
nor U2691 (N_2691,N_2611,N_2637);
and U2692 (N_2692,N_2638,N_2616);
nor U2693 (N_2693,N_2624,N_2642);
and U2694 (N_2694,N_2612,N_2644);
nand U2695 (N_2695,N_2608,N_2647);
nand U2696 (N_2696,N_2645,N_2612);
xnor U2697 (N_2697,N_2608,N_2636);
and U2698 (N_2698,N_2612,N_2633);
nor U2699 (N_2699,N_2622,N_2608);
and U2700 (N_2700,N_2676,N_2669);
and U2701 (N_2701,N_2696,N_2650);
xor U2702 (N_2702,N_2663,N_2699);
and U2703 (N_2703,N_2657,N_2688);
nor U2704 (N_2704,N_2667,N_2677);
nor U2705 (N_2705,N_2670,N_2674);
nor U2706 (N_2706,N_2671,N_2685);
nand U2707 (N_2707,N_2681,N_2675);
nor U2708 (N_2708,N_2656,N_2654);
xnor U2709 (N_2709,N_2662,N_2659);
and U2710 (N_2710,N_2682,N_2678);
and U2711 (N_2711,N_2664,N_2665);
nand U2712 (N_2712,N_2698,N_2652);
nor U2713 (N_2713,N_2673,N_2655);
and U2714 (N_2714,N_2668,N_2660);
or U2715 (N_2715,N_2661,N_2680);
nand U2716 (N_2716,N_2694,N_2684);
and U2717 (N_2717,N_2672,N_2695);
or U2718 (N_2718,N_2666,N_2653);
nor U2719 (N_2719,N_2697,N_2693);
or U2720 (N_2720,N_2658,N_2686);
nor U2721 (N_2721,N_2683,N_2679);
nand U2722 (N_2722,N_2687,N_2689);
and U2723 (N_2723,N_2691,N_2692);
or U2724 (N_2724,N_2651,N_2690);
and U2725 (N_2725,N_2682,N_2677);
and U2726 (N_2726,N_2677,N_2661);
nand U2727 (N_2727,N_2679,N_2667);
nor U2728 (N_2728,N_2657,N_2687);
and U2729 (N_2729,N_2674,N_2650);
and U2730 (N_2730,N_2685,N_2687);
nand U2731 (N_2731,N_2653,N_2699);
nand U2732 (N_2732,N_2698,N_2696);
and U2733 (N_2733,N_2695,N_2674);
or U2734 (N_2734,N_2652,N_2694);
and U2735 (N_2735,N_2698,N_2661);
nand U2736 (N_2736,N_2665,N_2663);
nand U2737 (N_2737,N_2671,N_2695);
nor U2738 (N_2738,N_2691,N_2678);
or U2739 (N_2739,N_2673,N_2674);
nor U2740 (N_2740,N_2666,N_2671);
xor U2741 (N_2741,N_2697,N_2653);
nor U2742 (N_2742,N_2675,N_2651);
or U2743 (N_2743,N_2687,N_2661);
or U2744 (N_2744,N_2660,N_2696);
nand U2745 (N_2745,N_2695,N_2658);
nand U2746 (N_2746,N_2652,N_2680);
or U2747 (N_2747,N_2686,N_2689);
nor U2748 (N_2748,N_2657,N_2677);
nor U2749 (N_2749,N_2677,N_2686);
nor U2750 (N_2750,N_2723,N_2726);
nor U2751 (N_2751,N_2739,N_2749);
xor U2752 (N_2752,N_2729,N_2701);
and U2753 (N_2753,N_2741,N_2716);
and U2754 (N_2754,N_2732,N_2721);
nor U2755 (N_2755,N_2713,N_2711);
nand U2756 (N_2756,N_2703,N_2747);
nand U2757 (N_2757,N_2706,N_2709);
and U2758 (N_2758,N_2717,N_2710);
nand U2759 (N_2759,N_2733,N_2724);
and U2760 (N_2760,N_2712,N_2728);
and U2761 (N_2761,N_2704,N_2745);
nand U2762 (N_2762,N_2746,N_2730);
and U2763 (N_2763,N_2702,N_2736);
or U2764 (N_2764,N_2725,N_2743);
and U2765 (N_2765,N_2708,N_2714);
or U2766 (N_2766,N_2718,N_2715);
nand U2767 (N_2767,N_2731,N_2700);
nor U2768 (N_2768,N_2705,N_2742);
or U2769 (N_2769,N_2727,N_2744);
xnor U2770 (N_2770,N_2737,N_2740);
and U2771 (N_2771,N_2735,N_2748);
nor U2772 (N_2772,N_2734,N_2707);
or U2773 (N_2773,N_2738,N_2719);
or U2774 (N_2774,N_2722,N_2720);
or U2775 (N_2775,N_2748,N_2726);
and U2776 (N_2776,N_2740,N_2727);
and U2777 (N_2777,N_2742,N_2709);
and U2778 (N_2778,N_2717,N_2744);
nor U2779 (N_2779,N_2711,N_2700);
or U2780 (N_2780,N_2749,N_2746);
nand U2781 (N_2781,N_2740,N_2749);
or U2782 (N_2782,N_2748,N_2729);
nand U2783 (N_2783,N_2734,N_2727);
xnor U2784 (N_2784,N_2744,N_2714);
and U2785 (N_2785,N_2705,N_2720);
nor U2786 (N_2786,N_2729,N_2705);
xor U2787 (N_2787,N_2719,N_2742);
nor U2788 (N_2788,N_2742,N_2704);
nor U2789 (N_2789,N_2744,N_2728);
and U2790 (N_2790,N_2737,N_2713);
and U2791 (N_2791,N_2709,N_2738);
nand U2792 (N_2792,N_2705,N_2708);
nand U2793 (N_2793,N_2744,N_2735);
nand U2794 (N_2794,N_2740,N_2709);
xor U2795 (N_2795,N_2749,N_2714);
xor U2796 (N_2796,N_2703,N_2740);
or U2797 (N_2797,N_2710,N_2712);
nor U2798 (N_2798,N_2710,N_2739);
nor U2799 (N_2799,N_2721,N_2714);
nand U2800 (N_2800,N_2753,N_2798);
nor U2801 (N_2801,N_2766,N_2785);
nor U2802 (N_2802,N_2768,N_2770);
nor U2803 (N_2803,N_2755,N_2752);
nand U2804 (N_2804,N_2791,N_2760);
and U2805 (N_2805,N_2782,N_2778);
and U2806 (N_2806,N_2796,N_2767);
nor U2807 (N_2807,N_2773,N_2771);
and U2808 (N_2808,N_2777,N_2775);
nor U2809 (N_2809,N_2799,N_2790);
or U2810 (N_2810,N_2769,N_2758);
or U2811 (N_2811,N_2750,N_2797);
xnor U2812 (N_2812,N_2774,N_2780);
nand U2813 (N_2813,N_2756,N_2793);
and U2814 (N_2814,N_2787,N_2794);
nand U2815 (N_2815,N_2776,N_2759);
or U2816 (N_2816,N_2792,N_2788);
nor U2817 (N_2817,N_2779,N_2751);
nor U2818 (N_2818,N_2789,N_2795);
xor U2819 (N_2819,N_2783,N_2786);
nor U2820 (N_2820,N_2764,N_2772);
xnor U2821 (N_2821,N_2784,N_2781);
xor U2822 (N_2822,N_2762,N_2754);
nand U2823 (N_2823,N_2761,N_2757);
and U2824 (N_2824,N_2763,N_2765);
or U2825 (N_2825,N_2755,N_2793);
or U2826 (N_2826,N_2753,N_2754);
and U2827 (N_2827,N_2797,N_2771);
nand U2828 (N_2828,N_2768,N_2775);
and U2829 (N_2829,N_2799,N_2791);
nand U2830 (N_2830,N_2793,N_2763);
or U2831 (N_2831,N_2771,N_2768);
or U2832 (N_2832,N_2790,N_2791);
nor U2833 (N_2833,N_2777,N_2754);
and U2834 (N_2834,N_2794,N_2779);
or U2835 (N_2835,N_2789,N_2766);
or U2836 (N_2836,N_2778,N_2757);
or U2837 (N_2837,N_2784,N_2792);
and U2838 (N_2838,N_2750,N_2783);
nand U2839 (N_2839,N_2778,N_2797);
nand U2840 (N_2840,N_2769,N_2785);
or U2841 (N_2841,N_2750,N_2774);
or U2842 (N_2842,N_2786,N_2753);
or U2843 (N_2843,N_2759,N_2758);
nor U2844 (N_2844,N_2784,N_2798);
nand U2845 (N_2845,N_2789,N_2771);
and U2846 (N_2846,N_2764,N_2784);
or U2847 (N_2847,N_2797,N_2763);
or U2848 (N_2848,N_2782,N_2799);
nand U2849 (N_2849,N_2794,N_2789);
and U2850 (N_2850,N_2813,N_2826);
nor U2851 (N_2851,N_2847,N_2810);
and U2852 (N_2852,N_2817,N_2841);
nand U2853 (N_2853,N_2825,N_2842);
or U2854 (N_2854,N_2836,N_2815);
or U2855 (N_2855,N_2829,N_2831);
and U2856 (N_2856,N_2803,N_2848);
nand U2857 (N_2857,N_2802,N_2820);
xor U2858 (N_2858,N_2814,N_2824);
or U2859 (N_2859,N_2818,N_2812);
and U2860 (N_2860,N_2830,N_2805);
and U2861 (N_2861,N_2833,N_2808);
and U2862 (N_2862,N_2800,N_2846);
nand U2863 (N_2863,N_2823,N_2809);
nor U2864 (N_2864,N_2822,N_2839);
or U2865 (N_2865,N_2845,N_2828);
nand U2866 (N_2866,N_2837,N_2843);
or U2867 (N_2867,N_2821,N_2827);
xor U2868 (N_2868,N_2816,N_2834);
nand U2869 (N_2869,N_2811,N_2806);
and U2870 (N_2870,N_2801,N_2807);
and U2871 (N_2871,N_2804,N_2838);
nor U2872 (N_2872,N_2840,N_2832);
nand U2873 (N_2873,N_2819,N_2849);
and U2874 (N_2874,N_2844,N_2835);
and U2875 (N_2875,N_2815,N_2832);
nand U2876 (N_2876,N_2830,N_2811);
and U2877 (N_2877,N_2834,N_2818);
xnor U2878 (N_2878,N_2826,N_2836);
nand U2879 (N_2879,N_2823,N_2813);
nor U2880 (N_2880,N_2800,N_2843);
nor U2881 (N_2881,N_2827,N_2818);
nand U2882 (N_2882,N_2813,N_2800);
nand U2883 (N_2883,N_2837,N_2807);
and U2884 (N_2884,N_2829,N_2848);
nor U2885 (N_2885,N_2808,N_2844);
nand U2886 (N_2886,N_2842,N_2803);
nor U2887 (N_2887,N_2823,N_2824);
xor U2888 (N_2888,N_2822,N_2842);
nand U2889 (N_2889,N_2839,N_2824);
and U2890 (N_2890,N_2834,N_2827);
nor U2891 (N_2891,N_2830,N_2817);
nor U2892 (N_2892,N_2808,N_2821);
and U2893 (N_2893,N_2830,N_2813);
and U2894 (N_2894,N_2843,N_2826);
nor U2895 (N_2895,N_2818,N_2840);
or U2896 (N_2896,N_2815,N_2820);
and U2897 (N_2897,N_2840,N_2823);
nor U2898 (N_2898,N_2829,N_2839);
nand U2899 (N_2899,N_2826,N_2816);
nand U2900 (N_2900,N_2875,N_2859);
and U2901 (N_2901,N_2884,N_2858);
nor U2902 (N_2902,N_2865,N_2893);
and U2903 (N_2903,N_2879,N_2895);
nand U2904 (N_2904,N_2885,N_2850);
or U2905 (N_2905,N_2890,N_2855);
nor U2906 (N_2906,N_2872,N_2869);
or U2907 (N_2907,N_2854,N_2876);
xnor U2908 (N_2908,N_2856,N_2857);
nor U2909 (N_2909,N_2898,N_2874);
nor U2910 (N_2910,N_2851,N_2897);
or U2911 (N_2911,N_2860,N_2878);
and U2912 (N_2912,N_2887,N_2896);
xnor U2913 (N_2913,N_2888,N_2881);
and U2914 (N_2914,N_2886,N_2868);
xor U2915 (N_2915,N_2871,N_2873);
xor U2916 (N_2916,N_2870,N_2861);
and U2917 (N_2917,N_2867,N_2892);
and U2918 (N_2918,N_2882,N_2866);
nand U2919 (N_2919,N_2877,N_2863);
or U2920 (N_2920,N_2880,N_2883);
and U2921 (N_2921,N_2852,N_2891);
nor U2922 (N_2922,N_2899,N_2864);
nor U2923 (N_2923,N_2862,N_2853);
or U2924 (N_2924,N_2889,N_2894);
nand U2925 (N_2925,N_2862,N_2855);
nand U2926 (N_2926,N_2850,N_2878);
nand U2927 (N_2927,N_2897,N_2881);
and U2928 (N_2928,N_2894,N_2850);
nor U2929 (N_2929,N_2878,N_2872);
nor U2930 (N_2930,N_2851,N_2894);
nor U2931 (N_2931,N_2892,N_2873);
nand U2932 (N_2932,N_2881,N_2860);
and U2933 (N_2933,N_2852,N_2859);
and U2934 (N_2934,N_2858,N_2890);
nor U2935 (N_2935,N_2877,N_2893);
nor U2936 (N_2936,N_2858,N_2852);
or U2937 (N_2937,N_2870,N_2869);
nor U2938 (N_2938,N_2877,N_2872);
and U2939 (N_2939,N_2892,N_2865);
xor U2940 (N_2940,N_2857,N_2860);
nand U2941 (N_2941,N_2882,N_2883);
and U2942 (N_2942,N_2888,N_2899);
xnor U2943 (N_2943,N_2878,N_2867);
nor U2944 (N_2944,N_2886,N_2870);
and U2945 (N_2945,N_2880,N_2886);
nand U2946 (N_2946,N_2871,N_2853);
or U2947 (N_2947,N_2857,N_2873);
or U2948 (N_2948,N_2886,N_2877);
or U2949 (N_2949,N_2867,N_2852);
or U2950 (N_2950,N_2904,N_2926);
or U2951 (N_2951,N_2924,N_2910);
nor U2952 (N_2952,N_2933,N_2945);
nor U2953 (N_2953,N_2917,N_2940);
or U2954 (N_2954,N_2909,N_2906);
nand U2955 (N_2955,N_2902,N_2915);
nand U2956 (N_2956,N_2948,N_2938);
or U2957 (N_2957,N_2932,N_2908);
nand U2958 (N_2958,N_2914,N_2912);
xnor U2959 (N_2959,N_2946,N_2928);
and U2960 (N_2960,N_2929,N_2911);
nand U2961 (N_2961,N_2947,N_2934);
and U2962 (N_2962,N_2944,N_2931);
and U2963 (N_2963,N_2916,N_2941);
nor U2964 (N_2964,N_2925,N_2918);
and U2965 (N_2965,N_2903,N_2927);
xor U2966 (N_2966,N_2930,N_2943);
nor U2967 (N_2967,N_2913,N_2923);
nor U2968 (N_2968,N_2936,N_2921);
nand U2969 (N_2969,N_2920,N_2905);
nor U2970 (N_2970,N_2939,N_2922);
nand U2971 (N_2971,N_2937,N_2907);
nand U2972 (N_2972,N_2942,N_2949);
xor U2973 (N_2973,N_2919,N_2900);
nand U2974 (N_2974,N_2901,N_2935);
nand U2975 (N_2975,N_2939,N_2943);
nand U2976 (N_2976,N_2906,N_2941);
or U2977 (N_2977,N_2928,N_2932);
and U2978 (N_2978,N_2930,N_2934);
nor U2979 (N_2979,N_2908,N_2901);
nand U2980 (N_2980,N_2920,N_2928);
xor U2981 (N_2981,N_2907,N_2911);
and U2982 (N_2982,N_2949,N_2922);
xnor U2983 (N_2983,N_2922,N_2921);
nor U2984 (N_2984,N_2925,N_2910);
and U2985 (N_2985,N_2929,N_2913);
nand U2986 (N_2986,N_2924,N_2909);
nor U2987 (N_2987,N_2929,N_2909);
nor U2988 (N_2988,N_2911,N_2940);
nor U2989 (N_2989,N_2949,N_2923);
nand U2990 (N_2990,N_2913,N_2920);
nand U2991 (N_2991,N_2946,N_2949);
and U2992 (N_2992,N_2930,N_2928);
nor U2993 (N_2993,N_2920,N_2914);
or U2994 (N_2994,N_2936,N_2909);
nand U2995 (N_2995,N_2916,N_2914);
nand U2996 (N_2996,N_2922,N_2927);
nor U2997 (N_2997,N_2902,N_2937);
nand U2998 (N_2998,N_2925,N_2919);
xor U2999 (N_2999,N_2948,N_2902);
and UO_0 (O_0,N_2966,N_2977);
nor UO_1 (O_1,N_2967,N_2976);
nor UO_2 (O_2,N_2981,N_2958);
nor UO_3 (O_3,N_2990,N_2956);
nor UO_4 (O_4,N_2971,N_2969);
nor UO_5 (O_5,N_2960,N_2972);
nand UO_6 (O_6,N_2964,N_2997);
nor UO_7 (O_7,N_2965,N_2985);
nand UO_8 (O_8,N_2952,N_2962);
and UO_9 (O_9,N_2979,N_2986);
and UO_10 (O_10,N_2951,N_2983);
and UO_11 (O_11,N_2980,N_2959);
xor UO_12 (O_12,N_2987,N_2995);
or UO_13 (O_13,N_2950,N_2970);
nand UO_14 (O_14,N_2996,N_2993);
nand UO_15 (O_15,N_2961,N_2955);
or UO_16 (O_16,N_2953,N_2991);
nand UO_17 (O_17,N_2978,N_2957);
and UO_18 (O_18,N_2999,N_2988);
nand UO_19 (O_19,N_2984,N_2989);
and UO_20 (O_20,N_2982,N_2994);
nand UO_21 (O_21,N_2974,N_2998);
or UO_22 (O_22,N_2954,N_2963);
nor UO_23 (O_23,N_2975,N_2968);
or UO_24 (O_24,N_2992,N_2973);
nand UO_25 (O_25,N_2970,N_2956);
or UO_26 (O_26,N_2975,N_2978);
and UO_27 (O_27,N_2966,N_2975);
and UO_28 (O_28,N_2963,N_2959);
and UO_29 (O_29,N_2980,N_2985);
nand UO_30 (O_30,N_2978,N_2973);
or UO_31 (O_31,N_2965,N_2979);
xnor UO_32 (O_32,N_2997,N_2956);
and UO_33 (O_33,N_2962,N_2992);
and UO_34 (O_34,N_2976,N_2970);
xor UO_35 (O_35,N_2962,N_2995);
nand UO_36 (O_36,N_2964,N_2979);
and UO_37 (O_37,N_2963,N_2957);
nand UO_38 (O_38,N_2958,N_2974);
nor UO_39 (O_39,N_2985,N_2972);
and UO_40 (O_40,N_2987,N_2955);
and UO_41 (O_41,N_2984,N_2979);
or UO_42 (O_42,N_2959,N_2967);
xor UO_43 (O_43,N_2991,N_2983);
nor UO_44 (O_44,N_2968,N_2974);
and UO_45 (O_45,N_2966,N_2967);
and UO_46 (O_46,N_2991,N_2994);
and UO_47 (O_47,N_2978,N_2982);
or UO_48 (O_48,N_2950,N_2979);
or UO_49 (O_49,N_2978,N_2990);
nor UO_50 (O_50,N_2997,N_2959);
or UO_51 (O_51,N_2954,N_2970);
xor UO_52 (O_52,N_2963,N_2988);
xor UO_53 (O_53,N_2987,N_2967);
nor UO_54 (O_54,N_2997,N_2998);
nor UO_55 (O_55,N_2990,N_2975);
nor UO_56 (O_56,N_2981,N_2968);
and UO_57 (O_57,N_2976,N_2983);
or UO_58 (O_58,N_2992,N_2985);
nor UO_59 (O_59,N_2976,N_2984);
nand UO_60 (O_60,N_2965,N_2980);
nand UO_61 (O_61,N_2976,N_2981);
xor UO_62 (O_62,N_2977,N_2961);
nand UO_63 (O_63,N_2993,N_2968);
nand UO_64 (O_64,N_2954,N_2964);
nor UO_65 (O_65,N_2974,N_2981);
nor UO_66 (O_66,N_2988,N_2991);
and UO_67 (O_67,N_2964,N_2994);
nor UO_68 (O_68,N_2952,N_2978);
nand UO_69 (O_69,N_2956,N_2966);
nor UO_70 (O_70,N_2952,N_2968);
and UO_71 (O_71,N_2969,N_2988);
or UO_72 (O_72,N_2967,N_2979);
nor UO_73 (O_73,N_2969,N_2952);
xnor UO_74 (O_74,N_2992,N_2995);
nand UO_75 (O_75,N_2988,N_2975);
nand UO_76 (O_76,N_2988,N_2950);
xor UO_77 (O_77,N_2980,N_2956);
or UO_78 (O_78,N_2979,N_2991);
nor UO_79 (O_79,N_2973,N_2988);
xor UO_80 (O_80,N_2984,N_2972);
nand UO_81 (O_81,N_2973,N_2965);
nand UO_82 (O_82,N_2955,N_2957);
xor UO_83 (O_83,N_2983,N_2950);
and UO_84 (O_84,N_2985,N_2983);
or UO_85 (O_85,N_2967,N_2992);
nand UO_86 (O_86,N_2967,N_2980);
and UO_87 (O_87,N_2984,N_2961);
and UO_88 (O_88,N_2981,N_2964);
nor UO_89 (O_89,N_2979,N_2957);
and UO_90 (O_90,N_2972,N_2976);
nand UO_91 (O_91,N_2999,N_2995);
and UO_92 (O_92,N_2951,N_2986);
nor UO_93 (O_93,N_2977,N_2968);
and UO_94 (O_94,N_2952,N_2981);
nand UO_95 (O_95,N_2986,N_2959);
nand UO_96 (O_96,N_2964,N_2961);
xnor UO_97 (O_97,N_2953,N_2995);
nand UO_98 (O_98,N_2967,N_2982);
and UO_99 (O_99,N_2987,N_2954);
or UO_100 (O_100,N_2983,N_2971);
or UO_101 (O_101,N_2998,N_2956);
or UO_102 (O_102,N_2961,N_2965);
nor UO_103 (O_103,N_2985,N_2957);
xnor UO_104 (O_104,N_2979,N_2966);
or UO_105 (O_105,N_2974,N_2953);
nand UO_106 (O_106,N_2984,N_2963);
nand UO_107 (O_107,N_2975,N_2986);
or UO_108 (O_108,N_2979,N_2989);
and UO_109 (O_109,N_2998,N_2970);
nand UO_110 (O_110,N_2952,N_2999);
nand UO_111 (O_111,N_2996,N_2966);
or UO_112 (O_112,N_2957,N_2964);
nor UO_113 (O_113,N_2981,N_2962);
and UO_114 (O_114,N_2982,N_2969);
nor UO_115 (O_115,N_2974,N_2954);
and UO_116 (O_116,N_2963,N_2974);
nand UO_117 (O_117,N_2964,N_2951);
or UO_118 (O_118,N_2951,N_2971);
or UO_119 (O_119,N_2997,N_2991);
or UO_120 (O_120,N_2986,N_2956);
nor UO_121 (O_121,N_2989,N_2974);
or UO_122 (O_122,N_2958,N_2983);
nor UO_123 (O_123,N_2961,N_2983);
and UO_124 (O_124,N_2994,N_2972);
nand UO_125 (O_125,N_2959,N_2983);
nor UO_126 (O_126,N_2993,N_2999);
xnor UO_127 (O_127,N_2954,N_2967);
nor UO_128 (O_128,N_2994,N_2966);
or UO_129 (O_129,N_2989,N_2965);
nand UO_130 (O_130,N_2966,N_2988);
nor UO_131 (O_131,N_2965,N_2991);
and UO_132 (O_132,N_2989,N_2960);
nand UO_133 (O_133,N_2984,N_2966);
and UO_134 (O_134,N_2976,N_2957);
or UO_135 (O_135,N_2969,N_2990);
and UO_136 (O_136,N_2954,N_2973);
or UO_137 (O_137,N_2951,N_2954);
nor UO_138 (O_138,N_2952,N_2995);
and UO_139 (O_139,N_2971,N_2966);
nor UO_140 (O_140,N_2952,N_2991);
and UO_141 (O_141,N_2991,N_2986);
nand UO_142 (O_142,N_2967,N_2981);
or UO_143 (O_143,N_2969,N_2967);
or UO_144 (O_144,N_2982,N_2956);
or UO_145 (O_145,N_2971,N_2950);
or UO_146 (O_146,N_2984,N_2974);
nor UO_147 (O_147,N_2997,N_2992);
nand UO_148 (O_148,N_2999,N_2969);
xnor UO_149 (O_149,N_2997,N_2967);
nor UO_150 (O_150,N_2982,N_2970);
or UO_151 (O_151,N_2962,N_2977);
or UO_152 (O_152,N_2959,N_2999);
nand UO_153 (O_153,N_2997,N_2962);
and UO_154 (O_154,N_2994,N_2996);
nor UO_155 (O_155,N_2959,N_2979);
or UO_156 (O_156,N_2985,N_2989);
and UO_157 (O_157,N_2977,N_2981);
or UO_158 (O_158,N_2991,N_2975);
nand UO_159 (O_159,N_2978,N_2956);
and UO_160 (O_160,N_2994,N_2990);
or UO_161 (O_161,N_2971,N_2998);
and UO_162 (O_162,N_2980,N_2955);
or UO_163 (O_163,N_2995,N_2997);
nand UO_164 (O_164,N_2952,N_2956);
or UO_165 (O_165,N_2963,N_2981);
nand UO_166 (O_166,N_2988,N_2965);
nor UO_167 (O_167,N_2987,N_2998);
or UO_168 (O_168,N_2976,N_2996);
nand UO_169 (O_169,N_2981,N_2970);
nand UO_170 (O_170,N_2977,N_2958);
xnor UO_171 (O_171,N_2979,N_2952);
and UO_172 (O_172,N_2969,N_2955);
nand UO_173 (O_173,N_2974,N_2967);
or UO_174 (O_174,N_2998,N_2955);
or UO_175 (O_175,N_2967,N_2956);
and UO_176 (O_176,N_2977,N_2957);
and UO_177 (O_177,N_2964,N_2962);
nand UO_178 (O_178,N_2975,N_2951);
nor UO_179 (O_179,N_2954,N_2985);
nor UO_180 (O_180,N_2974,N_2992);
xnor UO_181 (O_181,N_2979,N_2988);
nand UO_182 (O_182,N_2959,N_2952);
xnor UO_183 (O_183,N_2976,N_2991);
and UO_184 (O_184,N_2999,N_2961);
or UO_185 (O_185,N_2961,N_2952);
nand UO_186 (O_186,N_2970,N_2972);
xor UO_187 (O_187,N_2970,N_2993);
nand UO_188 (O_188,N_2976,N_2953);
nand UO_189 (O_189,N_2994,N_2986);
nor UO_190 (O_190,N_2993,N_2986);
or UO_191 (O_191,N_2959,N_2955);
xor UO_192 (O_192,N_2979,N_2978);
nor UO_193 (O_193,N_2960,N_2984);
xor UO_194 (O_194,N_2980,N_2950);
nor UO_195 (O_195,N_2980,N_2992);
and UO_196 (O_196,N_2977,N_2954);
nor UO_197 (O_197,N_2959,N_2998);
xor UO_198 (O_198,N_2989,N_2956);
or UO_199 (O_199,N_2978,N_2963);
and UO_200 (O_200,N_2974,N_2951);
and UO_201 (O_201,N_2973,N_2964);
xnor UO_202 (O_202,N_2982,N_2951);
or UO_203 (O_203,N_2988,N_2994);
nand UO_204 (O_204,N_2960,N_2961);
nor UO_205 (O_205,N_2969,N_2970);
or UO_206 (O_206,N_2977,N_2978);
nand UO_207 (O_207,N_2983,N_2964);
nand UO_208 (O_208,N_2984,N_2986);
and UO_209 (O_209,N_2982,N_2998);
and UO_210 (O_210,N_2956,N_2954);
and UO_211 (O_211,N_2997,N_2960);
xnor UO_212 (O_212,N_2987,N_2984);
and UO_213 (O_213,N_2951,N_2977);
nor UO_214 (O_214,N_2964,N_2987);
xnor UO_215 (O_215,N_2953,N_2970);
or UO_216 (O_216,N_2952,N_2976);
nor UO_217 (O_217,N_2987,N_2965);
nor UO_218 (O_218,N_2957,N_2984);
nand UO_219 (O_219,N_2953,N_2982);
or UO_220 (O_220,N_2983,N_2978);
nor UO_221 (O_221,N_2965,N_2993);
xnor UO_222 (O_222,N_2992,N_2999);
and UO_223 (O_223,N_2980,N_2979);
or UO_224 (O_224,N_2961,N_2966);
or UO_225 (O_225,N_2952,N_2975);
and UO_226 (O_226,N_2978,N_2961);
and UO_227 (O_227,N_2975,N_2979);
and UO_228 (O_228,N_2994,N_2967);
xor UO_229 (O_229,N_2992,N_2958);
and UO_230 (O_230,N_2993,N_2995);
nor UO_231 (O_231,N_2977,N_2998);
nand UO_232 (O_232,N_2965,N_2969);
nor UO_233 (O_233,N_2976,N_2968);
or UO_234 (O_234,N_2978,N_2987);
or UO_235 (O_235,N_2953,N_2984);
or UO_236 (O_236,N_2986,N_2966);
nand UO_237 (O_237,N_2989,N_2987);
nand UO_238 (O_238,N_2996,N_2979);
and UO_239 (O_239,N_2966,N_2952);
nand UO_240 (O_240,N_2989,N_2953);
nor UO_241 (O_241,N_2994,N_2951);
nand UO_242 (O_242,N_2957,N_2992);
nor UO_243 (O_243,N_2960,N_2957);
nand UO_244 (O_244,N_2964,N_2974);
and UO_245 (O_245,N_2978,N_2953);
or UO_246 (O_246,N_2971,N_2984);
nor UO_247 (O_247,N_2978,N_2968);
nand UO_248 (O_248,N_2992,N_2972);
or UO_249 (O_249,N_2999,N_2984);
nand UO_250 (O_250,N_2986,N_2961);
xor UO_251 (O_251,N_2970,N_2966);
or UO_252 (O_252,N_2982,N_2975);
nor UO_253 (O_253,N_2976,N_2985);
nand UO_254 (O_254,N_2989,N_2963);
nor UO_255 (O_255,N_2956,N_2984);
and UO_256 (O_256,N_2974,N_2959);
xor UO_257 (O_257,N_2979,N_2987);
nor UO_258 (O_258,N_2997,N_2957);
nor UO_259 (O_259,N_2990,N_2999);
or UO_260 (O_260,N_2958,N_2979);
nand UO_261 (O_261,N_2961,N_2990);
and UO_262 (O_262,N_2950,N_2974);
nor UO_263 (O_263,N_2982,N_2950);
and UO_264 (O_264,N_2986,N_2990);
or UO_265 (O_265,N_2990,N_2953);
nor UO_266 (O_266,N_2954,N_2958);
nand UO_267 (O_267,N_2982,N_2980);
and UO_268 (O_268,N_2958,N_2970);
xor UO_269 (O_269,N_2981,N_2994);
nand UO_270 (O_270,N_2973,N_2971);
and UO_271 (O_271,N_2983,N_2974);
nand UO_272 (O_272,N_2968,N_2992);
and UO_273 (O_273,N_2958,N_2973);
nor UO_274 (O_274,N_2977,N_2991);
or UO_275 (O_275,N_2963,N_2965);
nor UO_276 (O_276,N_2952,N_2974);
and UO_277 (O_277,N_2964,N_2956);
xor UO_278 (O_278,N_2953,N_2956);
and UO_279 (O_279,N_2972,N_2968);
or UO_280 (O_280,N_2994,N_2950);
or UO_281 (O_281,N_2958,N_2960);
xor UO_282 (O_282,N_2956,N_2951);
or UO_283 (O_283,N_2952,N_2970);
nor UO_284 (O_284,N_2999,N_2994);
nor UO_285 (O_285,N_2983,N_2957);
or UO_286 (O_286,N_2960,N_2966);
and UO_287 (O_287,N_2995,N_2955);
or UO_288 (O_288,N_2958,N_2986);
nor UO_289 (O_289,N_2969,N_2954);
nor UO_290 (O_290,N_2961,N_2989);
or UO_291 (O_291,N_2990,N_2992);
nor UO_292 (O_292,N_2998,N_2965);
and UO_293 (O_293,N_2991,N_2955);
nor UO_294 (O_294,N_2988,N_2997);
and UO_295 (O_295,N_2987,N_2956);
nor UO_296 (O_296,N_2987,N_2977);
nor UO_297 (O_297,N_2974,N_2979);
and UO_298 (O_298,N_2955,N_2985);
and UO_299 (O_299,N_2959,N_2957);
nor UO_300 (O_300,N_2954,N_2982);
and UO_301 (O_301,N_2964,N_2965);
nor UO_302 (O_302,N_2983,N_2998);
and UO_303 (O_303,N_2987,N_2961);
or UO_304 (O_304,N_2999,N_2971);
or UO_305 (O_305,N_2996,N_2968);
nand UO_306 (O_306,N_2958,N_2968);
nand UO_307 (O_307,N_2964,N_2955);
and UO_308 (O_308,N_2996,N_2953);
nand UO_309 (O_309,N_2971,N_2980);
nor UO_310 (O_310,N_2984,N_2967);
or UO_311 (O_311,N_2985,N_2963);
nor UO_312 (O_312,N_2958,N_2953);
or UO_313 (O_313,N_2955,N_2986);
and UO_314 (O_314,N_2992,N_2970);
nor UO_315 (O_315,N_2954,N_2986);
nor UO_316 (O_316,N_2978,N_2966);
nor UO_317 (O_317,N_2972,N_2995);
nor UO_318 (O_318,N_2956,N_2988);
and UO_319 (O_319,N_2964,N_2993);
and UO_320 (O_320,N_2957,N_2996);
or UO_321 (O_321,N_2995,N_2950);
and UO_322 (O_322,N_2977,N_2955);
nand UO_323 (O_323,N_2960,N_2975);
nand UO_324 (O_324,N_2964,N_2986);
nor UO_325 (O_325,N_2980,N_2990);
nor UO_326 (O_326,N_2960,N_2976);
nor UO_327 (O_327,N_2983,N_2973);
and UO_328 (O_328,N_2996,N_2952);
nor UO_329 (O_329,N_2958,N_2999);
or UO_330 (O_330,N_2994,N_2956);
or UO_331 (O_331,N_2985,N_2956);
and UO_332 (O_332,N_2969,N_2963);
nand UO_333 (O_333,N_2956,N_2973);
nand UO_334 (O_334,N_2979,N_2961);
nor UO_335 (O_335,N_2986,N_2950);
xor UO_336 (O_336,N_2980,N_2963);
and UO_337 (O_337,N_2975,N_2974);
and UO_338 (O_338,N_2994,N_2963);
nor UO_339 (O_339,N_2978,N_2986);
xor UO_340 (O_340,N_2965,N_2967);
xnor UO_341 (O_341,N_2955,N_2999);
nand UO_342 (O_342,N_2984,N_2993);
nor UO_343 (O_343,N_2980,N_2975);
nand UO_344 (O_344,N_2952,N_2960);
nor UO_345 (O_345,N_2978,N_2960);
xor UO_346 (O_346,N_2955,N_2963);
and UO_347 (O_347,N_2967,N_2986);
nand UO_348 (O_348,N_2963,N_2979);
nand UO_349 (O_349,N_2988,N_2953);
nor UO_350 (O_350,N_2996,N_2955);
nor UO_351 (O_351,N_2951,N_2968);
and UO_352 (O_352,N_2952,N_2992);
and UO_353 (O_353,N_2973,N_2991);
or UO_354 (O_354,N_2998,N_2988);
or UO_355 (O_355,N_2995,N_2973);
and UO_356 (O_356,N_2987,N_2962);
or UO_357 (O_357,N_2958,N_2951);
xor UO_358 (O_358,N_2970,N_2964);
nand UO_359 (O_359,N_2951,N_2970);
and UO_360 (O_360,N_2980,N_2988);
or UO_361 (O_361,N_2972,N_2966);
and UO_362 (O_362,N_2991,N_2956);
or UO_363 (O_363,N_2967,N_2999);
nor UO_364 (O_364,N_2985,N_2967);
and UO_365 (O_365,N_2954,N_2981);
or UO_366 (O_366,N_2990,N_2998);
nor UO_367 (O_367,N_2971,N_2978);
nand UO_368 (O_368,N_2963,N_2958);
and UO_369 (O_369,N_2985,N_2996);
nor UO_370 (O_370,N_2998,N_2951);
and UO_371 (O_371,N_2955,N_2956);
nand UO_372 (O_372,N_2990,N_2991);
nor UO_373 (O_373,N_2991,N_2982);
and UO_374 (O_374,N_2952,N_2972);
nor UO_375 (O_375,N_2954,N_2996);
nand UO_376 (O_376,N_2961,N_2950);
and UO_377 (O_377,N_2970,N_2979);
nand UO_378 (O_378,N_2962,N_2951);
and UO_379 (O_379,N_2958,N_2996);
and UO_380 (O_380,N_2970,N_2962);
nand UO_381 (O_381,N_2959,N_2993);
nor UO_382 (O_382,N_2996,N_2970);
or UO_383 (O_383,N_2996,N_2999);
or UO_384 (O_384,N_2960,N_2996);
nor UO_385 (O_385,N_2985,N_2950);
and UO_386 (O_386,N_2991,N_2984);
nor UO_387 (O_387,N_2955,N_2976);
nor UO_388 (O_388,N_2964,N_2969);
and UO_389 (O_389,N_2959,N_2994);
and UO_390 (O_390,N_2994,N_2980);
nor UO_391 (O_391,N_2953,N_2965);
nor UO_392 (O_392,N_2982,N_2985);
or UO_393 (O_393,N_2998,N_2994);
and UO_394 (O_394,N_2980,N_2970);
nand UO_395 (O_395,N_2997,N_2974);
nand UO_396 (O_396,N_2957,N_2990);
nor UO_397 (O_397,N_2999,N_2983);
or UO_398 (O_398,N_2963,N_2970);
nand UO_399 (O_399,N_2970,N_2965);
nand UO_400 (O_400,N_2957,N_2989);
nor UO_401 (O_401,N_2973,N_2986);
and UO_402 (O_402,N_2967,N_2972);
xnor UO_403 (O_403,N_2968,N_2991);
nand UO_404 (O_404,N_2998,N_2993);
nand UO_405 (O_405,N_2984,N_2959);
nand UO_406 (O_406,N_2964,N_2966);
nor UO_407 (O_407,N_2968,N_2986);
nand UO_408 (O_408,N_2956,N_2950);
and UO_409 (O_409,N_2977,N_2964);
and UO_410 (O_410,N_2967,N_2973);
and UO_411 (O_411,N_2988,N_2977);
or UO_412 (O_412,N_2978,N_2980);
and UO_413 (O_413,N_2994,N_2960);
and UO_414 (O_414,N_2980,N_2996);
nand UO_415 (O_415,N_2965,N_2983);
xor UO_416 (O_416,N_2971,N_2963);
nor UO_417 (O_417,N_2958,N_2957);
nand UO_418 (O_418,N_2999,N_2972);
nor UO_419 (O_419,N_2971,N_2952);
nor UO_420 (O_420,N_2996,N_2962);
and UO_421 (O_421,N_2990,N_2976);
xor UO_422 (O_422,N_2977,N_2993);
nand UO_423 (O_423,N_2982,N_2997);
nand UO_424 (O_424,N_2963,N_2982);
nand UO_425 (O_425,N_2992,N_2983);
nor UO_426 (O_426,N_2961,N_2974);
and UO_427 (O_427,N_2976,N_2989);
nor UO_428 (O_428,N_2959,N_2962);
and UO_429 (O_429,N_2969,N_2986);
nor UO_430 (O_430,N_2978,N_2954);
nand UO_431 (O_431,N_2961,N_2998);
and UO_432 (O_432,N_2979,N_2951);
or UO_433 (O_433,N_2978,N_2999);
nor UO_434 (O_434,N_2995,N_2989);
and UO_435 (O_435,N_2975,N_2981);
xnor UO_436 (O_436,N_2958,N_2972);
nor UO_437 (O_437,N_2976,N_2962);
and UO_438 (O_438,N_2952,N_2993);
or UO_439 (O_439,N_2985,N_2977);
nand UO_440 (O_440,N_2992,N_2981);
and UO_441 (O_441,N_2965,N_2978);
nand UO_442 (O_442,N_2970,N_2997);
nor UO_443 (O_443,N_2975,N_2999);
nor UO_444 (O_444,N_2960,N_2951);
xnor UO_445 (O_445,N_2992,N_2964);
or UO_446 (O_446,N_2969,N_2979);
and UO_447 (O_447,N_2971,N_2953);
or UO_448 (O_448,N_2958,N_2997);
and UO_449 (O_449,N_2953,N_2985);
nor UO_450 (O_450,N_2981,N_2972);
nor UO_451 (O_451,N_2987,N_2952);
and UO_452 (O_452,N_2988,N_2960);
nand UO_453 (O_453,N_2953,N_2968);
and UO_454 (O_454,N_2986,N_2974);
or UO_455 (O_455,N_2955,N_2979);
nand UO_456 (O_456,N_2983,N_2987);
nor UO_457 (O_457,N_2983,N_2979);
xor UO_458 (O_458,N_2989,N_2977);
nand UO_459 (O_459,N_2954,N_2994);
and UO_460 (O_460,N_2951,N_2980);
or UO_461 (O_461,N_2992,N_2986);
or UO_462 (O_462,N_2996,N_2988);
and UO_463 (O_463,N_2975,N_2994);
or UO_464 (O_464,N_2983,N_2982);
nor UO_465 (O_465,N_2997,N_2968);
nor UO_466 (O_466,N_2990,N_2973);
or UO_467 (O_467,N_2995,N_2967);
and UO_468 (O_468,N_2968,N_2967);
and UO_469 (O_469,N_2983,N_2989);
or UO_470 (O_470,N_2990,N_2960);
and UO_471 (O_471,N_2968,N_2966);
nor UO_472 (O_472,N_2990,N_2954);
nand UO_473 (O_473,N_2962,N_2963);
nor UO_474 (O_474,N_2987,N_2975);
and UO_475 (O_475,N_2976,N_2995);
nor UO_476 (O_476,N_2955,N_2950);
xnor UO_477 (O_477,N_2957,N_2980);
and UO_478 (O_478,N_2977,N_2950);
and UO_479 (O_479,N_2972,N_2983);
xor UO_480 (O_480,N_2999,N_2953);
xnor UO_481 (O_481,N_2997,N_2993);
and UO_482 (O_482,N_2973,N_2952);
and UO_483 (O_483,N_2976,N_2974);
and UO_484 (O_484,N_2971,N_2965);
nor UO_485 (O_485,N_2972,N_2965);
or UO_486 (O_486,N_2976,N_2987);
nand UO_487 (O_487,N_2953,N_2979);
and UO_488 (O_488,N_2997,N_2985);
nand UO_489 (O_489,N_2998,N_2960);
and UO_490 (O_490,N_2993,N_2953);
nor UO_491 (O_491,N_2950,N_2967);
or UO_492 (O_492,N_2982,N_2957);
nand UO_493 (O_493,N_2995,N_2964);
nand UO_494 (O_494,N_2985,N_2998);
nor UO_495 (O_495,N_2975,N_2997);
and UO_496 (O_496,N_2989,N_2990);
or UO_497 (O_497,N_2960,N_2967);
and UO_498 (O_498,N_2984,N_2988);
or UO_499 (O_499,N_2952,N_2982);
endmodule