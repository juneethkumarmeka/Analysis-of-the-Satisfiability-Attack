module basic_1000_10000_1500_10_levels_1xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
and U0 (N_0,In_418,In_835);
nand U1 (N_1,In_451,In_686);
or U2 (N_2,In_522,In_872);
and U3 (N_3,In_834,In_743);
or U4 (N_4,In_67,In_741);
and U5 (N_5,In_916,In_921);
and U6 (N_6,In_636,In_990);
and U7 (N_7,In_216,In_580);
or U8 (N_8,In_715,In_317);
nor U9 (N_9,In_876,In_670);
nand U10 (N_10,In_653,In_83);
nand U11 (N_11,In_77,In_744);
and U12 (N_12,In_80,In_548);
nor U13 (N_13,In_350,In_899);
or U14 (N_14,In_693,In_874);
nor U15 (N_15,In_824,In_544);
nor U16 (N_16,In_22,In_807);
nor U17 (N_17,In_752,In_10);
nand U18 (N_18,In_160,In_838);
and U19 (N_19,In_507,In_945);
or U20 (N_20,In_383,In_880);
or U21 (N_21,In_764,In_576);
and U22 (N_22,In_806,In_247);
nand U23 (N_23,In_612,In_738);
and U24 (N_24,In_542,In_812);
nor U25 (N_25,In_659,In_347);
nor U26 (N_26,In_272,In_658);
and U27 (N_27,In_655,In_570);
or U28 (N_28,In_914,In_155);
nor U29 (N_29,In_192,In_525);
and U30 (N_30,In_619,In_957);
nor U31 (N_31,In_447,In_203);
or U32 (N_32,In_815,In_931);
nand U33 (N_33,In_200,In_57);
nor U34 (N_34,In_257,In_113);
nor U35 (N_35,In_21,In_991);
and U36 (N_36,In_376,In_147);
and U37 (N_37,In_918,In_905);
or U38 (N_38,In_29,In_49);
and U39 (N_39,In_831,In_816);
or U40 (N_40,In_749,In_438);
and U41 (N_41,In_270,In_152);
nor U42 (N_42,In_818,In_59);
nand U43 (N_43,In_159,In_291);
nand U44 (N_44,In_162,In_556);
nand U45 (N_45,In_61,In_87);
nor U46 (N_46,In_201,In_372);
nand U47 (N_47,In_966,In_657);
and U48 (N_48,In_250,In_589);
or U49 (N_49,In_88,In_627);
nand U50 (N_50,In_742,In_712);
and U51 (N_51,In_615,In_193);
and U52 (N_52,In_364,In_236);
and U53 (N_53,In_706,In_645);
and U54 (N_54,In_930,In_707);
nor U55 (N_55,In_395,In_249);
nand U56 (N_56,In_341,In_198);
or U57 (N_57,In_898,In_52);
nor U58 (N_58,In_313,In_359);
or U59 (N_59,In_756,In_348);
nand U60 (N_60,In_660,In_3);
and U61 (N_61,In_593,In_256);
nor U62 (N_62,In_828,In_760);
nor U63 (N_63,In_410,In_448);
nand U64 (N_64,In_354,In_284);
or U65 (N_65,In_19,In_261);
or U66 (N_66,In_53,In_186);
nor U67 (N_67,In_702,In_301);
nand U68 (N_68,In_850,In_811);
nand U69 (N_69,In_477,In_911);
nand U70 (N_70,In_783,In_639);
nor U71 (N_71,In_392,In_778);
nor U72 (N_72,In_573,In_298);
nor U73 (N_73,In_732,In_475);
nand U74 (N_74,In_25,In_163);
and U75 (N_75,In_353,In_727);
nor U76 (N_76,In_759,In_146);
nand U77 (N_77,In_822,In_206);
nor U78 (N_78,In_43,In_987);
nand U79 (N_79,In_191,In_240);
nor U80 (N_80,In_863,In_690);
and U81 (N_81,In_889,In_757);
nor U82 (N_82,In_797,In_151);
nand U83 (N_83,In_409,In_369);
nor U84 (N_84,In_505,In_932);
nand U85 (N_85,In_394,In_70);
nor U86 (N_86,In_330,In_798);
nor U87 (N_87,In_583,In_865);
and U88 (N_88,In_747,In_517);
and U89 (N_89,In_569,In_729);
or U90 (N_90,In_169,In_998);
nor U91 (N_91,In_404,In_72);
nand U92 (N_92,In_745,In_319);
or U93 (N_93,In_515,In_417);
and U94 (N_94,In_672,In_93);
nor U95 (N_95,In_852,In_119);
and U96 (N_96,In_318,In_253);
nand U97 (N_97,In_652,In_793);
nor U98 (N_98,In_399,In_164);
and U99 (N_99,In_337,In_551);
or U100 (N_100,In_733,In_597);
nand U101 (N_101,In_927,In_893);
or U102 (N_102,In_156,In_509);
or U103 (N_103,In_195,In_944);
or U104 (N_104,In_260,In_278);
nor U105 (N_105,In_427,In_943);
nand U106 (N_106,In_158,In_843);
and U107 (N_107,In_76,In_56);
and U108 (N_108,In_237,In_763);
nor U109 (N_109,In_973,In_150);
and U110 (N_110,In_922,In_882);
nand U111 (N_111,In_609,In_772);
or U112 (N_112,In_558,In_141);
nand U113 (N_113,In_582,In_904);
nor U114 (N_114,In_224,In_205);
nor U115 (N_115,In_599,In_626);
nor U116 (N_116,In_232,In_997);
or U117 (N_117,In_685,In_820);
and U118 (N_118,In_452,In_327);
nand U119 (N_119,In_381,In_188);
and U120 (N_120,In_873,In_50);
or U121 (N_121,In_17,In_833);
or U122 (N_122,In_423,In_243);
nor U123 (N_123,In_94,In_817);
nor U124 (N_124,In_518,In_962);
or U125 (N_125,In_445,In_455);
nor U126 (N_126,In_12,In_913);
or U127 (N_127,In_197,In_830);
and U128 (N_128,In_993,In_912);
nand U129 (N_129,In_390,In_387);
and U130 (N_130,In_716,In_721);
nor U131 (N_131,In_40,In_634);
or U132 (N_132,In_459,In_994);
and U133 (N_133,In_934,In_799);
nor U134 (N_134,In_688,In_613);
and U135 (N_135,In_602,In_262);
and U136 (N_136,In_808,In_836);
and U137 (N_137,In_400,In_435);
or U138 (N_138,In_366,In_233);
nand U139 (N_139,In_111,In_391);
nor U140 (N_140,In_123,In_258);
and U141 (N_141,In_462,In_101);
or U142 (N_142,In_540,In_183);
or U143 (N_143,In_403,In_221);
nor U144 (N_144,In_283,In_65);
nand U145 (N_145,In_287,In_888);
nand U146 (N_146,In_125,In_575);
or U147 (N_147,In_981,In_802);
xor U148 (N_148,In_86,In_765);
and U149 (N_149,In_884,In_434);
and U150 (N_150,In_559,In_109);
or U151 (N_151,In_175,In_726);
or U152 (N_152,In_595,In_571);
and U153 (N_153,In_784,In_97);
or U154 (N_154,In_762,In_211);
or U155 (N_155,In_254,In_924);
nand U156 (N_156,In_338,In_398);
and U157 (N_157,In_11,In_648);
or U158 (N_158,In_116,In_803);
or U159 (N_159,In_442,In_414);
nand U160 (N_160,In_121,In_430);
or U161 (N_161,In_720,In_185);
and U162 (N_162,In_750,In_857);
and U163 (N_163,In_9,In_251);
or U164 (N_164,In_794,In_596);
and U165 (N_165,In_333,In_98);
or U166 (N_166,In_496,In_32);
nor U167 (N_167,In_265,In_826);
and U168 (N_168,In_207,In_578);
and U169 (N_169,In_241,In_413);
or U170 (N_170,In_345,In_290);
nand U171 (N_171,In_497,In_5);
and U172 (N_172,In_604,In_180);
and U173 (N_173,In_854,In_555);
nor U174 (N_174,In_524,In_878);
nor U175 (N_175,In_105,In_877);
nand U176 (N_176,In_506,In_138);
nor U177 (N_177,In_126,In_845);
or U178 (N_178,In_388,In_1);
or U179 (N_179,In_714,In_965);
nor U180 (N_180,In_946,In_47);
nor U181 (N_181,In_502,In_329);
nor U182 (N_182,In_220,In_304);
or U183 (N_183,In_697,In_63);
nor U184 (N_184,In_28,In_855);
nand U185 (N_185,In_621,In_286);
nor U186 (N_186,In_84,In_89);
and U187 (N_187,In_687,In_380);
or U188 (N_188,In_182,In_416);
nor U189 (N_189,In_199,In_374);
nand U190 (N_190,In_315,In_587);
and U191 (N_191,In_988,In_933);
and U192 (N_192,In_124,In_15);
or U193 (N_193,In_723,In_620);
or U194 (N_194,In_62,In_553);
nor U195 (N_195,In_300,In_791);
nor U196 (N_196,In_407,In_891);
nand U197 (N_197,In_173,In_919);
nor U198 (N_198,In_344,In_950);
or U199 (N_199,In_696,In_935);
or U200 (N_200,In_214,In_16);
nand U201 (N_201,In_635,In_566);
nor U202 (N_202,In_297,In_346);
and U203 (N_203,In_947,In_681);
or U204 (N_204,In_379,In_157);
or U205 (N_205,In_190,In_534);
or U206 (N_206,In_903,In_755);
nor U207 (N_207,In_643,In_585);
nand U208 (N_208,In_564,In_234);
nor U209 (N_209,In_736,In_669);
or U210 (N_210,In_777,In_143);
nor U211 (N_211,In_27,In_36);
or U212 (N_212,In_859,In_335);
nand U213 (N_213,In_875,In_871);
or U214 (N_214,In_360,In_795);
and U215 (N_215,In_885,In_801);
nand U216 (N_216,In_456,In_66);
or U217 (N_217,In_511,In_623);
nand U218 (N_218,In_149,In_724);
or U219 (N_219,In_73,In_557);
nand U220 (N_220,In_483,In_238);
nand U221 (N_221,In_968,In_554);
nor U222 (N_222,In_91,In_252);
nor U223 (N_223,In_481,In_881);
nand U224 (N_224,In_979,In_95);
and U225 (N_225,In_656,In_689);
and U226 (N_226,In_271,In_948);
nor U227 (N_227,In_68,In_242);
and U228 (N_228,In_420,In_897);
or U229 (N_229,In_739,In_731);
nand U230 (N_230,In_805,In_393);
and U231 (N_231,In_960,In_117);
and U232 (N_232,In_279,In_673);
and U233 (N_233,In_227,In_770);
or U234 (N_234,In_974,In_684);
nand U235 (N_235,In_970,In_30);
nor U236 (N_236,In_100,In_142);
xor U237 (N_237,In_137,In_969);
and U238 (N_238,In_560,In_225);
nand U239 (N_239,In_282,In_473);
and U240 (N_240,In_492,In_925);
or U241 (N_241,In_649,In_299);
nand U242 (N_242,In_625,In_135);
nand U243 (N_243,In_526,In_840);
or U244 (N_244,In_331,In_375);
and U245 (N_245,In_78,In_489);
nor U246 (N_246,In_980,In_144);
nor U247 (N_247,In_644,In_737);
nor U248 (N_248,In_154,In_491);
nor U249 (N_249,In_268,In_848);
nor U250 (N_250,In_132,In_470);
and U251 (N_251,In_118,In_230);
or U252 (N_252,In_907,In_972);
and U253 (N_253,In_773,In_426);
nor U254 (N_254,In_229,In_767);
or U255 (N_255,In_939,In_187);
nand U256 (N_256,In_532,In_222);
and U257 (N_257,In_54,In_787);
nand U258 (N_258,In_292,In_2);
or U259 (N_259,In_691,In_546);
and U260 (N_260,In_860,In_82);
nor U261 (N_261,In_901,In_754);
and U262 (N_262,In_894,In_485);
xor U263 (N_263,In_614,In_136);
xor U264 (N_264,In_281,In_129);
and U265 (N_265,In_479,In_472);
or U266 (N_266,In_929,In_717);
nor U267 (N_267,In_349,In_996);
and U268 (N_268,In_428,In_539);
or U269 (N_269,In_501,In_902);
nand U270 (N_270,In_630,In_39);
nor U271 (N_271,In_883,In_314);
nor U272 (N_272,In_577,In_246);
nor U273 (N_273,In_202,In_326);
and U274 (N_274,In_718,In_231);
nand U275 (N_275,In_196,In_273);
or U276 (N_276,In_303,In_305);
and U277 (N_277,In_320,In_786);
nor U278 (N_278,In_208,In_145);
and U279 (N_279,In_469,In_362);
and U280 (N_280,In_184,In_565);
or U281 (N_281,In_458,In_266);
nand U282 (N_282,In_923,In_306);
nor U283 (N_283,In_992,In_495);
nor U284 (N_284,In_44,In_468);
or U285 (N_285,In_425,In_926);
and U286 (N_286,In_140,In_971);
and U287 (N_287,In_464,In_975);
or U288 (N_288,In_959,In_35);
nor U289 (N_289,In_41,In_120);
or U290 (N_290,In_941,In_955);
or U291 (N_291,In_704,In_789);
nor U292 (N_292,In_790,In_309);
or U293 (N_293,In_521,In_267);
nor U294 (N_294,In_680,In_461);
and U295 (N_295,In_890,In_734);
nand U296 (N_296,In_699,In_983);
nand U297 (N_297,In_856,In_255);
nor U298 (N_298,In_999,In_868);
nand U299 (N_299,In_513,In_611);
nand U300 (N_300,In_520,In_170);
nor U301 (N_301,In_710,In_771);
nand U302 (N_302,In_694,In_788);
and U303 (N_303,In_600,In_568);
or U304 (N_304,In_844,In_753);
nor U305 (N_305,In_322,In_210);
nor U306 (N_306,In_79,In_370);
or U307 (N_307,In_377,In_864);
or U308 (N_308,In_722,In_168);
nand U309 (N_309,In_510,In_134);
nor U310 (N_310,In_295,In_24);
or U311 (N_311,In_851,In_829);
nor U312 (N_312,In_839,In_821);
or U313 (N_313,In_776,In_519);
nor U314 (N_314,In_512,In_406);
or U315 (N_315,In_746,In_244);
nor U316 (N_316,In_4,In_682);
nor U317 (N_317,In_13,In_535);
or U318 (N_318,In_751,In_478);
and U319 (N_319,In_429,In_343);
and U320 (N_320,In_340,In_617);
and U321 (N_321,In_668,In_415);
nor U322 (N_322,In_867,In_591);
nor U323 (N_323,In_740,In_665);
nor U324 (N_324,In_779,In_176);
nand U325 (N_325,In_480,In_536);
and U326 (N_326,In_274,In_529);
or U327 (N_327,In_910,In_647);
or U328 (N_328,In_954,In_385);
or U329 (N_329,In_289,In_949);
or U330 (N_330,In_581,In_976);
nor U331 (N_331,In_610,In_424);
xor U332 (N_332,In_701,In_165);
nand U333 (N_333,In_769,In_758);
or U334 (N_334,In_870,In_74);
or U335 (N_335,In_310,In_549);
xnor U336 (N_336,In_679,In_695);
nor U337 (N_337,In_0,In_115);
nor U338 (N_338,In_92,In_832);
nand U339 (N_339,In_90,In_561);
nor U340 (N_340,In_55,In_408);
and U341 (N_341,In_453,In_709);
nor U342 (N_342,In_705,In_547);
and U343 (N_343,In_352,In_23);
and U344 (N_344,In_153,In_766);
and U345 (N_345,In_841,In_642);
or U346 (N_346,In_523,In_213);
nor U347 (N_347,In_45,In_819);
nor U348 (N_348,In_58,In_606);
nor U349 (N_349,In_953,In_543);
and U350 (N_350,In_661,In_356);
or U351 (N_351,In_530,In_444);
nand U352 (N_352,In_174,In_248);
nor U353 (N_353,In_46,In_671);
nor U354 (N_354,In_6,In_900);
nor U355 (N_355,In_936,In_486);
or U356 (N_356,In_703,In_476);
and U357 (N_357,In_804,In_952);
nor U358 (N_358,In_294,In_674);
nand U359 (N_359,In_892,In_528);
and U360 (N_360,In_449,In_629);
nand U361 (N_361,In_412,In_713);
and U362 (N_362,In_504,In_107);
nor U363 (N_363,In_325,In_683);
nand U364 (N_364,In_110,In_454);
nor U365 (N_365,In_809,In_396);
xnor U366 (N_366,In_984,In_735);
or U367 (N_367,In_373,In_574);
nor U368 (N_368,In_796,In_48);
nand U369 (N_369,In_217,In_651);
or U370 (N_370,In_748,In_482);
nand U371 (N_371,In_460,In_989);
nor U372 (N_372,In_640,In_781);
and U373 (N_373,In_280,In_917);
nor U374 (N_374,In_128,In_616);
nor U375 (N_375,In_296,In_60);
and U376 (N_376,In_339,In_441);
or U377 (N_377,In_603,In_127);
nand U378 (N_378,In_887,In_321);
and U379 (N_379,In_328,In_956);
xor U380 (N_380,In_958,In_368);
or U381 (N_381,In_537,In_386);
nor U382 (N_382,In_940,In_26);
nor U383 (N_383,In_586,In_365);
nand U384 (N_384,In_814,In_148);
or U385 (N_385,In_235,In_293);
nand U386 (N_386,In_323,In_664);
nor U387 (N_387,In_432,In_792);
nand U388 (N_388,In_466,In_405);
or U389 (N_389,In_218,In_527);
nor U390 (N_390,In_308,In_928);
nor U391 (N_391,In_633,In_130);
or U392 (N_392,In_361,In_411);
and U393 (N_393,In_915,In_336);
or U394 (N_394,In_895,In_516);
nand U395 (N_395,In_862,In_288);
nor U396 (N_396,In_334,In_499);
and U397 (N_397,In_239,In_436);
nand U398 (N_398,In_20,In_909);
nand U399 (N_399,In_312,In_302);
nand U400 (N_400,In_269,In_842);
and U401 (N_401,In_768,In_650);
nand U402 (N_402,In_598,In_692);
or U403 (N_403,In_285,In_719);
nor U404 (N_404,In_624,In_133);
nand U405 (N_405,In_131,In_75);
or U406 (N_406,In_849,In_245);
nor U407 (N_407,In_584,In_450);
nor U408 (N_408,In_780,In_641);
nand U409 (N_409,In_178,In_774);
nor U410 (N_410,In_708,In_172);
nand U411 (N_411,In_550,In_14);
nand U412 (N_412,In_775,In_977);
nor U413 (N_413,In_995,In_963);
nand U414 (N_414,In_228,In_324);
and U415 (N_415,In_263,In_908);
and U416 (N_416,In_401,In_311);
or U417 (N_417,In_31,In_985);
and U418 (N_418,In_358,In_18);
and U419 (N_419,In_171,In_700);
or U420 (N_420,In_810,In_646);
nand U421 (N_421,In_99,In_419);
nand U422 (N_422,In_33,In_440);
or U423 (N_423,In_106,In_71);
nand U424 (N_424,In_938,In_638);
nor U425 (N_425,In_601,In_605);
and U426 (N_426,In_662,In_823);
nand U427 (N_427,In_7,In_886);
nand U428 (N_428,In_181,In_982);
nor U429 (N_429,In_104,In_667);
and U430 (N_430,In_42,In_920);
or U431 (N_431,In_122,In_446);
and U432 (N_432,In_457,In_34);
nand U433 (N_433,In_533,In_675);
or U434 (N_434,In_866,In_64);
nor U435 (N_435,In_223,In_471);
and U436 (N_436,In_467,In_166);
and U437 (N_437,In_572,In_531);
or U438 (N_438,In_677,In_179);
nor U439 (N_439,In_474,In_853);
nor U440 (N_440,In_632,In_563);
nor U441 (N_441,In_378,In_503);
nand U442 (N_442,In_189,In_397);
nor U443 (N_443,In_355,In_725);
nor U444 (N_444,In_307,In_332);
nor U445 (N_445,In_161,In_978);
nor U446 (N_446,In_514,In_847);
nor U447 (N_447,In_389,In_858);
or U448 (N_448,In_590,In_541);
or U449 (N_449,In_942,In_618);
nor U450 (N_450,In_562,In_215);
nand U451 (N_451,In_631,In_508);
nor U452 (N_452,In_967,In_421);
and U453 (N_453,In_484,In_363);
and U454 (N_454,In_567,In_488);
nor U455 (N_455,In_552,In_102);
nand U456 (N_456,In_204,In_607);
and U457 (N_457,In_342,In_951);
nor U458 (N_458,In_194,In_357);
nor U459 (N_459,In_433,In_114);
nand U460 (N_460,In_490,In_402);
and U461 (N_461,In_437,In_259);
or U462 (N_462,In_487,In_38);
nand U463 (N_463,In_608,In_209);
nand U464 (N_464,In_711,In_761);
nand U465 (N_465,In_69,In_678);
nor U466 (N_466,In_827,In_837);
and U467 (N_467,In_937,In_139);
nand U468 (N_468,In_316,In_896);
nand U469 (N_469,In_879,In_277);
nor U470 (N_470,In_219,In_371);
nor U471 (N_471,In_51,In_986);
or U472 (N_472,In_112,In_500);
nand U473 (N_473,In_785,In_698);
nand U474 (N_474,In_498,In_869);
nand U475 (N_475,In_81,In_961);
nand U476 (N_476,In_579,In_177);
and U477 (N_477,In_666,In_422);
and U478 (N_478,In_663,In_494);
and U479 (N_479,In_37,In_906);
nand U480 (N_480,In_813,In_730);
nor U481 (N_481,In_964,In_276);
nand U482 (N_482,In_545,In_212);
and U483 (N_483,In_676,In_588);
or U484 (N_484,In_443,In_439);
nand U485 (N_485,In_103,In_8);
and U486 (N_486,In_465,In_728);
and U487 (N_487,In_861,In_846);
nor U488 (N_488,In_538,In_654);
nand U489 (N_489,In_628,In_167);
and U490 (N_490,In_367,In_351);
nand U491 (N_491,In_85,In_594);
nand U492 (N_492,In_275,In_622);
xor U493 (N_493,In_782,In_382);
and U494 (N_494,In_800,In_592);
or U495 (N_495,In_108,In_431);
nor U496 (N_496,In_384,In_493);
or U497 (N_497,In_637,In_96);
or U498 (N_498,In_264,In_463);
nand U499 (N_499,In_226,In_825);
nand U500 (N_500,In_449,In_748);
and U501 (N_501,In_441,In_405);
nor U502 (N_502,In_518,In_283);
or U503 (N_503,In_229,In_805);
and U504 (N_504,In_198,In_650);
or U505 (N_505,In_866,In_644);
nor U506 (N_506,In_999,In_956);
nor U507 (N_507,In_72,In_631);
nor U508 (N_508,In_265,In_737);
xor U509 (N_509,In_898,In_328);
or U510 (N_510,In_361,In_343);
nand U511 (N_511,In_617,In_205);
nor U512 (N_512,In_197,In_711);
nor U513 (N_513,In_802,In_347);
or U514 (N_514,In_769,In_910);
nor U515 (N_515,In_796,In_790);
or U516 (N_516,In_984,In_980);
or U517 (N_517,In_161,In_194);
nand U518 (N_518,In_460,In_681);
and U519 (N_519,In_827,In_814);
nor U520 (N_520,In_376,In_778);
nand U521 (N_521,In_381,In_179);
and U522 (N_522,In_375,In_312);
or U523 (N_523,In_152,In_258);
or U524 (N_524,In_392,In_671);
or U525 (N_525,In_388,In_944);
nand U526 (N_526,In_606,In_1);
nor U527 (N_527,In_664,In_401);
and U528 (N_528,In_342,In_556);
xnor U529 (N_529,In_751,In_368);
nor U530 (N_530,In_590,In_115);
nor U531 (N_531,In_940,In_830);
nand U532 (N_532,In_427,In_354);
and U533 (N_533,In_601,In_315);
nand U534 (N_534,In_274,In_810);
nor U535 (N_535,In_124,In_693);
nand U536 (N_536,In_134,In_128);
and U537 (N_537,In_179,In_333);
and U538 (N_538,In_523,In_775);
nand U539 (N_539,In_245,In_839);
nand U540 (N_540,In_468,In_948);
nand U541 (N_541,In_751,In_703);
nand U542 (N_542,In_317,In_983);
or U543 (N_543,In_588,In_671);
nand U544 (N_544,In_43,In_718);
or U545 (N_545,In_522,In_545);
xnor U546 (N_546,In_631,In_520);
nor U547 (N_547,In_894,In_163);
and U548 (N_548,In_46,In_932);
or U549 (N_549,In_58,In_532);
and U550 (N_550,In_476,In_686);
nor U551 (N_551,In_283,In_861);
nand U552 (N_552,In_994,In_968);
and U553 (N_553,In_295,In_789);
nand U554 (N_554,In_54,In_669);
or U555 (N_555,In_766,In_723);
and U556 (N_556,In_446,In_889);
and U557 (N_557,In_945,In_367);
nor U558 (N_558,In_1,In_474);
and U559 (N_559,In_621,In_136);
nor U560 (N_560,In_72,In_597);
and U561 (N_561,In_77,In_411);
and U562 (N_562,In_600,In_314);
nor U563 (N_563,In_625,In_951);
nor U564 (N_564,In_185,In_735);
and U565 (N_565,In_149,In_254);
or U566 (N_566,In_276,In_553);
or U567 (N_567,In_521,In_325);
and U568 (N_568,In_174,In_189);
or U569 (N_569,In_672,In_600);
nand U570 (N_570,In_217,In_880);
or U571 (N_571,In_989,In_288);
and U572 (N_572,In_841,In_857);
or U573 (N_573,In_238,In_32);
nand U574 (N_574,In_50,In_611);
nand U575 (N_575,In_502,In_334);
nor U576 (N_576,In_41,In_297);
nor U577 (N_577,In_688,In_293);
nand U578 (N_578,In_437,In_757);
nand U579 (N_579,In_870,In_540);
nor U580 (N_580,In_192,In_923);
nand U581 (N_581,In_97,In_184);
and U582 (N_582,In_992,In_820);
or U583 (N_583,In_5,In_258);
or U584 (N_584,In_971,In_865);
or U585 (N_585,In_672,In_956);
nor U586 (N_586,In_845,In_283);
nor U587 (N_587,In_320,In_485);
nor U588 (N_588,In_348,In_198);
nor U589 (N_589,In_904,In_471);
and U590 (N_590,In_757,In_588);
and U591 (N_591,In_231,In_535);
nor U592 (N_592,In_267,In_180);
nor U593 (N_593,In_586,In_219);
nor U594 (N_594,In_407,In_231);
and U595 (N_595,In_504,In_945);
nor U596 (N_596,In_757,In_688);
nand U597 (N_597,In_34,In_421);
nor U598 (N_598,In_776,In_288);
nand U599 (N_599,In_635,In_701);
nor U600 (N_600,In_337,In_352);
nor U601 (N_601,In_698,In_297);
nor U602 (N_602,In_640,In_44);
nand U603 (N_603,In_611,In_371);
and U604 (N_604,In_952,In_665);
nand U605 (N_605,In_28,In_20);
nor U606 (N_606,In_753,In_785);
and U607 (N_607,In_382,In_685);
and U608 (N_608,In_191,In_457);
and U609 (N_609,In_225,In_816);
nand U610 (N_610,In_875,In_332);
nor U611 (N_611,In_450,In_199);
and U612 (N_612,In_372,In_929);
and U613 (N_613,In_850,In_652);
nand U614 (N_614,In_640,In_928);
or U615 (N_615,In_253,In_910);
or U616 (N_616,In_750,In_218);
nand U617 (N_617,In_806,In_678);
or U618 (N_618,In_670,In_555);
and U619 (N_619,In_999,In_818);
and U620 (N_620,In_394,In_321);
or U621 (N_621,In_714,In_499);
nor U622 (N_622,In_314,In_553);
and U623 (N_623,In_629,In_886);
and U624 (N_624,In_590,In_803);
nand U625 (N_625,In_668,In_957);
and U626 (N_626,In_932,In_854);
and U627 (N_627,In_258,In_216);
or U628 (N_628,In_132,In_978);
or U629 (N_629,In_949,In_576);
or U630 (N_630,In_738,In_93);
or U631 (N_631,In_112,In_856);
or U632 (N_632,In_866,In_144);
nor U633 (N_633,In_168,In_884);
nand U634 (N_634,In_283,In_766);
and U635 (N_635,In_401,In_457);
nor U636 (N_636,In_827,In_611);
nand U637 (N_637,In_123,In_153);
or U638 (N_638,In_455,In_309);
or U639 (N_639,In_334,In_133);
nor U640 (N_640,In_556,In_79);
nand U641 (N_641,In_569,In_715);
or U642 (N_642,In_460,In_107);
or U643 (N_643,In_877,In_933);
nand U644 (N_644,In_397,In_457);
nor U645 (N_645,In_510,In_77);
and U646 (N_646,In_424,In_162);
or U647 (N_647,In_821,In_208);
or U648 (N_648,In_176,In_496);
or U649 (N_649,In_210,In_178);
or U650 (N_650,In_77,In_694);
or U651 (N_651,In_72,In_330);
nand U652 (N_652,In_311,In_660);
nand U653 (N_653,In_354,In_4);
or U654 (N_654,In_137,In_796);
nand U655 (N_655,In_982,In_55);
or U656 (N_656,In_561,In_963);
nor U657 (N_657,In_324,In_615);
and U658 (N_658,In_514,In_187);
nand U659 (N_659,In_694,In_207);
and U660 (N_660,In_173,In_145);
nor U661 (N_661,In_282,In_310);
or U662 (N_662,In_596,In_480);
or U663 (N_663,In_531,In_160);
or U664 (N_664,In_450,In_90);
nor U665 (N_665,In_319,In_338);
nand U666 (N_666,In_104,In_698);
nor U667 (N_667,In_437,In_60);
nor U668 (N_668,In_751,In_385);
nand U669 (N_669,In_431,In_660);
and U670 (N_670,In_164,In_185);
nor U671 (N_671,In_276,In_15);
or U672 (N_672,In_958,In_859);
nor U673 (N_673,In_548,In_539);
nor U674 (N_674,In_48,In_834);
nor U675 (N_675,In_619,In_860);
nand U676 (N_676,In_140,In_1);
xor U677 (N_677,In_800,In_382);
or U678 (N_678,In_786,In_78);
nor U679 (N_679,In_465,In_837);
nand U680 (N_680,In_809,In_460);
nor U681 (N_681,In_760,In_326);
or U682 (N_682,In_368,In_548);
or U683 (N_683,In_512,In_888);
and U684 (N_684,In_303,In_668);
nand U685 (N_685,In_339,In_55);
and U686 (N_686,In_976,In_42);
nor U687 (N_687,In_115,In_964);
nand U688 (N_688,In_168,In_58);
nor U689 (N_689,In_432,In_646);
and U690 (N_690,In_365,In_65);
nand U691 (N_691,In_167,In_671);
nor U692 (N_692,In_444,In_702);
or U693 (N_693,In_487,In_766);
and U694 (N_694,In_492,In_971);
and U695 (N_695,In_124,In_248);
nand U696 (N_696,In_486,In_673);
nand U697 (N_697,In_230,In_349);
nor U698 (N_698,In_487,In_158);
nor U699 (N_699,In_735,In_871);
nor U700 (N_700,In_821,In_462);
nor U701 (N_701,In_502,In_973);
or U702 (N_702,In_997,In_889);
and U703 (N_703,In_841,In_868);
nor U704 (N_704,In_978,In_135);
or U705 (N_705,In_5,In_276);
and U706 (N_706,In_421,In_694);
or U707 (N_707,In_767,In_804);
nor U708 (N_708,In_737,In_991);
nor U709 (N_709,In_406,In_931);
nand U710 (N_710,In_245,In_784);
and U711 (N_711,In_327,In_39);
and U712 (N_712,In_812,In_343);
nand U713 (N_713,In_336,In_561);
or U714 (N_714,In_900,In_26);
nor U715 (N_715,In_313,In_106);
and U716 (N_716,In_155,In_922);
nor U717 (N_717,In_512,In_536);
xor U718 (N_718,In_524,In_498);
nand U719 (N_719,In_510,In_370);
nor U720 (N_720,In_901,In_415);
or U721 (N_721,In_587,In_920);
nor U722 (N_722,In_970,In_949);
nand U723 (N_723,In_581,In_564);
or U724 (N_724,In_847,In_658);
nand U725 (N_725,In_197,In_401);
and U726 (N_726,In_560,In_74);
nor U727 (N_727,In_65,In_520);
nand U728 (N_728,In_444,In_611);
nand U729 (N_729,In_108,In_738);
nor U730 (N_730,In_201,In_706);
nor U731 (N_731,In_82,In_426);
or U732 (N_732,In_769,In_536);
or U733 (N_733,In_269,In_724);
and U734 (N_734,In_909,In_799);
or U735 (N_735,In_451,In_660);
and U736 (N_736,In_811,In_295);
or U737 (N_737,In_553,In_246);
and U738 (N_738,In_159,In_26);
and U739 (N_739,In_128,In_611);
or U740 (N_740,In_310,In_498);
or U741 (N_741,In_291,In_452);
and U742 (N_742,In_145,In_62);
nand U743 (N_743,In_513,In_562);
and U744 (N_744,In_199,In_879);
or U745 (N_745,In_156,In_967);
nand U746 (N_746,In_887,In_186);
or U747 (N_747,In_533,In_577);
nor U748 (N_748,In_185,In_519);
or U749 (N_749,In_541,In_824);
or U750 (N_750,In_559,In_596);
or U751 (N_751,In_215,In_428);
nor U752 (N_752,In_761,In_399);
and U753 (N_753,In_532,In_986);
and U754 (N_754,In_650,In_391);
nand U755 (N_755,In_390,In_683);
nand U756 (N_756,In_219,In_370);
or U757 (N_757,In_878,In_901);
or U758 (N_758,In_69,In_271);
xor U759 (N_759,In_397,In_919);
and U760 (N_760,In_849,In_808);
xnor U761 (N_761,In_787,In_567);
nor U762 (N_762,In_206,In_119);
nand U763 (N_763,In_649,In_432);
or U764 (N_764,In_115,In_771);
nand U765 (N_765,In_617,In_745);
nand U766 (N_766,In_698,In_705);
or U767 (N_767,In_352,In_635);
nand U768 (N_768,In_224,In_913);
or U769 (N_769,In_820,In_295);
nand U770 (N_770,In_219,In_246);
or U771 (N_771,In_385,In_583);
nor U772 (N_772,In_87,In_380);
or U773 (N_773,In_927,In_512);
or U774 (N_774,In_954,In_766);
nor U775 (N_775,In_670,In_100);
and U776 (N_776,In_433,In_432);
nor U777 (N_777,In_641,In_501);
nand U778 (N_778,In_513,In_352);
nand U779 (N_779,In_97,In_832);
nand U780 (N_780,In_610,In_348);
nand U781 (N_781,In_927,In_354);
or U782 (N_782,In_191,In_433);
nor U783 (N_783,In_781,In_881);
and U784 (N_784,In_587,In_925);
or U785 (N_785,In_567,In_384);
and U786 (N_786,In_352,In_77);
nand U787 (N_787,In_692,In_805);
nand U788 (N_788,In_566,In_211);
and U789 (N_789,In_377,In_659);
or U790 (N_790,In_372,In_56);
and U791 (N_791,In_907,In_718);
nand U792 (N_792,In_981,In_625);
and U793 (N_793,In_527,In_894);
nor U794 (N_794,In_4,In_614);
nand U795 (N_795,In_914,In_395);
nor U796 (N_796,In_802,In_764);
nand U797 (N_797,In_537,In_346);
or U798 (N_798,In_60,In_595);
or U799 (N_799,In_255,In_35);
and U800 (N_800,In_654,In_444);
nand U801 (N_801,In_545,In_586);
and U802 (N_802,In_769,In_367);
and U803 (N_803,In_210,In_32);
and U804 (N_804,In_591,In_464);
and U805 (N_805,In_833,In_459);
and U806 (N_806,In_244,In_962);
nand U807 (N_807,In_843,In_556);
nand U808 (N_808,In_258,In_742);
nand U809 (N_809,In_923,In_619);
and U810 (N_810,In_324,In_60);
nor U811 (N_811,In_144,In_428);
nor U812 (N_812,In_179,In_669);
or U813 (N_813,In_742,In_300);
and U814 (N_814,In_126,In_99);
nor U815 (N_815,In_937,In_964);
nand U816 (N_816,In_351,In_240);
nor U817 (N_817,In_132,In_767);
and U818 (N_818,In_386,In_556);
nand U819 (N_819,In_673,In_235);
and U820 (N_820,In_827,In_445);
and U821 (N_821,In_968,In_955);
or U822 (N_822,In_777,In_518);
nor U823 (N_823,In_656,In_159);
and U824 (N_824,In_449,In_648);
nor U825 (N_825,In_34,In_158);
or U826 (N_826,In_664,In_972);
and U827 (N_827,In_780,In_655);
nor U828 (N_828,In_621,In_723);
or U829 (N_829,In_904,In_670);
nand U830 (N_830,In_39,In_464);
nor U831 (N_831,In_261,In_150);
or U832 (N_832,In_216,In_266);
nor U833 (N_833,In_899,In_366);
xor U834 (N_834,In_796,In_103);
nand U835 (N_835,In_920,In_480);
and U836 (N_836,In_681,In_282);
and U837 (N_837,In_957,In_736);
nand U838 (N_838,In_393,In_267);
nor U839 (N_839,In_953,In_191);
nand U840 (N_840,In_698,In_578);
nor U841 (N_841,In_563,In_162);
nand U842 (N_842,In_933,In_809);
nand U843 (N_843,In_276,In_171);
nor U844 (N_844,In_781,In_318);
or U845 (N_845,In_45,In_122);
xor U846 (N_846,In_909,In_597);
and U847 (N_847,In_882,In_22);
or U848 (N_848,In_409,In_878);
nor U849 (N_849,In_671,In_978);
nor U850 (N_850,In_766,In_362);
nand U851 (N_851,In_414,In_498);
and U852 (N_852,In_25,In_940);
and U853 (N_853,In_383,In_769);
and U854 (N_854,In_373,In_572);
and U855 (N_855,In_294,In_820);
and U856 (N_856,In_680,In_722);
nand U857 (N_857,In_775,In_895);
or U858 (N_858,In_543,In_974);
nor U859 (N_859,In_767,In_518);
nand U860 (N_860,In_565,In_838);
nand U861 (N_861,In_466,In_310);
and U862 (N_862,In_167,In_251);
or U863 (N_863,In_305,In_619);
nor U864 (N_864,In_547,In_644);
nand U865 (N_865,In_50,In_416);
or U866 (N_866,In_240,In_706);
or U867 (N_867,In_160,In_76);
and U868 (N_868,In_596,In_383);
nand U869 (N_869,In_982,In_571);
and U870 (N_870,In_533,In_772);
or U871 (N_871,In_415,In_232);
and U872 (N_872,In_33,In_115);
nor U873 (N_873,In_59,In_437);
or U874 (N_874,In_99,In_912);
and U875 (N_875,In_257,In_797);
or U876 (N_876,In_523,In_98);
or U877 (N_877,In_739,In_56);
nand U878 (N_878,In_364,In_901);
nand U879 (N_879,In_685,In_827);
nor U880 (N_880,In_784,In_153);
nand U881 (N_881,In_488,In_565);
nor U882 (N_882,In_45,In_156);
nor U883 (N_883,In_747,In_298);
or U884 (N_884,In_377,In_658);
nor U885 (N_885,In_948,In_156);
or U886 (N_886,In_647,In_517);
or U887 (N_887,In_528,In_150);
nor U888 (N_888,In_908,In_128);
or U889 (N_889,In_175,In_490);
and U890 (N_890,In_217,In_500);
nor U891 (N_891,In_275,In_991);
nor U892 (N_892,In_764,In_597);
or U893 (N_893,In_726,In_957);
and U894 (N_894,In_589,In_495);
nor U895 (N_895,In_67,In_499);
and U896 (N_896,In_113,In_358);
nand U897 (N_897,In_127,In_536);
nor U898 (N_898,In_808,In_381);
or U899 (N_899,In_860,In_972);
and U900 (N_900,In_816,In_170);
or U901 (N_901,In_164,In_978);
nor U902 (N_902,In_474,In_973);
or U903 (N_903,In_104,In_554);
nand U904 (N_904,In_326,In_726);
and U905 (N_905,In_887,In_876);
nand U906 (N_906,In_738,In_451);
nand U907 (N_907,In_564,In_392);
and U908 (N_908,In_451,In_140);
nand U909 (N_909,In_524,In_418);
and U910 (N_910,In_342,In_336);
or U911 (N_911,In_260,In_289);
nor U912 (N_912,In_439,In_566);
nor U913 (N_913,In_854,In_385);
or U914 (N_914,In_457,In_541);
or U915 (N_915,In_298,In_921);
nor U916 (N_916,In_973,In_263);
or U917 (N_917,In_318,In_379);
and U918 (N_918,In_630,In_161);
nor U919 (N_919,In_372,In_156);
nand U920 (N_920,In_850,In_307);
or U921 (N_921,In_590,In_785);
and U922 (N_922,In_315,In_494);
and U923 (N_923,In_615,In_38);
nand U924 (N_924,In_449,In_88);
or U925 (N_925,In_566,In_904);
or U926 (N_926,In_343,In_91);
nand U927 (N_927,In_501,In_617);
and U928 (N_928,In_661,In_695);
nand U929 (N_929,In_686,In_318);
nor U930 (N_930,In_900,In_893);
xor U931 (N_931,In_636,In_324);
nor U932 (N_932,In_428,In_315);
nor U933 (N_933,In_499,In_845);
and U934 (N_934,In_499,In_710);
nand U935 (N_935,In_803,In_110);
nor U936 (N_936,In_515,In_958);
and U937 (N_937,In_88,In_653);
nor U938 (N_938,In_988,In_37);
nand U939 (N_939,In_692,In_538);
nand U940 (N_940,In_442,In_701);
or U941 (N_941,In_471,In_95);
and U942 (N_942,In_120,In_223);
nor U943 (N_943,In_319,In_199);
nand U944 (N_944,In_124,In_576);
nand U945 (N_945,In_201,In_979);
and U946 (N_946,In_782,In_609);
nor U947 (N_947,In_989,In_167);
or U948 (N_948,In_883,In_480);
nand U949 (N_949,In_523,In_473);
or U950 (N_950,In_185,In_900);
nor U951 (N_951,In_467,In_137);
and U952 (N_952,In_450,In_265);
and U953 (N_953,In_916,In_138);
and U954 (N_954,In_359,In_433);
nor U955 (N_955,In_531,In_777);
or U956 (N_956,In_978,In_388);
and U957 (N_957,In_4,In_111);
nor U958 (N_958,In_757,In_63);
nor U959 (N_959,In_114,In_518);
and U960 (N_960,In_626,In_697);
and U961 (N_961,In_63,In_732);
nor U962 (N_962,In_830,In_738);
nor U963 (N_963,In_438,In_375);
nand U964 (N_964,In_323,In_383);
nand U965 (N_965,In_995,In_181);
nand U966 (N_966,In_54,In_335);
or U967 (N_967,In_187,In_974);
nor U968 (N_968,In_739,In_663);
and U969 (N_969,In_478,In_96);
nor U970 (N_970,In_468,In_43);
and U971 (N_971,In_223,In_343);
nand U972 (N_972,In_477,In_232);
or U973 (N_973,In_930,In_729);
nand U974 (N_974,In_91,In_78);
and U975 (N_975,In_737,In_729);
nor U976 (N_976,In_191,In_6);
and U977 (N_977,In_640,In_952);
or U978 (N_978,In_480,In_356);
nand U979 (N_979,In_672,In_961);
nand U980 (N_980,In_320,In_172);
and U981 (N_981,In_405,In_164);
and U982 (N_982,In_207,In_90);
and U983 (N_983,In_834,In_974);
or U984 (N_984,In_843,In_319);
nor U985 (N_985,In_558,In_525);
nand U986 (N_986,In_21,In_737);
and U987 (N_987,In_469,In_807);
or U988 (N_988,In_252,In_358);
nor U989 (N_989,In_750,In_272);
and U990 (N_990,In_986,In_522);
or U991 (N_991,In_800,In_614);
nor U992 (N_992,In_302,In_820);
or U993 (N_993,In_75,In_687);
or U994 (N_994,In_472,In_552);
nor U995 (N_995,In_344,In_479);
nand U996 (N_996,In_349,In_569);
nand U997 (N_997,In_213,In_395);
or U998 (N_998,In_372,In_66);
or U999 (N_999,In_344,In_273);
nor U1000 (N_1000,N_393,N_786);
nor U1001 (N_1001,N_396,N_859);
nand U1002 (N_1002,N_98,N_759);
or U1003 (N_1003,N_325,N_671);
nand U1004 (N_1004,N_417,N_8);
nor U1005 (N_1005,N_824,N_23);
or U1006 (N_1006,N_525,N_904);
nand U1007 (N_1007,N_157,N_494);
nor U1008 (N_1008,N_269,N_988);
and U1009 (N_1009,N_320,N_902);
and U1010 (N_1010,N_560,N_910);
or U1011 (N_1011,N_749,N_339);
nand U1012 (N_1012,N_57,N_827);
and U1013 (N_1013,N_272,N_893);
nor U1014 (N_1014,N_475,N_590);
or U1015 (N_1015,N_582,N_20);
and U1016 (N_1016,N_943,N_929);
nand U1017 (N_1017,N_68,N_561);
nand U1018 (N_1018,N_507,N_428);
nor U1019 (N_1019,N_956,N_241);
or U1020 (N_1020,N_826,N_932);
nand U1021 (N_1021,N_328,N_692);
nand U1022 (N_1022,N_481,N_687);
or U1023 (N_1023,N_331,N_406);
nor U1024 (N_1024,N_142,N_482);
nand U1025 (N_1025,N_657,N_354);
nor U1026 (N_1026,N_126,N_222);
nor U1027 (N_1027,N_338,N_849);
and U1028 (N_1028,N_350,N_413);
nand U1029 (N_1029,N_670,N_776);
and U1030 (N_1030,N_566,N_962);
and U1031 (N_1031,N_882,N_974);
nand U1032 (N_1032,N_872,N_65);
or U1033 (N_1033,N_4,N_123);
nand U1034 (N_1034,N_33,N_627);
or U1035 (N_1035,N_758,N_994);
or U1036 (N_1036,N_42,N_992);
or U1037 (N_1037,N_490,N_835);
or U1038 (N_1038,N_392,N_295);
or U1039 (N_1039,N_293,N_263);
xor U1040 (N_1040,N_517,N_258);
nand U1041 (N_1041,N_764,N_686);
and U1042 (N_1042,N_822,N_104);
nor U1043 (N_1043,N_616,N_281);
nor U1044 (N_1044,N_972,N_179);
nor U1045 (N_1045,N_573,N_506);
or U1046 (N_1046,N_909,N_397);
and U1047 (N_1047,N_153,N_92);
nand U1048 (N_1048,N_586,N_809);
and U1049 (N_1049,N_915,N_869);
nand U1050 (N_1050,N_619,N_343);
or U1051 (N_1051,N_21,N_923);
nor U1052 (N_1052,N_733,N_930);
nand U1053 (N_1053,N_989,N_543);
nor U1054 (N_1054,N_645,N_846);
nand U1055 (N_1055,N_300,N_301);
and U1056 (N_1056,N_926,N_27);
or U1057 (N_1057,N_850,N_399);
or U1058 (N_1058,N_219,N_287);
nand U1059 (N_1059,N_933,N_620);
and U1060 (N_1060,N_492,N_424);
nand U1061 (N_1061,N_961,N_866);
and U1062 (N_1062,N_87,N_792);
or U1063 (N_1063,N_650,N_177);
nand U1064 (N_1064,N_775,N_461);
or U1065 (N_1065,N_767,N_358);
nor U1066 (N_1066,N_878,N_407);
and U1067 (N_1067,N_444,N_836);
nand U1068 (N_1068,N_533,N_204);
nor U1069 (N_1069,N_9,N_430);
nor U1070 (N_1070,N_739,N_696);
nor U1071 (N_1071,N_435,N_556);
nor U1072 (N_1072,N_711,N_569);
or U1073 (N_1073,N_449,N_381);
nand U1074 (N_1074,N_372,N_508);
nand U1075 (N_1075,N_754,N_433);
nor U1076 (N_1076,N_519,N_538);
or U1077 (N_1077,N_986,N_110);
and U1078 (N_1078,N_160,N_732);
or U1079 (N_1079,N_515,N_385);
and U1080 (N_1080,N_292,N_924);
nor U1081 (N_1081,N_383,N_768);
nor U1082 (N_1082,N_638,N_441);
nand U1083 (N_1083,N_159,N_847);
and U1084 (N_1084,N_439,N_315);
and U1085 (N_1085,N_797,N_857);
or U1086 (N_1086,N_18,N_800);
nor U1087 (N_1087,N_855,N_744);
nor U1088 (N_1088,N_349,N_120);
and U1089 (N_1089,N_969,N_984);
or U1090 (N_1090,N_564,N_689);
nand U1091 (N_1091,N_52,N_361);
nand U1092 (N_1092,N_243,N_649);
nand U1093 (N_1093,N_636,N_679);
nand U1094 (N_1094,N_576,N_861);
and U1095 (N_1095,N_553,N_675);
and U1096 (N_1096,N_922,N_498);
nand U1097 (N_1097,N_359,N_410);
or U1098 (N_1098,N_753,N_997);
and U1099 (N_1099,N_114,N_39);
nor U1100 (N_1100,N_682,N_524);
and U1101 (N_1101,N_26,N_446);
nand U1102 (N_1102,N_523,N_728);
or U1103 (N_1103,N_587,N_617);
or U1104 (N_1104,N_874,N_427);
nand U1105 (N_1105,N_830,N_963);
and U1106 (N_1106,N_780,N_803);
nor U1107 (N_1107,N_939,N_966);
and U1108 (N_1108,N_752,N_970);
or U1109 (N_1109,N_256,N_408);
or U1110 (N_1110,N_979,N_594);
nor U1111 (N_1111,N_419,N_633);
and U1112 (N_1112,N_395,N_693);
nor U1113 (N_1113,N_379,N_337);
and U1114 (N_1114,N_40,N_355);
nor U1115 (N_1115,N_672,N_680);
nor U1116 (N_1116,N_94,N_56);
nand U1117 (N_1117,N_363,N_815);
nor U1118 (N_1118,N_278,N_255);
and U1119 (N_1119,N_409,N_388);
and U1120 (N_1120,N_17,N_314);
and U1121 (N_1121,N_676,N_163);
and U1122 (N_1122,N_335,N_290);
and U1123 (N_1123,N_511,N_225);
or U1124 (N_1124,N_734,N_28);
nor U1125 (N_1125,N_387,N_921);
nor U1126 (N_1126,N_11,N_181);
or U1127 (N_1127,N_852,N_390);
nand U1128 (N_1128,N_964,N_124);
nand U1129 (N_1129,N_199,N_602);
nor U1130 (N_1130,N_581,N_871);
nand U1131 (N_1131,N_109,N_164);
or U1132 (N_1132,N_371,N_274);
or U1133 (N_1133,N_660,N_210);
nand U1134 (N_1134,N_634,N_726);
and U1135 (N_1135,N_656,N_900);
nand U1136 (N_1136,N_832,N_356);
nor U1137 (N_1137,N_457,N_466);
or U1138 (N_1138,N_280,N_968);
or U1139 (N_1139,N_63,N_777);
nand U1140 (N_1140,N_112,N_260);
or U1141 (N_1141,N_230,N_863);
nor U1142 (N_1142,N_426,N_699);
nor U1143 (N_1143,N_738,N_931);
and U1144 (N_1144,N_389,N_25);
nor U1145 (N_1145,N_980,N_530);
or U1146 (N_1146,N_659,N_722);
nand U1147 (N_1147,N_705,N_249);
nand U1148 (N_1148,N_478,N_78);
or U1149 (N_1149,N_622,N_958);
or U1150 (N_1150,N_305,N_520);
or U1151 (N_1151,N_978,N_479);
or U1152 (N_1152,N_505,N_631);
and U1153 (N_1153,N_7,N_628);
nor U1154 (N_1154,N_80,N_61);
or U1155 (N_1155,N_366,N_845);
nor U1156 (N_1156,N_745,N_599);
nor U1157 (N_1157,N_470,N_833);
or U1158 (N_1158,N_129,N_575);
nand U1159 (N_1159,N_499,N_431);
nor U1160 (N_1160,N_373,N_196);
or U1161 (N_1161,N_595,N_510);
or U1162 (N_1162,N_724,N_664);
and U1163 (N_1163,N_546,N_171);
nand U1164 (N_1164,N_232,N_898);
or U1165 (N_1165,N_261,N_793);
or U1166 (N_1166,N_558,N_193);
and U1167 (N_1167,N_941,N_48);
and U1168 (N_1168,N_90,N_303);
nand U1169 (N_1169,N_844,N_116);
nand U1170 (N_1170,N_731,N_772);
and U1171 (N_1171,N_578,N_496);
or U1172 (N_1172,N_117,N_662);
or U1173 (N_1173,N_987,N_140);
nor U1174 (N_1174,N_999,N_486);
nand U1175 (N_1175,N_954,N_162);
nand U1176 (N_1176,N_405,N_240);
nand U1177 (N_1177,N_730,N_512);
nand U1178 (N_1178,N_125,N_54);
nor U1179 (N_1179,N_723,N_197);
xor U1180 (N_1180,N_115,N_97);
nand U1181 (N_1181,N_429,N_445);
and U1182 (N_1182,N_840,N_134);
nor U1183 (N_1183,N_531,N_853);
and U1184 (N_1184,N_59,N_465);
or U1185 (N_1185,N_837,N_237);
and U1186 (N_1186,N_357,N_995);
nand U1187 (N_1187,N_841,N_459);
nor U1188 (N_1188,N_100,N_217);
nand U1189 (N_1189,N_453,N_567);
or U1190 (N_1190,N_147,N_487);
nand U1191 (N_1191,N_598,N_86);
or U1192 (N_1192,N_542,N_299);
nand U1193 (N_1193,N_655,N_539);
or U1194 (N_1194,N_37,N_72);
and U1195 (N_1195,N_351,N_574);
nand U1196 (N_1196,N_600,N_514);
or U1197 (N_1197,N_294,N_654);
nor U1198 (N_1198,N_151,N_121);
nand U1199 (N_1199,N_469,N_176);
nor U1200 (N_1200,N_262,N_306);
nor U1201 (N_1201,N_534,N_990);
nor U1202 (N_1202,N_765,N_19);
nor U1203 (N_1203,N_808,N_206);
nor U1204 (N_1204,N_761,N_137);
or U1205 (N_1205,N_432,N_828);
and U1206 (N_1206,N_811,N_370);
and U1207 (N_1207,N_736,N_597);
or U1208 (N_1208,N_794,N_344);
and U1209 (N_1209,N_106,N_603);
or U1210 (N_1210,N_981,N_532);
and U1211 (N_1211,N_279,N_960);
or U1212 (N_1212,N_756,N_220);
nand U1213 (N_1213,N_681,N_161);
and U1214 (N_1214,N_875,N_288);
nand U1215 (N_1215,N_377,N_77);
or U1216 (N_1216,N_796,N_639);
nor U1217 (N_1217,N_813,N_75);
nand U1218 (N_1218,N_170,N_669);
and U1219 (N_1219,N_606,N_937);
nor U1220 (N_1220,N_697,N_685);
nor U1221 (N_1221,N_259,N_559);
or U1222 (N_1222,N_973,N_477);
nand U1223 (N_1223,N_580,N_942);
and U1224 (N_1224,N_302,N_326);
nand U1225 (N_1225,N_551,N_688);
or U1226 (N_1226,N_703,N_312);
nand U1227 (N_1227,N_491,N_577);
and U1228 (N_1228,N_952,N_899);
nand U1229 (N_1229,N_829,N_787);
or U1230 (N_1230,N_275,N_545);
nand U1231 (N_1231,N_950,N_795);
and U1232 (N_1232,N_601,N_493);
or U1233 (N_1233,N_69,N_721);
nand U1234 (N_1234,N_47,N_329);
nor U1235 (N_1235,N_651,N_239);
nor U1236 (N_1236,N_812,N_216);
and U1237 (N_1237,N_831,N_854);
or U1238 (N_1238,N_858,N_641);
nor U1239 (N_1239,N_43,N_485);
nor U1240 (N_1240,N_34,N_630);
and U1241 (N_1241,N_897,N_977);
nand U1242 (N_1242,N_423,N_884);
nand U1243 (N_1243,N_15,N_951);
or U1244 (N_1244,N_64,N_557);
and U1245 (N_1245,N_848,N_190);
nor U1246 (N_1246,N_165,N_127);
and U1247 (N_1247,N_903,N_865);
nand U1248 (N_1248,N_462,N_13);
and U1249 (N_1249,N_266,N_402);
nand U1250 (N_1250,N_476,N_3);
and U1251 (N_1251,N_653,N_905);
or U1252 (N_1252,N_130,N_332);
and U1253 (N_1253,N_113,N_548);
and U1254 (N_1254,N_149,N_746);
nand U1255 (N_1255,N_30,N_6);
or U1256 (N_1256,N_228,N_801);
or U1257 (N_1257,N_535,N_621);
nor U1258 (N_1258,N_509,N_626);
nand U1259 (N_1259,N_102,N_178);
nand U1260 (N_1260,N_788,N_414);
and U1261 (N_1261,N_713,N_484);
and U1262 (N_1262,N_362,N_513);
or U1263 (N_1263,N_296,N_319);
nor U1264 (N_1264,N_250,N_562);
nor U1265 (N_1265,N_825,N_760);
nand U1266 (N_1266,N_489,N_547);
nand U1267 (N_1267,N_234,N_781);
and U1268 (N_1268,N_73,N_145);
and U1269 (N_1269,N_702,N_136);
and U1270 (N_1270,N_707,N_76);
nand U1271 (N_1271,N_53,N_386);
and U1272 (N_1272,N_271,N_2);
and U1273 (N_1273,N_762,N_254);
nand U1274 (N_1274,N_82,N_890);
and U1275 (N_1275,N_782,N_246);
or U1276 (N_1276,N_183,N_483);
nand U1277 (N_1277,N_528,N_154);
or U1278 (N_1278,N_504,N_155);
nand U1279 (N_1279,N_919,N_471);
nand U1280 (N_1280,N_215,N_286);
nand U1281 (N_1281,N_62,N_174);
nor U1282 (N_1282,N_717,N_816);
nor U1283 (N_1283,N_32,N_404);
or U1284 (N_1284,N_224,N_527);
and U1285 (N_1285,N_152,N_273);
and U1286 (N_1286,N_500,N_438);
and U1287 (N_1287,N_544,N_265);
nor U1288 (N_1288,N_554,N_873);
nor U1289 (N_1289,N_862,N_0);
nor U1290 (N_1290,N_785,N_60);
or U1291 (N_1291,N_537,N_901);
nand U1292 (N_1292,N_743,N_85);
nand U1293 (N_1293,N_522,N_172);
and U1294 (N_1294,N_195,N_66);
nor U1295 (N_1295,N_755,N_341);
or U1296 (N_1296,N_322,N_189);
or U1297 (N_1297,N_516,N_695);
and U1298 (N_1298,N_253,N_623);
or U1299 (N_1299,N_823,N_360);
or U1300 (N_1300,N_367,N_211);
and U1301 (N_1301,N_188,N_173);
and U1302 (N_1302,N_235,N_70);
nand U1303 (N_1303,N_766,N_991);
nor U1304 (N_1304,N_742,N_593);
and U1305 (N_1305,N_105,N_16);
and U1306 (N_1306,N_447,N_276);
nor U1307 (N_1307,N_876,N_88);
nor U1308 (N_1308,N_985,N_229);
and U1309 (N_1309,N_497,N_297);
and U1310 (N_1310,N_867,N_169);
and U1311 (N_1311,N_944,N_690);
nor U1312 (N_1312,N_710,N_838);
and U1313 (N_1313,N_719,N_443);
nor U1314 (N_1314,N_84,N_5);
nor U1315 (N_1315,N_139,N_691);
or U1316 (N_1316,N_579,N_916);
nand U1317 (N_1317,N_378,N_187);
or U1318 (N_1318,N_818,N_913);
nand U1319 (N_1319,N_185,N_194);
and U1320 (N_1320,N_223,N_227);
or U1321 (N_1321,N_918,N_665);
or U1322 (N_1322,N_167,N_894);
nand U1323 (N_1323,N_394,N_868);
nand U1324 (N_1324,N_771,N_425);
and U1325 (N_1325,N_291,N_906);
and U1326 (N_1326,N_971,N_834);
nor U1327 (N_1327,N_365,N_46);
and U1328 (N_1328,N_436,N_624);
nand U1329 (N_1329,N_783,N_321);
nor U1330 (N_1330,N_678,N_198);
and U1331 (N_1331,N_463,N_442);
nand U1332 (N_1332,N_625,N_420);
nand U1333 (N_1333,N_474,N_309);
nor U1334 (N_1334,N_141,N_945);
nand U1335 (N_1335,N_632,N_150);
or U1336 (N_1336,N_928,N_311);
or U1337 (N_1337,N_454,N_652);
or U1338 (N_1338,N_244,N_403);
nor U1339 (N_1339,N_440,N_773);
nand U1340 (N_1340,N_208,N_552);
or U1341 (N_1341,N_45,N_99);
and U1342 (N_1342,N_422,N_851);
nor U1343 (N_1343,N_93,N_807);
nand U1344 (N_1344,N_938,N_375);
or U1345 (N_1345,N_608,N_468);
and U1346 (N_1346,N_864,N_698);
nand U1347 (N_1347,N_79,N_10);
and U1348 (N_1348,N_748,N_175);
and U1349 (N_1349,N_791,N_236);
nor U1350 (N_1350,N_247,N_317);
and U1351 (N_1351,N_648,N_646);
and U1352 (N_1352,N_750,N_975);
nor U1353 (N_1353,N_327,N_814);
nand U1354 (N_1354,N_38,N_666);
nor U1355 (N_1355,N_401,N_284);
or U1356 (N_1356,N_618,N_877);
nand U1357 (N_1357,N_89,N_612);
nor U1358 (N_1358,N_455,N_763);
and U1359 (N_1359,N_451,N_609);
and U1360 (N_1360,N_374,N_36);
or U1361 (N_1361,N_607,N_22);
and U1362 (N_1362,N_158,N_166);
nor U1363 (N_1363,N_12,N_983);
and U1364 (N_1364,N_71,N_316);
nor U1365 (N_1365,N_770,N_345);
or U1366 (N_1366,N_501,N_131);
nand U1367 (N_1367,N_668,N_885);
nand U1368 (N_1368,N_720,N_550);
and U1369 (N_1369,N_368,N_629);
nor U1370 (N_1370,N_448,N_572);
nand U1371 (N_1371,N_585,N_31);
nor U1372 (N_1372,N_207,N_996);
nand U1373 (N_1373,N_982,N_673);
xor U1374 (N_1374,N_596,N_143);
nand U1375 (N_1375,N_967,N_122);
and U1376 (N_1376,N_555,N_583);
nor U1377 (N_1377,N_310,N_146);
or U1378 (N_1378,N_267,N_503);
or U1379 (N_1379,N_464,N_103);
nor U1380 (N_1380,N_714,N_334);
or U1381 (N_1381,N_421,N_391);
or U1382 (N_1382,N_200,N_709);
nor U1383 (N_1383,N_128,N_398);
or U1384 (N_1384,N_589,N_49);
nand U1385 (N_1385,N_382,N_214);
and U1386 (N_1386,N_896,N_285);
or U1387 (N_1387,N_44,N_58);
or U1388 (N_1388,N_615,N_107);
nand U1389 (N_1389,N_456,N_96);
or U1390 (N_1390,N_584,N_257);
or U1391 (N_1391,N_434,N_270);
or U1392 (N_1392,N_614,N_252);
nand U1393 (N_1393,N_674,N_184);
or U1394 (N_1394,N_412,N_592);
nor U1395 (N_1395,N_737,N_415);
nand U1396 (N_1396,N_708,N_324);
nand U1397 (N_1397,N_998,N_218);
or U1398 (N_1398,N_101,N_144);
and U1399 (N_1399,N_330,N_135);
and U1400 (N_1400,N_238,N_821);
or U1401 (N_1401,N_908,N_799);
nand U1402 (N_1402,N_473,N_661);
or U1403 (N_1403,N_643,N_138);
or U1404 (N_1404,N_203,N_804);
nand U1405 (N_1405,N_307,N_571);
nand U1406 (N_1406,N_888,N_192);
nand U1407 (N_1407,N_226,N_340);
nor U1408 (N_1408,N_384,N_29);
or U1409 (N_1409,N_817,N_725);
nor U1410 (N_1410,N_502,N_955);
and U1411 (N_1411,N_935,N_55);
nor U1412 (N_1412,N_706,N_318);
nand U1413 (N_1413,N_283,N_488);
nor U1414 (N_1414,N_348,N_298);
or U1415 (N_1415,N_352,N_953);
nor U1416 (N_1416,N_191,N_936);
and U1417 (N_1417,N_346,N_540);
nor U1418 (N_1418,N_186,N_480);
or U1419 (N_1419,N_251,N_642);
or U1420 (N_1420,N_95,N_778);
or U1421 (N_1421,N_886,N_880);
xnor U1422 (N_1422,N_245,N_640);
or U1423 (N_1423,N_604,N_467);
nand U1424 (N_1424,N_289,N_336);
and U1425 (N_1425,N_774,N_111);
and U1426 (N_1426,N_458,N_380);
nand U1427 (N_1427,N_605,N_74);
and U1428 (N_1428,N_927,N_347);
nand U1429 (N_1429,N_213,N_91);
or U1430 (N_1430,N_323,N_934);
and U1431 (N_1431,N_565,N_735);
and U1432 (N_1432,N_637,N_148);
nand U1433 (N_1433,N_700,N_647);
nand U1434 (N_1434,N_839,N_677);
and U1435 (N_1435,N_304,N_51);
and U1436 (N_1436,N_83,N_920);
nor U1437 (N_1437,N_856,N_694);
nand U1438 (N_1438,N_883,N_993);
or U1439 (N_1439,N_518,N_820);
or U1440 (N_1440,N_221,N_369);
nand U1441 (N_1441,N_264,N_205);
or U1442 (N_1442,N_400,N_716);
nor U1443 (N_1443,N_570,N_715);
and U1444 (N_1444,N_959,N_747);
nor U1445 (N_1445,N_1,N_946);
nand U1446 (N_1446,N_891,N_805);
or U1447 (N_1447,N_683,N_156);
and U1448 (N_1448,N_118,N_976);
or U1449 (N_1449,N_907,N_757);
nor U1450 (N_1450,N_740,N_802);
nand U1451 (N_1451,N_282,N_843);
and U1452 (N_1452,N_806,N_119);
nor U1453 (N_1453,N_644,N_411);
nand U1454 (N_1454,N_889,N_712);
nand U1455 (N_1455,N_248,N_526);
nand U1456 (N_1456,N_308,N_212);
nand U1457 (N_1457,N_233,N_667);
nand U1458 (N_1458,N_789,N_704);
nor U1459 (N_1459,N_588,N_133);
or U1460 (N_1460,N_610,N_277);
and U1461 (N_1461,N_563,N_914);
and U1462 (N_1462,N_611,N_729);
or U1463 (N_1463,N_450,N_947);
nand U1464 (N_1464,N_613,N_741);
and U1465 (N_1465,N_231,N_940);
nand U1466 (N_1466,N_472,N_35);
nor U1467 (N_1467,N_549,N_168);
or U1468 (N_1468,N_810,N_591);
and U1469 (N_1469,N_881,N_658);
nor U1470 (N_1470,N_108,N_268);
nand U1471 (N_1471,N_701,N_541);
nand U1472 (N_1472,N_949,N_912);
or U1473 (N_1473,N_529,N_536);
and U1474 (N_1474,N_887,N_842);
or U1475 (N_1475,N_460,N_452);
or U1476 (N_1476,N_684,N_24);
and U1477 (N_1477,N_879,N_416);
and U1478 (N_1478,N_418,N_779);
nand U1479 (N_1479,N_860,N_769);
nand U1480 (N_1480,N_202,N_495);
or U1481 (N_1481,N_50,N_727);
nand U1482 (N_1482,N_568,N_751);
nor U1483 (N_1483,N_790,N_819);
nor U1484 (N_1484,N_635,N_333);
nand U1485 (N_1485,N_342,N_353);
or U1486 (N_1486,N_925,N_718);
and U1487 (N_1487,N_663,N_521);
nor U1488 (N_1488,N_870,N_895);
nand U1489 (N_1489,N_67,N_182);
or U1490 (N_1490,N_892,N_957);
nor U1491 (N_1491,N_313,N_132);
nand U1492 (N_1492,N_201,N_14);
and U1493 (N_1493,N_41,N_784);
nand U1494 (N_1494,N_364,N_81);
nor U1495 (N_1495,N_180,N_917);
or U1496 (N_1496,N_242,N_437);
or U1497 (N_1497,N_948,N_798);
nor U1498 (N_1498,N_209,N_911);
nor U1499 (N_1499,N_376,N_965);
or U1500 (N_1500,N_823,N_346);
and U1501 (N_1501,N_411,N_433);
and U1502 (N_1502,N_143,N_656);
and U1503 (N_1503,N_991,N_450);
or U1504 (N_1504,N_910,N_28);
nand U1505 (N_1505,N_135,N_767);
nand U1506 (N_1506,N_168,N_302);
or U1507 (N_1507,N_203,N_18);
xnor U1508 (N_1508,N_109,N_976);
xor U1509 (N_1509,N_743,N_187);
or U1510 (N_1510,N_575,N_62);
or U1511 (N_1511,N_14,N_485);
nand U1512 (N_1512,N_313,N_798);
xnor U1513 (N_1513,N_222,N_991);
or U1514 (N_1514,N_147,N_706);
nand U1515 (N_1515,N_833,N_860);
or U1516 (N_1516,N_160,N_610);
nand U1517 (N_1517,N_371,N_358);
and U1518 (N_1518,N_838,N_91);
nand U1519 (N_1519,N_302,N_311);
nor U1520 (N_1520,N_746,N_558);
nand U1521 (N_1521,N_147,N_215);
nor U1522 (N_1522,N_717,N_325);
nand U1523 (N_1523,N_958,N_238);
and U1524 (N_1524,N_725,N_574);
and U1525 (N_1525,N_516,N_460);
and U1526 (N_1526,N_326,N_969);
nor U1527 (N_1527,N_313,N_245);
nand U1528 (N_1528,N_949,N_864);
and U1529 (N_1529,N_363,N_834);
nand U1530 (N_1530,N_850,N_273);
and U1531 (N_1531,N_637,N_457);
and U1532 (N_1532,N_743,N_943);
nor U1533 (N_1533,N_711,N_3);
and U1534 (N_1534,N_100,N_337);
and U1535 (N_1535,N_416,N_254);
and U1536 (N_1536,N_233,N_633);
nor U1537 (N_1537,N_68,N_93);
nand U1538 (N_1538,N_133,N_995);
or U1539 (N_1539,N_68,N_942);
nand U1540 (N_1540,N_677,N_96);
nand U1541 (N_1541,N_748,N_273);
nor U1542 (N_1542,N_96,N_917);
nor U1543 (N_1543,N_946,N_467);
nand U1544 (N_1544,N_387,N_796);
or U1545 (N_1545,N_628,N_55);
or U1546 (N_1546,N_718,N_930);
or U1547 (N_1547,N_953,N_796);
or U1548 (N_1548,N_473,N_869);
or U1549 (N_1549,N_718,N_754);
or U1550 (N_1550,N_328,N_384);
and U1551 (N_1551,N_453,N_288);
and U1552 (N_1552,N_698,N_456);
nand U1553 (N_1553,N_153,N_226);
nand U1554 (N_1554,N_328,N_77);
nand U1555 (N_1555,N_258,N_636);
or U1556 (N_1556,N_408,N_432);
and U1557 (N_1557,N_468,N_752);
or U1558 (N_1558,N_530,N_681);
or U1559 (N_1559,N_664,N_316);
and U1560 (N_1560,N_649,N_511);
nand U1561 (N_1561,N_3,N_478);
and U1562 (N_1562,N_535,N_646);
and U1563 (N_1563,N_423,N_314);
and U1564 (N_1564,N_256,N_938);
nand U1565 (N_1565,N_336,N_627);
xnor U1566 (N_1566,N_146,N_159);
nand U1567 (N_1567,N_612,N_517);
nand U1568 (N_1568,N_523,N_28);
nor U1569 (N_1569,N_238,N_526);
and U1570 (N_1570,N_147,N_94);
or U1571 (N_1571,N_847,N_564);
nor U1572 (N_1572,N_927,N_62);
nor U1573 (N_1573,N_928,N_512);
or U1574 (N_1574,N_662,N_813);
or U1575 (N_1575,N_454,N_597);
and U1576 (N_1576,N_830,N_84);
or U1577 (N_1577,N_266,N_255);
and U1578 (N_1578,N_481,N_584);
xor U1579 (N_1579,N_561,N_437);
or U1580 (N_1580,N_229,N_52);
nor U1581 (N_1581,N_793,N_703);
or U1582 (N_1582,N_425,N_542);
and U1583 (N_1583,N_115,N_947);
nor U1584 (N_1584,N_572,N_637);
nor U1585 (N_1585,N_201,N_151);
or U1586 (N_1586,N_86,N_279);
nor U1587 (N_1587,N_970,N_873);
and U1588 (N_1588,N_287,N_72);
or U1589 (N_1589,N_363,N_233);
and U1590 (N_1590,N_558,N_94);
nor U1591 (N_1591,N_365,N_558);
nor U1592 (N_1592,N_937,N_70);
and U1593 (N_1593,N_147,N_861);
or U1594 (N_1594,N_262,N_5);
and U1595 (N_1595,N_648,N_856);
xnor U1596 (N_1596,N_907,N_453);
or U1597 (N_1597,N_783,N_577);
nor U1598 (N_1598,N_624,N_267);
and U1599 (N_1599,N_177,N_804);
nor U1600 (N_1600,N_129,N_398);
or U1601 (N_1601,N_749,N_977);
or U1602 (N_1602,N_67,N_686);
nand U1603 (N_1603,N_787,N_25);
nor U1604 (N_1604,N_931,N_601);
nor U1605 (N_1605,N_149,N_524);
or U1606 (N_1606,N_693,N_15);
and U1607 (N_1607,N_684,N_730);
nand U1608 (N_1608,N_584,N_389);
or U1609 (N_1609,N_210,N_992);
nor U1610 (N_1610,N_188,N_390);
nand U1611 (N_1611,N_165,N_750);
nand U1612 (N_1612,N_165,N_147);
nor U1613 (N_1613,N_78,N_118);
nor U1614 (N_1614,N_275,N_448);
and U1615 (N_1615,N_732,N_717);
or U1616 (N_1616,N_167,N_824);
or U1617 (N_1617,N_331,N_905);
and U1618 (N_1618,N_244,N_742);
xor U1619 (N_1619,N_445,N_618);
nand U1620 (N_1620,N_548,N_148);
and U1621 (N_1621,N_793,N_43);
or U1622 (N_1622,N_917,N_18);
or U1623 (N_1623,N_226,N_319);
nor U1624 (N_1624,N_370,N_820);
nand U1625 (N_1625,N_703,N_902);
or U1626 (N_1626,N_528,N_96);
nand U1627 (N_1627,N_854,N_681);
or U1628 (N_1628,N_874,N_51);
nor U1629 (N_1629,N_206,N_247);
or U1630 (N_1630,N_984,N_184);
or U1631 (N_1631,N_72,N_536);
nor U1632 (N_1632,N_774,N_810);
and U1633 (N_1633,N_713,N_115);
nand U1634 (N_1634,N_675,N_49);
and U1635 (N_1635,N_398,N_254);
nor U1636 (N_1636,N_198,N_286);
and U1637 (N_1637,N_39,N_680);
nand U1638 (N_1638,N_107,N_413);
or U1639 (N_1639,N_24,N_319);
nand U1640 (N_1640,N_761,N_461);
and U1641 (N_1641,N_151,N_262);
nor U1642 (N_1642,N_715,N_912);
nor U1643 (N_1643,N_557,N_871);
nand U1644 (N_1644,N_800,N_198);
nand U1645 (N_1645,N_708,N_572);
nor U1646 (N_1646,N_315,N_37);
and U1647 (N_1647,N_736,N_339);
and U1648 (N_1648,N_849,N_792);
nand U1649 (N_1649,N_54,N_513);
nor U1650 (N_1650,N_438,N_944);
and U1651 (N_1651,N_191,N_621);
or U1652 (N_1652,N_225,N_463);
nor U1653 (N_1653,N_471,N_983);
nor U1654 (N_1654,N_461,N_685);
or U1655 (N_1655,N_446,N_981);
nor U1656 (N_1656,N_61,N_587);
and U1657 (N_1657,N_760,N_182);
nand U1658 (N_1658,N_277,N_263);
nand U1659 (N_1659,N_835,N_334);
and U1660 (N_1660,N_810,N_745);
or U1661 (N_1661,N_561,N_729);
or U1662 (N_1662,N_558,N_178);
or U1663 (N_1663,N_134,N_273);
nor U1664 (N_1664,N_604,N_615);
or U1665 (N_1665,N_175,N_71);
and U1666 (N_1666,N_266,N_946);
and U1667 (N_1667,N_926,N_404);
and U1668 (N_1668,N_399,N_36);
or U1669 (N_1669,N_601,N_570);
nand U1670 (N_1670,N_511,N_510);
or U1671 (N_1671,N_314,N_413);
and U1672 (N_1672,N_955,N_699);
nand U1673 (N_1673,N_192,N_347);
nor U1674 (N_1674,N_451,N_241);
nand U1675 (N_1675,N_701,N_603);
nor U1676 (N_1676,N_324,N_783);
nand U1677 (N_1677,N_367,N_657);
or U1678 (N_1678,N_340,N_178);
nor U1679 (N_1679,N_57,N_699);
nor U1680 (N_1680,N_385,N_29);
and U1681 (N_1681,N_624,N_820);
or U1682 (N_1682,N_870,N_164);
nand U1683 (N_1683,N_940,N_639);
nand U1684 (N_1684,N_732,N_443);
nand U1685 (N_1685,N_449,N_526);
nor U1686 (N_1686,N_203,N_813);
and U1687 (N_1687,N_63,N_587);
and U1688 (N_1688,N_841,N_969);
nand U1689 (N_1689,N_708,N_448);
nor U1690 (N_1690,N_95,N_275);
nor U1691 (N_1691,N_19,N_780);
and U1692 (N_1692,N_393,N_299);
or U1693 (N_1693,N_138,N_431);
or U1694 (N_1694,N_332,N_616);
nor U1695 (N_1695,N_251,N_394);
xor U1696 (N_1696,N_485,N_777);
or U1697 (N_1697,N_937,N_589);
or U1698 (N_1698,N_751,N_67);
or U1699 (N_1699,N_833,N_864);
nor U1700 (N_1700,N_558,N_369);
or U1701 (N_1701,N_967,N_494);
nand U1702 (N_1702,N_301,N_860);
nor U1703 (N_1703,N_509,N_566);
nor U1704 (N_1704,N_780,N_3);
and U1705 (N_1705,N_994,N_662);
and U1706 (N_1706,N_671,N_740);
and U1707 (N_1707,N_584,N_87);
and U1708 (N_1708,N_783,N_454);
or U1709 (N_1709,N_768,N_453);
nand U1710 (N_1710,N_105,N_90);
nand U1711 (N_1711,N_486,N_690);
nand U1712 (N_1712,N_696,N_533);
or U1713 (N_1713,N_698,N_694);
nand U1714 (N_1714,N_947,N_566);
nor U1715 (N_1715,N_217,N_310);
or U1716 (N_1716,N_848,N_55);
nor U1717 (N_1717,N_848,N_414);
nand U1718 (N_1718,N_649,N_21);
and U1719 (N_1719,N_242,N_987);
or U1720 (N_1720,N_843,N_270);
xnor U1721 (N_1721,N_709,N_203);
nand U1722 (N_1722,N_587,N_579);
and U1723 (N_1723,N_252,N_280);
and U1724 (N_1724,N_844,N_157);
or U1725 (N_1725,N_177,N_482);
and U1726 (N_1726,N_305,N_664);
and U1727 (N_1727,N_537,N_479);
nor U1728 (N_1728,N_349,N_497);
or U1729 (N_1729,N_401,N_376);
nor U1730 (N_1730,N_430,N_608);
and U1731 (N_1731,N_92,N_612);
nand U1732 (N_1732,N_631,N_563);
nor U1733 (N_1733,N_588,N_62);
nand U1734 (N_1734,N_991,N_155);
and U1735 (N_1735,N_705,N_533);
nand U1736 (N_1736,N_486,N_852);
nor U1737 (N_1737,N_330,N_274);
or U1738 (N_1738,N_827,N_573);
and U1739 (N_1739,N_44,N_941);
nand U1740 (N_1740,N_803,N_788);
nor U1741 (N_1741,N_995,N_917);
nand U1742 (N_1742,N_444,N_114);
nor U1743 (N_1743,N_392,N_448);
nor U1744 (N_1744,N_766,N_689);
or U1745 (N_1745,N_866,N_266);
nor U1746 (N_1746,N_268,N_46);
and U1747 (N_1747,N_974,N_724);
nor U1748 (N_1748,N_267,N_467);
and U1749 (N_1749,N_984,N_950);
xnor U1750 (N_1750,N_675,N_293);
or U1751 (N_1751,N_325,N_890);
nand U1752 (N_1752,N_947,N_878);
and U1753 (N_1753,N_850,N_722);
or U1754 (N_1754,N_503,N_524);
nor U1755 (N_1755,N_602,N_644);
and U1756 (N_1756,N_453,N_265);
or U1757 (N_1757,N_559,N_521);
nand U1758 (N_1758,N_384,N_54);
nor U1759 (N_1759,N_370,N_653);
nor U1760 (N_1760,N_42,N_365);
or U1761 (N_1761,N_589,N_989);
nand U1762 (N_1762,N_881,N_516);
nand U1763 (N_1763,N_211,N_325);
or U1764 (N_1764,N_190,N_890);
nor U1765 (N_1765,N_547,N_119);
nand U1766 (N_1766,N_19,N_984);
nor U1767 (N_1767,N_828,N_402);
or U1768 (N_1768,N_306,N_662);
nor U1769 (N_1769,N_137,N_314);
or U1770 (N_1770,N_29,N_11);
nand U1771 (N_1771,N_821,N_772);
nand U1772 (N_1772,N_536,N_992);
nand U1773 (N_1773,N_675,N_193);
or U1774 (N_1774,N_917,N_395);
or U1775 (N_1775,N_163,N_46);
or U1776 (N_1776,N_87,N_698);
xnor U1777 (N_1777,N_249,N_897);
and U1778 (N_1778,N_529,N_392);
and U1779 (N_1779,N_522,N_741);
or U1780 (N_1780,N_749,N_746);
nor U1781 (N_1781,N_404,N_273);
and U1782 (N_1782,N_373,N_339);
nor U1783 (N_1783,N_312,N_552);
nand U1784 (N_1784,N_9,N_648);
or U1785 (N_1785,N_423,N_217);
nor U1786 (N_1786,N_892,N_417);
nand U1787 (N_1787,N_788,N_658);
nand U1788 (N_1788,N_359,N_200);
nor U1789 (N_1789,N_244,N_418);
and U1790 (N_1790,N_485,N_924);
or U1791 (N_1791,N_148,N_363);
nand U1792 (N_1792,N_399,N_522);
or U1793 (N_1793,N_642,N_674);
or U1794 (N_1794,N_191,N_416);
nand U1795 (N_1795,N_204,N_323);
nor U1796 (N_1796,N_349,N_570);
and U1797 (N_1797,N_962,N_767);
or U1798 (N_1798,N_361,N_342);
nand U1799 (N_1799,N_167,N_666);
or U1800 (N_1800,N_900,N_107);
nor U1801 (N_1801,N_487,N_171);
nor U1802 (N_1802,N_88,N_535);
nand U1803 (N_1803,N_428,N_19);
or U1804 (N_1804,N_256,N_129);
and U1805 (N_1805,N_12,N_332);
and U1806 (N_1806,N_966,N_392);
nor U1807 (N_1807,N_352,N_250);
or U1808 (N_1808,N_43,N_742);
and U1809 (N_1809,N_420,N_487);
and U1810 (N_1810,N_595,N_111);
nand U1811 (N_1811,N_594,N_60);
and U1812 (N_1812,N_575,N_797);
nand U1813 (N_1813,N_291,N_882);
nor U1814 (N_1814,N_943,N_603);
and U1815 (N_1815,N_952,N_30);
and U1816 (N_1816,N_735,N_321);
nor U1817 (N_1817,N_190,N_975);
and U1818 (N_1818,N_523,N_378);
and U1819 (N_1819,N_863,N_381);
or U1820 (N_1820,N_580,N_604);
nor U1821 (N_1821,N_939,N_342);
or U1822 (N_1822,N_361,N_100);
nor U1823 (N_1823,N_433,N_77);
and U1824 (N_1824,N_465,N_939);
nand U1825 (N_1825,N_589,N_906);
and U1826 (N_1826,N_595,N_309);
and U1827 (N_1827,N_247,N_125);
and U1828 (N_1828,N_869,N_403);
nor U1829 (N_1829,N_906,N_644);
nand U1830 (N_1830,N_717,N_393);
nor U1831 (N_1831,N_232,N_915);
or U1832 (N_1832,N_397,N_946);
or U1833 (N_1833,N_54,N_482);
and U1834 (N_1834,N_18,N_683);
xnor U1835 (N_1835,N_449,N_984);
and U1836 (N_1836,N_162,N_841);
nor U1837 (N_1837,N_397,N_145);
or U1838 (N_1838,N_997,N_609);
nor U1839 (N_1839,N_501,N_603);
and U1840 (N_1840,N_218,N_931);
and U1841 (N_1841,N_941,N_965);
nor U1842 (N_1842,N_127,N_720);
nand U1843 (N_1843,N_467,N_501);
and U1844 (N_1844,N_466,N_322);
nor U1845 (N_1845,N_173,N_402);
nand U1846 (N_1846,N_414,N_747);
and U1847 (N_1847,N_921,N_976);
and U1848 (N_1848,N_244,N_793);
or U1849 (N_1849,N_27,N_747);
nand U1850 (N_1850,N_304,N_387);
or U1851 (N_1851,N_670,N_997);
and U1852 (N_1852,N_760,N_241);
or U1853 (N_1853,N_982,N_189);
nand U1854 (N_1854,N_199,N_75);
or U1855 (N_1855,N_557,N_72);
nor U1856 (N_1856,N_28,N_450);
nand U1857 (N_1857,N_536,N_851);
nand U1858 (N_1858,N_548,N_912);
and U1859 (N_1859,N_679,N_361);
and U1860 (N_1860,N_437,N_939);
or U1861 (N_1861,N_156,N_490);
nand U1862 (N_1862,N_871,N_154);
and U1863 (N_1863,N_939,N_859);
nor U1864 (N_1864,N_140,N_133);
or U1865 (N_1865,N_460,N_586);
or U1866 (N_1866,N_915,N_198);
or U1867 (N_1867,N_321,N_527);
and U1868 (N_1868,N_411,N_41);
and U1869 (N_1869,N_305,N_508);
and U1870 (N_1870,N_51,N_90);
or U1871 (N_1871,N_723,N_532);
and U1872 (N_1872,N_856,N_954);
nor U1873 (N_1873,N_268,N_270);
or U1874 (N_1874,N_482,N_440);
or U1875 (N_1875,N_32,N_397);
xnor U1876 (N_1876,N_85,N_136);
or U1877 (N_1877,N_510,N_132);
nor U1878 (N_1878,N_852,N_706);
and U1879 (N_1879,N_885,N_193);
or U1880 (N_1880,N_417,N_845);
nand U1881 (N_1881,N_114,N_888);
or U1882 (N_1882,N_718,N_74);
nand U1883 (N_1883,N_618,N_898);
nor U1884 (N_1884,N_205,N_74);
nor U1885 (N_1885,N_12,N_840);
or U1886 (N_1886,N_338,N_887);
nor U1887 (N_1887,N_68,N_690);
and U1888 (N_1888,N_345,N_114);
nand U1889 (N_1889,N_356,N_652);
and U1890 (N_1890,N_167,N_813);
and U1891 (N_1891,N_973,N_481);
or U1892 (N_1892,N_990,N_37);
and U1893 (N_1893,N_144,N_14);
nand U1894 (N_1894,N_34,N_372);
and U1895 (N_1895,N_38,N_183);
nand U1896 (N_1896,N_462,N_493);
and U1897 (N_1897,N_101,N_864);
or U1898 (N_1898,N_933,N_17);
nor U1899 (N_1899,N_65,N_145);
nand U1900 (N_1900,N_157,N_758);
and U1901 (N_1901,N_365,N_993);
or U1902 (N_1902,N_827,N_919);
and U1903 (N_1903,N_17,N_214);
nand U1904 (N_1904,N_406,N_795);
and U1905 (N_1905,N_583,N_15);
nor U1906 (N_1906,N_865,N_836);
or U1907 (N_1907,N_551,N_584);
or U1908 (N_1908,N_344,N_278);
or U1909 (N_1909,N_851,N_885);
nor U1910 (N_1910,N_805,N_344);
or U1911 (N_1911,N_441,N_124);
nor U1912 (N_1912,N_621,N_626);
nand U1913 (N_1913,N_840,N_20);
or U1914 (N_1914,N_700,N_230);
and U1915 (N_1915,N_672,N_674);
and U1916 (N_1916,N_77,N_156);
nand U1917 (N_1917,N_330,N_291);
and U1918 (N_1918,N_795,N_847);
nand U1919 (N_1919,N_963,N_200);
and U1920 (N_1920,N_46,N_951);
nor U1921 (N_1921,N_684,N_303);
nor U1922 (N_1922,N_91,N_499);
or U1923 (N_1923,N_628,N_92);
and U1924 (N_1924,N_320,N_243);
and U1925 (N_1925,N_472,N_84);
or U1926 (N_1926,N_430,N_844);
or U1927 (N_1927,N_972,N_625);
nor U1928 (N_1928,N_780,N_651);
and U1929 (N_1929,N_675,N_510);
nand U1930 (N_1930,N_349,N_266);
or U1931 (N_1931,N_867,N_544);
nand U1932 (N_1932,N_437,N_483);
nand U1933 (N_1933,N_651,N_87);
nor U1934 (N_1934,N_811,N_2);
nand U1935 (N_1935,N_295,N_643);
nand U1936 (N_1936,N_267,N_950);
and U1937 (N_1937,N_434,N_32);
nand U1938 (N_1938,N_142,N_717);
and U1939 (N_1939,N_695,N_963);
nand U1940 (N_1940,N_156,N_439);
or U1941 (N_1941,N_382,N_472);
and U1942 (N_1942,N_574,N_343);
nand U1943 (N_1943,N_295,N_571);
nand U1944 (N_1944,N_657,N_675);
or U1945 (N_1945,N_200,N_669);
and U1946 (N_1946,N_28,N_729);
nor U1947 (N_1947,N_765,N_336);
nor U1948 (N_1948,N_102,N_220);
nor U1949 (N_1949,N_732,N_638);
and U1950 (N_1950,N_304,N_271);
or U1951 (N_1951,N_164,N_611);
and U1952 (N_1952,N_963,N_499);
or U1953 (N_1953,N_830,N_489);
nand U1954 (N_1954,N_452,N_620);
nand U1955 (N_1955,N_374,N_638);
and U1956 (N_1956,N_808,N_978);
nand U1957 (N_1957,N_8,N_66);
and U1958 (N_1958,N_468,N_67);
nor U1959 (N_1959,N_779,N_240);
or U1960 (N_1960,N_503,N_730);
and U1961 (N_1961,N_934,N_95);
nand U1962 (N_1962,N_958,N_441);
nand U1963 (N_1963,N_520,N_688);
nand U1964 (N_1964,N_544,N_31);
or U1965 (N_1965,N_886,N_221);
nor U1966 (N_1966,N_744,N_106);
nor U1967 (N_1967,N_499,N_202);
or U1968 (N_1968,N_851,N_813);
nor U1969 (N_1969,N_303,N_152);
and U1970 (N_1970,N_943,N_829);
and U1971 (N_1971,N_869,N_988);
and U1972 (N_1972,N_194,N_762);
nor U1973 (N_1973,N_926,N_460);
and U1974 (N_1974,N_659,N_618);
nand U1975 (N_1975,N_408,N_373);
and U1976 (N_1976,N_952,N_764);
or U1977 (N_1977,N_550,N_733);
or U1978 (N_1978,N_677,N_946);
nand U1979 (N_1979,N_460,N_117);
nor U1980 (N_1980,N_107,N_569);
nand U1981 (N_1981,N_707,N_273);
xnor U1982 (N_1982,N_344,N_886);
nand U1983 (N_1983,N_682,N_582);
or U1984 (N_1984,N_810,N_172);
nand U1985 (N_1985,N_378,N_652);
nor U1986 (N_1986,N_140,N_34);
nand U1987 (N_1987,N_456,N_218);
nand U1988 (N_1988,N_853,N_500);
nor U1989 (N_1989,N_774,N_975);
and U1990 (N_1990,N_395,N_508);
nor U1991 (N_1991,N_411,N_935);
nor U1992 (N_1992,N_308,N_728);
nand U1993 (N_1993,N_534,N_555);
and U1994 (N_1994,N_506,N_403);
nand U1995 (N_1995,N_789,N_154);
nand U1996 (N_1996,N_12,N_733);
nor U1997 (N_1997,N_140,N_449);
and U1998 (N_1998,N_496,N_466);
nor U1999 (N_1999,N_127,N_200);
or U2000 (N_2000,N_1592,N_1316);
nor U2001 (N_2001,N_1270,N_1852);
nor U2002 (N_2002,N_1729,N_1082);
or U2003 (N_2003,N_1177,N_1692);
nor U2004 (N_2004,N_1336,N_1639);
nor U2005 (N_2005,N_1241,N_1805);
nand U2006 (N_2006,N_1333,N_1123);
nand U2007 (N_2007,N_1772,N_1754);
or U2008 (N_2008,N_1344,N_1731);
nand U2009 (N_2009,N_1637,N_1682);
nand U2010 (N_2010,N_1785,N_1866);
nand U2011 (N_2011,N_1480,N_1933);
and U2012 (N_2012,N_1432,N_1341);
or U2013 (N_2013,N_1571,N_1519);
nand U2014 (N_2014,N_1018,N_1569);
nor U2015 (N_2015,N_1271,N_1445);
nand U2016 (N_2016,N_1141,N_1752);
or U2017 (N_2017,N_1273,N_1513);
and U2018 (N_2018,N_1358,N_1980);
nand U2019 (N_2019,N_1599,N_1088);
nand U2020 (N_2020,N_1957,N_1433);
nor U2021 (N_2021,N_1118,N_1414);
nand U2022 (N_2022,N_1281,N_1412);
or U2023 (N_2023,N_1265,N_1258);
nand U2024 (N_2024,N_1342,N_1434);
and U2025 (N_2025,N_1105,N_1911);
nor U2026 (N_2026,N_1255,N_1121);
nand U2027 (N_2027,N_1978,N_1797);
nand U2028 (N_2028,N_1961,N_1328);
and U2029 (N_2029,N_1645,N_1487);
and U2030 (N_2030,N_1556,N_1643);
or U2031 (N_2031,N_1824,N_1831);
nor U2032 (N_2032,N_1009,N_1074);
and U2033 (N_2033,N_1767,N_1810);
or U2034 (N_2034,N_1232,N_1804);
and U2035 (N_2035,N_1077,N_1894);
nand U2036 (N_2036,N_1944,N_1520);
nor U2037 (N_2037,N_1872,N_1460);
and U2038 (N_2038,N_1275,N_1129);
nor U2039 (N_2039,N_1180,N_1380);
or U2040 (N_2040,N_1788,N_1163);
and U2041 (N_2041,N_1753,N_1646);
and U2042 (N_2042,N_1026,N_1264);
and U2043 (N_2043,N_1755,N_1337);
nand U2044 (N_2044,N_1638,N_1188);
and U2045 (N_2045,N_1392,N_1442);
nor U2046 (N_2046,N_1763,N_1013);
nor U2047 (N_2047,N_1710,N_1798);
nand U2048 (N_2048,N_1555,N_1137);
nand U2049 (N_2049,N_1268,N_1076);
nor U2050 (N_2050,N_1959,N_1929);
nor U2051 (N_2051,N_1529,N_1078);
nand U2052 (N_2052,N_1476,N_1318);
nand U2053 (N_2053,N_1486,N_1998);
nand U2054 (N_2054,N_1764,N_1701);
and U2055 (N_2055,N_1693,N_1651);
nor U2056 (N_2056,N_1135,N_1041);
nor U2057 (N_2057,N_1491,N_1463);
or U2058 (N_2058,N_1923,N_1936);
nand U2059 (N_2059,N_1377,N_1705);
nand U2060 (N_2060,N_1097,N_1222);
nor U2061 (N_2061,N_1361,N_1372);
nand U2062 (N_2062,N_1406,N_1808);
nand U2063 (N_2063,N_1374,N_1606);
nand U2064 (N_2064,N_1469,N_1544);
nor U2065 (N_2065,N_1649,N_1090);
nand U2066 (N_2066,N_1526,N_1005);
xnor U2067 (N_2067,N_1220,N_1614);
nor U2068 (N_2068,N_1548,N_1941);
nand U2069 (N_2069,N_1827,N_1715);
nor U2070 (N_2070,N_1849,N_1300);
nand U2071 (N_2071,N_1427,N_1218);
nor U2072 (N_2072,N_1535,N_1898);
nand U2073 (N_2073,N_1350,N_1716);
nor U2074 (N_2074,N_1181,N_1679);
or U2075 (N_2075,N_1627,N_1540);
nand U2076 (N_2076,N_1055,N_1033);
nand U2077 (N_2077,N_1545,N_1794);
nor U2078 (N_2078,N_1738,N_1830);
and U2079 (N_2079,N_1413,N_1884);
or U2080 (N_2080,N_1751,N_1956);
or U2081 (N_2081,N_1305,N_1900);
and U2082 (N_2082,N_1518,N_1801);
nand U2083 (N_2083,N_1471,N_1550);
nand U2084 (N_2084,N_1883,N_1367);
or U2085 (N_2085,N_1613,N_1559);
nor U2086 (N_2086,N_1838,N_1766);
and U2087 (N_2087,N_1708,N_1388);
nand U2088 (N_2088,N_1932,N_1667);
or U2089 (N_2089,N_1176,N_1850);
nand U2090 (N_2090,N_1573,N_1977);
or U2091 (N_2091,N_1408,N_1813);
nor U2092 (N_2092,N_1953,N_1577);
or U2093 (N_2093,N_1290,N_1768);
nand U2094 (N_2094,N_1511,N_1481);
or U2095 (N_2095,N_1819,N_1095);
or U2096 (N_2096,N_1016,N_1672);
or U2097 (N_2097,N_1418,N_1765);
and U2098 (N_2098,N_1058,N_1100);
nor U2099 (N_2099,N_1946,N_1285);
nor U2100 (N_2100,N_1669,N_1029);
and U2101 (N_2101,N_1871,N_1541);
nor U2102 (N_2102,N_1175,N_1096);
xnor U2103 (N_2103,N_1576,N_1620);
and U2104 (N_2104,N_1484,N_1722);
or U2105 (N_2105,N_1046,N_1862);
and U2106 (N_2106,N_1204,N_1227);
nor U2107 (N_2107,N_1161,N_1942);
and U2108 (N_2108,N_1308,N_1157);
and U2109 (N_2109,N_1869,N_1295);
nor U2110 (N_2110,N_1549,N_1776);
nand U2111 (N_2111,N_1634,N_1391);
or U2112 (N_2112,N_1725,N_1587);
nor U2113 (N_2113,N_1488,N_1183);
nand U2114 (N_2114,N_1791,N_1254);
and U2115 (N_2115,N_1023,N_1379);
nor U2116 (N_2116,N_1186,N_1820);
nor U2117 (N_2117,N_1602,N_1122);
nand U2118 (N_2118,N_1952,N_1636);
or U2119 (N_2119,N_1043,N_1119);
nand U2120 (N_2120,N_1990,N_1190);
or U2121 (N_2121,N_1037,N_1728);
nand U2122 (N_2122,N_1818,N_1260);
nor U2123 (N_2123,N_1653,N_1604);
nand U2124 (N_2124,N_1162,N_1330);
or U2125 (N_2125,N_1187,N_1600);
nand U2126 (N_2126,N_1086,N_1796);
nor U2127 (N_2127,N_1732,N_1992);
nand U2128 (N_2128,N_1371,N_1044);
nand U2129 (N_2129,N_1893,N_1447);
or U2130 (N_2130,N_1938,N_1853);
nand U2131 (N_2131,N_1761,N_1995);
and U2132 (N_2132,N_1702,N_1904);
and U2133 (N_2133,N_1383,N_1173);
nor U2134 (N_2134,N_1861,N_1746);
nor U2135 (N_2135,N_1973,N_1823);
and U2136 (N_2136,N_1498,N_1574);
nand U2137 (N_2137,N_1283,N_1685);
nand U2138 (N_2138,N_1654,N_1865);
nand U2139 (N_2139,N_1207,N_1527);
nor U2140 (N_2140,N_1880,N_1661);
nand U2141 (N_2141,N_1224,N_1249);
and U2142 (N_2142,N_1138,N_1735);
nor U2143 (N_2143,N_1323,N_1863);
and U2144 (N_2144,N_1053,N_1324);
and U2145 (N_2145,N_1897,N_1102);
nor U2146 (N_2146,N_1069,N_1931);
and U2147 (N_2147,N_1322,N_1558);
and U2148 (N_2148,N_1899,N_1854);
or U2149 (N_2149,N_1107,N_1168);
nor U2150 (N_2150,N_1782,N_1212);
nand U2151 (N_2151,N_1398,N_1635);
nor U2152 (N_2152,N_1325,N_1816);
nand U2153 (N_2153,N_1083,N_1451);
or U2154 (N_2154,N_1809,N_1561);
nand U2155 (N_2155,N_1934,N_1595);
nand U2156 (N_2156,N_1126,N_1142);
or U2157 (N_2157,N_1233,N_1726);
nor U2158 (N_2158,N_1700,N_1879);
nand U2159 (N_2159,N_1937,N_1309);
and U2160 (N_2160,N_1048,N_1652);
nor U2161 (N_2161,N_1890,N_1094);
nor U2162 (N_2162,N_1826,N_1237);
and U2163 (N_2163,N_1658,N_1662);
or U2164 (N_2164,N_1152,N_1125);
nand U2165 (N_2165,N_1557,N_1533);
nand U2166 (N_2166,N_1274,N_1777);
or U2167 (N_2167,N_1873,N_1428);
nor U2168 (N_2168,N_1339,N_1165);
nand U2169 (N_2169,N_1628,N_1775);
and U2170 (N_2170,N_1140,N_1566);
nor U2171 (N_2171,N_1762,N_1607);
nor U2172 (N_2172,N_1200,N_1150);
nor U2173 (N_2173,N_1349,N_1874);
nand U2174 (N_2174,N_1008,N_1231);
or U2175 (N_2175,N_1892,N_1881);
nand U2176 (N_2176,N_1317,N_1219);
or U2177 (N_2177,N_1441,N_1038);
nor U2178 (N_2178,N_1151,N_1128);
nor U2179 (N_2179,N_1909,N_1523);
or U2180 (N_2180,N_1686,N_1981);
or U2181 (N_2181,N_1279,N_1192);
nor U2182 (N_2182,N_1331,N_1800);
nor U2183 (N_2183,N_1594,N_1477);
nor U2184 (N_2184,N_1745,N_1774);
nand U2185 (N_2185,N_1506,N_1012);
nand U2186 (N_2186,N_1538,N_1542);
and U2187 (N_2187,N_1582,N_1292);
nand U2188 (N_2188,N_1568,N_1783);
nand U2189 (N_2189,N_1299,N_1773);
and U2190 (N_2190,N_1311,N_1502);
and U2191 (N_2191,N_1665,N_1531);
and U2192 (N_2192,N_1457,N_1036);
nor U2193 (N_2193,N_1389,N_1920);
nand U2194 (N_2194,N_1734,N_1202);
or U2195 (N_2195,N_1886,N_1962);
or U2196 (N_2196,N_1963,N_1707);
or U2197 (N_2197,N_1532,N_1688);
nor U2198 (N_2198,N_1515,N_1760);
nand U2199 (N_2199,N_1727,N_1357);
and U2200 (N_2200,N_1655,N_1583);
nor U2201 (N_2201,N_1049,N_1698);
nor U2202 (N_2202,N_1875,N_1440);
and U2203 (N_2203,N_1603,N_1756);
nand U2204 (N_2204,N_1297,N_1116);
and U2205 (N_2205,N_1354,N_1803);
or U2206 (N_2206,N_1958,N_1737);
and U2207 (N_2207,N_1117,N_1028);
or U2208 (N_2208,N_1790,N_1355);
or U2209 (N_2209,N_1251,N_1997);
or U2210 (N_2210,N_1034,N_1799);
nor U2211 (N_2211,N_1972,N_1924);
and U2212 (N_2212,N_1509,N_1402);
and U2213 (N_2213,N_1877,N_1411);
nand U2214 (N_2214,N_1927,N_1741);
and U2215 (N_2215,N_1326,N_1492);
nor U2216 (N_2216,N_1905,N_1362);
nor U2217 (N_2217,N_1743,N_1489);
nand U2218 (N_2218,N_1882,N_1091);
nand U2219 (N_2219,N_1784,N_1841);
nand U2220 (N_2220,N_1148,N_1598);
or U2221 (N_2221,N_1832,N_1468);
nor U2222 (N_2222,N_1517,N_1626);
or U2223 (N_2223,N_1787,N_1429);
or U2224 (N_2224,N_1421,N_1209);
nor U2225 (N_2225,N_1430,N_1424);
or U2226 (N_2226,N_1618,N_1199);
or U2227 (N_2227,N_1610,N_1178);
nand U2228 (N_2228,N_1294,N_1913);
nor U2229 (N_2229,N_1591,N_1581);
nor U2230 (N_2230,N_1416,N_1621);
or U2231 (N_2231,N_1185,N_1153);
nand U2232 (N_2232,N_1236,N_1828);
and U2233 (N_2233,N_1111,N_1706);
and U2234 (N_2234,N_1969,N_1431);
xnor U2235 (N_2235,N_1844,N_1387);
and U2236 (N_2236,N_1678,N_1683);
and U2237 (N_2237,N_1666,N_1807);
and U2238 (N_2238,N_1612,N_1196);
or U2239 (N_2239,N_1608,N_1359);
or U2240 (N_2240,N_1001,N_1245);
nand U2241 (N_2241,N_1822,N_1530);
or U2242 (N_2242,N_1553,N_1101);
nor U2243 (N_2243,N_1771,N_1843);
and U2244 (N_2244,N_1885,N_1059);
nand U2245 (N_2245,N_1006,N_1588);
and U2246 (N_2246,N_1966,N_1779);
nand U2247 (N_2247,N_1758,N_1572);
nand U2248 (N_2248,N_1906,N_1315);
or U2249 (N_2249,N_1465,N_1132);
or U2250 (N_2250,N_1960,N_1466);
nor U2251 (N_2251,N_1982,N_1160);
and U2252 (N_2252,N_1250,N_1159);
nor U2253 (N_2253,N_1373,N_1903);
and U2254 (N_2254,N_1288,N_1017);
nor U2255 (N_2255,N_1313,N_1475);
nand U2256 (N_2256,N_1914,N_1439);
and U2257 (N_2257,N_1409,N_1052);
nor U2258 (N_2258,N_1855,N_1605);
and U2259 (N_2259,N_1719,N_1000);
or U2260 (N_2260,N_1410,N_1695);
or U2261 (N_2261,N_1239,N_1143);
nand U2262 (N_2262,N_1631,N_1689);
or U2263 (N_2263,N_1586,N_1022);
or U2264 (N_2264,N_1659,N_1443);
xor U2265 (N_2265,N_1723,N_1497);
or U2266 (N_2266,N_1174,N_1390);
and U2267 (N_2267,N_1448,N_1127);
nand U2268 (N_2268,N_1951,N_1584);
and U2269 (N_2269,N_1343,N_1993);
or U2270 (N_2270,N_1216,N_1114);
nor U2271 (N_2271,N_1590,N_1145);
or U2272 (N_2272,N_1108,N_1435);
and U2273 (N_2273,N_1184,N_1266);
nand U2274 (N_2274,N_1170,N_1240);
or U2275 (N_2275,N_1347,N_1919);
nor U2276 (N_2276,N_1182,N_1625);
or U2277 (N_2277,N_1110,N_1611);
nor U2278 (N_2278,N_1139,N_1986);
or U2279 (N_2279,N_1539,N_1149);
nor U2280 (N_2280,N_1304,N_1045);
nand U2281 (N_2281,N_1935,N_1656);
and U2282 (N_2282,N_1563,N_1479);
nand U2283 (N_2283,N_1696,N_1422);
or U2284 (N_2284,N_1622,N_1505);
or U2285 (N_2285,N_1856,N_1467);
nor U2286 (N_2286,N_1994,N_1019);
nand U2287 (N_2287,N_1267,N_1071);
nor U2288 (N_2288,N_1385,N_1320);
or U2289 (N_2289,N_1747,N_1848);
nor U2290 (N_2290,N_1641,N_1195);
xor U2291 (N_2291,N_1269,N_1930);
and U2292 (N_2292,N_1965,N_1057);
or U2293 (N_2293,N_1718,N_1133);
and U2294 (N_2294,N_1438,N_1353);
and U2295 (N_2295,N_1314,N_1039);
nor U2296 (N_2296,N_1205,N_1675);
nor U2297 (N_2297,N_1282,N_1147);
or U2298 (N_2298,N_1449,N_1172);
and U2299 (N_2299,N_1499,N_1534);
or U2300 (N_2300,N_1321,N_1375);
or U2301 (N_2301,N_1522,N_1042);
xnor U2302 (N_2302,N_1870,N_1221);
nor U2303 (N_2303,N_1901,N_1400);
or U2304 (N_2304,N_1235,N_1368);
and U2305 (N_2305,N_1947,N_1979);
and U2306 (N_2306,N_1405,N_1851);
and U2307 (N_2307,N_1419,N_1464);
nor U2308 (N_2308,N_1201,N_1436);
or U2309 (N_2309,N_1717,N_1002);
or U2310 (N_2310,N_1423,N_1455);
nor U2311 (N_2311,N_1462,N_1617);
nor U2312 (N_2312,N_1842,N_1397);
nand U2313 (N_2313,N_1940,N_1242);
nor U2314 (N_2314,N_1054,N_1007);
or U2315 (N_2315,N_1954,N_1806);
or U2316 (N_2316,N_1793,N_1724);
xnor U2317 (N_2317,N_1364,N_1365);
and U2318 (N_2318,N_1570,N_1167);
or U2319 (N_2319,N_1889,N_1130);
and U2320 (N_2320,N_1112,N_1454);
and U2321 (N_2321,N_1061,N_1757);
nor U2322 (N_2322,N_1648,N_1814);
nor U2323 (N_2323,N_1291,N_1742);
and U2324 (N_2324,N_1303,N_1472);
and U2325 (N_2325,N_1276,N_1459);
nor U2326 (N_2326,N_1370,N_1524);
nand U2327 (N_2327,N_1781,N_1453);
and U2328 (N_2328,N_1261,N_1704);
and U2329 (N_2329,N_1458,N_1327);
nor U2330 (N_2330,N_1335,N_1507);
nand U2331 (N_2331,N_1099,N_1922);
and U2332 (N_2332,N_1081,N_1759);
nand U2333 (N_2333,N_1684,N_1407);
nand U2334 (N_2334,N_1399,N_1021);
nor U2335 (N_2335,N_1902,N_1712);
and U2336 (N_2336,N_1115,N_1360);
or U2337 (N_2337,N_1068,N_1629);
or U2338 (N_2338,N_1835,N_1067);
and U2339 (N_2339,N_1144,N_1490);
nor U2340 (N_2340,N_1687,N_1596);
and U2341 (N_2341,N_1403,N_1287);
or U2342 (N_2342,N_1426,N_1918);
nand U2343 (N_2343,N_1503,N_1677);
or U2344 (N_2344,N_1340,N_1075);
nand U2345 (N_2345,N_1415,N_1720);
nand U2346 (N_2346,N_1896,N_1562);
nor U2347 (N_2347,N_1106,N_1286);
or U2348 (N_2348,N_1010,N_1949);
and U2349 (N_2349,N_1811,N_1644);
nand U2350 (N_2350,N_1615,N_1504);
and U2351 (N_2351,N_1496,N_1868);
and U2352 (N_2352,N_1730,N_1084);
nand U2353 (N_2353,N_1713,N_1395);
or U2354 (N_2354,N_1166,N_1836);
and U2355 (N_2355,N_1493,N_1450);
nand U2356 (N_2356,N_1396,N_1733);
nor U2357 (N_2357,N_1277,N_1660);
nand U2358 (N_2358,N_1296,N_1825);
or U2359 (N_2359,N_1833,N_1345);
or U2360 (N_2360,N_1051,N_1263);
nor U2361 (N_2361,N_1478,N_1351);
nor U2362 (N_2362,N_1280,N_1864);
and U2363 (N_2363,N_1070,N_1792);
or U2364 (N_2364,N_1674,N_1073);
nand U2365 (N_2365,N_1748,N_1146);
nand U2366 (N_2366,N_1714,N_1983);
nor U2367 (N_2367,N_1289,N_1035);
and U2368 (N_2368,N_1999,N_1366);
or U2369 (N_2369,N_1575,N_1846);
and U2370 (N_2370,N_1908,N_1821);
nand U2371 (N_2371,N_1376,N_1812);
and U2372 (N_2372,N_1027,N_1967);
and U2373 (N_2373,N_1516,N_1740);
nor U2374 (N_2374,N_1063,N_1134);
and U2375 (N_2375,N_1551,N_1749);
or U2376 (N_2376,N_1197,N_1786);
nand U2377 (N_2377,N_1939,N_1891);
or U2378 (N_2378,N_1352,N_1306);
nor U2379 (N_2379,N_1860,N_1925);
or U2380 (N_2380,N_1964,N_1943);
nand U2381 (N_2381,N_1624,N_1302);
nand U2382 (N_2382,N_1203,N_1062);
and U2383 (N_2383,N_1681,N_1837);
nand U2384 (N_2384,N_1680,N_1697);
nor U2385 (N_2385,N_1169,N_1543);
and U2386 (N_2386,N_1065,N_1156);
or U2387 (N_2387,N_1348,N_1064);
nand U2388 (N_2388,N_1120,N_1721);
or U2389 (N_2389,N_1470,N_1514);
nand U2390 (N_2390,N_1262,N_1014);
nor U2391 (N_2391,N_1580,N_1750);
nand U2392 (N_2392,N_1691,N_1597);
or U2393 (N_2393,N_1154,N_1298);
and U2394 (N_2394,N_1921,N_1632);
nor U2395 (N_2395,N_1092,N_1425);
and U2396 (N_2396,N_1198,N_1560);
or U2397 (N_2397,N_1089,N_1736);
nand U2398 (N_2398,N_1915,N_1378);
or U2399 (N_2399,N_1916,N_1546);
nor U2400 (N_2400,N_1694,N_1229);
nand U2401 (N_2401,N_1578,N_1401);
nand U2402 (N_2402,N_1031,N_1711);
nand U2403 (N_2403,N_1609,N_1647);
or U2404 (N_2404,N_1673,N_1194);
or U2405 (N_2405,N_1976,N_1971);
or U2406 (N_2406,N_1945,N_1437);
nor U2407 (N_2407,N_1179,N_1917);
and U2408 (N_2408,N_1579,N_1537);
or U2409 (N_2409,N_1839,N_1554);
nand U2410 (N_2410,N_1991,N_1223);
nor U2411 (N_2411,N_1124,N_1420);
nand U2412 (N_2412,N_1136,N_1093);
or U2413 (N_2413,N_1670,N_1225);
or U2414 (N_2414,N_1248,N_1552);
nand U2415 (N_2415,N_1601,N_1346);
nor U2416 (N_2416,N_1616,N_1802);
and U2417 (N_2417,N_1525,N_1912);
and U2418 (N_2418,N_1040,N_1955);
and U2419 (N_2419,N_1989,N_1113);
and U2420 (N_2420,N_1050,N_1907);
nor U2421 (N_2421,N_1080,N_1664);
nand U2422 (N_2422,N_1858,N_1393);
nor U2423 (N_2423,N_1334,N_1567);
xnor U2424 (N_2424,N_1501,N_1474);
and U2425 (N_2425,N_1386,N_1640);
or U2426 (N_2426,N_1536,N_1310);
or U2427 (N_2427,N_1657,N_1817);
nand U2428 (N_2428,N_1593,N_1384);
nand U2429 (N_2429,N_1623,N_1011);
nor U2430 (N_2430,N_1238,N_1020);
nor U2431 (N_2431,N_1417,N_1312);
and U2432 (N_2432,N_1508,N_1770);
xnor U2433 (N_2433,N_1996,N_1500);
or U2434 (N_2434,N_1452,N_1003);
nor U2435 (N_2435,N_1984,N_1214);
and U2436 (N_2436,N_1257,N_1158);
nand U2437 (N_2437,N_1404,N_1512);
nand U2438 (N_2438,N_1895,N_1676);
nor U2439 (N_2439,N_1030,N_1066);
nand U2440 (N_2440,N_1272,N_1564);
nor U2441 (N_2441,N_1987,N_1633);
and U2442 (N_2442,N_1363,N_1744);
nor U2443 (N_2443,N_1256,N_1193);
nand U2444 (N_2444,N_1619,N_1970);
xor U2445 (N_2445,N_1085,N_1495);
and U2446 (N_2446,N_1338,N_1381);
or U2447 (N_2447,N_1815,N_1985);
nor U2448 (N_2448,N_1098,N_1888);
and U2449 (N_2449,N_1876,N_1191);
nor U2450 (N_2450,N_1293,N_1259);
nor U2451 (N_2451,N_1630,N_1004);
nand U2452 (N_2452,N_1087,N_1456);
nor U2453 (N_2453,N_1473,N_1332);
nor U2454 (N_2454,N_1446,N_1585);
nand U2455 (N_2455,N_1510,N_1060);
nand U2456 (N_2456,N_1690,N_1703);
and U2457 (N_2457,N_1230,N_1301);
nand U2458 (N_2458,N_1857,N_1329);
and U2459 (N_2459,N_1278,N_1521);
xnor U2460 (N_2460,N_1988,N_1845);
or U2461 (N_2461,N_1968,N_1444);
nor U2462 (N_2462,N_1483,N_1974);
or U2463 (N_2463,N_1047,N_1211);
nor U2464 (N_2464,N_1829,N_1025);
nor U2465 (N_2465,N_1668,N_1015);
nor U2466 (N_2466,N_1024,N_1494);
nor U2467 (N_2467,N_1056,N_1709);
xnor U2468 (N_2468,N_1948,N_1032);
nand U2469 (N_2469,N_1834,N_1950);
nand U2470 (N_2470,N_1215,N_1975);
nand U2471 (N_2471,N_1840,N_1671);
or U2472 (N_2472,N_1482,N_1547);
and U2473 (N_2473,N_1589,N_1079);
and U2474 (N_2474,N_1650,N_1228);
nor U2475 (N_2475,N_1926,N_1663);
nand U2476 (N_2476,N_1565,N_1778);
nand U2477 (N_2477,N_1739,N_1528);
nand U2478 (N_2478,N_1307,N_1382);
or U2479 (N_2479,N_1104,N_1252);
or U2480 (N_2480,N_1642,N_1164);
nor U2481 (N_2481,N_1369,N_1356);
nor U2482 (N_2482,N_1244,N_1699);
or U2483 (N_2483,N_1072,N_1461);
and U2484 (N_2484,N_1847,N_1795);
nand U2485 (N_2485,N_1910,N_1319);
and U2486 (N_2486,N_1217,N_1394);
nand U2487 (N_2487,N_1171,N_1155);
nand U2488 (N_2488,N_1789,N_1887);
nand U2489 (N_2489,N_1103,N_1226);
or U2490 (N_2490,N_1780,N_1928);
nand U2491 (N_2491,N_1867,N_1246);
nor U2492 (N_2492,N_1253,N_1189);
nor U2493 (N_2493,N_1485,N_1769);
nor U2494 (N_2494,N_1131,N_1206);
nand U2495 (N_2495,N_1213,N_1210);
nor U2496 (N_2496,N_1109,N_1247);
or U2497 (N_2497,N_1859,N_1878);
or U2498 (N_2498,N_1208,N_1234);
nor U2499 (N_2499,N_1243,N_1284);
nand U2500 (N_2500,N_1832,N_1146);
or U2501 (N_2501,N_1201,N_1256);
nand U2502 (N_2502,N_1747,N_1757);
and U2503 (N_2503,N_1390,N_1568);
nand U2504 (N_2504,N_1301,N_1102);
and U2505 (N_2505,N_1835,N_1431);
nand U2506 (N_2506,N_1081,N_1414);
or U2507 (N_2507,N_1401,N_1005);
nor U2508 (N_2508,N_1279,N_1474);
and U2509 (N_2509,N_1681,N_1182);
and U2510 (N_2510,N_1785,N_1459);
nor U2511 (N_2511,N_1351,N_1071);
nor U2512 (N_2512,N_1915,N_1786);
nand U2513 (N_2513,N_1975,N_1029);
nor U2514 (N_2514,N_1371,N_1631);
nand U2515 (N_2515,N_1353,N_1952);
and U2516 (N_2516,N_1919,N_1689);
or U2517 (N_2517,N_1516,N_1769);
and U2518 (N_2518,N_1875,N_1599);
nor U2519 (N_2519,N_1135,N_1911);
nor U2520 (N_2520,N_1286,N_1019);
nand U2521 (N_2521,N_1619,N_1403);
or U2522 (N_2522,N_1145,N_1951);
and U2523 (N_2523,N_1106,N_1702);
or U2524 (N_2524,N_1170,N_1289);
nand U2525 (N_2525,N_1006,N_1446);
or U2526 (N_2526,N_1052,N_1847);
nor U2527 (N_2527,N_1597,N_1056);
and U2528 (N_2528,N_1781,N_1677);
nand U2529 (N_2529,N_1976,N_1514);
nand U2530 (N_2530,N_1712,N_1267);
or U2531 (N_2531,N_1097,N_1163);
nor U2532 (N_2532,N_1551,N_1414);
or U2533 (N_2533,N_1931,N_1963);
nand U2534 (N_2534,N_1197,N_1896);
nand U2535 (N_2535,N_1178,N_1908);
nand U2536 (N_2536,N_1448,N_1830);
and U2537 (N_2537,N_1839,N_1965);
nand U2538 (N_2538,N_1900,N_1259);
nor U2539 (N_2539,N_1469,N_1178);
and U2540 (N_2540,N_1787,N_1440);
nor U2541 (N_2541,N_1070,N_1794);
and U2542 (N_2542,N_1086,N_1724);
or U2543 (N_2543,N_1875,N_1015);
nand U2544 (N_2544,N_1535,N_1360);
nand U2545 (N_2545,N_1413,N_1080);
nor U2546 (N_2546,N_1778,N_1780);
and U2547 (N_2547,N_1936,N_1805);
or U2548 (N_2548,N_1153,N_1080);
nand U2549 (N_2549,N_1389,N_1751);
and U2550 (N_2550,N_1309,N_1298);
nor U2551 (N_2551,N_1275,N_1998);
nor U2552 (N_2552,N_1345,N_1052);
and U2553 (N_2553,N_1556,N_1086);
nand U2554 (N_2554,N_1589,N_1275);
or U2555 (N_2555,N_1928,N_1381);
nor U2556 (N_2556,N_1037,N_1223);
nor U2557 (N_2557,N_1086,N_1243);
nor U2558 (N_2558,N_1806,N_1363);
or U2559 (N_2559,N_1554,N_1043);
nand U2560 (N_2560,N_1310,N_1847);
or U2561 (N_2561,N_1973,N_1472);
nand U2562 (N_2562,N_1196,N_1509);
nand U2563 (N_2563,N_1782,N_1600);
nand U2564 (N_2564,N_1944,N_1743);
nor U2565 (N_2565,N_1710,N_1951);
and U2566 (N_2566,N_1624,N_1580);
nand U2567 (N_2567,N_1211,N_1668);
or U2568 (N_2568,N_1247,N_1736);
and U2569 (N_2569,N_1549,N_1860);
nand U2570 (N_2570,N_1738,N_1674);
nand U2571 (N_2571,N_1808,N_1215);
nor U2572 (N_2572,N_1191,N_1866);
and U2573 (N_2573,N_1057,N_1851);
or U2574 (N_2574,N_1406,N_1697);
nor U2575 (N_2575,N_1996,N_1169);
and U2576 (N_2576,N_1120,N_1516);
or U2577 (N_2577,N_1904,N_1569);
nor U2578 (N_2578,N_1223,N_1259);
or U2579 (N_2579,N_1177,N_1536);
and U2580 (N_2580,N_1342,N_1523);
nand U2581 (N_2581,N_1498,N_1476);
and U2582 (N_2582,N_1219,N_1090);
nand U2583 (N_2583,N_1366,N_1598);
or U2584 (N_2584,N_1616,N_1727);
and U2585 (N_2585,N_1430,N_1226);
nor U2586 (N_2586,N_1037,N_1518);
nand U2587 (N_2587,N_1359,N_1703);
nor U2588 (N_2588,N_1885,N_1442);
or U2589 (N_2589,N_1415,N_1075);
or U2590 (N_2590,N_1148,N_1089);
or U2591 (N_2591,N_1249,N_1443);
or U2592 (N_2592,N_1018,N_1559);
nor U2593 (N_2593,N_1255,N_1508);
nand U2594 (N_2594,N_1415,N_1691);
or U2595 (N_2595,N_1709,N_1974);
nand U2596 (N_2596,N_1336,N_1591);
and U2597 (N_2597,N_1112,N_1563);
or U2598 (N_2598,N_1101,N_1026);
nor U2599 (N_2599,N_1172,N_1758);
or U2600 (N_2600,N_1892,N_1724);
and U2601 (N_2601,N_1850,N_1225);
nand U2602 (N_2602,N_1178,N_1948);
nor U2603 (N_2603,N_1471,N_1776);
or U2604 (N_2604,N_1672,N_1634);
or U2605 (N_2605,N_1753,N_1290);
and U2606 (N_2606,N_1377,N_1511);
nor U2607 (N_2607,N_1175,N_1232);
or U2608 (N_2608,N_1946,N_1995);
nor U2609 (N_2609,N_1714,N_1523);
and U2610 (N_2610,N_1584,N_1560);
nand U2611 (N_2611,N_1842,N_1101);
and U2612 (N_2612,N_1286,N_1039);
nand U2613 (N_2613,N_1154,N_1753);
and U2614 (N_2614,N_1564,N_1638);
and U2615 (N_2615,N_1895,N_1168);
nand U2616 (N_2616,N_1497,N_1180);
nor U2617 (N_2617,N_1408,N_1687);
xor U2618 (N_2618,N_1471,N_1323);
or U2619 (N_2619,N_1324,N_1168);
or U2620 (N_2620,N_1979,N_1724);
nor U2621 (N_2621,N_1790,N_1789);
or U2622 (N_2622,N_1032,N_1353);
and U2623 (N_2623,N_1055,N_1724);
nand U2624 (N_2624,N_1176,N_1087);
nor U2625 (N_2625,N_1814,N_1255);
and U2626 (N_2626,N_1590,N_1351);
nor U2627 (N_2627,N_1523,N_1429);
or U2628 (N_2628,N_1517,N_1858);
nand U2629 (N_2629,N_1818,N_1573);
or U2630 (N_2630,N_1827,N_1738);
nor U2631 (N_2631,N_1898,N_1808);
or U2632 (N_2632,N_1206,N_1843);
nor U2633 (N_2633,N_1543,N_1385);
and U2634 (N_2634,N_1340,N_1474);
nor U2635 (N_2635,N_1771,N_1388);
nand U2636 (N_2636,N_1070,N_1486);
or U2637 (N_2637,N_1626,N_1910);
or U2638 (N_2638,N_1604,N_1883);
or U2639 (N_2639,N_1487,N_1268);
nor U2640 (N_2640,N_1337,N_1828);
nor U2641 (N_2641,N_1593,N_1627);
nor U2642 (N_2642,N_1023,N_1411);
nor U2643 (N_2643,N_1277,N_1171);
nand U2644 (N_2644,N_1901,N_1647);
and U2645 (N_2645,N_1081,N_1353);
nor U2646 (N_2646,N_1377,N_1274);
or U2647 (N_2647,N_1396,N_1595);
nand U2648 (N_2648,N_1339,N_1227);
nor U2649 (N_2649,N_1467,N_1351);
or U2650 (N_2650,N_1421,N_1139);
or U2651 (N_2651,N_1157,N_1960);
nand U2652 (N_2652,N_1353,N_1909);
xnor U2653 (N_2653,N_1449,N_1758);
nor U2654 (N_2654,N_1565,N_1145);
nand U2655 (N_2655,N_1028,N_1975);
nand U2656 (N_2656,N_1355,N_1882);
or U2657 (N_2657,N_1808,N_1517);
and U2658 (N_2658,N_1232,N_1179);
or U2659 (N_2659,N_1171,N_1243);
and U2660 (N_2660,N_1133,N_1380);
nand U2661 (N_2661,N_1041,N_1941);
or U2662 (N_2662,N_1632,N_1104);
nand U2663 (N_2663,N_1088,N_1121);
nor U2664 (N_2664,N_1314,N_1988);
or U2665 (N_2665,N_1544,N_1566);
nor U2666 (N_2666,N_1858,N_1112);
nand U2667 (N_2667,N_1821,N_1598);
nand U2668 (N_2668,N_1671,N_1350);
nor U2669 (N_2669,N_1365,N_1300);
nand U2670 (N_2670,N_1396,N_1880);
nand U2671 (N_2671,N_1634,N_1263);
nand U2672 (N_2672,N_1200,N_1738);
nor U2673 (N_2673,N_1348,N_1552);
nor U2674 (N_2674,N_1239,N_1847);
and U2675 (N_2675,N_1613,N_1817);
and U2676 (N_2676,N_1827,N_1761);
nor U2677 (N_2677,N_1018,N_1468);
or U2678 (N_2678,N_1362,N_1120);
nand U2679 (N_2679,N_1533,N_1601);
or U2680 (N_2680,N_1778,N_1120);
nor U2681 (N_2681,N_1256,N_1251);
nor U2682 (N_2682,N_1571,N_1167);
nor U2683 (N_2683,N_1867,N_1970);
or U2684 (N_2684,N_1354,N_1691);
nor U2685 (N_2685,N_1196,N_1052);
or U2686 (N_2686,N_1238,N_1373);
and U2687 (N_2687,N_1499,N_1936);
nand U2688 (N_2688,N_1379,N_1198);
nor U2689 (N_2689,N_1662,N_1881);
and U2690 (N_2690,N_1623,N_1714);
or U2691 (N_2691,N_1319,N_1487);
or U2692 (N_2692,N_1665,N_1934);
or U2693 (N_2693,N_1060,N_1806);
nand U2694 (N_2694,N_1302,N_1698);
or U2695 (N_2695,N_1153,N_1074);
or U2696 (N_2696,N_1763,N_1978);
or U2697 (N_2697,N_1510,N_1039);
and U2698 (N_2698,N_1904,N_1301);
or U2699 (N_2699,N_1782,N_1355);
nand U2700 (N_2700,N_1868,N_1457);
or U2701 (N_2701,N_1702,N_1680);
or U2702 (N_2702,N_1376,N_1225);
or U2703 (N_2703,N_1302,N_1309);
nor U2704 (N_2704,N_1810,N_1449);
nor U2705 (N_2705,N_1223,N_1828);
and U2706 (N_2706,N_1297,N_1065);
nand U2707 (N_2707,N_1346,N_1177);
and U2708 (N_2708,N_1355,N_1032);
nor U2709 (N_2709,N_1069,N_1765);
or U2710 (N_2710,N_1552,N_1607);
and U2711 (N_2711,N_1638,N_1018);
nor U2712 (N_2712,N_1328,N_1020);
nand U2713 (N_2713,N_1885,N_1366);
nor U2714 (N_2714,N_1453,N_1020);
nor U2715 (N_2715,N_1623,N_1947);
or U2716 (N_2716,N_1537,N_1189);
and U2717 (N_2717,N_1273,N_1803);
nand U2718 (N_2718,N_1017,N_1336);
or U2719 (N_2719,N_1153,N_1638);
nand U2720 (N_2720,N_1859,N_1465);
and U2721 (N_2721,N_1677,N_1761);
nor U2722 (N_2722,N_1332,N_1911);
nor U2723 (N_2723,N_1503,N_1861);
and U2724 (N_2724,N_1036,N_1086);
nor U2725 (N_2725,N_1136,N_1147);
nand U2726 (N_2726,N_1968,N_1789);
and U2727 (N_2727,N_1324,N_1870);
and U2728 (N_2728,N_1111,N_1468);
nand U2729 (N_2729,N_1192,N_1368);
nand U2730 (N_2730,N_1204,N_1319);
nor U2731 (N_2731,N_1776,N_1567);
and U2732 (N_2732,N_1316,N_1471);
nor U2733 (N_2733,N_1443,N_1801);
and U2734 (N_2734,N_1729,N_1118);
nand U2735 (N_2735,N_1623,N_1772);
and U2736 (N_2736,N_1355,N_1070);
nor U2737 (N_2737,N_1472,N_1828);
nand U2738 (N_2738,N_1333,N_1032);
nor U2739 (N_2739,N_1942,N_1395);
or U2740 (N_2740,N_1893,N_1171);
xnor U2741 (N_2741,N_1362,N_1474);
and U2742 (N_2742,N_1484,N_1830);
nand U2743 (N_2743,N_1726,N_1019);
and U2744 (N_2744,N_1378,N_1165);
and U2745 (N_2745,N_1339,N_1815);
or U2746 (N_2746,N_1485,N_1477);
or U2747 (N_2747,N_1463,N_1321);
or U2748 (N_2748,N_1686,N_1062);
and U2749 (N_2749,N_1925,N_1111);
or U2750 (N_2750,N_1597,N_1553);
and U2751 (N_2751,N_1954,N_1960);
or U2752 (N_2752,N_1325,N_1746);
and U2753 (N_2753,N_1952,N_1489);
nand U2754 (N_2754,N_1326,N_1931);
nand U2755 (N_2755,N_1544,N_1573);
or U2756 (N_2756,N_1951,N_1451);
nor U2757 (N_2757,N_1774,N_1397);
and U2758 (N_2758,N_1461,N_1820);
and U2759 (N_2759,N_1435,N_1740);
nand U2760 (N_2760,N_1420,N_1443);
nor U2761 (N_2761,N_1409,N_1321);
and U2762 (N_2762,N_1965,N_1703);
or U2763 (N_2763,N_1057,N_1735);
or U2764 (N_2764,N_1467,N_1277);
and U2765 (N_2765,N_1118,N_1304);
and U2766 (N_2766,N_1790,N_1262);
and U2767 (N_2767,N_1549,N_1390);
or U2768 (N_2768,N_1056,N_1956);
or U2769 (N_2769,N_1399,N_1257);
nor U2770 (N_2770,N_1795,N_1247);
nand U2771 (N_2771,N_1362,N_1535);
and U2772 (N_2772,N_1648,N_1367);
and U2773 (N_2773,N_1777,N_1603);
nand U2774 (N_2774,N_1292,N_1265);
and U2775 (N_2775,N_1953,N_1473);
nand U2776 (N_2776,N_1672,N_1795);
or U2777 (N_2777,N_1732,N_1401);
and U2778 (N_2778,N_1501,N_1002);
nor U2779 (N_2779,N_1113,N_1184);
nand U2780 (N_2780,N_1987,N_1357);
xor U2781 (N_2781,N_1583,N_1627);
or U2782 (N_2782,N_1856,N_1982);
and U2783 (N_2783,N_1375,N_1390);
or U2784 (N_2784,N_1664,N_1306);
nand U2785 (N_2785,N_1206,N_1896);
nor U2786 (N_2786,N_1775,N_1866);
or U2787 (N_2787,N_1081,N_1080);
and U2788 (N_2788,N_1817,N_1626);
and U2789 (N_2789,N_1709,N_1975);
and U2790 (N_2790,N_1664,N_1840);
and U2791 (N_2791,N_1600,N_1372);
nor U2792 (N_2792,N_1940,N_1635);
nand U2793 (N_2793,N_1452,N_1074);
or U2794 (N_2794,N_1951,N_1397);
and U2795 (N_2795,N_1165,N_1463);
and U2796 (N_2796,N_1217,N_1473);
nand U2797 (N_2797,N_1059,N_1673);
and U2798 (N_2798,N_1249,N_1736);
nand U2799 (N_2799,N_1070,N_1397);
or U2800 (N_2800,N_1257,N_1140);
or U2801 (N_2801,N_1929,N_1033);
nand U2802 (N_2802,N_1070,N_1423);
and U2803 (N_2803,N_1262,N_1839);
and U2804 (N_2804,N_1913,N_1892);
nand U2805 (N_2805,N_1848,N_1918);
nand U2806 (N_2806,N_1039,N_1135);
nor U2807 (N_2807,N_1276,N_1436);
nand U2808 (N_2808,N_1676,N_1588);
nor U2809 (N_2809,N_1452,N_1728);
nor U2810 (N_2810,N_1207,N_1332);
nor U2811 (N_2811,N_1122,N_1244);
nor U2812 (N_2812,N_1194,N_1702);
nor U2813 (N_2813,N_1092,N_1341);
or U2814 (N_2814,N_1694,N_1888);
or U2815 (N_2815,N_1833,N_1047);
or U2816 (N_2816,N_1722,N_1460);
nand U2817 (N_2817,N_1143,N_1690);
or U2818 (N_2818,N_1523,N_1377);
nand U2819 (N_2819,N_1807,N_1573);
or U2820 (N_2820,N_1607,N_1399);
or U2821 (N_2821,N_1966,N_1517);
or U2822 (N_2822,N_1726,N_1515);
and U2823 (N_2823,N_1452,N_1738);
nand U2824 (N_2824,N_1942,N_1030);
nand U2825 (N_2825,N_1746,N_1663);
nor U2826 (N_2826,N_1581,N_1618);
nand U2827 (N_2827,N_1874,N_1211);
or U2828 (N_2828,N_1227,N_1071);
and U2829 (N_2829,N_1756,N_1203);
and U2830 (N_2830,N_1884,N_1286);
nand U2831 (N_2831,N_1179,N_1464);
or U2832 (N_2832,N_1743,N_1517);
or U2833 (N_2833,N_1071,N_1751);
or U2834 (N_2834,N_1550,N_1181);
or U2835 (N_2835,N_1275,N_1846);
nand U2836 (N_2836,N_1644,N_1041);
nor U2837 (N_2837,N_1958,N_1527);
nor U2838 (N_2838,N_1057,N_1082);
xor U2839 (N_2839,N_1510,N_1879);
and U2840 (N_2840,N_1215,N_1818);
and U2841 (N_2841,N_1355,N_1166);
and U2842 (N_2842,N_1786,N_1052);
nand U2843 (N_2843,N_1245,N_1049);
or U2844 (N_2844,N_1823,N_1965);
nor U2845 (N_2845,N_1985,N_1196);
and U2846 (N_2846,N_1665,N_1325);
or U2847 (N_2847,N_1360,N_1702);
nand U2848 (N_2848,N_1089,N_1950);
nand U2849 (N_2849,N_1535,N_1468);
nor U2850 (N_2850,N_1713,N_1430);
xor U2851 (N_2851,N_1655,N_1340);
or U2852 (N_2852,N_1766,N_1498);
nor U2853 (N_2853,N_1663,N_1541);
nor U2854 (N_2854,N_1415,N_1733);
nor U2855 (N_2855,N_1180,N_1857);
or U2856 (N_2856,N_1977,N_1330);
nand U2857 (N_2857,N_1645,N_1416);
or U2858 (N_2858,N_1959,N_1968);
nand U2859 (N_2859,N_1463,N_1113);
or U2860 (N_2860,N_1324,N_1379);
or U2861 (N_2861,N_1193,N_1636);
nor U2862 (N_2862,N_1188,N_1000);
or U2863 (N_2863,N_1243,N_1958);
or U2864 (N_2864,N_1132,N_1014);
xnor U2865 (N_2865,N_1782,N_1921);
or U2866 (N_2866,N_1563,N_1389);
nand U2867 (N_2867,N_1263,N_1669);
nor U2868 (N_2868,N_1940,N_1432);
and U2869 (N_2869,N_1560,N_1717);
nand U2870 (N_2870,N_1787,N_1588);
nand U2871 (N_2871,N_1732,N_1132);
nand U2872 (N_2872,N_1256,N_1783);
or U2873 (N_2873,N_1980,N_1569);
nand U2874 (N_2874,N_1578,N_1393);
nand U2875 (N_2875,N_1312,N_1376);
nor U2876 (N_2876,N_1897,N_1012);
and U2877 (N_2877,N_1907,N_1553);
and U2878 (N_2878,N_1216,N_1283);
nand U2879 (N_2879,N_1546,N_1413);
nand U2880 (N_2880,N_1598,N_1376);
nor U2881 (N_2881,N_1589,N_1450);
nand U2882 (N_2882,N_1329,N_1954);
nand U2883 (N_2883,N_1240,N_1005);
nand U2884 (N_2884,N_1461,N_1338);
and U2885 (N_2885,N_1474,N_1112);
and U2886 (N_2886,N_1845,N_1965);
nor U2887 (N_2887,N_1324,N_1465);
nand U2888 (N_2888,N_1747,N_1309);
and U2889 (N_2889,N_1757,N_1847);
and U2890 (N_2890,N_1190,N_1751);
nand U2891 (N_2891,N_1140,N_1695);
and U2892 (N_2892,N_1186,N_1345);
or U2893 (N_2893,N_1779,N_1629);
and U2894 (N_2894,N_1217,N_1412);
nand U2895 (N_2895,N_1730,N_1764);
nor U2896 (N_2896,N_1151,N_1876);
nand U2897 (N_2897,N_1165,N_1616);
and U2898 (N_2898,N_1834,N_1441);
nor U2899 (N_2899,N_1171,N_1664);
and U2900 (N_2900,N_1148,N_1858);
nand U2901 (N_2901,N_1524,N_1474);
or U2902 (N_2902,N_1429,N_1488);
or U2903 (N_2903,N_1211,N_1044);
nand U2904 (N_2904,N_1564,N_1664);
or U2905 (N_2905,N_1668,N_1841);
nand U2906 (N_2906,N_1843,N_1400);
and U2907 (N_2907,N_1838,N_1219);
nand U2908 (N_2908,N_1826,N_1726);
nand U2909 (N_2909,N_1610,N_1009);
or U2910 (N_2910,N_1843,N_1994);
nand U2911 (N_2911,N_1770,N_1592);
and U2912 (N_2912,N_1435,N_1847);
nor U2913 (N_2913,N_1320,N_1857);
or U2914 (N_2914,N_1079,N_1971);
or U2915 (N_2915,N_1778,N_1953);
and U2916 (N_2916,N_1657,N_1648);
nand U2917 (N_2917,N_1469,N_1417);
nand U2918 (N_2918,N_1210,N_1793);
nand U2919 (N_2919,N_1960,N_1200);
nand U2920 (N_2920,N_1429,N_1691);
nand U2921 (N_2921,N_1100,N_1272);
nor U2922 (N_2922,N_1603,N_1555);
nor U2923 (N_2923,N_1333,N_1632);
nand U2924 (N_2924,N_1146,N_1923);
nand U2925 (N_2925,N_1996,N_1105);
and U2926 (N_2926,N_1313,N_1698);
nor U2927 (N_2927,N_1432,N_1346);
nand U2928 (N_2928,N_1021,N_1489);
and U2929 (N_2929,N_1624,N_1345);
nand U2930 (N_2930,N_1554,N_1110);
and U2931 (N_2931,N_1810,N_1669);
nor U2932 (N_2932,N_1150,N_1155);
and U2933 (N_2933,N_1477,N_1165);
or U2934 (N_2934,N_1511,N_1167);
nor U2935 (N_2935,N_1723,N_1392);
nor U2936 (N_2936,N_1307,N_1116);
nand U2937 (N_2937,N_1304,N_1038);
or U2938 (N_2938,N_1551,N_1759);
nand U2939 (N_2939,N_1797,N_1516);
nand U2940 (N_2940,N_1996,N_1896);
or U2941 (N_2941,N_1202,N_1516);
nand U2942 (N_2942,N_1058,N_1473);
nand U2943 (N_2943,N_1064,N_1412);
nor U2944 (N_2944,N_1736,N_1363);
or U2945 (N_2945,N_1395,N_1612);
nand U2946 (N_2946,N_1039,N_1742);
or U2947 (N_2947,N_1211,N_1328);
and U2948 (N_2948,N_1521,N_1343);
or U2949 (N_2949,N_1551,N_1924);
nand U2950 (N_2950,N_1292,N_1018);
nand U2951 (N_2951,N_1481,N_1120);
nand U2952 (N_2952,N_1655,N_1867);
or U2953 (N_2953,N_1568,N_1632);
and U2954 (N_2954,N_1416,N_1789);
or U2955 (N_2955,N_1893,N_1464);
nor U2956 (N_2956,N_1291,N_1962);
nor U2957 (N_2957,N_1107,N_1339);
nand U2958 (N_2958,N_1931,N_1723);
and U2959 (N_2959,N_1256,N_1020);
nand U2960 (N_2960,N_1531,N_1731);
nor U2961 (N_2961,N_1451,N_1580);
nor U2962 (N_2962,N_1905,N_1690);
nand U2963 (N_2963,N_1991,N_1383);
and U2964 (N_2964,N_1336,N_1811);
or U2965 (N_2965,N_1757,N_1476);
nand U2966 (N_2966,N_1836,N_1715);
or U2967 (N_2967,N_1915,N_1675);
or U2968 (N_2968,N_1388,N_1330);
nor U2969 (N_2969,N_1362,N_1125);
and U2970 (N_2970,N_1706,N_1453);
nand U2971 (N_2971,N_1656,N_1601);
nor U2972 (N_2972,N_1363,N_1931);
nand U2973 (N_2973,N_1821,N_1172);
and U2974 (N_2974,N_1757,N_1693);
nand U2975 (N_2975,N_1403,N_1120);
and U2976 (N_2976,N_1458,N_1600);
and U2977 (N_2977,N_1058,N_1115);
and U2978 (N_2978,N_1999,N_1071);
or U2979 (N_2979,N_1440,N_1505);
or U2980 (N_2980,N_1362,N_1546);
or U2981 (N_2981,N_1788,N_1416);
or U2982 (N_2982,N_1324,N_1137);
xor U2983 (N_2983,N_1221,N_1840);
nand U2984 (N_2984,N_1027,N_1956);
or U2985 (N_2985,N_1871,N_1300);
and U2986 (N_2986,N_1275,N_1806);
and U2987 (N_2987,N_1869,N_1855);
nor U2988 (N_2988,N_1092,N_1838);
or U2989 (N_2989,N_1200,N_1029);
or U2990 (N_2990,N_1473,N_1195);
or U2991 (N_2991,N_1690,N_1131);
nor U2992 (N_2992,N_1056,N_1481);
and U2993 (N_2993,N_1703,N_1691);
and U2994 (N_2994,N_1582,N_1641);
or U2995 (N_2995,N_1355,N_1196);
or U2996 (N_2996,N_1724,N_1613);
nand U2997 (N_2997,N_1499,N_1952);
and U2998 (N_2998,N_1983,N_1503);
and U2999 (N_2999,N_1150,N_1135);
and U3000 (N_3000,N_2474,N_2696);
nand U3001 (N_3001,N_2140,N_2220);
nor U3002 (N_3002,N_2229,N_2968);
or U3003 (N_3003,N_2961,N_2235);
and U3004 (N_3004,N_2701,N_2245);
nor U3005 (N_3005,N_2392,N_2174);
nor U3006 (N_3006,N_2539,N_2413);
nand U3007 (N_3007,N_2595,N_2818);
or U3008 (N_3008,N_2124,N_2391);
or U3009 (N_3009,N_2939,N_2500);
nand U3010 (N_3010,N_2209,N_2752);
nor U3011 (N_3011,N_2334,N_2768);
and U3012 (N_3012,N_2410,N_2181);
or U3013 (N_3013,N_2447,N_2036);
nor U3014 (N_3014,N_2812,N_2241);
and U3015 (N_3015,N_2657,N_2033);
or U3016 (N_3016,N_2353,N_2093);
nand U3017 (N_3017,N_2553,N_2148);
nand U3018 (N_3018,N_2007,N_2041);
nand U3019 (N_3019,N_2321,N_2848);
nand U3020 (N_3020,N_2785,N_2890);
nand U3021 (N_3021,N_2782,N_2015);
nor U3022 (N_3022,N_2921,N_2069);
nand U3023 (N_3023,N_2061,N_2099);
nor U3024 (N_3024,N_2804,N_2516);
nand U3025 (N_3025,N_2364,N_2826);
nand U3026 (N_3026,N_2359,N_2847);
nor U3027 (N_3027,N_2728,N_2686);
or U3028 (N_3028,N_2621,N_2540);
and U3029 (N_3029,N_2278,N_2313);
and U3030 (N_3030,N_2611,N_2569);
nand U3031 (N_3031,N_2233,N_2064);
and U3032 (N_3032,N_2024,N_2045);
nand U3033 (N_3033,N_2868,N_2947);
nand U3034 (N_3034,N_2135,N_2730);
or U3035 (N_3035,N_2593,N_2940);
nand U3036 (N_3036,N_2675,N_2488);
and U3037 (N_3037,N_2419,N_2892);
nand U3038 (N_3038,N_2107,N_2376);
and U3039 (N_3039,N_2133,N_2487);
nor U3040 (N_3040,N_2470,N_2435);
xnor U3041 (N_3041,N_2159,N_2213);
and U3042 (N_3042,N_2199,N_2417);
or U3043 (N_3043,N_2337,N_2663);
or U3044 (N_3044,N_2171,N_2034);
nand U3045 (N_3045,N_2508,N_2214);
nor U3046 (N_3046,N_2506,N_2741);
or U3047 (N_3047,N_2620,N_2832);
nand U3048 (N_3048,N_2923,N_2808);
and U3049 (N_3049,N_2018,N_2844);
nor U3050 (N_3050,N_2924,N_2941);
nand U3051 (N_3051,N_2716,N_2173);
or U3052 (N_3052,N_2772,N_2354);
nand U3053 (N_3053,N_2079,N_2601);
nor U3054 (N_3054,N_2745,N_2095);
and U3055 (N_3055,N_2212,N_2455);
xnor U3056 (N_3056,N_2617,N_2993);
nand U3057 (N_3057,N_2368,N_2971);
nor U3058 (N_3058,N_2268,N_2980);
nand U3059 (N_3059,N_2915,N_2551);
nor U3060 (N_3060,N_2907,N_2115);
nand U3061 (N_3061,N_2454,N_2048);
and U3062 (N_3062,N_2127,N_2951);
nand U3063 (N_3063,N_2533,N_2379);
xnor U3064 (N_3064,N_2709,N_2513);
nand U3065 (N_3065,N_2625,N_2706);
or U3066 (N_3066,N_2491,N_2906);
or U3067 (N_3067,N_2444,N_2913);
nand U3068 (N_3068,N_2096,N_2265);
or U3069 (N_3069,N_2217,N_2116);
and U3070 (N_3070,N_2332,N_2598);
nor U3071 (N_3071,N_2578,N_2074);
or U3072 (N_3072,N_2985,N_2824);
and U3073 (N_3073,N_2762,N_2527);
and U3074 (N_3074,N_2575,N_2777);
nand U3075 (N_3075,N_2280,N_2319);
and U3076 (N_3076,N_2662,N_2408);
nand U3077 (N_3077,N_2149,N_2560);
nor U3078 (N_3078,N_2386,N_2082);
nor U3079 (N_3079,N_2381,N_2342);
nand U3080 (N_3080,N_2006,N_2987);
nor U3081 (N_3081,N_2315,N_2628);
or U3082 (N_3082,N_2011,N_2218);
or U3083 (N_3083,N_2108,N_2434);
nor U3084 (N_3084,N_2727,N_2234);
and U3085 (N_3085,N_2712,N_2242);
nor U3086 (N_3086,N_2162,N_2729);
nor U3087 (N_3087,N_2534,N_2667);
and U3088 (N_3088,N_2883,N_2801);
or U3089 (N_3089,N_2432,N_2948);
nand U3090 (N_3090,N_2122,N_2900);
and U3091 (N_3091,N_2949,N_2813);
and U3092 (N_3092,N_2404,N_2990);
and U3093 (N_3093,N_2425,N_2552);
or U3094 (N_3094,N_2695,N_2749);
and U3095 (N_3095,N_2955,N_2823);
nor U3096 (N_3096,N_2161,N_2778);
and U3097 (N_3097,N_2277,N_2304);
nand U3098 (N_3098,N_2889,N_2713);
or U3099 (N_3099,N_2251,N_2618);
nand U3100 (N_3100,N_2458,N_2022);
nor U3101 (N_3101,N_2424,N_2867);
or U3102 (N_3102,N_2072,N_2091);
or U3103 (N_3103,N_2537,N_2839);
nor U3104 (N_3104,N_2751,N_2270);
and U3105 (N_3105,N_2158,N_2744);
nor U3106 (N_3106,N_2682,N_2292);
nor U3107 (N_3107,N_2333,N_2763);
nor U3108 (N_3108,N_2462,N_2030);
or U3109 (N_3109,N_2860,N_2274);
or U3110 (N_3110,N_2493,N_2232);
and U3111 (N_3111,N_2416,N_2360);
nor U3112 (N_3112,N_2739,N_2957);
or U3113 (N_3113,N_2509,N_2166);
nor U3114 (N_3114,N_2974,N_2450);
and U3115 (N_3115,N_2878,N_2001);
nor U3116 (N_3116,N_2597,N_2774);
and U3117 (N_3117,N_2666,N_2685);
or U3118 (N_3118,N_2723,N_2795);
or U3119 (N_3119,N_2572,N_2835);
nor U3120 (N_3120,N_2151,N_2336);
nand U3121 (N_3121,N_2576,N_2524);
or U3122 (N_3122,N_2427,N_2038);
and U3123 (N_3123,N_2347,N_2211);
nand U3124 (N_3124,N_2609,N_2515);
nand U3125 (N_3125,N_2880,N_2356);
and U3126 (N_3126,N_2914,N_2262);
nor U3127 (N_3127,N_2950,N_2440);
nand U3128 (N_3128,N_2719,N_2825);
nand U3129 (N_3129,N_2445,N_2718);
nand U3130 (N_3130,N_2542,N_2326);
and U3131 (N_3131,N_2479,N_2874);
and U3132 (N_3132,N_2363,N_2845);
and U3133 (N_3133,N_2571,N_2495);
and U3134 (N_3134,N_2786,N_2403);
or U3135 (N_3135,N_2201,N_2400);
nor U3136 (N_3136,N_2283,N_2550);
nor U3137 (N_3137,N_2766,N_2215);
nor U3138 (N_3138,N_2464,N_2699);
and U3139 (N_3139,N_2260,N_2514);
nand U3140 (N_3140,N_2700,N_2112);
nand U3141 (N_3141,N_2080,N_2358);
nor U3142 (N_3142,N_2991,N_2303);
and U3143 (N_3143,N_2518,N_2330);
nor U3144 (N_3144,N_2089,N_2769);
and U3145 (N_3145,N_2687,N_2545);
and U3146 (N_3146,N_2021,N_2743);
and U3147 (N_3147,N_2630,N_2637);
and U3148 (N_3148,N_2558,N_2796);
and U3149 (N_3149,N_2642,N_2849);
and U3150 (N_3150,N_2163,N_2840);
and U3151 (N_3151,N_2945,N_2480);
nor U3152 (N_3152,N_2067,N_2613);
and U3153 (N_3153,N_2028,N_2012);
or U3154 (N_3154,N_2643,N_2224);
or U3155 (N_3155,N_2760,N_2992);
nor U3156 (N_3156,N_2688,N_2589);
or U3157 (N_3157,N_2414,N_2075);
or U3158 (N_3158,N_2517,N_2903);
nor U3159 (N_3159,N_2126,N_2633);
nor U3160 (N_3160,N_2486,N_2371);
and U3161 (N_3161,N_2145,N_2930);
and U3162 (N_3162,N_2655,N_2136);
and U3163 (N_3163,N_2412,N_2721);
or U3164 (N_3164,N_2855,N_2255);
nor U3165 (N_3165,N_2918,N_2928);
or U3166 (N_3166,N_2014,N_2966);
nor U3167 (N_3167,N_2311,N_2559);
or U3168 (N_3168,N_2894,N_2624);
nor U3169 (N_3169,N_2714,N_2086);
and U3170 (N_3170,N_2398,N_2580);
nor U3171 (N_3171,N_2710,N_2120);
or U3172 (N_3172,N_2259,N_2473);
nand U3173 (N_3173,N_2600,N_2281);
and U3174 (N_3174,N_2908,N_2927);
nor U3175 (N_3175,N_2636,N_2429);
nor U3176 (N_3176,N_2887,N_2694);
and U3177 (N_3177,N_2053,N_2221);
nand U3178 (N_3178,N_2790,N_2563);
nand U3179 (N_3179,N_2415,N_2877);
nor U3180 (N_3180,N_2302,N_2037);
and U3181 (N_3181,N_2390,N_2426);
nor U3182 (N_3182,N_2168,N_2267);
nand U3183 (N_3183,N_2737,N_2969);
nand U3184 (N_3184,N_2736,N_2420);
and U3185 (N_3185,N_2640,N_2556);
xor U3186 (N_3186,N_2704,N_2791);
nand U3187 (N_3187,N_2626,N_2461);
or U3188 (N_3188,N_2372,N_2418);
or U3189 (N_3189,N_2943,N_2238);
and U3190 (N_3190,N_2100,N_2344);
nor U3191 (N_3191,N_2726,N_2809);
nand U3192 (N_3192,N_2627,N_2382);
or U3193 (N_3193,N_2060,N_2103);
nor U3194 (N_3194,N_2439,N_2073);
nand U3195 (N_3195,N_2216,N_2478);
or U3196 (N_3196,N_2183,N_2512);
and U3197 (N_3197,N_2044,N_2853);
nand U3198 (N_3198,N_2407,N_2223);
or U3199 (N_3199,N_2222,N_2562);
nand U3200 (N_3200,N_2557,N_2476);
or U3201 (N_3201,N_2240,N_2130);
nand U3202 (N_3202,N_2647,N_2972);
nor U3203 (N_3203,N_2606,N_2187);
or U3204 (N_3204,N_2423,N_2979);
nand U3205 (N_3205,N_2463,N_2361);
nor U3206 (N_3206,N_2443,N_2679);
nor U3207 (N_3207,N_2293,N_2206);
and U3208 (N_3208,N_2020,N_2841);
nor U3209 (N_3209,N_2922,N_2043);
nand U3210 (N_3210,N_2659,N_2471);
or U3211 (N_3211,N_2697,N_2494);
or U3212 (N_3212,N_2731,N_2873);
nor U3213 (N_3213,N_2816,N_2891);
and U3214 (N_3214,N_2905,N_2146);
and U3215 (N_3215,N_2573,N_2466);
or U3216 (N_3216,N_2733,N_2735);
and U3217 (N_3217,N_2094,N_2803);
or U3218 (N_3218,N_2585,N_2156);
and U3219 (N_3219,N_2071,N_2568);
nand U3220 (N_3220,N_2077,N_2665);
nor U3221 (N_3221,N_2169,N_2295);
nor U3222 (N_3222,N_2810,N_2190);
nor U3223 (N_3223,N_2180,N_2608);
nor U3224 (N_3224,N_2118,N_2370);
nor U3225 (N_3225,N_2482,N_2317);
nor U3226 (N_3226,N_2207,N_2884);
and U3227 (N_3227,N_2000,N_2680);
or U3228 (N_3228,N_2449,N_2062);
nand U3229 (N_3229,N_2155,N_2057);
or U3230 (N_3230,N_2324,N_2339);
and U3231 (N_3231,N_2097,N_2252);
and U3232 (N_3232,N_2586,N_2646);
xnor U3233 (N_3233,N_2997,N_2871);
nand U3234 (N_3234,N_2555,N_2910);
nor U3235 (N_3235,N_2904,N_2285);
nor U3236 (N_3236,N_2742,N_2465);
or U3237 (N_3237,N_2632,N_2055);
or U3238 (N_3238,N_2437,N_2588);
nor U3239 (N_3239,N_2362,N_2109);
nand U3240 (N_3240,N_2177,N_2561);
or U3241 (N_3241,N_2164,N_2203);
or U3242 (N_3242,N_2366,N_2978);
or U3243 (N_3243,N_2834,N_2895);
nor U3244 (N_3244,N_2674,N_2179);
nor U3245 (N_3245,N_2864,N_2554);
or U3246 (N_3246,N_2629,N_2225);
and U3247 (N_3247,N_2504,N_2092);
nand U3248 (N_3248,N_2248,N_2005);
or U3249 (N_3249,N_2670,N_2854);
nand U3250 (N_3250,N_2770,N_2389);
or U3251 (N_3251,N_2377,N_2289);
nand U3252 (N_3252,N_2639,N_2862);
or U3253 (N_3253,N_2101,N_2388);
or U3254 (N_3254,N_2702,N_2469);
or U3255 (N_3255,N_2811,N_2087);
or U3256 (N_3256,N_2638,N_2231);
nand U3257 (N_3257,N_2357,N_2049);
and U3258 (N_3258,N_2352,N_2689);
or U3259 (N_3259,N_2305,N_2129);
nand U3260 (N_3260,N_2119,N_2153);
nand U3261 (N_3261,N_2881,N_2615);
nor U3262 (N_3262,N_2150,N_2147);
and U3263 (N_3263,N_2802,N_2298);
nor U3264 (N_3264,N_2604,N_2652);
nor U3265 (N_3265,N_2226,N_2200);
or U3266 (N_3266,N_2959,N_2349);
or U3267 (N_3267,N_2128,N_2882);
and U3268 (N_3268,N_2720,N_2564);
nand U3269 (N_3269,N_2935,N_2658);
nor U3270 (N_3270,N_2793,N_2523);
and U3271 (N_3271,N_2228,N_2300);
nor U3272 (N_3272,N_2901,N_2975);
nand U3273 (N_3273,N_2771,N_2934);
or U3274 (N_3274,N_2227,N_2477);
and U3275 (N_3275,N_2986,N_2247);
or U3276 (N_3276,N_2837,N_2291);
and U3277 (N_3277,N_2648,N_2290);
nor U3278 (N_3278,N_2954,N_2995);
nand U3279 (N_3279,N_2063,N_2483);
nor U3280 (N_3280,N_2886,N_2195);
nor U3281 (N_3281,N_2936,N_2253);
and U3282 (N_3282,N_2931,N_2870);
or U3283 (N_3283,N_2170,N_2178);
xnor U3284 (N_3284,N_2110,N_2430);
and U3285 (N_3285,N_2409,N_2799);
nand U3286 (N_3286,N_2485,N_2467);
or U3287 (N_3287,N_2343,N_2567);
and U3288 (N_3288,N_2944,N_2896);
nand U3289 (N_3289,N_2788,N_2405);
nand U3290 (N_3290,N_2275,N_2387);
nand U3291 (N_3291,N_2775,N_2738);
nand U3292 (N_3292,N_2831,N_2898);
or U3293 (N_3293,N_2938,N_2269);
or U3294 (N_3294,N_2929,N_2032);
nor U3295 (N_3295,N_2258,N_2926);
nor U3296 (N_3296,N_2520,N_2186);
or U3297 (N_3297,N_2973,N_2098);
nand U3298 (N_3298,N_2401,N_2084);
and U3299 (N_3299,N_2876,N_2673);
or U3300 (N_3300,N_2152,N_2040);
xor U3301 (N_3301,N_2919,N_2605);
or U3302 (N_3302,N_2244,N_2917);
nor U3303 (N_3303,N_2350,N_2983);
nor U3304 (N_3304,N_2789,N_2711);
nand U3305 (N_3305,N_2393,N_2994);
nand U3306 (N_3306,N_2998,N_2088);
nand U3307 (N_3307,N_2916,N_2507);
nor U3308 (N_3308,N_2654,N_2396);
or U3309 (N_3309,N_2031,N_2590);
or U3310 (N_3310,N_2246,N_2602);
and U3311 (N_3311,N_2541,N_2182);
nand U3312 (N_3312,N_2003,N_2645);
or U3313 (N_3313,N_2607,N_2530);
xnor U3314 (N_3314,N_2599,N_2176);
and U3315 (N_3315,N_2838,N_2584);
and U3316 (N_3316,N_2406,N_2276);
nand U3317 (N_3317,N_2373,N_2902);
and U3318 (N_3318,N_2858,N_2671);
nor U3319 (N_3319,N_2622,N_2996);
or U3320 (N_3320,N_2411,N_2309);
or U3321 (N_3321,N_2861,N_2946);
or U3322 (N_3322,N_2510,N_2776);
nor U3323 (N_3323,N_2113,N_2457);
or U3324 (N_3324,N_2453,N_2594);
or U3325 (N_3325,N_2167,N_2348);
or U3326 (N_3326,N_2511,N_2820);
nand U3327 (N_3327,N_2833,N_2193);
or U3328 (N_3328,N_2002,N_2273);
and U3329 (N_3329,N_2338,N_2428);
nand U3330 (N_3330,N_2757,N_2165);
or U3331 (N_3331,N_2765,N_2528);
or U3332 (N_3332,N_2869,N_2956);
and U3333 (N_3333,N_2355,N_2684);
nand U3334 (N_3334,N_2829,N_2656);
nor U3335 (N_3335,N_2784,N_2197);
nand U3336 (N_3336,N_2397,N_2492);
nand U3337 (N_3337,N_2351,N_2341);
and U3338 (N_3338,N_2385,N_2017);
or U3339 (N_3339,N_2383,N_2123);
and U3340 (N_3340,N_2953,N_2335);
or U3341 (N_3341,N_2806,N_2787);
nand U3342 (N_3342,N_2800,N_2703);
and U3343 (N_3343,N_2192,N_2125);
and U3344 (N_3344,N_2677,N_2888);
nand U3345 (N_3345,N_2746,N_2436);
and U3346 (N_3346,N_2189,N_2548);
nor U3347 (N_3347,N_2284,N_2821);
nand U3348 (N_3348,N_2340,N_2962);
nor U3349 (N_3349,N_2256,N_2982);
nand U3350 (N_3350,N_2967,N_2346);
nor U3351 (N_3351,N_2066,N_2814);
nor U3352 (N_3352,N_2958,N_2016);
nand U3353 (N_3353,N_2433,N_2254);
nand U3354 (N_3354,N_2374,N_2933);
and U3355 (N_3355,N_2641,N_2104);
or U3356 (N_3356,N_2960,N_2724);
nor U3357 (N_3357,N_2549,N_2318);
or U3358 (N_3358,N_2664,N_2484);
nor U3359 (N_3359,N_2230,N_2591);
nand U3360 (N_3360,N_2239,N_2475);
nor U3361 (N_3361,N_2297,N_2807);
nor U3362 (N_3362,N_2631,N_2725);
nand U3363 (N_3363,N_2852,N_2767);
and U3364 (N_3364,N_2683,N_2764);
nand U3365 (N_3365,N_2644,N_2828);
or U3366 (N_3366,N_2085,N_2544);
xnor U3367 (N_3367,N_2013,N_2202);
and U3368 (N_3368,N_2911,N_2137);
nand U3369 (N_3369,N_2989,N_2117);
and U3370 (N_3370,N_2750,N_2328);
nor U3371 (N_3371,N_2025,N_2287);
nand U3372 (N_3372,N_2596,N_2008);
nor U3373 (N_3373,N_2587,N_2603);
and U3374 (N_3374,N_2144,N_2266);
nor U3375 (N_3375,N_2157,N_2312);
nor U3376 (N_3376,N_2984,N_2367);
or U3377 (N_3377,N_2431,N_2925);
or U3378 (N_3378,N_2472,N_2394);
or U3379 (N_3379,N_2131,N_2805);
or U3380 (N_3380,N_2532,N_2634);
nor U3381 (N_3381,N_2210,N_2830);
nand U3382 (N_3382,N_2649,N_2325);
and U3383 (N_3383,N_2866,N_2623);
nand U3384 (N_3384,N_2068,N_2138);
or U3385 (N_3385,N_2378,N_2384);
nor U3386 (N_3386,N_2740,N_2172);
and U3387 (N_3387,N_2441,N_2536);
and U3388 (N_3388,N_2204,N_2612);
nand U3389 (N_3389,N_2009,N_2365);
nand U3390 (N_3390,N_2660,N_2056);
or U3391 (N_3391,N_2759,N_2893);
or U3392 (N_3392,N_2574,N_2546);
nand U3393 (N_3393,N_2160,N_2083);
nand U3394 (N_3394,N_2219,N_2327);
nand U3395 (N_3395,N_2614,N_2754);
nand U3396 (N_3396,N_2827,N_2196);
or U3397 (N_3397,N_2942,N_2395);
nand U3398 (N_3398,N_2707,N_2619);
nor U3399 (N_3399,N_2236,N_2781);
nand U3400 (N_3400,N_2912,N_2308);
nand U3401 (N_3401,N_2154,N_2583);
and U3402 (N_3402,N_2143,N_2792);
or U3403 (N_3403,N_2375,N_2681);
and U3404 (N_3404,N_2846,N_2758);
or U3405 (N_3405,N_2314,N_2529);
and U3406 (N_3406,N_2970,N_2753);
nand U3407 (N_3407,N_2050,N_2191);
or U3408 (N_3408,N_2316,N_2208);
nand U3409 (N_3409,N_2322,N_2070);
and U3410 (N_3410,N_2748,N_2965);
and U3411 (N_3411,N_2422,N_2566);
nor U3412 (N_3412,N_2456,N_2460);
or U3413 (N_3413,N_2581,N_2650);
and U3414 (N_3414,N_2081,N_2819);
nor U3415 (N_3415,N_2761,N_2708);
or U3416 (N_3416,N_2198,N_2521);
nand U3417 (N_3417,N_2090,N_2565);
or U3418 (N_3418,N_2243,N_2451);
or U3419 (N_3419,N_2909,N_2286);
nand U3420 (N_3420,N_2981,N_2616);
and U3421 (N_3421,N_2857,N_2503);
or U3422 (N_3422,N_2184,N_2794);
nand U3423 (N_3423,N_2842,N_2132);
nand U3424 (N_3424,N_2279,N_2452);
nor U3425 (N_3425,N_2272,N_2052);
nand U3426 (N_3426,N_2299,N_2526);
nor U3427 (N_3427,N_2582,N_2592);
and U3428 (N_3428,N_2004,N_2773);
nor U3429 (N_3429,N_2047,N_2653);
or U3430 (N_3430,N_2734,N_2141);
and U3431 (N_3431,N_2489,N_2237);
nand U3432 (N_3432,N_2497,N_2635);
nor U3433 (N_3433,N_2693,N_2543);
or U3434 (N_3434,N_2519,N_2732);
or U3435 (N_3435,N_2023,N_2722);
or U3436 (N_3436,N_2747,N_2875);
nor U3437 (N_3437,N_2780,N_2977);
and U3438 (N_3438,N_2263,N_2964);
nand U3439 (N_3439,N_2194,N_2142);
nand U3440 (N_3440,N_2026,N_2698);
and U3441 (N_3441,N_2438,N_2668);
nor U3442 (N_3442,N_2897,N_2872);
or U3443 (N_3443,N_2496,N_2331);
nand U3444 (N_3444,N_2705,N_2783);
or U3445 (N_3445,N_2501,N_2345);
nand U3446 (N_3446,N_2815,N_2661);
or U3447 (N_3447,N_2817,N_2976);
or U3448 (N_3448,N_2651,N_2899);
or U3449 (N_3449,N_2271,N_2380);
nand U3450 (N_3450,N_2797,N_2920);
nand U3451 (N_3451,N_2421,N_2249);
or U3452 (N_3452,N_2859,N_2755);
or U3453 (N_3453,N_2850,N_2185);
nor U3454 (N_3454,N_2027,N_2856);
and U3455 (N_3455,N_2717,N_2019);
nor U3456 (N_3456,N_2522,N_2505);
or U3457 (N_3457,N_2525,N_2448);
nand U3458 (N_3458,N_2863,N_2282);
nand U3459 (N_3459,N_2121,N_2932);
nor U3460 (N_3460,N_2139,N_2952);
and U3461 (N_3461,N_2054,N_2134);
nand U3462 (N_3462,N_2264,N_2672);
and U3463 (N_3463,N_2690,N_2102);
and U3464 (N_3464,N_2879,N_2490);
or U3465 (N_3465,N_2547,N_2865);
nor U3466 (N_3466,N_2442,N_2307);
nor U3467 (N_3467,N_2468,N_2106);
or U3468 (N_3468,N_2058,N_2498);
and U3469 (N_3469,N_2296,N_2836);
nand U3470 (N_3470,N_2676,N_2250);
nor U3471 (N_3471,N_2310,N_2399);
or U3472 (N_3472,N_2261,N_2459);
or U3473 (N_3473,N_2039,N_2402);
or U3474 (N_3474,N_2010,N_2114);
and U3475 (N_3475,N_2306,N_2963);
or U3476 (N_3476,N_2329,N_2678);
and U3477 (N_3477,N_2538,N_2988);
nand U3478 (N_3478,N_2579,N_2288);
nand U3479 (N_3479,N_2756,N_2502);
and U3480 (N_3480,N_2059,N_2046);
or U3481 (N_3481,N_2065,N_2105);
or U3482 (N_3482,N_2779,N_2843);
and U3483 (N_3483,N_2999,N_2205);
nor U3484 (N_3484,N_2531,N_2570);
nand U3485 (N_3485,N_2691,N_2320);
or U3486 (N_3486,N_2294,N_2446);
nand U3487 (N_3487,N_2042,N_2851);
nor U3488 (N_3488,N_2369,N_2610);
or U3489 (N_3489,N_2535,N_2499);
nand U3490 (N_3490,N_2885,N_2798);
or U3491 (N_3491,N_2035,N_2111);
nor U3492 (N_3492,N_2257,N_2188);
or U3493 (N_3493,N_2029,N_2715);
nand U3494 (N_3494,N_2301,N_2078);
or U3495 (N_3495,N_2669,N_2937);
or U3496 (N_3496,N_2577,N_2822);
nand U3497 (N_3497,N_2481,N_2175);
nor U3498 (N_3498,N_2076,N_2323);
and U3499 (N_3499,N_2051,N_2692);
and U3500 (N_3500,N_2077,N_2262);
nand U3501 (N_3501,N_2002,N_2827);
nor U3502 (N_3502,N_2507,N_2079);
or U3503 (N_3503,N_2705,N_2382);
or U3504 (N_3504,N_2208,N_2498);
nand U3505 (N_3505,N_2701,N_2275);
or U3506 (N_3506,N_2236,N_2254);
nor U3507 (N_3507,N_2919,N_2954);
and U3508 (N_3508,N_2529,N_2764);
or U3509 (N_3509,N_2391,N_2756);
and U3510 (N_3510,N_2262,N_2078);
nand U3511 (N_3511,N_2328,N_2675);
and U3512 (N_3512,N_2811,N_2140);
nand U3513 (N_3513,N_2550,N_2900);
nand U3514 (N_3514,N_2642,N_2032);
and U3515 (N_3515,N_2653,N_2454);
nor U3516 (N_3516,N_2632,N_2709);
and U3517 (N_3517,N_2413,N_2071);
nor U3518 (N_3518,N_2781,N_2621);
and U3519 (N_3519,N_2411,N_2680);
nor U3520 (N_3520,N_2419,N_2741);
nor U3521 (N_3521,N_2684,N_2794);
nand U3522 (N_3522,N_2944,N_2531);
nand U3523 (N_3523,N_2203,N_2490);
nand U3524 (N_3524,N_2563,N_2696);
nand U3525 (N_3525,N_2573,N_2035);
nor U3526 (N_3526,N_2783,N_2119);
nand U3527 (N_3527,N_2591,N_2816);
and U3528 (N_3528,N_2682,N_2852);
or U3529 (N_3529,N_2486,N_2876);
nor U3530 (N_3530,N_2854,N_2727);
nor U3531 (N_3531,N_2240,N_2974);
nor U3532 (N_3532,N_2775,N_2768);
or U3533 (N_3533,N_2755,N_2557);
nand U3534 (N_3534,N_2475,N_2790);
nor U3535 (N_3535,N_2091,N_2705);
nor U3536 (N_3536,N_2118,N_2316);
or U3537 (N_3537,N_2373,N_2739);
xor U3538 (N_3538,N_2371,N_2279);
or U3539 (N_3539,N_2842,N_2820);
nand U3540 (N_3540,N_2422,N_2414);
and U3541 (N_3541,N_2966,N_2929);
nor U3542 (N_3542,N_2967,N_2634);
and U3543 (N_3543,N_2058,N_2141);
nor U3544 (N_3544,N_2708,N_2179);
or U3545 (N_3545,N_2926,N_2970);
nor U3546 (N_3546,N_2593,N_2713);
nor U3547 (N_3547,N_2483,N_2928);
or U3548 (N_3548,N_2852,N_2759);
nand U3549 (N_3549,N_2660,N_2835);
and U3550 (N_3550,N_2063,N_2340);
or U3551 (N_3551,N_2552,N_2837);
or U3552 (N_3552,N_2655,N_2587);
nand U3553 (N_3553,N_2523,N_2587);
or U3554 (N_3554,N_2433,N_2160);
nor U3555 (N_3555,N_2356,N_2494);
and U3556 (N_3556,N_2510,N_2039);
or U3557 (N_3557,N_2517,N_2547);
and U3558 (N_3558,N_2052,N_2562);
and U3559 (N_3559,N_2928,N_2349);
and U3560 (N_3560,N_2241,N_2073);
and U3561 (N_3561,N_2698,N_2478);
or U3562 (N_3562,N_2392,N_2245);
or U3563 (N_3563,N_2233,N_2857);
nor U3564 (N_3564,N_2272,N_2815);
and U3565 (N_3565,N_2631,N_2326);
or U3566 (N_3566,N_2623,N_2236);
nand U3567 (N_3567,N_2367,N_2696);
and U3568 (N_3568,N_2836,N_2411);
or U3569 (N_3569,N_2548,N_2841);
nand U3570 (N_3570,N_2344,N_2801);
nand U3571 (N_3571,N_2584,N_2215);
nand U3572 (N_3572,N_2623,N_2083);
or U3573 (N_3573,N_2314,N_2456);
or U3574 (N_3574,N_2312,N_2697);
nor U3575 (N_3575,N_2946,N_2970);
nor U3576 (N_3576,N_2530,N_2290);
or U3577 (N_3577,N_2178,N_2706);
or U3578 (N_3578,N_2980,N_2631);
nor U3579 (N_3579,N_2229,N_2390);
nand U3580 (N_3580,N_2377,N_2649);
and U3581 (N_3581,N_2826,N_2314);
nand U3582 (N_3582,N_2107,N_2464);
or U3583 (N_3583,N_2344,N_2797);
nand U3584 (N_3584,N_2128,N_2634);
nor U3585 (N_3585,N_2594,N_2910);
nor U3586 (N_3586,N_2261,N_2614);
or U3587 (N_3587,N_2691,N_2845);
nor U3588 (N_3588,N_2586,N_2727);
and U3589 (N_3589,N_2820,N_2272);
or U3590 (N_3590,N_2410,N_2044);
or U3591 (N_3591,N_2931,N_2978);
and U3592 (N_3592,N_2900,N_2952);
or U3593 (N_3593,N_2786,N_2529);
nand U3594 (N_3594,N_2748,N_2015);
nor U3595 (N_3595,N_2347,N_2310);
nor U3596 (N_3596,N_2113,N_2083);
or U3597 (N_3597,N_2087,N_2205);
or U3598 (N_3598,N_2147,N_2317);
and U3599 (N_3599,N_2981,N_2595);
or U3600 (N_3600,N_2782,N_2573);
and U3601 (N_3601,N_2555,N_2145);
or U3602 (N_3602,N_2379,N_2599);
and U3603 (N_3603,N_2495,N_2134);
or U3604 (N_3604,N_2696,N_2792);
nor U3605 (N_3605,N_2784,N_2747);
nor U3606 (N_3606,N_2777,N_2497);
and U3607 (N_3607,N_2097,N_2621);
nor U3608 (N_3608,N_2397,N_2622);
or U3609 (N_3609,N_2502,N_2999);
and U3610 (N_3610,N_2887,N_2708);
xnor U3611 (N_3611,N_2294,N_2908);
and U3612 (N_3612,N_2249,N_2315);
or U3613 (N_3613,N_2559,N_2254);
and U3614 (N_3614,N_2557,N_2341);
nor U3615 (N_3615,N_2294,N_2834);
and U3616 (N_3616,N_2535,N_2100);
nand U3617 (N_3617,N_2500,N_2252);
nand U3618 (N_3618,N_2581,N_2353);
nor U3619 (N_3619,N_2291,N_2879);
and U3620 (N_3620,N_2571,N_2646);
and U3621 (N_3621,N_2621,N_2578);
and U3622 (N_3622,N_2054,N_2129);
and U3623 (N_3623,N_2229,N_2144);
and U3624 (N_3624,N_2958,N_2061);
and U3625 (N_3625,N_2996,N_2072);
nor U3626 (N_3626,N_2814,N_2901);
and U3627 (N_3627,N_2611,N_2331);
nand U3628 (N_3628,N_2110,N_2409);
nand U3629 (N_3629,N_2943,N_2472);
or U3630 (N_3630,N_2661,N_2971);
nand U3631 (N_3631,N_2041,N_2432);
and U3632 (N_3632,N_2750,N_2191);
nand U3633 (N_3633,N_2402,N_2051);
or U3634 (N_3634,N_2408,N_2475);
nand U3635 (N_3635,N_2578,N_2952);
or U3636 (N_3636,N_2706,N_2621);
and U3637 (N_3637,N_2976,N_2512);
or U3638 (N_3638,N_2548,N_2482);
or U3639 (N_3639,N_2694,N_2227);
and U3640 (N_3640,N_2055,N_2197);
or U3641 (N_3641,N_2626,N_2019);
nor U3642 (N_3642,N_2523,N_2978);
nand U3643 (N_3643,N_2117,N_2850);
or U3644 (N_3644,N_2562,N_2542);
or U3645 (N_3645,N_2359,N_2347);
and U3646 (N_3646,N_2586,N_2490);
nor U3647 (N_3647,N_2070,N_2727);
and U3648 (N_3648,N_2537,N_2575);
or U3649 (N_3649,N_2851,N_2543);
or U3650 (N_3650,N_2272,N_2790);
or U3651 (N_3651,N_2429,N_2752);
nand U3652 (N_3652,N_2001,N_2422);
xor U3653 (N_3653,N_2969,N_2503);
nor U3654 (N_3654,N_2947,N_2930);
or U3655 (N_3655,N_2915,N_2074);
nand U3656 (N_3656,N_2297,N_2315);
nor U3657 (N_3657,N_2586,N_2635);
and U3658 (N_3658,N_2678,N_2358);
nand U3659 (N_3659,N_2606,N_2301);
nor U3660 (N_3660,N_2959,N_2483);
and U3661 (N_3661,N_2013,N_2458);
and U3662 (N_3662,N_2140,N_2475);
nor U3663 (N_3663,N_2344,N_2398);
or U3664 (N_3664,N_2593,N_2333);
or U3665 (N_3665,N_2294,N_2841);
or U3666 (N_3666,N_2018,N_2971);
nand U3667 (N_3667,N_2582,N_2214);
nand U3668 (N_3668,N_2421,N_2637);
or U3669 (N_3669,N_2367,N_2084);
nand U3670 (N_3670,N_2583,N_2821);
and U3671 (N_3671,N_2347,N_2963);
or U3672 (N_3672,N_2937,N_2486);
or U3673 (N_3673,N_2860,N_2644);
xor U3674 (N_3674,N_2394,N_2850);
or U3675 (N_3675,N_2367,N_2790);
and U3676 (N_3676,N_2027,N_2266);
or U3677 (N_3677,N_2415,N_2803);
nand U3678 (N_3678,N_2543,N_2237);
or U3679 (N_3679,N_2310,N_2127);
or U3680 (N_3680,N_2488,N_2057);
and U3681 (N_3681,N_2934,N_2485);
and U3682 (N_3682,N_2104,N_2452);
nor U3683 (N_3683,N_2405,N_2559);
nor U3684 (N_3684,N_2453,N_2873);
nand U3685 (N_3685,N_2422,N_2388);
nor U3686 (N_3686,N_2191,N_2273);
or U3687 (N_3687,N_2307,N_2942);
or U3688 (N_3688,N_2553,N_2545);
nor U3689 (N_3689,N_2575,N_2761);
and U3690 (N_3690,N_2887,N_2381);
nor U3691 (N_3691,N_2663,N_2896);
nand U3692 (N_3692,N_2955,N_2845);
or U3693 (N_3693,N_2376,N_2572);
nor U3694 (N_3694,N_2803,N_2411);
nand U3695 (N_3695,N_2838,N_2886);
nor U3696 (N_3696,N_2077,N_2876);
nand U3697 (N_3697,N_2707,N_2821);
or U3698 (N_3698,N_2760,N_2837);
nand U3699 (N_3699,N_2447,N_2715);
nor U3700 (N_3700,N_2108,N_2572);
and U3701 (N_3701,N_2042,N_2457);
or U3702 (N_3702,N_2608,N_2819);
nand U3703 (N_3703,N_2560,N_2112);
nor U3704 (N_3704,N_2186,N_2318);
nor U3705 (N_3705,N_2502,N_2099);
nor U3706 (N_3706,N_2025,N_2597);
nor U3707 (N_3707,N_2925,N_2484);
and U3708 (N_3708,N_2237,N_2247);
or U3709 (N_3709,N_2689,N_2381);
or U3710 (N_3710,N_2584,N_2441);
or U3711 (N_3711,N_2981,N_2211);
and U3712 (N_3712,N_2048,N_2620);
or U3713 (N_3713,N_2870,N_2530);
or U3714 (N_3714,N_2064,N_2157);
nor U3715 (N_3715,N_2739,N_2567);
or U3716 (N_3716,N_2350,N_2288);
or U3717 (N_3717,N_2306,N_2944);
nor U3718 (N_3718,N_2224,N_2516);
or U3719 (N_3719,N_2449,N_2165);
nand U3720 (N_3720,N_2632,N_2848);
nor U3721 (N_3721,N_2589,N_2339);
or U3722 (N_3722,N_2328,N_2121);
nand U3723 (N_3723,N_2594,N_2940);
and U3724 (N_3724,N_2201,N_2428);
nand U3725 (N_3725,N_2231,N_2544);
and U3726 (N_3726,N_2496,N_2850);
and U3727 (N_3727,N_2372,N_2361);
nor U3728 (N_3728,N_2759,N_2593);
and U3729 (N_3729,N_2326,N_2750);
or U3730 (N_3730,N_2798,N_2536);
or U3731 (N_3731,N_2074,N_2623);
nand U3732 (N_3732,N_2967,N_2635);
nand U3733 (N_3733,N_2233,N_2424);
and U3734 (N_3734,N_2591,N_2596);
and U3735 (N_3735,N_2551,N_2224);
or U3736 (N_3736,N_2644,N_2799);
nor U3737 (N_3737,N_2318,N_2247);
and U3738 (N_3738,N_2592,N_2365);
or U3739 (N_3739,N_2840,N_2152);
nor U3740 (N_3740,N_2256,N_2610);
and U3741 (N_3741,N_2961,N_2494);
nor U3742 (N_3742,N_2490,N_2643);
and U3743 (N_3743,N_2300,N_2852);
nor U3744 (N_3744,N_2139,N_2436);
or U3745 (N_3745,N_2457,N_2011);
nor U3746 (N_3746,N_2504,N_2395);
and U3747 (N_3747,N_2810,N_2532);
and U3748 (N_3748,N_2407,N_2732);
nand U3749 (N_3749,N_2838,N_2040);
nor U3750 (N_3750,N_2804,N_2689);
and U3751 (N_3751,N_2158,N_2477);
nor U3752 (N_3752,N_2391,N_2028);
and U3753 (N_3753,N_2444,N_2839);
nand U3754 (N_3754,N_2749,N_2220);
nor U3755 (N_3755,N_2814,N_2761);
and U3756 (N_3756,N_2090,N_2515);
or U3757 (N_3757,N_2115,N_2970);
or U3758 (N_3758,N_2153,N_2016);
nand U3759 (N_3759,N_2549,N_2326);
or U3760 (N_3760,N_2294,N_2836);
nand U3761 (N_3761,N_2517,N_2533);
nor U3762 (N_3762,N_2726,N_2851);
and U3763 (N_3763,N_2796,N_2187);
nand U3764 (N_3764,N_2112,N_2684);
nand U3765 (N_3765,N_2727,N_2905);
and U3766 (N_3766,N_2627,N_2959);
nand U3767 (N_3767,N_2095,N_2415);
nand U3768 (N_3768,N_2241,N_2397);
nor U3769 (N_3769,N_2942,N_2481);
nor U3770 (N_3770,N_2374,N_2893);
or U3771 (N_3771,N_2773,N_2425);
and U3772 (N_3772,N_2738,N_2009);
and U3773 (N_3773,N_2792,N_2920);
or U3774 (N_3774,N_2519,N_2113);
and U3775 (N_3775,N_2701,N_2347);
or U3776 (N_3776,N_2583,N_2551);
nand U3777 (N_3777,N_2996,N_2229);
nor U3778 (N_3778,N_2401,N_2144);
nand U3779 (N_3779,N_2631,N_2676);
and U3780 (N_3780,N_2624,N_2375);
nor U3781 (N_3781,N_2682,N_2398);
and U3782 (N_3782,N_2652,N_2912);
nand U3783 (N_3783,N_2817,N_2924);
or U3784 (N_3784,N_2693,N_2947);
or U3785 (N_3785,N_2043,N_2298);
nand U3786 (N_3786,N_2797,N_2982);
nand U3787 (N_3787,N_2405,N_2890);
or U3788 (N_3788,N_2463,N_2349);
and U3789 (N_3789,N_2610,N_2768);
nor U3790 (N_3790,N_2398,N_2994);
and U3791 (N_3791,N_2101,N_2545);
and U3792 (N_3792,N_2486,N_2192);
nand U3793 (N_3793,N_2150,N_2157);
and U3794 (N_3794,N_2399,N_2796);
or U3795 (N_3795,N_2226,N_2231);
nor U3796 (N_3796,N_2202,N_2957);
nor U3797 (N_3797,N_2376,N_2922);
nand U3798 (N_3798,N_2512,N_2037);
and U3799 (N_3799,N_2296,N_2284);
nor U3800 (N_3800,N_2214,N_2447);
and U3801 (N_3801,N_2998,N_2149);
nor U3802 (N_3802,N_2617,N_2930);
xnor U3803 (N_3803,N_2915,N_2647);
or U3804 (N_3804,N_2897,N_2118);
nand U3805 (N_3805,N_2722,N_2570);
nor U3806 (N_3806,N_2692,N_2503);
nor U3807 (N_3807,N_2712,N_2626);
or U3808 (N_3808,N_2049,N_2058);
and U3809 (N_3809,N_2601,N_2757);
nor U3810 (N_3810,N_2232,N_2120);
or U3811 (N_3811,N_2402,N_2231);
or U3812 (N_3812,N_2326,N_2288);
nor U3813 (N_3813,N_2136,N_2421);
nand U3814 (N_3814,N_2651,N_2448);
nand U3815 (N_3815,N_2680,N_2432);
nor U3816 (N_3816,N_2661,N_2409);
nor U3817 (N_3817,N_2400,N_2941);
or U3818 (N_3818,N_2174,N_2917);
or U3819 (N_3819,N_2912,N_2251);
and U3820 (N_3820,N_2605,N_2310);
or U3821 (N_3821,N_2426,N_2407);
nor U3822 (N_3822,N_2224,N_2375);
or U3823 (N_3823,N_2021,N_2197);
or U3824 (N_3824,N_2271,N_2819);
or U3825 (N_3825,N_2244,N_2065);
and U3826 (N_3826,N_2469,N_2957);
nand U3827 (N_3827,N_2923,N_2944);
nor U3828 (N_3828,N_2635,N_2881);
nand U3829 (N_3829,N_2865,N_2212);
and U3830 (N_3830,N_2266,N_2394);
and U3831 (N_3831,N_2357,N_2163);
and U3832 (N_3832,N_2847,N_2669);
nand U3833 (N_3833,N_2519,N_2502);
nor U3834 (N_3834,N_2717,N_2209);
nand U3835 (N_3835,N_2513,N_2945);
and U3836 (N_3836,N_2547,N_2531);
nand U3837 (N_3837,N_2945,N_2740);
nand U3838 (N_3838,N_2009,N_2608);
nand U3839 (N_3839,N_2693,N_2458);
or U3840 (N_3840,N_2429,N_2538);
and U3841 (N_3841,N_2615,N_2346);
or U3842 (N_3842,N_2566,N_2087);
and U3843 (N_3843,N_2001,N_2170);
nor U3844 (N_3844,N_2605,N_2874);
nand U3845 (N_3845,N_2575,N_2249);
nor U3846 (N_3846,N_2264,N_2708);
nand U3847 (N_3847,N_2537,N_2252);
nor U3848 (N_3848,N_2275,N_2061);
nand U3849 (N_3849,N_2583,N_2029);
or U3850 (N_3850,N_2072,N_2082);
nand U3851 (N_3851,N_2005,N_2704);
and U3852 (N_3852,N_2630,N_2114);
and U3853 (N_3853,N_2567,N_2839);
or U3854 (N_3854,N_2557,N_2914);
nand U3855 (N_3855,N_2543,N_2441);
or U3856 (N_3856,N_2777,N_2890);
nor U3857 (N_3857,N_2445,N_2255);
nor U3858 (N_3858,N_2153,N_2760);
or U3859 (N_3859,N_2407,N_2672);
or U3860 (N_3860,N_2527,N_2753);
nor U3861 (N_3861,N_2010,N_2492);
or U3862 (N_3862,N_2087,N_2679);
and U3863 (N_3863,N_2707,N_2279);
nand U3864 (N_3864,N_2019,N_2147);
or U3865 (N_3865,N_2633,N_2267);
and U3866 (N_3866,N_2210,N_2254);
nand U3867 (N_3867,N_2145,N_2722);
nand U3868 (N_3868,N_2453,N_2376);
or U3869 (N_3869,N_2524,N_2436);
or U3870 (N_3870,N_2814,N_2948);
nand U3871 (N_3871,N_2844,N_2444);
and U3872 (N_3872,N_2389,N_2789);
and U3873 (N_3873,N_2195,N_2506);
and U3874 (N_3874,N_2259,N_2661);
nand U3875 (N_3875,N_2225,N_2758);
nor U3876 (N_3876,N_2225,N_2247);
nor U3877 (N_3877,N_2525,N_2457);
nand U3878 (N_3878,N_2504,N_2638);
nand U3879 (N_3879,N_2246,N_2578);
or U3880 (N_3880,N_2051,N_2721);
or U3881 (N_3881,N_2890,N_2418);
or U3882 (N_3882,N_2029,N_2857);
nor U3883 (N_3883,N_2372,N_2925);
nor U3884 (N_3884,N_2089,N_2050);
and U3885 (N_3885,N_2930,N_2408);
and U3886 (N_3886,N_2138,N_2649);
nand U3887 (N_3887,N_2253,N_2009);
nor U3888 (N_3888,N_2158,N_2901);
nand U3889 (N_3889,N_2121,N_2453);
or U3890 (N_3890,N_2115,N_2029);
nand U3891 (N_3891,N_2175,N_2825);
or U3892 (N_3892,N_2790,N_2466);
and U3893 (N_3893,N_2294,N_2488);
nor U3894 (N_3894,N_2756,N_2191);
and U3895 (N_3895,N_2789,N_2054);
nand U3896 (N_3896,N_2975,N_2828);
and U3897 (N_3897,N_2244,N_2252);
nor U3898 (N_3898,N_2195,N_2945);
nand U3899 (N_3899,N_2562,N_2213);
nor U3900 (N_3900,N_2107,N_2885);
or U3901 (N_3901,N_2235,N_2574);
nor U3902 (N_3902,N_2021,N_2842);
nor U3903 (N_3903,N_2201,N_2137);
nor U3904 (N_3904,N_2598,N_2739);
and U3905 (N_3905,N_2712,N_2446);
or U3906 (N_3906,N_2629,N_2139);
nand U3907 (N_3907,N_2216,N_2276);
or U3908 (N_3908,N_2923,N_2149);
nor U3909 (N_3909,N_2956,N_2750);
nor U3910 (N_3910,N_2023,N_2878);
nor U3911 (N_3911,N_2545,N_2226);
and U3912 (N_3912,N_2616,N_2236);
or U3913 (N_3913,N_2047,N_2310);
nand U3914 (N_3914,N_2385,N_2665);
nor U3915 (N_3915,N_2512,N_2978);
and U3916 (N_3916,N_2142,N_2880);
or U3917 (N_3917,N_2760,N_2705);
or U3918 (N_3918,N_2255,N_2274);
or U3919 (N_3919,N_2767,N_2468);
nand U3920 (N_3920,N_2885,N_2245);
or U3921 (N_3921,N_2492,N_2168);
nor U3922 (N_3922,N_2761,N_2034);
nand U3923 (N_3923,N_2403,N_2073);
nor U3924 (N_3924,N_2895,N_2922);
nand U3925 (N_3925,N_2815,N_2062);
or U3926 (N_3926,N_2131,N_2436);
and U3927 (N_3927,N_2147,N_2248);
or U3928 (N_3928,N_2399,N_2023);
nor U3929 (N_3929,N_2276,N_2833);
nand U3930 (N_3930,N_2084,N_2087);
nor U3931 (N_3931,N_2083,N_2153);
nand U3932 (N_3932,N_2752,N_2162);
and U3933 (N_3933,N_2130,N_2556);
and U3934 (N_3934,N_2486,N_2143);
nor U3935 (N_3935,N_2096,N_2851);
nand U3936 (N_3936,N_2468,N_2489);
and U3937 (N_3937,N_2719,N_2357);
nor U3938 (N_3938,N_2476,N_2857);
nand U3939 (N_3939,N_2299,N_2478);
or U3940 (N_3940,N_2875,N_2225);
nor U3941 (N_3941,N_2872,N_2180);
and U3942 (N_3942,N_2606,N_2372);
or U3943 (N_3943,N_2502,N_2038);
and U3944 (N_3944,N_2603,N_2002);
and U3945 (N_3945,N_2544,N_2533);
and U3946 (N_3946,N_2842,N_2575);
and U3947 (N_3947,N_2662,N_2504);
and U3948 (N_3948,N_2493,N_2834);
nor U3949 (N_3949,N_2290,N_2246);
and U3950 (N_3950,N_2930,N_2989);
nand U3951 (N_3951,N_2789,N_2609);
or U3952 (N_3952,N_2620,N_2402);
nor U3953 (N_3953,N_2415,N_2444);
and U3954 (N_3954,N_2423,N_2075);
and U3955 (N_3955,N_2556,N_2008);
or U3956 (N_3956,N_2557,N_2581);
nand U3957 (N_3957,N_2320,N_2653);
and U3958 (N_3958,N_2451,N_2416);
nor U3959 (N_3959,N_2098,N_2076);
or U3960 (N_3960,N_2532,N_2595);
and U3961 (N_3961,N_2011,N_2827);
nand U3962 (N_3962,N_2732,N_2822);
nand U3963 (N_3963,N_2057,N_2994);
and U3964 (N_3964,N_2391,N_2548);
and U3965 (N_3965,N_2739,N_2485);
nand U3966 (N_3966,N_2701,N_2964);
nor U3967 (N_3967,N_2646,N_2688);
nor U3968 (N_3968,N_2879,N_2728);
nand U3969 (N_3969,N_2678,N_2471);
xor U3970 (N_3970,N_2712,N_2560);
nor U3971 (N_3971,N_2733,N_2621);
nor U3972 (N_3972,N_2064,N_2908);
nor U3973 (N_3973,N_2395,N_2303);
nand U3974 (N_3974,N_2797,N_2837);
or U3975 (N_3975,N_2961,N_2814);
and U3976 (N_3976,N_2491,N_2294);
nor U3977 (N_3977,N_2743,N_2871);
nor U3978 (N_3978,N_2672,N_2382);
and U3979 (N_3979,N_2298,N_2527);
xor U3980 (N_3980,N_2873,N_2523);
nand U3981 (N_3981,N_2416,N_2800);
or U3982 (N_3982,N_2085,N_2741);
and U3983 (N_3983,N_2009,N_2202);
nor U3984 (N_3984,N_2565,N_2198);
nor U3985 (N_3985,N_2867,N_2806);
nor U3986 (N_3986,N_2584,N_2540);
nor U3987 (N_3987,N_2312,N_2513);
nor U3988 (N_3988,N_2243,N_2828);
nand U3989 (N_3989,N_2006,N_2893);
and U3990 (N_3990,N_2963,N_2364);
and U3991 (N_3991,N_2378,N_2720);
and U3992 (N_3992,N_2272,N_2060);
or U3993 (N_3993,N_2993,N_2259);
nor U3994 (N_3994,N_2154,N_2565);
nand U3995 (N_3995,N_2785,N_2874);
nor U3996 (N_3996,N_2076,N_2840);
and U3997 (N_3997,N_2018,N_2908);
nor U3998 (N_3998,N_2597,N_2373);
nor U3999 (N_3999,N_2721,N_2017);
nand U4000 (N_4000,N_3140,N_3977);
nand U4001 (N_4001,N_3208,N_3354);
or U4002 (N_4002,N_3804,N_3382);
nand U4003 (N_4003,N_3993,N_3246);
and U4004 (N_4004,N_3723,N_3846);
and U4005 (N_4005,N_3758,N_3563);
or U4006 (N_4006,N_3111,N_3269);
and U4007 (N_4007,N_3272,N_3948);
and U4008 (N_4008,N_3837,N_3787);
or U4009 (N_4009,N_3765,N_3194);
or U4010 (N_4010,N_3964,N_3971);
nand U4011 (N_4011,N_3931,N_3090);
nor U4012 (N_4012,N_3982,N_3626);
nor U4013 (N_4013,N_3395,N_3682);
or U4014 (N_4014,N_3568,N_3475);
or U4015 (N_4015,N_3615,N_3457);
nand U4016 (N_4016,N_3887,N_3730);
xnor U4017 (N_4017,N_3679,N_3461);
nor U4018 (N_4018,N_3956,N_3227);
and U4019 (N_4019,N_3996,N_3824);
and U4020 (N_4020,N_3391,N_3707);
or U4021 (N_4021,N_3476,N_3443);
and U4022 (N_4022,N_3381,N_3703);
and U4023 (N_4023,N_3125,N_3734);
or U4024 (N_4024,N_3625,N_3132);
nor U4025 (N_4025,N_3434,N_3264);
and U4026 (N_4026,N_3712,N_3932);
nor U4027 (N_4027,N_3327,N_3583);
nor U4028 (N_4028,N_3684,N_3581);
nand U4029 (N_4029,N_3627,N_3018);
and U4030 (N_4030,N_3153,N_3023);
or U4031 (N_4031,N_3046,N_3522);
and U4032 (N_4032,N_3501,N_3812);
and U4033 (N_4033,N_3740,N_3291);
or U4034 (N_4034,N_3172,N_3429);
nand U4035 (N_4035,N_3148,N_3176);
nor U4036 (N_4036,N_3918,N_3388);
or U4037 (N_4037,N_3049,N_3845);
or U4038 (N_4038,N_3944,N_3534);
and U4039 (N_4039,N_3375,N_3916);
nor U4040 (N_4040,N_3784,N_3867);
nand U4041 (N_4041,N_3464,N_3805);
nor U4042 (N_4042,N_3618,N_3997);
and U4043 (N_4043,N_3348,N_3743);
or U4044 (N_4044,N_3753,N_3098);
nand U4045 (N_4045,N_3386,N_3197);
and U4046 (N_4046,N_3649,N_3565);
and U4047 (N_4047,N_3899,N_3135);
or U4048 (N_4048,N_3319,N_3080);
nand U4049 (N_4049,N_3667,N_3069);
or U4050 (N_4050,N_3007,N_3260);
xor U4051 (N_4051,N_3822,N_3590);
nor U4052 (N_4052,N_3187,N_3589);
and U4053 (N_4053,N_3518,N_3513);
and U4054 (N_4054,N_3092,N_3324);
nor U4055 (N_4055,N_3431,N_3751);
nand U4056 (N_4056,N_3778,N_3735);
nand U4057 (N_4057,N_3117,N_3142);
or U4058 (N_4058,N_3862,N_3481);
or U4059 (N_4059,N_3509,N_3396);
nor U4060 (N_4060,N_3575,N_3803);
and U4061 (N_4061,N_3392,N_3234);
nand U4062 (N_4062,N_3196,N_3315);
or U4063 (N_4063,N_3529,N_3584);
nand U4064 (N_4064,N_3926,N_3442);
nand U4065 (N_4065,N_3756,N_3341);
or U4066 (N_4066,N_3326,N_3219);
and U4067 (N_4067,N_3611,N_3441);
nor U4068 (N_4068,N_3598,N_3124);
and U4069 (N_4069,N_3585,N_3383);
or U4070 (N_4070,N_3953,N_3817);
nor U4071 (N_4071,N_3737,N_3314);
nand U4072 (N_4072,N_3651,N_3594);
and U4073 (N_4073,N_3550,N_3718);
or U4074 (N_4074,N_3504,N_3939);
nand U4075 (N_4075,N_3722,N_3256);
nor U4076 (N_4076,N_3379,N_3281);
nand U4077 (N_4077,N_3167,N_3890);
and U4078 (N_4078,N_3793,N_3818);
and U4079 (N_4079,N_3211,N_3795);
or U4080 (N_4080,N_3500,N_3059);
nand U4081 (N_4081,N_3791,N_3448);
or U4082 (N_4082,N_3545,N_3232);
and U4083 (N_4083,N_3782,N_3498);
nor U4084 (N_4084,N_3493,N_3366);
nand U4085 (N_4085,N_3826,N_3012);
or U4086 (N_4086,N_3733,N_3732);
or U4087 (N_4087,N_3571,N_3278);
or U4088 (N_4088,N_3162,N_3631);
nor U4089 (N_4089,N_3605,N_3008);
nor U4090 (N_4090,N_3928,N_3151);
or U4091 (N_4091,N_3149,N_3970);
nor U4092 (N_4092,N_3489,N_3749);
nand U4093 (N_4093,N_3164,N_3917);
nand U4094 (N_4094,N_3108,N_3295);
or U4095 (N_4095,N_3469,N_3159);
or U4096 (N_4096,N_3335,N_3236);
nand U4097 (N_4097,N_3548,N_3178);
and U4098 (N_4098,N_3633,N_3171);
nand U4099 (N_4099,N_3599,N_3919);
and U4100 (N_4100,N_3901,N_3898);
nor U4101 (N_4101,N_3138,N_3698);
and U4102 (N_4102,N_3497,N_3025);
and U4103 (N_4103,N_3222,N_3864);
nand U4104 (N_4104,N_3405,N_3847);
and U4105 (N_4105,N_3305,N_3933);
nor U4106 (N_4106,N_3680,N_3639);
or U4107 (N_4107,N_3681,N_3658);
or U4108 (N_4108,N_3569,N_3853);
or U4109 (N_4109,N_3717,N_3607);
nor U4110 (N_4110,N_3225,N_3249);
or U4111 (N_4111,N_3774,N_3367);
nor U4112 (N_4112,N_3202,N_3426);
and U4113 (N_4113,N_3022,N_3959);
nor U4114 (N_4114,N_3700,N_3419);
and U4115 (N_4115,N_3346,N_3988);
and U4116 (N_4116,N_3073,N_3378);
and U4117 (N_4117,N_3248,N_3000);
or U4118 (N_4118,N_3713,N_3866);
or U4119 (N_4119,N_3075,N_3237);
nor U4120 (N_4120,N_3850,N_3458);
nor U4121 (N_4121,N_3333,N_3685);
and U4122 (N_4122,N_3216,N_3965);
or U4123 (N_4123,N_3129,N_3871);
nor U4124 (N_4124,N_3384,N_3438);
or U4125 (N_4125,N_3861,N_3994);
and U4126 (N_4126,N_3277,N_3353);
or U4127 (N_4127,N_3958,N_3621);
and U4128 (N_4128,N_3413,N_3851);
and U4129 (N_4129,N_3825,N_3728);
or U4130 (N_4130,N_3056,N_3455);
or U4131 (N_4131,N_3173,N_3582);
and U4132 (N_4132,N_3990,N_3478);
nand U4133 (N_4133,N_3473,N_3293);
nand U4134 (N_4134,N_3537,N_3244);
or U4135 (N_4135,N_3286,N_3935);
or U4136 (N_4136,N_3450,N_3838);
nor U4137 (N_4137,N_3533,N_3863);
nand U4138 (N_4138,N_3891,N_3711);
or U4139 (N_4139,N_3066,N_3636);
nand U4140 (N_4140,N_3699,N_3035);
and U4141 (N_4141,N_3224,N_3811);
nor U4142 (N_4142,N_3266,N_3910);
or U4143 (N_4143,N_3859,N_3528);
nor U4144 (N_4144,N_3350,N_3430);
nor U4145 (N_4145,N_3016,N_3688);
and U4146 (N_4146,N_3666,N_3609);
nor U4147 (N_4147,N_3045,N_3296);
nand U4148 (N_4148,N_3542,N_3253);
xnor U4149 (N_4149,N_3654,N_3963);
nor U4150 (N_4150,N_3978,N_3297);
or U4151 (N_4151,N_3562,N_3676);
and U4152 (N_4152,N_3947,N_3109);
or U4153 (N_4153,N_3410,N_3815);
nor U4154 (N_4154,N_3245,N_3759);
and U4155 (N_4155,N_3689,N_3033);
nand U4156 (N_4156,N_3198,N_3002);
or U4157 (N_4157,N_3029,N_3868);
and U4158 (N_4158,N_3058,N_3706);
nand U4159 (N_4159,N_3084,N_3468);
or U4160 (N_4160,N_3349,N_3945);
and U4161 (N_4161,N_3601,N_3054);
or U4162 (N_4162,N_3792,N_3628);
or U4163 (N_4163,N_3215,N_3311);
and U4164 (N_4164,N_3100,N_3201);
nand U4165 (N_4165,N_3067,N_3347);
nand U4166 (N_4166,N_3377,N_3229);
and U4167 (N_4167,N_3189,N_3247);
nand U4168 (N_4168,N_3083,N_3492);
or U4169 (N_4169,N_3702,N_3114);
or U4170 (N_4170,N_3320,N_3042);
or U4171 (N_4171,N_3781,N_3608);
nand U4172 (N_4172,N_3727,N_3950);
nand U4173 (N_4173,N_3870,N_3554);
nand U4174 (N_4174,N_3188,N_3652);
nand U4175 (N_4175,N_3827,N_3401);
nand U4176 (N_4176,N_3725,N_3486);
nor U4177 (N_4177,N_3263,N_3465);
or U4178 (N_4178,N_3112,N_3337);
or U4179 (N_4179,N_3516,N_3449);
nor U4180 (N_4180,N_3421,N_3339);
nor U4181 (N_4181,N_3287,N_3510);
and U4182 (N_4182,N_3640,N_3009);
or U4183 (N_4183,N_3034,N_3619);
and U4184 (N_4184,N_3436,N_3664);
xnor U4185 (N_4185,N_3409,N_3252);
nand U4186 (N_4186,N_3356,N_3484);
nand U4187 (N_4187,N_3397,N_3612);
nor U4188 (N_4188,N_3404,N_3549);
or U4189 (N_4189,N_3610,N_3031);
nand U4190 (N_4190,N_3437,N_3788);
and U4191 (N_4191,N_3318,N_3446);
nor U4192 (N_4192,N_3230,N_3217);
or U4193 (N_4193,N_3491,N_3243);
nor U4194 (N_4194,N_3139,N_3980);
and U4195 (N_4195,N_3313,N_3301);
and U4196 (N_4196,N_3720,N_3331);
nor U4197 (N_4197,N_3808,N_3488);
or U4198 (N_4198,N_3573,N_3721);
or U4199 (N_4199,N_3686,N_3168);
nand U4200 (N_4200,N_3329,N_3370);
nor U4201 (N_4201,N_3250,N_3041);
and U4202 (N_4202,N_3694,N_3422);
or U4203 (N_4203,N_3677,N_3163);
or U4204 (N_4204,N_3538,N_3906);
nand U4205 (N_4205,N_3072,N_3028);
nand U4206 (N_4206,N_3960,N_3647);
or U4207 (N_4207,N_3102,N_3907);
or U4208 (N_4208,N_3223,N_3360);
nand U4209 (N_4209,N_3466,N_3883);
or U4210 (N_4210,N_3143,N_3472);
or U4211 (N_4211,N_3494,N_3527);
nor U4212 (N_4212,N_3981,N_3574);
nand U4213 (N_4213,N_3506,N_3558);
and U4214 (N_4214,N_3719,N_3536);
nand U4215 (N_4215,N_3043,N_3453);
nand U4216 (N_4216,N_3943,N_3844);
nor U4217 (N_4217,N_3284,N_3869);
and U4218 (N_4218,N_3524,N_3519);
or U4219 (N_4219,N_3181,N_3662);
nor U4220 (N_4220,N_3641,N_3695);
nand U4221 (N_4221,N_3136,N_3710);
nor U4222 (N_4222,N_3690,N_3412);
nand U4223 (N_4223,N_3345,N_3439);
nor U4224 (N_4224,N_3929,N_3755);
nor U4225 (N_4225,N_3570,N_3340);
and U4226 (N_4226,N_3687,N_3860);
or U4227 (N_4227,N_3507,N_3130);
and U4228 (N_4228,N_3579,N_3802);
nand U4229 (N_4229,N_3423,N_3128);
nor U4230 (N_4230,N_3062,N_3220);
and U4231 (N_4231,N_3499,N_3955);
xnor U4232 (N_4232,N_3203,N_3362);
nor U4233 (N_4233,N_3294,N_3177);
nand U4234 (N_4234,N_3540,N_3146);
or U4235 (N_4235,N_3357,N_3338);
or U4236 (N_4236,N_3544,N_3828);
and U4237 (N_4237,N_3769,N_3359);
or U4238 (N_4238,N_3897,N_3195);
nor U4239 (N_4239,N_3592,N_3637);
and U4240 (N_4240,N_3772,N_3814);
or U4241 (N_4241,N_3076,N_3079);
nand U4242 (N_4242,N_3986,N_3060);
nor U4243 (N_4243,N_3400,N_3038);
and U4244 (N_4244,N_3752,N_3741);
and U4245 (N_4245,N_3071,N_3303);
nor U4246 (N_4246,N_3704,N_3954);
nand U4247 (N_4247,N_3322,N_3192);
nand U4248 (N_4248,N_3089,N_3334);
and U4249 (N_4249,N_3632,N_3403);
and U4250 (N_4250,N_3279,N_3290);
nor U4251 (N_4251,N_3806,N_3231);
or U4252 (N_4252,N_3646,N_3014);
and U4253 (N_4253,N_3643,N_3675);
or U4254 (N_4254,N_3044,N_3113);
nor U4255 (N_4255,N_3952,N_3179);
nor U4256 (N_4256,N_3979,N_3801);
nand U4257 (N_4257,N_3270,N_3505);
nor U4258 (N_4258,N_3880,N_3670);
and U4259 (N_4259,N_3665,N_3004);
or U4260 (N_4260,N_3921,N_3376);
nor U4261 (N_4261,N_3145,N_3927);
or U4262 (N_4262,N_3739,N_3744);
nor U4263 (N_4263,N_3766,N_3776);
nand U4264 (N_4264,N_3039,N_3040);
or U4265 (N_4265,N_3526,N_3551);
nand U4266 (N_4266,N_3726,N_3399);
or U4267 (N_4267,N_3030,N_3914);
and U4268 (N_4268,N_3560,N_3393);
and U4269 (N_4269,N_3515,N_3839);
or U4270 (N_4270,N_3555,N_3051);
xnor U4271 (N_4271,N_3779,N_3158);
nand U4272 (N_4272,N_3483,N_3474);
and U4273 (N_4273,N_3693,N_3156);
nor U4274 (N_4274,N_3174,N_3622);
and U4275 (N_4275,N_3794,N_3973);
nor U4276 (N_4276,N_3332,N_3175);
nand U4277 (N_4277,N_3521,N_3411);
or U4278 (N_4278,N_3099,N_3026);
xor U4279 (N_4279,N_3904,N_3487);
nand U4280 (N_4280,N_3729,N_3613);
and U4281 (N_4281,N_3559,N_3255);
nand U4282 (N_4282,N_3161,N_3127);
nor U4283 (N_4283,N_3104,N_3095);
nor U4284 (N_4284,N_3508,N_3541);
and U4285 (N_4285,N_3561,N_3661);
nor U4286 (N_4286,N_3152,N_3205);
nor U4287 (N_4287,N_3330,N_3742);
and U4288 (N_4288,N_3961,N_3616);
nor U4289 (N_4289,N_3900,N_3432);
nor U4290 (N_4290,N_3586,N_3226);
or U4291 (N_4291,N_3819,N_3701);
nand U4292 (N_4292,N_3660,N_3941);
and U4293 (N_4293,N_3160,N_3325);
nor U4294 (N_4294,N_3088,N_3836);
nor U4295 (N_4295,N_3275,N_3995);
nand U4296 (N_4296,N_3876,N_3134);
and U4297 (N_4297,N_3539,N_3015);
or U4298 (N_4298,N_3180,N_3514);
or U4299 (N_4299,N_3480,N_3663);
and U4300 (N_4300,N_3922,N_3656);
nor U4301 (N_4301,N_3520,N_3417);
nand U4302 (N_4302,N_3240,N_3271);
nor U4303 (N_4303,N_3934,N_3708);
or U4304 (N_4304,N_3209,N_3445);
nor U4305 (N_4305,N_3485,N_3343);
and U4306 (N_4306,N_3535,N_3849);
and U4307 (N_4307,N_3428,N_3617);
nor U4308 (N_4308,N_3830,N_3942);
nand U4309 (N_4309,N_3107,N_3094);
and U4310 (N_4310,N_3987,N_3920);
or U4311 (N_4311,N_3886,N_3967);
and U4312 (N_4312,N_3074,N_3047);
or U4313 (N_4313,N_3697,N_3052);
and U4314 (N_4314,N_3714,N_3502);
xor U4315 (N_4315,N_3451,N_3895);
nor U4316 (N_4316,N_3757,N_3169);
and U4317 (N_4317,N_3241,N_3050);
and U4318 (N_4318,N_3800,N_3055);
nand U4319 (N_4319,N_3604,N_3414);
or U4320 (N_4320,N_3593,N_3358);
nand U4321 (N_4321,N_3238,N_3829);
or U4322 (N_4322,N_3771,N_3302);
and U4323 (N_4323,N_3523,N_3003);
and U4324 (N_4324,N_3150,N_3299);
nand U4325 (N_4325,N_3655,N_3207);
nand U4326 (N_4326,N_3764,N_3328);
nor U4327 (N_4327,N_3760,N_3634);
nand U4328 (N_4328,N_3402,N_3966);
nand U4329 (N_4329,N_3091,N_3011);
or U4330 (N_4330,N_3783,N_3832);
nand U4331 (N_4331,N_3915,N_3444);
nand U4332 (N_4332,N_3239,N_3893);
or U4333 (N_4333,N_3036,N_3731);
and U4334 (N_4334,N_3857,N_3261);
and U4335 (N_4335,N_3930,N_3892);
nand U4336 (N_4336,N_3972,N_3603);
nor U4337 (N_4337,N_3085,N_3191);
nor U4338 (N_4338,N_3736,N_3659);
or U4339 (N_4339,N_3137,N_3233);
and U4340 (N_4340,N_3490,N_3775);
or U4341 (N_4341,N_3365,N_3877);
and U4342 (N_4342,N_3093,N_3975);
or U4343 (N_4343,N_3543,N_3495);
or U4344 (N_4344,N_3452,N_3267);
or U4345 (N_4345,N_3553,N_3283);
and U4346 (N_4346,N_3602,N_3983);
nor U4347 (N_4347,N_3144,N_3065);
and U4348 (N_4348,N_3323,N_3373);
nand U4349 (N_4349,N_3447,N_3309);
nand U4350 (N_4350,N_3556,N_3768);
and U4351 (N_4351,N_3304,N_3912);
nor U4352 (N_4352,N_3407,N_3874);
nor U4353 (N_4353,N_3566,N_3511);
or U4354 (N_4354,N_3116,N_3576);
and U4355 (N_4355,N_3678,N_3342);
and U4356 (N_4356,N_3767,N_3355);
nand U4357 (N_4357,N_3282,N_3268);
or U4358 (N_4358,N_3923,N_3259);
or U4359 (N_4359,N_3463,N_3110);
nor U4360 (N_4360,N_3336,N_3848);
and U4361 (N_4361,N_3770,N_3858);
nand U4362 (N_4362,N_3154,N_3258);
or U4363 (N_4363,N_3816,N_3389);
and U4364 (N_4364,N_3894,N_3369);
and U4365 (N_4365,N_3200,N_3385);
nand U4366 (N_4366,N_3213,N_3024);
nand U4367 (N_4367,N_3969,N_3242);
and U4368 (N_4368,N_3597,N_3840);
or U4369 (N_4369,N_3668,N_3097);
nand U4370 (N_4370,N_3087,N_3754);
nand U4371 (N_4371,N_3937,N_3620);
or U4372 (N_4372,N_3673,N_3101);
nand U4373 (N_4373,N_3063,N_3810);
and U4374 (N_4374,N_3418,N_3118);
nand U4375 (N_4375,N_3962,N_3193);
or U4376 (N_4376,N_3946,N_3186);
and U4377 (N_4377,N_3856,N_3440);
or U4378 (N_4378,N_3517,N_3773);
and U4379 (N_4379,N_3408,N_3019);
and U4380 (N_4380,N_3459,N_3913);
and U4381 (N_4381,N_3477,N_3021);
nor U4382 (N_4382,N_3165,N_3057);
nand U4383 (N_4383,N_3155,N_3999);
and U4384 (N_4384,N_3635,N_3985);
and U4385 (N_4385,N_3882,N_3317);
nor U4386 (N_4386,N_3471,N_3361);
nor U4387 (N_4387,N_3068,N_3889);
nor U4388 (N_4388,N_3235,N_3798);
nor U4389 (N_4389,N_3218,N_3709);
and U4390 (N_4390,N_3761,N_3027);
nand U4391 (N_4391,N_3909,N_3600);
and U4392 (N_4392,N_3671,N_3885);
and U4393 (N_4393,N_3064,N_3131);
and U4394 (N_4394,N_3300,N_3949);
or U4395 (N_4395,N_3745,N_3017);
nand U4396 (N_4396,N_3435,N_3276);
or U4397 (N_4397,N_3228,N_3307);
or U4398 (N_4398,N_3119,N_3976);
and U4399 (N_4399,N_3053,N_3790);
nor U4400 (N_4400,N_3061,N_3936);
and U4401 (N_4401,N_3121,N_3762);
and U4402 (N_4402,N_3298,N_3274);
and U4403 (N_4403,N_3624,N_3462);
nor U4404 (N_4404,N_3683,N_3420);
and U4405 (N_4405,N_3479,N_3968);
or U4406 (N_4406,N_3878,N_3273);
nor U4407 (N_4407,N_3390,N_3105);
and U4408 (N_4408,N_3292,N_3564);
and U4409 (N_4409,N_3873,N_3896);
nand U4410 (N_4410,N_3210,N_3081);
and U4411 (N_4411,N_3394,N_3424);
or U4412 (N_4412,N_3746,N_3813);
and U4413 (N_4413,N_3833,N_3842);
nand U4414 (N_4414,N_3289,N_3789);
nand U4415 (N_4415,N_3454,N_3831);
nand U4416 (N_4416,N_3696,N_3750);
nor U4417 (N_4417,N_3123,N_3908);
or U4418 (N_4418,N_3316,N_3374);
nor U4419 (N_4419,N_3120,N_3991);
or U4420 (N_4420,N_3221,N_3070);
and U4421 (N_4421,N_3799,N_3310);
nor U4422 (N_4422,N_3747,N_3588);
or U4423 (N_4423,N_3005,N_3855);
and U4424 (N_4424,N_3823,N_3372);
or U4425 (N_4425,N_3780,N_3427);
and U4426 (N_4426,N_3482,N_3881);
and U4427 (N_4427,N_3648,N_3580);
nor U4428 (N_4428,N_3470,N_3925);
and U4429 (N_4429,N_3371,N_3503);
nand U4430 (N_4430,N_3199,N_3777);
and U4431 (N_4431,N_3763,N_3531);
and U4432 (N_4432,N_3530,N_3352);
and U4433 (N_4433,N_3786,N_3126);
nand U4434 (N_4434,N_3578,N_3037);
and U4435 (N_4435,N_3425,N_3077);
and U4436 (N_4436,N_3032,N_3546);
or U4437 (N_4437,N_3204,N_3957);
and U4438 (N_4438,N_3020,N_3496);
and U4439 (N_4439,N_3285,N_3312);
nand U4440 (N_4440,N_3623,N_3001);
and U4441 (N_4441,N_3595,N_3596);
nor U4442 (N_4442,N_3190,N_3872);
nor U4443 (N_4443,N_3879,N_3865);
nand U4444 (N_4444,N_3629,N_3748);
nor U4445 (N_4445,N_3809,N_3460);
nor U4446 (N_4446,N_3415,N_3467);
xnor U4447 (N_4447,N_3854,N_3938);
nand U4448 (N_4448,N_3852,N_3013);
or U4449 (N_4449,N_3096,N_3398);
nor U4450 (N_4450,N_3433,N_3416);
and U4451 (N_4451,N_3653,N_3905);
nor U4452 (N_4452,N_3724,N_3078);
or U4453 (N_4453,N_3716,N_3841);
or U4454 (N_4454,N_3525,N_3974);
nor U4455 (N_4455,N_3406,N_3606);
nand U4456 (N_4456,N_3321,N_3821);
and U4457 (N_4457,N_3984,N_3257);
or U4458 (N_4458,N_3262,N_3797);
nand U4459 (N_4459,N_3715,N_3835);
or U4460 (N_4460,N_3820,N_3182);
or U4461 (N_4461,N_3884,N_3567);
nand U4462 (N_4462,N_3992,N_3785);
and U4463 (N_4463,N_3115,N_3368);
nor U4464 (N_4464,N_3456,N_3380);
xnor U4465 (N_4465,N_3364,N_3552);
nand U4466 (N_4466,N_3206,N_3642);
and U4467 (N_4467,N_3630,N_3572);
or U4468 (N_4468,N_3924,N_3644);
and U4469 (N_4469,N_3587,N_3989);
or U4470 (N_4470,N_3157,N_3103);
xor U4471 (N_4471,N_3254,N_3577);
or U4472 (N_4472,N_3265,N_3387);
and U4473 (N_4473,N_3591,N_3669);
nand U4474 (N_4474,N_3657,N_3951);
and U4475 (N_4475,N_3512,N_3214);
nor U4476 (N_4476,N_3911,N_3166);
nor U4477 (N_4477,N_3796,N_3006);
and U4478 (N_4478,N_3363,N_3557);
and U4479 (N_4479,N_3738,N_3692);
nor U4480 (N_4480,N_3705,N_3834);
nor U4481 (N_4481,N_3183,N_3638);
nand U4482 (N_4482,N_3888,N_3902);
nand U4483 (N_4483,N_3547,N_3185);
nor U4484 (N_4484,N_3308,N_3048);
nor U4485 (N_4485,N_3106,N_3672);
nand U4486 (N_4486,N_3691,N_3170);
nor U4487 (N_4487,N_3843,N_3532);
and U4488 (N_4488,N_3998,N_3614);
nor U4489 (N_4489,N_3212,N_3344);
and U4490 (N_4490,N_3133,N_3807);
and U4491 (N_4491,N_3650,N_3875);
or U4492 (N_4492,N_3082,N_3903);
or U4493 (N_4493,N_3288,N_3010);
nand U4494 (N_4494,N_3141,N_3351);
and U4495 (N_4495,N_3645,N_3674);
nand U4496 (N_4496,N_3940,N_3122);
and U4497 (N_4497,N_3147,N_3184);
nor U4498 (N_4498,N_3086,N_3280);
nand U4499 (N_4499,N_3306,N_3251);
nand U4500 (N_4500,N_3402,N_3083);
and U4501 (N_4501,N_3642,N_3749);
and U4502 (N_4502,N_3484,N_3131);
nor U4503 (N_4503,N_3150,N_3612);
or U4504 (N_4504,N_3941,N_3837);
nor U4505 (N_4505,N_3291,N_3060);
nand U4506 (N_4506,N_3845,N_3378);
nand U4507 (N_4507,N_3593,N_3383);
and U4508 (N_4508,N_3695,N_3050);
and U4509 (N_4509,N_3270,N_3308);
nor U4510 (N_4510,N_3050,N_3129);
nor U4511 (N_4511,N_3979,N_3278);
and U4512 (N_4512,N_3365,N_3795);
or U4513 (N_4513,N_3597,N_3712);
or U4514 (N_4514,N_3367,N_3447);
or U4515 (N_4515,N_3910,N_3166);
nand U4516 (N_4516,N_3268,N_3664);
nor U4517 (N_4517,N_3670,N_3527);
or U4518 (N_4518,N_3346,N_3401);
xor U4519 (N_4519,N_3371,N_3045);
and U4520 (N_4520,N_3469,N_3840);
or U4521 (N_4521,N_3389,N_3979);
nor U4522 (N_4522,N_3636,N_3114);
and U4523 (N_4523,N_3724,N_3338);
nand U4524 (N_4524,N_3701,N_3025);
or U4525 (N_4525,N_3286,N_3983);
and U4526 (N_4526,N_3900,N_3385);
nand U4527 (N_4527,N_3959,N_3526);
and U4528 (N_4528,N_3950,N_3445);
or U4529 (N_4529,N_3484,N_3809);
nor U4530 (N_4530,N_3202,N_3720);
or U4531 (N_4531,N_3319,N_3512);
and U4532 (N_4532,N_3091,N_3155);
and U4533 (N_4533,N_3519,N_3223);
nand U4534 (N_4534,N_3433,N_3674);
nand U4535 (N_4535,N_3782,N_3473);
or U4536 (N_4536,N_3727,N_3290);
nor U4537 (N_4537,N_3754,N_3140);
or U4538 (N_4538,N_3013,N_3083);
nor U4539 (N_4539,N_3940,N_3091);
nor U4540 (N_4540,N_3594,N_3939);
nor U4541 (N_4541,N_3253,N_3663);
or U4542 (N_4542,N_3669,N_3965);
nor U4543 (N_4543,N_3343,N_3705);
nor U4544 (N_4544,N_3047,N_3596);
nand U4545 (N_4545,N_3508,N_3964);
and U4546 (N_4546,N_3041,N_3007);
or U4547 (N_4547,N_3625,N_3930);
or U4548 (N_4548,N_3769,N_3351);
and U4549 (N_4549,N_3570,N_3555);
nand U4550 (N_4550,N_3679,N_3551);
nand U4551 (N_4551,N_3262,N_3090);
nor U4552 (N_4552,N_3426,N_3086);
nand U4553 (N_4553,N_3419,N_3878);
or U4554 (N_4554,N_3671,N_3981);
and U4555 (N_4555,N_3385,N_3322);
nand U4556 (N_4556,N_3351,N_3607);
nor U4557 (N_4557,N_3174,N_3844);
or U4558 (N_4558,N_3174,N_3697);
nand U4559 (N_4559,N_3650,N_3816);
nand U4560 (N_4560,N_3406,N_3535);
and U4561 (N_4561,N_3147,N_3252);
and U4562 (N_4562,N_3842,N_3259);
nor U4563 (N_4563,N_3319,N_3310);
nand U4564 (N_4564,N_3389,N_3013);
and U4565 (N_4565,N_3816,N_3745);
nor U4566 (N_4566,N_3516,N_3961);
xor U4567 (N_4567,N_3536,N_3435);
or U4568 (N_4568,N_3940,N_3934);
nand U4569 (N_4569,N_3077,N_3293);
xnor U4570 (N_4570,N_3168,N_3953);
nor U4571 (N_4571,N_3136,N_3592);
and U4572 (N_4572,N_3584,N_3897);
nor U4573 (N_4573,N_3498,N_3287);
and U4574 (N_4574,N_3709,N_3922);
or U4575 (N_4575,N_3838,N_3711);
nand U4576 (N_4576,N_3243,N_3907);
nor U4577 (N_4577,N_3018,N_3738);
nand U4578 (N_4578,N_3819,N_3078);
nor U4579 (N_4579,N_3242,N_3754);
nand U4580 (N_4580,N_3282,N_3541);
nand U4581 (N_4581,N_3301,N_3191);
nand U4582 (N_4582,N_3173,N_3610);
nand U4583 (N_4583,N_3830,N_3046);
or U4584 (N_4584,N_3421,N_3433);
nor U4585 (N_4585,N_3517,N_3089);
or U4586 (N_4586,N_3048,N_3152);
and U4587 (N_4587,N_3991,N_3834);
nand U4588 (N_4588,N_3134,N_3774);
nand U4589 (N_4589,N_3317,N_3952);
and U4590 (N_4590,N_3061,N_3543);
nor U4591 (N_4591,N_3023,N_3858);
or U4592 (N_4592,N_3684,N_3269);
nor U4593 (N_4593,N_3283,N_3562);
or U4594 (N_4594,N_3336,N_3403);
nor U4595 (N_4595,N_3354,N_3353);
and U4596 (N_4596,N_3047,N_3466);
nor U4597 (N_4597,N_3301,N_3143);
or U4598 (N_4598,N_3071,N_3301);
or U4599 (N_4599,N_3245,N_3008);
and U4600 (N_4600,N_3421,N_3013);
nand U4601 (N_4601,N_3877,N_3300);
or U4602 (N_4602,N_3037,N_3558);
or U4603 (N_4603,N_3297,N_3179);
or U4604 (N_4604,N_3350,N_3848);
nand U4605 (N_4605,N_3401,N_3525);
and U4606 (N_4606,N_3584,N_3456);
nand U4607 (N_4607,N_3734,N_3655);
and U4608 (N_4608,N_3047,N_3621);
or U4609 (N_4609,N_3758,N_3479);
nor U4610 (N_4610,N_3275,N_3656);
nor U4611 (N_4611,N_3687,N_3419);
or U4612 (N_4612,N_3177,N_3009);
nand U4613 (N_4613,N_3313,N_3007);
nand U4614 (N_4614,N_3104,N_3328);
nor U4615 (N_4615,N_3396,N_3613);
or U4616 (N_4616,N_3369,N_3979);
nor U4617 (N_4617,N_3625,N_3326);
nor U4618 (N_4618,N_3608,N_3949);
and U4619 (N_4619,N_3709,N_3952);
and U4620 (N_4620,N_3681,N_3019);
or U4621 (N_4621,N_3509,N_3680);
nand U4622 (N_4622,N_3367,N_3943);
nor U4623 (N_4623,N_3161,N_3495);
nand U4624 (N_4624,N_3007,N_3075);
and U4625 (N_4625,N_3032,N_3641);
and U4626 (N_4626,N_3462,N_3278);
nand U4627 (N_4627,N_3711,N_3285);
and U4628 (N_4628,N_3496,N_3300);
or U4629 (N_4629,N_3287,N_3107);
or U4630 (N_4630,N_3372,N_3532);
and U4631 (N_4631,N_3690,N_3960);
nor U4632 (N_4632,N_3053,N_3460);
nand U4633 (N_4633,N_3367,N_3995);
nand U4634 (N_4634,N_3989,N_3190);
or U4635 (N_4635,N_3236,N_3379);
and U4636 (N_4636,N_3028,N_3731);
nand U4637 (N_4637,N_3425,N_3655);
nand U4638 (N_4638,N_3188,N_3340);
or U4639 (N_4639,N_3690,N_3492);
or U4640 (N_4640,N_3079,N_3970);
nand U4641 (N_4641,N_3043,N_3614);
or U4642 (N_4642,N_3779,N_3145);
xnor U4643 (N_4643,N_3366,N_3705);
nor U4644 (N_4644,N_3692,N_3349);
and U4645 (N_4645,N_3018,N_3607);
nor U4646 (N_4646,N_3197,N_3590);
or U4647 (N_4647,N_3563,N_3128);
nand U4648 (N_4648,N_3640,N_3150);
and U4649 (N_4649,N_3539,N_3082);
or U4650 (N_4650,N_3432,N_3970);
or U4651 (N_4651,N_3603,N_3636);
nand U4652 (N_4652,N_3559,N_3162);
nor U4653 (N_4653,N_3489,N_3540);
and U4654 (N_4654,N_3010,N_3336);
nor U4655 (N_4655,N_3704,N_3712);
or U4656 (N_4656,N_3492,N_3485);
nand U4657 (N_4657,N_3727,N_3209);
or U4658 (N_4658,N_3032,N_3055);
nand U4659 (N_4659,N_3661,N_3014);
and U4660 (N_4660,N_3822,N_3805);
nand U4661 (N_4661,N_3902,N_3556);
or U4662 (N_4662,N_3214,N_3788);
nor U4663 (N_4663,N_3078,N_3648);
or U4664 (N_4664,N_3463,N_3718);
nand U4665 (N_4665,N_3983,N_3748);
and U4666 (N_4666,N_3492,N_3160);
and U4667 (N_4667,N_3970,N_3512);
and U4668 (N_4668,N_3246,N_3196);
nor U4669 (N_4669,N_3168,N_3535);
and U4670 (N_4670,N_3655,N_3193);
and U4671 (N_4671,N_3581,N_3412);
nand U4672 (N_4672,N_3864,N_3391);
nor U4673 (N_4673,N_3629,N_3092);
and U4674 (N_4674,N_3176,N_3425);
or U4675 (N_4675,N_3336,N_3327);
and U4676 (N_4676,N_3427,N_3339);
and U4677 (N_4677,N_3761,N_3976);
nor U4678 (N_4678,N_3793,N_3707);
nand U4679 (N_4679,N_3281,N_3678);
nand U4680 (N_4680,N_3442,N_3311);
nand U4681 (N_4681,N_3516,N_3708);
nor U4682 (N_4682,N_3379,N_3859);
nor U4683 (N_4683,N_3930,N_3840);
and U4684 (N_4684,N_3779,N_3913);
and U4685 (N_4685,N_3206,N_3783);
nor U4686 (N_4686,N_3242,N_3407);
nand U4687 (N_4687,N_3302,N_3677);
nor U4688 (N_4688,N_3047,N_3303);
or U4689 (N_4689,N_3418,N_3475);
nor U4690 (N_4690,N_3169,N_3529);
nand U4691 (N_4691,N_3257,N_3606);
nor U4692 (N_4692,N_3795,N_3298);
and U4693 (N_4693,N_3900,N_3642);
and U4694 (N_4694,N_3916,N_3530);
nor U4695 (N_4695,N_3118,N_3401);
or U4696 (N_4696,N_3250,N_3660);
and U4697 (N_4697,N_3370,N_3384);
or U4698 (N_4698,N_3237,N_3024);
or U4699 (N_4699,N_3986,N_3133);
nand U4700 (N_4700,N_3971,N_3980);
nand U4701 (N_4701,N_3868,N_3534);
and U4702 (N_4702,N_3436,N_3030);
nor U4703 (N_4703,N_3218,N_3065);
or U4704 (N_4704,N_3951,N_3443);
nor U4705 (N_4705,N_3841,N_3359);
or U4706 (N_4706,N_3662,N_3585);
nand U4707 (N_4707,N_3396,N_3297);
or U4708 (N_4708,N_3498,N_3173);
nand U4709 (N_4709,N_3452,N_3610);
or U4710 (N_4710,N_3609,N_3620);
nor U4711 (N_4711,N_3691,N_3845);
nor U4712 (N_4712,N_3816,N_3400);
or U4713 (N_4713,N_3313,N_3824);
nor U4714 (N_4714,N_3525,N_3556);
nand U4715 (N_4715,N_3328,N_3068);
nand U4716 (N_4716,N_3745,N_3149);
nand U4717 (N_4717,N_3898,N_3142);
nand U4718 (N_4718,N_3289,N_3317);
nor U4719 (N_4719,N_3285,N_3813);
nand U4720 (N_4720,N_3594,N_3426);
nand U4721 (N_4721,N_3822,N_3119);
nor U4722 (N_4722,N_3740,N_3478);
nor U4723 (N_4723,N_3864,N_3418);
nand U4724 (N_4724,N_3866,N_3213);
nor U4725 (N_4725,N_3644,N_3303);
nor U4726 (N_4726,N_3887,N_3113);
nand U4727 (N_4727,N_3401,N_3385);
or U4728 (N_4728,N_3851,N_3167);
nor U4729 (N_4729,N_3913,N_3673);
and U4730 (N_4730,N_3915,N_3470);
nand U4731 (N_4731,N_3145,N_3516);
or U4732 (N_4732,N_3802,N_3785);
or U4733 (N_4733,N_3396,N_3944);
nor U4734 (N_4734,N_3011,N_3253);
nor U4735 (N_4735,N_3301,N_3338);
nand U4736 (N_4736,N_3751,N_3839);
nand U4737 (N_4737,N_3244,N_3915);
nor U4738 (N_4738,N_3094,N_3720);
or U4739 (N_4739,N_3105,N_3694);
nor U4740 (N_4740,N_3365,N_3549);
nand U4741 (N_4741,N_3201,N_3356);
nand U4742 (N_4742,N_3442,N_3872);
and U4743 (N_4743,N_3216,N_3118);
or U4744 (N_4744,N_3177,N_3216);
and U4745 (N_4745,N_3621,N_3439);
or U4746 (N_4746,N_3334,N_3243);
nor U4747 (N_4747,N_3916,N_3514);
nor U4748 (N_4748,N_3856,N_3506);
and U4749 (N_4749,N_3736,N_3727);
and U4750 (N_4750,N_3315,N_3633);
or U4751 (N_4751,N_3572,N_3390);
nand U4752 (N_4752,N_3106,N_3957);
nand U4753 (N_4753,N_3108,N_3466);
and U4754 (N_4754,N_3255,N_3962);
and U4755 (N_4755,N_3707,N_3014);
nand U4756 (N_4756,N_3972,N_3709);
nand U4757 (N_4757,N_3798,N_3677);
nand U4758 (N_4758,N_3305,N_3844);
nand U4759 (N_4759,N_3340,N_3225);
and U4760 (N_4760,N_3811,N_3469);
nor U4761 (N_4761,N_3499,N_3449);
nor U4762 (N_4762,N_3389,N_3878);
or U4763 (N_4763,N_3168,N_3042);
and U4764 (N_4764,N_3952,N_3369);
nor U4765 (N_4765,N_3917,N_3069);
nand U4766 (N_4766,N_3149,N_3873);
and U4767 (N_4767,N_3676,N_3178);
nand U4768 (N_4768,N_3168,N_3882);
nor U4769 (N_4769,N_3432,N_3732);
or U4770 (N_4770,N_3490,N_3171);
or U4771 (N_4771,N_3466,N_3028);
nand U4772 (N_4772,N_3575,N_3944);
or U4773 (N_4773,N_3887,N_3897);
nor U4774 (N_4774,N_3101,N_3645);
nand U4775 (N_4775,N_3454,N_3914);
nand U4776 (N_4776,N_3882,N_3803);
nor U4777 (N_4777,N_3619,N_3408);
and U4778 (N_4778,N_3733,N_3503);
or U4779 (N_4779,N_3526,N_3686);
and U4780 (N_4780,N_3435,N_3203);
and U4781 (N_4781,N_3338,N_3655);
and U4782 (N_4782,N_3039,N_3378);
nand U4783 (N_4783,N_3489,N_3611);
xnor U4784 (N_4784,N_3681,N_3514);
and U4785 (N_4785,N_3933,N_3543);
or U4786 (N_4786,N_3173,N_3350);
or U4787 (N_4787,N_3827,N_3566);
and U4788 (N_4788,N_3010,N_3625);
nor U4789 (N_4789,N_3896,N_3751);
or U4790 (N_4790,N_3907,N_3457);
xor U4791 (N_4791,N_3843,N_3876);
and U4792 (N_4792,N_3092,N_3979);
nor U4793 (N_4793,N_3958,N_3486);
nand U4794 (N_4794,N_3294,N_3615);
nor U4795 (N_4795,N_3435,N_3234);
nor U4796 (N_4796,N_3618,N_3549);
nor U4797 (N_4797,N_3108,N_3882);
and U4798 (N_4798,N_3671,N_3687);
nand U4799 (N_4799,N_3929,N_3734);
or U4800 (N_4800,N_3900,N_3829);
and U4801 (N_4801,N_3179,N_3615);
nor U4802 (N_4802,N_3091,N_3586);
nor U4803 (N_4803,N_3382,N_3912);
nand U4804 (N_4804,N_3796,N_3320);
nand U4805 (N_4805,N_3128,N_3785);
nand U4806 (N_4806,N_3072,N_3163);
nor U4807 (N_4807,N_3997,N_3666);
nor U4808 (N_4808,N_3975,N_3487);
nor U4809 (N_4809,N_3954,N_3768);
and U4810 (N_4810,N_3468,N_3872);
nor U4811 (N_4811,N_3989,N_3792);
and U4812 (N_4812,N_3664,N_3293);
or U4813 (N_4813,N_3955,N_3205);
or U4814 (N_4814,N_3960,N_3591);
or U4815 (N_4815,N_3517,N_3533);
or U4816 (N_4816,N_3610,N_3336);
nand U4817 (N_4817,N_3833,N_3050);
or U4818 (N_4818,N_3322,N_3249);
nand U4819 (N_4819,N_3628,N_3204);
or U4820 (N_4820,N_3077,N_3349);
nand U4821 (N_4821,N_3008,N_3640);
nand U4822 (N_4822,N_3254,N_3324);
or U4823 (N_4823,N_3159,N_3975);
nor U4824 (N_4824,N_3118,N_3669);
nor U4825 (N_4825,N_3615,N_3184);
and U4826 (N_4826,N_3832,N_3336);
or U4827 (N_4827,N_3181,N_3244);
nand U4828 (N_4828,N_3431,N_3330);
nor U4829 (N_4829,N_3930,N_3041);
and U4830 (N_4830,N_3504,N_3316);
and U4831 (N_4831,N_3846,N_3244);
nand U4832 (N_4832,N_3280,N_3514);
nand U4833 (N_4833,N_3962,N_3268);
nor U4834 (N_4834,N_3341,N_3524);
or U4835 (N_4835,N_3291,N_3629);
nor U4836 (N_4836,N_3984,N_3998);
nand U4837 (N_4837,N_3833,N_3319);
nor U4838 (N_4838,N_3585,N_3526);
or U4839 (N_4839,N_3745,N_3983);
and U4840 (N_4840,N_3958,N_3345);
or U4841 (N_4841,N_3205,N_3607);
and U4842 (N_4842,N_3873,N_3007);
or U4843 (N_4843,N_3723,N_3543);
nand U4844 (N_4844,N_3151,N_3178);
nand U4845 (N_4845,N_3453,N_3079);
nor U4846 (N_4846,N_3887,N_3253);
nand U4847 (N_4847,N_3505,N_3781);
nor U4848 (N_4848,N_3128,N_3358);
nor U4849 (N_4849,N_3917,N_3719);
nand U4850 (N_4850,N_3528,N_3842);
nand U4851 (N_4851,N_3560,N_3647);
nand U4852 (N_4852,N_3516,N_3446);
xor U4853 (N_4853,N_3127,N_3149);
and U4854 (N_4854,N_3511,N_3956);
nand U4855 (N_4855,N_3984,N_3589);
and U4856 (N_4856,N_3171,N_3661);
or U4857 (N_4857,N_3448,N_3173);
nand U4858 (N_4858,N_3619,N_3675);
and U4859 (N_4859,N_3921,N_3960);
and U4860 (N_4860,N_3672,N_3393);
nor U4861 (N_4861,N_3495,N_3165);
and U4862 (N_4862,N_3251,N_3083);
and U4863 (N_4863,N_3163,N_3473);
or U4864 (N_4864,N_3539,N_3551);
or U4865 (N_4865,N_3140,N_3437);
nand U4866 (N_4866,N_3985,N_3389);
or U4867 (N_4867,N_3490,N_3840);
nor U4868 (N_4868,N_3560,N_3737);
or U4869 (N_4869,N_3261,N_3891);
and U4870 (N_4870,N_3376,N_3766);
nand U4871 (N_4871,N_3363,N_3811);
or U4872 (N_4872,N_3403,N_3449);
or U4873 (N_4873,N_3582,N_3009);
nor U4874 (N_4874,N_3871,N_3981);
nand U4875 (N_4875,N_3402,N_3809);
and U4876 (N_4876,N_3566,N_3618);
nor U4877 (N_4877,N_3557,N_3643);
nand U4878 (N_4878,N_3922,N_3045);
or U4879 (N_4879,N_3246,N_3329);
nand U4880 (N_4880,N_3128,N_3592);
and U4881 (N_4881,N_3573,N_3030);
and U4882 (N_4882,N_3807,N_3519);
or U4883 (N_4883,N_3748,N_3744);
nor U4884 (N_4884,N_3043,N_3643);
nor U4885 (N_4885,N_3208,N_3280);
or U4886 (N_4886,N_3531,N_3650);
nor U4887 (N_4887,N_3858,N_3708);
or U4888 (N_4888,N_3119,N_3352);
nor U4889 (N_4889,N_3335,N_3859);
nor U4890 (N_4890,N_3942,N_3968);
or U4891 (N_4891,N_3037,N_3191);
or U4892 (N_4892,N_3779,N_3776);
and U4893 (N_4893,N_3283,N_3118);
or U4894 (N_4894,N_3860,N_3380);
xnor U4895 (N_4895,N_3548,N_3943);
or U4896 (N_4896,N_3567,N_3690);
or U4897 (N_4897,N_3314,N_3818);
nor U4898 (N_4898,N_3932,N_3682);
and U4899 (N_4899,N_3210,N_3828);
nand U4900 (N_4900,N_3114,N_3040);
nor U4901 (N_4901,N_3768,N_3020);
nor U4902 (N_4902,N_3209,N_3613);
or U4903 (N_4903,N_3864,N_3194);
and U4904 (N_4904,N_3654,N_3269);
nor U4905 (N_4905,N_3166,N_3787);
nand U4906 (N_4906,N_3802,N_3510);
and U4907 (N_4907,N_3936,N_3090);
and U4908 (N_4908,N_3126,N_3298);
nor U4909 (N_4909,N_3517,N_3660);
and U4910 (N_4910,N_3397,N_3790);
and U4911 (N_4911,N_3848,N_3414);
and U4912 (N_4912,N_3108,N_3794);
and U4913 (N_4913,N_3890,N_3074);
nor U4914 (N_4914,N_3565,N_3872);
and U4915 (N_4915,N_3279,N_3094);
nand U4916 (N_4916,N_3871,N_3822);
or U4917 (N_4917,N_3203,N_3312);
nand U4918 (N_4918,N_3666,N_3319);
nand U4919 (N_4919,N_3173,N_3367);
or U4920 (N_4920,N_3113,N_3578);
and U4921 (N_4921,N_3226,N_3779);
or U4922 (N_4922,N_3837,N_3948);
nor U4923 (N_4923,N_3042,N_3470);
and U4924 (N_4924,N_3610,N_3393);
and U4925 (N_4925,N_3439,N_3264);
nand U4926 (N_4926,N_3135,N_3436);
nor U4927 (N_4927,N_3023,N_3479);
and U4928 (N_4928,N_3425,N_3078);
nor U4929 (N_4929,N_3235,N_3890);
nand U4930 (N_4930,N_3459,N_3296);
or U4931 (N_4931,N_3298,N_3627);
or U4932 (N_4932,N_3054,N_3792);
and U4933 (N_4933,N_3440,N_3563);
nor U4934 (N_4934,N_3576,N_3673);
nor U4935 (N_4935,N_3536,N_3631);
and U4936 (N_4936,N_3772,N_3353);
xor U4937 (N_4937,N_3709,N_3009);
and U4938 (N_4938,N_3699,N_3254);
nand U4939 (N_4939,N_3329,N_3536);
or U4940 (N_4940,N_3446,N_3517);
or U4941 (N_4941,N_3662,N_3357);
and U4942 (N_4942,N_3215,N_3916);
nor U4943 (N_4943,N_3681,N_3911);
nor U4944 (N_4944,N_3656,N_3914);
and U4945 (N_4945,N_3718,N_3805);
nor U4946 (N_4946,N_3831,N_3890);
xnor U4947 (N_4947,N_3831,N_3763);
nor U4948 (N_4948,N_3042,N_3423);
and U4949 (N_4949,N_3001,N_3032);
nor U4950 (N_4950,N_3223,N_3264);
and U4951 (N_4951,N_3771,N_3441);
nand U4952 (N_4952,N_3703,N_3345);
and U4953 (N_4953,N_3775,N_3136);
nor U4954 (N_4954,N_3086,N_3810);
nor U4955 (N_4955,N_3010,N_3043);
and U4956 (N_4956,N_3665,N_3190);
or U4957 (N_4957,N_3772,N_3118);
nand U4958 (N_4958,N_3755,N_3604);
or U4959 (N_4959,N_3403,N_3290);
nor U4960 (N_4960,N_3155,N_3192);
or U4961 (N_4961,N_3501,N_3380);
nand U4962 (N_4962,N_3251,N_3608);
and U4963 (N_4963,N_3486,N_3326);
or U4964 (N_4964,N_3184,N_3950);
and U4965 (N_4965,N_3129,N_3593);
nor U4966 (N_4966,N_3749,N_3245);
or U4967 (N_4967,N_3090,N_3985);
nand U4968 (N_4968,N_3745,N_3781);
nor U4969 (N_4969,N_3967,N_3999);
or U4970 (N_4970,N_3582,N_3553);
and U4971 (N_4971,N_3093,N_3642);
nand U4972 (N_4972,N_3391,N_3694);
nand U4973 (N_4973,N_3509,N_3516);
nand U4974 (N_4974,N_3162,N_3044);
and U4975 (N_4975,N_3369,N_3912);
or U4976 (N_4976,N_3908,N_3258);
and U4977 (N_4977,N_3706,N_3802);
nand U4978 (N_4978,N_3927,N_3082);
and U4979 (N_4979,N_3464,N_3244);
and U4980 (N_4980,N_3607,N_3196);
nor U4981 (N_4981,N_3354,N_3528);
nor U4982 (N_4982,N_3702,N_3008);
nor U4983 (N_4983,N_3716,N_3545);
nor U4984 (N_4984,N_3797,N_3728);
nor U4985 (N_4985,N_3267,N_3375);
nand U4986 (N_4986,N_3420,N_3796);
and U4987 (N_4987,N_3762,N_3528);
nand U4988 (N_4988,N_3941,N_3640);
nor U4989 (N_4989,N_3422,N_3502);
nor U4990 (N_4990,N_3410,N_3380);
and U4991 (N_4991,N_3877,N_3211);
nand U4992 (N_4992,N_3263,N_3192);
nor U4993 (N_4993,N_3177,N_3513);
nand U4994 (N_4994,N_3531,N_3724);
and U4995 (N_4995,N_3125,N_3908);
and U4996 (N_4996,N_3810,N_3809);
nand U4997 (N_4997,N_3904,N_3775);
nand U4998 (N_4998,N_3359,N_3287);
or U4999 (N_4999,N_3285,N_3229);
or U5000 (N_5000,N_4455,N_4418);
nand U5001 (N_5001,N_4001,N_4436);
nor U5002 (N_5002,N_4952,N_4621);
and U5003 (N_5003,N_4800,N_4341);
or U5004 (N_5004,N_4324,N_4350);
or U5005 (N_5005,N_4853,N_4470);
nor U5006 (N_5006,N_4877,N_4162);
or U5007 (N_5007,N_4799,N_4101);
nand U5008 (N_5008,N_4511,N_4863);
nor U5009 (N_5009,N_4122,N_4238);
nor U5010 (N_5010,N_4038,N_4339);
nor U5011 (N_5011,N_4267,N_4434);
nand U5012 (N_5012,N_4012,N_4165);
nand U5013 (N_5013,N_4944,N_4253);
nand U5014 (N_5014,N_4115,N_4018);
or U5015 (N_5015,N_4219,N_4599);
or U5016 (N_5016,N_4456,N_4929);
nor U5017 (N_5017,N_4426,N_4995);
or U5018 (N_5018,N_4871,N_4246);
nand U5019 (N_5019,N_4521,N_4232);
nand U5020 (N_5020,N_4340,N_4626);
or U5021 (N_5021,N_4728,N_4619);
nor U5022 (N_5022,N_4093,N_4309);
or U5023 (N_5023,N_4475,N_4243);
xor U5024 (N_5024,N_4723,N_4110);
nand U5025 (N_5025,N_4379,N_4605);
or U5026 (N_5026,N_4941,N_4123);
and U5027 (N_5027,N_4380,N_4789);
nand U5028 (N_5028,N_4450,N_4580);
or U5029 (N_5029,N_4722,N_4003);
or U5030 (N_5030,N_4473,N_4355);
nor U5031 (N_5031,N_4199,N_4260);
nor U5032 (N_5032,N_4490,N_4888);
or U5033 (N_5033,N_4480,N_4215);
nor U5034 (N_5034,N_4827,N_4264);
nor U5035 (N_5035,N_4988,N_4277);
nor U5036 (N_5036,N_4601,N_4532);
nor U5037 (N_5037,N_4642,N_4903);
nand U5038 (N_5038,N_4058,N_4420);
or U5039 (N_5039,N_4501,N_4977);
and U5040 (N_5040,N_4907,N_4411);
nor U5041 (N_5041,N_4374,N_4329);
and U5042 (N_5042,N_4416,N_4275);
nand U5043 (N_5043,N_4064,N_4106);
and U5044 (N_5044,N_4760,N_4709);
nand U5045 (N_5045,N_4421,N_4000);
or U5046 (N_5046,N_4075,N_4125);
or U5047 (N_5047,N_4936,N_4160);
and U5048 (N_5048,N_4478,N_4690);
or U5049 (N_5049,N_4507,N_4498);
nor U5050 (N_5050,N_4677,N_4306);
and U5051 (N_5051,N_4033,N_4778);
nand U5052 (N_5052,N_4195,N_4831);
or U5053 (N_5053,N_4155,N_4039);
and U5054 (N_5054,N_4856,N_4183);
nor U5055 (N_5055,N_4116,N_4625);
nand U5056 (N_5056,N_4196,N_4210);
nor U5057 (N_5057,N_4323,N_4504);
and U5058 (N_5058,N_4011,N_4112);
nor U5059 (N_5059,N_4527,N_4131);
or U5060 (N_5060,N_4793,N_4274);
nand U5061 (N_5061,N_4537,N_4235);
or U5062 (N_5062,N_4497,N_4540);
and U5063 (N_5063,N_4556,N_4717);
or U5064 (N_5064,N_4515,N_4213);
or U5065 (N_5065,N_4797,N_4710);
nand U5066 (N_5066,N_4822,N_4136);
nand U5067 (N_5067,N_4749,N_4188);
nor U5068 (N_5068,N_4686,N_4041);
and U5069 (N_5069,N_4975,N_4399);
and U5070 (N_5070,N_4454,N_4865);
nand U5071 (N_5071,N_4387,N_4792);
and U5072 (N_5072,N_4807,N_4342);
nor U5073 (N_5073,N_4163,N_4998);
nor U5074 (N_5074,N_4653,N_4970);
xnor U5075 (N_5075,N_4627,N_4826);
nor U5076 (N_5076,N_4356,N_4948);
or U5077 (N_5077,N_4588,N_4146);
nand U5078 (N_5078,N_4631,N_4730);
or U5079 (N_5079,N_4885,N_4102);
nor U5080 (N_5080,N_4539,N_4816);
and U5081 (N_5081,N_4180,N_4549);
or U5082 (N_5082,N_4397,N_4230);
or U5083 (N_5083,N_4485,N_4844);
or U5084 (N_5084,N_4933,N_4185);
or U5085 (N_5085,N_4014,N_4758);
and U5086 (N_5086,N_4996,N_4472);
nand U5087 (N_5087,N_4629,N_4296);
nor U5088 (N_5088,N_4139,N_4770);
and U5089 (N_5089,N_4972,N_4207);
nand U5090 (N_5090,N_4942,N_4283);
and U5091 (N_5091,N_4285,N_4810);
or U5092 (N_5092,N_4422,N_4652);
nor U5093 (N_5093,N_4451,N_4688);
or U5094 (N_5094,N_4834,N_4239);
nor U5095 (N_5095,N_4665,N_4325);
nor U5096 (N_5096,N_4392,N_4755);
nor U5097 (N_5097,N_4425,N_4693);
nor U5098 (N_5098,N_4320,N_4555);
or U5099 (N_5099,N_4365,N_4233);
and U5100 (N_5100,N_4358,N_4674);
and U5101 (N_5101,N_4271,N_4567);
or U5102 (N_5102,N_4600,N_4869);
or U5103 (N_5103,N_4939,N_4591);
nor U5104 (N_5104,N_4985,N_4724);
and U5105 (N_5105,N_4109,N_4026);
nor U5106 (N_5106,N_4638,N_4250);
nor U5107 (N_5107,N_4214,N_4337);
or U5108 (N_5108,N_4432,N_4280);
nor U5109 (N_5109,N_4510,N_4276);
nor U5110 (N_5110,N_4444,N_4587);
nor U5111 (N_5111,N_4494,N_4171);
nor U5112 (N_5112,N_4303,N_4801);
nand U5113 (N_5113,N_4153,N_4804);
nor U5114 (N_5114,N_4345,N_4767);
nor U5115 (N_5115,N_4299,N_4791);
nand U5116 (N_5116,N_4366,N_4209);
or U5117 (N_5117,N_4842,N_4570);
nor U5118 (N_5118,N_4773,N_4828);
and U5119 (N_5119,N_4746,N_4229);
and U5120 (N_5120,N_4083,N_4937);
nand U5121 (N_5121,N_4095,N_4569);
or U5122 (N_5122,N_4646,N_4928);
or U5123 (N_5123,N_4911,N_4389);
and U5124 (N_5124,N_4062,N_4634);
nand U5125 (N_5125,N_4533,N_4304);
nand U5126 (N_5126,N_4817,N_4986);
nor U5127 (N_5127,N_4245,N_4419);
nand U5128 (N_5128,N_4874,N_4013);
and U5129 (N_5129,N_4137,N_4071);
nand U5130 (N_5130,N_4658,N_4811);
nor U5131 (N_5131,N_4481,N_4117);
and U5132 (N_5132,N_4585,N_4441);
nor U5133 (N_5133,N_4097,N_4343);
nand U5134 (N_5134,N_4133,N_4896);
xnor U5135 (N_5135,N_4595,N_4734);
and U5136 (N_5136,N_4108,N_4035);
and U5137 (N_5137,N_4057,N_4573);
and U5138 (N_5138,N_4346,N_4484);
or U5139 (N_5139,N_4782,N_4173);
nor U5140 (N_5140,N_4904,N_4543);
nor U5141 (N_5141,N_4876,N_4545);
and U5142 (N_5142,N_4920,N_4187);
nand U5143 (N_5143,N_4649,N_4669);
and U5144 (N_5144,N_4186,N_4524);
and U5145 (N_5145,N_4316,N_4505);
nor U5146 (N_5146,N_4868,N_4336);
nor U5147 (N_5147,N_4417,N_4733);
or U5148 (N_5148,N_4025,N_4708);
and U5149 (N_5149,N_4630,N_4667);
or U5150 (N_5150,N_4881,N_4007);
or U5151 (N_5151,N_4697,N_4867);
and U5152 (N_5152,N_4034,N_4766);
or U5153 (N_5153,N_4568,N_4247);
nand U5154 (N_5154,N_4616,N_4575);
nor U5155 (N_5155,N_4613,N_4221);
and U5156 (N_5156,N_4564,N_4546);
and U5157 (N_5157,N_4732,N_4381);
or U5158 (N_5158,N_4086,N_4819);
nor U5159 (N_5159,N_4692,N_4976);
or U5160 (N_5160,N_4287,N_4583);
nor U5161 (N_5161,N_4503,N_4774);
and U5162 (N_5162,N_4973,N_4256);
nand U5163 (N_5163,N_4447,N_4360);
and U5164 (N_5164,N_4302,N_4242);
nor U5165 (N_5165,N_4938,N_4969);
nor U5166 (N_5166,N_4307,N_4037);
nor U5167 (N_5167,N_4500,N_4783);
or U5168 (N_5168,N_4496,N_4886);
or U5169 (N_5169,N_4184,N_4678);
nor U5170 (N_5170,N_4716,N_4368);
and U5171 (N_5171,N_4319,N_4582);
and U5172 (N_5172,N_4428,N_4781);
nor U5173 (N_5173,N_4081,N_4676);
or U5174 (N_5174,N_4482,N_4747);
and U5175 (N_5175,N_4956,N_4148);
nand U5176 (N_5176,N_4502,N_4872);
nand U5177 (N_5177,N_4963,N_4802);
and U5178 (N_5178,N_4633,N_4855);
or U5179 (N_5179,N_4427,N_4182);
nand U5180 (N_5180,N_4407,N_4359);
nor U5181 (N_5181,N_4618,N_4166);
nand U5182 (N_5182,N_4405,N_4236);
and U5183 (N_5183,N_4918,N_4517);
nand U5184 (N_5184,N_4351,N_4400);
nand U5185 (N_5185,N_4413,N_4852);
nand U5186 (N_5186,N_4523,N_4449);
nor U5187 (N_5187,N_4906,N_4396);
or U5188 (N_5188,N_4795,N_4541);
and U5189 (N_5189,N_4661,N_4949);
nand U5190 (N_5190,N_4921,N_4679);
and U5191 (N_5191,N_4964,N_4909);
or U5192 (N_5192,N_4477,N_4061);
nand U5193 (N_5193,N_4735,N_4032);
nand U5194 (N_5194,N_4823,N_4887);
nor U5195 (N_5195,N_4771,N_4009);
or U5196 (N_5196,N_4288,N_4689);
and U5197 (N_5197,N_4495,N_4435);
and U5198 (N_5198,N_4980,N_4189);
nand U5199 (N_5199,N_4635,N_4445);
or U5200 (N_5200,N_4409,N_4005);
and U5201 (N_5201,N_4286,N_4803);
or U5202 (N_5202,N_4753,N_4310);
nand U5203 (N_5203,N_4790,N_4111);
or U5204 (N_5204,N_4281,N_4848);
nand U5205 (N_5205,N_4947,N_4684);
and U5206 (N_5206,N_4741,N_4703);
or U5207 (N_5207,N_4094,N_4002);
or U5208 (N_5208,N_4377,N_4893);
and U5209 (N_5209,N_4592,N_4135);
nor U5210 (N_5210,N_4363,N_4727);
and U5211 (N_5211,N_4934,N_4483);
or U5212 (N_5212,N_4464,N_4751);
nand U5213 (N_5213,N_4401,N_4654);
nand U5214 (N_5214,N_4089,N_4114);
or U5215 (N_5215,N_4547,N_4718);
nand U5216 (N_5216,N_4344,N_4408);
nand U5217 (N_5217,N_4327,N_4971);
nor U5218 (N_5218,N_4042,N_4784);
and U5219 (N_5219,N_4141,N_4491);
nor U5220 (N_5220,N_4895,N_4206);
nor U5221 (N_5221,N_4590,N_4237);
nand U5222 (N_5222,N_4958,N_4151);
nand U5223 (N_5223,N_4251,N_4768);
nand U5224 (N_5224,N_4489,N_4147);
or U5225 (N_5225,N_4048,N_4130);
nand U5226 (N_5226,N_4530,N_4090);
or U5227 (N_5227,N_4092,N_4552);
nand U5228 (N_5228,N_4073,N_4036);
nor U5229 (N_5229,N_4809,N_4258);
nand U5230 (N_5230,N_4702,N_4301);
or U5231 (N_5231,N_4371,N_4082);
nand U5232 (N_5232,N_4712,N_4586);
and U5233 (N_5233,N_4177,N_4047);
or U5234 (N_5234,N_4891,N_4596);
nor U5235 (N_5235,N_4597,N_4651);
nor U5236 (N_5236,N_4950,N_4312);
and U5237 (N_5237,N_4443,N_4467);
nand U5238 (N_5238,N_4538,N_4143);
nor U5239 (N_5239,N_4640,N_4923);
nor U5240 (N_5240,N_4067,N_4338);
nand U5241 (N_5241,N_4284,N_4334);
nand U5242 (N_5242,N_4813,N_4333);
or U5243 (N_5243,N_4721,N_4265);
nand U5244 (N_5244,N_4927,N_4015);
nor U5245 (N_5245,N_4750,N_4328);
nor U5246 (N_5246,N_4765,N_4020);
nand U5247 (N_5247,N_4528,N_4412);
nor U5248 (N_5248,N_4068,N_4987);
and U5249 (N_5249,N_4706,N_4926);
and U5250 (N_5250,N_4119,N_4022);
nor U5251 (N_5251,N_4922,N_4332);
nor U5252 (N_5252,N_4992,N_4897);
and U5253 (N_5253,N_4305,N_4694);
nand U5254 (N_5254,N_4311,N_4562);
nand U5255 (N_5255,N_4049,N_4925);
or U5256 (N_5256,N_4474,N_4979);
nand U5257 (N_5257,N_4096,N_4079);
nor U5258 (N_5258,N_4668,N_4691);
nor U5259 (N_5259,N_4168,N_4846);
nor U5260 (N_5260,N_4225,N_4492);
or U5261 (N_5261,N_4269,N_4849);
nor U5262 (N_5262,N_4603,N_4589);
and U5263 (N_5263,N_4118,N_4879);
and U5264 (N_5264,N_4606,N_4211);
and U5265 (N_5265,N_4255,N_4430);
nor U5266 (N_5266,N_4318,N_4632);
nor U5267 (N_5267,N_4650,N_4152);
or U5268 (N_5268,N_4272,N_4901);
nand U5269 (N_5269,N_4157,N_4617);
nor U5270 (N_5270,N_4989,N_4442);
and U5271 (N_5271,N_4685,N_4628);
nand U5272 (N_5272,N_4699,N_4369);
nor U5273 (N_5273,N_4981,N_4839);
nand U5274 (N_5274,N_4719,N_4832);
and U5275 (N_5275,N_4382,N_4860);
nor U5276 (N_5276,N_4913,N_4637);
and U5277 (N_5277,N_4990,N_4814);
or U5278 (N_5278,N_4295,N_4683);
and U5279 (N_5279,N_4493,N_4469);
nand U5280 (N_5280,N_4720,N_4598);
or U5281 (N_5281,N_4191,N_4244);
or U5282 (N_5282,N_4076,N_4576);
or U5283 (N_5283,N_4818,N_4088);
nand U5284 (N_5284,N_4931,N_4608);
or U5285 (N_5285,N_4257,N_4330);
or U5286 (N_5286,N_4508,N_4912);
or U5287 (N_5287,N_4223,N_4704);
and U5288 (N_5288,N_4357,N_4806);
nand U5289 (N_5289,N_4935,N_4390);
and U5290 (N_5290,N_4660,N_4349);
and U5291 (N_5291,N_4103,N_4200);
or U5292 (N_5292,N_4824,N_4615);
and U5293 (N_5293,N_4252,N_4056);
and U5294 (N_5294,N_4203,N_4205);
nand U5295 (N_5295,N_4880,N_4461);
or U5296 (N_5296,N_4065,N_4763);
nor U5297 (N_5297,N_4574,N_4870);
and U5298 (N_5298,N_4959,N_4087);
and U5299 (N_5299,N_4140,N_4446);
nand U5300 (N_5300,N_4940,N_4584);
nor U5301 (N_5301,N_4393,N_4282);
nand U5302 (N_5302,N_4883,N_4466);
or U5303 (N_5303,N_4840,N_4966);
and U5304 (N_5304,N_4170,N_4965);
or U5305 (N_5305,N_4178,N_4748);
or U5306 (N_5306,N_4620,N_4074);
nand U5307 (N_5307,N_4080,N_4815);
or U5308 (N_5308,N_4978,N_4391);
and U5309 (N_5309,N_4594,N_4394);
and U5310 (N_5310,N_4051,N_4268);
nor U5311 (N_5311,N_4006,N_4534);
nor U5312 (N_5312,N_4156,N_4991);
and U5313 (N_5313,N_4217,N_4623);
nor U5314 (N_5314,N_4462,N_4725);
nor U5315 (N_5315,N_4529,N_4259);
or U5316 (N_5316,N_4270,N_4577);
and U5317 (N_5317,N_4664,N_4046);
nor U5318 (N_5318,N_4463,N_4054);
and U5319 (N_5319,N_4579,N_4019);
nor U5320 (N_5320,N_4297,N_4604);
nor U5321 (N_5321,N_4614,N_4031);
nand U5322 (N_5322,N_4878,N_4231);
or U5323 (N_5323,N_4127,N_4898);
and U5324 (N_5324,N_4439,N_4460);
nand U5325 (N_5325,N_4314,N_4645);
nor U5326 (N_5326,N_4657,N_4364);
or U5327 (N_5327,N_4943,N_4794);
nand U5328 (N_5328,N_4077,N_4370);
and U5329 (N_5329,N_4100,N_4851);
nor U5330 (N_5330,N_4861,N_4729);
and U5331 (N_5331,N_4375,N_4465);
nand U5332 (N_5332,N_4085,N_4107);
or U5333 (N_5333,N_4662,N_4731);
nor U5334 (N_5334,N_4053,N_4999);
nand U5335 (N_5335,N_4776,N_4593);
nand U5336 (N_5336,N_4957,N_4278);
or U5337 (N_5337,N_4315,N_4362);
or U5338 (N_5338,N_4698,N_4908);
and U5339 (N_5339,N_4565,N_4754);
nand U5340 (N_5340,N_4044,N_4542);
nor U5341 (N_5341,N_4761,N_4841);
nand U5342 (N_5342,N_4994,N_4403);
nand U5343 (N_5343,N_4671,N_4429);
and U5344 (N_5344,N_4675,N_4670);
or U5345 (N_5345,N_4805,N_4739);
nand U5346 (N_5346,N_4930,N_4571);
nor U5347 (N_5347,N_4352,N_4993);
or U5348 (N_5348,N_4641,N_4138);
or U5349 (N_5349,N_4967,N_4202);
and U5350 (N_5350,N_4572,N_4738);
nor U5351 (N_5351,N_4820,N_4149);
and U5352 (N_5352,N_4701,N_4643);
nand U5353 (N_5353,N_4150,N_4300);
and U5354 (N_5354,N_4663,N_4932);
or U5355 (N_5355,N_4845,N_4946);
and U5356 (N_5356,N_4129,N_4535);
nand U5357 (N_5357,N_4759,N_4864);
nand U5358 (N_5358,N_4513,N_4821);
nor U5359 (N_5359,N_4084,N_4241);
and U5360 (N_5360,N_4953,N_4028);
and U5361 (N_5361,N_4326,N_4126);
nor U5362 (N_5362,N_4559,N_4762);
or U5363 (N_5363,N_4273,N_4175);
nand U5364 (N_5364,N_4681,N_4737);
or U5365 (N_5365,N_4955,N_4059);
nor U5366 (N_5366,N_4779,N_4752);
nand U5367 (N_5367,N_4383,N_4960);
nor U5368 (N_5368,N_4910,N_4438);
nor U5369 (N_5369,N_4248,N_4027);
and U5370 (N_5370,N_4968,N_4558);
nor U5371 (N_5371,N_4289,N_4070);
or U5372 (N_5372,N_4843,N_4566);
nand U5373 (N_5373,N_4164,N_4226);
and U5374 (N_5374,N_4764,N_4487);
and U5375 (N_5375,N_4373,N_4388);
and U5376 (N_5376,N_4372,N_4673);
or U5377 (N_5377,N_4548,N_4395);
nand U5378 (N_5378,N_4700,N_4866);
nand U5379 (N_5379,N_4402,N_4424);
and U5380 (N_5380,N_4894,N_4982);
and U5381 (N_5381,N_4197,N_4040);
or U5382 (N_5382,N_4847,N_4004);
or U5383 (N_5383,N_4829,N_4120);
nand U5384 (N_5384,N_4655,N_4458);
nor U5385 (N_5385,N_4105,N_4249);
nand U5386 (N_5386,N_4132,N_4208);
and U5387 (N_5387,N_4376,N_4914);
nand U5388 (N_5388,N_4190,N_4335);
nand U5389 (N_5389,N_4581,N_4744);
nor U5390 (N_5390,N_4578,N_4290);
and U5391 (N_5391,N_4899,N_4945);
and U5392 (N_5392,N_4398,N_4974);
and U5393 (N_5393,N_4361,N_4008);
nor U5394 (N_5394,N_4404,N_4179);
or U5395 (N_5395,N_4726,N_4854);
nand U5396 (N_5396,N_4780,N_4917);
nor U5397 (N_5397,N_4551,N_4261);
and U5398 (N_5398,N_4788,N_4951);
and U5399 (N_5399,N_4757,N_4743);
and U5400 (N_5400,N_4715,N_4769);
nand U5401 (N_5401,N_4410,N_4181);
nand U5402 (N_5402,N_4499,N_4526);
nand U5403 (N_5403,N_4666,N_4218);
and U5404 (N_5404,N_4516,N_4159);
nor U5405 (N_5405,N_4525,N_4837);
and U5406 (N_5406,N_4322,N_4063);
and U5407 (N_5407,N_4984,N_4128);
nand U5408 (N_5408,N_4777,N_4563);
nor U5409 (N_5409,N_4055,N_4321);
or U5410 (N_5410,N_4317,N_4385);
nor U5411 (N_5411,N_4468,N_4682);
nor U5412 (N_5412,N_4506,N_4142);
or U5413 (N_5413,N_4154,N_4518);
nor U5414 (N_5414,N_4017,N_4557);
nor U5415 (N_5415,N_4212,N_4648);
nor U5416 (N_5416,N_4622,N_4415);
nor U5417 (N_5417,N_4113,N_4656);
and U5418 (N_5418,N_4194,N_4636);
nand U5419 (N_5419,N_4787,N_4602);
nor U5420 (N_5420,N_4890,N_4161);
nand U5421 (N_5421,N_4023,N_4220);
nand U5422 (N_5422,N_4386,N_4121);
or U5423 (N_5423,N_4030,N_4266);
nor U5424 (N_5424,N_4512,N_4354);
nand U5425 (N_5425,N_4240,N_4672);
and U5426 (N_5426,N_4553,N_4263);
or U5427 (N_5427,N_4192,N_4850);
and U5428 (N_5428,N_4687,N_4291);
nor U5429 (N_5429,N_4124,N_4786);
nor U5430 (N_5430,N_4262,N_4457);
and U5431 (N_5431,N_4775,N_4833);
nor U5432 (N_5432,N_4459,N_4104);
nor U5433 (N_5433,N_4772,N_4607);
nor U5434 (N_5434,N_4448,N_4902);
or U5435 (N_5435,N_4954,N_4875);
or U5436 (N_5436,N_4962,N_4367);
nor U5437 (N_5437,N_4134,N_4544);
or U5438 (N_5438,N_4384,N_4091);
and U5439 (N_5439,N_4167,N_4045);
nor U5440 (N_5440,N_4889,N_4293);
nand U5441 (N_5441,N_4452,N_4644);
nor U5442 (N_5442,N_4216,N_4016);
nor U5443 (N_5443,N_4740,N_4915);
nand U5444 (N_5444,N_4331,N_4695);
or U5445 (N_5445,N_4078,N_4234);
or U5446 (N_5446,N_4158,N_4659);
and U5447 (N_5447,N_4924,N_4835);
nand U5448 (N_5448,N_4997,N_4098);
nor U5449 (N_5449,N_4476,N_4414);
nand U5450 (N_5450,N_4560,N_4072);
nor U5451 (N_5451,N_4292,N_4254);
and U5452 (N_5452,N_4193,N_4224);
nand U5453 (N_5453,N_4825,N_4812);
and U5454 (N_5454,N_4021,N_4440);
and U5455 (N_5455,N_4858,N_4900);
or U5456 (N_5456,N_4531,N_4857);
nor U5457 (N_5457,N_4169,N_4882);
nor U5458 (N_5458,N_4204,N_4279);
and U5459 (N_5459,N_4961,N_4522);
and U5460 (N_5460,N_4479,N_4010);
nor U5461 (N_5461,N_4808,N_4519);
nor U5462 (N_5462,N_4714,N_4043);
nor U5463 (N_5463,N_4099,N_4836);
or U5464 (N_5464,N_4680,N_4144);
nor U5465 (N_5465,N_4308,N_4611);
nor U5466 (N_5466,N_4647,N_4222);
nor U5467 (N_5467,N_4610,N_4198);
nand U5468 (N_5468,N_4536,N_4069);
and U5469 (N_5469,N_4639,N_4029);
nand U5470 (N_5470,N_4423,N_4453);
or U5471 (N_5471,N_4520,N_4798);
nor U5472 (N_5472,N_4707,N_4294);
nand U5473 (N_5473,N_4052,N_4554);
nor U5474 (N_5474,N_4347,N_4983);
and U5475 (N_5475,N_4919,N_4431);
nand U5476 (N_5476,N_4313,N_4488);
and U5477 (N_5477,N_4378,N_4609);
nor U5478 (N_5478,N_4705,N_4873);
and U5479 (N_5479,N_4050,N_4916);
and U5480 (N_5480,N_4745,N_4838);
nand U5481 (N_5481,N_4227,N_4859);
nand U5482 (N_5482,N_4612,N_4201);
or U5483 (N_5483,N_4437,N_4624);
nand U5484 (N_5484,N_4796,N_4884);
and U5485 (N_5485,N_4348,N_4486);
nand U5486 (N_5486,N_4696,N_4145);
and U5487 (N_5487,N_4550,N_4433);
or U5488 (N_5488,N_4060,N_4711);
nand U5489 (N_5489,N_4785,N_4892);
or U5490 (N_5490,N_4228,N_4176);
nand U5491 (N_5491,N_4172,N_4514);
and U5492 (N_5492,N_4471,N_4756);
or U5493 (N_5493,N_4174,N_4353);
nand U5494 (N_5494,N_4561,N_4862);
nand U5495 (N_5495,N_4742,N_4736);
nand U5496 (N_5496,N_4509,N_4024);
nand U5497 (N_5497,N_4406,N_4905);
nand U5498 (N_5498,N_4830,N_4713);
or U5499 (N_5499,N_4066,N_4298);
and U5500 (N_5500,N_4455,N_4780);
nand U5501 (N_5501,N_4272,N_4848);
and U5502 (N_5502,N_4817,N_4266);
nor U5503 (N_5503,N_4678,N_4091);
and U5504 (N_5504,N_4097,N_4259);
and U5505 (N_5505,N_4207,N_4257);
nand U5506 (N_5506,N_4709,N_4497);
and U5507 (N_5507,N_4855,N_4903);
and U5508 (N_5508,N_4700,N_4565);
or U5509 (N_5509,N_4168,N_4767);
nor U5510 (N_5510,N_4709,N_4955);
nand U5511 (N_5511,N_4158,N_4880);
and U5512 (N_5512,N_4996,N_4937);
nand U5513 (N_5513,N_4568,N_4242);
nor U5514 (N_5514,N_4094,N_4524);
and U5515 (N_5515,N_4717,N_4140);
and U5516 (N_5516,N_4846,N_4435);
nor U5517 (N_5517,N_4723,N_4885);
or U5518 (N_5518,N_4741,N_4392);
nor U5519 (N_5519,N_4311,N_4305);
nand U5520 (N_5520,N_4082,N_4578);
nand U5521 (N_5521,N_4450,N_4244);
nor U5522 (N_5522,N_4843,N_4374);
nor U5523 (N_5523,N_4415,N_4346);
and U5524 (N_5524,N_4272,N_4717);
and U5525 (N_5525,N_4481,N_4967);
nor U5526 (N_5526,N_4923,N_4644);
nor U5527 (N_5527,N_4459,N_4576);
nand U5528 (N_5528,N_4195,N_4730);
and U5529 (N_5529,N_4484,N_4796);
nor U5530 (N_5530,N_4003,N_4341);
or U5531 (N_5531,N_4466,N_4041);
nand U5532 (N_5532,N_4173,N_4608);
nand U5533 (N_5533,N_4589,N_4038);
nand U5534 (N_5534,N_4310,N_4636);
xnor U5535 (N_5535,N_4752,N_4477);
nand U5536 (N_5536,N_4257,N_4684);
nand U5537 (N_5537,N_4881,N_4792);
nand U5538 (N_5538,N_4957,N_4942);
or U5539 (N_5539,N_4104,N_4288);
and U5540 (N_5540,N_4481,N_4698);
xor U5541 (N_5541,N_4921,N_4309);
nand U5542 (N_5542,N_4389,N_4414);
nand U5543 (N_5543,N_4792,N_4356);
or U5544 (N_5544,N_4407,N_4939);
nor U5545 (N_5545,N_4326,N_4415);
and U5546 (N_5546,N_4652,N_4715);
and U5547 (N_5547,N_4321,N_4466);
and U5548 (N_5548,N_4172,N_4970);
nand U5549 (N_5549,N_4570,N_4965);
nand U5550 (N_5550,N_4081,N_4647);
or U5551 (N_5551,N_4455,N_4435);
or U5552 (N_5552,N_4256,N_4883);
and U5553 (N_5553,N_4655,N_4173);
nand U5554 (N_5554,N_4718,N_4923);
nand U5555 (N_5555,N_4686,N_4700);
and U5556 (N_5556,N_4461,N_4246);
and U5557 (N_5557,N_4352,N_4849);
and U5558 (N_5558,N_4558,N_4215);
or U5559 (N_5559,N_4063,N_4810);
nor U5560 (N_5560,N_4198,N_4486);
nand U5561 (N_5561,N_4615,N_4527);
or U5562 (N_5562,N_4497,N_4972);
or U5563 (N_5563,N_4884,N_4675);
nand U5564 (N_5564,N_4657,N_4800);
nor U5565 (N_5565,N_4414,N_4492);
nor U5566 (N_5566,N_4224,N_4462);
or U5567 (N_5567,N_4145,N_4873);
nand U5568 (N_5568,N_4674,N_4112);
and U5569 (N_5569,N_4550,N_4936);
nand U5570 (N_5570,N_4256,N_4931);
and U5571 (N_5571,N_4827,N_4808);
or U5572 (N_5572,N_4521,N_4381);
and U5573 (N_5573,N_4779,N_4991);
and U5574 (N_5574,N_4216,N_4355);
or U5575 (N_5575,N_4487,N_4817);
nor U5576 (N_5576,N_4479,N_4088);
and U5577 (N_5577,N_4705,N_4957);
nand U5578 (N_5578,N_4839,N_4044);
and U5579 (N_5579,N_4276,N_4560);
and U5580 (N_5580,N_4021,N_4800);
and U5581 (N_5581,N_4712,N_4101);
or U5582 (N_5582,N_4797,N_4550);
nor U5583 (N_5583,N_4665,N_4175);
nand U5584 (N_5584,N_4247,N_4103);
or U5585 (N_5585,N_4488,N_4012);
and U5586 (N_5586,N_4041,N_4788);
nor U5587 (N_5587,N_4496,N_4433);
or U5588 (N_5588,N_4860,N_4788);
and U5589 (N_5589,N_4965,N_4388);
or U5590 (N_5590,N_4277,N_4062);
or U5591 (N_5591,N_4396,N_4374);
or U5592 (N_5592,N_4497,N_4660);
nor U5593 (N_5593,N_4187,N_4855);
or U5594 (N_5594,N_4923,N_4539);
and U5595 (N_5595,N_4749,N_4705);
or U5596 (N_5596,N_4830,N_4387);
or U5597 (N_5597,N_4734,N_4263);
and U5598 (N_5598,N_4285,N_4231);
and U5599 (N_5599,N_4477,N_4376);
and U5600 (N_5600,N_4323,N_4949);
nand U5601 (N_5601,N_4831,N_4099);
or U5602 (N_5602,N_4284,N_4766);
nand U5603 (N_5603,N_4047,N_4733);
or U5604 (N_5604,N_4487,N_4769);
nand U5605 (N_5605,N_4808,N_4043);
nand U5606 (N_5606,N_4029,N_4094);
nor U5607 (N_5607,N_4475,N_4250);
and U5608 (N_5608,N_4405,N_4009);
nand U5609 (N_5609,N_4439,N_4185);
nand U5610 (N_5610,N_4342,N_4757);
nor U5611 (N_5611,N_4369,N_4007);
nor U5612 (N_5612,N_4633,N_4021);
and U5613 (N_5613,N_4299,N_4883);
or U5614 (N_5614,N_4024,N_4749);
and U5615 (N_5615,N_4378,N_4985);
and U5616 (N_5616,N_4984,N_4533);
and U5617 (N_5617,N_4941,N_4197);
and U5618 (N_5618,N_4367,N_4547);
nor U5619 (N_5619,N_4173,N_4414);
nor U5620 (N_5620,N_4201,N_4814);
or U5621 (N_5621,N_4789,N_4883);
and U5622 (N_5622,N_4653,N_4415);
nor U5623 (N_5623,N_4064,N_4421);
nor U5624 (N_5624,N_4399,N_4987);
or U5625 (N_5625,N_4537,N_4995);
and U5626 (N_5626,N_4723,N_4142);
or U5627 (N_5627,N_4387,N_4565);
and U5628 (N_5628,N_4658,N_4136);
and U5629 (N_5629,N_4969,N_4031);
or U5630 (N_5630,N_4910,N_4086);
or U5631 (N_5631,N_4147,N_4008);
or U5632 (N_5632,N_4232,N_4923);
nand U5633 (N_5633,N_4019,N_4509);
or U5634 (N_5634,N_4645,N_4289);
nand U5635 (N_5635,N_4783,N_4964);
nand U5636 (N_5636,N_4096,N_4811);
nor U5637 (N_5637,N_4431,N_4689);
or U5638 (N_5638,N_4103,N_4590);
and U5639 (N_5639,N_4076,N_4639);
or U5640 (N_5640,N_4474,N_4542);
and U5641 (N_5641,N_4963,N_4511);
or U5642 (N_5642,N_4097,N_4523);
and U5643 (N_5643,N_4829,N_4462);
or U5644 (N_5644,N_4846,N_4996);
or U5645 (N_5645,N_4412,N_4340);
and U5646 (N_5646,N_4351,N_4705);
nor U5647 (N_5647,N_4748,N_4255);
or U5648 (N_5648,N_4000,N_4053);
and U5649 (N_5649,N_4696,N_4133);
and U5650 (N_5650,N_4616,N_4736);
and U5651 (N_5651,N_4159,N_4335);
nand U5652 (N_5652,N_4803,N_4752);
or U5653 (N_5653,N_4429,N_4596);
and U5654 (N_5654,N_4432,N_4419);
and U5655 (N_5655,N_4370,N_4768);
xor U5656 (N_5656,N_4262,N_4120);
nand U5657 (N_5657,N_4160,N_4641);
and U5658 (N_5658,N_4961,N_4982);
nand U5659 (N_5659,N_4395,N_4455);
nand U5660 (N_5660,N_4551,N_4999);
nand U5661 (N_5661,N_4594,N_4622);
nor U5662 (N_5662,N_4050,N_4533);
or U5663 (N_5663,N_4454,N_4509);
nor U5664 (N_5664,N_4218,N_4796);
or U5665 (N_5665,N_4124,N_4374);
nand U5666 (N_5666,N_4128,N_4245);
or U5667 (N_5667,N_4001,N_4977);
and U5668 (N_5668,N_4325,N_4090);
or U5669 (N_5669,N_4972,N_4821);
nand U5670 (N_5670,N_4026,N_4383);
and U5671 (N_5671,N_4194,N_4993);
or U5672 (N_5672,N_4517,N_4743);
and U5673 (N_5673,N_4573,N_4497);
nor U5674 (N_5674,N_4332,N_4784);
and U5675 (N_5675,N_4199,N_4820);
nor U5676 (N_5676,N_4851,N_4989);
nand U5677 (N_5677,N_4419,N_4847);
nand U5678 (N_5678,N_4581,N_4084);
nor U5679 (N_5679,N_4608,N_4697);
nor U5680 (N_5680,N_4993,N_4373);
nor U5681 (N_5681,N_4167,N_4583);
nand U5682 (N_5682,N_4511,N_4067);
nand U5683 (N_5683,N_4863,N_4062);
or U5684 (N_5684,N_4274,N_4559);
nor U5685 (N_5685,N_4945,N_4730);
nand U5686 (N_5686,N_4449,N_4355);
nor U5687 (N_5687,N_4885,N_4165);
or U5688 (N_5688,N_4012,N_4315);
nor U5689 (N_5689,N_4959,N_4751);
and U5690 (N_5690,N_4289,N_4295);
nand U5691 (N_5691,N_4350,N_4274);
xnor U5692 (N_5692,N_4121,N_4150);
or U5693 (N_5693,N_4134,N_4996);
or U5694 (N_5694,N_4088,N_4722);
and U5695 (N_5695,N_4230,N_4529);
and U5696 (N_5696,N_4650,N_4103);
nand U5697 (N_5697,N_4349,N_4110);
and U5698 (N_5698,N_4309,N_4039);
or U5699 (N_5699,N_4219,N_4589);
nand U5700 (N_5700,N_4592,N_4255);
nor U5701 (N_5701,N_4048,N_4886);
nor U5702 (N_5702,N_4951,N_4216);
and U5703 (N_5703,N_4527,N_4112);
or U5704 (N_5704,N_4160,N_4230);
or U5705 (N_5705,N_4745,N_4561);
nand U5706 (N_5706,N_4221,N_4681);
nand U5707 (N_5707,N_4981,N_4702);
and U5708 (N_5708,N_4369,N_4856);
and U5709 (N_5709,N_4836,N_4627);
and U5710 (N_5710,N_4448,N_4433);
nand U5711 (N_5711,N_4763,N_4527);
or U5712 (N_5712,N_4102,N_4561);
and U5713 (N_5713,N_4598,N_4301);
or U5714 (N_5714,N_4878,N_4513);
and U5715 (N_5715,N_4708,N_4443);
nand U5716 (N_5716,N_4000,N_4126);
and U5717 (N_5717,N_4832,N_4594);
nand U5718 (N_5718,N_4962,N_4623);
or U5719 (N_5719,N_4354,N_4111);
and U5720 (N_5720,N_4710,N_4877);
and U5721 (N_5721,N_4099,N_4534);
nand U5722 (N_5722,N_4868,N_4278);
nor U5723 (N_5723,N_4302,N_4734);
and U5724 (N_5724,N_4718,N_4137);
nand U5725 (N_5725,N_4829,N_4232);
nand U5726 (N_5726,N_4152,N_4835);
nand U5727 (N_5727,N_4884,N_4053);
or U5728 (N_5728,N_4839,N_4618);
and U5729 (N_5729,N_4082,N_4768);
and U5730 (N_5730,N_4255,N_4519);
and U5731 (N_5731,N_4179,N_4191);
nor U5732 (N_5732,N_4111,N_4656);
nand U5733 (N_5733,N_4793,N_4602);
or U5734 (N_5734,N_4982,N_4339);
or U5735 (N_5735,N_4879,N_4605);
and U5736 (N_5736,N_4236,N_4591);
and U5737 (N_5737,N_4214,N_4859);
and U5738 (N_5738,N_4043,N_4190);
nor U5739 (N_5739,N_4094,N_4288);
nor U5740 (N_5740,N_4150,N_4216);
nand U5741 (N_5741,N_4201,N_4241);
nand U5742 (N_5742,N_4281,N_4136);
or U5743 (N_5743,N_4208,N_4590);
xor U5744 (N_5744,N_4023,N_4398);
nor U5745 (N_5745,N_4797,N_4011);
nor U5746 (N_5746,N_4083,N_4383);
nand U5747 (N_5747,N_4116,N_4717);
or U5748 (N_5748,N_4541,N_4646);
xor U5749 (N_5749,N_4613,N_4229);
nand U5750 (N_5750,N_4089,N_4335);
nand U5751 (N_5751,N_4618,N_4705);
and U5752 (N_5752,N_4956,N_4096);
and U5753 (N_5753,N_4420,N_4448);
nand U5754 (N_5754,N_4172,N_4537);
nor U5755 (N_5755,N_4998,N_4223);
or U5756 (N_5756,N_4110,N_4609);
or U5757 (N_5757,N_4132,N_4608);
and U5758 (N_5758,N_4499,N_4264);
or U5759 (N_5759,N_4640,N_4501);
or U5760 (N_5760,N_4628,N_4049);
nor U5761 (N_5761,N_4329,N_4056);
nand U5762 (N_5762,N_4690,N_4256);
or U5763 (N_5763,N_4662,N_4647);
xnor U5764 (N_5764,N_4029,N_4036);
or U5765 (N_5765,N_4567,N_4531);
or U5766 (N_5766,N_4999,N_4369);
nor U5767 (N_5767,N_4208,N_4023);
nor U5768 (N_5768,N_4742,N_4172);
nand U5769 (N_5769,N_4552,N_4148);
or U5770 (N_5770,N_4230,N_4100);
nand U5771 (N_5771,N_4505,N_4793);
nand U5772 (N_5772,N_4840,N_4176);
or U5773 (N_5773,N_4001,N_4937);
nor U5774 (N_5774,N_4312,N_4205);
nor U5775 (N_5775,N_4476,N_4212);
or U5776 (N_5776,N_4503,N_4661);
and U5777 (N_5777,N_4160,N_4152);
nor U5778 (N_5778,N_4247,N_4052);
nor U5779 (N_5779,N_4702,N_4923);
nand U5780 (N_5780,N_4278,N_4900);
nand U5781 (N_5781,N_4413,N_4457);
or U5782 (N_5782,N_4365,N_4169);
nand U5783 (N_5783,N_4396,N_4006);
nor U5784 (N_5784,N_4386,N_4228);
nand U5785 (N_5785,N_4215,N_4145);
nor U5786 (N_5786,N_4326,N_4226);
nand U5787 (N_5787,N_4409,N_4415);
nand U5788 (N_5788,N_4372,N_4149);
and U5789 (N_5789,N_4906,N_4073);
nor U5790 (N_5790,N_4115,N_4355);
or U5791 (N_5791,N_4706,N_4281);
nand U5792 (N_5792,N_4958,N_4273);
nand U5793 (N_5793,N_4668,N_4366);
and U5794 (N_5794,N_4452,N_4922);
nor U5795 (N_5795,N_4212,N_4790);
and U5796 (N_5796,N_4524,N_4402);
nor U5797 (N_5797,N_4419,N_4028);
nor U5798 (N_5798,N_4662,N_4930);
nor U5799 (N_5799,N_4608,N_4946);
nand U5800 (N_5800,N_4589,N_4249);
and U5801 (N_5801,N_4660,N_4884);
nand U5802 (N_5802,N_4038,N_4563);
or U5803 (N_5803,N_4393,N_4438);
and U5804 (N_5804,N_4260,N_4425);
and U5805 (N_5805,N_4606,N_4140);
or U5806 (N_5806,N_4762,N_4397);
and U5807 (N_5807,N_4396,N_4279);
nand U5808 (N_5808,N_4525,N_4894);
nor U5809 (N_5809,N_4320,N_4478);
nor U5810 (N_5810,N_4007,N_4067);
and U5811 (N_5811,N_4412,N_4611);
nand U5812 (N_5812,N_4178,N_4425);
nor U5813 (N_5813,N_4013,N_4373);
nor U5814 (N_5814,N_4309,N_4209);
or U5815 (N_5815,N_4049,N_4812);
nand U5816 (N_5816,N_4947,N_4608);
and U5817 (N_5817,N_4973,N_4114);
or U5818 (N_5818,N_4757,N_4109);
or U5819 (N_5819,N_4261,N_4588);
nor U5820 (N_5820,N_4329,N_4822);
or U5821 (N_5821,N_4745,N_4619);
or U5822 (N_5822,N_4471,N_4179);
or U5823 (N_5823,N_4151,N_4906);
xnor U5824 (N_5824,N_4393,N_4721);
or U5825 (N_5825,N_4123,N_4232);
and U5826 (N_5826,N_4589,N_4851);
xor U5827 (N_5827,N_4929,N_4977);
nor U5828 (N_5828,N_4091,N_4114);
and U5829 (N_5829,N_4800,N_4877);
and U5830 (N_5830,N_4089,N_4789);
nor U5831 (N_5831,N_4171,N_4713);
nor U5832 (N_5832,N_4420,N_4819);
nand U5833 (N_5833,N_4487,N_4302);
nor U5834 (N_5834,N_4371,N_4620);
and U5835 (N_5835,N_4468,N_4648);
nand U5836 (N_5836,N_4050,N_4678);
and U5837 (N_5837,N_4198,N_4289);
and U5838 (N_5838,N_4464,N_4595);
and U5839 (N_5839,N_4931,N_4409);
and U5840 (N_5840,N_4551,N_4944);
and U5841 (N_5841,N_4592,N_4407);
and U5842 (N_5842,N_4797,N_4663);
and U5843 (N_5843,N_4682,N_4433);
or U5844 (N_5844,N_4765,N_4693);
nor U5845 (N_5845,N_4558,N_4598);
and U5846 (N_5846,N_4268,N_4351);
nor U5847 (N_5847,N_4496,N_4952);
or U5848 (N_5848,N_4888,N_4178);
nor U5849 (N_5849,N_4200,N_4952);
and U5850 (N_5850,N_4290,N_4725);
nor U5851 (N_5851,N_4799,N_4776);
nand U5852 (N_5852,N_4387,N_4029);
and U5853 (N_5853,N_4073,N_4331);
and U5854 (N_5854,N_4497,N_4172);
and U5855 (N_5855,N_4346,N_4312);
nor U5856 (N_5856,N_4912,N_4698);
nand U5857 (N_5857,N_4277,N_4761);
and U5858 (N_5858,N_4764,N_4059);
nand U5859 (N_5859,N_4239,N_4948);
nand U5860 (N_5860,N_4090,N_4254);
or U5861 (N_5861,N_4693,N_4217);
and U5862 (N_5862,N_4445,N_4539);
and U5863 (N_5863,N_4456,N_4204);
and U5864 (N_5864,N_4084,N_4350);
or U5865 (N_5865,N_4577,N_4883);
or U5866 (N_5866,N_4169,N_4021);
nor U5867 (N_5867,N_4612,N_4782);
or U5868 (N_5868,N_4878,N_4112);
nand U5869 (N_5869,N_4380,N_4162);
nand U5870 (N_5870,N_4168,N_4115);
nor U5871 (N_5871,N_4171,N_4633);
and U5872 (N_5872,N_4209,N_4071);
nor U5873 (N_5873,N_4955,N_4374);
and U5874 (N_5874,N_4926,N_4585);
xnor U5875 (N_5875,N_4560,N_4617);
and U5876 (N_5876,N_4996,N_4582);
and U5877 (N_5877,N_4355,N_4849);
or U5878 (N_5878,N_4592,N_4648);
or U5879 (N_5879,N_4482,N_4654);
and U5880 (N_5880,N_4620,N_4394);
and U5881 (N_5881,N_4953,N_4509);
nor U5882 (N_5882,N_4708,N_4404);
or U5883 (N_5883,N_4820,N_4411);
nand U5884 (N_5884,N_4819,N_4010);
or U5885 (N_5885,N_4834,N_4890);
nand U5886 (N_5886,N_4619,N_4004);
and U5887 (N_5887,N_4637,N_4895);
and U5888 (N_5888,N_4953,N_4906);
or U5889 (N_5889,N_4375,N_4827);
or U5890 (N_5890,N_4244,N_4291);
and U5891 (N_5891,N_4590,N_4597);
or U5892 (N_5892,N_4100,N_4713);
and U5893 (N_5893,N_4686,N_4456);
and U5894 (N_5894,N_4003,N_4365);
and U5895 (N_5895,N_4795,N_4348);
xnor U5896 (N_5896,N_4316,N_4332);
nand U5897 (N_5897,N_4173,N_4776);
nand U5898 (N_5898,N_4399,N_4589);
nor U5899 (N_5899,N_4575,N_4887);
or U5900 (N_5900,N_4745,N_4775);
or U5901 (N_5901,N_4180,N_4762);
or U5902 (N_5902,N_4608,N_4826);
nand U5903 (N_5903,N_4931,N_4699);
nand U5904 (N_5904,N_4110,N_4060);
nand U5905 (N_5905,N_4113,N_4731);
and U5906 (N_5906,N_4568,N_4814);
or U5907 (N_5907,N_4001,N_4629);
or U5908 (N_5908,N_4819,N_4156);
and U5909 (N_5909,N_4510,N_4188);
nor U5910 (N_5910,N_4993,N_4920);
nand U5911 (N_5911,N_4981,N_4362);
xor U5912 (N_5912,N_4322,N_4185);
nand U5913 (N_5913,N_4185,N_4133);
nor U5914 (N_5914,N_4352,N_4022);
nand U5915 (N_5915,N_4400,N_4313);
or U5916 (N_5916,N_4021,N_4456);
or U5917 (N_5917,N_4286,N_4577);
or U5918 (N_5918,N_4165,N_4814);
nor U5919 (N_5919,N_4175,N_4908);
nor U5920 (N_5920,N_4607,N_4868);
or U5921 (N_5921,N_4360,N_4286);
nor U5922 (N_5922,N_4231,N_4778);
nand U5923 (N_5923,N_4684,N_4767);
nand U5924 (N_5924,N_4975,N_4058);
nor U5925 (N_5925,N_4354,N_4933);
or U5926 (N_5926,N_4540,N_4215);
nor U5927 (N_5927,N_4346,N_4756);
or U5928 (N_5928,N_4576,N_4196);
nor U5929 (N_5929,N_4721,N_4937);
and U5930 (N_5930,N_4175,N_4891);
nor U5931 (N_5931,N_4759,N_4935);
nor U5932 (N_5932,N_4727,N_4639);
nand U5933 (N_5933,N_4026,N_4893);
and U5934 (N_5934,N_4365,N_4214);
nand U5935 (N_5935,N_4686,N_4177);
nand U5936 (N_5936,N_4572,N_4706);
nor U5937 (N_5937,N_4065,N_4185);
nand U5938 (N_5938,N_4093,N_4493);
or U5939 (N_5939,N_4031,N_4107);
nand U5940 (N_5940,N_4650,N_4421);
nor U5941 (N_5941,N_4081,N_4787);
nand U5942 (N_5942,N_4105,N_4101);
nand U5943 (N_5943,N_4344,N_4742);
and U5944 (N_5944,N_4347,N_4426);
nand U5945 (N_5945,N_4111,N_4209);
or U5946 (N_5946,N_4240,N_4755);
and U5947 (N_5947,N_4089,N_4368);
and U5948 (N_5948,N_4588,N_4649);
nor U5949 (N_5949,N_4689,N_4956);
nand U5950 (N_5950,N_4399,N_4237);
or U5951 (N_5951,N_4716,N_4899);
nand U5952 (N_5952,N_4648,N_4273);
nand U5953 (N_5953,N_4512,N_4237);
or U5954 (N_5954,N_4289,N_4807);
and U5955 (N_5955,N_4640,N_4271);
nor U5956 (N_5956,N_4466,N_4902);
and U5957 (N_5957,N_4305,N_4598);
nor U5958 (N_5958,N_4603,N_4272);
nand U5959 (N_5959,N_4595,N_4112);
and U5960 (N_5960,N_4961,N_4323);
and U5961 (N_5961,N_4467,N_4508);
and U5962 (N_5962,N_4928,N_4611);
nand U5963 (N_5963,N_4283,N_4212);
and U5964 (N_5964,N_4454,N_4366);
nand U5965 (N_5965,N_4774,N_4343);
nand U5966 (N_5966,N_4658,N_4366);
nor U5967 (N_5967,N_4926,N_4985);
and U5968 (N_5968,N_4343,N_4318);
or U5969 (N_5969,N_4457,N_4998);
nor U5970 (N_5970,N_4216,N_4468);
nor U5971 (N_5971,N_4600,N_4958);
and U5972 (N_5972,N_4778,N_4683);
nand U5973 (N_5973,N_4951,N_4857);
or U5974 (N_5974,N_4742,N_4555);
and U5975 (N_5975,N_4586,N_4213);
nand U5976 (N_5976,N_4520,N_4360);
nor U5977 (N_5977,N_4847,N_4668);
nand U5978 (N_5978,N_4483,N_4776);
or U5979 (N_5979,N_4718,N_4710);
nor U5980 (N_5980,N_4351,N_4330);
or U5981 (N_5981,N_4953,N_4602);
or U5982 (N_5982,N_4485,N_4728);
nor U5983 (N_5983,N_4413,N_4745);
and U5984 (N_5984,N_4836,N_4868);
nor U5985 (N_5985,N_4958,N_4200);
and U5986 (N_5986,N_4874,N_4227);
and U5987 (N_5987,N_4110,N_4036);
or U5988 (N_5988,N_4823,N_4619);
and U5989 (N_5989,N_4855,N_4599);
or U5990 (N_5990,N_4768,N_4369);
and U5991 (N_5991,N_4967,N_4777);
or U5992 (N_5992,N_4638,N_4651);
and U5993 (N_5993,N_4937,N_4541);
or U5994 (N_5994,N_4778,N_4019);
or U5995 (N_5995,N_4545,N_4860);
nand U5996 (N_5996,N_4966,N_4686);
or U5997 (N_5997,N_4933,N_4894);
nor U5998 (N_5998,N_4107,N_4932);
nor U5999 (N_5999,N_4270,N_4720);
and U6000 (N_6000,N_5166,N_5240);
nand U6001 (N_6001,N_5974,N_5326);
nand U6002 (N_6002,N_5594,N_5820);
or U6003 (N_6003,N_5484,N_5328);
and U6004 (N_6004,N_5323,N_5712);
and U6005 (N_6005,N_5063,N_5543);
or U6006 (N_6006,N_5727,N_5443);
and U6007 (N_6007,N_5968,N_5438);
nor U6008 (N_6008,N_5315,N_5486);
nand U6009 (N_6009,N_5124,N_5874);
or U6010 (N_6010,N_5203,N_5773);
nor U6011 (N_6011,N_5197,N_5214);
or U6012 (N_6012,N_5939,N_5029);
and U6013 (N_6013,N_5038,N_5905);
nor U6014 (N_6014,N_5147,N_5653);
nor U6015 (N_6015,N_5338,N_5117);
nor U6016 (N_6016,N_5418,N_5944);
nor U6017 (N_6017,N_5686,N_5473);
or U6018 (N_6018,N_5632,N_5841);
and U6019 (N_6019,N_5250,N_5190);
nand U6020 (N_6020,N_5886,N_5591);
nor U6021 (N_6021,N_5707,N_5532);
nor U6022 (N_6022,N_5836,N_5081);
nand U6023 (N_6023,N_5458,N_5657);
and U6024 (N_6024,N_5239,N_5355);
or U6025 (N_6025,N_5281,N_5284);
or U6026 (N_6026,N_5756,N_5131);
and U6027 (N_6027,N_5389,N_5376);
or U6028 (N_6028,N_5118,N_5390);
nor U6029 (N_6029,N_5526,N_5781);
or U6030 (N_6030,N_5701,N_5372);
nor U6031 (N_6031,N_5011,N_5554);
or U6032 (N_6032,N_5784,N_5674);
nor U6033 (N_6033,N_5083,N_5044);
and U6034 (N_6034,N_5794,N_5845);
and U6035 (N_6035,N_5741,N_5377);
or U6036 (N_6036,N_5912,N_5742);
nor U6037 (N_6037,N_5075,N_5154);
and U6038 (N_6038,N_5157,N_5538);
nor U6039 (N_6039,N_5206,N_5425);
and U6040 (N_6040,N_5351,N_5631);
and U6041 (N_6041,N_5960,N_5415);
or U6042 (N_6042,N_5346,N_5212);
or U6043 (N_6043,N_5243,N_5790);
and U6044 (N_6044,N_5204,N_5915);
nand U6045 (N_6045,N_5465,N_5432);
nor U6046 (N_6046,N_5302,N_5942);
or U6047 (N_6047,N_5463,N_5614);
and U6048 (N_6048,N_5381,N_5142);
nor U6049 (N_6049,N_5347,N_5812);
and U6050 (N_6050,N_5217,N_5667);
nand U6051 (N_6051,N_5881,N_5399);
and U6052 (N_6052,N_5004,N_5472);
nor U6053 (N_6053,N_5468,N_5109);
or U6054 (N_6054,N_5609,N_5548);
and U6055 (N_6055,N_5183,N_5477);
or U6056 (N_6056,N_5179,N_5344);
or U6057 (N_6057,N_5625,N_5489);
nor U6058 (N_6058,N_5870,N_5890);
nor U6059 (N_6059,N_5746,N_5151);
nor U6060 (N_6060,N_5138,N_5963);
and U6061 (N_6061,N_5551,N_5534);
nor U6062 (N_6062,N_5184,N_5170);
nand U6063 (N_6063,N_5518,N_5656);
nor U6064 (N_6064,N_5012,N_5149);
nand U6065 (N_6065,N_5034,N_5134);
nor U6066 (N_6066,N_5815,N_5775);
and U6067 (N_6067,N_5826,N_5491);
nand U6068 (N_6068,N_5878,N_5860);
or U6069 (N_6069,N_5635,N_5037);
or U6070 (N_6070,N_5041,N_5076);
or U6071 (N_6071,N_5242,N_5854);
or U6072 (N_6072,N_5357,N_5530);
nand U6073 (N_6073,N_5201,N_5174);
nor U6074 (N_6074,N_5867,N_5764);
or U6075 (N_6075,N_5414,N_5064);
nand U6076 (N_6076,N_5908,N_5492);
nand U6077 (N_6077,N_5618,N_5364);
or U6078 (N_6078,N_5226,N_5132);
or U6079 (N_6079,N_5630,N_5622);
nand U6080 (N_6080,N_5261,N_5977);
or U6081 (N_6081,N_5780,N_5430);
and U6082 (N_6082,N_5036,N_5280);
and U6083 (N_6083,N_5649,N_5298);
nor U6084 (N_6084,N_5487,N_5767);
nor U6085 (N_6085,N_5506,N_5545);
nand U6086 (N_6086,N_5439,N_5366);
nand U6087 (N_6087,N_5185,N_5453);
and U6088 (N_6088,N_5804,N_5525);
or U6089 (N_6089,N_5039,N_5988);
and U6090 (N_6090,N_5019,N_5168);
nor U6091 (N_6091,N_5795,N_5792);
and U6092 (N_6092,N_5768,N_5931);
or U6093 (N_6093,N_5807,N_5195);
nand U6094 (N_6094,N_5521,N_5313);
nand U6095 (N_6095,N_5398,N_5803);
xnor U6096 (N_6096,N_5749,N_5650);
and U6097 (N_6097,N_5309,N_5289);
or U6098 (N_6098,N_5581,N_5924);
or U6099 (N_6099,N_5842,N_5436);
nor U6100 (N_6100,N_5215,N_5579);
or U6101 (N_6101,N_5175,N_5838);
or U6102 (N_6102,N_5735,N_5725);
or U6103 (N_6103,N_5176,N_5615);
and U6104 (N_6104,N_5702,N_5995);
or U6105 (N_6105,N_5342,N_5213);
or U6106 (N_6106,N_5028,N_5847);
or U6107 (N_6107,N_5208,N_5013);
or U6108 (N_6108,N_5139,N_5646);
or U6109 (N_6109,N_5852,N_5816);
and U6110 (N_6110,N_5503,N_5979);
and U6111 (N_6111,N_5726,N_5071);
and U6112 (N_6112,N_5613,N_5504);
nor U6113 (N_6113,N_5937,N_5736);
nor U6114 (N_6114,N_5483,N_5370);
nand U6115 (N_6115,N_5222,N_5435);
nand U6116 (N_6116,N_5066,N_5994);
nand U6117 (N_6117,N_5909,N_5638);
nand U6118 (N_6118,N_5893,N_5959);
nor U6119 (N_6119,N_5588,N_5100);
and U6120 (N_6120,N_5047,N_5691);
nor U6121 (N_6121,N_5368,N_5456);
or U6122 (N_6122,N_5745,N_5099);
nand U6123 (N_6123,N_5282,N_5546);
nor U6124 (N_6124,N_5297,N_5263);
or U6125 (N_6125,N_5798,N_5003);
nor U6126 (N_6126,N_5050,N_5896);
and U6127 (N_6127,N_5200,N_5428);
nand U6128 (N_6128,N_5868,N_5125);
and U6129 (N_6129,N_5395,N_5835);
and U6130 (N_6130,N_5286,N_5998);
and U6131 (N_6131,N_5837,N_5306);
or U6132 (N_6132,N_5949,N_5394);
and U6133 (N_6133,N_5008,N_5021);
or U6134 (N_6134,N_5945,N_5528);
and U6135 (N_6135,N_5152,N_5000);
and U6136 (N_6136,N_5058,N_5387);
and U6137 (N_6137,N_5252,N_5855);
nor U6138 (N_6138,N_5605,N_5552);
or U6139 (N_6139,N_5336,N_5329);
nor U6140 (N_6140,N_5556,N_5163);
nand U6141 (N_6141,N_5007,N_5762);
nand U6142 (N_6142,N_5822,N_5333);
or U6143 (N_6143,N_5469,N_5073);
nor U6144 (N_6144,N_5207,N_5694);
nor U6145 (N_6145,N_5724,N_5412);
or U6146 (N_6146,N_5950,N_5692);
or U6147 (N_6147,N_5516,N_5661);
or U6148 (N_6148,N_5902,N_5951);
and U6149 (N_6149,N_5771,N_5916);
nor U6150 (N_6150,N_5713,N_5062);
nand U6151 (N_6151,N_5573,N_5763);
nand U6152 (N_6152,N_5932,N_5311);
nor U6153 (N_6153,N_5723,N_5734);
xnor U6154 (N_6154,N_5660,N_5305);
nor U6155 (N_6155,N_5512,N_5940);
xnor U6156 (N_6156,N_5006,N_5269);
or U6157 (N_6157,N_5885,N_5666);
nor U6158 (N_6158,N_5793,N_5259);
nand U6159 (N_6159,N_5380,N_5113);
and U6160 (N_6160,N_5017,N_5777);
nor U6161 (N_6161,N_5172,N_5408);
nand U6162 (N_6162,N_5108,N_5929);
and U6163 (N_6163,N_5522,N_5900);
nand U6164 (N_6164,N_5189,N_5400);
nor U6165 (N_6165,N_5907,N_5730);
and U6166 (N_6166,N_5230,N_5975);
nor U6167 (N_6167,N_5218,N_5043);
xnor U6168 (N_6168,N_5301,N_5386);
and U6169 (N_6169,N_5488,N_5110);
nand U6170 (N_6170,N_5446,N_5859);
nand U6171 (N_6171,N_5140,N_5508);
nor U6172 (N_6172,N_5085,N_5608);
nor U6173 (N_6173,N_5757,N_5426);
nand U6174 (N_6174,N_5153,N_5875);
or U6175 (N_6175,N_5843,N_5278);
nor U6176 (N_6176,N_5105,N_5801);
and U6177 (N_6177,N_5126,N_5624);
and U6178 (N_6178,N_5930,N_5397);
nand U6179 (N_6179,N_5920,N_5334);
and U6180 (N_6180,N_5884,N_5481);
or U6181 (N_6181,N_5211,N_5514);
nor U6182 (N_6182,N_5987,N_5090);
nand U6183 (N_6183,N_5722,N_5580);
nand U6184 (N_6184,N_5232,N_5541);
or U6185 (N_6185,N_5349,N_5634);
nor U6186 (N_6186,N_5621,N_5510);
or U6187 (N_6187,N_5403,N_5533);
and U6188 (N_6188,N_5059,N_5283);
and U6189 (N_6189,N_5501,N_5671);
nand U6190 (N_6190,N_5141,N_5866);
or U6191 (N_6191,N_5655,N_5693);
nand U6192 (N_6192,N_5084,N_5448);
and U6193 (N_6193,N_5358,N_5561);
or U6194 (N_6194,N_5231,N_5562);
or U6195 (N_6195,N_5070,N_5602);
nand U6196 (N_6196,N_5955,N_5619);
nor U6197 (N_6197,N_5547,N_5848);
nor U6198 (N_6198,N_5310,N_5558);
and U6199 (N_6199,N_5502,N_5479);
and U6200 (N_6200,N_5799,N_5710);
nand U6201 (N_6201,N_5873,N_5620);
nand U6202 (N_6202,N_5894,N_5679);
nor U6203 (N_6203,N_5889,N_5941);
nand U6204 (N_6204,N_5228,N_5042);
nor U6205 (N_6205,N_5511,N_5500);
nor U6206 (N_6206,N_5193,N_5402);
or U6207 (N_6207,N_5341,N_5367);
nand U6208 (N_6208,N_5985,N_5589);
nand U6209 (N_6209,N_5288,N_5449);
or U6210 (N_6210,N_5419,N_5753);
or U6211 (N_6211,N_5715,N_5160);
nor U6212 (N_6212,N_5169,N_5352);
nor U6213 (N_6213,N_5583,N_5564);
and U6214 (N_6214,N_5524,N_5089);
or U6215 (N_6215,N_5292,N_5743);
nor U6216 (N_6216,N_5056,N_5300);
nor U6217 (N_6217,N_5237,N_5122);
and U6218 (N_6218,N_5354,N_5485);
nand U6219 (N_6219,N_5652,N_5221);
or U6220 (N_6220,N_5143,N_5965);
nand U6221 (N_6221,N_5135,N_5892);
nor U6222 (N_6222,N_5628,N_5586);
and U6223 (N_6223,N_5369,N_5235);
and U6224 (N_6224,N_5331,N_5277);
and U6225 (N_6225,N_5274,N_5279);
nor U6226 (N_6226,N_5199,N_5791);
nand U6227 (N_6227,N_5429,N_5382);
nand U6228 (N_6228,N_5891,N_5356);
and U6229 (N_6229,N_5769,N_5265);
and U6230 (N_6230,N_5392,N_5688);
nor U6231 (N_6231,N_5180,N_5427);
nor U6232 (N_6232,N_5009,N_5244);
nand U6233 (N_6233,N_5721,N_5754);
nand U6234 (N_6234,N_5928,N_5317);
or U6235 (N_6235,N_5079,N_5680);
nor U6236 (N_6236,N_5923,N_5695);
nor U6237 (N_6237,N_5805,N_5496);
and U6238 (N_6238,N_5598,N_5747);
or U6239 (N_6239,N_5321,N_5636);
or U6240 (N_6240,N_5840,N_5434);
nand U6241 (N_6241,N_5689,N_5708);
nand U6242 (N_6242,N_5010,N_5751);
nor U6243 (N_6243,N_5953,N_5895);
or U6244 (N_6244,N_5360,N_5457);
and U6245 (N_6245,N_5922,N_5054);
nand U6246 (N_6246,N_5999,N_5146);
nor U6247 (N_6247,N_5103,N_5729);
or U6248 (N_6248,N_5983,N_5626);
nand U6249 (N_6249,N_5061,N_5563);
nor U6250 (N_6250,N_5971,N_5032);
nor U6251 (N_6251,N_5603,N_5952);
and U6252 (N_6252,N_5850,N_5474);
or U6253 (N_6253,N_5253,N_5567);
nor U6254 (N_6254,N_5844,N_5452);
nor U6255 (N_6255,N_5744,N_5188);
nor U6256 (N_6256,N_5171,N_5460);
and U6257 (N_6257,N_5264,N_5353);
and U6258 (N_6258,N_5993,N_5023);
and U6259 (N_6259,N_5320,N_5144);
or U6260 (N_6260,N_5832,N_5828);
and U6261 (N_6261,N_5196,N_5925);
and U6262 (N_6262,N_5102,N_5610);
or U6263 (N_6263,N_5719,N_5733);
nand U6264 (N_6264,N_5248,N_5121);
and U6265 (N_6265,N_5943,N_5165);
or U6266 (N_6266,N_5833,N_5571);
or U6267 (N_6267,N_5779,N_5304);
nand U6268 (N_6268,N_5969,N_5879);
or U6269 (N_6269,N_5527,N_5093);
and U6270 (N_6270,N_5665,N_5825);
and U6271 (N_6271,N_5440,N_5823);
xnor U6272 (N_6272,N_5480,N_5967);
nor U6273 (N_6273,N_5623,N_5576);
xor U6274 (N_6274,N_5658,N_5542);
nor U6275 (N_6275,N_5883,N_5027);
or U6276 (N_6276,N_5130,N_5475);
nor U6277 (N_6277,N_5509,N_5187);
and U6278 (N_6278,N_5557,N_5216);
and U6279 (N_6279,N_5470,N_5464);
or U6280 (N_6280,N_5536,N_5568);
and U6281 (N_6281,N_5919,N_5155);
or U6282 (N_6282,N_5574,N_5572);
or U6283 (N_6283,N_5441,N_5830);
nor U6284 (N_6284,N_5811,N_5544);
nand U6285 (N_6285,N_5645,N_5150);
nand U6286 (N_6286,N_5690,N_5220);
and U6287 (N_6287,N_5072,N_5926);
nand U6288 (N_6288,N_5782,N_5015);
nand U6289 (N_6289,N_5080,N_5651);
or U6290 (N_6290,N_5864,N_5587);
nor U6291 (N_6291,N_5194,N_5114);
or U6292 (N_6292,N_5697,N_5405);
nor U6293 (N_6293,N_5271,N_5851);
nor U6294 (N_6294,N_5770,N_5772);
or U6295 (N_6295,N_5976,N_5225);
nor U6296 (N_6296,N_5560,N_5322);
nor U6297 (N_6297,N_5810,N_5787);
or U6298 (N_6298,N_5290,N_5716);
and U6299 (N_6299,N_5330,N_5343);
nand U6300 (N_6300,N_5664,N_5888);
and U6301 (N_6301,N_5997,N_5123);
nor U6302 (N_6302,N_5391,N_5378);
and U6303 (N_6303,N_5684,N_5094);
or U6304 (N_6304,N_5299,N_5088);
or U6305 (N_6305,N_5128,N_5934);
and U6306 (N_6306,N_5540,N_5324);
xor U6307 (N_6307,N_5565,N_5026);
nor U6308 (N_6308,N_5872,N_5633);
xor U6309 (N_6309,N_5296,N_5956);
or U6310 (N_6310,N_5946,N_5120);
nand U6311 (N_6311,N_5858,N_5936);
nor U6312 (N_6312,N_5682,N_5910);
nor U6313 (N_6313,N_5535,N_5307);
or U6314 (N_6314,N_5383,N_5115);
and U6315 (N_6315,N_5601,N_5853);
nand U6316 (N_6316,N_5992,N_5025);
or U6317 (N_6317,N_5861,N_5752);
nor U6318 (N_6318,N_5709,N_5718);
nor U6319 (N_6319,N_5363,N_5046);
or U6320 (N_6320,N_5494,N_5857);
or U6321 (N_6321,N_5670,N_5732);
nand U6322 (N_6322,N_5318,N_5935);
nand U6323 (N_6323,N_5549,N_5877);
nor U6324 (N_6324,N_5871,N_5700);
nor U6325 (N_6325,N_5880,N_5906);
nand U6326 (N_6326,N_5566,N_5433);
nand U6327 (N_6327,N_5814,N_5611);
and U6328 (N_6328,N_5173,N_5086);
nand U6329 (N_6329,N_5761,N_5918);
nand U6330 (N_6330,N_5824,N_5164);
or U6331 (N_6331,N_5699,N_5629);
nor U6332 (N_6332,N_5437,N_5097);
or U6333 (N_6333,N_5839,N_5785);
nand U6334 (N_6334,N_5681,N_5249);
or U6335 (N_6335,N_5531,N_5595);
and U6336 (N_6336,N_5597,N_5158);
nand U6337 (N_6337,N_5031,N_5495);
or U6338 (N_6338,N_5018,N_5033);
nand U6339 (N_6339,N_5766,N_5513);
nor U6340 (N_6340,N_5466,N_5731);
nor U6341 (N_6341,N_5182,N_5800);
or U6342 (N_6342,N_5238,N_5698);
and U6343 (N_6343,N_5933,N_5467);
or U6344 (N_6344,N_5233,N_5789);
and U6345 (N_6345,N_5325,N_5584);
nor U6346 (N_6346,N_5001,N_5846);
xor U6347 (N_6347,N_5648,N_5676);
or U6348 (N_6348,N_5388,N_5738);
and U6349 (N_6349,N_5964,N_5234);
or U6350 (N_6350,N_5593,N_5641);
and U6351 (N_6351,N_5411,N_5592);
or U6352 (N_6352,N_5981,N_5616);
or U6353 (N_6353,N_5303,N_5984);
and U6354 (N_6354,N_5074,N_5393);
and U6355 (N_6355,N_5817,N_5519);
or U6356 (N_6356,N_5654,N_5406);
or U6357 (N_6357,N_5555,N_5339);
nand U6358 (N_6358,N_5396,N_5260);
or U6359 (N_6359,N_5258,N_5424);
nand U6360 (N_6360,N_5312,N_5821);
nand U6361 (N_6361,N_5482,N_5082);
nand U6362 (N_6362,N_5161,N_5760);
nor U6363 (N_6363,N_5314,N_5087);
nor U6364 (N_6364,N_5783,N_5365);
nand U6365 (N_6365,N_5947,N_5268);
and U6366 (N_6366,N_5499,N_5717);
nand U6367 (N_6367,N_5578,N_5060);
and U6368 (N_6368,N_5737,N_5181);
nand U6369 (N_6369,N_5903,N_5529);
or U6370 (N_6370,N_5991,N_5921);
nand U6371 (N_6371,N_5416,N_5219);
or U6372 (N_6372,N_5714,N_5677);
nand U6373 (N_6373,N_5678,N_5270);
nand U6374 (N_6374,N_5672,N_5319);
or U6375 (N_6375,N_5711,N_5407);
nor U6376 (N_6376,N_5178,N_5797);
nand U6377 (N_6377,N_5927,N_5639);
or U6378 (N_6378,N_5030,N_5246);
or U6379 (N_6379,N_5740,N_5668);
nor U6380 (N_6380,N_5644,N_5198);
nor U6381 (N_6381,N_5640,N_5241);
nand U6382 (N_6382,N_5040,N_5119);
and U6383 (N_6383,N_5162,N_5459);
or U6384 (N_6384,N_5673,N_5014);
and U6385 (N_6385,N_5917,N_5765);
and U6386 (N_6386,N_5254,N_5167);
or U6387 (N_6387,N_5361,N_5862);
nor U6388 (N_6388,N_5539,N_5111);
nand U6389 (N_6389,N_5148,N_5016);
nand U6390 (N_6390,N_5335,N_5266);
nor U6391 (N_6391,N_5092,N_5819);
nand U6392 (N_6392,N_5421,N_5829);
nand U6393 (N_6393,N_5970,N_5505);
nand U6394 (N_6394,N_5451,N_5444);
or U6395 (N_6395,N_5057,N_5642);
and U6396 (N_6396,N_5982,N_5827);
and U6397 (N_6397,N_5116,N_5156);
nand U6398 (N_6398,N_5582,N_5091);
nor U6399 (N_6399,N_5759,N_5989);
nor U6400 (N_6400,N_5461,N_5256);
and U6401 (N_6401,N_5683,N_5024);
or U6402 (N_6402,N_5869,N_5192);
nor U6403 (N_6403,N_5275,N_5898);
or U6404 (N_6404,N_5055,N_5758);
and U6405 (N_6405,N_5417,N_5209);
or U6406 (N_6406,N_5020,N_5669);
or U6407 (N_6407,N_5276,N_5604);
xnor U6408 (N_6408,N_5786,N_5515);
nand U6409 (N_6409,N_5136,N_5617);
nand U6410 (N_6410,N_5447,N_5612);
nor U6411 (N_6411,N_5590,N_5863);
nor U6412 (N_6412,N_5308,N_5607);
nand U6413 (N_6413,N_5569,N_5413);
xnor U6414 (N_6414,N_5384,N_5454);
and U6415 (N_6415,N_5938,N_5455);
or U6416 (N_6416,N_5647,N_5813);
nor U6417 (N_6417,N_5112,N_5005);
nor U6418 (N_6418,N_5159,N_5954);
and U6419 (N_6419,N_5065,N_5223);
or U6420 (N_6420,N_5101,N_5627);
or U6421 (N_6421,N_5901,N_5049);
nand U6422 (N_6422,N_5808,N_5887);
nor U6423 (N_6423,N_5606,N_5705);
nand U6424 (N_6424,N_5051,N_5996);
or U6425 (N_6425,N_5359,N_5137);
or U6426 (N_6426,N_5267,N_5078);
nand U6427 (N_6427,N_5599,N_5273);
or U6428 (N_6428,N_5404,N_5520);
and U6429 (N_6429,N_5778,N_5776);
nand U6430 (N_6430,N_5373,N_5272);
and U6431 (N_6431,N_5553,N_5913);
nor U6432 (N_6432,N_5507,N_5973);
and U6433 (N_6433,N_5471,N_5236);
or U6434 (N_6434,N_5362,N_5659);
xor U6435 (N_6435,N_5077,N_5327);
xor U6436 (N_6436,N_5002,N_5637);
and U6437 (N_6437,N_5375,N_5145);
or U6438 (N_6438,N_5053,N_5247);
nor U6439 (N_6439,N_5420,N_5685);
nand U6440 (N_6440,N_5911,N_5497);
or U6441 (N_6441,N_5127,N_5035);
nor U6442 (N_6442,N_5834,N_5229);
and U6443 (N_6443,N_5914,N_5739);
or U6444 (N_6444,N_5978,N_5202);
nor U6445 (N_6445,N_5098,N_5818);
nand U6446 (N_6446,N_5423,N_5774);
nand U6447 (N_6447,N_5980,N_5227);
or U6448 (N_6448,N_5831,N_5962);
nand U6449 (N_6449,N_5374,N_5191);
or U6450 (N_6450,N_5720,N_5663);
and U6451 (N_6451,N_5517,N_5177);
or U6452 (N_6452,N_5133,N_5245);
and U6453 (N_6453,N_5899,N_5550);
and U6454 (N_6454,N_5350,N_5961);
or U6455 (N_6455,N_5728,N_5379);
nand U6456 (N_6456,N_5431,N_5210);
nand U6457 (N_6457,N_5643,N_5371);
nor U6458 (N_6458,N_5291,N_5285);
or U6459 (N_6459,N_5255,N_5957);
nor U6460 (N_6460,N_5069,N_5972);
nor U6461 (N_6461,N_5490,N_5048);
and U6462 (N_6462,N_5107,N_5704);
nor U6463 (N_6463,N_5401,N_5600);
and U6464 (N_6464,N_5570,N_5445);
xor U6465 (N_6465,N_5340,N_5293);
or U6466 (N_6466,N_5748,N_5675);
nor U6467 (N_6467,N_5948,N_5068);
nand U6468 (N_6468,N_5865,N_5493);
and U6469 (N_6469,N_5856,N_5287);
nand U6470 (N_6470,N_5523,N_5958);
nor U6471 (N_6471,N_5966,N_5257);
nand U6472 (N_6472,N_5385,N_5990);
nor U6473 (N_6473,N_5095,N_5696);
or U6474 (N_6474,N_5849,N_5802);
nor U6475 (N_6475,N_5410,N_5332);
nand U6476 (N_6476,N_5662,N_5755);
and U6477 (N_6477,N_5462,N_5205);
or U6478 (N_6478,N_5904,N_5345);
or U6479 (N_6479,N_5294,N_5045);
and U6480 (N_6480,N_5251,N_5897);
or U6481 (N_6481,N_5096,N_5806);
or U6482 (N_6482,N_5067,N_5596);
nor U6483 (N_6483,N_5262,N_5788);
and U6484 (N_6484,N_5295,N_5348);
and U6485 (N_6485,N_5478,N_5104);
or U6486 (N_6486,N_5316,N_5129);
nor U6487 (N_6487,N_5337,N_5986);
or U6488 (N_6488,N_5703,N_5224);
nand U6489 (N_6489,N_5585,N_5106);
and U6490 (N_6490,N_5575,N_5422);
or U6491 (N_6491,N_5559,N_5882);
nand U6492 (N_6492,N_5442,N_5409);
nand U6493 (N_6493,N_5186,N_5476);
or U6494 (N_6494,N_5706,N_5809);
or U6495 (N_6495,N_5687,N_5577);
nor U6496 (N_6496,N_5498,N_5022);
or U6497 (N_6497,N_5876,N_5750);
nand U6498 (N_6498,N_5796,N_5052);
or U6499 (N_6499,N_5537,N_5450);
or U6500 (N_6500,N_5811,N_5661);
and U6501 (N_6501,N_5301,N_5605);
and U6502 (N_6502,N_5321,N_5697);
nor U6503 (N_6503,N_5886,N_5912);
or U6504 (N_6504,N_5956,N_5634);
or U6505 (N_6505,N_5313,N_5569);
nand U6506 (N_6506,N_5038,N_5352);
nand U6507 (N_6507,N_5853,N_5729);
nor U6508 (N_6508,N_5117,N_5686);
or U6509 (N_6509,N_5133,N_5072);
and U6510 (N_6510,N_5607,N_5085);
or U6511 (N_6511,N_5198,N_5849);
and U6512 (N_6512,N_5604,N_5175);
nor U6513 (N_6513,N_5908,N_5375);
and U6514 (N_6514,N_5971,N_5775);
and U6515 (N_6515,N_5099,N_5416);
or U6516 (N_6516,N_5210,N_5948);
nor U6517 (N_6517,N_5043,N_5839);
and U6518 (N_6518,N_5384,N_5636);
nand U6519 (N_6519,N_5896,N_5261);
and U6520 (N_6520,N_5111,N_5359);
and U6521 (N_6521,N_5256,N_5102);
nand U6522 (N_6522,N_5261,N_5745);
and U6523 (N_6523,N_5481,N_5888);
nand U6524 (N_6524,N_5663,N_5919);
nand U6525 (N_6525,N_5674,N_5321);
nand U6526 (N_6526,N_5659,N_5484);
and U6527 (N_6527,N_5334,N_5855);
nor U6528 (N_6528,N_5046,N_5879);
or U6529 (N_6529,N_5044,N_5931);
nor U6530 (N_6530,N_5830,N_5840);
nor U6531 (N_6531,N_5274,N_5658);
or U6532 (N_6532,N_5392,N_5090);
and U6533 (N_6533,N_5367,N_5340);
or U6534 (N_6534,N_5001,N_5538);
and U6535 (N_6535,N_5863,N_5156);
and U6536 (N_6536,N_5796,N_5394);
and U6537 (N_6537,N_5523,N_5280);
and U6538 (N_6538,N_5074,N_5709);
and U6539 (N_6539,N_5442,N_5046);
nand U6540 (N_6540,N_5446,N_5131);
nor U6541 (N_6541,N_5946,N_5087);
and U6542 (N_6542,N_5002,N_5287);
and U6543 (N_6543,N_5708,N_5173);
xnor U6544 (N_6544,N_5084,N_5008);
nand U6545 (N_6545,N_5587,N_5821);
nor U6546 (N_6546,N_5503,N_5889);
and U6547 (N_6547,N_5280,N_5606);
nor U6548 (N_6548,N_5351,N_5013);
and U6549 (N_6549,N_5379,N_5057);
and U6550 (N_6550,N_5403,N_5135);
and U6551 (N_6551,N_5535,N_5244);
or U6552 (N_6552,N_5776,N_5654);
xnor U6553 (N_6553,N_5779,N_5699);
or U6554 (N_6554,N_5916,N_5453);
and U6555 (N_6555,N_5960,N_5815);
nand U6556 (N_6556,N_5829,N_5082);
nand U6557 (N_6557,N_5638,N_5677);
nand U6558 (N_6558,N_5215,N_5016);
nand U6559 (N_6559,N_5064,N_5240);
nand U6560 (N_6560,N_5175,N_5068);
nand U6561 (N_6561,N_5590,N_5726);
and U6562 (N_6562,N_5283,N_5966);
nand U6563 (N_6563,N_5294,N_5878);
or U6564 (N_6564,N_5815,N_5414);
or U6565 (N_6565,N_5374,N_5037);
nor U6566 (N_6566,N_5078,N_5407);
nor U6567 (N_6567,N_5936,N_5318);
nor U6568 (N_6568,N_5047,N_5185);
and U6569 (N_6569,N_5636,N_5609);
nand U6570 (N_6570,N_5129,N_5574);
or U6571 (N_6571,N_5833,N_5630);
nor U6572 (N_6572,N_5610,N_5885);
nand U6573 (N_6573,N_5489,N_5245);
or U6574 (N_6574,N_5085,N_5349);
nor U6575 (N_6575,N_5543,N_5435);
xor U6576 (N_6576,N_5196,N_5100);
nor U6577 (N_6577,N_5442,N_5679);
and U6578 (N_6578,N_5557,N_5111);
nor U6579 (N_6579,N_5537,N_5885);
nor U6580 (N_6580,N_5464,N_5504);
or U6581 (N_6581,N_5490,N_5810);
or U6582 (N_6582,N_5657,N_5953);
or U6583 (N_6583,N_5135,N_5097);
nor U6584 (N_6584,N_5129,N_5602);
nor U6585 (N_6585,N_5620,N_5582);
nand U6586 (N_6586,N_5623,N_5703);
nor U6587 (N_6587,N_5376,N_5380);
or U6588 (N_6588,N_5721,N_5085);
or U6589 (N_6589,N_5087,N_5376);
or U6590 (N_6590,N_5274,N_5213);
nor U6591 (N_6591,N_5689,N_5754);
nand U6592 (N_6592,N_5174,N_5227);
or U6593 (N_6593,N_5220,N_5891);
or U6594 (N_6594,N_5963,N_5596);
and U6595 (N_6595,N_5519,N_5268);
nor U6596 (N_6596,N_5750,N_5828);
or U6597 (N_6597,N_5157,N_5435);
and U6598 (N_6598,N_5317,N_5015);
or U6599 (N_6599,N_5804,N_5241);
or U6600 (N_6600,N_5139,N_5713);
and U6601 (N_6601,N_5110,N_5449);
and U6602 (N_6602,N_5368,N_5403);
nand U6603 (N_6603,N_5781,N_5549);
and U6604 (N_6604,N_5195,N_5237);
or U6605 (N_6605,N_5624,N_5788);
nor U6606 (N_6606,N_5374,N_5073);
or U6607 (N_6607,N_5781,N_5872);
nor U6608 (N_6608,N_5844,N_5666);
and U6609 (N_6609,N_5700,N_5737);
and U6610 (N_6610,N_5192,N_5642);
nor U6611 (N_6611,N_5357,N_5747);
and U6612 (N_6612,N_5066,N_5230);
nand U6613 (N_6613,N_5611,N_5840);
nand U6614 (N_6614,N_5039,N_5340);
or U6615 (N_6615,N_5299,N_5774);
nor U6616 (N_6616,N_5698,N_5616);
and U6617 (N_6617,N_5705,N_5894);
nor U6618 (N_6618,N_5784,N_5783);
or U6619 (N_6619,N_5552,N_5578);
or U6620 (N_6620,N_5767,N_5810);
nor U6621 (N_6621,N_5561,N_5810);
nand U6622 (N_6622,N_5202,N_5226);
and U6623 (N_6623,N_5292,N_5788);
and U6624 (N_6624,N_5689,N_5673);
and U6625 (N_6625,N_5486,N_5431);
nand U6626 (N_6626,N_5626,N_5514);
nor U6627 (N_6627,N_5822,N_5421);
or U6628 (N_6628,N_5382,N_5477);
nand U6629 (N_6629,N_5353,N_5251);
nor U6630 (N_6630,N_5968,N_5523);
and U6631 (N_6631,N_5553,N_5117);
nor U6632 (N_6632,N_5281,N_5452);
and U6633 (N_6633,N_5950,N_5670);
or U6634 (N_6634,N_5141,N_5482);
nand U6635 (N_6635,N_5245,N_5626);
and U6636 (N_6636,N_5977,N_5036);
and U6637 (N_6637,N_5870,N_5940);
or U6638 (N_6638,N_5248,N_5615);
nor U6639 (N_6639,N_5188,N_5231);
or U6640 (N_6640,N_5039,N_5761);
nand U6641 (N_6641,N_5967,N_5763);
nor U6642 (N_6642,N_5717,N_5113);
nor U6643 (N_6643,N_5739,N_5614);
and U6644 (N_6644,N_5549,N_5448);
nand U6645 (N_6645,N_5233,N_5834);
nor U6646 (N_6646,N_5934,N_5805);
and U6647 (N_6647,N_5863,N_5565);
xor U6648 (N_6648,N_5536,N_5010);
xor U6649 (N_6649,N_5870,N_5982);
nand U6650 (N_6650,N_5491,N_5587);
and U6651 (N_6651,N_5773,N_5782);
nor U6652 (N_6652,N_5244,N_5766);
nand U6653 (N_6653,N_5131,N_5311);
and U6654 (N_6654,N_5689,N_5734);
or U6655 (N_6655,N_5451,N_5022);
nand U6656 (N_6656,N_5790,N_5170);
or U6657 (N_6657,N_5222,N_5520);
and U6658 (N_6658,N_5981,N_5180);
and U6659 (N_6659,N_5895,N_5540);
or U6660 (N_6660,N_5556,N_5860);
nand U6661 (N_6661,N_5985,N_5586);
or U6662 (N_6662,N_5608,N_5750);
or U6663 (N_6663,N_5732,N_5011);
or U6664 (N_6664,N_5778,N_5154);
and U6665 (N_6665,N_5567,N_5950);
or U6666 (N_6666,N_5272,N_5748);
nand U6667 (N_6667,N_5285,N_5917);
nand U6668 (N_6668,N_5290,N_5000);
or U6669 (N_6669,N_5575,N_5221);
or U6670 (N_6670,N_5451,N_5537);
nor U6671 (N_6671,N_5623,N_5544);
or U6672 (N_6672,N_5007,N_5042);
and U6673 (N_6673,N_5421,N_5141);
nand U6674 (N_6674,N_5552,N_5295);
or U6675 (N_6675,N_5639,N_5913);
nor U6676 (N_6676,N_5289,N_5415);
or U6677 (N_6677,N_5930,N_5906);
and U6678 (N_6678,N_5701,N_5797);
nand U6679 (N_6679,N_5109,N_5808);
and U6680 (N_6680,N_5119,N_5413);
and U6681 (N_6681,N_5091,N_5161);
and U6682 (N_6682,N_5977,N_5999);
nor U6683 (N_6683,N_5650,N_5933);
or U6684 (N_6684,N_5838,N_5493);
or U6685 (N_6685,N_5200,N_5440);
nor U6686 (N_6686,N_5050,N_5103);
or U6687 (N_6687,N_5363,N_5562);
nand U6688 (N_6688,N_5809,N_5303);
nand U6689 (N_6689,N_5577,N_5620);
nand U6690 (N_6690,N_5882,N_5964);
nand U6691 (N_6691,N_5444,N_5387);
and U6692 (N_6692,N_5663,N_5788);
nor U6693 (N_6693,N_5815,N_5402);
or U6694 (N_6694,N_5625,N_5022);
nand U6695 (N_6695,N_5543,N_5117);
or U6696 (N_6696,N_5988,N_5941);
nand U6697 (N_6697,N_5048,N_5964);
nor U6698 (N_6698,N_5931,N_5388);
nor U6699 (N_6699,N_5596,N_5826);
nand U6700 (N_6700,N_5021,N_5159);
nand U6701 (N_6701,N_5391,N_5321);
and U6702 (N_6702,N_5671,N_5127);
nor U6703 (N_6703,N_5712,N_5378);
or U6704 (N_6704,N_5058,N_5004);
nand U6705 (N_6705,N_5890,N_5964);
nor U6706 (N_6706,N_5810,N_5257);
nand U6707 (N_6707,N_5154,N_5614);
or U6708 (N_6708,N_5924,N_5964);
and U6709 (N_6709,N_5317,N_5999);
or U6710 (N_6710,N_5357,N_5143);
xor U6711 (N_6711,N_5791,N_5822);
nand U6712 (N_6712,N_5168,N_5840);
or U6713 (N_6713,N_5523,N_5947);
and U6714 (N_6714,N_5472,N_5936);
nor U6715 (N_6715,N_5212,N_5572);
and U6716 (N_6716,N_5742,N_5691);
nand U6717 (N_6717,N_5056,N_5481);
and U6718 (N_6718,N_5627,N_5074);
or U6719 (N_6719,N_5051,N_5915);
or U6720 (N_6720,N_5985,N_5775);
nor U6721 (N_6721,N_5868,N_5421);
or U6722 (N_6722,N_5828,N_5766);
and U6723 (N_6723,N_5278,N_5331);
and U6724 (N_6724,N_5317,N_5177);
nand U6725 (N_6725,N_5491,N_5082);
and U6726 (N_6726,N_5400,N_5967);
and U6727 (N_6727,N_5469,N_5589);
nor U6728 (N_6728,N_5216,N_5207);
or U6729 (N_6729,N_5179,N_5833);
or U6730 (N_6730,N_5694,N_5000);
and U6731 (N_6731,N_5085,N_5533);
and U6732 (N_6732,N_5398,N_5122);
and U6733 (N_6733,N_5637,N_5785);
nand U6734 (N_6734,N_5540,N_5239);
nand U6735 (N_6735,N_5279,N_5108);
nor U6736 (N_6736,N_5559,N_5046);
nor U6737 (N_6737,N_5177,N_5034);
and U6738 (N_6738,N_5814,N_5761);
nand U6739 (N_6739,N_5107,N_5335);
or U6740 (N_6740,N_5956,N_5834);
nand U6741 (N_6741,N_5879,N_5307);
or U6742 (N_6742,N_5176,N_5146);
nand U6743 (N_6743,N_5896,N_5152);
nor U6744 (N_6744,N_5560,N_5124);
nand U6745 (N_6745,N_5309,N_5243);
nand U6746 (N_6746,N_5256,N_5370);
nor U6747 (N_6747,N_5886,N_5392);
nand U6748 (N_6748,N_5155,N_5358);
nor U6749 (N_6749,N_5220,N_5737);
and U6750 (N_6750,N_5365,N_5733);
nor U6751 (N_6751,N_5066,N_5799);
and U6752 (N_6752,N_5543,N_5425);
and U6753 (N_6753,N_5828,N_5005);
and U6754 (N_6754,N_5337,N_5616);
nand U6755 (N_6755,N_5870,N_5280);
xor U6756 (N_6756,N_5686,N_5347);
and U6757 (N_6757,N_5472,N_5830);
nor U6758 (N_6758,N_5835,N_5120);
nand U6759 (N_6759,N_5997,N_5711);
nand U6760 (N_6760,N_5092,N_5185);
nor U6761 (N_6761,N_5859,N_5027);
nand U6762 (N_6762,N_5477,N_5748);
nand U6763 (N_6763,N_5776,N_5856);
or U6764 (N_6764,N_5622,N_5316);
or U6765 (N_6765,N_5209,N_5728);
nand U6766 (N_6766,N_5617,N_5072);
or U6767 (N_6767,N_5652,N_5978);
nor U6768 (N_6768,N_5128,N_5982);
and U6769 (N_6769,N_5284,N_5154);
and U6770 (N_6770,N_5874,N_5212);
nor U6771 (N_6771,N_5550,N_5895);
nor U6772 (N_6772,N_5399,N_5604);
nor U6773 (N_6773,N_5183,N_5691);
nand U6774 (N_6774,N_5159,N_5924);
or U6775 (N_6775,N_5336,N_5479);
or U6776 (N_6776,N_5705,N_5548);
and U6777 (N_6777,N_5213,N_5736);
nand U6778 (N_6778,N_5836,N_5204);
or U6779 (N_6779,N_5871,N_5634);
nor U6780 (N_6780,N_5685,N_5030);
or U6781 (N_6781,N_5417,N_5309);
and U6782 (N_6782,N_5543,N_5953);
nand U6783 (N_6783,N_5507,N_5314);
and U6784 (N_6784,N_5425,N_5564);
and U6785 (N_6785,N_5618,N_5144);
nand U6786 (N_6786,N_5383,N_5118);
nand U6787 (N_6787,N_5627,N_5798);
nand U6788 (N_6788,N_5876,N_5892);
nor U6789 (N_6789,N_5046,N_5578);
nor U6790 (N_6790,N_5486,N_5365);
and U6791 (N_6791,N_5744,N_5085);
nor U6792 (N_6792,N_5578,N_5193);
xor U6793 (N_6793,N_5049,N_5460);
or U6794 (N_6794,N_5015,N_5295);
or U6795 (N_6795,N_5354,N_5525);
or U6796 (N_6796,N_5791,N_5340);
and U6797 (N_6797,N_5235,N_5907);
nor U6798 (N_6798,N_5338,N_5531);
nand U6799 (N_6799,N_5585,N_5188);
or U6800 (N_6800,N_5938,N_5531);
or U6801 (N_6801,N_5850,N_5692);
or U6802 (N_6802,N_5111,N_5172);
or U6803 (N_6803,N_5816,N_5533);
and U6804 (N_6804,N_5010,N_5143);
nor U6805 (N_6805,N_5793,N_5005);
nor U6806 (N_6806,N_5772,N_5932);
nor U6807 (N_6807,N_5220,N_5187);
nand U6808 (N_6808,N_5489,N_5880);
and U6809 (N_6809,N_5737,N_5767);
and U6810 (N_6810,N_5203,N_5512);
nor U6811 (N_6811,N_5532,N_5471);
and U6812 (N_6812,N_5119,N_5649);
or U6813 (N_6813,N_5607,N_5553);
and U6814 (N_6814,N_5903,N_5737);
nor U6815 (N_6815,N_5155,N_5037);
nor U6816 (N_6816,N_5650,N_5440);
nand U6817 (N_6817,N_5593,N_5065);
nor U6818 (N_6818,N_5993,N_5771);
and U6819 (N_6819,N_5521,N_5436);
nand U6820 (N_6820,N_5212,N_5872);
and U6821 (N_6821,N_5096,N_5952);
or U6822 (N_6822,N_5749,N_5799);
nor U6823 (N_6823,N_5221,N_5149);
and U6824 (N_6824,N_5762,N_5867);
nand U6825 (N_6825,N_5754,N_5380);
and U6826 (N_6826,N_5719,N_5155);
nor U6827 (N_6827,N_5954,N_5841);
and U6828 (N_6828,N_5400,N_5196);
nand U6829 (N_6829,N_5447,N_5357);
nor U6830 (N_6830,N_5251,N_5893);
or U6831 (N_6831,N_5383,N_5581);
and U6832 (N_6832,N_5351,N_5261);
nor U6833 (N_6833,N_5109,N_5026);
nor U6834 (N_6834,N_5353,N_5125);
or U6835 (N_6835,N_5076,N_5685);
nand U6836 (N_6836,N_5804,N_5037);
nor U6837 (N_6837,N_5780,N_5966);
or U6838 (N_6838,N_5049,N_5884);
nor U6839 (N_6839,N_5611,N_5861);
nor U6840 (N_6840,N_5441,N_5899);
xor U6841 (N_6841,N_5260,N_5509);
and U6842 (N_6842,N_5392,N_5148);
nor U6843 (N_6843,N_5364,N_5320);
nor U6844 (N_6844,N_5402,N_5495);
and U6845 (N_6845,N_5869,N_5272);
or U6846 (N_6846,N_5224,N_5210);
and U6847 (N_6847,N_5383,N_5830);
and U6848 (N_6848,N_5375,N_5940);
nand U6849 (N_6849,N_5722,N_5859);
and U6850 (N_6850,N_5547,N_5787);
or U6851 (N_6851,N_5538,N_5418);
and U6852 (N_6852,N_5708,N_5119);
or U6853 (N_6853,N_5459,N_5778);
nor U6854 (N_6854,N_5178,N_5749);
and U6855 (N_6855,N_5711,N_5334);
and U6856 (N_6856,N_5337,N_5388);
and U6857 (N_6857,N_5852,N_5650);
nor U6858 (N_6858,N_5958,N_5092);
or U6859 (N_6859,N_5344,N_5972);
nor U6860 (N_6860,N_5650,N_5101);
and U6861 (N_6861,N_5255,N_5575);
nand U6862 (N_6862,N_5490,N_5498);
and U6863 (N_6863,N_5771,N_5261);
or U6864 (N_6864,N_5114,N_5752);
nand U6865 (N_6865,N_5297,N_5609);
and U6866 (N_6866,N_5327,N_5682);
or U6867 (N_6867,N_5472,N_5046);
and U6868 (N_6868,N_5803,N_5734);
nand U6869 (N_6869,N_5118,N_5190);
or U6870 (N_6870,N_5352,N_5861);
and U6871 (N_6871,N_5000,N_5691);
nor U6872 (N_6872,N_5727,N_5366);
nand U6873 (N_6873,N_5841,N_5769);
or U6874 (N_6874,N_5863,N_5968);
nand U6875 (N_6875,N_5405,N_5046);
or U6876 (N_6876,N_5341,N_5326);
or U6877 (N_6877,N_5122,N_5415);
nor U6878 (N_6878,N_5910,N_5599);
and U6879 (N_6879,N_5943,N_5312);
nand U6880 (N_6880,N_5806,N_5655);
nor U6881 (N_6881,N_5958,N_5957);
or U6882 (N_6882,N_5873,N_5411);
nor U6883 (N_6883,N_5816,N_5030);
nor U6884 (N_6884,N_5027,N_5036);
nor U6885 (N_6885,N_5013,N_5449);
or U6886 (N_6886,N_5610,N_5701);
nand U6887 (N_6887,N_5251,N_5896);
and U6888 (N_6888,N_5962,N_5507);
xor U6889 (N_6889,N_5022,N_5587);
nand U6890 (N_6890,N_5685,N_5815);
and U6891 (N_6891,N_5233,N_5150);
xor U6892 (N_6892,N_5580,N_5284);
nand U6893 (N_6893,N_5402,N_5519);
and U6894 (N_6894,N_5647,N_5642);
and U6895 (N_6895,N_5923,N_5321);
nor U6896 (N_6896,N_5317,N_5226);
and U6897 (N_6897,N_5365,N_5103);
nor U6898 (N_6898,N_5295,N_5860);
nand U6899 (N_6899,N_5611,N_5046);
nand U6900 (N_6900,N_5745,N_5184);
or U6901 (N_6901,N_5531,N_5981);
or U6902 (N_6902,N_5194,N_5521);
or U6903 (N_6903,N_5913,N_5843);
nor U6904 (N_6904,N_5231,N_5263);
xor U6905 (N_6905,N_5635,N_5521);
nand U6906 (N_6906,N_5174,N_5759);
or U6907 (N_6907,N_5505,N_5873);
or U6908 (N_6908,N_5722,N_5363);
nor U6909 (N_6909,N_5380,N_5094);
nor U6910 (N_6910,N_5321,N_5993);
nor U6911 (N_6911,N_5362,N_5178);
and U6912 (N_6912,N_5389,N_5335);
nand U6913 (N_6913,N_5132,N_5814);
and U6914 (N_6914,N_5803,N_5166);
nand U6915 (N_6915,N_5537,N_5126);
nand U6916 (N_6916,N_5274,N_5275);
or U6917 (N_6917,N_5666,N_5271);
nor U6918 (N_6918,N_5306,N_5933);
nand U6919 (N_6919,N_5091,N_5209);
nor U6920 (N_6920,N_5468,N_5401);
nand U6921 (N_6921,N_5606,N_5955);
and U6922 (N_6922,N_5663,N_5391);
nand U6923 (N_6923,N_5017,N_5601);
and U6924 (N_6924,N_5994,N_5135);
nor U6925 (N_6925,N_5378,N_5862);
nor U6926 (N_6926,N_5124,N_5624);
and U6927 (N_6927,N_5523,N_5643);
nand U6928 (N_6928,N_5250,N_5784);
nand U6929 (N_6929,N_5693,N_5812);
nor U6930 (N_6930,N_5255,N_5534);
nand U6931 (N_6931,N_5694,N_5397);
or U6932 (N_6932,N_5390,N_5402);
and U6933 (N_6933,N_5133,N_5648);
nor U6934 (N_6934,N_5206,N_5741);
nand U6935 (N_6935,N_5198,N_5412);
nand U6936 (N_6936,N_5046,N_5441);
nand U6937 (N_6937,N_5740,N_5879);
or U6938 (N_6938,N_5516,N_5677);
or U6939 (N_6939,N_5520,N_5162);
or U6940 (N_6940,N_5060,N_5257);
and U6941 (N_6941,N_5942,N_5540);
and U6942 (N_6942,N_5397,N_5773);
or U6943 (N_6943,N_5228,N_5003);
nor U6944 (N_6944,N_5249,N_5537);
nor U6945 (N_6945,N_5948,N_5333);
nor U6946 (N_6946,N_5798,N_5556);
and U6947 (N_6947,N_5940,N_5699);
and U6948 (N_6948,N_5187,N_5448);
nand U6949 (N_6949,N_5614,N_5422);
and U6950 (N_6950,N_5404,N_5014);
nand U6951 (N_6951,N_5058,N_5769);
or U6952 (N_6952,N_5521,N_5267);
or U6953 (N_6953,N_5545,N_5713);
nor U6954 (N_6954,N_5361,N_5172);
or U6955 (N_6955,N_5284,N_5255);
nor U6956 (N_6956,N_5897,N_5419);
or U6957 (N_6957,N_5245,N_5487);
or U6958 (N_6958,N_5761,N_5568);
or U6959 (N_6959,N_5510,N_5837);
nand U6960 (N_6960,N_5854,N_5222);
and U6961 (N_6961,N_5949,N_5176);
or U6962 (N_6962,N_5830,N_5279);
and U6963 (N_6963,N_5075,N_5892);
nand U6964 (N_6964,N_5804,N_5841);
and U6965 (N_6965,N_5560,N_5721);
nor U6966 (N_6966,N_5508,N_5434);
or U6967 (N_6967,N_5700,N_5142);
nor U6968 (N_6968,N_5957,N_5385);
or U6969 (N_6969,N_5256,N_5139);
or U6970 (N_6970,N_5498,N_5272);
nor U6971 (N_6971,N_5077,N_5460);
or U6972 (N_6972,N_5489,N_5859);
and U6973 (N_6973,N_5606,N_5646);
or U6974 (N_6974,N_5641,N_5416);
or U6975 (N_6975,N_5951,N_5950);
nor U6976 (N_6976,N_5643,N_5685);
and U6977 (N_6977,N_5760,N_5049);
nand U6978 (N_6978,N_5446,N_5724);
or U6979 (N_6979,N_5776,N_5705);
or U6980 (N_6980,N_5098,N_5577);
or U6981 (N_6981,N_5683,N_5531);
and U6982 (N_6982,N_5431,N_5584);
nor U6983 (N_6983,N_5747,N_5169);
nand U6984 (N_6984,N_5194,N_5453);
nor U6985 (N_6985,N_5825,N_5494);
nor U6986 (N_6986,N_5757,N_5001);
nand U6987 (N_6987,N_5436,N_5838);
nor U6988 (N_6988,N_5983,N_5347);
nor U6989 (N_6989,N_5189,N_5038);
or U6990 (N_6990,N_5851,N_5304);
or U6991 (N_6991,N_5847,N_5661);
nand U6992 (N_6992,N_5195,N_5752);
or U6993 (N_6993,N_5001,N_5879);
nor U6994 (N_6994,N_5980,N_5043);
nor U6995 (N_6995,N_5083,N_5254);
and U6996 (N_6996,N_5582,N_5155);
nor U6997 (N_6997,N_5990,N_5208);
nand U6998 (N_6998,N_5500,N_5632);
or U6999 (N_6999,N_5860,N_5948);
nor U7000 (N_7000,N_6571,N_6330);
or U7001 (N_7001,N_6155,N_6914);
or U7002 (N_7002,N_6227,N_6030);
nand U7003 (N_7003,N_6469,N_6923);
or U7004 (N_7004,N_6134,N_6592);
nor U7005 (N_7005,N_6891,N_6577);
and U7006 (N_7006,N_6312,N_6302);
and U7007 (N_7007,N_6282,N_6277);
nand U7008 (N_7008,N_6096,N_6388);
and U7009 (N_7009,N_6257,N_6678);
or U7010 (N_7010,N_6797,N_6912);
or U7011 (N_7011,N_6174,N_6296);
and U7012 (N_7012,N_6769,N_6660);
nor U7013 (N_7013,N_6074,N_6793);
or U7014 (N_7014,N_6634,N_6029);
and U7015 (N_7015,N_6798,N_6364);
nor U7016 (N_7016,N_6421,N_6256);
or U7017 (N_7017,N_6832,N_6360);
or U7018 (N_7018,N_6412,N_6309);
and U7019 (N_7019,N_6645,N_6075);
or U7020 (N_7020,N_6380,N_6056);
nand U7021 (N_7021,N_6119,N_6274);
nor U7022 (N_7022,N_6345,N_6117);
nor U7023 (N_7023,N_6325,N_6034);
and U7024 (N_7024,N_6992,N_6584);
and U7025 (N_7025,N_6605,N_6014);
nand U7026 (N_7026,N_6445,N_6062);
or U7027 (N_7027,N_6899,N_6591);
or U7028 (N_7028,N_6852,N_6949);
or U7029 (N_7029,N_6858,N_6960);
nor U7030 (N_7030,N_6252,N_6067);
or U7031 (N_7031,N_6479,N_6483);
or U7032 (N_7032,N_6422,N_6272);
nor U7033 (N_7033,N_6481,N_6893);
nor U7034 (N_7034,N_6970,N_6642);
and U7035 (N_7035,N_6694,N_6083);
nor U7036 (N_7036,N_6962,N_6619);
or U7037 (N_7037,N_6974,N_6526);
and U7038 (N_7038,N_6452,N_6488);
and U7039 (N_7039,N_6513,N_6885);
or U7040 (N_7040,N_6219,N_6443);
and U7041 (N_7041,N_6465,N_6983);
and U7042 (N_7042,N_6040,N_6509);
nor U7043 (N_7043,N_6763,N_6341);
nor U7044 (N_7044,N_6868,N_6944);
and U7045 (N_7045,N_6870,N_6672);
and U7046 (N_7046,N_6831,N_6265);
nor U7047 (N_7047,N_6299,N_6281);
nand U7048 (N_7048,N_6808,N_6218);
xnor U7049 (N_7049,N_6984,N_6264);
nor U7050 (N_7050,N_6175,N_6095);
nor U7051 (N_7051,N_6298,N_6140);
nor U7052 (N_7052,N_6856,N_6215);
and U7053 (N_7053,N_6574,N_6021);
or U7054 (N_7054,N_6965,N_6730);
or U7055 (N_7055,N_6186,N_6639);
nor U7056 (N_7056,N_6123,N_6196);
or U7057 (N_7057,N_6743,N_6118);
or U7058 (N_7058,N_6401,N_6582);
nor U7059 (N_7059,N_6512,N_6379);
nand U7060 (N_7060,N_6587,N_6644);
nor U7061 (N_7061,N_6036,N_6776);
nor U7062 (N_7062,N_6935,N_6648);
or U7063 (N_7063,N_6113,N_6154);
and U7064 (N_7064,N_6597,N_6342);
or U7065 (N_7065,N_6843,N_6514);
or U7066 (N_7066,N_6403,N_6551);
or U7067 (N_7067,N_6669,N_6573);
nor U7068 (N_7068,N_6127,N_6522);
nor U7069 (N_7069,N_6092,N_6413);
or U7070 (N_7070,N_6623,N_6718);
or U7071 (N_7071,N_6037,N_6842);
nand U7072 (N_7072,N_6815,N_6789);
nand U7073 (N_7073,N_6911,N_6076);
or U7074 (N_7074,N_6745,N_6951);
or U7075 (N_7075,N_6316,N_6724);
nand U7076 (N_7076,N_6505,N_6959);
or U7077 (N_7077,N_6437,N_6916);
nand U7078 (N_7078,N_6759,N_6781);
nor U7079 (N_7079,N_6225,N_6658);
nand U7080 (N_7080,N_6816,N_6071);
and U7081 (N_7081,N_6840,N_6384);
nor U7082 (N_7082,N_6354,N_6957);
or U7083 (N_7083,N_6011,N_6996);
and U7084 (N_7084,N_6482,N_6480);
or U7085 (N_7085,N_6601,N_6251);
nand U7086 (N_7086,N_6953,N_6129);
nor U7087 (N_7087,N_6667,N_6449);
or U7088 (N_7088,N_6552,N_6841);
nor U7089 (N_7089,N_6518,N_6824);
and U7090 (N_7090,N_6979,N_6833);
nand U7091 (N_7091,N_6487,N_6566);
nor U7092 (N_7092,N_6968,N_6359);
nand U7093 (N_7093,N_6908,N_6019);
and U7094 (N_7094,N_6429,N_6801);
and U7095 (N_7095,N_6244,N_6922);
and U7096 (N_7096,N_6693,N_6652);
and U7097 (N_7097,N_6041,N_6976);
nor U7098 (N_7098,N_6270,N_6268);
or U7099 (N_7099,N_6416,N_6398);
and U7100 (N_7100,N_6839,N_6973);
or U7101 (N_7101,N_6098,N_6042);
nor U7102 (N_7102,N_6451,N_6865);
and U7103 (N_7103,N_6077,N_6150);
or U7104 (N_7104,N_6521,N_6002);
nor U7105 (N_7105,N_6246,N_6611);
nor U7106 (N_7106,N_6440,N_6685);
nand U7107 (N_7107,N_6564,N_6696);
or U7108 (N_7108,N_6989,N_6245);
or U7109 (N_7109,N_6527,N_6160);
or U7110 (N_7110,N_6131,N_6448);
and U7111 (N_7111,N_6598,N_6016);
nand U7112 (N_7112,N_6236,N_6144);
nor U7113 (N_7113,N_6603,N_6431);
nor U7114 (N_7114,N_6604,N_6169);
nor U7115 (N_7115,N_6762,N_6723);
and U7116 (N_7116,N_6321,N_6085);
and U7117 (N_7117,N_6570,N_6136);
nand U7118 (N_7118,N_6947,N_6758);
and U7119 (N_7119,N_6837,N_6927);
nor U7120 (N_7120,N_6269,N_6609);
nand U7121 (N_7121,N_6541,N_6322);
nor U7122 (N_7122,N_6365,N_6751);
nand U7123 (N_7123,N_6662,N_6569);
nand U7124 (N_7124,N_6862,N_6241);
and U7125 (N_7125,N_6222,N_6708);
and U7126 (N_7126,N_6640,N_6934);
nand U7127 (N_7127,N_6361,N_6247);
nand U7128 (N_7128,N_6814,N_6060);
nor U7129 (N_7129,N_6271,N_6905);
or U7130 (N_7130,N_6059,N_6727);
nand U7131 (N_7131,N_6779,N_6120);
nand U7132 (N_7132,N_6687,N_6647);
nand U7133 (N_7133,N_6627,N_6790);
nand U7134 (N_7134,N_6020,N_6133);
nand U7135 (N_7135,N_6803,N_6765);
or U7136 (N_7136,N_6884,N_6677);
and U7137 (N_7137,N_6917,N_6494);
and U7138 (N_7138,N_6848,N_6371);
nand U7139 (N_7139,N_6819,N_6520);
or U7140 (N_7140,N_6007,N_6346);
nand U7141 (N_7141,N_6100,N_6877);
and U7142 (N_7142,N_6532,N_6612);
and U7143 (N_7143,N_6396,N_6475);
nand U7144 (N_7144,N_6213,N_6210);
nor U7145 (N_7145,N_6882,N_6430);
or U7146 (N_7146,N_6702,N_6954);
xor U7147 (N_7147,N_6317,N_6048);
and U7148 (N_7148,N_6046,N_6990);
nor U7149 (N_7149,N_6279,N_6802);
nor U7150 (N_7150,N_6108,N_6641);
nand U7151 (N_7151,N_6539,N_6772);
and U7152 (N_7152,N_6871,N_6284);
and U7153 (N_7153,N_6999,N_6301);
nand U7154 (N_7154,N_6378,N_6557);
and U7155 (N_7155,N_6939,N_6435);
nand U7156 (N_7156,N_6050,N_6446);
or U7157 (N_7157,N_6664,N_6796);
nor U7158 (N_7158,N_6065,N_6909);
nor U7159 (N_7159,N_6516,N_6988);
or U7160 (N_7160,N_6757,N_6242);
nor U7161 (N_7161,N_6670,N_6495);
and U7162 (N_7162,N_6419,N_6635);
or U7163 (N_7163,N_6053,N_6580);
or U7164 (N_7164,N_6504,N_6528);
and U7165 (N_7165,N_6358,N_6233);
nor U7166 (N_7166,N_6190,N_6069);
nand U7167 (N_7167,N_6397,N_6561);
and U7168 (N_7168,N_6375,N_6286);
or U7169 (N_7169,N_6332,N_6485);
xor U7170 (N_7170,N_6918,N_6187);
or U7171 (N_7171,N_6283,N_6054);
nor U7172 (N_7172,N_6148,N_6051);
nor U7173 (N_7173,N_6982,N_6945);
or U7174 (N_7174,N_6964,N_6139);
and U7175 (N_7175,N_6825,N_6567);
and U7176 (N_7176,N_6699,N_6867);
nand U7177 (N_7177,N_6239,N_6903);
nand U7178 (N_7178,N_6300,N_6936);
nand U7179 (N_7179,N_6207,N_6863);
nor U7180 (N_7180,N_6890,N_6544);
and U7181 (N_7181,N_6860,N_6220);
nand U7182 (N_7182,N_6695,N_6826);
nand U7183 (N_7183,N_6761,N_6315);
or U7184 (N_7184,N_6807,N_6637);
or U7185 (N_7185,N_6084,N_6439);
nand U7186 (N_7186,N_6478,N_6904);
or U7187 (N_7187,N_6058,N_6854);
or U7188 (N_7188,N_6313,N_6173);
nand U7189 (N_7189,N_6700,N_6209);
nor U7190 (N_7190,N_6369,N_6583);
or U7191 (N_7191,N_6333,N_6367);
nor U7192 (N_7192,N_6955,N_6472);
nor U7193 (N_7193,N_6921,N_6529);
nor U7194 (N_7194,N_6698,N_6755);
nand U7195 (N_7195,N_6156,N_6292);
nor U7196 (N_7196,N_6460,N_6686);
nand U7197 (N_7197,N_6515,N_6436);
nand U7198 (N_7198,N_6203,N_6079);
nand U7199 (N_7199,N_6829,N_6794);
nor U7200 (N_7200,N_6946,N_6651);
nor U7201 (N_7201,N_6656,N_6303);
or U7202 (N_7202,N_6255,N_6760);
nor U7203 (N_7203,N_6188,N_6864);
and U7204 (N_7204,N_6602,N_6559);
and U7205 (N_7205,N_6705,N_6082);
nand U7206 (N_7206,N_6850,N_6625);
and U7207 (N_7207,N_6978,N_6971);
or U7208 (N_7208,N_6287,N_6106);
nand U7209 (N_7209,N_6896,N_6237);
or U7210 (N_7210,N_6942,N_6463);
nor U7211 (N_7211,N_6734,N_6809);
nand U7212 (N_7212,N_6356,N_6746);
or U7213 (N_7213,N_6261,N_6943);
nor U7214 (N_7214,N_6950,N_6250);
nand U7215 (N_7215,N_6128,N_6327);
nor U7216 (N_7216,N_6170,N_6399);
nor U7217 (N_7217,N_6417,N_6434);
nor U7218 (N_7218,N_6748,N_6726);
nor U7219 (N_7219,N_6097,N_6613);
nand U7220 (N_7220,N_6895,N_6786);
nor U7221 (N_7221,N_6307,N_6035);
nand U7222 (N_7222,N_6558,N_6044);
or U7223 (N_7223,N_6105,N_6400);
and U7224 (N_7224,N_6766,N_6919);
or U7225 (N_7225,N_6110,N_6116);
and U7226 (N_7226,N_6510,N_6859);
nand U7227 (N_7227,N_6366,N_6590);
nand U7228 (N_7228,N_6608,N_6381);
nand U7229 (N_7229,N_6783,N_6107);
and U7230 (N_7230,N_6663,N_6703);
and U7231 (N_7231,N_6370,N_6392);
nand U7232 (N_7232,N_6579,N_6178);
and U7233 (N_7233,N_6800,N_6249);
and U7234 (N_7234,N_6047,N_6986);
or U7235 (N_7235,N_6376,N_6151);
nand U7236 (N_7236,N_6471,N_6818);
and U7237 (N_7237,N_6238,N_6888);
and U7238 (N_7238,N_6735,N_6719);
nor U7239 (N_7239,N_6661,N_6621);
or U7240 (N_7240,N_6428,N_6620);
and U7241 (N_7241,N_6349,N_6638);
nand U7242 (N_7242,N_6081,N_6103);
and U7243 (N_7243,N_6070,N_6486);
nor U7244 (N_7244,N_6273,N_6545);
or U7245 (N_7245,N_6424,N_6458);
nor U7246 (N_7246,N_6866,N_6183);
or U7247 (N_7247,N_6254,N_6711);
and U7248 (N_7248,N_6997,N_6845);
nor U7249 (N_7249,N_6624,N_6088);
and U7250 (N_7250,N_6288,N_6229);
and U7251 (N_7251,N_6683,N_6519);
nand U7252 (N_7252,N_6828,N_6650);
nor U7253 (N_7253,N_6453,N_6985);
xnor U7254 (N_7254,N_6336,N_6750);
nand U7255 (N_7255,N_6524,N_6501);
or U7256 (N_7256,N_6872,N_6130);
nor U7257 (N_7257,N_6844,N_6147);
nand U7258 (N_7258,N_6122,N_6967);
and U7259 (N_7259,N_6740,N_6290);
nand U7260 (N_7260,N_6963,N_6351);
nor U7261 (N_7261,N_6023,N_6474);
and U7262 (N_7262,N_6142,N_6172);
nand U7263 (N_7263,N_6061,N_6956);
xor U7264 (N_7264,N_6291,N_6163);
nor U7265 (N_7265,N_6900,N_6659);
and U7266 (N_7266,N_6715,N_6224);
nand U7267 (N_7267,N_6792,N_6243);
nand U7268 (N_7268,N_6933,N_6024);
or U7269 (N_7269,N_6576,N_6338);
nor U7270 (N_7270,N_6555,N_6861);
nor U7271 (N_7271,N_6668,N_6937);
and U7272 (N_7272,N_6714,N_6994);
nor U7273 (N_7273,N_6427,N_6733);
and U7274 (N_7274,N_6414,N_6348);
nand U7275 (N_7275,N_6262,N_6771);
and U7276 (N_7276,N_6208,N_6595);
nor U7277 (N_7277,N_6340,N_6200);
nor U7278 (N_7278,N_6628,N_6805);
nor U7279 (N_7279,N_6198,N_6138);
nand U7280 (N_7280,N_6770,N_6892);
and U7281 (N_7281,N_6467,N_6217);
nor U7282 (N_7282,N_6897,N_6390);
and U7283 (N_7283,N_6876,N_6423);
nand U7284 (N_7284,N_6902,N_6906);
nand U7285 (N_7285,N_6682,N_6033);
nand U7286 (N_7286,N_6588,N_6143);
nor U7287 (N_7287,N_6560,N_6407);
nand U7288 (N_7288,N_6673,N_6847);
or U7289 (N_7289,N_6226,N_6523);
xor U7290 (N_7290,N_6199,N_6630);
or U7291 (N_7291,N_6649,N_6838);
and U7292 (N_7292,N_6055,N_6491);
and U7293 (N_7293,N_6806,N_6631);
nor U7294 (N_7294,N_6846,N_6575);
nor U7295 (N_7295,N_6910,N_6738);
or U7296 (N_7296,N_6032,N_6260);
and U7297 (N_7297,N_6402,N_6812);
nand U7298 (N_7298,N_6804,N_6450);
nor U7299 (N_7299,N_6464,N_6907);
nand U7300 (N_7300,N_6420,N_6438);
or U7301 (N_7301,N_6126,N_6318);
and U7302 (N_7302,N_6995,N_6537);
and U7303 (N_7303,N_6599,N_6409);
nor U7304 (N_7304,N_6607,N_6194);
nor U7305 (N_7305,N_6655,N_6159);
nand U7306 (N_7306,N_6774,N_6610);
nor U7307 (N_7307,N_6689,N_6498);
nor U7308 (N_7308,N_6493,N_6830);
or U7309 (N_7309,N_6869,N_6554);
nand U7310 (N_7310,N_6005,N_6881);
nand U7311 (N_7311,N_6404,N_6386);
nor U7312 (N_7312,N_6679,N_6878);
nand U7313 (N_7313,N_6164,N_6606);
or U7314 (N_7314,N_6001,N_6228);
nand U7315 (N_7315,N_6991,N_6089);
and U7316 (N_7316,N_6006,N_6572);
and U7317 (N_7317,N_6185,N_6177);
and U7318 (N_7318,N_6295,N_6731);
nor U7319 (N_7319,N_6328,N_6114);
xnor U7320 (N_7320,N_6232,N_6728);
nor U7321 (N_7321,N_6004,N_6530);
nor U7322 (N_7322,N_6276,N_6924);
nand U7323 (N_7323,N_6353,N_6820);
nor U7324 (N_7324,N_6179,N_6152);
nand U7325 (N_7325,N_6433,N_6168);
nor U7326 (N_7326,N_6556,N_6344);
nand U7327 (N_7327,N_6548,N_6101);
nor U7328 (N_7328,N_6094,N_6879);
and U7329 (N_7329,N_6952,N_6025);
and U7330 (N_7330,N_6767,N_6461);
nor U7331 (N_7331,N_6387,N_6615);
nand U7332 (N_7332,N_6240,N_6444);
and U7333 (N_7333,N_6454,N_6003);
or U7334 (N_7334,N_6618,N_6216);
or U7335 (N_7335,N_6886,N_6742);
nor U7336 (N_7336,N_6235,N_6182);
nand U7337 (N_7337,N_6553,N_6263);
or U7338 (N_7338,N_6915,N_6857);
nand U7339 (N_7339,N_6500,N_6442);
and U7340 (N_7340,N_6459,N_6851);
nor U7341 (N_7341,N_6517,N_6093);
or U7342 (N_7342,N_6626,N_6115);
nand U7343 (N_7343,N_6080,N_6455);
and U7344 (N_7344,N_6331,N_6940);
nor U7345 (N_7345,N_6739,N_6674);
nor U7346 (N_7346,N_6535,N_6355);
nor U7347 (N_7347,N_6109,N_6646);
and U7348 (N_7348,N_6280,N_6204);
nand U7349 (N_7349,N_6785,N_6010);
nand U7350 (N_7350,N_6121,N_6880);
and U7351 (N_7351,N_6665,N_6675);
nor U7352 (N_7352,N_6202,N_6206);
and U7353 (N_7353,N_6536,N_6395);
nor U7354 (N_7354,N_6230,N_6657);
nor U7355 (N_7355,N_6310,N_6720);
nor U7356 (N_7356,N_6275,N_6320);
nor U7357 (N_7357,N_6343,N_6594);
or U7358 (N_7358,N_6267,N_6432);
nor U7359 (N_7359,N_6339,N_6617);
nor U7360 (N_7360,N_6810,N_6408);
and U7361 (N_7361,N_6931,N_6932);
nand U7362 (N_7362,N_6546,N_6784);
nor U7363 (N_7363,N_6031,N_6543);
or U7364 (N_7364,N_6362,N_6191);
and U7365 (N_7365,N_6181,N_6072);
nand U7366 (N_7366,N_6319,N_6889);
nand U7367 (N_7367,N_6335,N_6063);
or U7368 (N_7368,N_6057,N_6141);
nor U7369 (N_7369,N_6064,N_6490);
and U7370 (N_7370,N_6166,N_6104);
nor U7371 (N_7371,N_6920,N_6925);
nor U7372 (N_7372,N_6966,N_6167);
nor U7373 (N_7373,N_6780,N_6489);
and U7374 (N_7374,N_6052,N_6087);
and U7375 (N_7375,N_6135,N_6171);
nand U7376 (N_7376,N_6531,N_6898);
nor U7377 (N_7377,N_6393,N_6690);
nor U7378 (N_7378,N_6773,N_6015);
nand U7379 (N_7379,N_6600,N_6542);
nand U7380 (N_7380,N_6722,N_6124);
and U7381 (N_7381,N_6323,N_6180);
nand U7382 (N_7382,N_6749,N_6248);
or U7383 (N_7383,N_6294,N_6680);
or U7384 (N_7384,N_6221,N_6855);
nand U7385 (N_7385,N_6534,N_6496);
and U7386 (N_7386,N_6913,N_6707);
nand U7387 (N_7387,N_6314,N_6347);
nand U7388 (N_7388,N_6737,N_6716);
nor U7389 (N_7389,N_6525,N_6149);
nor U7390 (N_7390,N_6499,N_6091);
or U7391 (N_7391,N_6578,N_6508);
nor U7392 (N_7392,N_6132,N_6350);
and U7393 (N_7393,N_6297,N_6258);
or U7394 (N_7394,N_6980,N_6972);
or U7395 (N_7395,N_6017,N_6285);
or U7396 (N_7396,N_6326,N_6157);
and U7397 (N_7397,N_6470,N_6629);
or U7398 (N_7398,N_6028,N_6456);
nand U7399 (N_7399,N_6813,N_6926);
and U7400 (N_7400,N_6732,N_6993);
or U7401 (N_7401,N_6468,N_6756);
and U7402 (N_7402,N_6506,N_6883);
and U7403 (N_7403,N_6836,N_6622);
nor U7404 (N_7404,N_6441,N_6176);
nand U7405 (N_7405,N_6636,N_6589);
and U7406 (N_7406,N_6125,N_6259);
and U7407 (N_7407,N_6616,N_6352);
nor U7408 (N_7408,N_6073,N_6305);
nand U7409 (N_7409,N_6596,N_6411);
and U7410 (N_7410,N_6391,N_6383);
and U7411 (N_7411,N_6975,N_6568);
and U7412 (N_7412,N_6713,N_6747);
and U7413 (N_7413,N_6214,N_6811);
nand U7414 (N_7414,N_6009,N_6234);
nand U7415 (N_7415,N_6266,N_6278);
or U7416 (N_7416,N_6145,N_6562);
or U7417 (N_7417,N_6357,N_6835);
or U7418 (N_7418,N_6410,N_6692);
or U7419 (N_7419,N_6507,N_6146);
nand U7420 (N_7420,N_6654,N_6068);
and U7421 (N_7421,N_6195,N_6363);
xor U7422 (N_7422,N_6764,N_6928);
or U7423 (N_7423,N_6827,N_6744);
or U7424 (N_7424,N_6008,N_6503);
and U7425 (N_7425,N_6643,N_6415);
and U7426 (N_7426,N_6875,N_6045);
or U7427 (N_7427,N_6334,N_6153);
nand U7428 (N_7428,N_6165,N_6477);
and U7429 (N_7429,N_6688,N_6538);
or U7430 (N_7430,N_6676,N_6775);
and U7431 (N_7431,N_6729,N_6308);
or U7432 (N_7432,N_6373,N_6377);
and U7433 (N_7433,N_6043,N_6701);
and U7434 (N_7434,N_6102,N_6511);
or U7435 (N_7435,N_6706,N_6549);
nor U7436 (N_7436,N_6653,N_6026);
and U7437 (N_7437,N_6887,N_6853);
nand U7438 (N_7438,N_6681,N_6473);
and U7439 (N_7439,N_6337,N_6184);
and U7440 (N_7440,N_6709,N_6018);
and U7441 (N_7441,N_6788,N_6476);
nand U7442 (N_7442,N_6484,N_6581);
nor U7443 (N_7443,N_6752,N_6158);
nor U7444 (N_7444,N_6012,N_6930);
and U7445 (N_7445,N_6768,N_6585);
and U7446 (N_7446,N_6374,N_6563);
and U7447 (N_7447,N_6704,N_6078);
nand U7448 (N_7448,N_6712,N_6389);
and U7449 (N_7449,N_6632,N_6961);
or U7450 (N_7450,N_6193,N_6137);
or U7451 (N_7451,N_6721,N_6736);
nand U7452 (N_7452,N_6741,N_6874);
or U7453 (N_7453,N_6684,N_6394);
nand U7454 (N_7454,N_6717,N_6948);
and U7455 (N_7455,N_6197,N_6192);
and U7456 (N_7456,N_6791,N_6754);
and U7457 (N_7457,N_6998,N_6372);
nand U7458 (N_7458,N_6823,N_6466);
nand U7459 (N_7459,N_6586,N_6565);
nor U7460 (N_7460,N_6969,N_6189);
or U7461 (N_7461,N_6834,N_6253);
nor U7462 (N_7462,N_6666,N_6112);
nand U7463 (N_7463,N_6049,N_6426);
and U7464 (N_7464,N_6671,N_6593);
nand U7465 (N_7465,N_6013,N_6457);
or U7466 (N_7466,N_6614,N_6231);
or U7467 (N_7467,N_6550,N_6938);
nor U7468 (N_7468,N_6894,N_6368);
or U7469 (N_7469,N_6697,N_6405);
or U7470 (N_7470,N_6385,N_6795);
and U7471 (N_7471,N_6691,N_6633);
nor U7472 (N_7472,N_6090,N_6211);
and U7473 (N_7473,N_6425,N_6289);
nand U7474 (N_7474,N_6782,N_6497);
or U7475 (N_7475,N_6540,N_6161);
nand U7476 (N_7476,N_6205,N_6849);
nor U7477 (N_7477,N_6223,N_6901);
nor U7478 (N_7478,N_6039,N_6778);
nor U7479 (N_7479,N_6941,N_6753);
or U7480 (N_7480,N_6311,N_6304);
nor U7481 (N_7481,N_6492,N_6710);
or U7482 (N_7482,N_6777,N_6418);
nand U7483 (N_7483,N_6000,N_6817);
or U7484 (N_7484,N_6533,N_6873);
nand U7485 (N_7485,N_6201,N_6027);
and U7486 (N_7486,N_6382,N_6038);
nand U7487 (N_7487,N_6725,N_6406);
and U7488 (N_7488,N_6502,N_6958);
nor U7489 (N_7489,N_6977,N_6162);
or U7490 (N_7490,N_6822,N_6324);
and U7491 (N_7491,N_6447,N_6022);
or U7492 (N_7492,N_6066,N_6821);
nand U7493 (N_7493,N_6086,N_6987);
nor U7494 (N_7494,N_6099,N_6799);
and U7495 (N_7495,N_6547,N_6462);
nor U7496 (N_7496,N_6981,N_6787);
and U7497 (N_7497,N_6929,N_6306);
or U7498 (N_7498,N_6329,N_6111);
and U7499 (N_7499,N_6293,N_6212);
or U7500 (N_7500,N_6511,N_6085);
or U7501 (N_7501,N_6972,N_6403);
nor U7502 (N_7502,N_6283,N_6838);
or U7503 (N_7503,N_6824,N_6867);
nand U7504 (N_7504,N_6600,N_6383);
or U7505 (N_7505,N_6034,N_6717);
and U7506 (N_7506,N_6537,N_6444);
nor U7507 (N_7507,N_6141,N_6654);
and U7508 (N_7508,N_6443,N_6240);
nand U7509 (N_7509,N_6543,N_6388);
nand U7510 (N_7510,N_6130,N_6734);
and U7511 (N_7511,N_6636,N_6296);
or U7512 (N_7512,N_6575,N_6912);
or U7513 (N_7513,N_6092,N_6160);
xor U7514 (N_7514,N_6381,N_6213);
nor U7515 (N_7515,N_6178,N_6249);
nor U7516 (N_7516,N_6813,N_6775);
nor U7517 (N_7517,N_6305,N_6493);
and U7518 (N_7518,N_6637,N_6065);
nor U7519 (N_7519,N_6861,N_6830);
nand U7520 (N_7520,N_6842,N_6144);
and U7521 (N_7521,N_6236,N_6677);
nand U7522 (N_7522,N_6509,N_6638);
or U7523 (N_7523,N_6934,N_6271);
nand U7524 (N_7524,N_6458,N_6621);
nand U7525 (N_7525,N_6647,N_6426);
and U7526 (N_7526,N_6318,N_6887);
or U7527 (N_7527,N_6357,N_6472);
or U7528 (N_7528,N_6318,N_6615);
or U7529 (N_7529,N_6613,N_6642);
nand U7530 (N_7530,N_6878,N_6770);
or U7531 (N_7531,N_6878,N_6647);
nor U7532 (N_7532,N_6404,N_6984);
nor U7533 (N_7533,N_6499,N_6007);
or U7534 (N_7534,N_6989,N_6396);
nor U7535 (N_7535,N_6756,N_6479);
nand U7536 (N_7536,N_6603,N_6259);
nand U7537 (N_7537,N_6821,N_6357);
nand U7538 (N_7538,N_6510,N_6115);
nand U7539 (N_7539,N_6192,N_6054);
nand U7540 (N_7540,N_6978,N_6962);
nand U7541 (N_7541,N_6086,N_6123);
and U7542 (N_7542,N_6507,N_6171);
nand U7543 (N_7543,N_6925,N_6661);
nand U7544 (N_7544,N_6303,N_6975);
nor U7545 (N_7545,N_6455,N_6148);
or U7546 (N_7546,N_6485,N_6499);
xnor U7547 (N_7547,N_6377,N_6706);
nand U7548 (N_7548,N_6621,N_6037);
nor U7549 (N_7549,N_6508,N_6217);
nor U7550 (N_7550,N_6862,N_6356);
or U7551 (N_7551,N_6082,N_6501);
and U7552 (N_7552,N_6853,N_6038);
nor U7553 (N_7553,N_6196,N_6770);
or U7554 (N_7554,N_6975,N_6037);
nor U7555 (N_7555,N_6840,N_6111);
or U7556 (N_7556,N_6922,N_6593);
or U7557 (N_7557,N_6051,N_6483);
nand U7558 (N_7558,N_6378,N_6699);
and U7559 (N_7559,N_6829,N_6217);
nand U7560 (N_7560,N_6734,N_6851);
and U7561 (N_7561,N_6240,N_6281);
and U7562 (N_7562,N_6588,N_6054);
nor U7563 (N_7563,N_6893,N_6364);
nand U7564 (N_7564,N_6605,N_6617);
nor U7565 (N_7565,N_6413,N_6629);
nand U7566 (N_7566,N_6414,N_6716);
nand U7567 (N_7567,N_6988,N_6986);
nand U7568 (N_7568,N_6055,N_6577);
nand U7569 (N_7569,N_6672,N_6358);
nor U7570 (N_7570,N_6856,N_6377);
nand U7571 (N_7571,N_6671,N_6322);
or U7572 (N_7572,N_6717,N_6757);
nor U7573 (N_7573,N_6173,N_6720);
and U7574 (N_7574,N_6423,N_6128);
and U7575 (N_7575,N_6071,N_6558);
and U7576 (N_7576,N_6466,N_6810);
or U7577 (N_7577,N_6207,N_6553);
nor U7578 (N_7578,N_6503,N_6090);
nand U7579 (N_7579,N_6205,N_6387);
nor U7580 (N_7580,N_6096,N_6384);
or U7581 (N_7581,N_6224,N_6007);
and U7582 (N_7582,N_6507,N_6519);
nor U7583 (N_7583,N_6585,N_6292);
and U7584 (N_7584,N_6389,N_6105);
nor U7585 (N_7585,N_6499,N_6704);
nand U7586 (N_7586,N_6345,N_6630);
nor U7587 (N_7587,N_6703,N_6278);
and U7588 (N_7588,N_6817,N_6434);
nand U7589 (N_7589,N_6698,N_6893);
and U7590 (N_7590,N_6968,N_6626);
nor U7591 (N_7591,N_6281,N_6637);
or U7592 (N_7592,N_6197,N_6764);
nor U7593 (N_7593,N_6425,N_6829);
or U7594 (N_7594,N_6291,N_6317);
nand U7595 (N_7595,N_6163,N_6520);
and U7596 (N_7596,N_6656,N_6894);
nor U7597 (N_7597,N_6541,N_6179);
or U7598 (N_7598,N_6262,N_6922);
nand U7599 (N_7599,N_6052,N_6777);
and U7600 (N_7600,N_6092,N_6001);
or U7601 (N_7601,N_6743,N_6605);
nand U7602 (N_7602,N_6170,N_6231);
nor U7603 (N_7603,N_6039,N_6460);
nor U7604 (N_7604,N_6693,N_6760);
or U7605 (N_7605,N_6153,N_6456);
nor U7606 (N_7606,N_6454,N_6392);
or U7607 (N_7607,N_6568,N_6417);
or U7608 (N_7608,N_6176,N_6292);
and U7609 (N_7609,N_6747,N_6012);
nor U7610 (N_7610,N_6003,N_6648);
nor U7611 (N_7611,N_6373,N_6650);
or U7612 (N_7612,N_6305,N_6548);
nand U7613 (N_7613,N_6532,N_6674);
nand U7614 (N_7614,N_6333,N_6608);
nand U7615 (N_7615,N_6954,N_6417);
nand U7616 (N_7616,N_6547,N_6237);
or U7617 (N_7617,N_6669,N_6000);
or U7618 (N_7618,N_6489,N_6016);
or U7619 (N_7619,N_6041,N_6275);
or U7620 (N_7620,N_6434,N_6586);
nor U7621 (N_7621,N_6918,N_6401);
or U7622 (N_7622,N_6015,N_6019);
or U7623 (N_7623,N_6654,N_6824);
or U7624 (N_7624,N_6475,N_6416);
or U7625 (N_7625,N_6817,N_6636);
or U7626 (N_7626,N_6563,N_6360);
nand U7627 (N_7627,N_6967,N_6109);
or U7628 (N_7628,N_6561,N_6549);
and U7629 (N_7629,N_6795,N_6497);
and U7630 (N_7630,N_6652,N_6657);
nor U7631 (N_7631,N_6641,N_6998);
nand U7632 (N_7632,N_6230,N_6598);
or U7633 (N_7633,N_6239,N_6619);
and U7634 (N_7634,N_6627,N_6110);
or U7635 (N_7635,N_6655,N_6562);
or U7636 (N_7636,N_6622,N_6030);
nand U7637 (N_7637,N_6301,N_6977);
nor U7638 (N_7638,N_6621,N_6912);
and U7639 (N_7639,N_6170,N_6902);
or U7640 (N_7640,N_6646,N_6561);
and U7641 (N_7641,N_6573,N_6490);
or U7642 (N_7642,N_6237,N_6305);
nor U7643 (N_7643,N_6812,N_6230);
nand U7644 (N_7644,N_6011,N_6155);
and U7645 (N_7645,N_6915,N_6457);
nor U7646 (N_7646,N_6452,N_6799);
nand U7647 (N_7647,N_6709,N_6891);
nand U7648 (N_7648,N_6366,N_6813);
nand U7649 (N_7649,N_6957,N_6478);
or U7650 (N_7650,N_6010,N_6788);
or U7651 (N_7651,N_6208,N_6171);
xnor U7652 (N_7652,N_6064,N_6739);
or U7653 (N_7653,N_6535,N_6920);
nor U7654 (N_7654,N_6869,N_6401);
nor U7655 (N_7655,N_6775,N_6674);
and U7656 (N_7656,N_6072,N_6193);
nand U7657 (N_7657,N_6004,N_6636);
nor U7658 (N_7658,N_6659,N_6207);
and U7659 (N_7659,N_6667,N_6231);
or U7660 (N_7660,N_6132,N_6572);
or U7661 (N_7661,N_6910,N_6432);
nand U7662 (N_7662,N_6513,N_6202);
and U7663 (N_7663,N_6131,N_6047);
nor U7664 (N_7664,N_6145,N_6380);
nor U7665 (N_7665,N_6140,N_6534);
xnor U7666 (N_7666,N_6227,N_6146);
nand U7667 (N_7667,N_6561,N_6190);
nand U7668 (N_7668,N_6792,N_6204);
and U7669 (N_7669,N_6416,N_6174);
and U7670 (N_7670,N_6105,N_6097);
or U7671 (N_7671,N_6244,N_6510);
nor U7672 (N_7672,N_6184,N_6713);
and U7673 (N_7673,N_6902,N_6171);
or U7674 (N_7674,N_6243,N_6183);
nor U7675 (N_7675,N_6627,N_6113);
nor U7676 (N_7676,N_6684,N_6121);
or U7677 (N_7677,N_6439,N_6222);
or U7678 (N_7678,N_6614,N_6271);
xnor U7679 (N_7679,N_6874,N_6882);
nand U7680 (N_7680,N_6957,N_6602);
nor U7681 (N_7681,N_6775,N_6264);
nand U7682 (N_7682,N_6110,N_6461);
or U7683 (N_7683,N_6752,N_6153);
xnor U7684 (N_7684,N_6014,N_6638);
nand U7685 (N_7685,N_6603,N_6670);
and U7686 (N_7686,N_6370,N_6046);
or U7687 (N_7687,N_6246,N_6166);
and U7688 (N_7688,N_6114,N_6917);
nor U7689 (N_7689,N_6493,N_6744);
nor U7690 (N_7690,N_6378,N_6402);
nor U7691 (N_7691,N_6422,N_6902);
or U7692 (N_7692,N_6461,N_6226);
nor U7693 (N_7693,N_6688,N_6552);
or U7694 (N_7694,N_6141,N_6189);
nor U7695 (N_7695,N_6427,N_6792);
nand U7696 (N_7696,N_6144,N_6901);
nand U7697 (N_7697,N_6769,N_6130);
and U7698 (N_7698,N_6928,N_6064);
nor U7699 (N_7699,N_6663,N_6569);
nor U7700 (N_7700,N_6304,N_6890);
and U7701 (N_7701,N_6674,N_6589);
or U7702 (N_7702,N_6405,N_6085);
nand U7703 (N_7703,N_6697,N_6765);
and U7704 (N_7704,N_6267,N_6111);
or U7705 (N_7705,N_6272,N_6538);
and U7706 (N_7706,N_6886,N_6491);
nand U7707 (N_7707,N_6143,N_6893);
and U7708 (N_7708,N_6465,N_6000);
and U7709 (N_7709,N_6120,N_6668);
and U7710 (N_7710,N_6304,N_6406);
nand U7711 (N_7711,N_6580,N_6114);
or U7712 (N_7712,N_6298,N_6121);
nor U7713 (N_7713,N_6924,N_6038);
nor U7714 (N_7714,N_6294,N_6777);
nand U7715 (N_7715,N_6794,N_6174);
nand U7716 (N_7716,N_6899,N_6171);
and U7717 (N_7717,N_6141,N_6405);
nor U7718 (N_7718,N_6497,N_6023);
nand U7719 (N_7719,N_6859,N_6456);
nor U7720 (N_7720,N_6368,N_6567);
and U7721 (N_7721,N_6862,N_6239);
and U7722 (N_7722,N_6587,N_6449);
nor U7723 (N_7723,N_6173,N_6330);
and U7724 (N_7724,N_6043,N_6194);
or U7725 (N_7725,N_6174,N_6716);
or U7726 (N_7726,N_6227,N_6210);
or U7727 (N_7727,N_6044,N_6874);
or U7728 (N_7728,N_6454,N_6770);
or U7729 (N_7729,N_6728,N_6157);
or U7730 (N_7730,N_6649,N_6006);
and U7731 (N_7731,N_6692,N_6528);
or U7732 (N_7732,N_6356,N_6263);
or U7733 (N_7733,N_6426,N_6862);
nor U7734 (N_7734,N_6559,N_6832);
or U7735 (N_7735,N_6529,N_6631);
nand U7736 (N_7736,N_6316,N_6594);
nand U7737 (N_7737,N_6321,N_6762);
nor U7738 (N_7738,N_6618,N_6014);
and U7739 (N_7739,N_6002,N_6578);
nand U7740 (N_7740,N_6258,N_6422);
nand U7741 (N_7741,N_6146,N_6352);
nor U7742 (N_7742,N_6563,N_6464);
nand U7743 (N_7743,N_6011,N_6820);
or U7744 (N_7744,N_6266,N_6372);
and U7745 (N_7745,N_6695,N_6084);
or U7746 (N_7746,N_6671,N_6347);
nor U7747 (N_7747,N_6263,N_6119);
nor U7748 (N_7748,N_6467,N_6972);
or U7749 (N_7749,N_6082,N_6351);
nor U7750 (N_7750,N_6407,N_6433);
or U7751 (N_7751,N_6738,N_6620);
or U7752 (N_7752,N_6818,N_6039);
nor U7753 (N_7753,N_6734,N_6911);
and U7754 (N_7754,N_6150,N_6816);
nor U7755 (N_7755,N_6393,N_6948);
or U7756 (N_7756,N_6039,N_6701);
or U7757 (N_7757,N_6586,N_6633);
or U7758 (N_7758,N_6532,N_6076);
nor U7759 (N_7759,N_6483,N_6985);
nor U7760 (N_7760,N_6813,N_6071);
nor U7761 (N_7761,N_6297,N_6595);
and U7762 (N_7762,N_6645,N_6322);
nor U7763 (N_7763,N_6190,N_6148);
or U7764 (N_7764,N_6021,N_6987);
and U7765 (N_7765,N_6426,N_6519);
or U7766 (N_7766,N_6461,N_6282);
or U7767 (N_7767,N_6278,N_6845);
or U7768 (N_7768,N_6760,N_6020);
nand U7769 (N_7769,N_6570,N_6695);
nand U7770 (N_7770,N_6773,N_6233);
nor U7771 (N_7771,N_6641,N_6090);
and U7772 (N_7772,N_6275,N_6794);
nand U7773 (N_7773,N_6854,N_6451);
nor U7774 (N_7774,N_6058,N_6363);
nor U7775 (N_7775,N_6149,N_6441);
or U7776 (N_7776,N_6300,N_6123);
nand U7777 (N_7777,N_6522,N_6271);
nand U7778 (N_7778,N_6994,N_6451);
and U7779 (N_7779,N_6953,N_6979);
or U7780 (N_7780,N_6835,N_6775);
or U7781 (N_7781,N_6166,N_6705);
xor U7782 (N_7782,N_6181,N_6660);
or U7783 (N_7783,N_6431,N_6750);
and U7784 (N_7784,N_6840,N_6236);
and U7785 (N_7785,N_6779,N_6835);
or U7786 (N_7786,N_6953,N_6851);
and U7787 (N_7787,N_6059,N_6701);
or U7788 (N_7788,N_6053,N_6347);
and U7789 (N_7789,N_6355,N_6828);
and U7790 (N_7790,N_6311,N_6066);
nor U7791 (N_7791,N_6735,N_6392);
or U7792 (N_7792,N_6729,N_6817);
nand U7793 (N_7793,N_6501,N_6218);
nand U7794 (N_7794,N_6032,N_6450);
nand U7795 (N_7795,N_6679,N_6138);
or U7796 (N_7796,N_6078,N_6804);
or U7797 (N_7797,N_6513,N_6281);
or U7798 (N_7798,N_6242,N_6005);
or U7799 (N_7799,N_6171,N_6434);
or U7800 (N_7800,N_6762,N_6217);
xor U7801 (N_7801,N_6899,N_6994);
nor U7802 (N_7802,N_6984,N_6804);
or U7803 (N_7803,N_6155,N_6920);
nor U7804 (N_7804,N_6050,N_6441);
and U7805 (N_7805,N_6466,N_6461);
xor U7806 (N_7806,N_6513,N_6990);
nor U7807 (N_7807,N_6387,N_6341);
or U7808 (N_7808,N_6674,N_6059);
or U7809 (N_7809,N_6474,N_6448);
and U7810 (N_7810,N_6548,N_6170);
nor U7811 (N_7811,N_6643,N_6007);
and U7812 (N_7812,N_6097,N_6608);
or U7813 (N_7813,N_6656,N_6132);
nor U7814 (N_7814,N_6578,N_6224);
nor U7815 (N_7815,N_6284,N_6148);
nor U7816 (N_7816,N_6843,N_6178);
nand U7817 (N_7817,N_6418,N_6730);
or U7818 (N_7818,N_6777,N_6466);
and U7819 (N_7819,N_6388,N_6706);
or U7820 (N_7820,N_6303,N_6229);
and U7821 (N_7821,N_6439,N_6367);
and U7822 (N_7822,N_6938,N_6197);
nand U7823 (N_7823,N_6723,N_6989);
nor U7824 (N_7824,N_6074,N_6231);
nand U7825 (N_7825,N_6863,N_6989);
nor U7826 (N_7826,N_6952,N_6104);
nand U7827 (N_7827,N_6187,N_6368);
nor U7828 (N_7828,N_6325,N_6867);
nor U7829 (N_7829,N_6216,N_6142);
and U7830 (N_7830,N_6542,N_6947);
or U7831 (N_7831,N_6755,N_6196);
nor U7832 (N_7832,N_6895,N_6185);
xor U7833 (N_7833,N_6242,N_6608);
or U7834 (N_7834,N_6280,N_6975);
or U7835 (N_7835,N_6186,N_6013);
nand U7836 (N_7836,N_6683,N_6370);
nor U7837 (N_7837,N_6203,N_6052);
nor U7838 (N_7838,N_6165,N_6767);
and U7839 (N_7839,N_6687,N_6225);
or U7840 (N_7840,N_6435,N_6866);
and U7841 (N_7841,N_6988,N_6778);
nand U7842 (N_7842,N_6685,N_6288);
nor U7843 (N_7843,N_6346,N_6805);
and U7844 (N_7844,N_6745,N_6088);
or U7845 (N_7845,N_6133,N_6406);
nand U7846 (N_7846,N_6142,N_6998);
nand U7847 (N_7847,N_6149,N_6075);
and U7848 (N_7848,N_6926,N_6117);
or U7849 (N_7849,N_6361,N_6065);
or U7850 (N_7850,N_6555,N_6512);
nand U7851 (N_7851,N_6402,N_6728);
nand U7852 (N_7852,N_6735,N_6229);
nor U7853 (N_7853,N_6511,N_6770);
nand U7854 (N_7854,N_6684,N_6010);
nand U7855 (N_7855,N_6631,N_6716);
and U7856 (N_7856,N_6304,N_6192);
and U7857 (N_7857,N_6036,N_6843);
or U7858 (N_7858,N_6074,N_6041);
nand U7859 (N_7859,N_6784,N_6343);
nor U7860 (N_7860,N_6530,N_6550);
nand U7861 (N_7861,N_6005,N_6536);
nor U7862 (N_7862,N_6422,N_6006);
or U7863 (N_7863,N_6289,N_6345);
and U7864 (N_7864,N_6877,N_6103);
or U7865 (N_7865,N_6447,N_6885);
nand U7866 (N_7866,N_6217,N_6873);
nand U7867 (N_7867,N_6771,N_6875);
nand U7868 (N_7868,N_6104,N_6802);
xor U7869 (N_7869,N_6044,N_6698);
nand U7870 (N_7870,N_6362,N_6622);
nand U7871 (N_7871,N_6071,N_6780);
or U7872 (N_7872,N_6008,N_6315);
nor U7873 (N_7873,N_6201,N_6737);
or U7874 (N_7874,N_6262,N_6365);
and U7875 (N_7875,N_6952,N_6717);
nand U7876 (N_7876,N_6072,N_6936);
or U7877 (N_7877,N_6395,N_6910);
nor U7878 (N_7878,N_6672,N_6263);
and U7879 (N_7879,N_6031,N_6300);
nor U7880 (N_7880,N_6190,N_6378);
or U7881 (N_7881,N_6032,N_6851);
nand U7882 (N_7882,N_6821,N_6248);
and U7883 (N_7883,N_6591,N_6486);
nor U7884 (N_7884,N_6816,N_6929);
nand U7885 (N_7885,N_6259,N_6683);
nor U7886 (N_7886,N_6851,N_6714);
and U7887 (N_7887,N_6484,N_6288);
and U7888 (N_7888,N_6559,N_6251);
nand U7889 (N_7889,N_6999,N_6099);
nand U7890 (N_7890,N_6729,N_6005);
nor U7891 (N_7891,N_6008,N_6004);
or U7892 (N_7892,N_6959,N_6252);
or U7893 (N_7893,N_6126,N_6340);
nand U7894 (N_7894,N_6450,N_6541);
or U7895 (N_7895,N_6451,N_6878);
and U7896 (N_7896,N_6237,N_6640);
and U7897 (N_7897,N_6893,N_6708);
and U7898 (N_7898,N_6453,N_6312);
or U7899 (N_7899,N_6780,N_6496);
and U7900 (N_7900,N_6545,N_6469);
nand U7901 (N_7901,N_6634,N_6556);
nand U7902 (N_7902,N_6104,N_6644);
and U7903 (N_7903,N_6535,N_6388);
or U7904 (N_7904,N_6999,N_6410);
or U7905 (N_7905,N_6108,N_6520);
nand U7906 (N_7906,N_6741,N_6501);
and U7907 (N_7907,N_6976,N_6756);
xor U7908 (N_7908,N_6073,N_6540);
or U7909 (N_7909,N_6134,N_6583);
nor U7910 (N_7910,N_6096,N_6850);
nand U7911 (N_7911,N_6834,N_6002);
nand U7912 (N_7912,N_6214,N_6979);
or U7913 (N_7913,N_6853,N_6792);
nand U7914 (N_7914,N_6588,N_6169);
and U7915 (N_7915,N_6943,N_6819);
or U7916 (N_7916,N_6775,N_6987);
nor U7917 (N_7917,N_6779,N_6243);
nor U7918 (N_7918,N_6122,N_6426);
or U7919 (N_7919,N_6628,N_6377);
or U7920 (N_7920,N_6549,N_6660);
nor U7921 (N_7921,N_6674,N_6835);
nor U7922 (N_7922,N_6718,N_6008);
nor U7923 (N_7923,N_6735,N_6596);
nand U7924 (N_7924,N_6249,N_6958);
nor U7925 (N_7925,N_6786,N_6258);
and U7926 (N_7926,N_6377,N_6235);
xnor U7927 (N_7927,N_6837,N_6053);
and U7928 (N_7928,N_6809,N_6849);
nand U7929 (N_7929,N_6101,N_6822);
nand U7930 (N_7930,N_6233,N_6042);
nor U7931 (N_7931,N_6449,N_6030);
nor U7932 (N_7932,N_6440,N_6999);
nand U7933 (N_7933,N_6053,N_6304);
nor U7934 (N_7934,N_6364,N_6295);
and U7935 (N_7935,N_6241,N_6042);
or U7936 (N_7936,N_6231,N_6865);
nor U7937 (N_7937,N_6789,N_6802);
nor U7938 (N_7938,N_6506,N_6672);
nor U7939 (N_7939,N_6633,N_6932);
nand U7940 (N_7940,N_6895,N_6208);
nor U7941 (N_7941,N_6454,N_6474);
nor U7942 (N_7942,N_6494,N_6908);
and U7943 (N_7943,N_6044,N_6368);
nand U7944 (N_7944,N_6405,N_6443);
nand U7945 (N_7945,N_6524,N_6128);
nand U7946 (N_7946,N_6500,N_6252);
nand U7947 (N_7947,N_6372,N_6265);
nor U7948 (N_7948,N_6010,N_6678);
nor U7949 (N_7949,N_6319,N_6081);
or U7950 (N_7950,N_6465,N_6257);
and U7951 (N_7951,N_6072,N_6329);
nor U7952 (N_7952,N_6478,N_6934);
or U7953 (N_7953,N_6093,N_6668);
or U7954 (N_7954,N_6041,N_6354);
or U7955 (N_7955,N_6676,N_6650);
or U7956 (N_7956,N_6883,N_6923);
and U7957 (N_7957,N_6829,N_6077);
nand U7958 (N_7958,N_6508,N_6196);
nand U7959 (N_7959,N_6318,N_6285);
or U7960 (N_7960,N_6681,N_6263);
and U7961 (N_7961,N_6857,N_6400);
nand U7962 (N_7962,N_6866,N_6845);
and U7963 (N_7963,N_6674,N_6009);
and U7964 (N_7964,N_6588,N_6985);
and U7965 (N_7965,N_6054,N_6029);
nand U7966 (N_7966,N_6094,N_6622);
nor U7967 (N_7967,N_6798,N_6704);
or U7968 (N_7968,N_6518,N_6798);
and U7969 (N_7969,N_6730,N_6221);
nor U7970 (N_7970,N_6095,N_6849);
xnor U7971 (N_7971,N_6439,N_6260);
and U7972 (N_7972,N_6176,N_6009);
and U7973 (N_7973,N_6192,N_6254);
nor U7974 (N_7974,N_6902,N_6285);
nor U7975 (N_7975,N_6198,N_6244);
or U7976 (N_7976,N_6495,N_6315);
nor U7977 (N_7977,N_6125,N_6979);
and U7978 (N_7978,N_6049,N_6700);
nand U7979 (N_7979,N_6198,N_6282);
nand U7980 (N_7980,N_6169,N_6179);
or U7981 (N_7981,N_6142,N_6792);
and U7982 (N_7982,N_6364,N_6583);
nor U7983 (N_7983,N_6550,N_6850);
and U7984 (N_7984,N_6043,N_6252);
or U7985 (N_7985,N_6951,N_6733);
nand U7986 (N_7986,N_6118,N_6077);
or U7987 (N_7987,N_6221,N_6986);
or U7988 (N_7988,N_6547,N_6212);
nand U7989 (N_7989,N_6505,N_6215);
and U7990 (N_7990,N_6987,N_6412);
nand U7991 (N_7991,N_6169,N_6469);
and U7992 (N_7992,N_6443,N_6886);
nor U7993 (N_7993,N_6966,N_6302);
nor U7994 (N_7994,N_6122,N_6822);
nand U7995 (N_7995,N_6395,N_6306);
and U7996 (N_7996,N_6779,N_6353);
and U7997 (N_7997,N_6598,N_6747);
or U7998 (N_7998,N_6660,N_6012);
xor U7999 (N_7999,N_6556,N_6363);
or U8000 (N_8000,N_7180,N_7991);
and U8001 (N_8001,N_7225,N_7556);
nand U8002 (N_8002,N_7072,N_7677);
nand U8003 (N_8003,N_7578,N_7674);
nand U8004 (N_8004,N_7142,N_7678);
nand U8005 (N_8005,N_7586,N_7730);
xor U8006 (N_8006,N_7226,N_7116);
nand U8007 (N_8007,N_7296,N_7319);
and U8008 (N_8008,N_7244,N_7601);
and U8009 (N_8009,N_7168,N_7326);
and U8010 (N_8010,N_7111,N_7502);
or U8011 (N_8011,N_7020,N_7394);
nor U8012 (N_8012,N_7806,N_7830);
and U8013 (N_8013,N_7918,N_7937);
and U8014 (N_8014,N_7763,N_7602);
nand U8015 (N_8015,N_7755,N_7553);
nand U8016 (N_8016,N_7949,N_7420);
nor U8017 (N_8017,N_7542,N_7143);
nand U8018 (N_8018,N_7236,N_7006);
nand U8019 (N_8019,N_7384,N_7560);
and U8020 (N_8020,N_7575,N_7768);
nor U8021 (N_8021,N_7695,N_7077);
and U8022 (N_8022,N_7365,N_7805);
nor U8023 (N_8023,N_7503,N_7290);
nand U8024 (N_8024,N_7467,N_7446);
nand U8025 (N_8025,N_7130,N_7416);
nor U8026 (N_8026,N_7252,N_7270);
nand U8027 (N_8027,N_7411,N_7689);
nor U8028 (N_8028,N_7486,N_7884);
and U8029 (N_8029,N_7975,N_7257);
nand U8030 (N_8030,N_7698,N_7623);
and U8031 (N_8031,N_7105,N_7259);
and U8032 (N_8032,N_7992,N_7759);
and U8033 (N_8033,N_7109,N_7375);
nor U8034 (N_8034,N_7412,N_7335);
nand U8035 (N_8035,N_7315,N_7426);
nand U8036 (N_8036,N_7841,N_7247);
or U8037 (N_8037,N_7620,N_7627);
and U8038 (N_8038,N_7559,N_7219);
nand U8039 (N_8039,N_7134,N_7612);
nand U8040 (N_8040,N_7320,N_7260);
and U8041 (N_8041,N_7492,N_7816);
or U8042 (N_8042,N_7714,N_7582);
nor U8043 (N_8043,N_7308,N_7484);
nand U8044 (N_8044,N_7428,N_7980);
and U8045 (N_8045,N_7908,N_7838);
or U8046 (N_8046,N_7849,N_7986);
or U8047 (N_8047,N_7670,N_7004);
nor U8048 (N_8048,N_7403,N_7432);
nor U8049 (N_8049,N_7833,N_7165);
and U8050 (N_8050,N_7039,N_7987);
nor U8051 (N_8051,N_7189,N_7699);
nand U8052 (N_8052,N_7463,N_7147);
nand U8053 (N_8053,N_7124,N_7464);
and U8054 (N_8054,N_7353,N_7438);
nand U8055 (N_8055,N_7622,N_7897);
or U8056 (N_8056,N_7187,N_7048);
or U8057 (N_8057,N_7227,N_7826);
nand U8058 (N_8058,N_7697,N_7823);
or U8059 (N_8059,N_7898,N_7241);
nand U8060 (N_8060,N_7842,N_7715);
and U8061 (N_8061,N_7812,N_7362);
and U8062 (N_8062,N_7984,N_7632);
nor U8063 (N_8063,N_7658,N_7572);
xor U8064 (N_8064,N_7704,N_7414);
xnor U8065 (N_8065,N_7899,N_7676);
nand U8066 (N_8066,N_7780,N_7835);
nand U8067 (N_8067,N_7358,N_7961);
or U8068 (N_8068,N_7756,N_7691);
nor U8069 (N_8069,N_7639,N_7700);
and U8070 (N_8070,N_7324,N_7153);
or U8071 (N_8071,N_7073,N_7558);
nor U8072 (N_8072,N_7643,N_7799);
or U8073 (N_8073,N_7907,N_7679);
nand U8074 (N_8074,N_7901,N_7278);
nor U8075 (N_8075,N_7728,N_7589);
and U8076 (N_8076,N_7435,N_7748);
or U8077 (N_8077,N_7204,N_7146);
nor U8078 (N_8078,N_7313,N_7138);
or U8079 (N_8079,N_7051,N_7212);
or U8080 (N_8080,N_7047,N_7211);
nor U8081 (N_8081,N_7738,N_7292);
and U8082 (N_8082,N_7186,N_7857);
or U8083 (N_8083,N_7177,N_7520);
nand U8084 (N_8084,N_7163,N_7543);
or U8085 (N_8085,N_7318,N_7500);
and U8086 (N_8086,N_7036,N_7644);
or U8087 (N_8087,N_7951,N_7049);
nor U8088 (N_8088,N_7333,N_7158);
and U8089 (N_8089,N_7108,N_7648);
or U8090 (N_8090,N_7652,N_7996);
nand U8091 (N_8091,N_7757,N_7417);
and U8092 (N_8092,N_7062,N_7911);
nor U8093 (N_8093,N_7903,N_7206);
nand U8094 (N_8094,N_7149,N_7303);
nand U8095 (N_8095,N_7924,N_7683);
or U8096 (N_8096,N_7374,N_7169);
or U8097 (N_8097,N_7409,N_7673);
nand U8098 (N_8098,N_7485,N_7473);
nand U8099 (N_8099,N_7793,N_7536);
and U8100 (N_8100,N_7468,N_7444);
or U8101 (N_8101,N_7462,N_7958);
nor U8102 (N_8102,N_7330,N_7282);
nor U8103 (N_8103,N_7990,N_7954);
nand U8104 (N_8104,N_7339,N_7203);
and U8105 (N_8105,N_7068,N_7064);
nand U8106 (N_8106,N_7499,N_7086);
and U8107 (N_8107,N_7224,N_7916);
and U8108 (N_8108,N_7494,N_7171);
and U8109 (N_8109,N_7367,N_7495);
nor U8110 (N_8110,N_7865,N_7873);
nor U8111 (N_8111,N_7406,N_7630);
or U8112 (N_8112,N_7571,N_7779);
xnor U8113 (N_8113,N_7915,N_7110);
or U8114 (N_8114,N_7482,N_7321);
and U8115 (N_8115,N_7496,N_7377);
nor U8116 (N_8116,N_7882,N_7708);
and U8117 (N_8117,N_7091,N_7803);
nand U8118 (N_8118,N_7606,N_7938);
or U8119 (N_8119,N_7385,N_7242);
nand U8120 (N_8120,N_7727,N_7968);
or U8121 (N_8121,N_7790,N_7490);
nand U8122 (N_8122,N_7526,N_7610);
or U8123 (N_8123,N_7185,N_7316);
nor U8124 (N_8124,N_7568,N_7513);
nor U8125 (N_8125,N_7096,N_7289);
nor U8126 (N_8126,N_7075,N_7533);
nand U8127 (N_8127,N_7076,N_7925);
nor U8128 (N_8128,N_7810,N_7624);
nor U8129 (N_8129,N_7767,N_7713);
nand U8130 (N_8130,N_7782,N_7523);
and U8131 (N_8131,N_7969,N_7722);
nor U8132 (N_8132,N_7262,N_7887);
and U8133 (N_8133,N_7564,N_7210);
or U8134 (N_8134,N_7030,N_7376);
nand U8135 (N_8135,N_7796,N_7245);
or U8136 (N_8136,N_7976,N_7615);
or U8137 (N_8137,N_7524,N_7607);
or U8138 (N_8138,N_7393,N_7354);
nand U8139 (N_8139,N_7479,N_7046);
or U8140 (N_8140,N_7232,N_7939);
or U8141 (N_8141,N_7603,N_7457);
or U8142 (N_8142,N_7345,N_7170);
or U8143 (N_8143,N_7735,N_7477);
nor U8144 (N_8144,N_7514,N_7650);
nor U8145 (N_8145,N_7044,N_7010);
nand U8146 (N_8146,N_7382,N_7867);
or U8147 (N_8147,N_7504,N_7974);
nand U8148 (N_8148,N_7295,N_7408);
or U8149 (N_8149,N_7703,N_7645);
or U8150 (N_8150,N_7709,N_7476);
or U8151 (N_8151,N_7660,N_7126);
and U8152 (N_8152,N_7929,N_7668);
nor U8153 (N_8153,N_7002,N_7593);
and U8154 (N_8154,N_7035,N_7363);
nand U8155 (N_8155,N_7872,N_7861);
nor U8156 (N_8156,N_7041,N_7877);
nor U8157 (N_8157,N_7264,N_7058);
nand U8158 (N_8158,N_7117,N_7253);
nand U8159 (N_8159,N_7856,N_7018);
or U8160 (N_8160,N_7285,N_7173);
or U8161 (N_8161,N_7718,N_7940);
and U8162 (N_8162,N_7979,N_7815);
and U8163 (N_8163,N_7251,N_7519);
nor U8164 (N_8164,N_7113,N_7896);
or U8165 (N_8165,N_7087,N_7478);
and U8166 (N_8166,N_7711,N_7263);
or U8167 (N_8167,N_7784,N_7902);
xor U8168 (N_8168,N_7125,N_7972);
nand U8169 (N_8169,N_7395,N_7577);
or U8170 (N_8170,N_7583,N_7405);
nand U8171 (N_8171,N_7088,N_7846);
or U8172 (N_8172,N_7818,N_7827);
or U8173 (N_8173,N_7100,N_7013);
nor U8174 (N_8174,N_7092,N_7066);
and U8175 (N_8175,N_7552,N_7864);
and U8176 (N_8176,N_7716,N_7380);
nor U8177 (N_8177,N_7063,N_7631);
nor U8178 (N_8178,N_7135,N_7895);
or U8179 (N_8179,N_7407,N_7913);
and U8180 (N_8180,N_7538,N_7923);
nand U8181 (N_8181,N_7137,N_7885);
or U8182 (N_8182,N_7122,N_7136);
nand U8183 (N_8183,N_7389,N_7928);
nor U8184 (N_8184,N_7860,N_7655);
or U8185 (N_8185,N_7014,N_7231);
nor U8186 (N_8186,N_7119,N_7300);
nand U8187 (N_8187,N_7009,N_7999);
nor U8188 (N_8188,N_7215,N_7447);
nand U8189 (N_8189,N_7297,N_7317);
nor U8190 (N_8190,N_7981,N_7220);
or U8191 (N_8191,N_7894,N_7900);
or U8192 (N_8192,N_7530,N_7466);
nand U8193 (N_8193,N_7343,N_7741);
or U8194 (N_8194,N_7788,N_7957);
and U8195 (N_8195,N_7982,N_7201);
nor U8196 (N_8196,N_7619,N_7331);
and U8197 (N_8197,N_7166,N_7555);
nor U8198 (N_8198,N_7207,N_7657);
nand U8199 (N_8199,N_7956,N_7754);
and U8200 (N_8200,N_7269,N_7007);
xnor U8201 (N_8201,N_7230,N_7917);
nor U8202 (N_8202,N_7256,N_7875);
nor U8203 (N_8203,N_7581,N_7717);
nand U8204 (N_8204,N_7775,N_7356);
nand U8205 (N_8205,N_7167,N_7022);
nor U8206 (N_8206,N_7946,N_7172);
nand U8207 (N_8207,N_7760,N_7618);
or U8208 (N_8208,N_7181,N_7789);
or U8209 (N_8209,N_7952,N_7346);
and U8210 (N_8210,N_7129,N_7539);
nand U8211 (N_8211,N_7995,N_7684);
and U8212 (N_8212,N_7766,N_7962);
or U8213 (N_8213,N_7642,N_7688);
or U8214 (N_8214,N_7104,N_7390);
nand U8215 (N_8215,N_7569,N_7919);
or U8216 (N_8216,N_7507,N_7712);
and U8217 (N_8217,N_7240,N_7156);
nor U8218 (N_8218,N_7521,N_7617);
nor U8219 (N_8219,N_7591,N_7460);
and U8220 (N_8220,N_7587,N_7157);
nor U8221 (N_8221,N_7505,N_7774);
nor U8222 (N_8222,N_7598,N_7840);
or U8223 (N_8223,N_7144,N_7629);
and U8224 (N_8224,N_7016,N_7792);
and U8225 (N_8225,N_7440,N_7011);
nand U8226 (N_8226,N_7123,N_7474);
and U8227 (N_8227,N_7566,N_7943);
nand U8228 (N_8228,N_7585,N_7509);
nand U8229 (N_8229,N_7855,N_7261);
nor U8230 (N_8230,N_7944,N_7284);
nor U8231 (N_8231,N_7419,N_7522);
or U8232 (N_8232,N_7848,N_7302);
nor U8233 (N_8233,N_7942,N_7905);
nor U8234 (N_8234,N_7445,N_7557);
nand U8235 (N_8235,N_7069,N_7879);
and U8236 (N_8236,N_7874,N_7150);
or U8237 (N_8237,N_7613,N_7233);
nand U8238 (N_8238,N_7489,N_7997);
or U8239 (N_8239,N_7636,N_7537);
and U8240 (N_8240,N_7311,N_7890);
nor U8241 (N_8241,N_7265,N_7139);
xor U8242 (N_8242,N_7732,N_7941);
nor U8243 (N_8243,N_7690,N_7360);
and U8244 (N_8244,N_7800,N_7675);
or U8245 (N_8245,N_7055,N_7026);
nand U8246 (N_8246,N_7392,N_7831);
or U8247 (N_8247,N_7776,N_7851);
and U8248 (N_8248,N_7191,N_7205);
and U8249 (N_8249,N_7439,N_7344);
and U8250 (N_8250,N_7948,N_7028);
nor U8251 (N_8251,N_7229,N_7825);
or U8252 (N_8252,N_7945,N_7854);
nor U8253 (N_8253,N_7054,N_7272);
and U8254 (N_8254,N_7162,N_7038);
and U8255 (N_8255,N_7071,N_7822);
nand U8256 (N_8256,N_7280,N_7305);
nor U8257 (N_8257,N_7950,N_7661);
or U8258 (N_8258,N_7294,N_7043);
nor U8259 (N_8259,N_7931,N_7880);
nor U8260 (N_8260,N_7588,N_7646);
nor U8261 (N_8261,N_7074,N_7930);
nor U8262 (N_8262,N_7740,N_7025);
and U8263 (N_8263,N_7037,N_7031);
nor U8264 (N_8264,N_7527,N_7161);
nor U8265 (N_8265,N_7634,N_7341);
and U8266 (N_8266,N_7275,N_7449);
and U8267 (N_8267,N_7199,N_7298);
and U8268 (N_8268,N_7239,N_7337);
and U8269 (N_8269,N_7659,N_7770);
nand U8270 (N_8270,N_7140,N_7761);
nand U8271 (N_8271,N_7508,N_7084);
and U8272 (N_8272,N_7461,N_7608);
nor U8273 (N_8273,N_7535,N_7706);
or U8274 (N_8274,N_7985,N_7567);
nand U8275 (N_8275,N_7510,N_7785);
or U8276 (N_8276,N_7451,N_7425);
nor U8277 (N_8277,N_7798,N_7746);
and U8278 (N_8278,N_7693,N_7621);
nand U8279 (N_8279,N_7744,N_7807);
nand U8280 (N_8280,N_7531,N_7596);
and U8281 (N_8281,N_7966,N_7115);
nor U8282 (N_8282,N_7164,N_7291);
or U8283 (N_8283,N_7663,N_7254);
nor U8284 (N_8284,N_7604,N_7102);
or U8285 (N_8285,N_7769,N_7131);
or U8286 (N_8286,N_7057,N_7061);
nand U8287 (N_8287,N_7085,N_7065);
nand U8288 (N_8288,N_7762,N_7914);
nor U8289 (N_8289,N_7743,N_7379);
nor U8290 (N_8290,N_7179,N_7029);
nor U8291 (N_8291,N_7921,N_7506);
or U8292 (N_8292,N_7863,N_7352);
or U8293 (N_8293,N_7633,N_7828);
or U8294 (N_8294,N_7758,N_7200);
and U8295 (N_8295,N_7368,N_7731);
nand U8296 (N_8296,N_7332,N_7653);
nand U8297 (N_8297,N_7483,N_7042);
nor U8298 (N_8298,N_7024,N_7853);
and U8299 (N_8299,N_7176,N_7196);
nor U8300 (N_8300,N_7101,N_7594);
and U8301 (N_8301,N_7198,N_7097);
and U8302 (N_8302,N_7431,N_7488);
nor U8303 (N_8303,N_7491,N_7306);
and U8304 (N_8304,N_7248,N_7751);
or U8305 (N_8305,N_7934,N_7310);
or U8306 (N_8306,N_7859,N_7733);
nand U8307 (N_8307,N_7920,N_7933);
nor U8308 (N_8308,N_7843,N_7223);
and U8309 (N_8309,N_7283,N_7402);
nor U8310 (N_8310,N_7287,N_7059);
nand U8311 (N_8311,N_7103,N_7373);
nand U8312 (N_8312,N_7288,N_7081);
and U8313 (N_8313,N_7237,N_7813);
nand U8314 (N_8314,N_7183,N_7545);
or U8315 (N_8315,N_7145,N_7960);
and U8316 (N_8316,N_7834,N_7672);
or U8317 (N_8317,N_7197,N_7436);
nor U8318 (N_8318,N_7702,N_7692);
nor U8319 (N_8319,N_7396,N_7079);
nor U8320 (N_8320,N_7753,N_7616);
and U8321 (N_8321,N_7450,N_7573);
nor U8322 (N_8322,N_7953,N_7935);
nand U8323 (N_8323,N_7628,N_7970);
nor U8324 (N_8324,N_7654,N_7366);
nor U8325 (N_8325,N_7973,N_7551);
or U8326 (N_8326,N_7993,N_7094);
and U8327 (N_8327,N_7437,N_7600);
nand U8328 (N_8328,N_7750,N_7497);
xnor U8329 (N_8329,N_7312,N_7737);
or U8330 (N_8330,N_7133,N_7347);
or U8331 (N_8331,N_7955,N_7481);
or U8332 (N_8332,N_7534,N_7413);
nor U8333 (N_8333,N_7994,N_7216);
or U8334 (N_8334,N_7487,N_7787);
nor U8335 (N_8335,N_7829,N_7794);
nor U8336 (N_8336,N_7682,N_7400);
and U8337 (N_8337,N_7977,N_7511);
nand U8338 (N_8338,N_7355,N_7404);
or U8339 (N_8339,N_7273,N_7371);
nor U8340 (N_8340,N_7584,N_7562);
or U8341 (N_8341,N_7340,N_7391);
nand U8342 (N_8342,N_7095,N_7926);
nor U8343 (N_8343,N_7881,N_7082);
or U8344 (N_8344,N_7141,N_7736);
nand U8345 (N_8345,N_7370,N_7745);
and U8346 (N_8346,N_7434,N_7597);
or U8347 (N_8347,N_7611,N_7155);
and U8348 (N_8348,N_7023,N_7008);
nor U8349 (N_8349,N_7192,N_7878);
or U8350 (N_8350,N_7554,N_7299);
and U8351 (N_8351,N_7458,N_7070);
nor U8352 (N_8352,N_7429,N_7060);
nor U8353 (N_8353,N_7871,N_7705);
nor U8354 (N_8354,N_7868,N_7862);
nand U8355 (N_8355,N_7228,N_7824);
and U8356 (N_8356,N_7837,N_7387);
nor U8357 (N_8357,N_7327,N_7338);
and U8358 (N_8358,N_7786,N_7415);
nand U8359 (N_8359,N_7563,N_7032);
or U8360 (N_8360,N_7614,N_7114);
or U8361 (N_8361,N_7217,N_7040);
nor U8362 (N_8362,N_7243,N_7817);
and U8363 (N_8363,N_7012,N_7640);
or U8364 (N_8364,N_7369,N_7529);
or U8365 (N_8365,N_7729,N_7719);
nor U8366 (N_8366,N_7361,N_7080);
nand U8367 (N_8367,N_7099,N_7869);
and U8368 (N_8368,N_7765,N_7399);
nand U8369 (N_8369,N_7430,N_7681);
and U8370 (N_8370,N_7696,N_7159);
nor U8371 (N_8371,N_7329,N_7238);
nand U8372 (N_8372,N_7423,N_7725);
or U8373 (N_8373,N_7307,N_7809);
nor U8374 (N_8374,N_7067,N_7132);
nand U8375 (N_8375,N_7246,N_7574);
nor U8376 (N_8376,N_7772,N_7194);
nand U8377 (N_8377,N_7221,N_7107);
nand U8378 (N_8378,N_7271,N_7286);
or U8379 (N_8379,N_7590,N_7561);
nand U8380 (N_8380,N_7249,N_7469);
or U8381 (N_8381,N_7421,N_7443);
or U8382 (N_8382,N_7184,N_7541);
or U8383 (N_8383,N_7322,N_7255);
and U8384 (N_8384,N_7532,N_7005);
or U8385 (N_8385,N_7625,N_7418);
and U8386 (N_8386,N_7671,N_7666);
or U8387 (N_8387,N_7193,N_7680);
or U8388 (N_8388,N_7027,N_7664);
nor U8389 (N_8389,N_7098,N_7250);
or U8390 (N_8390,N_7304,N_7342);
and U8391 (N_8391,N_7971,N_7154);
nand U8392 (N_8392,N_7638,N_7988);
or U8393 (N_8393,N_7819,N_7349);
or U8394 (N_8394,N_7267,N_7876);
and U8395 (N_8395,N_7963,N_7820);
nand U8396 (N_8396,N_7093,N_7427);
or U8397 (N_8397,N_7364,N_7752);
and U8398 (N_8398,N_7351,N_7381);
nand U8399 (N_8399,N_7936,N_7540);
nand U8400 (N_8400,N_7323,N_7626);
nand U8401 (N_8401,N_7001,N_7802);
and U8402 (N_8402,N_7281,N_7148);
or U8403 (N_8403,N_7442,N_7685);
nand U8404 (N_8404,N_7325,N_7662);
nand U8405 (N_8405,N_7127,N_7647);
nand U8406 (N_8406,N_7605,N_7512);
nor U8407 (N_8407,N_7383,N_7850);
or U8408 (N_8408,N_7694,N_7964);
or U8409 (N_8409,N_7637,N_7866);
and U8410 (N_8410,N_7309,N_7359);
nand U8411 (N_8411,N_7795,N_7083);
nor U8412 (N_8412,N_7019,N_7889);
or U8413 (N_8413,N_7544,N_7465);
and U8414 (N_8414,N_7797,N_7386);
nand U8415 (N_8415,N_7045,N_7651);
or U8416 (N_8416,N_7517,N_7978);
and U8417 (N_8417,N_7839,N_7515);
nand U8418 (N_8418,N_7764,N_7274);
nor U8419 (N_8419,N_7175,N_7279);
nand U8420 (N_8420,N_7471,N_7214);
nor U8421 (N_8421,N_7773,N_7410);
nand U8422 (N_8422,N_7548,N_7965);
nor U8423 (N_8423,N_7433,N_7456);
nor U8424 (N_8424,N_7152,N_7053);
nand U8425 (N_8425,N_7348,N_7003);
nor U8426 (N_8426,N_7998,N_7493);
or U8427 (N_8427,N_7777,N_7334);
nand U8428 (N_8428,N_7922,N_7470);
and U8429 (N_8429,N_7641,N_7821);
nand U8430 (N_8430,N_7547,N_7480);
nor U8431 (N_8431,N_7720,N_7665);
nor U8432 (N_8432,N_7277,N_7128);
or U8433 (N_8433,N_7814,N_7870);
nor U8434 (N_8434,N_7090,N_7858);
or U8435 (N_8435,N_7742,N_7452);
nor U8436 (N_8436,N_7906,N_7441);
or U8437 (N_8437,N_7888,N_7686);
and U8438 (N_8438,N_7182,N_7707);
nor U8439 (N_8439,N_7579,N_7580);
nor U8440 (N_8440,N_7845,N_7844);
nor U8441 (N_8441,N_7378,N_7771);
nand U8442 (N_8442,N_7314,N_7208);
nand U8443 (N_8443,N_7448,N_7983);
xor U8444 (N_8444,N_7190,N_7893);
or U8445 (N_8445,N_7932,N_7687);
nor U8446 (N_8446,N_7576,N_7218);
or U8447 (N_8447,N_7886,N_7266);
and U8448 (N_8448,N_7609,N_7565);
or U8449 (N_8449,N_7202,N_7398);
nor U8450 (N_8450,N_7120,N_7160);
or U8451 (N_8451,N_7089,N_7669);
nand U8452 (N_8452,N_7516,N_7454);
nand U8453 (N_8453,N_7017,N_7546);
or U8454 (N_8454,N_7832,N_7891);
or U8455 (N_8455,N_7453,N_7422);
or U8456 (N_8456,N_7724,N_7501);
and U8457 (N_8457,N_7549,N_7989);
nor U8458 (N_8458,N_7912,N_7293);
or U8459 (N_8459,N_7112,N_7710);
nand U8460 (N_8460,N_7947,N_7424);
and U8461 (N_8461,N_7472,N_7749);
or U8462 (N_8462,N_7301,N_7667);
nand U8463 (N_8463,N_7892,N_7967);
nor U8464 (N_8464,N_7276,N_7151);
nor U8465 (N_8465,N_7525,N_7778);
or U8466 (N_8466,N_7078,N_7213);
nor U8467 (N_8467,N_7033,N_7235);
nor U8468 (N_8468,N_7804,N_7927);
nand U8469 (N_8469,N_7015,N_7328);
nor U8470 (N_8470,N_7388,N_7550);
nor U8471 (N_8471,N_7372,N_7350);
or U8472 (N_8472,N_7781,N_7498);
nor U8473 (N_8473,N_7726,N_7050);
nand U8474 (N_8474,N_7883,N_7739);
nor U8475 (N_8475,N_7847,N_7397);
nand U8476 (N_8476,N_7121,N_7052);
nand U8477 (N_8477,N_7528,N_7357);
nand U8478 (N_8478,N_7701,N_7401);
nand U8479 (N_8479,N_7904,N_7808);
or U8480 (N_8480,N_7209,N_7455);
or U8481 (N_8481,N_7909,N_7118);
and U8482 (N_8482,N_7910,N_7595);
nand U8483 (N_8483,N_7836,N_7459);
or U8484 (N_8484,N_7178,N_7222);
nand U8485 (N_8485,N_7635,N_7475);
or U8486 (N_8486,N_7592,N_7195);
nand U8487 (N_8487,N_7518,N_7599);
nand U8488 (N_8488,N_7656,N_7234);
or U8489 (N_8489,N_7811,N_7000);
nand U8490 (N_8490,N_7056,N_7336);
and U8491 (N_8491,N_7747,N_7106);
nand U8492 (N_8492,N_7734,N_7723);
or U8493 (N_8493,N_7021,N_7570);
or U8494 (N_8494,N_7783,N_7791);
and U8495 (N_8495,N_7801,N_7649);
and U8496 (N_8496,N_7268,N_7959);
nor U8497 (N_8497,N_7034,N_7721);
nand U8498 (N_8498,N_7188,N_7174);
nand U8499 (N_8499,N_7258,N_7852);
or U8500 (N_8500,N_7984,N_7722);
and U8501 (N_8501,N_7918,N_7883);
and U8502 (N_8502,N_7536,N_7543);
or U8503 (N_8503,N_7355,N_7387);
nand U8504 (N_8504,N_7310,N_7764);
nor U8505 (N_8505,N_7231,N_7757);
nor U8506 (N_8506,N_7898,N_7665);
and U8507 (N_8507,N_7014,N_7591);
nor U8508 (N_8508,N_7398,N_7447);
nor U8509 (N_8509,N_7255,N_7333);
and U8510 (N_8510,N_7798,N_7374);
or U8511 (N_8511,N_7956,N_7409);
nand U8512 (N_8512,N_7928,N_7979);
and U8513 (N_8513,N_7539,N_7121);
nor U8514 (N_8514,N_7837,N_7422);
or U8515 (N_8515,N_7951,N_7548);
nand U8516 (N_8516,N_7228,N_7510);
nand U8517 (N_8517,N_7777,N_7725);
or U8518 (N_8518,N_7092,N_7563);
nor U8519 (N_8519,N_7347,N_7961);
nor U8520 (N_8520,N_7146,N_7071);
and U8521 (N_8521,N_7795,N_7713);
nor U8522 (N_8522,N_7961,N_7033);
nor U8523 (N_8523,N_7677,N_7959);
nand U8524 (N_8524,N_7554,N_7631);
and U8525 (N_8525,N_7793,N_7092);
nand U8526 (N_8526,N_7366,N_7227);
and U8527 (N_8527,N_7958,N_7811);
nor U8528 (N_8528,N_7359,N_7123);
and U8529 (N_8529,N_7711,N_7498);
and U8530 (N_8530,N_7978,N_7257);
and U8531 (N_8531,N_7334,N_7757);
nor U8532 (N_8532,N_7876,N_7745);
and U8533 (N_8533,N_7620,N_7718);
nor U8534 (N_8534,N_7864,N_7738);
or U8535 (N_8535,N_7435,N_7845);
and U8536 (N_8536,N_7421,N_7586);
and U8537 (N_8537,N_7178,N_7495);
nor U8538 (N_8538,N_7399,N_7229);
nor U8539 (N_8539,N_7840,N_7718);
nand U8540 (N_8540,N_7931,N_7679);
nor U8541 (N_8541,N_7227,N_7361);
nor U8542 (N_8542,N_7018,N_7049);
and U8543 (N_8543,N_7981,N_7002);
and U8544 (N_8544,N_7920,N_7117);
and U8545 (N_8545,N_7434,N_7294);
nor U8546 (N_8546,N_7421,N_7346);
and U8547 (N_8547,N_7441,N_7933);
and U8548 (N_8548,N_7622,N_7620);
nand U8549 (N_8549,N_7407,N_7518);
nor U8550 (N_8550,N_7720,N_7010);
or U8551 (N_8551,N_7105,N_7909);
nand U8552 (N_8552,N_7977,N_7261);
or U8553 (N_8553,N_7393,N_7333);
nand U8554 (N_8554,N_7122,N_7770);
nand U8555 (N_8555,N_7153,N_7563);
or U8556 (N_8556,N_7598,N_7694);
nand U8557 (N_8557,N_7827,N_7890);
and U8558 (N_8558,N_7175,N_7540);
or U8559 (N_8559,N_7299,N_7890);
nand U8560 (N_8560,N_7569,N_7252);
or U8561 (N_8561,N_7401,N_7081);
nand U8562 (N_8562,N_7228,N_7158);
nand U8563 (N_8563,N_7805,N_7588);
nand U8564 (N_8564,N_7946,N_7793);
or U8565 (N_8565,N_7695,N_7448);
nand U8566 (N_8566,N_7331,N_7510);
or U8567 (N_8567,N_7913,N_7966);
and U8568 (N_8568,N_7303,N_7109);
or U8569 (N_8569,N_7418,N_7824);
nor U8570 (N_8570,N_7674,N_7167);
or U8571 (N_8571,N_7624,N_7594);
nand U8572 (N_8572,N_7089,N_7578);
or U8573 (N_8573,N_7662,N_7467);
nand U8574 (N_8574,N_7720,N_7778);
nand U8575 (N_8575,N_7431,N_7209);
and U8576 (N_8576,N_7045,N_7830);
or U8577 (N_8577,N_7180,N_7763);
nand U8578 (N_8578,N_7941,N_7284);
nor U8579 (N_8579,N_7079,N_7137);
and U8580 (N_8580,N_7623,N_7881);
nor U8581 (N_8581,N_7837,N_7093);
nor U8582 (N_8582,N_7252,N_7278);
nand U8583 (N_8583,N_7736,N_7386);
nand U8584 (N_8584,N_7607,N_7288);
nor U8585 (N_8585,N_7738,N_7798);
or U8586 (N_8586,N_7890,N_7883);
nor U8587 (N_8587,N_7834,N_7969);
nand U8588 (N_8588,N_7463,N_7593);
or U8589 (N_8589,N_7125,N_7042);
and U8590 (N_8590,N_7889,N_7962);
or U8591 (N_8591,N_7664,N_7450);
or U8592 (N_8592,N_7520,N_7554);
or U8593 (N_8593,N_7460,N_7817);
nor U8594 (N_8594,N_7434,N_7666);
nand U8595 (N_8595,N_7678,N_7016);
or U8596 (N_8596,N_7919,N_7061);
and U8597 (N_8597,N_7776,N_7461);
nor U8598 (N_8598,N_7072,N_7321);
nor U8599 (N_8599,N_7375,N_7393);
xnor U8600 (N_8600,N_7690,N_7071);
nor U8601 (N_8601,N_7938,N_7217);
nor U8602 (N_8602,N_7462,N_7448);
or U8603 (N_8603,N_7390,N_7725);
nor U8604 (N_8604,N_7419,N_7521);
nand U8605 (N_8605,N_7619,N_7774);
or U8606 (N_8606,N_7660,N_7382);
nand U8607 (N_8607,N_7872,N_7189);
nor U8608 (N_8608,N_7605,N_7341);
nor U8609 (N_8609,N_7014,N_7335);
nor U8610 (N_8610,N_7483,N_7036);
or U8611 (N_8611,N_7096,N_7478);
nor U8612 (N_8612,N_7113,N_7765);
nor U8613 (N_8613,N_7574,N_7085);
or U8614 (N_8614,N_7155,N_7428);
or U8615 (N_8615,N_7293,N_7722);
xnor U8616 (N_8616,N_7220,N_7048);
and U8617 (N_8617,N_7021,N_7935);
and U8618 (N_8618,N_7492,N_7936);
or U8619 (N_8619,N_7687,N_7637);
or U8620 (N_8620,N_7507,N_7751);
or U8621 (N_8621,N_7435,N_7264);
or U8622 (N_8622,N_7271,N_7029);
and U8623 (N_8623,N_7756,N_7121);
nand U8624 (N_8624,N_7628,N_7159);
xor U8625 (N_8625,N_7610,N_7695);
nor U8626 (N_8626,N_7194,N_7274);
nor U8627 (N_8627,N_7843,N_7326);
nor U8628 (N_8628,N_7934,N_7700);
nand U8629 (N_8629,N_7070,N_7309);
nor U8630 (N_8630,N_7255,N_7795);
and U8631 (N_8631,N_7138,N_7645);
nor U8632 (N_8632,N_7595,N_7040);
and U8633 (N_8633,N_7916,N_7154);
nor U8634 (N_8634,N_7828,N_7453);
nor U8635 (N_8635,N_7924,N_7356);
and U8636 (N_8636,N_7459,N_7727);
nor U8637 (N_8637,N_7926,N_7148);
nor U8638 (N_8638,N_7391,N_7347);
or U8639 (N_8639,N_7224,N_7787);
or U8640 (N_8640,N_7077,N_7027);
and U8641 (N_8641,N_7000,N_7470);
nand U8642 (N_8642,N_7727,N_7408);
or U8643 (N_8643,N_7982,N_7050);
nor U8644 (N_8644,N_7641,N_7305);
nand U8645 (N_8645,N_7811,N_7386);
nand U8646 (N_8646,N_7990,N_7756);
nor U8647 (N_8647,N_7286,N_7068);
nand U8648 (N_8648,N_7823,N_7995);
nor U8649 (N_8649,N_7237,N_7505);
nand U8650 (N_8650,N_7927,N_7822);
nand U8651 (N_8651,N_7041,N_7530);
or U8652 (N_8652,N_7509,N_7701);
or U8653 (N_8653,N_7173,N_7720);
nor U8654 (N_8654,N_7006,N_7122);
nand U8655 (N_8655,N_7881,N_7457);
or U8656 (N_8656,N_7514,N_7092);
nand U8657 (N_8657,N_7100,N_7227);
nand U8658 (N_8658,N_7765,N_7220);
nand U8659 (N_8659,N_7750,N_7821);
nand U8660 (N_8660,N_7152,N_7538);
nand U8661 (N_8661,N_7908,N_7145);
and U8662 (N_8662,N_7650,N_7855);
or U8663 (N_8663,N_7468,N_7639);
xor U8664 (N_8664,N_7329,N_7205);
and U8665 (N_8665,N_7872,N_7887);
and U8666 (N_8666,N_7559,N_7639);
nand U8667 (N_8667,N_7691,N_7602);
or U8668 (N_8668,N_7777,N_7355);
nand U8669 (N_8669,N_7609,N_7185);
and U8670 (N_8670,N_7612,N_7111);
and U8671 (N_8671,N_7260,N_7949);
nor U8672 (N_8672,N_7172,N_7074);
nor U8673 (N_8673,N_7575,N_7512);
nor U8674 (N_8674,N_7053,N_7741);
nor U8675 (N_8675,N_7437,N_7598);
nor U8676 (N_8676,N_7194,N_7280);
or U8677 (N_8677,N_7480,N_7464);
nand U8678 (N_8678,N_7163,N_7571);
nor U8679 (N_8679,N_7837,N_7105);
nand U8680 (N_8680,N_7946,N_7807);
and U8681 (N_8681,N_7755,N_7156);
nor U8682 (N_8682,N_7655,N_7010);
nor U8683 (N_8683,N_7792,N_7169);
or U8684 (N_8684,N_7077,N_7159);
nor U8685 (N_8685,N_7426,N_7952);
nand U8686 (N_8686,N_7166,N_7971);
or U8687 (N_8687,N_7396,N_7433);
nand U8688 (N_8688,N_7306,N_7150);
and U8689 (N_8689,N_7425,N_7671);
nand U8690 (N_8690,N_7785,N_7306);
nor U8691 (N_8691,N_7200,N_7870);
nor U8692 (N_8692,N_7937,N_7813);
nand U8693 (N_8693,N_7781,N_7453);
nand U8694 (N_8694,N_7726,N_7480);
nor U8695 (N_8695,N_7634,N_7113);
nand U8696 (N_8696,N_7740,N_7158);
or U8697 (N_8697,N_7471,N_7858);
nand U8698 (N_8698,N_7728,N_7733);
and U8699 (N_8699,N_7942,N_7931);
and U8700 (N_8700,N_7340,N_7734);
and U8701 (N_8701,N_7469,N_7221);
or U8702 (N_8702,N_7554,N_7561);
and U8703 (N_8703,N_7003,N_7822);
or U8704 (N_8704,N_7048,N_7151);
or U8705 (N_8705,N_7475,N_7601);
or U8706 (N_8706,N_7605,N_7839);
or U8707 (N_8707,N_7766,N_7336);
nand U8708 (N_8708,N_7642,N_7310);
nor U8709 (N_8709,N_7579,N_7438);
and U8710 (N_8710,N_7688,N_7008);
or U8711 (N_8711,N_7033,N_7850);
and U8712 (N_8712,N_7083,N_7273);
and U8713 (N_8713,N_7592,N_7803);
and U8714 (N_8714,N_7629,N_7572);
nand U8715 (N_8715,N_7261,N_7904);
nor U8716 (N_8716,N_7458,N_7014);
or U8717 (N_8717,N_7685,N_7676);
and U8718 (N_8718,N_7538,N_7100);
nor U8719 (N_8719,N_7929,N_7418);
nor U8720 (N_8720,N_7831,N_7824);
or U8721 (N_8721,N_7732,N_7933);
nand U8722 (N_8722,N_7302,N_7376);
xor U8723 (N_8723,N_7304,N_7750);
or U8724 (N_8724,N_7682,N_7922);
or U8725 (N_8725,N_7822,N_7219);
and U8726 (N_8726,N_7075,N_7738);
nand U8727 (N_8727,N_7747,N_7844);
or U8728 (N_8728,N_7616,N_7908);
or U8729 (N_8729,N_7770,N_7702);
or U8730 (N_8730,N_7437,N_7679);
nand U8731 (N_8731,N_7695,N_7842);
nand U8732 (N_8732,N_7342,N_7887);
nor U8733 (N_8733,N_7747,N_7124);
xor U8734 (N_8734,N_7357,N_7121);
and U8735 (N_8735,N_7352,N_7867);
or U8736 (N_8736,N_7819,N_7102);
or U8737 (N_8737,N_7489,N_7691);
nor U8738 (N_8738,N_7678,N_7277);
nor U8739 (N_8739,N_7751,N_7630);
nand U8740 (N_8740,N_7582,N_7164);
nor U8741 (N_8741,N_7361,N_7189);
nor U8742 (N_8742,N_7919,N_7314);
nor U8743 (N_8743,N_7786,N_7541);
and U8744 (N_8744,N_7421,N_7513);
or U8745 (N_8745,N_7663,N_7511);
or U8746 (N_8746,N_7452,N_7009);
and U8747 (N_8747,N_7264,N_7918);
nor U8748 (N_8748,N_7959,N_7688);
and U8749 (N_8749,N_7084,N_7221);
or U8750 (N_8750,N_7760,N_7044);
nor U8751 (N_8751,N_7899,N_7258);
nand U8752 (N_8752,N_7624,N_7572);
and U8753 (N_8753,N_7642,N_7473);
and U8754 (N_8754,N_7095,N_7414);
nand U8755 (N_8755,N_7228,N_7247);
nand U8756 (N_8756,N_7771,N_7250);
nor U8757 (N_8757,N_7783,N_7255);
nand U8758 (N_8758,N_7926,N_7950);
or U8759 (N_8759,N_7400,N_7798);
nand U8760 (N_8760,N_7189,N_7080);
and U8761 (N_8761,N_7792,N_7241);
and U8762 (N_8762,N_7932,N_7715);
nor U8763 (N_8763,N_7487,N_7743);
nor U8764 (N_8764,N_7016,N_7818);
nand U8765 (N_8765,N_7379,N_7471);
nor U8766 (N_8766,N_7673,N_7020);
nand U8767 (N_8767,N_7732,N_7676);
and U8768 (N_8768,N_7533,N_7492);
nand U8769 (N_8769,N_7321,N_7135);
nor U8770 (N_8770,N_7050,N_7458);
nand U8771 (N_8771,N_7986,N_7255);
nand U8772 (N_8772,N_7381,N_7762);
nand U8773 (N_8773,N_7718,N_7609);
xor U8774 (N_8774,N_7709,N_7182);
or U8775 (N_8775,N_7833,N_7568);
and U8776 (N_8776,N_7509,N_7439);
nand U8777 (N_8777,N_7516,N_7094);
or U8778 (N_8778,N_7272,N_7926);
or U8779 (N_8779,N_7308,N_7193);
and U8780 (N_8780,N_7717,N_7176);
nand U8781 (N_8781,N_7584,N_7024);
nand U8782 (N_8782,N_7186,N_7905);
nand U8783 (N_8783,N_7880,N_7993);
and U8784 (N_8784,N_7968,N_7567);
nor U8785 (N_8785,N_7068,N_7399);
or U8786 (N_8786,N_7487,N_7778);
nand U8787 (N_8787,N_7346,N_7262);
and U8788 (N_8788,N_7840,N_7907);
or U8789 (N_8789,N_7722,N_7675);
or U8790 (N_8790,N_7900,N_7059);
nor U8791 (N_8791,N_7382,N_7756);
nand U8792 (N_8792,N_7762,N_7109);
and U8793 (N_8793,N_7633,N_7799);
nor U8794 (N_8794,N_7016,N_7018);
or U8795 (N_8795,N_7220,N_7844);
and U8796 (N_8796,N_7605,N_7834);
nand U8797 (N_8797,N_7492,N_7709);
nand U8798 (N_8798,N_7705,N_7494);
and U8799 (N_8799,N_7779,N_7430);
nor U8800 (N_8800,N_7407,N_7691);
nand U8801 (N_8801,N_7848,N_7027);
or U8802 (N_8802,N_7939,N_7692);
nor U8803 (N_8803,N_7940,N_7467);
nand U8804 (N_8804,N_7310,N_7175);
nand U8805 (N_8805,N_7389,N_7734);
xnor U8806 (N_8806,N_7888,N_7564);
and U8807 (N_8807,N_7789,N_7453);
nand U8808 (N_8808,N_7483,N_7965);
or U8809 (N_8809,N_7158,N_7884);
nor U8810 (N_8810,N_7359,N_7886);
nand U8811 (N_8811,N_7532,N_7755);
and U8812 (N_8812,N_7139,N_7083);
nor U8813 (N_8813,N_7341,N_7534);
or U8814 (N_8814,N_7354,N_7578);
and U8815 (N_8815,N_7633,N_7189);
and U8816 (N_8816,N_7361,N_7074);
nand U8817 (N_8817,N_7608,N_7830);
and U8818 (N_8818,N_7138,N_7406);
and U8819 (N_8819,N_7334,N_7485);
or U8820 (N_8820,N_7736,N_7262);
and U8821 (N_8821,N_7437,N_7556);
nand U8822 (N_8822,N_7793,N_7762);
nand U8823 (N_8823,N_7264,N_7121);
nor U8824 (N_8824,N_7656,N_7377);
nand U8825 (N_8825,N_7475,N_7913);
or U8826 (N_8826,N_7578,N_7161);
or U8827 (N_8827,N_7425,N_7308);
nand U8828 (N_8828,N_7989,N_7243);
nand U8829 (N_8829,N_7163,N_7600);
and U8830 (N_8830,N_7633,N_7844);
or U8831 (N_8831,N_7948,N_7244);
nor U8832 (N_8832,N_7256,N_7955);
nor U8833 (N_8833,N_7687,N_7137);
or U8834 (N_8834,N_7860,N_7235);
and U8835 (N_8835,N_7256,N_7383);
and U8836 (N_8836,N_7244,N_7083);
nand U8837 (N_8837,N_7342,N_7383);
and U8838 (N_8838,N_7444,N_7062);
or U8839 (N_8839,N_7232,N_7303);
nor U8840 (N_8840,N_7371,N_7026);
nor U8841 (N_8841,N_7002,N_7020);
and U8842 (N_8842,N_7740,N_7461);
or U8843 (N_8843,N_7543,N_7178);
nor U8844 (N_8844,N_7096,N_7749);
or U8845 (N_8845,N_7552,N_7542);
nor U8846 (N_8846,N_7182,N_7055);
nand U8847 (N_8847,N_7592,N_7018);
or U8848 (N_8848,N_7577,N_7921);
or U8849 (N_8849,N_7973,N_7390);
nor U8850 (N_8850,N_7144,N_7600);
and U8851 (N_8851,N_7748,N_7219);
nor U8852 (N_8852,N_7404,N_7059);
or U8853 (N_8853,N_7677,N_7081);
or U8854 (N_8854,N_7791,N_7817);
and U8855 (N_8855,N_7916,N_7820);
or U8856 (N_8856,N_7658,N_7880);
and U8857 (N_8857,N_7850,N_7525);
and U8858 (N_8858,N_7428,N_7504);
or U8859 (N_8859,N_7414,N_7074);
nand U8860 (N_8860,N_7689,N_7256);
and U8861 (N_8861,N_7985,N_7725);
or U8862 (N_8862,N_7638,N_7488);
and U8863 (N_8863,N_7023,N_7478);
and U8864 (N_8864,N_7852,N_7583);
nand U8865 (N_8865,N_7611,N_7714);
nor U8866 (N_8866,N_7208,N_7895);
nand U8867 (N_8867,N_7163,N_7919);
or U8868 (N_8868,N_7757,N_7262);
nor U8869 (N_8869,N_7042,N_7257);
nand U8870 (N_8870,N_7186,N_7410);
nand U8871 (N_8871,N_7513,N_7995);
or U8872 (N_8872,N_7269,N_7613);
nand U8873 (N_8873,N_7452,N_7333);
nand U8874 (N_8874,N_7718,N_7900);
and U8875 (N_8875,N_7200,N_7464);
nand U8876 (N_8876,N_7085,N_7058);
or U8877 (N_8877,N_7778,N_7662);
nand U8878 (N_8878,N_7645,N_7426);
or U8879 (N_8879,N_7482,N_7036);
and U8880 (N_8880,N_7746,N_7078);
nand U8881 (N_8881,N_7208,N_7030);
or U8882 (N_8882,N_7250,N_7081);
or U8883 (N_8883,N_7656,N_7806);
or U8884 (N_8884,N_7264,N_7220);
or U8885 (N_8885,N_7465,N_7298);
nand U8886 (N_8886,N_7699,N_7191);
nor U8887 (N_8887,N_7607,N_7320);
or U8888 (N_8888,N_7592,N_7854);
and U8889 (N_8889,N_7149,N_7878);
or U8890 (N_8890,N_7199,N_7821);
or U8891 (N_8891,N_7170,N_7407);
or U8892 (N_8892,N_7296,N_7034);
nor U8893 (N_8893,N_7449,N_7466);
nand U8894 (N_8894,N_7603,N_7333);
and U8895 (N_8895,N_7177,N_7903);
or U8896 (N_8896,N_7531,N_7267);
nand U8897 (N_8897,N_7426,N_7705);
nor U8898 (N_8898,N_7263,N_7998);
nor U8899 (N_8899,N_7674,N_7758);
and U8900 (N_8900,N_7772,N_7323);
nor U8901 (N_8901,N_7957,N_7005);
or U8902 (N_8902,N_7675,N_7969);
and U8903 (N_8903,N_7250,N_7915);
and U8904 (N_8904,N_7584,N_7908);
and U8905 (N_8905,N_7377,N_7220);
nand U8906 (N_8906,N_7474,N_7388);
and U8907 (N_8907,N_7387,N_7328);
nor U8908 (N_8908,N_7556,N_7801);
or U8909 (N_8909,N_7529,N_7685);
nor U8910 (N_8910,N_7509,N_7971);
and U8911 (N_8911,N_7003,N_7751);
nand U8912 (N_8912,N_7535,N_7893);
or U8913 (N_8913,N_7239,N_7461);
or U8914 (N_8914,N_7711,N_7405);
and U8915 (N_8915,N_7520,N_7345);
or U8916 (N_8916,N_7732,N_7044);
or U8917 (N_8917,N_7792,N_7311);
or U8918 (N_8918,N_7561,N_7028);
nor U8919 (N_8919,N_7274,N_7677);
or U8920 (N_8920,N_7280,N_7809);
nand U8921 (N_8921,N_7130,N_7602);
and U8922 (N_8922,N_7806,N_7176);
nor U8923 (N_8923,N_7921,N_7533);
nor U8924 (N_8924,N_7940,N_7389);
or U8925 (N_8925,N_7850,N_7875);
nor U8926 (N_8926,N_7189,N_7780);
and U8927 (N_8927,N_7652,N_7849);
or U8928 (N_8928,N_7874,N_7151);
and U8929 (N_8929,N_7932,N_7255);
nor U8930 (N_8930,N_7150,N_7165);
nand U8931 (N_8931,N_7067,N_7836);
and U8932 (N_8932,N_7096,N_7769);
nand U8933 (N_8933,N_7215,N_7265);
nor U8934 (N_8934,N_7508,N_7090);
and U8935 (N_8935,N_7996,N_7763);
nand U8936 (N_8936,N_7888,N_7702);
nand U8937 (N_8937,N_7244,N_7341);
nand U8938 (N_8938,N_7309,N_7312);
or U8939 (N_8939,N_7596,N_7794);
and U8940 (N_8940,N_7977,N_7679);
xor U8941 (N_8941,N_7107,N_7413);
and U8942 (N_8942,N_7090,N_7078);
and U8943 (N_8943,N_7100,N_7898);
nand U8944 (N_8944,N_7191,N_7042);
nand U8945 (N_8945,N_7188,N_7243);
nor U8946 (N_8946,N_7526,N_7983);
or U8947 (N_8947,N_7052,N_7915);
or U8948 (N_8948,N_7344,N_7302);
nand U8949 (N_8949,N_7010,N_7877);
or U8950 (N_8950,N_7787,N_7054);
and U8951 (N_8951,N_7797,N_7459);
nor U8952 (N_8952,N_7522,N_7361);
and U8953 (N_8953,N_7191,N_7858);
nand U8954 (N_8954,N_7997,N_7664);
nor U8955 (N_8955,N_7108,N_7996);
nor U8956 (N_8956,N_7792,N_7935);
and U8957 (N_8957,N_7097,N_7334);
nor U8958 (N_8958,N_7615,N_7363);
nor U8959 (N_8959,N_7150,N_7405);
or U8960 (N_8960,N_7458,N_7868);
nor U8961 (N_8961,N_7757,N_7637);
or U8962 (N_8962,N_7391,N_7037);
and U8963 (N_8963,N_7137,N_7795);
and U8964 (N_8964,N_7311,N_7139);
nand U8965 (N_8965,N_7227,N_7723);
or U8966 (N_8966,N_7386,N_7366);
nand U8967 (N_8967,N_7302,N_7341);
or U8968 (N_8968,N_7682,N_7535);
or U8969 (N_8969,N_7305,N_7190);
nor U8970 (N_8970,N_7144,N_7577);
and U8971 (N_8971,N_7378,N_7709);
and U8972 (N_8972,N_7120,N_7107);
and U8973 (N_8973,N_7238,N_7589);
and U8974 (N_8974,N_7883,N_7249);
and U8975 (N_8975,N_7728,N_7746);
nor U8976 (N_8976,N_7291,N_7173);
or U8977 (N_8977,N_7873,N_7835);
nor U8978 (N_8978,N_7142,N_7800);
or U8979 (N_8979,N_7672,N_7390);
nand U8980 (N_8980,N_7710,N_7441);
or U8981 (N_8981,N_7687,N_7249);
or U8982 (N_8982,N_7115,N_7582);
or U8983 (N_8983,N_7856,N_7991);
nand U8984 (N_8984,N_7412,N_7373);
and U8985 (N_8985,N_7785,N_7424);
nor U8986 (N_8986,N_7668,N_7464);
nand U8987 (N_8987,N_7206,N_7406);
or U8988 (N_8988,N_7269,N_7457);
or U8989 (N_8989,N_7998,N_7830);
and U8990 (N_8990,N_7225,N_7373);
and U8991 (N_8991,N_7182,N_7845);
and U8992 (N_8992,N_7507,N_7041);
nand U8993 (N_8993,N_7209,N_7999);
nand U8994 (N_8994,N_7991,N_7101);
nand U8995 (N_8995,N_7745,N_7934);
and U8996 (N_8996,N_7644,N_7537);
nor U8997 (N_8997,N_7940,N_7432);
nand U8998 (N_8998,N_7862,N_7839);
and U8999 (N_8999,N_7467,N_7119);
and U9000 (N_9000,N_8114,N_8978);
or U9001 (N_9001,N_8753,N_8318);
nand U9002 (N_9002,N_8795,N_8980);
and U9003 (N_9003,N_8561,N_8793);
or U9004 (N_9004,N_8000,N_8189);
and U9005 (N_9005,N_8348,N_8226);
or U9006 (N_9006,N_8073,N_8860);
or U9007 (N_9007,N_8542,N_8733);
nor U9008 (N_9008,N_8258,N_8293);
nor U9009 (N_9009,N_8620,N_8074);
nor U9010 (N_9010,N_8387,N_8842);
nor U9011 (N_9011,N_8922,N_8637);
and U9012 (N_9012,N_8631,N_8392);
nand U9013 (N_9013,N_8076,N_8791);
or U9014 (N_9014,N_8736,N_8004);
and U9015 (N_9015,N_8589,N_8823);
and U9016 (N_9016,N_8035,N_8916);
or U9017 (N_9017,N_8200,N_8996);
nor U9018 (N_9018,N_8085,N_8810);
nand U9019 (N_9019,N_8523,N_8134);
or U9020 (N_9020,N_8500,N_8877);
or U9021 (N_9021,N_8297,N_8895);
and U9022 (N_9022,N_8368,N_8956);
nand U9023 (N_9023,N_8011,N_8636);
nor U9024 (N_9024,N_8016,N_8448);
nor U9025 (N_9025,N_8694,N_8121);
or U9026 (N_9026,N_8755,N_8147);
nand U9027 (N_9027,N_8816,N_8477);
or U9028 (N_9028,N_8682,N_8516);
and U9029 (N_9029,N_8774,N_8760);
nand U9030 (N_9030,N_8543,N_8897);
and U9031 (N_9031,N_8855,N_8556);
and U9032 (N_9032,N_8170,N_8867);
nand U9033 (N_9033,N_8946,N_8140);
nand U9034 (N_9034,N_8399,N_8827);
or U9035 (N_9035,N_8115,N_8580);
nor U9036 (N_9036,N_8982,N_8030);
or U9037 (N_9037,N_8447,N_8741);
and U9038 (N_9038,N_8811,N_8782);
and U9039 (N_9039,N_8911,N_8410);
nor U9040 (N_9040,N_8369,N_8779);
and U9041 (N_9041,N_8290,N_8781);
and U9042 (N_9042,N_8272,N_8048);
or U9043 (N_9043,N_8175,N_8906);
or U9044 (N_9044,N_8717,N_8788);
or U9045 (N_9045,N_8110,N_8427);
or U9046 (N_9046,N_8798,N_8449);
and U9047 (N_9047,N_8057,N_8645);
nand U9048 (N_9048,N_8202,N_8591);
and U9049 (N_9049,N_8187,N_8949);
nor U9050 (N_9050,N_8541,N_8100);
and U9051 (N_9051,N_8910,N_8098);
nor U9052 (N_9052,N_8773,N_8455);
and U9053 (N_9053,N_8245,N_8193);
or U9054 (N_9054,N_8548,N_8436);
or U9055 (N_9055,N_8767,N_8721);
and U9056 (N_9056,N_8322,N_8987);
nand U9057 (N_9057,N_8619,N_8931);
or U9058 (N_9058,N_8353,N_8787);
or U9059 (N_9059,N_8994,N_8878);
or U9060 (N_9060,N_8233,N_8285);
or U9061 (N_9061,N_8444,N_8567);
nand U9062 (N_9062,N_8959,N_8920);
nand U9063 (N_9063,N_8428,N_8169);
nor U9064 (N_9064,N_8903,N_8466);
and U9065 (N_9065,N_8754,N_8406);
and U9066 (N_9066,N_8805,N_8157);
and U9067 (N_9067,N_8985,N_8062);
nor U9068 (N_9068,N_8735,N_8087);
nand U9069 (N_9069,N_8845,N_8874);
nand U9070 (N_9070,N_8283,N_8067);
nor U9071 (N_9071,N_8314,N_8598);
nor U9072 (N_9072,N_8102,N_8613);
nand U9073 (N_9073,N_8858,N_8416);
or U9074 (N_9074,N_8995,N_8396);
and U9075 (N_9075,N_8021,N_8208);
nor U9076 (N_9076,N_8780,N_8264);
or U9077 (N_9077,N_8586,N_8834);
or U9078 (N_9078,N_8966,N_8199);
nor U9079 (N_9079,N_8653,N_8148);
or U9080 (N_9080,N_8853,N_8641);
nor U9081 (N_9081,N_8190,N_8109);
nand U9082 (N_9082,N_8316,N_8622);
and U9083 (N_9083,N_8677,N_8330);
nand U9084 (N_9084,N_8808,N_8332);
and U9085 (N_9085,N_8761,N_8521);
nor U9086 (N_9086,N_8326,N_8469);
or U9087 (N_9087,N_8219,N_8043);
nor U9088 (N_9088,N_8390,N_8618);
nand U9089 (N_9089,N_8594,N_8889);
nand U9090 (N_9090,N_8703,N_8128);
nor U9091 (N_9091,N_8388,N_8433);
nor U9092 (N_9092,N_8441,N_8470);
nor U9093 (N_9093,N_8003,N_8431);
nand U9094 (N_9094,N_8010,N_8551);
nand U9095 (N_9095,N_8349,N_8864);
or U9096 (N_9096,N_8592,N_8487);
nor U9097 (N_9097,N_8304,N_8132);
and U9098 (N_9098,N_8524,N_8090);
and U9099 (N_9099,N_8565,N_8749);
or U9100 (N_9100,N_8014,N_8738);
and U9101 (N_9101,N_8601,N_8674);
nand U9102 (N_9102,N_8558,N_8796);
or U9103 (N_9103,N_8496,N_8023);
nand U9104 (N_9104,N_8154,N_8092);
or U9105 (N_9105,N_8711,N_8149);
and U9106 (N_9106,N_8254,N_8731);
nand U9107 (N_9107,N_8778,N_8400);
or U9108 (N_9108,N_8282,N_8244);
or U9109 (N_9109,N_8381,N_8847);
and U9110 (N_9110,N_8861,N_8953);
and U9111 (N_9111,N_8331,N_8686);
and U9112 (N_9112,N_8667,N_8403);
nor U9113 (N_9113,N_8367,N_8344);
nand U9114 (N_9114,N_8958,N_8859);
or U9115 (N_9115,N_8902,N_8530);
nand U9116 (N_9116,N_8484,N_8358);
nor U9117 (N_9117,N_8955,N_8256);
or U9118 (N_9118,N_8405,N_8361);
nor U9119 (N_9119,N_8497,N_8585);
nor U9120 (N_9120,N_8588,N_8270);
nand U9121 (N_9121,N_8746,N_8950);
and U9122 (N_9122,N_8952,N_8714);
or U9123 (N_9123,N_8882,N_8616);
nor U9124 (N_9124,N_8355,N_8395);
nand U9125 (N_9125,N_8311,N_8183);
and U9126 (N_9126,N_8380,N_8777);
nand U9127 (N_9127,N_8207,N_8852);
or U9128 (N_9128,N_8770,N_8826);
and U9129 (N_9129,N_8309,N_8573);
nand U9130 (N_9130,N_8172,N_8655);
nor U9131 (N_9131,N_8243,N_8513);
nor U9132 (N_9132,N_8769,N_8841);
nand U9133 (N_9133,N_8634,N_8607);
nor U9134 (N_9134,N_8462,N_8130);
nand U9135 (N_9135,N_8156,N_8943);
or U9136 (N_9136,N_8532,N_8206);
or U9137 (N_9137,N_8216,N_8701);
and U9138 (N_9138,N_8918,N_8514);
and U9139 (N_9139,N_8739,N_8537);
and U9140 (N_9140,N_8710,N_8397);
nor U9141 (N_9141,N_8101,N_8215);
nand U9142 (N_9142,N_8732,N_8263);
or U9143 (N_9143,N_8800,N_8596);
nand U9144 (N_9144,N_8070,N_8357);
and U9145 (N_9145,N_8450,N_8893);
nor U9146 (N_9146,N_8471,N_8602);
nand U9147 (N_9147,N_8376,N_8512);
and U9148 (N_9148,N_8040,N_8197);
nor U9149 (N_9149,N_8255,N_8231);
nor U9150 (N_9150,N_8609,N_8482);
nand U9151 (N_9151,N_8338,N_8941);
or U9152 (N_9152,N_8784,N_8252);
nand U9153 (N_9153,N_8965,N_8693);
nand U9154 (N_9154,N_8923,N_8993);
and U9155 (N_9155,N_8209,N_8006);
nor U9156 (N_9156,N_8974,N_8454);
and U9157 (N_9157,N_8547,N_8865);
nand U9158 (N_9158,N_8574,N_8518);
or U9159 (N_9159,N_8086,N_8379);
and U9160 (N_9160,N_8196,N_8107);
or U9161 (N_9161,N_8302,N_8179);
or U9162 (N_9162,N_8013,N_8099);
or U9163 (N_9163,N_8989,N_8564);
and U9164 (N_9164,N_8813,N_8480);
nand U9165 (N_9165,N_8743,N_8072);
or U9166 (N_9166,N_8398,N_8772);
nand U9167 (N_9167,N_8075,N_8069);
nor U9168 (N_9168,N_8323,N_8061);
or U9169 (N_9169,N_8205,N_8663);
nand U9170 (N_9170,N_8894,N_8123);
nand U9171 (N_9171,N_8881,N_8786);
nand U9172 (N_9172,N_8198,N_8578);
nand U9173 (N_9173,N_8131,N_8650);
and U9174 (N_9174,N_8942,N_8135);
nor U9175 (N_9175,N_8563,N_8643);
nand U9176 (N_9176,N_8463,N_8539);
or U9177 (N_9177,N_8790,N_8136);
nand U9178 (N_9178,N_8127,N_8981);
and U9179 (N_9179,N_8590,N_8756);
and U9180 (N_9180,N_8167,N_8235);
xnor U9181 (N_9181,N_8583,N_8873);
and U9182 (N_9182,N_8153,N_8232);
nand U9183 (N_9183,N_8915,N_8673);
or U9184 (N_9184,N_8220,N_8194);
nand U9185 (N_9185,N_8697,N_8624);
nand U9186 (N_9186,N_8654,N_8005);
and U9187 (N_9187,N_8051,N_8990);
or U9188 (N_9188,N_8414,N_8105);
nand U9189 (N_9189,N_8831,N_8527);
and U9190 (N_9190,N_8476,N_8844);
and U9191 (N_9191,N_8928,N_8522);
nand U9192 (N_9192,N_8181,N_8825);
and U9193 (N_9193,N_8820,N_8045);
or U9194 (N_9194,N_8579,N_8164);
and U9195 (N_9195,N_8603,N_8288);
nor U9196 (N_9196,N_8230,N_8875);
nand U9197 (N_9197,N_8716,N_8015);
and U9198 (N_9198,N_8507,N_8247);
nor U9199 (N_9199,N_8992,N_8765);
and U9200 (N_9200,N_8327,N_8412);
and U9201 (N_9201,N_8423,N_8939);
and U9202 (N_9202,N_8120,N_8064);
and U9203 (N_9203,N_8708,N_8227);
and U9204 (N_9204,N_8824,N_8821);
and U9205 (N_9205,N_8896,N_8696);
nand U9206 (N_9206,N_8520,N_8529);
or U9207 (N_9207,N_8575,N_8660);
or U9208 (N_9208,N_8662,N_8934);
nor U9209 (N_9209,N_8659,N_8913);
nand U9210 (N_9210,N_8486,N_8020);
or U9211 (N_9211,N_8386,N_8017);
nor U9212 (N_9212,N_8600,N_8287);
or U9213 (N_9213,N_8335,N_8041);
nor U9214 (N_9214,N_8633,N_8037);
xor U9215 (N_9215,N_8666,N_8550);
nor U9216 (N_9216,N_8528,N_8722);
or U9217 (N_9217,N_8345,N_8028);
nor U9218 (N_9218,N_8509,N_8248);
and U9219 (N_9219,N_8999,N_8933);
nor U9220 (N_9220,N_8737,N_8748);
nor U9221 (N_9221,N_8126,N_8569);
and U9222 (N_9222,N_8411,N_8321);
nand U9223 (N_9223,N_8740,N_8088);
nor U9224 (N_9224,N_8060,N_8310);
or U9225 (N_9225,N_8690,N_8122);
and U9226 (N_9226,N_8623,N_8803);
or U9227 (N_9227,N_8242,N_8036);
nand U9228 (N_9228,N_8689,N_8262);
or U9229 (N_9229,N_8108,N_8174);
or U9230 (N_9230,N_8794,N_8246);
nand U9231 (N_9231,N_8295,N_8239);
xnor U9232 (N_9232,N_8445,N_8453);
nor U9233 (N_9233,N_8425,N_8642);
and U9234 (N_9234,N_8300,N_8026);
nand U9235 (N_9235,N_8320,N_8472);
or U9236 (N_9236,N_8728,N_8336);
nor U9237 (N_9237,N_8033,N_8328);
nor U9238 (N_9238,N_8143,N_8888);
or U9239 (N_9239,N_8401,N_8176);
nand U9240 (N_9240,N_8342,N_8203);
nor U9241 (N_9241,N_8912,N_8201);
or U9242 (N_9242,N_8555,N_8764);
nand U9243 (N_9243,N_8862,N_8250);
nand U9244 (N_9244,N_8751,N_8566);
nor U9245 (N_9245,N_8267,N_8094);
and U9246 (N_9246,N_8251,N_8757);
nor U9247 (N_9247,N_8467,N_8341);
and U9248 (N_9248,N_8534,N_8079);
nor U9249 (N_9249,N_8807,N_8475);
or U9250 (N_9250,N_8442,N_8935);
and U9251 (N_9251,N_8621,N_8649);
or U9252 (N_9252,N_8229,N_8526);
and U9253 (N_9253,N_8812,N_8818);
nor U9254 (N_9254,N_8093,N_8365);
and U9255 (N_9255,N_8763,N_8370);
or U9256 (N_9256,N_8511,N_8052);
or U9257 (N_9257,N_8658,N_8138);
nor U9258 (N_9258,N_8426,N_8917);
nand U9259 (N_9259,N_8678,N_8402);
nor U9260 (N_9260,N_8253,N_8927);
or U9261 (N_9261,N_8829,N_8281);
and U9262 (N_9262,N_8907,N_8439);
nand U9263 (N_9263,N_8880,N_8819);
nor U9264 (N_9264,N_8744,N_8479);
nand U9265 (N_9265,N_8089,N_8571);
nand U9266 (N_9266,N_8970,N_8277);
and U9267 (N_9267,N_8891,N_8605);
or U9268 (N_9268,N_8452,N_8651);
nor U9269 (N_9269,N_8544,N_8625);
nor U9270 (N_9270,N_8814,N_8635);
nand U9271 (N_9271,N_8413,N_8404);
and U9272 (N_9272,N_8078,N_8315);
or U9273 (N_9273,N_8991,N_8599);
or U9274 (N_9274,N_8068,N_8192);
nand U9275 (N_9275,N_8593,N_8485);
nand U9276 (N_9276,N_8185,N_8887);
nor U9277 (N_9277,N_8418,N_8804);
nand U9278 (N_9278,N_8675,N_8681);
nor U9279 (N_9279,N_8615,N_8223);
or U9280 (N_9280,N_8065,N_8626);
nand U9281 (N_9281,N_8885,N_8266);
nand U9282 (N_9282,N_8166,N_8019);
and U9283 (N_9283,N_8799,N_8071);
nor U9284 (N_9284,N_8630,N_8776);
nand U9285 (N_9285,N_8871,N_8178);
nor U9286 (N_9286,N_8611,N_8545);
xnor U9287 (N_9287,N_8298,N_8260);
and U9288 (N_9288,N_8604,N_8726);
and U9289 (N_9289,N_8382,N_8560);
nand U9290 (N_9290,N_8919,N_8313);
nand U9291 (N_9291,N_8464,N_8727);
nand U9292 (N_9292,N_8142,N_8025);
nor U9293 (N_9293,N_8775,N_8458);
or U9294 (N_9294,N_8173,N_8945);
or U9295 (N_9295,N_8184,N_8032);
and U9296 (N_9296,N_8222,N_8113);
xnor U9297 (N_9297,N_8366,N_8840);
or U9298 (N_9298,N_8280,N_8271);
or U9299 (N_9299,N_8951,N_8116);
nor U9300 (N_9300,N_8683,N_8967);
and U9301 (N_9301,N_8329,N_8627);
nor U9302 (N_9302,N_8533,N_8312);
nand U9303 (N_9303,N_8211,N_8119);
nor U9304 (N_9304,N_8077,N_8163);
or U9305 (N_9305,N_8237,N_8461);
or U9306 (N_9306,N_8286,N_8608);
and U9307 (N_9307,N_8284,N_8553);
nor U9308 (N_9308,N_8289,N_8162);
or U9309 (N_9309,N_8771,N_8238);
or U9310 (N_9310,N_8224,N_8870);
or U9311 (N_9311,N_8815,N_8047);
and U9312 (N_9312,N_8212,N_8789);
or U9313 (N_9313,N_8901,N_8639);
or U9314 (N_9314,N_8718,N_8656);
nand U9315 (N_9315,N_8671,N_8117);
and U9316 (N_9316,N_8360,N_8519);
nand U9317 (N_9317,N_8712,N_8009);
and U9318 (N_9318,N_8698,N_8325);
nand U9319 (N_9319,N_8940,N_8279);
nand U9320 (N_9320,N_8986,N_8837);
or U9321 (N_9321,N_8540,N_8435);
or U9322 (N_9322,N_8408,N_8930);
or U9323 (N_9323,N_8095,N_8407);
nor U9324 (N_9324,N_8876,N_8029);
nand U9325 (N_9325,N_8221,N_8747);
nand U9326 (N_9326,N_8356,N_8056);
or U9327 (N_9327,N_8661,N_8278);
nand U9328 (N_9328,N_8988,N_8129);
or U9329 (N_9329,N_8339,N_8856);
nand U9330 (N_9330,N_8457,N_8493);
nor U9331 (N_9331,N_8872,N_8848);
nor U9332 (N_9332,N_8165,N_8024);
and U9333 (N_9333,N_8680,N_8758);
and U9334 (N_9334,N_8228,N_8261);
and U9335 (N_9335,N_8415,N_8139);
or U9336 (N_9336,N_8091,N_8350);
nand U9337 (N_9337,N_8490,N_8617);
and U9338 (N_9338,N_8505,N_8160);
nor U9339 (N_9339,N_8857,N_8954);
nand U9340 (N_9340,N_8393,N_8745);
or U9341 (N_9341,N_8707,N_8692);
or U9342 (N_9342,N_8039,N_8042);
and U9343 (N_9343,N_8843,N_8614);
and U9344 (N_9344,N_8451,N_8421);
and U9345 (N_9345,N_8141,N_8879);
and U9346 (N_9346,N_8587,N_8979);
or U9347 (N_9347,N_8234,N_8801);
nor U9348 (N_9348,N_8424,N_8063);
and U9349 (N_9349,N_8557,N_8146);
and U9350 (N_9350,N_8822,N_8299);
nand U9351 (N_9351,N_8863,N_8351);
nor U9352 (N_9352,N_8050,N_8515);
nand U9353 (N_9353,N_8525,N_8629);
and U9354 (N_9354,N_8171,N_8151);
and U9355 (N_9355,N_8577,N_8306);
nor U9356 (N_9356,N_8438,N_8417);
nand U9357 (N_9357,N_8506,N_8976);
or U9358 (N_9358,N_8002,N_8670);
nand U9359 (N_9359,N_8503,N_8374);
and U9360 (N_9360,N_8549,N_8730);
and U9361 (N_9361,N_8640,N_8066);
nand U9362 (N_9362,N_8495,N_8652);
nand U9363 (N_9363,N_8430,N_8275);
nand U9364 (N_9364,N_8898,N_8054);
or U9365 (N_9365,N_8606,N_8492);
nand U9366 (N_9366,N_8612,N_8582);
nor U9367 (N_9367,N_8576,N_8983);
or U9368 (N_9368,N_8854,N_8481);
nor U9369 (N_9369,N_8685,N_8383);
nand U9370 (N_9370,N_8968,N_8308);
nor U9371 (N_9371,N_8468,N_8610);
nor U9372 (N_9372,N_8572,N_8429);
nor U9373 (N_9373,N_8925,N_8676);
nor U9374 (N_9374,N_8699,N_8762);
and U9375 (N_9375,N_8038,N_8489);
nor U9376 (N_9376,N_8937,N_8538);
or U9377 (N_9377,N_8103,N_8504);
nor U9378 (N_9378,N_8268,N_8097);
nor U9379 (N_9379,N_8473,N_8352);
or U9380 (N_9380,N_8155,N_8723);
nand U9381 (N_9381,N_8904,N_8301);
or U9382 (N_9382,N_8494,N_8783);
and U9383 (N_9383,N_8672,N_8241);
nand U9384 (N_9384,N_8111,N_8307);
nand U9385 (N_9385,N_8971,N_8502);
and U9386 (N_9386,N_8044,N_8715);
xnor U9387 (N_9387,N_8446,N_8719);
nor U9388 (N_9388,N_8018,N_8150);
nor U9389 (N_9389,N_8665,N_8535);
nand U9390 (N_9390,N_8836,N_8646);
nand U9391 (N_9391,N_8001,N_8944);
and U9392 (N_9392,N_8145,N_8276);
or U9393 (N_9393,N_8570,N_8962);
or U9394 (N_9394,N_8975,N_8884);
nand U9395 (N_9395,N_8213,N_8552);
and U9396 (N_9396,N_8456,N_8768);
nand U9397 (N_9397,N_8240,N_8081);
nor U9398 (N_9398,N_8972,N_8084);
or U9399 (N_9399,N_8249,N_8998);
nand U9400 (N_9400,N_8724,N_8378);
and U9401 (N_9401,N_8055,N_8459);
nor U9402 (N_9402,N_8317,N_8568);
or U9403 (N_9403,N_8647,N_8936);
and U9404 (N_9404,N_8914,N_8225);
nand U9405 (N_9405,N_8296,N_8188);
nor U9406 (N_9406,N_8319,N_8562);
and U9407 (N_9407,N_8218,N_8832);
and U9408 (N_9408,N_8359,N_8343);
or U9409 (N_9409,N_8501,N_8409);
nor U9410 (N_9410,N_8385,N_8363);
nand U9411 (N_9411,N_8394,N_8833);
or U9412 (N_9412,N_8182,N_8759);
or U9413 (N_9413,N_8498,N_8691);
nand U9414 (N_9414,N_8706,N_8303);
nor U9415 (N_9415,N_8177,N_8908);
nand U9416 (N_9416,N_8973,N_8729);
or U9417 (N_9417,N_8269,N_8734);
or U9418 (N_9418,N_8362,N_8008);
nand U9419 (N_9419,N_8305,N_8389);
and U9420 (N_9420,N_8273,N_8977);
nor U9421 (N_9421,N_8419,N_8460);
nand U9422 (N_9422,N_8096,N_8644);
nor U9423 (N_9423,N_8713,N_8802);
or U9424 (N_9424,N_8892,N_8900);
and U9425 (N_9425,N_8488,N_8124);
nand U9426 (N_9426,N_8905,N_8478);
or U9427 (N_9427,N_8371,N_8702);
nand U9428 (N_9428,N_8932,N_8082);
nand U9429 (N_9429,N_8375,N_8809);
or U9430 (N_9430,N_8373,N_8684);
nand U9431 (N_9431,N_8866,N_8559);
nand U9432 (N_9432,N_8688,N_8053);
nor U9433 (N_9433,N_8391,N_8112);
nor U9434 (N_9434,N_8725,N_8118);
and U9435 (N_9435,N_8628,N_8664);
or U9436 (N_9436,N_8420,N_8909);
nor U9437 (N_9437,N_8938,N_8947);
nand U9438 (N_9438,N_8687,N_8929);
or U9439 (N_9439,N_8531,N_8274);
nor U9440 (N_9440,N_8957,N_8080);
nand U9441 (N_9441,N_8963,N_8546);
nand U9442 (N_9442,N_8839,N_8186);
or U9443 (N_9443,N_8027,N_8752);
or U9444 (N_9444,N_8483,N_8106);
nor U9445 (N_9445,N_8152,N_8828);
nor U9446 (N_9446,N_8869,N_8632);
or U9447 (N_9447,N_8536,N_8432);
nand U9448 (N_9448,N_8334,N_8850);
nand U9449 (N_9449,N_8668,N_8750);
nor U9450 (N_9450,N_8554,N_8742);
or U9451 (N_9451,N_8034,N_8584);
and U9452 (N_9452,N_8333,N_8049);
nor U9453 (N_9453,N_8257,N_8785);
nand U9454 (N_9454,N_8797,N_8377);
or U9455 (N_9455,N_8437,N_8434);
and U9456 (N_9456,N_8059,N_8104);
and U9457 (N_9457,N_8265,N_8517);
or U9458 (N_9458,N_8294,N_8846);
nor U9459 (N_9459,N_8886,N_8161);
and U9460 (N_9460,N_8158,N_8669);
and U9461 (N_9461,N_8499,N_8384);
and U9462 (N_9462,N_8926,N_8291);
or U9463 (N_9463,N_8838,N_8058);
and U9464 (N_9464,N_8948,N_8210);
or U9465 (N_9465,N_8443,N_8491);
and U9466 (N_9466,N_8679,N_8595);
nor U9467 (N_9467,N_8214,N_8806);
or U9468 (N_9468,N_8657,N_8372);
nand U9469 (N_9469,N_8997,N_8191);
nand U9470 (N_9470,N_8031,N_8851);
nor U9471 (N_9471,N_8899,N_8259);
or U9472 (N_9472,N_8921,N_8964);
or U9473 (N_9473,N_8695,N_8597);
nand U9474 (N_9474,N_8354,N_8709);
or U9475 (N_9475,N_8883,N_8581);
and U9476 (N_9476,N_8022,N_8465);
xor U9477 (N_9477,N_8340,N_8422);
nand U9478 (N_9478,N_8924,N_8144);
nor U9479 (N_9479,N_8217,N_8180);
nor U9480 (N_9480,N_8440,N_8648);
nor U9481 (N_9481,N_8292,N_8337);
or U9482 (N_9482,N_8849,N_8766);
and U9483 (N_9483,N_8638,N_8984);
and U9484 (N_9484,N_8830,N_8720);
or U9485 (N_9485,N_8347,N_8868);
and U9486 (N_9486,N_8137,N_8324);
or U9487 (N_9487,N_8969,N_8364);
or U9488 (N_9488,N_8792,N_8236);
or U9489 (N_9489,N_8083,N_8510);
or U9490 (N_9490,N_8346,N_8704);
and U9491 (N_9491,N_8133,N_8817);
or U9492 (N_9492,N_8835,N_8700);
and U9493 (N_9493,N_8046,N_8890);
and U9494 (N_9494,N_8195,N_8474);
nand U9495 (N_9495,N_8012,N_8961);
and U9496 (N_9496,N_8508,N_8125);
and U9497 (N_9497,N_8705,N_8007);
or U9498 (N_9498,N_8960,N_8159);
and U9499 (N_9499,N_8168,N_8204);
and U9500 (N_9500,N_8665,N_8069);
or U9501 (N_9501,N_8600,N_8295);
nor U9502 (N_9502,N_8190,N_8381);
and U9503 (N_9503,N_8092,N_8258);
or U9504 (N_9504,N_8909,N_8143);
and U9505 (N_9505,N_8531,N_8650);
or U9506 (N_9506,N_8421,N_8616);
or U9507 (N_9507,N_8464,N_8292);
nand U9508 (N_9508,N_8213,N_8136);
or U9509 (N_9509,N_8025,N_8272);
nand U9510 (N_9510,N_8086,N_8113);
nand U9511 (N_9511,N_8816,N_8557);
and U9512 (N_9512,N_8467,N_8879);
nor U9513 (N_9513,N_8666,N_8522);
nand U9514 (N_9514,N_8121,N_8104);
or U9515 (N_9515,N_8300,N_8070);
nor U9516 (N_9516,N_8163,N_8322);
or U9517 (N_9517,N_8999,N_8745);
or U9518 (N_9518,N_8431,N_8740);
nor U9519 (N_9519,N_8310,N_8934);
nand U9520 (N_9520,N_8554,N_8875);
nor U9521 (N_9521,N_8558,N_8624);
and U9522 (N_9522,N_8210,N_8351);
nand U9523 (N_9523,N_8361,N_8611);
or U9524 (N_9524,N_8818,N_8651);
or U9525 (N_9525,N_8779,N_8585);
nand U9526 (N_9526,N_8811,N_8490);
or U9527 (N_9527,N_8371,N_8451);
or U9528 (N_9528,N_8311,N_8989);
nor U9529 (N_9529,N_8881,N_8862);
nor U9530 (N_9530,N_8495,N_8172);
nand U9531 (N_9531,N_8243,N_8482);
nand U9532 (N_9532,N_8722,N_8966);
nor U9533 (N_9533,N_8135,N_8841);
or U9534 (N_9534,N_8242,N_8840);
or U9535 (N_9535,N_8410,N_8192);
xnor U9536 (N_9536,N_8091,N_8671);
nor U9537 (N_9537,N_8616,N_8044);
or U9538 (N_9538,N_8656,N_8304);
nor U9539 (N_9539,N_8870,N_8850);
or U9540 (N_9540,N_8413,N_8771);
or U9541 (N_9541,N_8185,N_8483);
xnor U9542 (N_9542,N_8808,N_8325);
nor U9543 (N_9543,N_8841,N_8878);
nand U9544 (N_9544,N_8764,N_8290);
or U9545 (N_9545,N_8083,N_8301);
and U9546 (N_9546,N_8790,N_8708);
nand U9547 (N_9547,N_8165,N_8153);
or U9548 (N_9548,N_8324,N_8359);
and U9549 (N_9549,N_8219,N_8531);
and U9550 (N_9550,N_8472,N_8018);
nor U9551 (N_9551,N_8264,N_8727);
nor U9552 (N_9552,N_8572,N_8190);
and U9553 (N_9553,N_8998,N_8519);
or U9554 (N_9554,N_8842,N_8361);
nand U9555 (N_9555,N_8545,N_8478);
or U9556 (N_9556,N_8805,N_8491);
or U9557 (N_9557,N_8022,N_8209);
or U9558 (N_9558,N_8309,N_8692);
nor U9559 (N_9559,N_8189,N_8291);
nor U9560 (N_9560,N_8676,N_8017);
or U9561 (N_9561,N_8720,N_8389);
nand U9562 (N_9562,N_8326,N_8325);
nand U9563 (N_9563,N_8824,N_8169);
nand U9564 (N_9564,N_8877,N_8626);
and U9565 (N_9565,N_8636,N_8545);
nor U9566 (N_9566,N_8578,N_8972);
nand U9567 (N_9567,N_8409,N_8367);
nor U9568 (N_9568,N_8707,N_8630);
or U9569 (N_9569,N_8489,N_8855);
and U9570 (N_9570,N_8412,N_8568);
nand U9571 (N_9571,N_8601,N_8711);
xor U9572 (N_9572,N_8588,N_8926);
nor U9573 (N_9573,N_8945,N_8853);
or U9574 (N_9574,N_8413,N_8735);
or U9575 (N_9575,N_8112,N_8687);
nor U9576 (N_9576,N_8615,N_8852);
or U9577 (N_9577,N_8495,N_8733);
nor U9578 (N_9578,N_8049,N_8258);
nor U9579 (N_9579,N_8892,N_8919);
and U9580 (N_9580,N_8041,N_8364);
or U9581 (N_9581,N_8097,N_8075);
nand U9582 (N_9582,N_8556,N_8018);
nand U9583 (N_9583,N_8394,N_8882);
and U9584 (N_9584,N_8405,N_8238);
or U9585 (N_9585,N_8461,N_8663);
nor U9586 (N_9586,N_8350,N_8591);
nor U9587 (N_9587,N_8706,N_8189);
or U9588 (N_9588,N_8210,N_8042);
nand U9589 (N_9589,N_8154,N_8578);
xor U9590 (N_9590,N_8503,N_8364);
nor U9591 (N_9591,N_8826,N_8354);
nand U9592 (N_9592,N_8642,N_8961);
and U9593 (N_9593,N_8133,N_8082);
or U9594 (N_9594,N_8904,N_8251);
nor U9595 (N_9595,N_8671,N_8208);
or U9596 (N_9596,N_8336,N_8668);
or U9597 (N_9597,N_8597,N_8993);
nand U9598 (N_9598,N_8672,N_8351);
and U9599 (N_9599,N_8886,N_8845);
nor U9600 (N_9600,N_8403,N_8802);
and U9601 (N_9601,N_8922,N_8211);
or U9602 (N_9602,N_8154,N_8198);
or U9603 (N_9603,N_8744,N_8149);
nand U9604 (N_9604,N_8693,N_8280);
or U9605 (N_9605,N_8859,N_8657);
and U9606 (N_9606,N_8420,N_8412);
and U9607 (N_9607,N_8195,N_8814);
or U9608 (N_9608,N_8942,N_8511);
nand U9609 (N_9609,N_8471,N_8263);
nor U9610 (N_9610,N_8344,N_8610);
and U9611 (N_9611,N_8961,N_8117);
nand U9612 (N_9612,N_8097,N_8796);
nand U9613 (N_9613,N_8968,N_8982);
nand U9614 (N_9614,N_8286,N_8943);
nand U9615 (N_9615,N_8905,N_8541);
and U9616 (N_9616,N_8991,N_8361);
nor U9617 (N_9617,N_8538,N_8262);
and U9618 (N_9618,N_8462,N_8767);
or U9619 (N_9619,N_8972,N_8534);
nor U9620 (N_9620,N_8259,N_8955);
or U9621 (N_9621,N_8010,N_8045);
or U9622 (N_9622,N_8489,N_8992);
nor U9623 (N_9623,N_8063,N_8787);
nand U9624 (N_9624,N_8086,N_8834);
or U9625 (N_9625,N_8007,N_8232);
nand U9626 (N_9626,N_8143,N_8053);
nand U9627 (N_9627,N_8332,N_8452);
nor U9628 (N_9628,N_8627,N_8365);
and U9629 (N_9629,N_8761,N_8794);
nor U9630 (N_9630,N_8465,N_8425);
nand U9631 (N_9631,N_8566,N_8702);
nor U9632 (N_9632,N_8224,N_8014);
nand U9633 (N_9633,N_8385,N_8626);
nand U9634 (N_9634,N_8525,N_8538);
nor U9635 (N_9635,N_8457,N_8913);
nor U9636 (N_9636,N_8177,N_8877);
nand U9637 (N_9637,N_8045,N_8658);
and U9638 (N_9638,N_8640,N_8069);
or U9639 (N_9639,N_8805,N_8935);
nor U9640 (N_9640,N_8215,N_8061);
or U9641 (N_9641,N_8305,N_8696);
nor U9642 (N_9642,N_8474,N_8664);
and U9643 (N_9643,N_8231,N_8020);
or U9644 (N_9644,N_8453,N_8590);
nor U9645 (N_9645,N_8585,N_8839);
nand U9646 (N_9646,N_8469,N_8973);
and U9647 (N_9647,N_8477,N_8120);
or U9648 (N_9648,N_8545,N_8673);
or U9649 (N_9649,N_8343,N_8888);
nand U9650 (N_9650,N_8435,N_8299);
nand U9651 (N_9651,N_8350,N_8626);
nor U9652 (N_9652,N_8187,N_8806);
nand U9653 (N_9653,N_8399,N_8864);
and U9654 (N_9654,N_8421,N_8397);
nand U9655 (N_9655,N_8679,N_8063);
nand U9656 (N_9656,N_8078,N_8439);
nand U9657 (N_9657,N_8986,N_8948);
nor U9658 (N_9658,N_8590,N_8185);
and U9659 (N_9659,N_8284,N_8671);
and U9660 (N_9660,N_8439,N_8679);
and U9661 (N_9661,N_8304,N_8520);
nor U9662 (N_9662,N_8575,N_8909);
or U9663 (N_9663,N_8059,N_8979);
or U9664 (N_9664,N_8013,N_8259);
nand U9665 (N_9665,N_8832,N_8248);
nand U9666 (N_9666,N_8977,N_8113);
nand U9667 (N_9667,N_8477,N_8158);
or U9668 (N_9668,N_8708,N_8703);
and U9669 (N_9669,N_8190,N_8836);
nor U9670 (N_9670,N_8897,N_8859);
and U9671 (N_9671,N_8387,N_8562);
xor U9672 (N_9672,N_8736,N_8492);
nand U9673 (N_9673,N_8484,N_8459);
and U9674 (N_9674,N_8492,N_8793);
nand U9675 (N_9675,N_8514,N_8497);
and U9676 (N_9676,N_8614,N_8497);
nor U9677 (N_9677,N_8091,N_8340);
and U9678 (N_9678,N_8378,N_8916);
nor U9679 (N_9679,N_8538,N_8758);
and U9680 (N_9680,N_8084,N_8026);
and U9681 (N_9681,N_8967,N_8804);
nand U9682 (N_9682,N_8518,N_8276);
nand U9683 (N_9683,N_8530,N_8386);
nand U9684 (N_9684,N_8241,N_8660);
and U9685 (N_9685,N_8489,N_8066);
nand U9686 (N_9686,N_8555,N_8474);
or U9687 (N_9687,N_8997,N_8946);
nand U9688 (N_9688,N_8605,N_8970);
nor U9689 (N_9689,N_8257,N_8818);
and U9690 (N_9690,N_8749,N_8635);
or U9691 (N_9691,N_8126,N_8597);
or U9692 (N_9692,N_8165,N_8238);
nor U9693 (N_9693,N_8838,N_8414);
nand U9694 (N_9694,N_8510,N_8237);
and U9695 (N_9695,N_8909,N_8207);
and U9696 (N_9696,N_8595,N_8463);
or U9697 (N_9697,N_8928,N_8169);
and U9698 (N_9698,N_8128,N_8951);
and U9699 (N_9699,N_8157,N_8814);
or U9700 (N_9700,N_8982,N_8130);
nand U9701 (N_9701,N_8014,N_8464);
and U9702 (N_9702,N_8613,N_8907);
nand U9703 (N_9703,N_8261,N_8474);
nor U9704 (N_9704,N_8407,N_8840);
nand U9705 (N_9705,N_8234,N_8822);
nor U9706 (N_9706,N_8690,N_8906);
or U9707 (N_9707,N_8792,N_8794);
and U9708 (N_9708,N_8012,N_8099);
nand U9709 (N_9709,N_8407,N_8007);
nor U9710 (N_9710,N_8557,N_8061);
or U9711 (N_9711,N_8895,N_8426);
nand U9712 (N_9712,N_8211,N_8500);
nand U9713 (N_9713,N_8790,N_8822);
nand U9714 (N_9714,N_8636,N_8352);
or U9715 (N_9715,N_8929,N_8266);
or U9716 (N_9716,N_8874,N_8566);
nor U9717 (N_9717,N_8575,N_8520);
xor U9718 (N_9718,N_8426,N_8161);
or U9719 (N_9719,N_8938,N_8514);
or U9720 (N_9720,N_8423,N_8086);
nor U9721 (N_9721,N_8396,N_8488);
nor U9722 (N_9722,N_8234,N_8870);
nor U9723 (N_9723,N_8473,N_8498);
nor U9724 (N_9724,N_8627,N_8752);
and U9725 (N_9725,N_8861,N_8804);
and U9726 (N_9726,N_8238,N_8468);
nor U9727 (N_9727,N_8153,N_8200);
nor U9728 (N_9728,N_8378,N_8750);
xor U9729 (N_9729,N_8956,N_8928);
and U9730 (N_9730,N_8387,N_8508);
or U9731 (N_9731,N_8487,N_8875);
and U9732 (N_9732,N_8208,N_8153);
or U9733 (N_9733,N_8241,N_8493);
or U9734 (N_9734,N_8906,N_8819);
or U9735 (N_9735,N_8539,N_8447);
and U9736 (N_9736,N_8284,N_8030);
nand U9737 (N_9737,N_8546,N_8891);
or U9738 (N_9738,N_8302,N_8525);
and U9739 (N_9739,N_8299,N_8771);
and U9740 (N_9740,N_8513,N_8927);
and U9741 (N_9741,N_8124,N_8993);
or U9742 (N_9742,N_8719,N_8110);
nand U9743 (N_9743,N_8238,N_8958);
or U9744 (N_9744,N_8162,N_8229);
nand U9745 (N_9745,N_8234,N_8630);
and U9746 (N_9746,N_8907,N_8784);
nor U9747 (N_9747,N_8958,N_8042);
nand U9748 (N_9748,N_8858,N_8329);
and U9749 (N_9749,N_8578,N_8017);
nor U9750 (N_9750,N_8344,N_8661);
nand U9751 (N_9751,N_8819,N_8031);
nor U9752 (N_9752,N_8981,N_8532);
nand U9753 (N_9753,N_8732,N_8142);
nand U9754 (N_9754,N_8682,N_8370);
nand U9755 (N_9755,N_8537,N_8125);
nor U9756 (N_9756,N_8311,N_8830);
nor U9757 (N_9757,N_8430,N_8463);
and U9758 (N_9758,N_8447,N_8842);
nor U9759 (N_9759,N_8302,N_8406);
nand U9760 (N_9760,N_8341,N_8427);
nand U9761 (N_9761,N_8087,N_8716);
nand U9762 (N_9762,N_8815,N_8489);
nand U9763 (N_9763,N_8296,N_8643);
nor U9764 (N_9764,N_8710,N_8440);
nor U9765 (N_9765,N_8546,N_8208);
or U9766 (N_9766,N_8620,N_8747);
nor U9767 (N_9767,N_8210,N_8893);
and U9768 (N_9768,N_8045,N_8851);
or U9769 (N_9769,N_8350,N_8187);
nand U9770 (N_9770,N_8750,N_8477);
nand U9771 (N_9771,N_8160,N_8491);
and U9772 (N_9772,N_8074,N_8306);
nor U9773 (N_9773,N_8980,N_8899);
nand U9774 (N_9774,N_8579,N_8345);
xor U9775 (N_9775,N_8315,N_8522);
nand U9776 (N_9776,N_8929,N_8835);
nor U9777 (N_9777,N_8852,N_8413);
and U9778 (N_9778,N_8851,N_8087);
and U9779 (N_9779,N_8817,N_8496);
nor U9780 (N_9780,N_8856,N_8393);
and U9781 (N_9781,N_8874,N_8514);
nand U9782 (N_9782,N_8138,N_8598);
nor U9783 (N_9783,N_8732,N_8318);
nor U9784 (N_9784,N_8507,N_8238);
and U9785 (N_9785,N_8262,N_8041);
nand U9786 (N_9786,N_8648,N_8951);
nand U9787 (N_9787,N_8638,N_8887);
and U9788 (N_9788,N_8854,N_8626);
nand U9789 (N_9789,N_8109,N_8706);
and U9790 (N_9790,N_8181,N_8646);
or U9791 (N_9791,N_8848,N_8169);
or U9792 (N_9792,N_8145,N_8448);
nor U9793 (N_9793,N_8749,N_8784);
nor U9794 (N_9794,N_8350,N_8254);
or U9795 (N_9795,N_8422,N_8093);
nand U9796 (N_9796,N_8503,N_8987);
or U9797 (N_9797,N_8732,N_8029);
or U9798 (N_9798,N_8943,N_8821);
or U9799 (N_9799,N_8291,N_8316);
or U9800 (N_9800,N_8794,N_8491);
nor U9801 (N_9801,N_8201,N_8944);
or U9802 (N_9802,N_8879,N_8500);
or U9803 (N_9803,N_8351,N_8623);
nor U9804 (N_9804,N_8459,N_8234);
and U9805 (N_9805,N_8910,N_8795);
nand U9806 (N_9806,N_8063,N_8604);
and U9807 (N_9807,N_8295,N_8696);
nand U9808 (N_9808,N_8736,N_8642);
nand U9809 (N_9809,N_8962,N_8245);
or U9810 (N_9810,N_8546,N_8391);
nand U9811 (N_9811,N_8943,N_8583);
nor U9812 (N_9812,N_8896,N_8935);
nand U9813 (N_9813,N_8473,N_8704);
or U9814 (N_9814,N_8583,N_8746);
and U9815 (N_9815,N_8062,N_8161);
nor U9816 (N_9816,N_8311,N_8654);
and U9817 (N_9817,N_8770,N_8338);
nand U9818 (N_9818,N_8871,N_8309);
nand U9819 (N_9819,N_8005,N_8622);
and U9820 (N_9820,N_8532,N_8432);
and U9821 (N_9821,N_8525,N_8368);
and U9822 (N_9822,N_8804,N_8380);
nand U9823 (N_9823,N_8237,N_8242);
and U9824 (N_9824,N_8726,N_8420);
nand U9825 (N_9825,N_8747,N_8020);
nand U9826 (N_9826,N_8399,N_8373);
or U9827 (N_9827,N_8880,N_8950);
nand U9828 (N_9828,N_8333,N_8995);
or U9829 (N_9829,N_8420,N_8855);
nor U9830 (N_9830,N_8493,N_8733);
nand U9831 (N_9831,N_8895,N_8594);
or U9832 (N_9832,N_8813,N_8081);
nor U9833 (N_9833,N_8025,N_8394);
and U9834 (N_9834,N_8034,N_8106);
or U9835 (N_9835,N_8039,N_8784);
nand U9836 (N_9836,N_8664,N_8730);
and U9837 (N_9837,N_8176,N_8954);
nand U9838 (N_9838,N_8196,N_8339);
nand U9839 (N_9839,N_8120,N_8151);
and U9840 (N_9840,N_8272,N_8506);
nor U9841 (N_9841,N_8182,N_8636);
nor U9842 (N_9842,N_8493,N_8391);
nor U9843 (N_9843,N_8138,N_8377);
or U9844 (N_9844,N_8704,N_8630);
nand U9845 (N_9845,N_8316,N_8461);
nor U9846 (N_9846,N_8323,N_8557);
or U9847 (N_9847,N_8521,N_8273);
or U9848 (N_9848,N_8374,N_8592);
nor U9849 (N_9849,N_8468,N_8407);
nand U9850 (N_9850,N_8597,N_8830);
nor U9851 (N_9851,N_8645,N_8462);
nor U9852 (N_9852,N_8317,N_8719);
or U9853 (N_9853,N_8941,N_8529);
nor U9854 (N_9854,N_8661,N_8321);
and U9855 (N_9855,N_8482,N_8470);
or U9856 (N_9856,N_8214,N_8913);
and U9857 (N_9857,N_8437,N_8952);
or U9858 (N_9858,N_8407,N_8629);
or U9859 (N_9859,N_8007,N_8307);
nand U9860 (N_9860,N_8263,N_8012);
nor U9861 (N_9861,N_8160,N_8387);
or U9862 (N_9862,N_8690,N_8821);
nand U9863 (N_9863,N_8126,N_8957);
nand U9864 (N_9864,N_8478,N_8175);
nor U9865 (N_9865,N_8327,N_8723);
nand U9866 (N_9866,N_8097,N_8633);
and U9867 (N_9867,N_8156,N_8176);
or U9868 (N_9868,N_8821,N_8180);
and U9869 (N_9869,N_8100,N_8689);
nor U9870 (N_9870,N_8589,N_8517);
or U9871 (N_9871,N_8251,N_8214);
and U9872 (N_9872,N_8409,N_8714);
nor U9873 (N_9873,N_8173,N_8012);
nand U9874 (N_9874,N_8621,N_8192);
or U9875 (N_9875,N_8721,N_8987);
nand U9876 (N_9876,N_8794,N_8935);
nor U9877 (N_9877,N_8033,N_8055);
nor U9878 (N_9878,N_8192,N_8341);
nand U9879 (N_9879,N_8917,N_8192);
xor U9880 (N_9880,N_8385,N_8240);
nand U9881 (N_9881,N_8581,N_8381);
nand U9882 (N_9882,N_8913,N_8371);
and U9883 (N_9883,N_8106,N_8685);
or U9884 (N_9884,N_8538,N_8356);
and U9885 (N_9885,N_8254,N_8201);
and U9886 (N_9886,N_8134,N_8832);
nand U9887 (N_9887,N_8859,N_8372);
or U9888 (N_9888,N_8266,N_8113);
xor U9889 (N_9889,N_8145,N_8255);
nor U9890 (N_9890,N_8703,N_8883);
nor U9891 (N_9891,N_8857,N_8443);
and U9892 (N_9892,N_8387,N_8327);
and U9893 (N_9893,N_8529,N_8512);
nor U9894 (N_9894,N_8342,N_8948);
nand U9895 (N_9895,N_8842,N_8849);
nand U9896 (N_9896,N_8849,N_8828);
and U9897 (N_9897,N_8784,N_8401);
nand U9898 (N_9898,N_8223,N_8641);
or U9899 (N_9899,N_8645,N_8429);
and U9900 (N_9900,N_8821,N_8564);
nand U9901 (N_9901,N_8006,N_8455);
nand U9902 (N_9902,N_8893,N_8545);
and U9903 (N_9903,N_8979,N_8931);
and U9904 (N_9904,N_8995,N_8996);
and U9905 (N_9905,N_8508,N_8702);
nand U9906 (N_9906,N_8606,N_8545);
and U9907 (N_9907,N_8955,N_8457);
or U9908 (N_9908,N_8124,N_8604);
and U9909 (N_9909,N_8712,N_8000);
and U9910 (N_9910,N_8555,N_8952);
nor U9911 (N_9911,N_8032,N_8247);
and U9912 (N_9912,N_8103,N_8840);
and U9913 (N_9913,N_8030,N_8302);
nor U9914 (N_9914,N_8171,N_8136);
nor U9915 (N_9915,N_8673,N_8387);
nand U9916 (N_9916,N_8269,N_8530);
and U9917 (N_9917,N_8980,N_8495);
or U9918 (N_9918,N_8260,N_8830);
xor U9919 (N_9919,N_8891,N_8975);
nand U9920 (N_9920,N_8330,N_8204);
or U9921 (N_9921,N_8846,N_8319);
or U9922 (N_9922,N_8344,N_8056);
nand U9923 (N_9923,N_8367,N_8394);
nor U9924 (N_9924,N_8726,N_8273);
nor U9925 (N_9925,N_8271,N_8624);
nand U9926 (N_9926,N_8911,N_8730);
nand U9927 (N_9927,N_8745,N_8891);
nor U9928 (N_9928,N_8132,N_8222);
and U9929 (N_9929,N_8238,N_8606);
nor U9930 (N_9930,N_8735,N_8990);
or U9931 (N_9931,N_8188,N_8643);
nand U9932 (N_9932,N_8870,N_8347);
nor U9933 (N_9933,N_8097,N_8501);
nor U9934 (N_9934,N_8870,N_8054);
nor U9935 (N_9935,N_8245,N_8927);
or U9936 (N_9936,N_8690,N_8955);
nand U9937 (N_9937,N_8405,N_8528);
and U9938 (N_9938,N_8357,N_8096);
xor U9939 (N_9939,N_8004,N_8647);
nor U9940 (N_9940,N_8403,N_8825);
nand U9941 (N_9941,N_8688,N_8913);
or U9942 (N_9942,N_8325,N_8951);
and U9943 (N_9943,N_8911,N_8291);
nand U9944 (N_9944,N_8957,N_8603);
and U9945 (N_9945,N_8041,N_8076);
and U9946 (N_9946,N_8722,N_8127);
nor U9947 (N_9947,N_8820,N_8010);
and U9948 (N_9948,N_8590,N_8190);
nor U9949 (N_9949,N_8512,N_8159);
or U9950 (N_9950,N_8689,N_8530);
and U9951 (N_9951,N_8375,N_8081);
nand U9952 (N_9952,N_8538,N_8045);
and U9953 (N_9953,N_8366,N_8106);
nand U9954 (N_9954,N_8659,N_8849);
nand U9955 (N_9955,N_8970,N_8828);
and U9956 (N_9956,N_8142,N_8258);
nor U9957 (N_9957,N_8289,N_8165);
and U9958 (N_9958,N_8755,N_8255);
nand U9959 (N_9959,N_8933,N_8823);
and U9960 (N_9960,N_8213,N_8109);
or U9961 (N_9961,N_8252,N_8485);
and U9962 (N_9962,N_8360,N_8918);
and U9963 (N_9963,N_8602,N_8084);
nand U9964 (N_9964,N_8947,N_8473);
nor U9965 (N_9965,N_8853,N_8488);
or U9966 (N_9966,N_8914,N_8116);
or U9967 (N_9967,N_8926,N_8461);
nand U9968 (N_9968,N_8059,N_8853);
and U9969 (N_9969,N_8047,N_8522);
or U9970 (N_9970,N_8135,N_8457);
nand U9971 (N_9971,N_8698,N_8513);
or U9972 (N_9972,N_8678,N_8486);
nand U9973 (N_9973,N_8235,N_8041);
nor U9974 (N_9974,N_8771,N_8117);
or U9975 (N_9975,N_8717,N_8576);
nor U9976 (N_9976,N_8403,N_8181);
nor U9977 (N_9977,N_8229,N_8428);
or U9978 (N_9978,N_8285,N_8750);
nor U9979 (N_9979,N_8933,N_8739);
nor U9980 (N_9980,N_8918,N_8983);
and U9981 (N_9981,N_8675,N_8515);
or U9982 (N_9982,N_8065,N_8035);
and U9983 (N_9983,N_8962,N_8893);
and U9984 (N_9984,N_8270,N_8724);
or U9985 (N_9985,N_8408,N_8389);
and U9986 (N_9986,N_8637,N_8060);
nor U9987 (N_9987,N_8516,N_8989);
nor U9988 (N_9988,N_8582,N_8971);
or U9989 (N_9989,N_8354,N_8174);
or U9990 (N_9990,N_8923,N_8548);
or U9991 (N_9991,N_8659,N_8686);
or U9992 (N_9992,N_8833,N_8344);
and U9993 (N_9993,N_8608,N_8151);
and U9994 (N_9994,N_8921,N_8568);
or U9995 (N_9995,N_8043,N_8780);
nor U9996 (N_9996,N_8869,N_8040);
and U9997 (N_9997,N_8721,N_8560);
nand U9998 (N_9998,N_8345,N_8015);
and U9999 (N_9999,N_8120,N_8556);
nor UO_0 (O_0,N_9290,N_9623);
and UO_1 (O_1,N_9027,N_9598);
nand UO_2 (O_2,N_9133,N_9094);
and UO_3 (O_3,N_9003,N_9801);
or UO_4 (O_4,N_9779,N_9681);
and UO_5 (O_5,N_9359,N_9233);
or UO_6 (O_6,N_9826,N_9562);
and UO_7 (O_7,N_9506,N_9538);
nand UO_8 (O_8,N_9706,N_9237);
or UO_9 (O_9,N_9356,N_9453);
nand UO_10 (O_10,N_9895,N_9261);
or UO_11 (O_11,N_9047,N_9467);
nor UO_12 (O_12,N_9867,N_9567);
nor UO_13 (O_13,N_9518,N_9182);
or UO_14 (O_14,N_9395,N_9303);
nor UO_15 (O_15,N_9054,N_9025);
and UO_16 (O_16,N_9455,N_9354);
or UO_17 (O_17,N_9044,N_9199);
or UO_18 (O_18,N_9206,N_9722);
nor UO_19 (O_19,N_9529,N_9390);
or UO_20 (O_20,N_9600,N_9240);
nand UO_21 (O_21,N_9447,N_9316);
nand UO_22 (O_22,N_9160,N_9350);
nand UO_23 (O_23,N_9621,N_9231);
nand UO_24 (O_24,N_9573,N_9211);
and UO_25 (O_25,N_9507,N_9281);
and UO_26 (O_26,N_9406,N_9088);
or UO_27 (O_27,N_9011,N_9682);
or UO_28 (O_28,N_9360,N_9139);
nand UO_29 (O_29,N_9658,N_9012);
and UO_30 (O_30,N_9483,N_9148);
nand UO_31 (O_31,N_9813,N_9659);
xnor UO_32 (O_32,N_9664,N_9505);
or UO_33 (O_33,N_9421,N_9437);
and UO_34 (O_34,N_9570,N_9585);
and UO_35 (O_35,N_9524,N_9663);
or UO_36 (O_36,N_9081,N_9920);
nand UO_37 (O_37,N_9517,N_9549);
nor UO_38 (O_38,N_9343,N_9975);
and UO_39 (O_39,N_9187,N_9117);
nand UO_40 (O_40,N_9642,N_9721);
or UO_41 (O_41,N_9050,N_9137);
nand UO_42 (O_42,N_9900,N_9302);
nor UO_43 (O_43,N_9164,N_9781);
or UO_44 (O_44,N_9917,N_9858);
or UO_45 (O_45,N_9935,N_9702);
and UO_46 (O_46,N_9687,N_9400);
and UO_47 (O_47,N_9171,N_9479);
and UO_48 (O_48,N_9545,N_9819);
and UO_49 (O_49,N_9512,N_9926);
and UO_50 (O_50,N_9533,N_9167);
nor UO_51 (O_51,N_9474,N_9734);
and UO_52 (O_52,N_9662,N_9785);
and UO_53 (O_53,N_9454,N_9821);
nand UO_54 (O_54,N_9898,N_9970);
nand UO_55 (O_55,N_9023,N_9615);
and UO_56 (O_56,N_9030,N_9887);
or UO_57 (O_57,N_9924,N_9837);
nand UO_58 (O_58,N_9057,N_9367);
nand UO_59 (O_59,N_9019,N_9763);
and UO_60 (O_60,N_9697,N_9141);
nor UO_61 (O_61,N_9212,N_9607);
and UO_62 (O_62,N_9203,N_9449);
nor UO_63 (O_63,N_9990,N_9045);
and UO_64 (O_64,N_9296,N_9002);
nor UO_65 (O_65,N_9864,N_9803);
nor UO_66 (O_66,N_9724,N_9192);
or UO_67 (O_67,N_9641,N_9080);
nand UO_68 (O_68,N_9910,N_9964);
or UO_69 (O_69,N_9024,N_9745);
nand UO_70 (O_70,N_9105,N_9756);
or UO_71 (O_71,N_9056,N_9635);
nand UO_72 (O_72,N_9280,N_9995);
nor UO_73 (O_73,N_9099,N_9742);
or UO_74 (O_74,N_9863,N_9918);
nor UO_75 (O_75,N_9547,N_9961);
nand UO_76 (O_76,N_9005,N_9156);
and UO_77 (O_77,N_9059,N_9010);
or UO_78 (O_78,N_9413,N_9346);
and UO_79 (O_79,N_9614,N_9569);
nor UO_80 (O_80,N_9186,N_9272);
nand UO_81 (O_81,N_9960,N_9210);
or UO_82 (O_82,N_9006,N_9448);
or UO_83 (O_83,N_9202,N_9078);
or UO_84 (O_84,N_9311,N_9034);
and UO_85 (O_85,N_9852,N_9865);
and UO_86 (O_86,N_9994,N_9786);
nor UO_87 (O_87,N_9107,N_9739);
nor UO_88 (O_88,N_9124,N_9608);
and UO_89 (O_89,N_9140,N_9992);
and UO_90 (O_90,N_9007,N_9481);
or UO_91 (O_91,N_9339,N_9872);
nor UO_92 (O_92,N_9589,N_9723);
and UO_93 (O_93,N_9731,N_9844);
nand UO_94 (O_94,N_9443,N_9333);
and UO_95 (O_95,N_9675,N_9767);
and UO_96 (O_96,N_9869,N_9193);
and UO_97 (O_97,N_9435,N_9546);
nand UO_98 (O_98,N_9254,N_9725);
nand UO_99 (O_99,N_9230,N_9618);
or UO_100 (O_100,N_9520,N_9564);
nor UO_101 (O_101,N_9521,N_9499);
or UO_102 (O_102,N_9309,N_9176);
nor UO_103 (O_103,N_9277,N_9808);
and UO_104 (O_104,N_9847,N_9076);
and UO_105 (O_105,N_9065,N_9070);
or UO_106 (O_106,N_9241,N_9227);
or UO_107 (O_107,N_9735,N_9314);
or UO_108 (O_108,N_9695,N_9438);
or UO_109 (O_109,N_9669,N_9824);
and UO_110 (O_110,N_9408,N_9679);
nand UO_111 (O_111,N_9285,N_9265);
or UO_112 (O_112,N_9183,N_9509);
or UO_113 (O_113,N_9282,N_9972);
nand UO_114 (O_114,N_9415,N_9369);
nand UO_115 (O_115,N_9049,N_9266);
nor UO_116 (O_116,N_9306,N_9480);
nor UO_117 (O_117,N_9250,N_9610);
nand UO_118 (O_118,N_9829,N_9515);
and UO_119 (O_119,N_9541,N_9072);
and UO_120 (O_120,N_9357,N_9519);
nand UO_121 (O_121,N_9783,N_9861);
or UO_122 (O_122,N_9856,N_9613);
and UO_123 (O_123,N_9158,N_9712);
nor UO_124 (O_124,N_9670,N_9028);
nand UO_125 (O_125,N_9477,N_9755);
nor UO_126 (O_126,N_9778,N_9118);
nand UO_127 (O_127,N_9226,N_9322);
nand UO_128 (O_128,N_9419,N_9544);
nand UO_129 (O_129,N_9996,N_9629);
or UO_130 (O_130,N_9068,N_9301);
and UO_131 (O_131,N_9840,N_9765);
and UO_132 (O_132,N_9750,N_9175);
nand UO_133 (O_133,N_9699,N_9949);
nor UO_134 (O_134,N_9248,N_9729);
nor UO_135 (O_135,N_9827,N_9685);
or UO_136 (O_136,N_9113,N_9032);
nor UO_137 (O_137,N_9560,N_9905);
or UO_138 (O_138,N_9267,N_9096);
or UO_139 (O_139,N_9789,N_9292);
nand UO_140 (O_140,N_9436,N_9442);
or UO_141 (O_141,N_9033,N_9582);
nand UO_142 (O_142,N_9255,N_9914);
or UO_143 (O_143,N_9692,N_9643);
nor UO_144 (O_144,N_9262,N_9040);
or UO_145 (O_145,N_9458,N_9351);
nand UO_146 (O_146,N_9557,N_9283);
or UO_147 (O_147,N_9934,N_9901);
or UO_148 (O_148,N_9177,N_9603);
or UO_149 (O_149,N_9672,N_9084);
nor UO_150 (O_150,N_9784,N_9835);
nand UO_151 (O_151,N_9397,N_9403);
and UO_152 (O_152,N_9656,N_9434);
nand UO_153 (O_153,N_9691,N_9768);
or UO_154 (O_154,N_9119,N_9195);
or UO_155 (O_155,N_9200,N_9649);
nor UO_156 (O_156,N_9748,N_9074);
or UO_157 (O_157,N_9576,N_9851);
nand UO_158 (O_158,N_9432,N_9191);
or UO_159 (O_159,N_9109,N_9540);
nand UO_160 (O_160,N_9622,N_9252);
or UO_161 (O_161,N_9720,N_9606);
nor UO_162 (O_162,N_9143,N_9973);
and UO_163 (O_163,N_9657,N_9665);
nand UO_164 (O_164,N_9341,N_9147);
nand UO_165 (O_165,N_9501,N_9575);
nor UO_166 (O_166,N_9222,N_9348);
nand UO_167 (O_167,N_9583,N_9365);
nand UO_168 (O_168,N_9022,N_9769);
nor UO_169 (O_169,N_9700,N_9539);
or UO_170 (O_170,N_9381,N_9451);
nand UO_171 (O_171,N_9843,N_9269);
and UO_172 (O_172,N_9795,N_9636);
or UO_173 (O_173,N_9605,N_9980);
nand UO_174 (O_174,N_9325,N_9161);
or UO_175 (O_175,N_9839,N_9873);
nand UO_176 (O_176,N_9998,N_9071);
and UO_177 (O_177,N_9940,N_9014);
nand UO_178 (O_178,N_9198,N_9168);
nand UO_179 (O_179,N_9159,N_9761);
nor UO_180 (O_180,N_9468,N_9135);
and UO_181 (O_181,N_9718,N_9184);
or UO_182 (O_182,N_9979,N_9806);
and UO_183 (O_183,N_9411,N_9881);
or UO_184 (O_184,N_9746,N_9441);
or UO_185 (O_185,N_9812,N_9150);
nand UO_186 (O_186,N_9410,N_9379);
and UO_187 (O_187,N_9758,N_9352);
or UO_188 (O_188,N_9899,N_9897);
nand UO_189 (O_189,N_9937,N_9668);
and UO_190 (O_190,N_9083,N_9108);
and UO_191 (O_191,N_9429,N_9497);
and UO_192 (O_192,N_9792,N_9445);
and UO_193 (O_193,N_9836,N_9305);
nor UO_194 (O_194,N_9157,N_9991);
and UO_195 (O_195,N_9271,N_9149);
nor UO_196 (O_196,N_9110,N_9038);
and UO_197 (O_197,N_9207,N_9087);
nand UO_198 (O_198,N_9568,N_9772);
or UO_199 (O_199,N_9327,N_9082);
nor UO_200 (O_200,N_9661,N_9418);
or UO_201 (O_201,N_9880,N_9737);
nand UO_202 (O_202,N_9263,N_9950);
nor UO_203 (O_203,N_9300,N_9707);
and UO_204 (O_204,N_9239,N_9604);
or UO_205 (O_205,N_9152,N_9402);
and UO_206 (O_206,N_9754,N_9336);
nand UO_207 (O_207,N_9624,N_9491);
and UO_208 (O_208,N_9466,N_9091);
or UO_209 (O_209,N_9115,N_9977);
and UO_210 (O_210,N_9247,N_9104);
nand UO_211 (O_211,N_9275,N_9730);
and UO_212 (O_212,N_9586,N_9823);
and UO_213 (O_213,N_9698,N_9075);
or UO_214 (O_214,N_9951,N_9776);
and UO_215 (O_215,N_9279,N_9079);
or UO_216 (O_216,N_9578,N_9759);
nand UO_217 (O_217,N_9425,N_9253);
and UO_218 (O_218,N_9154,N_9417);
nor UO_219 (O_219,N_9422,N_9470);
nor UO_220 (O_220,N_9896,N_9132);
nor UO_221 (O_221,N_9052,N_9828);
nand UO_222 (O_222,N_9450,N_9751);
nand UO_223 (O_223,N_9749,N_9249);
nor UO_224 (O_224,N_9554,N_9955);
nor UO_225 (O_225,N_9787,N_9256);
nor UO_226 (O_226,N_9609,N_9324);
or UO_227 (O_227,N_9018,N_9845);
nor UO_228 (O_228,N_9764,N_9220);
nor UO_229 (O_229,N_9085,N_9475);
or UO_230 (O_230,N_9891,N_9185);
nor UO_231 (O_231,N_9911,N_9138);
and UO_232 (O_232,N_9457,N_9883);
nor UO_233 (O_233,N_9962,N_9811);
nand UO_234 (O_234,N_9574,N_9871);
or UO_235 (O_235,N_9958,N_9988);
or UO_236 (O_236,N_9055,N_9294);
or UO_237 (O_237,N_9594,N_9375);
nor UO_238 (O_238,N_9903,N_9342);
nor UO_239 (O_239,N_9577,N_9602);
or UO_240 (O_240,N_9331,N_9486);
or UO_241 (O_241,N_9719,N_9259);
or UO_242 (O_242,N_9671,N_9634);
or UO_243 (O_243,N_9654,N_9162);
and UO_244 (O_244,N_9209,N_9217);
or UO_245 (O_245,N_9771,N_9092);
or UO_246 (O_246,N_9144,N_9472);
nand UO_247 (O_247,N_9894,N_9553);
and UO_248 (O_248,N_9460,N_9944);
nor UO_249 (O_249,N_9705,N_9987);
or UO_250 (O_250,N_9974,N_9713);
and UO_251 (O_251,N_9216,N_9062);
and UO_252 (O_252,N_9584,N_9116);
nor UO_253 (O_253,N_9374,N_9295);
nand UO_254 (O_254,N_9304,N_9503);
nor UO_255 (O_255,N_9798,N_9368);
and UO_256 (O_256,N_9627,N_9537);
nand UO_257 (O_257,N_9464,N_9915);
nor UO_258 (O_258,N_9444,N_9525);
or UO_259 (O_259,N_9593,N_9923);
or UO_260 (O_260,N_9978,N_9257);
and UO_261 (O_261,N_9572,N_9715);
nand UO_262 (O_262,N_9617,N_9596);
and UO_263 (O_263,N_9888,N_9630);
and UO_264 (O_264,N_9373,N_9726);
nand UO_265 (O_265,N_9985,N_9932);
and UO_266 (O_266,N_9652,N_9245);
nand UO_267 (O_267,N_9362,N_9041);
nand UO_268 (O_268,N_9592,N_9875);
nor UO_269 (O_269,N_9879,N_9551);
or UO_270 (O_270,N_9225,N_9482);
nand UO_271 (O_271,N_9866,N_9361);
and UO_272 (O_272,N_9743,N_9939);
nor UO_273 (O_273,N_9640,N_9244);
and UO_274 (O_274,N_9841,N_9163);
nor UO_275 (O_275,N_9552,N_9588);
nor UO_276 (O_276,N_9431,N_9371);
or UO_277 (O_277,N_9462,N_9153);
xor UO_278 (O_278,N_9077,N_9051);
or UO_279 (O_279,N_9859,N_9831);
and UO_280 (O_280,N_9456,N_9407);
nand UO_281 (O_281,N_9439,N_9902);
or UO_282 (O_282,N_9571,N_9676);
or UO_283 (O_283,N_9126,N_9967);
nand UO_284 (O_284,N_9794,N_9580);
nor UO_285 (O_285,N_9326,N_9928);
nor UO_286 (O_286,N_9619,N_9878);
and UO_287 (O_287,N_9293,N_9971);
and UO_288 (O_288,N_9101,N_9814);
nor UO_289 (O_289,N_9732,N_9733);
nor UO_290 (O_290,N_9969,N_9550);
nand UO_291 (O_291,N_9953,N_9908);
nand UO_292 (O_292,N_9492,N_9264);
or UO_293 (O_293,N_9416,N_9031);
nor UO_294 (O_294,N_9907,N_9377);
and UO_295 (O_295,N_9334,N_9633);
nand UO_296 (O_296,N_9744,N_9016);
or UO_297 (O_297,N_9628,N_9892);
and UO_298 (O_298,N_9531,N_9963);
or UO_299 (O_299,N_9493,N_9204);
and UO_300 (O_300,N_9516,N_9678);
or UO_301 (O_301,N_9136,N_9461);
nand UO_302 (O_302,N_9535,N_9142);
nand UO_303 (O_303,N_9412,N_9850);
nand UO_304 (O_304,N_9922,N_9004);
and UO_305 (O_305,N_9484,N_9830);
nand UO_306 (O_306,N_9386,N_9906);
and UO_307 (O_307,N_9433,N_9223);
nand UO_308 (O_308,N_9876,N_9297);
and UO_309 (O_309,N_9620,N_9612);
or UO_310 (O_310,N_9145,N_9999);
or UO_311 (O_311,N_9810,N_9009);
and UO_312 (O_312,N_9638,N_9542);
nor UO_313 (O_313,N_9208,N_9921);
nand UO_314 (O_314,N_9860,N_9563);
nor UO_315 (O_315,N_9793,N_9965);
or UO_316 (O_316,N_9340,N_9762);
nor UO_317 (O_317,N_9766,N_9655);
nand UO_318 (O_318,N_9258,N_9982);
or UO_319 (O_319,N_9561,N_9423);
nor UO_320 (O_320,N_9318,N_9349);
nand UO_321 (O_321,N_9180,N_9114);
and UO_322 (O_322,N_9328,N_9215);
nor UO_323 (O_323,N_9409,N_9120);
or UO_324 (O_324,N_9355,N_9129);
nand UO_325 (O_325,N_9067,N_9853);
nor UO_326 (O_326,N_9854,N_9882);
and UO_327 (O_327,N_9112,N_9488);
nor UO_328 (O_328,N_9674,N_9173);
or UO_329 (O_329,N_9530,N_9774);
and UO_330 (O_330,N_9338,N_9945);
nor UO_331 (O_331,N_9645,N_9727);
nand UO_332 (O_332,N_9452,N_9708);
nor UO_333 (O_333,N_9399,N_9644);
or UO_334 (O_334,N_9363,N_9378);
and UO_335 (O_335,N_9036,N_9274);
or UO_336 (O_336,N_9048,N_9639);
and UO_337 (O_337,N_9251,N_9807);
or UO_338 (O_338,N_9565,N_9337);
nor UO_339 (O_339,N_9490,N_9086);
nand UO_340 (O_340,N_9956,N_9205);
nand UO_341 (O_341,N_9816,N_9330);
and UO_342 (O_342,N_9242,N_9268);
and UO_343 (O_343,N_9221,N_9376);
nor UO_344 (O_344,N_9782,N_9959);
nor UO_345 (O_345,N_9832,N_9201);
nor UO_346 (O_346,N_9246,N_9260);
nor UO_347 (O_347,N_9401,N_9601);
nand UO_348 (O_348,N_9757,N_9954);
nor UO_349 (O_349,N_9273,N_9465);
nand UO_350 (O_350,N_9849,N_9666);
and UO_351 (O_351,N_9913,N_9947);
and UO_352 (O_352,N_9653,N_9820);
nand UO_353 (O_353,N_9893,N_9952);
or UO_354 (O_354,N_9123,N_9693);
nor UO_355 (O_355,N_9232,N_9428);
nor UO_356 (O_356,N_9064,N_9389);
nand UO_357 (O_357,N_9799,N_9696);
and UO_358 (O_358,N_9008,N_9513);
nand UO_359 (O_359,N_9528,N_9728);
nand UO_360 (O_360,N_9625,N_9134);
and UO_361 (O_361,N_9889,N_9276);
or UO_362 (O_362,N_9741,N_9393);
and UO_363 (O_363,N_9286,N_9523);
and UO_364 (O_364,N_9353,N_9704);
or UO_365 (O_365,N_9058,N_9485);
and UO_366 (O_366,N_9556,N_9214);
nand UO_367 (O_367,N_9380,N_9777);
and UO_368 (O_368,N_9637,N_9414);
and UO_369 (O_369,N_9647,N_9838);
and UO_370 (O_370,N_9877,N_9364);
nor UO_371 (O_371,N_9155,N_9308);
or UO_372 (O_372,N_9405,N_9502);
and UO_373 (O_373,N_9536,N_9121);
nor UO_374 (O_374,N_9329,N_9013);
nor UO_375 (O_375,N_9870,N_9494);
and UO_376 (O_376,N_9775,N_9689);
and UO_377 (O_377,N_9287,N_9815);
or UO_378 (O_378,N_9335,N_9976);
and UO_379 (O_379,N_9714,N_9650);
nand UO_380 (O_380,N_9151,N_9857);
nor UO_381 (O_381,N_9344,N_9595);
nand UO_382 (O_382,N_9886,N_9463);
nor UO_383 (O_383,N_9919,N_9738);
and UO_384 (O_384,N_9802,N_9385);
or UO_385 (O_385,N_9053,N_9818);
or UO_386 (O_386,N_9760,N_9319);
nand UO_387 (O_387,N_9066,N_9825);
or UO_388 (O_388,N_9098,N_9383);
nand UO_389 (O_389,N_9703,N_9788);
nand UO_390 (O_390,N_9504,N_9912);
and UO_391 (O_391,N_9218,N_9420);
nor UO_392 (O_392,N_9511,N_9868);
or UO_393 (O_393,N_9424,N_9986);
or UO_394 (O_394,N_9194,N_9370);
and UO_395 (O_395,N_9904,N_9646);
nand UO_396 (O_396,N_9291,N_9323);
nor UO_397 (O_397,N_9234,N_9073);
and UO_398 (O_398,N_9943,N_9046);
and UO_399 (O_399,N_9931,N_9299);
nor UO_400 (O_400,N_9968,N_9235);
and UO_401 (O_401,N_9189,N_9270);
and UO_402 (O_402,N_9885,N_9229);
and UO_403 (O_403,N_9347,N_9042);
or UO_404 (O_404,N_9688,N_9809);
nand UO_405 (O_405,N_9566,N_9398);
nor UO_406 (O_406,N_9446,N_9833);
nor UO_407 (O_407,N_9862,N_9938);
and UO_408 (O_408,N_9890,N_9927);
nand UO_409 (O_409,N_9473,N_9307);
or UO_410 (O_410,N_9984,N_9321);
or UO_411 (O_411,N_9496,N_9532);
nand UO_412 (O_412,N_9489,N_9320);
and UO_413 (O_413,N_9579,N_9534);
or UO_414 (O_414,N_9061,N_9800);
or UO_415 (O_415,N_9855,N_9315);
nor UO_416 (O_416,N_9243,N_9174);
nand UO_417 (O_417,N_9916,N_9558);
or UO_418 (O_418,N_9372,N_9817);
nor UO_419 (O_419,N_9312,N_9394);
xnor UO_420 (O_420,N_9667,N_9948);
and UO_421 (O_421,N_9111,N_9165);
or UO_422 (O_422,N_9093,N_9581);
or UO_423 (O_423,N_9000,N_9966);
and UO_424 (O_424,N_9993,N_9514);
or UO_425 (O_425,N_9128,N_9392);
nand UO_426 (O_426,N_9037,N_9805);
and UO_427 (O_427,N_9021,N_9543);
nor UO_428 (O_428,N_9178,N_9611);
nand UO_429 (O_429,N_9063,N_9388);
and UO_430 (O_430,N_9382,N_9317);
or UO_431 (O_431,N_9471,N_9020);
xnor UO_432 (O_432,N_9500,N_9122);
and UO_433 (O_433,N_9701,N_9387);
and UO_434 (O_434,N_9957,N_9170);
or UO_435 (O_435,N_9941,N_9790);
and UO_436 (O_436,N_9289,N_9213);
and UO_437 (O_437,N_9591,N_9780);
and UO_438 (O_438,N_9228,N_9469);
nor UO_439 (O_439,N_9770,N_9555);
nand UO_440 (O_440,N_9660,N_9190);
and UO_441 (O_441,N_9396,N_9060);
and UO_442 (O_442,N_9100,N_9404);
or UO_443 (O_443,N_9773,N_9478);
nor UO_444 (O_444,N_9278,N_9172);
and UO_445 (O_445,N_9527,N_9196);
nand UO_446 (O_446,N_9616,N_9933);
nand UO_447 (O_447,N_9587,N_9391);
or UO_448 (O_448,N_9874,N_9834);
nand UO_449 (O_449,N_9332,N_9043);
nor UO_450 (O_450,N_9288,N_9179);
nor UO_451 (O_451,N_9102,N_9752);
or UO_452 (O_452,N_9313,N_9476);
or UO_453 (O_453,N_9804,N_9181);
nand UO_454 (O_454,N_9753,N_9236);
nor UO_455 (O_455,N_9711,N_9736);
nand UO_456 (O_456,N_9690,N_9526);
or UO_457 (O_457,N_9632,N_9626);
and UO_458 (O_458,N_9197,N_9716);
or UO_459 (O_459,N_9125,N_9131);
or UO_460 (O_460,N_9842,N_9942);
nand UO_461 (O_461,N_9946,N_9683);
nand UO_462 (O_462,N_9680,N_9169);
or UO_463 (O_463,N_9686,N_9345);
nor UO_464 (O_464,N_9599,N_9188);
or UO_465 (O_465,N_9310,N_9366);
or UO_466 (O_466,N_9936,N_9358);
and UO_467 (O_467,N_9797,N_9747);
nor UO_468 (O_468,N_9498,N_9740);
and UO_469 (O_469,N_9548,N_9035);
nor UO_470 (O_470,N_9284,N_9384);
nand UO_471 (O_471,N_9069,N_9130);
or UO_472 (O_472,N_9981,N_9459);
and UO_473 (O_473,N_9426,N_9106);
nor UO_474 (O_474,N_9590,N_9709);
or UO_475 (O_475,N_9648,N_9029);
nor UO_476 (O_476,N_9146,N_9015);
nor UO_477 (O_477,N_9694,N_9929);
and UO_478 (O_478,N_9846,N_9983);
and UO_479 (O_479,N_9224,N_9430);
and UO_480 (O_480,N_9522,N_9039);
xor UO_481 (O_481,N_9095,N_9127);
nor UO_482 (O_482,N_9791,N_9298);
and UO_483 (O_483,N_9427,N_9884);
or UO_484 (O_484,N_9090,N_9717);
and UO_485 (O_485,N_9097,N_9238);
nor UO_486 (O_486,N_9559,N_9508);
or UO_487 (O_487,N_9822,N_9930);
or UO_488 (O_488,N_9026,N_9651);
nand UO_489 (O_489,N_9997,N_9684);
nand UO_490 (O_490,N_9710,N_9017);
nand UO_491 (O_491,N_9597,N_9001);
and UO_492 (O_492,N_9909,N_9677);
nand UO_493 (O_493,N_9219,N_9103);
and UO_494 (O_494,N_9495,N_9166);
or UO_495 (O_495,N_9510,N_9848);
nor UO_496 (O_496,N_9487,N_9440);
nor UO_497 (O_497,N_9673,N_9796);
or UO_498 (O_498,N_9089,N_9631);
nor UO_499 (O_499,N_9989,N_9925);
nand UO_500 (O_500,N_9112,N_9118);
and UO_501 (O_501,N_9051,N_9221);
or UO_502 (O_502,N_9613,N_9183);
nor UO_503 (O_503,N_9960,N_9471);
and UO_504 (O_504,N_9953,N_9840);
and UO_505 (O_505,N_9968,N_9956);
nor UO_506 (O_506,N_9733,N_9279);
nor UO_507 (O_507,N_9092,N_9730);
nand UO_508 (O_508,N_9714,N_9230);
and UO_509 (O_509,N_9967,N_9872);
nand UO_510 (O_510,N_9288,N_9575);
nand UO_511 (O_511,N_9203,N_9506);
or UO_512 (O_512,N_9936,N_9240);
xor UO_513 (O_513,N_9502,N_9995);
or UO_514 (O_514,N_9710,N_9550);
and UO_515 (O_515,N_9319,N_9420);
nor UO_516 (O_516,N_9108,N_9131);
or UO_517 (O_517,N_9549,N_9510);
nor UO_518 (O_518,N_9408,N_9159);
nor UO_519 (O_519,N_9235,N_9481);
or UO_520 (O_520,N_9382,N_9226);
nor UO_521 (O_521,N_9117,N_9858);
or UO_522 (O_522,N_9973,N_9981);
and UO_523 (O_523,N_9449,N_9298);
or UO_524 (O_524,N_9068,N_9723);
or UO_525 (O_525,N_9873,N_9351);
nor UO_526 (O_526,N_9090,N_9172);
or UO_527 (O_527,N_9887,N_9582);
nor UO_528 (O_528,N_9607,N_9162);
and UO_529 (O_529,N_9174,N_9936);
or UO_530 (O_530,N_9633,N_9447);
nand UO_531 (O_531,N_9933,N_9090);
and UO_532 (O_532,N_9386,N_9405);
nand UO_533 (O_533,N_9400,N_9229);
or UO_534 (O_534,N_9083,N_9727);
and UO_535 (O_535,N_9000,N_9185);
nor UO_536 (O_536,N_9650,N_9594);
nand UO_537 (O_537,N_9438,N_9192);
nor UO_538 (O_538,N_9110,N_9530);
and UO_539 (O_539,N_9240,N_9237);
and UO_540 (O_540,N_9507,N_9513);
and UO_541 (O_541,N_9032,N_9656);
nand UO_542 (O_542,N_9415,N_9615);
nor UO_543 (O_543,N_9338,N_9427);
and UO_544 (O_544,N_9263,N_9167);
and UO_545 (O_545,N_9349,N_9772);
or UO_546 (O_546,N_9806,N_9763);
or UO_547 (O_547,N_9067,N_9839);
and UO_548 (O_548,N_9822,N_9251);
nand UO_549 (O_549,N_9828,N_9848);
and UO_550 (O_550,N_9997,N_9100);
or UO_551 (O_551,N_9890,N_9539);
nand UO_552 (O_552,N_9544,N_9417);
nor UO_553 (O_553,N_9495,N_9431);
nand UO_554 (O_554,N_9412,N_9503);
or UO_555 (O_555,N_9220,N_9955);
or UO_556 (O_556,N_9151,N_9288);
or UO_557 (O_557,N_9539,N_9288);
and UO_558 (O_558,N_9143,N_9315);
or UO_559 (O_559,N_9972,N_9489);
and UO_560 (O_560,N_9882,N_9597);
nand UO_561 (O_561,N_9803,N_9929);
and UO_562 (O_562,N_9726,N_9795);
nor UO_563 (O_563,N_9209,N_9278);
or UO_564 (O_564,N_9545,N_9614);
nor UO_565 (O_565,N_9908,N_9354);
and UO_566 (O_566,N_9478,N_9367);
nand UO_567 (O_567,N_9069,N_9949);
nand UO_568 (O_568,N_9178,N_9003);
or UO_569 (O_569,N_9726,N_9648);
and UO_570 (O_570,N_9678,N_9345);
and UO_571 (O_571,N_9707,N_9690);
or UO_572 (O_572,N_9637,N_9585);
nand UO_573 (O_573,N_9871,N_9297);
nand UO_574 (O_574,N_9343,N_9484);
or UO_575 (O_575,N_9488,N_9109);
and UO_576 (O_576,N_9167,N_9702);
nand UO_577 (O_577,N_9515,N_9876);
and UO_578 (O_578,N_9495,N_9738);
nor UO_579 (O_579,N_9329,N_9671);
nand UO_580 (O_580,N_9618,N_9867);
and UO_581 (O_581,N_9627,N_9176);
nor UO_582 (O_582,N_9520,N_9861);
and UO_583 (O_583,N_9524,N_9350);
and UO_584 (O_584,N_9391,N_9964);
and UO_585 (O_585,N_9925,N_9354);
nor UO_586 (O_586,N_9577,N_9275);
or UO_587 (O_587,N_9813,N_9845);
xnor UO_588 (O_588,N_9497,N_9563);
and UO_589 (O_589,N_9307,N_9960);
xnor UO_590 (O_590,N_9391,N_9835);
and UO_591 (O_591,N_9659,N_9980);
and UO_592 (O_592,N_9158,N_9913);
nand UO_593 (O_593,N_9761,N_9561);
and UO_594 (O_594,N_9751,N_9159);
and UO_595 (O_595,N_9158,N_9459);
and UO_596 (O_596,N_9731,N_9105);
or UO_597 (O_597,N_9376,N_9346);
and UO_598 (O_598,N_9448,N_9242);
or UO_599 (O_599,N_9478,N_9383);
and UO_600 (O_600,N_9224,N_9696);
or UO_601 (O_601,N_9948,N_9601);
nand UO_602 (O_602,N_9939,N_9890);
or UO_603 (O_603,N_9958,N_9900);
nand UO_604 (O_604,N_9776,N_9716);
and UO_605 (O_605,N_9568,N_9327);
nand UO_606 (O_606,N_9968,N_9178);
and UO_607 (O_607,N_9385,N_9211);
xor UO_608 (O_608,N_9482,N_9539);
nand UO_609 (O_609,N_9961,N_9644);
and UO_610 (O_610,N_9593,N_9601);
nor UO_611 (O_611,N_9776,N_9796);
and UO_612 (O_612,N_9002,N_9050);
nor UO_613 (O_613,N_9692,N_9737);
and UO_614 (O_614,N_9806,N_9253);
or UO_615 (O_615,N_9754,N_9021);
and UO_616 (O_616,N_9219,N_9720);
or UO_617 (O_617,N_9820,N_9963);
nand UO_618 (O_618,N_9115,N_9689);
and UO_619 (O_619,N_9351,N_9145);
and UO_620 (O_620,N_9761,N_9259);
or UO_621 (O_621,N_9133,N_9376);
or UO_622 (O_622,N_9538,N_9236);
and UO_623 (O_623,N_9316,N_9059);
and UO_624 (O_624,N_9810,N_9941);
nor UO_625 (O_625,N_9561,N_9389);
nand UO_626 (O_626,N_9952,N_9897);
nor UO_627 (O_627,N_9050,N_9967);
or UO_628 (O_628,N_9206,N_9108);
nand UO_629 (O_629,N_9928,N_9998);
nor UO_630 (O_630,N_9294,N_9466);
nand UO_631 (O_631,N_9546,N_9849);
nand UO_632 (O_632,N_9136,N_9251);
nor UO_633 (O_633,N_9843,N_9225);
nor UO_634 (O_634,N_9838,N_9924);
nand UO_635 (O_635,N_9407,N_9327);
and UO_636 (O_636,N_9675,N_9649);
nor UO_637 (O_637,N_9034,N_9932);
nor UO_638 (O_638,N_9066,N_9442);
nor UO_639 (O_639,N_9782,N_9456);
nand UO_640 (O_640,N_9460,N_9243);
or UO_641 (O_641,N_9462,N_9069);
and UO_642 (O_642,N_9210,N_9203);
nor UO_643 (O_643,N_9314,N_9851);
nor UO_644 (O_644,N_9998,N_9512);
and UO_645 (O_645,N_9612,N_9953);
nor UO_646 (O_646,N_9934,N_9625);
nand UO_647 (O_647,N_9461,N_9372);
and UO_648 (O_648,N_9613,N_9004);
nor UO_649 (O_649,N_9447,N_9828);
or UO_650 (O_650,N_9886,N_9249);
or UO_651 (O_651,N_9547,N_9936);
or UO_652 (O_652,N_9367,N_9274);
nor UO_653 (O_653,N_9369,N_9956);
and UO_654 (O_654,N_9911,N_9862);
nand UO_655 (O_655,N_9882,N_9309);
and UO_656 (O_656,N_9201,N_9365);
nand UO_657 (O_657,N_9492,N_9031);
or UO_658 (O_658,N_9756,N_9199);
nand UO_659 (O_659,N_9514,N_9257);
nor UO_660 (O_660,N_9928,N_9602);
nor UO_661 (O_661,N_9756,N_9094);
and UO_662 (O_662,N_9881,N_9875);
nor UO_663 (O_663,N_9786,N_9291);
nor UO_664 (O_664,N_9842,N_9225);
or UO_665 (O_665,N_9301,N_9412);
nand UO_666 (O_666,N_9824,N_9935);
nand UO_667 (O_667,N_9610,N_9074);
nor UO_668 (O_668,N_9228,N_9215);
nor UO_669 (O_669,N_9313,N_9273);
nand UO_670 (O_670,N_9614,N_9407);
and UO_671 (O_671,N_9579,N_9189);
nor UO_672 (O_672,N_9007,N_9610);
nand UO_673 (O_673,N_9102,N_9610);
or UO_674 (O_674,N_9963,N_9538);
and UO_675 (O_675,N_9234,N_9387);
and UO_676 (O_676,N_9090,N_9177);
nor UO_677 (O_677,N_9884,N_9908);
and UO_678 (O_678,N_9010,N_9086);
or UO_679 (O_679,N_9181,N_9078);
nor UO_680 (O_680,N_9606,N_9016);
nor UO_681 (O_681,N_9118,N_9998);
nor UO_682 (O_682,N_9128,N_9559);
or UO_683 (O_683,N_9554,N_9570);
or UO_684 (O_684,N_9280,N_9377);
nor UO_685 (O_685,N_9674,N_9916);
nand UO_686 (O_686,N_9843,N_9969);
nor UO_687 (O_687,N_9286,N_9437);
and UO_688 (O_688,N_9163,N_9287);
or UO_689 (O_689,N_9173,N_9451);
and UO_690 (O_690,N_9505,N_9981);
and UO_691 (O_691,N_9774,N_9430);
xor UO_692 (O_692,N_9334,N_9620);
nor UO_693 (O_693,N_9512,N_9033);
nor UO_694 (O_694,N_9414,N_9277);
or UO_695 (O_695,N_9266,N_9828);
or UO_696 (O_696,N_9045,N_9114);
nand UO_697 (O_697,N_9473,N_9201);
or UO_698 (O_698,N_9164,N_9285);
or UO_699 (O_699,N_9351,N_9857);
nand UO_700 (O_700,N_9310,N_9399);
and UO_701 (O_701,N_9852,N_9576);
and UO_702 (O_702,N_9210,N_9613);
and UO_703 (O_703,N_9245,N_9581);
or UO_704 (O_704,N_9347,N_9859);
or UO_705 (O_705,N_9085,N_9155);
and UO_706 (O_706,N_9054,N_9487);
and UO_707 (O_707,N_9847,N_9948);
nor UO_708 (O_708,N_9454,N_9340);
nor UO_709 (O_709,N_9761,N_9486);
nand UO_710 (O_710,N_9482,N_9463);
and UO_711 (O_711,N_9177,N_9642);
nor UO_712 (O_712,N_9907,N_9422);
nand UO_713 (O_713,N_9433,N_9638);
or UO_714 (O_714,N_9785,N_9550);
and UO_715 (O_715,N_9306,N_9323);
nor UO_716 (O_716,N_9317,N_9629);
nand UO_717 (O_717,N_9552,N_9719);
nand UO_718 (O_718,N_9999,N_9048);
nand UO_719 (O_719,N_9517,N_9673);
nand UO_720 (O_720,N_9274,N_9042);
nor UO_721 (O_721,N_9145,N_9816);
and UO_722 (O_722,N_9499,N_9019);
or UO_723 (O_723,N_9166,N_9391);
and UO_724 (O_724,N_9773,N_9576);
nand UO_725 (O_725,N_9495,N_9581);
nand UO_726 (O_726,N_9306,N_9201);
nand UO_727 (O_727,N_9899,N_9432);
and UO_728 (O_728,N_9018,N_9816);
nand UO_729 (O_729,N_9353,N_9323);
nor UO_730 (O_730,N_9966,N_9497);
nand UO_731 (O_731,N_9816,N_9672);
nor UO_732 (O_732,N_9652,N_9817);
nand UO_733 (O_733,N_9695,N_9117);
and UO_734 (O_734,N_9403,N_9146);
or UO_735 (O_735,N_9695,N_9431);
or UO_736 (O_736,N_9396,N_9620);
and UO_737 (O_737,N_9383,N_9797);
nor UO_738 (O_738,N_9995,N_9346);
nor UO_739 (O_739,N_9669,N_9024);
nand UO_740 (O_740,N_9991,N_9177);
or UO_741 (O_741,N_9546,N_9170);
and UO_742 (O_742,N_9859,N_9306);
and UO_743 (O_743,N_9781,N_9021);
and UO_744 (O_744,N_9805,N_9234);
nor UO_745 (O_745,N_9080,N_9883);
nand UO_746 (O_746,N_9051,N_9697);
and UO_747 (O_747,N_9477,N_9107);
nand UO_748 (O_748,N_9948,N_9250);
nor UO_749 (O_749,N_9839,N_9127);
and UO_750 (O_750,N_9929,N_9956);
nor UO_751 (O_751,N_9561,N_9811);
and UO_752 (O_752,N_9745,N_9940);
nand UO_753 (O_753,N_9413,N_9496);
nor UO_754 (O_754,N_9994,N_9283);
nor UO_755 (O_755,N_9898,N_9946);
nand UO_756 (O_756,N_9985,N_9277);
and UO_757 (O_757,N_9668,N_9923);
nor UO_758 (O_758,N_9146,N_9581);
or UO_759 (O_759,N_9510,N_9304);
nand UO_760 (O_760,N_9864,N_9924);
or UO_761 (O_761,N_9803,N_9664);
nand UO_762 (O_762,N_9053,N_9257);
nor UO_763 (O_763,N_9715,N_9029);
nor UO_764 (O_764,N_9391,N_9056);
nand UO_765 (O_765,N_9923,N_9095);
or UO_766 (O_766,N_9514,N_9098);
nor UO_767 (O_767,N_9600,N_9799);
nor UO_768 (O_768,N_9065,N_9486);
and UO_769 (O_769,N_9792,N_9023);
nand UO_770 (O_770,N_9460,N_9476);
nor UO_771 (O_771,N_9572,N_9603);
and UO_772 (O_772,N_9093,N_9954);
or UO_773 (O_773,N_9379,N_9682);
or UO_774 (O_774,N_9275,N_9431);
or UO_775 (O_775,N_9044,N_9547);
and UO_776 (O_776,N_9857,N_9252);
and UO_777 (O_777,N_9340,N_9739);
nor UO_778 (O_778,N_9193,N_9514);
or UO_779 (O_779,N_9052,N_9240);
nor UO_780 (O_780,N_9415,N_9190);
nor UO_781 (O_781,N_9615,N_9425);
nor UO_782 (O_782,N_9928,N_9917);
and UO_783 (O_783,N_9919,N_9434);
or UO_784 (O_784,N_9911,N_9028);
or UO_785 (O_785,N_9359,N_9897);
and UO_786 (O_786,N_9672,N_9002);
and UO_787 (O_787,N_9098,N_9061);
nand UO_788 (O_788,N_9244,N_9212);
nor UO_789 (O_789,N_9057,N_9981);
nor UO_790 (O_790,N_9463,N_9752);
nand UO_791 (O_791,N_9843,N_9526);
nor UO_792 (O_792,N_9924,N_9801);
nor UO_793 (O_793,N_9404,N_9287);
or UO_794 (O_794,N_9751,N_9708);
and UO_795 (O_795,N_9381,N_9227);
or UO_796 (O_796,N_9788,N_9486);
or UO_797 (O_797,N_9055,N_9385);
or UO_798 (O_798,N_9559,N_9613);
nand UO_799 (O_799,N_9250,N_9917);
nor UO_800 (O_800,N_9901,N_9503);
and UO_801 (O_801,N_9572,N_9534);
and UO_802 (O_802,N_9657,N_9406);
nand UO_803 (O_803,N_9743,N_9252);
and UO_804 (O_804,N_9128,N_9524);
nor UO_805 (O_805,N_9970,N_9683);
and UO_806 (O_806,N_9041,N_9788);
nor UO_807 (O_807,N_9711,N_9414);
and UO_808 (O_808,N_9826,N_9564);
nor UO_809 (O_809,N_9637,N_9492);
or UO_810 (O_810,N_9886,N_9922);
or UO_811 (O_811,N_9535,N_9279);
or UO_812 (O_812,N_9620,N_9154);
nand UO_813 (O_813,N_9300,N_9019);
nor UO_814 (O_814,N_9682,N_9343);
or UO_815 (O_815,N_9162,N_9249);
nand UO_816 (O_816,N_9990,N_9617);
nand UO_817 (O_817,N_9722,N_9486);
or UO_818 (O_818,N_9685,N_9756);
or UO_819 (O_819,N_9392,N_9895);
nand UO_820 (O_820,N_9557,N_9646);
or UO_821 (O_821,N_9948,N_9950);
or UO_822 (O_822,N_9358,N_9834);
nor UO_823 (O_823,N_9960,N_9830);
nor UO_824 (O_824,N_9961,N_9663);
and UO_825 (O_825,N_9923,N_9098);
nor UO_826 (O_826,N_9298,N_9052);
nor UO_827 (O_827,N_9503,N_9121);
or UO_828 (O_828,N_9315,N_9660);
nand UO_829 (O_829,N_9373,N_9079);
nand UO_830 (O_830,N_9774,N_9560);
and UO_831 (O_831,N_9572,N_9294);
or UO_832 (O_832,N_9636,N_9996);
and UO_833 (O_833,N_9564,N_9736);
nor UO_834 (O_834,N_9021,N_9965);
nor UO_835 (O_835,N_9867,N_9003);
or UO_836 (O_836,N_9144,N_9211);
or UO_837 (O_837,N_9281,N_9138);
nor UO_838 (O_838,N_9063,N_9176);
or UO_839 (O_839,N_9264,N_9842);
and UO_840 (O_840,N_9858,N_9390);
nor UO_841 (O_841,N_9046,N_9948);
nand UO_842 (O_842,N_9642,N_9334);
or UO_843 (O_843,N_9650,N_9138);
or UO_844 (O_844,N_9532,N_9447);
nand UO_845 (O_845,N_9615,N_9551);
and UO_846 (O_846,N_9711,N_9692);
and UO_847 (O_847,N_9821,N_9715);
nor UO_848 (O_848,N_9737,N_9646);
and UO_849 (O_849,N_9620,N_9647);
nand UO_850 (O_850,N_9620,N_9486);
nand UO_851 (O_851,N_9857,N_9578);
nand UO_852 (O_852,N_9308,N_9972);
xor UO_853 (O_853,N_9787,N_9276);
nand UO_854 (O_854,N_9757,N_9998);
or UO_855 (O_855,N_9717,N_9169);
or UO_856 (O_856,N_9148,N_9777);
nor UO_857 (O_857,N_9250,N_9574);
nor UO_858 (O_858,N_9375,N_9026);
and UO_859 (O_859,N_9902,N_9512);
and UO_860 (O_860,N_9277,N_9145);
or UO_861 (O_861,N_9860,N_9206);
or UO_862 (O_862,N_9817,N_9798);
and UO_863 (O_863,N_9990,N_9753);
nand UO_864 (O_864,N_9506,N_9972);
nor UO_865 (O_865,N_9208,N_9802);
nor UO_866 (O_866,N_9099,N_9700);
or UO_867 (O_867,N_9018,N_9711);
or UO_868 (O_868,N_9170,N_9431);
and UO_869 (O_869,N_9301,N_9211);
and UO_870 (O_870,N_9886,N_9207);
nor UO_871 (O_871,N_9769,N_9265);
nand UO_872 (O_872,N_9040,N_9647);
nor UO_873 (O_873,N_9098,N_9689);
and UO_874 (O_874,N_9068,N_9789);
nor UO_875 (O_875,N_9920,N_9041);
or UO_876 (O_876,N_9600,N_9009);
nor UO_877 (O_877,N_9725,N_9942);
nand UO_878 (O_878,N_9871,N_9972);
or UO_879 (O_879,N_9390,N_9376);
or UO_880 (O_880,N_9657,N_9621);
nand UO_881 (O_881,N_9688,N_9607);
or UO_882 (O_882,N_9179,N_9424);
or UO_883 (O_883,N_9977,N_9517);
and UO_884 (O_884,N_9431,N_9556);
nor UO_885 (O_885,N_9018,N_9562);
or UO_886 (O_886,N_9886,N_9944);
or UO_887 (O_887,N_9299,N_9911);
nor UO_888 (O_888,N_9818,N_9155);
nand UO_889 (O_889,N_9387,N_9259);
and UO_890 (O_890,N_9071,N_9622);
nor UO_891 (O_891,N_9038,N_9904);
nor UO_892 (O_892,N_9419,N_9963);
nor UO_893 (O_893,N_9811,N_9004);
and UO_894 (O_894,N_9640,N_9491);
xnor UO_895 (O_895,N_9859,N_9071);
and UO_896 (O_896,N_9649,N_9970);
nor UO_897 (O_897,N_9054,N_9916);
nand UO_898 (O_898,N_9773,N_9320);
nor UO_899 (O_899,N_9146,N_9915);
or UO_900 (O_900,N_9836,N_9517);
or UO_901 (O_901,N_9955,N_9878);
nand UO_902 (O_902,N_9823,N_9284);
nor UO_903 (O_903,N_9590,N_9323);
or UO_904 (O_904,N_9944,N_9170);
and UO_905 (O_905,N_9510,N_9912);
nor UO_906 (O_906,N_9572,N_9825);
or UO_907 (O_907,N_9369,N_9440);
nor UO_908 (O_908,N_9797,N_9039);
or UO_909 (O_909,N_9580,N_9246);
nor UO_910 (O_910,N_9157,N_9731);
and UO_911 (O_911,N_9877,N_9644);
or UO_912 (O_912,N_9621,N_9458);
or UO_913 (O_913,N_9507,N_9996);
and UO_914 (O_914,N_9571,N_9170);
nor UO_915 (O_915,N_9764,N_9796);
nand UO_916 (O_916,N_9360,N_9712);
nand UO_917 (O_917,N_9276,N_9438);
nor UO_918 (O_918,N_9756,N_9010);
nand UO_919 (O_919,N_9322,N_9881);
and UO_920 (O_920,N_9704,N_9291);
nand UO_921 (O_921,N_9691,N_9788);
and UO_922 (O_922,N_9889,N_9159);
nor UO_923 (O_923,N_9141,N_9394);
and UO_924 (O_924,N_9521,N_9906);
nor UO_925 (O_925,N_9519,N_9768);
nor UO_926 (O_926,N_9946,N_9534);
xor UO_927 (O_927,N_9468,N_9911);
and UO_928 (O_928,N_9292,N_9872);
nor UO_929 (O_929,N_9299,N_9848);
nand UO_930 (O_930,N_9761,N_9034);
nor UO_931 (O_931,N_9619,N_9049);
nor UO_932 (O_932,N_9320,N_9205);
nand UO_933 (O_933,N_9363,N_9581);
and UO_934 (O_934,N_9625,N_9491);
or UO_935 (O_935,N_9391,N_9200);
nand UO_936 (O_936,N_9954,N_9652);
nor UO_937 (O_937,N_9447,N_9399);
nand UO_938 (O_938,N_9026,N_9456);
and UO_939 (O_939,N_9256,N_9674);
and UO_940 (O_940,N_9964,N_9701);
and UO_941 (O_941,N_9133,N_9630);
and UO_942 (O_942,N_9201,N_9857);
nand UO_943 (O_943,N_9127,N_9677);
nor UO_944 (O_944,N_9527,N_9558);
nand UO_945 (O_945,N_9630,N_9716);
xor UO_946 (O_946,N_9038,N_9435);
nor UO_947 (O_947,N_9109,N_9562);
nor UO_948 (O_948,N_9462,N_9150);
nand UO_949 (O_949,N_9335,N_9359);
nand UO_950 (O_950,N_9557,N_9772);
and UO_951 (O_951,N_9421,N_9415);
and UO_952 (O_952,N_9271,N_9477);
nor UO_953 (O_953,N_9139,N_9105);
and UO_954 (O_954,N_9126,N_9778);
nor UO_955 (O_955,N_9213,N_9623);
or UO_956 (O_956,N_9474,N_9096);
or UO_957 (O_957,N_9769,N_9647);
or UO_958 (O_958,N_9620,N_9965);
or UO_959 (O_959,N_9464,N_9639);
and UO_960 (O_960,N_9433,N_9904);
nor UO_961 (O_961,N_9794,N_9820);
and UO_962 (O_962,N_9714,N_9770);
nor UO_963 (O_963,N_9365,N_9112);
nor UO_964 (O_964,N_9288,N_9857);
or UO_965 (O_965,N_9843,N_9049);
and UO_966 (O_966,N_9969,N_9168);
and UO_967 (O_967,N_9328,N_9007);
and UO_968 (O_968,N_9114,N_9392);
nand UO_969 (O_969,N_9807,N_9399);
and UO_970 (O_970,N_9642,N_9783);
and UO_971 (O_971,N_9816,N_9531);
nand UO_972 (O_972,N_9487,N_9101);
or UO_973 (O_973,N_9583,N_9341);
or UO_974 (O_974,N_9290,N_9187);
nor UO_975 (O_975,N_9648,N_9039);
nand UO_976 (O_976,N_9931,N_9447);
and UO_977 (O_977,N_9159,N_9258);
nand UO_978 (O_978,N_9810,N_9754);
and UO_979 (O_979,N_9925,N_9542);
and UO_980 (O_980,N_9848,N_9653);
nor UO_981 (O_981,N_9405,N_9051);
nand UO_982 (O_982,N_9273,N_9054);
or UO_983 (O_983,N_9345,N_9071);
nand UO_984 (O_984,N_9591,N_9837);
and UO_985 (O_985,N_9927,N_9799);
and UO_986 (O_986,N_9087,N_9512);
or UO_987 (O_987,N_9199,N_9636);
nor UO_988 (O_988,N_9306,N_9560);
nand UO_989 (O_989,N_9384,N_9148);
or UO_990 (O_990,N_9835,N_9903);
and UO_991 (O_991,N_9224,N_9359);
and UO_992 (O_992,N_9140,N_9692);
nor UO_993 (O_993,N_9465,N_9259);
or UO_994 (O_994,N_9932,N_9608);
or UO_995 (O_995,N_9168,N_9968);
nand UO_996 (O_996,N_9485,N_9608);
nand UO_997 (O_997,N_9619,N_9426);
xor UO_998 (O_998,N_9150,N_9191);
and UO_999 (O_999,N_9327,N_9012);
nand UO_1000 (O_1000,N_9010,N_9558);
nor UO_1001 (O_1001,N_9700,N_9426);
nor UO_1002 (O_1002,N_9494,N_9889);
nand UO_1003 (O_1003,N_9163,N_9239);
nor UO_1004 (O_1004,N_9035,N_9369);
or UO_1005 (O_1005,N_9106,N_9769);
nor UO_1006 (O_1006,N_9924,N_9152);
nor UO_1007 (O_1007,N_9930,N_9378);
or UO_1008 (O_1008,N_9037,N_9244);
or UO_1009 (O_1009,N_9804,N_9143);
or UO_1010 (O_1010,N_9618,N_9270);
xnor UO_1011 (O_1011,N_9364,N_9183);
nand UO_1012 (O_1012,N_9381,N_9254);
nor UO_1013 (O_1013,N_9014,N_9281);
or UO_1014 (O_1014,N_9797,N_9421);
nand UO_1015 (O_1015,N_9702,N_9833);
nor UO_1016 (O_1016,N_9210,N_9470);
nor UO_1017 (O_1017,N_9117,N_9362);
or UO_1018 (O_1018,N_9904,N_9264);
nor UO_1019 (O_1019,N_9849,N_9520);
nand UO_1020 (O_1020,N_9712,N_9395);
or UO_1021 (O_1021,N_9852,N_9690);
nor UO_1022 (O_1022,N_9714,N_9582);
or UO_1023 (O_1023,N_9257,N_9741);
and UO_1024 (O_1024,N_9845,N_9529);
nor UO_1025 (O_1025,N_9461,N_9657);
or UO_1026 (O_1026,N_9803,N_9979);
nand UO_1027 (O_1027,N_9965,N_9670);
nor UO_1028 (O_1028,N_9550,N_9741);
nor UO_1029 (O_1029,N_9412,N_9193);
nand UO_1030 (O_1030,N_9451,N_9273);
or UO_1031 (O_1031,N_9060,N_9537);
nand UO_1032 (O_1032,N_9702,N_9817);
nand UO_1033 (O_1033,N_9283,N_9174);
nand UO_1034 (O_1034,N_9144,N_9976);
and UO_1035 (O_1035,N_9923,N_9026);
or UO_1036 (O_1036,N_9289,N_9322);
or UO_1037 (O_1037,N_9171,N_9636);
nand UO_1038 (O_1038,N_9853,N_9578);
nand UO_1039 (O_1039,N_9407,N_9782);
nor UO_1040 (O_1040,N_9129,N_9366);
nand UO_1041 (O_1041,N_9873,N_9699);
or UO_1042 (O_1042,N_9989,N_9899);
nand UO_1043 (O_1043,N_9135,N_9156);
nor UO_1044 (O_1044,N_9795,N_9912);
or UO_1045 (O_1045,N_9579,N_9510);
or UO_1046 (O_1046,N_9096,N_9862);
and UO_1047 (O_1047,N_9672,N_9873);
nor UO_1048 (O_1048,N_9777,N_9124);
nand UO_1049 (O_1049,N_9053,N_9422);
or UO_1050 (O_1050,N_9045,N_9217);
nand UO_1051 (O_1051,N_9173,N_9015);
or UO_1052 (O_1052,N_9916,N_9313);
or UO_1053 (O_1053,N_9788,N_9182);
and UO_1054 (O_1054,N_9085,N_9059);
and UO_1055 (O_1055,N_9135,N_9716);
and UO_1056 (O_1056,N_9329,N_9263);
nor UO_1057 (O_1057,N_9487,N_9752);
nor UO_1058 (O_1058,N_9817,N_9063);
and UO_1059 (O_1059,N_9441,N_9271);
nand UO_1060 (O_1060,N_9785,N_9092);
and UO_1061 (O_1061,N_9719,N_9953);
nor UO_1062 (O_1062,N_9309,N_9903);
or UO_1063 (O_1063,N_9517,N_9704);
or UO_1064 (O_1064,N_9126,N_9070);
or UO_1065 (O_1065,N_9699,N_9673);
or UO_1066 (O_1066,N_9143,N_9533);
or UO_1067 (O_1067,N_9075,N_9996);
and UO_1068 (O_1068,N_9821,N_9455);
nor UO_1069 (O_1069,N_9945,N_9726);
and UO_1070 (O_1070,N_9725,N_9322);
nand UO_1071 (O_1071,N_9147,N_9301);
nor UO_1072 (O_1072,N_9633,N_9790);
nor UO_1073 (O_1073,N_9625,N_9303);
nand UO_1074 (O_1074,N_9262,N_9027);
or UO_1075 (O_1075,N_9996,N_9960);
and UO_1076 (O_1076,N_9462,N_9211);
nand UO_1077 (O_1077,N_9089,N_9327);
nand UO_1078 (O_1078,N_9342,N_9517);
nor UO_1079 (O_1079,N_9271,N_9812);
and UO_1080 (O_1080,N_9588,N_9520);
or UO_1081 (O_1081,N_9337,N_9772);
nand UO_1082 (O_1082,N_9875,N_9622);
nor UO_1083 (O_1083,N_9404,N_9229);
nor UO_1084 (O_1084,N_9342,N_9808);
nor UO_1085 (O_1085,N_9296,N_9731);
nor UO_1086 (O_1086,N_9475,N_9060);
and UO_1087 (O_1087,N_9141,N_9756);
nor UO_1088 (O_1088,N_9277,N_9914);
xnor UO_1089 (O_1089,N_9312,N_9598);
nand UO_1090 (O_1090,N_9946,N_9169);
nor UO_1091 (O_1091,N_9389,N_9326);
nand UO_1092 (O_1092,N_9505,N_9878);
nand UO_1093 (O_1093,N_9716,N_9809);
xnor UO_1094 (O_1094,N_9028,N_9275);
and UO_1095 (O_1095,N_9693,N_9139);
nand UO_1096 (O_1096,N_9589,N_9756);
nor UO_1097 (O_1097,N_9603,N_9541);
and UO_1098 (O_1098,N_9859,N_9801);
or UO_1099 (O_1099,N_9461,N_9042);
nand UO_1100 (O_1100,N_9512,N_9452);
or UO_1101 (O_1101,N_9659,N_9712);
nor UO_1102 (O_1102,N_9273,N_9721);
nor UO_1103 (O_1103,N_9839,N_9069);
nand UO_1104 (O_1104,N_9954,N_9126);
or UO_1105 (O_1105,N_9438,N_9919);
and UO_1106 (O_1106,N_9681,N_9823);
nand UO_1107 (O_1107,N_9070,N_9688);
or UO_1108 (O_1108,N_9416,N_9537);
xnor UO_1109 (O_1109,N_9800,N_9462);
nor UO_1110 (O_1110,N_9493,N_9142);
nor UO_1111 (O_1111,N_9576,N_9254);
nand UO_1112 (O_1112,N_9945,N_9573);
and UO_1113 (O_1113,N_9666,N_9213);
and UO_1114 (O_1114,N_9421,N_9358);
or UO_1115 (O_1115,N_9262,N_9860);
or UO_1116 (O_1116,N_9649,N_9245);
nand UO_1117 (O_1117,N_9656,N_9125);
and UO_1118 (O_1118,N_9216,N_9781);
nor UO_1119 (O_1119,N_9080,N_9875);
nand UO_1120 (O_1120,N_9523,N_9781);
nand UO_1121 (O_1121,N_9573,N_9427);
nor UO_1122 (O_1122,N_9441,N_9414);
and UO_1123 (O_1123,N_9465,N_9601);
nor UO_1124 (O_1124,N_9216,N_9117);
and UO_1125 (O_1125,N_9434,N_9786);
nand UO_1126 (O_1126,N_9000,N_9952);
or UO_1127 (O_1127,N_9845,N_9414);
or UO_1128 (O_1128,N_9615,N_9954);
nor UO_1129 (O_1129,N_9605,N_9521);
and UO_1130 (O_1130,N_9012,N_9330);
nand UO_1131 (O_1131,N_9890,N_9608);
nand UO_1132 (O_1132,N_9140,N_9350);
nand UO_1133 (O_1133,N_9441,N_9530);
and UO_1134 (O_1134,N_9122,N_9229);
or UO_1135 (O_1135,N_9807,N_9571);
and UO_1136 (O_1136,N_9441,N_9187);
or UO_1137 (O_1137,N_9658,N_9964);
and UO_1138 (O_1138,N_9392,N_9678);
nand UO_1139 (O_1139,N_9008,N_9537);
nand UO_1140 (O_1140,N_9533,N_9262);
or UO_1141 (O_1141,N_9072,N_9321);
and UO_1142 (O_1142,N_9505,N_9097);
nand UO_1143 (O_1143,N_9530,N_9231);
nand UO_1144 (O_1144,N_9399,N_9749);
nand UO_1145 (O_1145,N_9014,N_9498);
nor UO_1146 (O_1146,N_9690,N_9525);
or UO_1147 (O_1147,N_9359,N_9008);
nand UO_1148 (O_1148,N_9631,N_9626);
or UO_1149 (O_1149,N_9428,N_9868);
or UO_1150 (O_1150,N_9937,N_9044);
nor UO_1151 (O_1151,N_9584,N_9201);
and UO_1152 (O_1152,N_9965,N_9346);
nand UO_1153 (O_1153,N_9908,N_9665);
or UO_1154 (O_1154,N_9370,N_9052);
nor UO_1155 (O_1155,N_9538,N_9472);
nor UO_1156 (O_1156,N_9689,N_9359);
or UO_1157 (O_1157,N_9715,N_9852);
nor UO_1158 (O_1158,N_9100,N_9751);
nor UO_1159 (O_1159,N_9237,N_9484);
or UO_1160 (O_1160,N_9879,N_9402);
nor UO_1161 (O_1161,N_9492,N_9151);
and UO_1162 (O_1162,N_9419,N_9403);
or UO_1163 (O_1163,N_9903,N_9974);
nand UO_1164 (O_1164,N_9978,N_9228);
and UO_1165 (O_1165,N_9842,N_9122);
nor UO_1166 (O_1166,N_9420,N_9235);
nor UO_1167 (O_1167,N_9402,N_9154);
or UO_1168 (O_1168,N_9075,N_9365);
nor UO_1169 (O_1169,N_9619,N_9670);
nor UO_1170 (O_1170,N_9207,N_9346);
nand UO_1171 (O_1171,N_9201,N_9902);
and UO_1172 (O_1172,N_9769,N_9800);
and UO_1173 (O_1173,N_9778,N_9500);
nand UO_1174 (O_1174,N_9067,N_9632);
or UO_1175 (O_1175,N_9828,N_9691);
nand UO_1176 (O_1176,N_9789,N_9512);
nor UO_1177 (O_1177,N_9313,N_9610);
nor UO_1178 (O_1178,N_9171,N_9210);
and UO_1179 (O_1179,N_9463,N_9496);
and UO_1180 (O_1180,N_9492,N_9287);
nor UO_1181 (O_1181,N_9396,N_9441);
nor UO_1182 (O_1182,N_9204,N_9045);
nand UO_1183 (O_1183,N_9030,N_9366);
nand UO_1184 (O_1184,N_9203,N_9095);
nand UO_1185 (O_1185,N_9498,N_9928);
nor UO_1186 (O_1186,N_9182,N_9262);
and UO_1187 (O_1187,N_9905,N_9932);
and UO_1188 (O_1188,N_9261,N_9841);
nand UO_1189 (O_1189,N_9533,N_9477);
and UO_1190 (O_1190,N_9506,N_9606);
and UO_1191 (O_1191,N_9959,N_9559);
nor UO_1192 (O_1192,N_9925,N_9555);
nor UO_1193 (O_1193,N_9425,N_9095);
nand UO_1194 (O_1194,N_9413,N_9056);
nor UO_1195 (O_1195,N_9473,N_9166);
nand UO_1196 (O_1196,N_9674,N_9787);
and UO_1197 (O_1197,N_9919,N_9710);
or UO_1198 (O_1198,N_9461,N_9370);
nand UO_1199 (O_1199,N_9617,N_9358);
or UO_1200 (O_1200,N_9838,N_9678);
nand UO_1201 (O_1201,N_9714,N_9008);
xor UO_1202 (O_1202,N_9242,N_9550);
nand UO_1203 (O_1203,N_9458,N_9225);
and UO_1204 (O_1204,N_9726,N_9078);
nor UO_1205 (O_1205,N_9977,N_9615);
and UO_1206 (O_1206,N_9733,N_9559);
or UO_1207 (O_1207,N_9094,N_9233);
and UO_1208 (O_1208,N_9260,N_9126);
or UO_1209 (O_1209,N_9278,N_9139);
nor UO_1210 (O_1210,N_9686,N_9198);
and UO_1211 (O_1211,N_9751,N_9819);
nand UO_1212 (O_1212,N_9581,N_9587);
and UO_1213 (O_1213,N_9722,N_9263);
nand UO_1214 (O_1214,N_9457,N_9227);
nand UO_1215 (O_1215,N_9020,N_9887);
nand UO_1216 (O_1216,N_9394,N_9119);
and UO_1217 (O_1217,N_9973,N_9560);
nand UO_1218 (O_1218,N_9306,N_9545);
or UO_1219 (O_1219,N_9393,N_9849);
and UO_1220 (O_1220,N_9076,N_9147);
nor UO_1221 (O_1221,N_9928,N_9737);
nand UO_1222 (O_1222,N_9760,N_9719);
and UO_1223 (O_1223,N_9133,N_9304);
nor UO_1224 (O_1224,N_9349,N_9976);
and UO_1225 (O_1225,N_9981,N_9360);
nor UO_1226 (O_1226,N_9399,N_9692);
nand UO_1227 (O_1227,N_9780,N_9675);
nand UO_1228 (O_1228,N_9748,N_9112);
nor UO_1229 (O_1229,N_9779,N_9543);
nand UO_1230 (O_1230,N_9948,N_9642);
nor UO_1231 (O_1231,N_9061,N_9047);
nand UO_1232 (O_1232,N_9946,N_9045);
nor UO_1233 (O_1233,N_9599,N_9976);
or UO_1234 (O_1234,N_9806,N_9196);
nand UO_1235 (O_1235,N_9796,N_9705);
nor UO_1236 (O_1236,N_9597,N_9576);
nor UO_1237 (O_1237,N_9728,N_9109);
and UO_1238 (O_1238,N_9417,N_9657);
or UO_1239 (O_1239,N_9096,N_9895);
nand UO_1240 (O_1240,N_9061,N_9211);
or UO_1241 (O_1241,N_9951,N_9873);
nor UO_1242 (O_1242,N_9240,N_9379);
nand UO_1243 (O_1243,N_9241,N_9894);
and UO_1244 (O_1244,N_9001,N_9451);
or UO_1245 (O_1245,N_9811,N_9821);
nor UO_1246 (O_1246,N_9422,N_9154);
nand UO_1247 (O_1247,N_9959,N_9129);
or UO_1248 (O_1248,N_9281,N_9852);
or UO_1249 (O_1249,N_9427,N_9484);
or UO_1250 (O_1250,N_9104,N_9296);
and UO_1251 (O_1251,N_9615,N_9264);
nor UO_1252 (O_1252,N_9857,N_9343);
nor UO_1253 (O_1253,N_9666,N_9221);
and UO_1254 (O_1254,N_9799,N_9177);
nor UO_1255 (O_1255,N_9755,N_9498);
or UO_1256 (O_1256,N_9210,N_9602);
and UO_1257 (O_1257,N_9196,N_9488);
and UO_1258 (O_1258,N_9084,N_9293);
or UO_1259 (O_1259,N_9474,N_9978);
nand UO_1260 (O_1260,N_9319,N_9787);
and UO_1261 (O_1261,N_9564,N_9302);
and UO_1262 (O_1262,N_9136,N_9016);
or UO_1263 (O_1263,N_9997,N_9043);
nor UO_1264 (O_1264,N_9601,N_9287);
nor UO_1265 (O_1265,N_9604,N_9886);
or UO_1266 (O_1266,N_9648,N_9056);
or UO_1267 (O_1267,N_9466,N_9784);
and UO_1268 (O_1268,N_9219,N_9485);
and UO_1269 (O_1269,N_9694,N_9033);
and UO_1270 (O_1270,N_9459,N_9582);
nor UO_1271 (O_1271,N_9946,N_9254);
nand UO_1272 (O_1272,N_9809,N_9921);
and UO_1273 (O_1273,N_9391,N_9293);
or UO_1274 (O_1274,N_9485,N_9356);
or UO_1275 (O_1275,N_9716,N_9718);
and UO_1276 (O_1276,N_9973,N_9292);
nor UO_1277 (O_1277,N_9779,N_9178);
nand UO_1278 (O_1278,N_9013,N_9284);
or UO_1279 (O_1279,N_9073,N_9660);
nand UO_1280 (O_1280,N_9738,N_9853);
nand UO_1281 (O_1281,N_9782,N_9180);
or UO_1282 (O_1282,N_9188,N_9240);
or UO_1283 (O_1283,N_9942,N_9471);
nand UO_1284 (O_1284,N_9815,N_9635);
and UO_1285 (O_1285,N_9318,N_9717);
nor UO_1286 (O_1286,N_9348,N_9784);
or UO_1287 (O_1287,N_9677,N_9730);
nor UO_1288 (O_1288,N_9191,N_9141);
or UO_1289 (O_1289,N_9642,N_9131);
or UO_1290 (O_1290,N_9263,N_9746);
nor UO_1291 (O_1291,N_9091,N_9171);
and UO_1292 (O_1292,N_9647,N_9424);
nor UO_1293 (O_1293,N_9112,N_9695);
and UO_1294 (O_1294,N_9062,N_9320);
and UO_1295 (O_1295,N_9238,N_9230);
and UO_1296 (O_1296,N_9995,N_9198);
or UO_1297 (O_1297,N_9616,N_9783);
and UO_1298 (O_1298,N_9773,N_9499);
and UO_1299 (O_1299,N_9990,N_9069);
nand UO_1300 (O_1300,N_9026,N_9077);
or UO_1301 (O_1301,N_9177,N_9481);
and UO_1302 (O_1302,N_9565,N_9538);
or UO_1303 (O_1303,N_9638,N_9454);
nand UO_1304 (O_1304,N_9661,N_9314);
nand UO_1305 (O_1305,N_9177,N_9035);
nor UO_1306 (O_1306,N_9122,N_9939);
or UO_1307 (O_1307,N_9431,N_9687);
nor UO_1308 (O_1308,N_9132,N_9426);
or UO_1309 (O_1309,N_9155,N_9524);
nor UO_1310 (O_1310,N_9742,N_9729);
or UO_1311 (O_1311,N_9769,N_9045);
nor UO_1312 (O_1312,N_9265,N_9493);
or UO_1313 (O_1313,N_9867,N_9934);
or UO_1314 (O_1314,N_9597,N_9695);
and UO_1315 (O_1315,N_9614,N_9063);
and UO_1316 (O_1316,N_9458,N_9876);
nor UO_1317 (O_1317,N_9165,N_9541);
nand UO_1318 (O_1318,N_9758,N_9414);
and UO_1319 (O_1319,N_9315,N_9525);
or UO_1320 (O_1320,N_9101,N_9608);
xnor UO_1321 (O_1321,N_9994,N_9907);
and UO_1322 (O_1322,N_9345,N_9748);
nand UO_1323 (O_1323,N_9827,N_9859);
nor UO_1324 (O_1324,N_9725,N_9527);
and UO_1325 (O_1325,N_9331,N_9367);
and UO_1326 (O_1326,N_9637,N_9876);
or UO_1327 (O_1327,N_9225,N_9049);
nor UO_1328 (O_1328,N_9071,N_9872);
or UO_1329 (O_1329,N_9870,N_9082);
and UO_1330 (O_1330,N_9955,N_9325);
nor UO_1331 (O_1331,N_9459,N_9378);
and UO_1332 (O_1332,N_9058,N_9945);
nand UO_1333 (O_1333,N_9133,N_9477);
or UO_1334 (O_1334,N_9519,N_9499);
nor UO_1335 (O_1335,N_9298,N_9554);
and UO_1336 (O_1336,N_9326,N_9886);
or UO_1337 (O_1337,N_9614,N_9578);
nand UO_1338 (O_1338,N_9490,N_9489);
nand UO_1339 (O_1339,N_9286,N_9388);
or UO_1340 (O_1340,N_9929,N_9693);
and UO_1341 (O_1341,N_9252,N_9485);
or UO_1342 (O_1342,N_9477,N_9361);
or UO_1343 (O_1343,N_9815,N_9769);
nand UO_1344 (O_1344,N_9857,N_9599);
or UO_1345 (O_1345,N_9352,N_9083);
or UO_1346 (O_1346,N_9619,N_9061);
nand UO_1347 (O_1347,N_9567,N_9610);
and UO_1348 (O_1348,N_9696,N_9757);
or UO_1349 (O_1349,N_9738,N_9543);
and UO_1350 (O_1350,N_9216,N_9875);
nand UO_1351 (O_1351,N_9463,N_9296);
or UO_1352 (O_1352,N_9987,N_9181);
or UO_1353 (O_1353,N_9178,N_9364);
and UO_1354 (O_1354,N_9495,N_9040);
nand UO_1355 (O_1355,N_9729,N_9454);
or UO_1356 (O_1356,N_9345,N_9751);
or UO_1357 (O_1357,N_9973,N_9582);
or UO_1358 (O_1358,N_9628,N_9083);
nor UO_1359 (O_1359,N_9444,N_9869);
and UO_1360 (O_1360,N_9034,N_9234);
nor UO_1361 (O_1361,N_9315,N_9584);
and UO_1362 (O_1362,N_9930,N_9276);
and UO_1363 (O_1363,N_9837,N_9404);
nor UO_1364 (O_1364,N_9851,N_9709);
or UO_1365 (O_1365,N_9351,N_9154);
and UO_1366 (O_1366,N_9327,N_9021);
nor UO_1367 (O_1367,N_9307,N_9134);
nor UO_1368 (O_1368,N_9338,N_9476);
or UO_1369 (O_1369,N_9240,N_9124);
or UO_1370 (O_1370,N_9264,N_9962);
and UO_1371 (O_1371,N_9347,N_9991);
nor UO_1372 (O_1372,N_9816,N_9433);
and UO_1373 (O_1373,N_9491,N_9817);
and UO_1374 (O_1374,N_9540,N_9118);
and UO_1375 (O_1375,N_9327,N_9957);
or UO_1376 (O_1376,N_9681,N_9118);
nand UO_1377 (O_1377,N_9213,N_9401);
or UO_1378 (O_1378,N_9146,N_9653);
or UO_1379 (O_1379,N_9145,N_9515);
nor UO_1380 (O_1380,N_9148,N_9132);
nand UO_1381 (O_1381,N_9532,N_9335);
and UO_1382 (O_1382,N_9451,N_9757);
and UO_1383 (O_1383,N_9295,N_9684);
nand UO_1384 (O_1384,N_9139,N_9455);
nor UO_1385 (O_1385,N_9143,N_9793);
or UO_1386 (O_1386,N_9792,N_9322);
and UO_1387 (O_1387,N_9396,N_9159);
nand UO_1388 (O_1388,N_9269,N_9872);
or UO_1389 (O_1389,N_9347,N_9415);
or UO_1390 (O_1390,N_9346,N_9108);
and UO_1391 (O_1391,N_9683,N_9235);
nor UO_1392 (O_1392,N_9268,N_9281);
nand UO_1393 (O_1393,N_9737,N_9005);
and UO_1394 (O_1394,N_9119,N_9387);
or UO_1395 (O_1395,N_9979,N_9380);
or UO_1396 (O_1396,N_9603,N_9906);
nor UO_1397 (O_1397,N_9908,N_9599);
or UO_1398 (O_1398,N_9791,N_9723);
and UO_1399 (O_1399,N_9284,N_9489);
or UO_1400 (O_1400,N_9541,N_9533);
or UO_1401 (O_1401,N_9762,N_9661);
and UO_1402 (O_1402,N_9296,N_9804);
or UO_1403 (O_1403,N_9778,N_9909);
and UO_1404 (O_1404,N_9349,N_9187);
or UO_1405 (O_1405,N_9781,N_9047);
nand UO_1406 (O_1406,N_9629,N_9804);
or UO_1407 (O_1407,N_9948,N_9863);
nand UO_1408 (O_1408,N_9285,N_9949);
nor UO_1409 (O_1409,N_9025,N_9249);
and UO_1410 (O_1410,N_9924,N_9720);
or UO_1411 (O_1411,N_9102,N_9617);
or UO_1412 (O_1412,N_9268,N_9527);
nand UO_1413 (O_1413,N_9583,N_9028);
or UO_1414 (O_1414,N_9543,N_9472);
and UO_1415 (O_1415,N_9747,N_9834);
nor UO_1416 (O_1416,N_9240,N_9641);
and UO_1417 (O_1417,N_9508,N_9733);
nand UO_1418 (O_1418,N_9524,N_9944);
nor UO_1419 (O_1419,N_9479,N_9170);
nand UO_1420 (O_1420,N_9817,N_9856);
nand UO_1421 (O_1421,N_9711,N_9699);
nor UO_1422 (O_1422,N_9882,N_9090);
nor UO_1423 (O_1423,N_9302,N_9582);
or UO_1424 (O_1424,N_9907,N_9320);
nor UO_1425 (O_1425,N_9283,N_9890);
nor UO_1426 (O_1426,N_9456,N_9431);
nand UO_1427 (O_1427,N_9674,N_9406);
or UO_1428 (O_1428,N_9283,N_9041);
xnor UO_1429 (O_1429,N_9685,N_9314);
nor UO_1430 (O_1430,N_9144,N_9859);
nor UO_1431 (O_1431,N_9242,N_9310);
nor UO_1432 (O_1432,N_9852,N_9696);
or UO_1433 (O_1433,N_9757,N_9687);
and UO_1434 (O_1434,N_9122,N_9950);
and UO_1435 (O_1435,N_9963,N_9028);
and UO_1436 (O_1436,N_9762,N_9409);
nor UO_1437 (O_1437,N_9837,N_9823);
nor UO_1438 (O_1438,N_9484,N_9324);
and UO_1439 (O_1439,N_9760,N_9374);
and UO_1440 (O_1440,N_9436,N_9054);
nor UO_1441 (O_1441,N_9812,N_9879);
and UO_1442 (O_1442,N_9485,N_9456);
or UO_1443 (O_1443,N_9567,N_9509);
and UO_1444 (O_1444,N_9529,N_9353);
and UO_1445 (O_1445,N_9301,N_9351);
nand UO_1446 (O_1446,N_9734,N_9048);
nand UO_1447 (O_1447,N_9499,N_9131);
nand UO_1448 (O_1448,N_9062,N_9113);
or UO_1449 (O_1449,N_9212,N_9097);
nand UO_1450 (O_1450,N_9448,N_9036);
nand UO_1451 (O_1451,N_9352,N_9707);
nand UO_1452 (O_1452,N_9237,N_9994);
nand UO_1453 (O_1453,N_9240,N_9504);
nor UO_1454 (O_1454,N_9728,N_9749);
or UO_1455 (O_1455,N_9872,N_9615);
and UO_1456 (O_1456,N_9218,N_9766);
or UO_1457 (O_1457,N_9601,N_9099);
nand UO_1458 (O_1458,N_9400,N_9068);
or UO_1459 (O_1459,N_9073,N_9726);
or UO_1460 (O_1460,N_9760,N_9526);
and UO_1461 (O_1461,N_9058,N_9770);
nor UO_1462 (O_1462,N_9485,N_9040);
xor UO_1463 (O_1463,N_9545,N_9792);
nand UO_1464 (O_1464,N_9747,N_9174);
or UO_1465 (O_1465,N_9535,N_9361);
nor UO_1466 (O_1466,N_9561,N_9938);
or UO_1467 (O_1467,N_9315,N_9220);
nand UO_1468 (O_1468,N_9744,N_9395);
and UO_1469 (O_1469,N_9692,N_9596);
or UO_1470 (O_1470,N_9495,N_9821);
and UO_1471 (O_1471,N_9900,N_9057);
or UO_1472 (O_1472,N_9200,N_9245);
nand UO_1473 (O_1473,N_9438,N_9738);
nor UO_1474 (O_1474,N_9664,N_9501);
and UO_1475 (O_1475,N_9259,N_9109);
or UO_1476 (O_1476,N_9119,N_9876);
or UO_1477 (O_1477,N_9898,N_9532);
nor UO_1478 (O_1478,N_9800,N_9988);
nand UO_1479 (O_1479,N_9240,N_9995);
nand UO_1480 (O_1480,N_9853,N_9334);
and UO_1481 (O_1481,N_9304,N_9618);
and UO_1482 (O_1482,N_9475,N_9463);
nand UO_1483 (O_1483,N_9920,N_9535);
and UO_1484 (O_1484,N_9910,N_9623);
and UO_1485 (O_1485,N_9455,N_9642);
nor UO_1486 (O_1486,N_9315,N_9340);
or UO_1487 (O_1487,N_9551,N_9224);
nor UO_1488 (O_1488,N_9533,N_9616);
nand UO_1489 (O_1489,N_9037,N_9851);
nor UO_1490 (O_1490,N_9005,N_9773);
nor UO_1491 (O_1491,N_9580,N_9067);
nor UO_1492 (O_1492,N_9144,N_9704);
or UO_1493 (O_1493,N_9510,N_9948);
or UO_1494 (O_1494,N_9627,N_9933);
or UO_1495 (O_1495,N_9781,N_9818);
and UO_1496 (O_1496,N_9280,N_9346);
nor UO_1497 (O_1497,N_9474,N_9358);
nand UO_1498 (O_1498,N_9625,N_9589);
and UO_1499 (O_1499,N_9554,N_9879);
endmodule