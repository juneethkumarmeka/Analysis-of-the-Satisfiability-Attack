module basic_750_5000_1000_10_levels_2xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
and U0 (N_0,In_596,In_726);
or U1 (N_1,In_64,In_406);
nor U2 (N_2,In_656,In_706);
or U3 (N_3,In_649,In_164);
or U4 (N_4,In_683,In_542);
and U5 (N_5,In_432,In_90);
nor U6 (N_6,In_484,In_343);
nand U7 (N_7,In_518,In_268);
nor U8 (N_8,In_203,In_18);
or U9 (N_9,In_492,In_326);
xor U10 (N_10,In_449,In_208);
nor U11 (N_11,In_462,In_604);
nand U12 (N_12,In_737,In_503);
xnor U13 (N_13,In_357,In_283);
nor U14 (N_14,In_354,In_516);
or U15 (N_15,In_332,In_273);
nor U16 (N_16,In_439,In_337);
nand U17 (N_17,In_426,In_393);
nor U18 (N_18,In_670,In_468);
and U19 (N_19,In_317,In_544);
nor U20 (N_20,In_188,In_504);
nor U21 (N_21,In_632,In_315);
nor U22 (N_22,In_733,In_394);
and U23 (N_23,In_240,In_392);
or U24 (N_24,In_689,In_586);
or U25 (N_25,In_366,In_175);
nand U26 (N_26,In_299,In_230);
nor U27 (N_27,In_271,In_150);
and U28 (N_28,In_454,In_385);
or U29 (N_29,In_697,In_42);
nor U30 (N_30,In_154,In_163);
nor U31 (N_31,In_75,In_94);
or U32 (N_32,In_7,In_641);
nor U33 (N_33,In_585,In_118);
or U34 (N_34,In_571,In_251);
nand U35 (N_35,In_651,In_113);
or U36 (N_36,In_309,In_265);
xor U37 (N_37,In_704,In_573);
or U38 (N_38,In_347,In_124);
nor U39 (N_39,In_3,In_691);
and U40 (N_40,In_471,In_184);
nor U41 (N_41,In_27,In_625);
or U42 (N_42,In_535,In_609);
nand U43 (N_43,In_555,In_517);
or U44 (N_44,In_146,In_145);
nor U45 (N_45,In_296,In_568);
nor U46 (N_46,In_16,In_152);
nor U47 (N_47,In_636,In_436);
or U48 (N_48,In_681,In_721);
nand U49 (N_49,In_287,In_14);
nor U50 (N_50,In_156,In_738);
nand U51 (N_51,In_709,In_615);
and U52 (N_52,In_143,In_565);
and U53 (N_53,In_358,In_532);
nand U54 (N_54,In_493,In_618);
nand U55 (N_55,In_576,In_599);
and U56 (N_56,In_639,In_664);
or U57 (N_57,In_458,In_659);
or U58 (N_58,In_82,In_252);
nor U59 (N_59,In_375,In_259);
or U60 (N_60,In_226,In_258);
or U61 (N_61,In_212,In_266);
and U62 (N_62,In_74,In_291);
nor U63 (N_63,In_514,In_144);
or U64 (N_64,In_215,In_102);
nand U65 (N_65,In_80,In_229);
nor U66 (N_66,In_86,In_658);
nand U67 (N_67,In_54,In_151);
nand U68 (N_68,In_421,In_340);
or U69 (N_69,In_710,In_483);
and U70 (N_70,In_20,In_480);
nand U71 (N_71,In_333,In_735);
nor U72 (N_72,In_668,In_722);
or U73 (N_73,In_399,In_589);
and U74 (N_74,In_679,In_490);
nand U75 (N_75,In_570,In_37);
xor U76 (N_76,In_174,In_114);
nand U77 (N_77,In_257,In_467);
or U78 (N_78,In_727,In_384);
nand U79 (N_79,In_370,In_523);
nor U80 (N_80,In_682,In_349);
and U81 (N_81,In_593,In_137);
and U82 (N_82,In_566,In_624);
or U83 (N_83,In_457,In_598);
nor U84 (N_84,In_141,In_429);
nand U85 (N_85,In_536,In_607);
and U86 (N_86,In_136,In_43);
nor U87 (N_87,In_254,In_717);
or U88 (N_88,In_142,In_65);
and U89 (N_89,In_386,In_374);
nor U90 (N_90,In_635,In_183);
nand U91 (N_91,In_614,In_667);
or U92 (N_92,In_556,In_88);
nor U93 (N_93,In_637,In_494);
or U94 (N_94,In_638,In_172);
and U95 (N_95,In_502,In_407);
nor U96 (N_96,In_509,In_351);
or U97 (N_97,In_671,In_631);
and U98 (N_98,In_250,In_228);
nand U99 (N_99,In_459,In_372);
nor U100 (N_100,In_83,In_93);
nor U101 (N_101,In_466,In_197);
or U102 (N_102,In_654,In_70);
nand U103 (N_103,In_613,In_371);
or U104 (N_104,In_295,In_246);
nand U105 (N_105,In_108,In_498);
or U106 (N_106,In_403,In_474);
or U107 (N_107,In_119,In_218);
nor U108 (N_108,In_307,In_269);
nor U109 (N_109,In_718,In_546);
nand U110 (N_110,In_311,In_234);
nor U111 (N_111,In_647,In_328);
nor U112 (N_112,In_25,In_131);
or U113 (N_113,In_437,In_262);
and U114 (N_114,In_182,In_220);
and U115 (N_115,In_100,In_103);
or U116 (N_116,In_158,In_91);
nand U117 (N_117,In_742,In_313);
or U118 (N_118,In_626,In_198);
or U119 (N_119,In_104,In_499);
nand U120 (N_120,In_460,In_248);
or U121 (N_121,In_213,In_52);
and U122 (N_122,In_341,In_67);
or U123 (N_123,In_540,In_711);
nand U124 (N_124,In_714,In_206);
or U125 (N_125,In_741,In_389);
or U126 (N_126,In_40,In_256);
or U127 (N_127,In_648,In_98);
nor U128 (N_128,In_12,In_496);
and U129 (N_129,In_33,In_552);
and U130 (N_130,In_562,In_410);
nor U131 (N_131,In_23,In_415);
and U132 (N_132,In_379,In_601);
or U133 (N_133,In_270,In_708);
and U134 (N_134,In_507,In_322);
nor U135 (N_135,In_422,In_644);
nor U136 (N_136,In_186,In_425);
nor U137 (N_137,In_686,In_643);
nand U138 (N_138,In_189,In_655);
nor U139 (N_139,In_600,In_456);
and U140 (N_140,In_115,In_486);
or U141 (N_141,In_284,In_744);
nand U142 (N_142,In_304,In_612);
nand U143 (N_143,In_272,In_62);
nor U144 (N_144,In_34,In_723);
or U145 (N_145,In_702,In_699);
nand U146 (N_146,In_690,In_650);
or U147 (N_147,In_587,In_713);
or U148 (N_148,In_633,In_352);
and U149 (N_149,In_110,In_235);
nand U150 (N_150,In_531,In_325);
and U151 (N_151,In_120,In_550);
and U152 (N_152,In_619,In_39);
and U153 (N_153,In_303,In_133);
or U154 (N_154,In_528,In_0);
or U155 (N_155,In_448,In_376);
nand U156 (N_156,In_719,In_348);
and U157 (N_157,In_391,In_581);
nand U158 (N_158,In_675,In_167);
or U159 (N_159,In_255,In_253);
nand U160 (N_160,In_31,In_378);
and U161 (N_161,In_560,In_380);
or U162 (N_162,In_334,In_314);
nand U163 (N_163,In_36,In_530);
nor U164 (N_164,In_703,In_580);
nor U165 (N_165,In_748,In_72);
nor U166 (N_166,In_548,In_305);
nand U167 (N_167,In_8,In_173);
nor U168 (N_168,In_730,In_746);
nand U169 (N_169,In_640,In_588);
nor U170 (N_170,In_382,In_264);
nand U171 (N_171,In_430,In_594);
and U172 (N_172,In_396,In_97);
nand U173 (N_173,In_126,In_522);
and U174 (N_174,In_491,In_720);
and U175 (N_175,In_435,In_127);
or U176 (N_176,In_282,In_543);
and U177 (N_177,In_53,In_400);
nor U178 (N_178,In_73,In_111);
nor U179 (N_179,In_60,In_2);
and U180 (N_180,In_569,In_729);
nor U181 (N_181,In_165,In_477);
xnor U182 (N_182,In_319,In_574);
or U183 (N_183,In_176,In_324);
nor U184 (N_184,In_545,In_673);
or U185 (N_185,In_427,In_563);
nor U186 (N_186,In_628,In_222);
nand U187 (N_187,In_132,In_591);
or U188 (N_188,In_179,In_21);
xor U189 (N_189,In_244,In_464);
or U190 (N_190,In_424,In_672);
xnor U191 (N_191,In_6,In_99);
xnor U192 (N_192,In_211,In_301);
xor U193 (N_193,In_237,In_292);
or U194 (N_194,In_520,In_745);
nor U195 (N_195,In_463,In_185);
and U196 (N_196,In_290,In_177);
nand U197 (N_197,In_68,In_390);
and U198 (N_198,In_572,In_715);
and U199 (N_199,In_685,In_168);
nor U200 (N_200,In_280,In_245);
xnor U201 (N_201,In_318,In_696);
or U202 (N_202,In_321,In_109);
nand U203 (N_203,In_153,In_217);
nor U204 (N_204,In_433,In_238);
nand U205 (N_205,In_95,In_293);
nand U206 (N_206,In_105,In_661);
nor U207 (N_207,In_734,In_17);
and U208 (N_208,In_455,In_350);
or U209 (N_209,In_652,In_28);
and U210 (N_210,In_346,In_181);
nor U211 (N_211,In_582,In_428);
nand U212 (N_212,In_192,In_279);
or U213 (N_213,In_564,In_320);
or U214 (N_214,In_461,In_395);
and U215 (N_215,In_162,In_653);
nor U216 (N_216,In_694,In_533);
nand U217 (N_217,In_221,In_166);
or U218 (N_218,In_701,In_216);
or U219 (N_219,In_78,In_29);
nand U220 (N_220,In_583,In_362);
nor U221 (N_221,In_81,In_465);
and U222 (N_222,In_450,In_125);
or U223 (N_223,In_278,In_479);
or U224 (N_224,In_302,In_9);
xnor U225 (N_225,In_214,In_662);
nor U226 (N_226,In_327,In_342);
nand U227 (N_227,In_495,In_207);
nor U228 (N_228,In_116,In_657);
and U229 (N_229,In_50,In_170);
or U230 (N_230,In_71,In_205);
nand U231 (N_231,In_684,In_242);
nor U232 (N_232,In_549,In_482);
or U233 (N_233,In_687,In_408);
or U234 (N_234,In_56,In_547);
nand U235 (N_235,In_377,In_478);
nand U236 (N_236,In_294,In_49);
or U237 (N_237,In_551,In_381);
nor U238 (N_238,In_335,In_610);
and U239 (N_239,In_515,In_112);
nand U240 (N_240,In_194,In_660);
nand U241 (N_241,In_336,In_510);
and U242 (N_242,In_611,In_524);
nand U243 (N_243,In_473,In_512);
nand U244 (N_244,In_329,In_501);
nand U245 (N_245,In_621,In_169);
nand U246 (N_246,In_312,In_595);
nor U247 (N_247,In_645,In_414);
and U248 (N_248,In_338,In_209);
and U249 (N_249,In_260,In_559);
and U250 (N_250,In_525,In_716);
or U251 (N_251,In_196,In_231);
or U252 (N_252,In_526,In_202);
nor U253 (N_253,In_663,In_261);
and U254 (N_254,In_360,In_130);
and U255 (N_255,In_676,In_700);
nand U256 (N_256,In_511,In_431);
and U257 (N_257,In_233,In_739);
and U258 (N_258,In_4,In_606);
and U259 (N_259,In_411,In_447);
nor U260 (N_260,In_698,In_267);
and U261 (N_261,In_646,In_608);
nand U262 (N_262,In_692,In_409);
nor U263 (N_263,In_101,In_308);
or U264 (N_264,In_159,In_161);
and U265 (N_265,In_241,In_59);
xnor U266 (N_266,In_368,In_434);
or U267 (N_267,In_578,In_344);
nor U268 (N_268,In_44,In_623);
and U269 (N_269,In_87,In_420);
or U270 (N_270,In_135,In_387);
nand U271 (N_271,In_243,In_193);
nor U272 (N_272,In_69,In_289);
nor U273 (N_273,In_286,In_359);
nand U274 (N_274,In_597,In_5);
and U275 (N_275,In_140,In_191);
xnor U276 (N_276,In_732,In_627);
or U277 (N_277,In_634,In_160);
or U278 (N_278,In_227,In_677);
nor U279 (N_279,In_725,In_605);
nand U280 (N_280,In_355,In_541);
nand U281 (N_281,In_443,In_77);
or U282 (N_282,In_451,In_740);
nor U283 (N_283,In_47,In_225);
or U284 (N_284,In_353,In_239);
nand U285 (N_285,In_412,In_630);
xnor U286 (N_286,In_413,In_356);
or U287 (N_287,In_534,In_274);
or U288 (N_288,In_731,In_470);
or U289 (N_289,In_401,In_666);
nand U290 (N_290,In_148,In_508);
and U291 (N_291,In_45,In_224);
or U292 (N_292,In_339,In_180);
and U293 (N_293,In_497,In_561);
or U294 (N_294,In_51,In_10);
nand U295 (N_295,In_603,In_361);
and U296 (N_296,In_418,In_513);
and U297 (N_297,In_46,In_405);
or U298 (N_298,In_481,In_398);
nor U299 (N_299,In_345,In_92);
nand U300 (N_300,In_590,In_452);
or U301 (N_301,In_204,In_123);
or U302 (N_302,In_680,In_500);
nor U303 (N_303,In_55,In_688);
or U304 (N_304,In_210,In_199);
nor U305 (N_305,In_32,In_200);
and U306 (N_306,In_592,In_453);
nand U307 (N_307,In_15,In_76);
nand U308 (N_308,In_505,In_404);
nand U309 (N_309,In_58,In_297);
or U310 (N_310,In_223,In_288);
or U311 (N_311,In_579,In_149);
and U312 (N_312,In_620,In_300);
nor U313 (N_313,In_539,In_629);
or U314 (N_314,In_38,In_402);
nand U315 (N_315,In_472,In_584);
and U316 (N_316,In_416,In_275);
and U317 (N_317,In_57,In_11);
nand U318 (N_318,In_277,In_249);
or U319 (N_319,In_419,In_476);
nand U320 (N_320,In_575,In_117);
and U321 (N_321,In_310,In_678);
and U322 (N_322,In_61,In_79);
and U323 (N_323,In_388,In_707);
and U324 (N_324,In_129,In_417);
or U325 (N_325,In_519,In_695);
nand U326 (N_326,In_247,In_323);
and U327 (N_327,In_577,In_622);
and U328 (N_328,In_232,In_367);
nand U329 (N_329,In_485,In_567);
or U330 (N_330,In_469,In_693);
and U331 (N_331,In_48,In_538);
and U332 (N_332,In_30,In_712);
and U333 (N_333,In_1,In_363);
nand U334 (N_334,In_423,In_26);
or U335 (N_335,In_527,In_85);
or U336 (N_336,In_190,In_330);
and U337 (N_337,In_383,In_35);
or U338 (N_338,In_281,In_442);
nor U339 (N_339,In_316,In_178);
nand U340 (N_340,In_139,In_128);
nor U341 (N_341,In_529,In_521);
nand U342 (N_342,In_22,In_554);
and U343 (N_343,In_736,In_84);
nand U344 (N_344,In_195,In_444);
nand U345 (N_345,In_445,In_155);
and U346 (N_346,In_138,In_89);
and U347 (N_347,In_122,In_642);
nand U348 (N_348,In_728,In_475);
xnor U349 (N_349,In_276,In_96);
and U350 (N_350,In_743,In_441);
nand U351 (N_351,In_19,In_557);
nand U352 (N_352,In_397,In_63);
nand U353 (N_353,In_489,In_747);
nor U354 (N_354,In_669,In_369);
and U355 (N_355,In_665,In_285);
and U356 (N_356,In_724,In_446);
and U357 (N_357,In_365,In_306);
nand U358 (N_358,In_373,In_66);
or U359 (N_359,In_487,In_616);
or U360 (N_360,In_705,In_537);
nand U361 (N_361,In_106,In_263);
nand U362 (N_362,In_236,In_157);
and U363 (N_363,In_440,In_147);
and U364 (N_364,In_171,In_364);
or U365 (N_365,In_121,In_134);
and U366 (N_366,In_107,In_553);
xnor U367 (N_367,In_602,In_506);
nand U368 (N_368,In_298,In_674);
or U369 (N_369,In_13,In_438);
and U370 (N_370,In_488,In_219);
or U371 (N_371,In_558,In_749);
and U372 (N_372,In_201,In_41);
nand U373 (N_373,In_24,In_331);
nand U374 (N_374,In_187,In_617);
xor U375 (N_375,In_23,In_9);
nand U376 (N_376,In_715,In_484);
nand U377 (N_377,In_672,In_241);
nor U378 (N_378,In_726,In_50);
and U379 (N_379,In_120,In_400);
and U380 (N_380,In_445,In_711);
nand U381 (N_381,In_749,In_452);
xnor U382 (N_382,In_652,In_373);
nor U383 (N_383,In_390,In_410);
or U384 (N_384,In_228,In_705);
xnor U385 (N_385,In_532,In_410);
xnor U386 (N_386,In_142,In_109);
and U387 (N_387,In_59,In_528);
or U388 (N_388,In_478,In_187);
and U389 (N_389,In_326,In_710);
nand U390 (N_390,In_417,In_629);
nand U391 (N_391,In_413,In_653);
nand U392 (N_392,In_207,In_312);
or U393 (N_393,In_5,In_267);
nor U394 (N_394,In_315,In_702);
xnor U395 (N_395,In_404,In_225);
nor U396 (N_396,In_500,In_228);
nand U397 (N_397,In_732,In_590);
nand U398 (N_398,In_171,In_156);
or U399 (N_399,In_227,In_345);
nand U400 (N_400,In_232,In_652);
or U401 (N_401,In_417,In_41);
and U402 (N_402,In_731,In_269);
nor U403 (N_403,In_710,In_701);
nand U404 (N_404,In_259,In_722);
nand U405 (N_405,In_515,In_43);
and U406 (N_406,In_511,In_365);
nor U407 (N_407,In_196,In_526);
nand U408 (N_408,In_641,In_269);
and U409 (N_409,In_644,In_559);
and U410 (N_410,In_345,In_535);
or U411 (N_411,In_144,In_93);
or U412 (N_412,In_531,In_510);
and U413 (N_413,In_672,In_645);
or U414 (N_414,In_594,In_625);
and U415 (N_415,In_206,In_189);
or U416 (N_416,In_685,In_551);
nor U417 (N_417,In_26,In_311);
nor U418 (N_418,In_273,In_597);
nand U419 (N_419,In_735,In_315);
or U420 (N_420,In_265,In_452);
nand U421 (N_421,In_351,In_723);
nor U422 (N_422,In_343,In_356);
or U423 (N_423,In_566,In_308);
and U424 (N_424,In_487,In_155);
nand U425 (N_425,In_548,In_673);
nand U426 (N_426,In_285,In_130);
or U427 (N_427,In_551,In_524);
or U428 (N_428,In_102,In_397);
xnor U429 (N_429,In_583,In_267);
nor U430 (N_430,In_5,In_510);
nand U431 (N_431,In_332,In_538);
and U432 (N_432,In_446,In_159);
nor U433 (N_433,In_736,In_698);
nand U434 (N_434,In_256,In_642);
nor U435 (N_435,In_150,In_83);
nor U436 (N_436,In_463,In_18);
and U437 (N_437,In_68,In_409);
or U438 (N_438,In_528,In_731);
xnor U439 (N_439,In_392,In_375);
or U440 (N_440,In_370,In_687);
or U441 (N_441,In_439,In_255);
nor U442 (N_442,In_670,In_599);
and U443 (N_443,In_698,In_79);
and U444 (N_444,In_699,In_236);
and U445 (N_445,In_637,In_475);
or U446 (N_446,In_525,In_116);
nand U447 (N_447,In_251,In_717);
or U448 (N_448,In_702,In_583);
nand U449 (N_449,In_596,In_520);
nor U450 (N_450,In_738,In_94);
nor U451 (N_451,In_142,In_518);
nand U452 (N_452,In_148,In_175);
nor U453 (N_453,In_725,In_430);
or U454 (N_454,In_383,In_422);
and U455 (N_455,In_290,In_312);
and U456 (N_456,In_228,In_669);
nor U457 (N_457,In_410,In_567);
nor U458 (N_458,In_334,In_180);
and U459 (N_459,In_317,In_182);
nand U460 (N_460,In_114,In_99);
or U461 (N_461,In_117,In_680);
nor U462 (N_462,In_246,In_3);
nor U463 (N_463,In_568,In_491);
or U464 (N_464,In_207,In_624);
xnor U465 (N_465,In_374,In_501);
nand U466 (N_466,In_257,In_648);
or U467 (N_467,In_572,In_137);
nor U468 (N_468,In_556,In_732);
or U469 (N_469,In_213,In_462);
nor U470 (N_470,In_164,In_433);
nor U471 (N_471,In_114,In_451);
nor U472 (N_472,In_274,In_189);
nor U473 (N_473,In_172,In_216);
nand U474 (N_474,In_444,In_636);
and U475 (N_475,In_63,In_511);
nor U476 (N_476,In_189,In_628);
nand U477 (N_477,In_293,In_44);
nor U478 (N_478,In_27,In_126);
nand U479 (N_479,In_635,In_289);
or U480 (N_480,In_113,In_366);
nand U481 (N_481,In_349,In_122);
nor U482 (N_482,In_231,In_368);
nand U483 (N_483,In_45,In_85);
nor U484 (N_484,In_10,In_533);
xor U485 (N_485,In_299,In_74);
xnor U486 (N_486,In_393,In_567);
and U487 (N_487,In_236,In_600);
or U488 (N_488,In_182,In_88);
nand U489 (N_489,In_434,In_580);
nor U490 (N_490,In_617,In_286);
and U491 (N_491,In_584,In_173);
nand U492 (N_492,In_50,In_694);
nor U493 (N_493,In_406,In_167);
nor U494 (N_494,In_735,In_188);
nand U495 (N_495,In_159,In_413);
nor U496 (N_496,In_65,In_709);
and U497 (N_497,In_643,In_719);
or U498 (N_498,In_102,In_436);
nand U499 (N_499,In_508,In_277);
and U500 (N_500,N_60,N_221);
nor U501 (N_501,N_205,N_431);
nand U502 (N_502,N_196,N_136);
or U503 (N_503,N_24,N_63);
and U504 (N_504,N_39,N_386);
nand U505 (N_505,N_295,N_401);
and U506 (N_506,N_365,N_255);
nor U507 (N_507,N_347,N_204);
and U508 (N_508,N_174,N_184);
or U509 (N_509,N_469,N_310);
or U510 (N_510,N_300,N_170);
and U511 (N_511,N_16,N_473);
and U512 (N_512,N_46,N_351);
nand U513 (N_513,N_165,N_207);
nand U514 (N_514,N_292,N_408);
and U515 (N_515,N_82,N_225);
and U516 (N_516,N_102,N_139);
nand U517 (N_517,N_360,N_297);
nor U518 (N_518,N_135,N_324);
and U519 (N_519,N_433,N_305);
or U520 (N_520,N_419,N_450);
and U521 (N_521,N_229,N_114);
nand U522 (N_522,N_220,N_329);
and U523 (N_523,N_238,N_141);
nand U524 (N_524,N_234,N_390);
and U525 (N_525,N_402,N_302);
nor U526 (N_526,N_12,N_296);
and U527 (N_527,N_458,N_421);
nand U528 (N_528,N_110,N_298);
and U529 (N_529,N_389,N_308);
nor U530 (N_530,N_363,N_479);
and U531 (N_531,N_407,N_263);
nand U532 (N_532,N_166,N_59);
nand U533 (N_533,N_427,N_45);
nor U534 (N_534,N_1,N_465);
and U535 (N_535,N_118,N_32);
nor U536 (N_536,N_357,N_333);
nand U537 (N_537,N_299,N_482);
nor U538 (N_538,N_154,N_335);
nand U539 (N_539,N_151,N_105);
or U540 (N_540,N_303,N_278);
or U541 (N_541,N_9,N_442);
nand U542 (N_542,N_31,N_285);
nand U543 (N_543,N_98,N_89);
and U544 (N_544,N_287,N_273);
nand U545 (N_545,N_80,N_288);
nand U546 (N_546,N_157,N_35);
xor U547 (N_547,N_282,N_168);
xor U548 (N_548,N_11,N_8);
nor U549 (N_549,N_199,N_200);
or U550 (N_550,N_256,N_131);
nor U551 (N_551,N_384,N_396);
nand U552 (N_552,N_393,N_489);
nor U553 (N_553,N_249,N_474);
or U554 (N_554,N_178,N_435);
and U555 (N_555,N_180,N_499);
nand U556 (N_556,N_337,N_439);
and U557 (N_557,N_19,N_491);
nor U558 (N_558,N_179,N_159);
nand U559 (N_559,N_284,N_3);
or U560 (N_560,N_22,N_124);
or U561 (N_561,N_270,N_72);
nor U562 (N_562,N_466,N_93);
xnor U563 (N_563,N_190,N_133);
nor U564 (N_564,N_475,N_422);
nand U565 (N_565,N_283,N_91);
or U566 (N_566,N_368,N_173);
and U567 (N_567,N_428,N_318);
nor U568 (N_568,N_275,N_158);
or U569 (N_569,N_84,N_240);
nand U570 (N_570,N_29,N_241);
and U571 (N_571,N_254,N_252);
or U572 (N_572,N_239,N_334);
nand U573 (N_573,N_486,N_494);
nor U574 (N_574,N_65,N_88);
nand U575 (N_575,N_2,N_152);
nor U576 (N_576,N_478,N_20);
nand U577 (N_577,N_456,N_370);
nor U578 (N_578,N_484,N_113);
or U579 (N_579,N_194,N_79);
or U580 (N_580,N_392,N_28);
nor U581 (N_581,N_201,N_211);
and U582 (N_582,N_155,N_423);
and U583 (N_583,N_50,N_230);
and U584 (N_584,N_411,N_359);
nand U585 (N_585,N_18,N_78);
and U586 (N_586,N_100,N_235);
nor U587 (N_587,N_62,N_150);
and U588 (N_588,N_214,N_380);
nor U589 (N_589,N_14,N_243);
nor U590 (N_590,N_438,N_76);
or U591 (N_591,N_485,N_497);
or U592 (N_592,N_344,N_189);
nor U593 (N_593,N_463,N_391);
nand U594 (N_594,N_148,N_25);
and U595 (N_595,N_128,N_232);
and U596 (N_596,N_259,N_352);
and U597 (N_597,N_58,N_228);
or U598 (N_598,N_341,N_245);
nor U599 (N_599,N_195,N_217);
and U600 (N_600,N_52,N_33);
nor U601 (N_601,N_187,N_26);
or U602 (N_602,N_403,N_247);
nand U603 (N_603,N_446,N_440);
nand U604 (N_604,N_317,N_361);
nor U605 (N_605,N_425,N_413);
or U606 (N_606,N_362,N_77);
nor U607 (N_607,N_345,N_452);
nor U608 (N_608,N_67,N_304);
nand U609 (N_609,N_371,N_289);
nor U610 (N_610,N_294,N_0);
and U611 (N_611,N_429,N_400);
and U612 (N_612,N_115,N_129);
and U613 (N_613,N_472,N_13);
or U614 (N_614,N_40,N_346);
nand U615 (N_615,N_350,N_197);
and U616 (N_616,N_117,N_41);
nor U617 (N_617,N_258,N_264);
and U618 (N_618,N_379,N_426);
nand U619 (N_619,N_164,N_260);
nand U620 (N_620,N_281,N_87);
nor U621 (N_621,N_343,N_175);
and U622 (N_622,N_138,N_274);
or U623 (N_623,N_309,N_147);
and U624 (N_624,N_97,N_387);
or U625 (N_625,N_444,N_301);
nand U626 (N_626,N_276,N_216);
or U627 (N_627,N_161,N_315);
or U628 (N_628,N_325,N_464);
nand U629 (N_629,N_470,N_74);
or U630 (N_630,N_353,N_55);
and U631 (N_631,N_376,N_443);
and U632 (N_632,N_412,N_64);
nor U633 (N_633,N_85,N_107);
nor U634 (N_634,N_468,N_261);
nand U635 (N_635,N_23,N_244);
and U636 (N_636,N_354,N_434);
or U637 (N_637,N_323,N_42);
nand U638 (N_638,N_126,N_206);
nand U639 (N_639,N_231,N_405);
nor U640 (N_640,N_348,N_457);
nor U641 (N_641,N_373,N_218);
or U642 (N_642,N_48,N_108);
nor U643 (N_643,N_417,N_43);
and U644 (N_644,N_415,N_449);
nand U645 (N_645,N_103,N_210);
nand U646 (N_646,N_153,N_459);
or U647 (N_647,N_382,N_383);
nor U648 (N_648,N_34,N_242);
or U649 (N_649,N_92,N_492);
or U650 (N_650,N_219,N_330);
nor U651 (N_651,N_375,N_462);
nor U652 (N_652,N_251,N_293);
nand U653 (N_653,N_266,N_83);
and U654 (N_654,N_71,N_101);
nand U655 (N_655,N_253,N_476);
nand U656 (N_656,N_398,N_163);
and U657 (N_657,N_146,N_208);
or U658 (N_658,N_54,N_445);
or U659 (N_659,N_185,N_377);
and U660 (N_660,N_339,N_306);
or U661 (N_661,N_191,N_81);
or U662 (N_662,N_495,N_156);
nor U663 (N_663,N_268,N_224);
and U664 (N_664,N_467,N_149);
or U665 (N_665,N_112,N_49);
nand U666 (N_666,N_336,N_192);
xor U667 (N_667,N_409,N_183);
nand U668 (N_668,N_436,N_483);
or U669 (N_669,N_397,N_202);
or U670 (N_670,N_420,N_327);
and U671 (N_671,N_496,N_73);
nand U672 (N_672,N_291,N_132);
and U673 (N_673,N_6,N_314);
and U674 (N_674,N_290,N_320);
nor U675 (N_675,N_21,N_56);
nand U676 (N_676,N_342,N_328);
nor U677 (N_677,N_262,N_250);
nor U678 (N_678,N_367,N_271);
nor U679 (N_679,N_86,N_374);
or U680 (N_680,N_280,N_441);
nand U681 (N_681,N_277,N_319);
nand U682 (N_682,N_246,N_142);
or U683 (N_683,N_188,N_57);
nor U684 (N_684,N_487,N_104);
and U685 (N_685,N_404,N_223);
nor U686 (N_686,N_167,N_455);
or U687 (N_687,N_203,N_477);
xor U688 (N_688,N_460,N_182);
or U689 (N_689,N_171,N_414);
and U690 (N_690,N_169,N_447);
nand U691 (N_691,N_237,N_316);
or U692 (N_692,N_338,N_36);
or U693 (N_693,N_257,N_61);
nor U694 (N_694,N_222,N_448);
and U695 (N_695,N_68,N_358);
nand U696 (N_696,N_481,N_140);
or U697 (N_697,N_137,N_215);
nor U698 (N_698,N_134,N_498);
or U699 (N_699,N_322,N_176);
nand U700 (N_700,N_332,N_286);
or U701 (N_701,N_10,N_488);
and U702 (N_702,N_99,N_5);
or U703 (N_703,N_395,N_130);
and U704 (N_704,N_17,N_27);
and U705 (N_705,N_418,N_490);
nand U706 (N_706,N_127,N_480);
nor U707 (N_707,N_172,N_53);
nor U708 (N_708,N_461,N_209);
or U709 (N_709,N_95,N_66);
or U710 (N_710,N_378,N_437);
and U711 (N_711,N_96,N_4);
nand U712 (N_712,N_424,N_15);
nor U713 (N_713,N_7,N_122);
and U714 (N_714,N_111,N_51);
or U715 (N_715,N_227,N_356);
or U716 (N_716,N_410,N_44);
nand U717 (N_717,N_70,N_331);
and U718 (N_718,N_366,N_453);
and U719 (N_719,N_451,N_116);
xor U720 (N_720,N_121,N_181);
or U721 (N_721,N_406,N_269);
and U722 (N_722,N_388,N_381);
and U723 (N_723,N_144,N_38);
nor U724 (N_724,N_119,N_236);
and U725 (N_725,N_369,N_265);
nand U726 (N_726,N_372,N_313);
nor U727 (N_727,N_94,N_471);
nor U728 (N_728,N_340,N_364);
nor U729 (N_729,N_106,N_233);
or U730 (N_730,N_267,N_430);
nand U731 (N_731,N_37,N_394);
nand U732 (N_732,N_432,N_90);
or U733 (N_733,N_125,N_109);
or U734 (N_734,N_75,N_162);
nand U735 (N_735,N_272,N_454);
or U736 (N_736,N_143,N_307);
or U737 (N_737,N_30,N_212);
nand U738 (N_738,N_349,N_385);
and U739 (N_739,N_69,N_145);
nand U740 (N_740,N_326,N_47);
nor U741 (N_741,N_355,N_120);
nand U742 (N_742,N_248,N_493);
or U743 (N_743,N_160,N_226);
nand U744 (N_744,N_177,N_311);
or U745 (N_745,N_123,N_279);
or U746 (N_746,N_399,N_321);
nor U747 (N_747,N_416,N_198);
or U748 (N_748,N_312,N_186);
or U749 (N_749,N_193,N_213);
or U750 (N_750,N_226,N_147);
nand U751 (N_751,N_28,N_444);
nor U752 (N_752,N_495,N_59);
or U753 (N_753,N_387,N_462);
nor U754 (N_754,N_98,N_35);
and U755 (N_755,N_77,N_404);
and U756 (N_756,N_154,N_93);
nor U757 (N_757,N_475,N_433);
and U758 (N_758,N_295,N_147);
and U759 (N_759,N_351,N_283);
nand U760 (N_760,N_438,N_283);
or U761 (N_761,N_249,N_413);
or U762 (N_762,N_117,N_61);
and U763 (N_763,N_390,N_83);
or U764 (N_764,N_324,N_112);
and U765 (N_765,N_467,N_177);
nand U766 (N_766,N_419,N_441);
nor U767 (N_767,N_13,N_439);
and U768 (N_768,N_195,N_280);
nand U769 (N_769,N_163,N_240);
or U770 (N_770,N_255,N_89);
and U771 (N_771,N_186,N_482);
and U772 (N_772,N_416,N_352);
nor U773 (N_773,N_369,N_308);
and U774 (N_774,N_165,N_33);
nor U775 (N_775,N_322,N_109);
nand U776 (N_776,N_308,N_138);
nand U777 (N_777,N_221,N_192);
or U778 (N_778,N_306,N_424);
or U779 (N_779,N_258,N_18);
or U780 (N_780,N_215,N_280);
and U781 (N_781,N_192,N_262);
nand U782 (N_782,N_411,N_188);
nor U783 (N_783,N_469,N_260);
or U784 (N_784,N_66,N_57);
nor U785 (N_785,N_254,N_303);
nor U786 (N_786,N_315,N_278);
nor U787 (N_787,N_474,N_419);
and U788 (N_788,N_342,N_372);
and U789 (N_789,N_407,N_318);
nand U790 (N_790,N_57,N_484);
or U791 (N_791,N_203,N_250);
nor U792 (N_792,N_448,N_380);
nand U793 (N_793,N_15,N_247);
nand U794 (N_794,N_15,N_13);
or U795 (N_795,N_279,N_443);
and U796 (N_796,N_231,N_494);
or U797 (N_797,N_451,N_296);
and U798 (N_798,N_293,N_19);
or U799 (N_799,N_61,N_249);
or U800 (N_800,N_320,N_378);
and U801 (N_801,N_463,N_394);
nor U802 (N_802,N_353,N_424);
and U803 (N_803,N_30,N_304);
and U804 (N_804,N_287,N_143);
and U805 (N_805,N_73,N_483);
and U806 (N_806,N_80,N_119);
nand U807 (N_807,N_481,N_48);
and U808 (N_808,N_138,N_253);
or U809 (N_809,N_92,N_9);
nand U810 (N_810,N_492,N_273);
xnor U811 (N_811,N_116,N_417);
nor U812 (N_812,N_270,N_124);
and U813 (N_813,N_409,N_389);
nor U814 (N_814,N_290,N_330);
nand U815 (N_815,N_59,N_387);
and U816 (N_816,N_395,N_286);
or U817 (N_817,N_63,N_376);
and U818 (N_818,N_77,N_136);
nand U819 (N_819,N_227,N_220);
or U820 (N_820,N_236,N_106);
nand U821 (N_821,N_161,N_426);
or U822 (N_822,N_159,N_211);
or U823 (N_823,N_173,N_91);
and U824 (N_824,N_339,N_499);
and U825 (N_825,N_294,N_265);
and U826 (N_826,N_341,N_453);
nand U827 (N_827,N_249,N_43);
nor U828 (N_828,N_127,N_108);
or U829 (N_829,N_191,N_186);
nor U830 (N_830,N_40,N_118);
nand U831 (N_831,N_484,N_450);
and U832 (N_832,N_139,N_299);
or U833 (N_833,N_355,N_252);
nor U834 (N_834,N_361,N_475);
and U835 (N_835,N_269,N_247);
nor U836 (N_836,N_342,N_387);
nand U837 (N_837,N_41,N_9);
and U838 (N_838,N_489,N_243);
or U839 (N_839,N_33,N_282);
or U840 (N_840,N_407,N_119);
nand U841 (N_841,N_448,N_348);
nand U842 (N_842,N_388,N_375);
nand U843 (N_843,N_92,N_374);
xnor U844 (N_844,N_340,N_206);
nand U845 (N_845,N_113,N_446);
or U846 (N_846,N_94,N_224);
xnor U847 (N_847,N_355,N_229);
nand U848 (N_848,N_21,N_22);
or U849 (N_849,N_405,N_336);
nor U850 (N_850,N_207,N_483);
xnor U851 (N_851,N_473,N_237);
or U852 (N_852,N_325,N_221);
nand U853 (N_853,N_152,N_139);
and U854 (N_854,N_240,N_484);
xnor U855 (N_855,N_102,N_353);
and U856 (N_856,N_253,N_356);
nand U857 (N_857,N_134,N_193);
nor U858 (N_858,N_25,N_362);
nand U859 (N_859,N_455,N_209);
or U860 (N_860,N_199,N_394);
and U861 (N_861,N_343,N_378);
and U862 (N_862,N_445,N_290);
nor U863 (N_863,N_458,N_213);
and U864 (N_864,N_474,N_126);
nand U865 (N_865,N_467,N_132);
and U866 (N_866,N_427,N_244);
nor U867 (N_867,N_220,N_393);
xor U868 (N_868,N_379,N_364);
and U869 (N_869,N_31,N_244);
nand U870 (N_870,N_314,N_422);
nor U871 (N_871,N_289,N_22);
nor U872 (N_872,N_277,N_38);
and U873 (N_873,N_348,N_272);
nand U874 (N_874,N_225,N_296);
xnor U875 (N_875,N_493,N_318);
nor U876 (N_876,N_245,N_108);
and U877 (N_877,N_335,N_75);
nand U878 (N_878,N_181,N_393);
nand U879 (N_879,N_181,N_8);
xor U880 (N_880,N_115,N_59);
nand U881 (N_881,N_301,N_499);
nor U882 (N_882,N_194,N_126);
or U883 (N_883,N_354,N_23);
or U884 (N_884,N_148,N_284);
and U885 (N_885,N_431,N_261);
nand U886 (N_886,N_173,N_385);
or U887 (N_887,N_37,N_213);
and U888 (N_888,N_211,N_307);
or U889 (N_889,N_96,N_74);
or U890 (N_890,N_432,N_324);
nand U891 (N_891,N_334,N_274);
nor U892 (N_892,N_154,N_393);
or U893 (N_893,N_119,N_391);
nand U894 (N_894,N_443,N_119);
nand U895 (N_895,N_109,N_237);
or U896 (N_896,N_181,N_107);
or U897 (N_897,N_485,N_399);
nand U898 (N_898,N_233,N_171);
or U899 (N_899,N_128,N_237);
nand U900 (N_900,N_33,N_188);
nand U901 (N_901,N_461,N_412);
nor U902 (N_902,N_289,N_50);
nand U903 (N_903,N_465,N_325);
xnor U904 (N_904,N_327,N_32);
nor U905 (N_905,N_343,N_25);
or U906 (N_906,N_207,N_142);
and U907 (N_907,N_119,N_113);
nor U908 (N_908,N_3,N_18);
and U909 (N_909,N_411,N_221);
nand U910 (N_910,N_367,N_134);
nand U911 (N_911,N_179,N_430);
nand U912 (N_912,N_435,N_360);
nor U913 (N_913,N_451,N_381);
or U914 (N_914,N_379,N_279);
nand U915 (N_915,N_269,N_81);
nor U916 (N_916,N_80,N_266);
or U917 (N_917,N_253,N_193);
or U918 (N_918,N_234,N_178);
nor U919 (N_919,N_326,N_356);
or U920 (N_920,N_277,N_172);
nand U921 (N_921,N_478,N_67);
or U922 (N_922,N_99,N_233);
nor U923 (N_923,N_283,N_291);
and U924 (N_924,N_241,N_384);
xor U925 (N_925,N_182,N_210);
or U926 (N_926,N_104,N_465);
xnor U927 (N_927,N_106,N_435);
nor U928 (N_928,N_300,N_133);
nand U929 (N_929,N_460,N_498);
nand U930 (N_930,N_469,N_214);
nand U931 (N_931,N_362,N_255);
or U932 (N_932,N_51,N_474);
nand U933 (N_933,N_140,N_447);
nand U934 (N_934,N_216,N_297);
or U935 (N_935,N_351,N_284);
and U936 (N_936,N_433,N_170);
or U937 (N_937,N_468,N_36);
and U938 (N_938,N_459,N_280);
and U939 (N_939,N_58,N_265);
nand U940 (N_940,N_65,N_212);
nor U941 (N_941,N_298,N_361);
or U942 (N_942,N_23,N_201);
nand U943 (N_943,N_273,N_333);
nor U944 (N_944,N_339,N_105);
nand U945 (N_945,N_364,N_497);
nor U946 (N_946,N_80,N_323);
nand U947 (N_947,N_370,N_492);
and U948 (N_948,N_331,N_246);
and U949 (N_949,N_466,N_259);
or U950 (N_950,N_65,N_184);
nand U951 (N_951,N_122,N_493);
nand U952 (N_952,N_472,N_18);
and U953 (N_953,N_410,N_381);
and U954 (N_954,N_174,N_250);
and U955 (N_955,N_466,N_155);
nand U956 (N_956,N_124,N_149);
nand U957 (N_957,N_452,N_113);
or U958 (N_958,N_253,N_53);
nand U959 (N_959,N_133,N_198);
and U960 (N_960,N_422,N_249);
nand U961 (N_961,N_406,N_199);
and U962 (N_962,N_271,N_1);
or U963 (N_963,N_54,N_386);
or U964 (N_964,N_458,N_286);
nor U965 (N_965,N_151,N_33);
and U966 (N_966,N_318,N_197);
nor U967 (N_967,N_392,N_236);
nand U968 (N_968,N_40,N_406);
and U969 (N_969,N_263,N_82);
nand U970 (N_970,N_88,N_19);
or U971 (N_971,N_360,N_32);
or U972 (N_972,N_307,N_355);
nand U973 (N_973,N_399,N_464);
and U974 (N_974,N_62,N_213);
nor U975 (N_975,N_55,N_199);
nand U976 (N_976,N_227,N_116);
nor U977 (N_977,N_243,N_24);
or U978 (N_978,N_413,N_12);
and U979 (N_979,N_182,N_171);
nand U980 (N_980,N_230,N_52);
and U981 (N_981,N_169,N_295);
and U982 (N_982,N_273,N_348);
xnor U983 (N_983,N_401,N_332);
or U984 (N_984,N_435,N_344);
nor U985 (N_985,N_198,N_127);
or U986 (N_986,N_39,N_343);
nor U987 (N_987,N_426,N_194);
and U988 (N_988,N_267,N_244);
nand U989 (N_989,N_47,N_176);
and U990 (N_990,N_179,N_62);
nor U991 (N_991,N_431,N_485);
nand U992 (N_992,N_446,N_296);
and U993 (N_993,N_394,N_438);
or U994 (N_994,N_165,N_297);
nor U995 (N_995,N_330,N_363);
nor U996 (N_996,N_354,N_42);
or U997 (N_997,N_451,N_234);
nand U998 (N_998,N_270,N_46);
or U999 (N_999,N_462,N_267);
or U1000 (N_1000,N_694,N_782);
nor U1001 (N_1001,N_703,N_581);
and U1002 (N_1002,N_851,N_614);
nand U1003 (N_1003,N_714,N_546);
nor U1004 (N_1004,N_684,N_661);
or U1005 (N_1005,N_855,N_665);
nand U1006 (N_1006,N_504,N_867);
and U1007 (N_1007,N_557,N_635);
or U1008 (N_1008,N_746,N_956);
nand U1009 (N_1009,N_599,N_869);
nor U1010 (N_1010,N_908,N_821);
and U1011 (N_1011,N_965,N_912);
nor U1012 (N_1012,N_553,N_626);
nor U1013 (N_1013,N_894,N_536);
nor U1014 (N_1014,N_976,N_803);
and U1015 (N_1015,N_566,N_818);
nor U1016 (N_1016,N_530,N_570);
or U1017 (N_1017,N_957,N_528);
nor U1018 (N_1018,N_556,N_751);
and U1019 (N_1019,N_892,N_507);
or U1020 (N_1020,N_659,N_651);
nand U1021 (N_1021,N_757,N_545);
and U1022 (N_1022,N_799,N_940);
or U1023 (N_1023,N_549,N_909);
or U1024 (N_1024,N_878,N_750);
nor U1025 (N_1025,N_730,N_834);
and U1026 (N_1026,N_502,N_796);
and U1027 (N_1027,N_766,N_920);
and U1028 (N_1028,N_575,N_736);
and U1029 (N_1029,N_781,N_786);
and U1030 (N_1030,N_603,N_945);
nand U1031 (N_1031,N_563,N_721);
nor U1032 (N_1032,N_817,N_939);
or U1033 (N_1033,N_697,N_875);
or U1034 (N_1034,N_512,N_764);
or U1035 (N_1035,N_726,N_707);
or U1036 (N_1036,N_578,N_858);
nor U1037 (N_1037,N_637,N_889);
nor U1038 (N_1038,N_706,N_871);
or U1039 (N_1039,N_668,N_623);
nand U1040 (N_1040,N_552,N_601);
and U1041 (N_1041,N_806,N_934);
or U1042 (N_1042,N_738,N_833);
and U1043 (N_1043,N_516,N_579);
and U1044 (N_1044,N_845,N_759);
and U1045 (N_1045,N_692,N_854);
nand U1046 (N_1046,N_655,N_744);
or U1047 (N_1047,N_591,N_704);
nor U1048 (N_1048,N_784,N_633);
nor U1049 (N_1049,N_961,N_667);
and U1050 (N_1050,N_761,N_977);
nand U1051 (N_1051,N_802,N_792);
and U1052 (N_1052,N_804,N_815);
nor U1053 (N_1053,N_526,N_723);
nor U1054 (N_1054,N_779,N_571);
or U1055 (N_1055,N_644,N_699);
or U1056 (N_1056,N_636,N_540);
xnor U1057 (N_1057,N_505,N_922);
and U1058 (N_1058,N_735,N_612);
nand U1059 (N_1059,N_943,N_535);
nand U1060 (N_1060,N_793,N_836);
nor U1061 (N_1061,N_564,N_510);
nor U1062 (N_1062,N_893,N_754);
nor U1063 (N_1063,N_605,N_890);
and U1064 (N_1064,N_868,N_853);
or U1065 (N_1065,N_646,N_944);
nand U1066 (N_1066,N_740,N_967);
xnor U1067 (N_1067,N_884,N_620);
nor U1068 (N_1068,N_525,N_995);
and U1069 (N_1069,N_963,N_715);
nand U1070 (N_1070,N_598,N_518);
or U1071 (N_1071,N_882,N_508);
nor U1072 (N_1072,N_596,N_992);
or U1073 (N_1073,N_600,N_568);
nor U1074 (N_1074,N_835,N_808);
or U1075 (N_1075,N_933,N_594);
and U1076 (N_1076,N_900,N_631);
xnor U1077 (N_1077,N_671,N_517);
or U1078 (N_1078,N_639,N_917);
nor U1079 (N_1079,N_844,N_687);
and U1080 (N_1080,N_617,N_700);
nand U1081 (N_1081,N_787,N_606);
and U1082 (N_1082,N_653,N_569);
or U1083 (N_1083,N_732,N_883);
or U1084 (N_1084,N_968,N_662);
xnor U1085 (N_1085,N_515,N_627);
nor U1086 (N_1086,N_805,N_901);
nor U1087 (N_1087,N_899,N_743);
and U1088 (N_1088,N_728,N_980);
nor U1089 (N_1089,N_885,N_597);
nor U1090 (N_1090,N_725,N_790);
and U1091 (N_1091,N_860,N_755);
or U1092 (N_1092,N_708,N_576);
and U1093 (N_1093,N_775,N_865);
or U1094 (N_1094,N_921,N_826);
nand U1095 (N_1095,N_814,N_816);
or U1096 (N_1096,N_820,N_769);
and U1097 (N_1097,N_717,N_688);
nor U1098 (N_1098,N_710,N_773);
nor U1099 (N_1099,N_991,N_734);
nand U1100 (N_1100,N_749,N_999);
nand U1101 (N_1101,N_788,N_770);
and U1102 (N_1102,N_513,N_765);
or U1103 (N_1103,N_543,N_693);
xor U1104 (N_1104,N_807,N_670);
or U1105 (N_1105,N_645,N_918);
or U1106 (N_1106,N_932,N_955);
nor U1107 (N_1107,N_610,N_829);
nor U1108 (N_1108,N_998,N_837);
nand U1109 (N_1109,N_698,N_970);
nor U1110 (N_1110,N_685,N_642);
nor U1111 (N_1111,N_979,N_953);
nand U1112 (N_1112,N_705,N_827);
nand U1113 (N_1113,N_959,N_663);
and U1114 (N_1114,N_501,N_866);
nor U1115 (N_1115,N_539,N_511);
or U1116 (N_1116,N_586,N_810);
and U1117 (N_1117,N_873,N_771);
and U1118 (N_1118,N_843,N_630);
nor U1119 (N_1119,N_548,N_647);
nor U1120 (N_1120,N_621,N_842);
and U1121 (N_1121,N_971,N_652);
or U1122 (N_1122,N_941,N_811);
nand U1123 (N_1123,N_729,N_949);
and U1124 (N_1124,N_628,N_972);
nor U1125 (N_1125,N_733,N_896);
nand U1126 (N_1126,N_731,N_924);
or U1127 (N_1127,N_862,N_607);
nand U1128 (N_1128,N_574,N_824);
or U1129 (N_1129,N_506,N_903);
nor U1130 (N_1130,N_696,N_783);
nor U1131 (N_1131,N_947,N_776);
nor U1132 (N_1132,N_712,N_825);
nor U1133 (N_1133,N_672,N_919);
nand U1134 (N_1134,N_881,N_519);
or U1135 (N_1135,N_859,N_602);
or U1136 (N_1136,N_928,N_915);
and U1137 (N_1137,N_679,N_994);
and U1138 (N_1138,N_969,N_916);
nor U1139 (N_1139,N_529,N_709);
nand U1140 (N_1140,N_978,N_819);
and U1141 (N_1141,N_931,N_532);
and U1142 (N_1142,N_774,N_509);
nor U1143 (N_1143,N_643,N_849);
nand U1144 (N_1144,N_906,N_938);
or U1145 (N_1145,N_577,N_641);
or U1146 (N_1146,N_780,N_624);
nor U1147 (N_1147,N_946,N_534);
and U1148 (N_1148,N_622,N_907);
or U1149 (N_1149,N_974,N_711);
nor U1150 (N_1150,N_555,N_996);
nor U1151 (N_1151,N_905,N_608);
nand U1152 (N_1152,N_554,N_966);
nor U1153 (N_1153,N_531,N_935);
or U1154 (N_1154,N_960,N_632);
nand U1155 (N_1155,N_936,N_742);
or U1156 (N_1156,N_544,N_822);
nand U1157 (N_1157,N_616,N_657);
or U1158 (N_1158,N_852,N_739);
and U1159 (N_1159,N_879,N_520);
or U1160 (N_1160,N_745,N_990);
nor U1161 (N_1161,N_649,N_986);
nor U1162 (N_1162,N_841,N_888);
or U1163 (N_1163,N_595,N_923);
nor U1164 (N_1164,N_791,N_611);
or U1165 (N_1165,N_690,N_981);
nor U1166 (N_1166,N_795,N_997);
or U1167 (N_1167,N_942,N_737);
or U1168 (N_1168,N_660,N_948);
and U1169 (N_1169,N_718,N_547);
or U1170 (N_1170,N_588,N_801);
and U1171 (N_1171,N_951,N_800);
or U1172 (N_1172,N_925,N_584);
nand U1173 (N_1173,N_678,N_590);
nand U1174 (N_1174,N_987,N_656);
nand U1175 (N_1175,N_777,N_870);
nand U1176 (N_1176,N_929,N_898);
or U1177 (N_1177,N_560,N_983);
nor U1178 (N_1178,N_830,N_551);
and U1179 (N_1179,N_989,N_832);
nand U1180 (N_1180,N_887,N_702);
nor U1181 (N_1181,N_686,N_582);
and U1182 (N_1182,N_831,N_580);
and U1183 (N_1183,N_625,N_619);
and U1184 (N_1184,N_681,N_701);
or U1185 (N_1185,N_993,N_719);
nand U1186 (N_1186,N_863,N_975);
nor U1187 (N_1187,N_658,N_877);
and U1188 (N_1188,N_813,N_926);
and U1189 (N_1189,N_985,N_675);
and U1190 (N_1190,N_604,N_524);
and U1191 (N_1191,N_798,N_895);
nor U1192 (N_1192,N_772,N_542);
nor U1193 (N_1193,N_741,N_550);
nor U1194 (N_1194,N_558,N_861);
nand U1195 (N_1195,N_695,N_716);
and U1196 (N_1196,N_891,N_812);
nor U1197 (N_1197,N_880,N_864);
and U1198 (N_1198,N_984,N_654);
or U1199 (N_1199,N_914,N_911);
or U1200 (N_1200,N_847,N_973);
nand U1201 (N_1201,N_838,N_629);
nor U1202 (N_1202,N_572,N_682);
or U1203 (N_1203,N_762,N_538);
nand U1204 (N_1204,N_857,N_958);
and U1205 (N_1205,N_565,N_615);
or U1206 (N_1206,N_541,N_573);
or U1207 (N_1207,N_856,N_930);
nand U1208 (N_1208,N_567,N_587);
or U1209 (N_1209,N_676,N_724);
nand U1210 (N_1210,N_794,N_562);
and U1211 (N_1211,N_613,N_522);
nor U1212 (N_1212,N_982,N_527);
xnor U1213 (N_1213,N_674,N_648);
nor U1214 (N_1214,N_823,N_954);
and U1215 (N_1215,N_673,N_683);
nand U1216 (N_1216,N_713,N_876);
xnor U1217 (N_1217,N_846,N_747);
nand U1218 (N_1218,N_886,N_618);
and U1219 (N_1219,N_758,N_839);
nand U1220 (N_1220,N_727,N_634);
and U1221 (N_1221,N_500,N_680);
or U1222 (N_1222,N_797,N_760);
nand U1223 (N_1223,N_872,N_897);
nand U1224 (N_1224,N_720,N_561);
nand U1225 (N_1225,N_514,N_521);
or U1226 (N_1226,N_638,N_593);
and U1227 (N_1227,N_848,N_669);
or U1228 (N_1228,N_559,N_650);
nand U1229 (N_1229,N_850,N_523);
nand U1230 (N_1230,N_768,N_689);
or U1231 (N_1231,N_583,N_537);
xnor U1232 (N_1232,N_748,N_666);
and U1233 (N_1233,N_691,N_964);
nand U1234 (N_1234,N_664,N_753);
nand U1235 (N_1235,N_785,N_763);
nor U1236 (N_1236,N_913,N_902);
or U1237 (N_1237,N_840,N_904);
and U1238 (N_1238,N_789,N_828);
and U1239 (N_1239,N_533,N_962);
and U1240 (N_1240,N_809,N_640);
or U1241 (N_1241,N_722,N_609);
nand U1242 (N_1242,N_950,N_767);
xor U1243 (N_1243,N_937,N_756);
and U1244 (N_1244,N_910,N_874);
or U1245 (N_1245,N_952,N_752);
nand U1246 (N_1246,N_592,N_677);
nor U1247 (N_1247,N_589,N_585);
nor U1248 (N_1248,N_503,N_778);
nand U1249 (N_1249,N_988,N_927);
nor U1250 (N_1250,N_779,N_985);
nand U1251 (N_1251,N_820,N_904);
nor U1252 (N_1252,N_869,N_995);
and U1253 (N_1253,N_832,N_638);
and U1254 (N_1254,N_616,N_942);
nand U1255 (N_1255,N_911,N_559);
nand U1256 (N_1256,N_953,N_727);
nor U1257 (N_1257,N_567,N_991);
and U1258 (N_1258,N_511,N_816);
nor U1259 (N_1259,N_548,N_535);
nand U1260 (N_1260,N_819,N_934);
nand U1261 (N_1261,N_535,N_557);
nand U1262 (N_1262,N_578,N_911);
nand U1263 (N_1263,N_850,N_772);
and U1264 (N_1264,N_765,N_710);
or U1265 (N_1265,N_865,N_838);
nor U1266 (N_1266,N_745,N_593);
nand U1267 (N_1267,N_653,N_999);
nand U1268 (N_1268,N_528,N_602);
nor U1269 (N_1269,N_749,N_968);
nor U1270 (N_1270,N_687,N_710);
nor U1271 (N_1271,N_616,N_627);
and U1272 (N_1272,N_899,N_939);
nand U1273 (N_1273,N_592,N_662);
or U1274 (N_1274,N_891,N_589);
nor U1275 (N_1275,N_850,N_998);
nor U1276 (N_1276,N_888,N_683);
nor U1277 (N_1277,N_791,N_533);
nor U1278 (N_1278,N_663,N_591);
xnor U1279 (N_1279,N_547,N_572);
nand U1280 (N_1280,N_885,N_870);
or U1281 (N_1281,N_902,N_511);
and U1282 (N_1282,N_676,N_867);
nor U1283 (N_1283,N_928,N_520);
and U1284 (N_1284,N_803,N_914);
and U1285 (N_1285,N_615,N_825);
nand U1286 (N_1286,N_947,N_980);
or U1287 (N_1287,N_652,N_791);
nor U1288 (N_1288,N_851,N_692);
nand U1289 (N_1289,N_945,N_836);
nor U1290 (N_1290,N_648,N_785);
nand U1291 (N_1291,N_547,N_563);
nand U1292 (N_1292,N_774,N_584);
or U1293 (N_1293,N_817,N_922);
nor U1294 (N_1294,N_818,N_879);
and U1295 (N_1295,N_806,N_631);
nor U1296 (N_1296,N_632,N_558);
or U1297 (N_1297,N_744,N_687);
or U1298 (N_1298,N_945,N_732);
nand U1299 (N_1299,N_723,N_781);
nor U1300 (N_1300,N_964,N_893);
nand U1301 (N_1301,N_532,N_884);
nand U1302 (N_1302,N_851,N_717);
and U1303 (N_1303,N_582,N_886);
nand U1304 (N_1304,N_774,N_910);
xnor U1305 (N_1305,N_940,N_623);
nor U1306 (N_1306,N_919,N_845);
nand U1307 (N_1307,N_563,N_637);
and U1308 (N_1308,N_883,N_650);
nor U1309 (N_1309,N_657,N_510);
nand U1310 (N_1310,N_636,N_606);
and U1311 (N_1311,N_923,N_701);
and U1312 (N_1312,N_888,N_933);
or U1313 (N_1313,N_653,N_947);
nand U1314 (N_1314,N_685,N_630);
and U1315 (N_1315,N_843,N_731);
and U1316 (N_1316,N_740,N_732);
nand U1317 (N_1317,N_781,N_646);
and U1318 (N_1318,N_953,N_572);
or U1319 (N_1319,N_858,N_973);
or U1320 (N_1320,N_952,N_895);
nor U1321 (N_1321,N_949,N_621);
nor U1322 (N_1322,N_938,N_781);
or U1323 (N_1323,N_661,N_888);
nand U1324 (N_1324,N_524,N_659);
nor U1325 (N_1325,N_695,N_831);
or U1326 (N_1326,N_763,N_754);
and U1327 (N_1327,N_851,N_963);
or U1328 (N_1328,N_786,N_686);
nor U1329 (N_1329,N_565,N_717);
nand U1330 (N_1330,N_885,N_651);
nand U1331 (N_1331,N_569,N_716);
nor U1332 (N_1332,N_964,N_560);
nor U1333 (N_1333,N_530,N_941);
nor U1334 (N_1334,N_954,N_940);
nor U1335 (N_1335,N_548,N_855);
and U1336 (N_1336,N_835,N_736);
or U1337 (N_1337,N_559,N_672);
nor U1338 (N_1338,N_881,N_837);
or U1339 (N_1339,N_673,N_556);
and U1340 (N_1340,N_632,N_580);
and U1341 (N_1341,N_619,N_878);
nor U1342 (N_1342,N_729,N_512);
or U1343 (N_1343,N_918,N_745);
nor U1344 (N_1344,N_579,N_998);
and U1345 (N_1345,N_961,N_630);
nor U1346 (N_1346,N_835,N_758);
nor U1347 (N_1347,N_900,N_740);
nand U1348 (N_1348,N_777,N_742);
and U1349 (N_1349,N_666,N_949);
nor U1350 (N_1350,N_953,N_964);
nand U1351 (N_1351,N_524,N_780);
or U1352 (N_1352,N_719,N_872);
nand U1353 (N_1353,N_700,N_749);
nand U1354 (N_1354,N_932,N_634);
and U1355 (N_1355,N_574,N_601);
nor U1356 (N_1356,N_794,N_963);
and U1357 (N_1357,N_872,N_567);
and U1358 (N_1358,N_659,N_504);
and U1359 (N_1359,N_988,N_920);
nor U1360 (N_1360,N_844,N_961);
or U1361 (N_1361,N_619,N_918);
or U1362 (N_1362,N_857,N_819);
or U1363 (N_1363,N_520,N_872);
or U1364 (N_1364,N_979,N_726);
nor U1365 (N_1365,N_867,N_549);
xnor U1366 (N_1366,N_774,N_700);
and U1367 (N_1367,N_825,N_984);
nor U1368 (N_1368,N_737,N_725);
and U1369 (N_1369,N_520,N_585);
nand U1370 (N_1370,N_847,N_937);
or U1371 (N_1371,N_537,N_715);
nor U1372 (N_1372,N_933,N_568);
and U1373 (N_1373,N_577,N_549);
or U1374 (N_1374,N_724,N_683);
nand U1375 (N_1375,N_923,N_952);
nand U1376 (N_1376,N_613,N_880);
and U1377 (N_1377,N_978,N_694);
and U1378 (N_1378,N_774,N_758);
or U1379 (N_1379,N_695,N_730);
and U1380 (N_1380,N_958,N_659);
or U1381 (N_1381,N_517,N_917);
nand U1382 (N_1382,N_994,N_861);
nor U1383 (N_1383,N_677,N_821);
or U1384 (N_1384,N_693,N_847);
nor U1385 (N_1385,N_553,N_656);
or U1386 (N_1386,N_730,N_779);
xnor U1387 (N_1387,N_900,N_552);
or U1388 (N_1388,N_843,N_563);
or U1389 (N_1389,N_836,N_750);
and U1390 (N_1390,N_825,N_626);
nand U1391 (N_1391,N_782,N_695);
nand U1392 (N_1392,N_578,N_559);
nor U1393 (N_1393,N_993,N_654);
or U1394 (N_1394,N_875,N_660);
nor U1395 (N_1395,N_637,N_500);
and U1396 (N_1396,N_847,N_957);
nand U1397 (N_1397,N_540,N_660);
xnor U1398 (N_1398,N_847,N_948);
nand U1399 (N_1399,N_707,N_962);
or U1400 (N_1400,N_566,N_643);
and U1401 (N_1401,N_839,N_664);
nor U1402 (N_1402,N_776,N_610);
or U1403 (N_1403,N_822,N_993);
and U1404 (N_1404,N_774,N_582);
nor U1405 (N_1405,N_719,N_953);
or U1406 (N_1406,N_521,N_791);
nand U1407 (N_1407,N_574,N_657);
and U1408 (N_1408,N_978,N_762);
nor U1409 (N_1409,N_852,N_939);
and U1410 (N_1410,N_603,N_634);
and U1411 (N_1411,N_531,N_765);
nand U1412 (N_1412,N_998,N_629);
and U1413 (N_1413,N_934,N_999);
nand U1414 (N_1414,N_983,N_514);
or U1415 (N_1415,N_794,N_570);
and U1416 (N_1416,N_500,N_700);
and U1417 (N_1417,N_958,N_847);
or U1418 (N_1418,N_770,N_797);
or U1419 (N_1419,N_859,N_788);
or U1420 (N_1420,N_534,N_803);
nor U1421 (N_1421,N_595,N_677);
nor U1422 (N_1422,N_631,N_831);
and U1423 (N_1423,N_760,N_829);
nor U1424 (N_1424,N_865,N_943);
nor U1425 (N_1425,N_642,N_835);
nor U1426 (N_1426,N_868,N_513);
or U1427 (N_1427,N_988,N_880);
or U1428 (N_1428,N_718,N_822);
or U1429 (N_1429,N_978,N_783);
or U1430 (N_1430,N_634,N_599);
nor U1431 (N_1431,N_592,N_646);
nor U1432 (N_1432,N_502,N_984);
nor U1433 (N_1433,N_613,N_658);
and U1434 (N_1434,N_964,N_939);
nand U1435 (N_1435,N_864,N_645);
and U1436 (N_1436,N_602,N_697);
and U1437 (N_1437,N_922,N_616);
nand U1438 (N_1438,N_989,N_741);
nor U1439 (N_1439,N_622,N_989);
and U1440 (N_1440,N_868,N_690);
or U1441 (N_1441,N_566,N_963);
nand U1442 (N_1442,N_828,N_766);
and U1443 (N_1443,N_900,N_927);
nor U1444 (N_1444,N_993,N_998);
nand U1445 (N_1445,N_564,N_995);
xor U1446 (N_1446,N_989,N_572);
or U1447 (N_1447,N_880,N_773);
nand U1448 (N_1448,N_857,N_620);
and U1449 (N_1449,N_664,N_904);
and U1450 (N_1450,N_701,N_892);
and U1451 (N_1451,N_505,N_923);
and U1452 (N_1452,N_562,N_991);
or U1453 (N_1453,N_794,N_645);
or U1454 (N_1454,N_964,N_641);
and U1455 (N_1455,N_500,N_562);
nor U1456 (N_1456,N_611,N_737);
or U1457 (N_1457,N_551,N_824);
nand U1458 (N_1458,N_981,N_581);
and U1459 (N_1459,N_894,N_924);
or U1460 (N_1460,N_738,N_916);
and U1461 (N_1461,N_601,N_908);
or U1462 (N_1462,N_692,N_686);
nand U1463 (N_1463,N_741,N_995);
or U1464 (N_1464,N_760,N_822);
nor U1465 (N_1465,N_734,N_769);
or U1466 (N_1466,N_751,N_667);
nor U1467 (N_1467,N_983,N_524);
nand U1468 (N_1468,N_885,N_874);
nand U1469 (N_1469,N_629,N_902);
or U1470 (N_1470,N_516,N_839);
and U1471 (N_1471,N_999,N_942);
nor U1472 (N_1472,N_863,N_531);
nor U1473 (N_1473,N_518,N_777);
and U1474 (N_1474,N_855,N_797);
or U1475 (N_1475,N_819,N_909);
nand U1476 (N_1476,N_847,N_730);
and U1477 (N_1477,N_798,N_698);
nor U1478 (N_1478,N_561,N_529);
and U1479 (N_1479,N_527,N_521);
nand U1480 (N_1480,N_775,N_846);
nand U1481 (N_1481,N_805,N_839);
or U1482 (N_1482,N_626,N_500);
nand U1483 (N_1483,N_879,N_957);
nor U1484 (N_1484,N_510,N_675);
and U1485 (N_1485,N_800,N_538);
nand U1486 (N_1486,N_787,N_915);
or U1487 (N_1487,N_834,N_503);
or U1488 (N_1488,N_927,N_526);
and U1489 (N_1489,N_631,N_653);
xor U1490 (N_1490,N_622,N_674);
or U1491 (N_1491,N_676,N_928);
or U1492 (N_1492,N_728,N_510);
nor U1493 (N_1493,N_946,N_727);
nand U1494 (N_1494,N_803,N_938);
nor U1495 (N_1495,N_517,N_787);
and U1496 (N_1496,N_779,N_890);
and U1497 (N_1497,N_717,N_800);
or U1498 (N_1498,N_511,N_516);
nor U1499 (N_1499,N_640,N_794);
and U1500 (N_1500,N_1226,N_1307);
or U1501 (N_1501,N_1156,N_1193);
nand U1502 (N_1502,N_1013,N_1315);
and U1503 (N_1503,N_1477,N_1475);
or U1504 (N_1504,N_1035,N_1478);
and U1505 (N_1505,N_1474,N_1020);
or U1506 (N_1506,N_1048,N_1420);
or U1507 (N_1507,N_1301,N_1245);
or U1508 (N_1508,N_1361,N_1004);
nand U1509 (N_1509,N_1014,N_1489);
and U1510 (N_1510,N_1170,N_1227);
and U1511 (N_1511,N_1340,N_1370);
nor U1512 (N_1512,N_1224,N_1120);
nand U1513 (N_1513,N_1068,N_1395);
nor U1514 (N_1514,N_1184,N_1263);
nand U1515 (N_1515,N_1481,N_1183);
nor U1516 (N_1516,N_1221,N_1202);
nor U1517 (N_1517,N_1488,N_1169);
and U1518 (N_1518,N_1312,N_1348);
nand U1519 (N_1519,N_1476,N_1285);
nor U1520 (N_1520,N_1492,N_1334);
and U1521 (N_1521,N_1306,N_1253);
nor U1522 (N_1522,N_1335,N_1145);
or U1523 (N_1523,N_1311,N_1103);
and U1524 (N_1524,N_1444,N_1409);
or U1525 (N_1525,N_1007,N_1490);
nor U1526 (N_1526,N_1251,N_1254);
and U1527 (N_1527,N_1295,N_1276);
nand U1528 (N_1528,N_1451,N_1376);
nor U1529 (N_1529,N_1163,N_1213);
nand U1530 (N_1530,N_1327,N_1408);
and U1531 (N_1531,N_1175,N_1282);
and U1532 (N_1532,N_1000,N_1287);
and U1533 (N_1533,N_1324,N_1345);
and U1534 (N_1534,N_1441,N_1344);
xnor U1535 (N_1535,N_1223,N_1003);
and U1536 (N_1536,N_1211,N_1038);
or U1537 (N_1537,N_1450,N_1012);
and U1538 (N_1538,N_1364,N_1466);
nor U1539 (N_1539,N_1473,N_1069);
nand U1540 (N_1540,N_1382,N_1387);
xnor U1541 (N_1541,N_1192,N_1233);
or U1542 (N_1542,N_1375,N_1355);
nor U1543 (N_1543,N_1422,N_1142);
nor U1544 (N_1544,N_1102,N_1427);
or U1545 (N_1545,N_1131,N_1416);
nor U1546 (N_1546,N_1110,N_1021);
nand U1547 (N_1547,N_1162,N_1284);
nand U1548 (N_1548,N_1027,N_1434);
nand U1549 (N_1549,N_1423,N_1132);
and U1550 (N_1550,N_1467,N_1430);
nor U1551 (N_1551,N_1234,N_1199);
and U1552 (N_1552,N_1469,N_1191);
nor U1553 (N_1553,N_1269,N_1201);
nand U1554 (N_1554,N_1052,N_1219);
and U1555 (N_1555,N_1299,N_1290);
and U1556 (N_1556,N_1333,N_1198);
nand U1557 (N_1557,N_1380,N_1262);
nor U1558 (N_1558,N_1238,N_1497);
nor U1559 (N_1559,N_1055,N_1394);
or U1560 (N_1560,N_1229,N_1207);
nand U1561 (N_1561,N_1122,N_1465);
or U1562 (N_1562,N_1124,N_1092);
or U1563 (N_1563,N_1241,N_1030);
xnor U1564 (N_1564,N_1025,N_1396);
nor U1565 (N_1565,N_1417,N_1281);
and U1566 (N_1566,N_1483,N_1329);
or U1567 (N_1567,N_1305,N_1138);
and U1568 (N_1568,N_1240,N_1248);
nand U1569 (N_1569,N_1414,N_1220);
nand U1570 (N_1570,N_1083,N_1051);
nor U1571 (N_1571,N_1249,N_1403);
and U1572 (N_1572,N_1437,N_1339);
nand U1573 (N_1573,N_1017,N_1093);
and U1574 (N_1574,N_1379,N_1082);
and U1575 (N_1575,N_1426,N_1126);
and U1576 (N_1576,N_1112,N_1143);
and U1577 (N_1577,N_1039,N_1428);
nor U1578 (N_1578,N_1129,N_1098);
nor U1579 (N_1579,N_1458,N_1400);
or U1580 (N_1580,N_1010,N_1034);
or U1581 (N_1581,N_1174,N_1018);
nor U1582 (N_1582,N_1372,N_1147);
or U1583 (N_1583,N_1206,N_1009);
or U1584 (N_1584,N_1390,N_1029);
or U1585 (N_1585,N_1040,N_1369);
nand U1586 (N_1586,N_1429,N_1108);
or U1587 (N_1587,N_1036,N_1316);
nand U1588 (N_1588,N_1128,N_1074);
nand U1589 (N_1589,N_1383,N_1259);
and U1590 (N_1590,N_1354,N_1413);
nor U1591 (N_1591,N_1391,N_1065);
and U1592 (N_1592,N_1480,N_1002);
nand U1593 (N_1593,N_1215,N_1117);
and U1594 (N_1594,N_1062,N_1454);
xnor U1595 (N_1595,N_1255,N_1178);
or U1596 (N_1596,N_1288,N_1078);
nor U1597 (N_1597,N_1067,N_1137);
nand U1598 (N_1598,N_1101,N_1231);
nand U1599 (N_1599,N_1165,N_1471);
nand U1600 (N_1600,N_1398,N_1419);
nand U1601 (N_1601,N_1270,N_1278);
and U1602 (N_1602,N_1022,N_1043);
nor U1603 (N_1603,N_1257,N_1144);
nor U1604 (N_1604,N_1080,N_1159);
nor U1605 (N_1605,N_1019,N_1341);
nand U1606 (N_1606,N_1006,N_1059);
nand U1607 (N_1607,N_1457,N_1188);
or U1608 (N_1608,N_1077,N_1258);
nor U1609 (N_1609,N_1111,N_1271);
nor U1610 (N_1610,N_1140,N_1094);
nor U1611 (N_1611,N_1261,N_1182);
and U1612 (N_1612,N_1032,N_1325);
nor U1613 (N_1613,N_1195,N_1001);
and U1614 (N_1614,N_1453,N_1499);
nand U1615 (N_1615,N_1479,N_1304);
and U1616 (N_1616,N_1150,N_1421);
nand U1617 (N_1617,N_1496,N_1113);
or U1618 (N_1618,N_1446,N_1146);
nor U1619 (N_1619,N_1037,N_1330);
nand U1620 (N_1620,N_1091,N_1109);
nor U1621 (N_1621,N_1431,N_1107);
or U1622 (N_1622,N_1296,N_1384);
nor U1623 (N_1623,N_1378,N_1486);
nor U1624 (N_1624,N_1189,N_1320);
and U1625 (N_1625,N_1358,N_1024);
or U1626 (N_1626,N_1141,N_1374);
nand U1627 (N_1627,N_1064,N_1366);
or U1628 (N_1628,N_1106,N_1470);
nand U1629 (N_1629,N_1464,N_1168);
and U1630 (N_1630,N_1205,N_1187);
and U1631 (N_1631,N_1095,N_1468);
or U1632 (N_1632,N_1050,N_1045);
and U1633 (N_1633,N_1256,N_1115);
or U1634 (N_1634,N_1114,N_1322);
and U1635 (N_1635,N_1289,N_1267);
nand U1636 (N_1636,N_1455,N_1432);
nor U1637 (N_1637,N_1268,N_1081);
and U1638 (N_1638,N_1439,N_1151);
or U1639 (N_1639,N_1365,N_1100);
nand U1640 (N_1640,N_1368,N_1237);
and U1641 (N_1641,N_1209,N_1171);
nor U1642 (N_1642,N_1217,N_1449);
or U1643 (N_1643,N_1208,N_1415);
or U1644 (N_1644,N_1389,N_1442);
and U1645 (N_1645,N_1484,N_1196);
nor U1646 (N_1646,N_1186,N_1346);
nand U1647 (N_1647,N_1347,N_1054);
nor U1648 (N_1648,N_1152,N_1338);
or U1649 (N_1649,N_1298,N_1047);
nand U1650 (N_1650,N_1360,N_1185);
nand U1651 (N_1651,N_1090,N_1023);
and U1652 (N_1652,N_1392,N_1216);
nand U1653 (N_1653,N_1239,N_1167);
and U1654 (N_1654,N_1130,N_1097);
nor U1655 (N_1655,N_1359,N_1194);
and U1656 (N_1656,N_1166,N_1046);
nor U1657 (N_1657,N_1401,N_1393);
and U1658 (N_1658,N_1044,N_1066);
or U1659 (N_1659,N_1318,N_1367);
or U1660 (N_1660,N_1272,N_1406);
and U1661 (N_1661,N_1123,N_1433);
nor U1662 (N_1662,N_1008,N_1425);
nor U1663 (N_1663,N_1385,N_1309);
nor U1664 (N_1664,N_1356,N_1179);
nor U1665 (N_1665,N_1149,N_1049);
or U1666 (N_1666,N_1319,N_1321);
nand U1667 (N_1667,N_1031,N_1397);
nand U1668 (N_1668,N_1242,N_1172);
nand U1669 (N_1669,N_1448,N_1214);
nand U1670 (N_1670,N_1134,N_1160);
or U1671 (N_1671,N_1352,N_1063);
or U1672 (N_1672,N_1314,N_1087);
or U1673 (N_1673,N_1088,N_1399);
nand U1674 (N_1674,N_1494,N_1294);
xnor U1675 (N_1675,N_1228,N_1181);
xor U1676 (N_1676,N_1438,N_1323);
or U1677 (N_1677,N_1053,N_1212);
nand U1678 (N_1678,N_1243,N_1161);
or U1679 (N_1679,N_1084,N_1412);
nand U1680 (N_1680,N_1332,N_1197);
nand U1681 (N_1681,N_1061,N_1337);
nand U1682 (N_1682,N_1459,N_1353);
nor U1683 (N_1683,N_1070,N_1203);
nor U1684 (N_1684,N_1073,N_1351);
nor U1685 (N_1685,N_1292,N_1099);
nor U1686 (N_1686,N_1157,N_1498);
or U1687 (N_1687,N_1283,N_1447);
or U1688 (N_1688,N_1331,N_1440);
nand U1689 (N_1689,N_1461,N_1300);
nand U1690 (N_1690,N_1279,N_1176);
nand U1691 (N_1691,N_1072,N_1487);
or U1692 (N_1692,N_1033,N_1133);
nor U1693 (N_1693,N_1005,N_1028);
and U1694 (N_1694,N_1491,N_1139);
xor U1695 (N_1695,N_1404,N_1230);
or U1696 (N_1696,N_1302,N_1058);
or U1697 (N_1697,N_1011,N_1472);
nand U1698 (N_1698,N_1244,N_1260);
or U1699 (N_1699,N_1264,N_1158);
or U1700 (N_1700,N_1411,N_1357);
or U1701 (N_1701,N_1456,N_1291);
and U1702 (N_1702,N_1200,N_1342);
nor U1703 (N_1703,N_1155,N_1060);
nor U1704 (N_1704,N_1086,N_1085);
or U1705 (N_1705,N_1293,N_1362);
nand U1706 (N_1706,N_1460,N_1273);
and U1707 (N_1707,N_1326,N_1116);
xnor U1708 (N_1708,N_1232,N_1445);
nor U1709 (N_1709,N_1328,N_1482);
nor U1710 (N_1710,N_1435,N_1317);
and U1711 (N_1711,N_1225,N_1042);
and U1712 (N_1712,N_1096,N_1056);
and U1713 (N_1713,N_1218,N_1173);
and U1714 (N_1714,N_1308,N_1075);
nor U1715 (N_1715,N_1121,N_1371);
or U1716 (N_1716,N_1136,N_1105);
nor U1717 (N_1717,N_1089,N_1127);
nor U1718 (N_1718,N_1015,N_1402);
nor U1719 (N_1719,N_1462,N_1280);
nand U1720 (N_1720,N_1071,N_1222);
or U1721 (N_1721,N_1016,N_1373);
nand U1722 (N_1722,N_1154,N_1235);
and U1723 (N_1723,N_1204,N_1310);
xor U1724 (N_1724,N_1125,N_1135);
nor U1725 (N_1725,N_1407,N_1119);
nand U1726 (N_1726,N_1436,N_1493);
and U1727 (N_1727,N_1041,N_1313);
or U1728 (N_1728,N_1190,N_1265);
nand U1729 (N_1729,N_1343,N_1303);
nand U1730 (N_1730,N_1388,N_1452);
nand U1731 (N_1731,N_1118,N_1252);
nand U1732 (N_1732,N_1349,N_1405);
and U1733 (N_1733,N_1079,N_1286);
nor U1734 (N_1734,N_1418,N_1495);
and U1735 (N_1735,N_1424,N_1210);
nand U1736 (N_1736,N_1410,N_1386);
and U1737 (N_1737,N_1236,N_1266);
or U1738 (N_1738,N_1485,N_1246);
nand U1739 (N_1739,N_1297,N_1463);
or U1740 (N_1740,N_1350,N_1177);
and U1741 (N_1741,N_1057,N_1336);
nor U1742 (N_1742,N_1180,N_1153);
or U1743 (N_1743,N_1076,N_1148);
and U1744 (N_1744,N_1274,N_1250);
nand U1745 (N_1745,N_1443,N_1363);
and U1746 (N_1746,N_1247,N_1104);
or U1747 (N_1747,N_1164,N_1275);
or U1748 (N_1748,N_1277,N_1381);
nor U1749 (N_1749,N_1026,N_1377);
and U1750 (N_1750,N_1484,N_1288);
and U1751 (N_1751,N_1163,N_1395);
nor U1752 (N_1752,N_1063,N_1054);
or U1753 (N_1753,N_1167,N_1353);
nand U1754 (N_1754,N_1041,N_1286);
and U1755 (N_1755,N_1140,N_1119);
and U1756 (N_1756,N_1483,N_1127);
and U1757 (N_1757,N_1142,N_1252);
and U1758 (N_1758,N_1173,N_1419);
nand U1759 (N_1759,N_1368,N_1334);
nand U1760 (N_1760,N_1494,N_1195);
nor U1761 (N_1761,N_1290,N_1106);
nand U1762 (N_1762,N_1378,N_1146);
and U1763 (N_1763,N_1009,N_1197);
nor U1764 (N_1764,N_1197,N_1022);
or U1765 (N_1765,N_1304,N_1156);
xnor U1766 (N_1766,N_1304,N_1237);
nor U1767 (N_1767,N_1381,N_1379);
and U1768 (N_1768,N_1086,N_1040);
nand U1769 (N_1769,N_1162,N_1042);
and U1770 (N_1770,N_1019,N_1301);
or U1771 (N_1771,N_1391,N_1142);
nand U1772 (N_1772,N_1474,N_1140);
or U1773 (N_1773,N_1160,N_1046);
nor U1774 (N_1774,N_1492,N_1037);
or U1775 (N_1775,N_1371,N_1451);
or U1776 (N_1776,N_1164,N_1369);
and U1777 (N_1777,N_1127,N_1466);
and U1778 (N_1778,N_1342,N_1201);
and U1779 (N_1779,N_1131,N_1268);
or U1780 (N_1780,N_1086,N_1460);
nor U1781 (N_1781,N_1435,N_1165);
or U1782 (N_1782,N_1015,N_1312);
xnor U1783 (N_1783,N_1190,N_1419);
and U1784 (N_1784,N_1007,N_1001);
nor U1785 (N_1785,N_1153,N_1319);
and U1786 (N_1786,N_1415,N_1292);
nor U1787 (N_1787,N_1179,N_1125);
and U1788 (N_1788,N_1393,N_1293);
nand U1789 (N_1789,N_1365,N_1004);
and U1790 (N_1790,N_1076,N_1490);
nand U1791 (N_1791,N_1094,N_1190);
nand U1792 (N_1792,N_1339,N_1406);
nand U1793 (N_1793,N_1409,N_1387);
and U1794 (N_1794,N_1472,N_1058);
xnor U1795 (N_1795,N_1014,N_1480);
and U1796 (N_1796,N_1384,N_1387);
nand U1797 (N_1797,N_1347,N_1223);
or U1798 (N_1798,N_1480,N_1460);
nor U1799 (N_1799,N_1155,N_1440);
and U1800 (N_1800,N_1287,N_1217);
or U1801 (N_1801,N_1435,N_1480);
nor U1802 (N_1802,N_1337,N_1139);
xnor U1803 (N_1803,N_1012,N_1116);
and U1804 (N_1804,N_1491,N_1486);
nor U1805 (N_1805,N_1458,N_1179);
xnor U1806 (N_1806,N_1236,N_1330);
nand U1807 (N_1807,N_1120,N_1236);
nor U1808 (N_1808,N_1201,N_1145);
and U1809 (N_1809,N_1249,N_1067);
or U1810 (N_1810,N_1124,N_1228);
or U1811 (N_1811,N_1447,N_1344);
nor U1812 (N_1812,N_1340,N_1249);
nor U1813 (N_1813,N_1088,N_1026);
and U1814 (N_1814,N_1407,N_1040);
or U1815 (N_1815,N_1000,N_1022);
nor U1816 (N_1816,N_1150,N_1320);
and U1817 (N_1817,N_1380,N_1077);
nand U1818 (N_1818,N_1065,N_1119);
and U1819 (N_1819,N_1360,N_1201);
and U1820 (N_1820,N_1490,N_1091);
or U1821 (N_1821,N_1049,N_1186);
nand U1822 (N_1822,N_1149,N_1295);
and U1823 (N_1823,N_1310,N_1381);
nor U1824 (N_1824,N_1189,N_1104);
nor U1825 (N_1825,N_1233,N_1310);
nand U1826 (N_1826,N_1339,N_1491);
nor U1827 (N_1827,N_1093,N_1171);
nand U1828 (N_1828,N_1339,N_1307);
nand U1829 (N_1829,N_1036,N_1384);
nand U1830 (N_1830,N_1127,N_1479);
nor U1831 (N_1831,N_1095,N_1331);
nand U1832 (N_1832,N_1205,N_1459);
nand U1833 (N_1833,N_1061,N_1166);
nor U1834 (N_1834,N_1150,N_1039);
and U1835 (N_1835,N_1420,N_1319);
and U1836 (N_1836,N_1345,N_1159);
and U1837 (N_1837,N_1421,N_1242);
and U1838 (N_1838,N_1362,N_1023);
or U1839 (N_1839,N_1049,N_1012);
nand U1840 (N_1840,N_1484,N_1057);
and U1841 (N_1841,N_1070,N_1465);
nand U1842 (N_1842,N_1053,N_1313);
and U1843 (N_1843,N_1375,N_1230);
and U1844 (N_1844,N_1392,N_1294);
nand U1845 (N_1845,N_1024,N_1008);
and U1846 (N_1846,N_1262,N_1371);
and U1847 (N_1847,N_1122,N_1010);
nand U1848 (N_1848,N_1208,N_1032);
xor U1849 (N_1849,N_1050,N_1235);
and U1850 (N_1850,N_1194,N_1261);
nand U1851 (N_1851,N_1402,N_1428);
nand U1852 (N_1852,N_1427,N_1275);
and U1853 (N_1853,N_1491,N_1377);
nand U1854 (N_1854,N_1128,N_1000);
and U1855 (N_1855,N_1111,N_1108);
and U1856 (N_1856,N_1045,N_1182);
nand U1857 (N_1857,N_1003,N_1465);
nor U1858 (N_1858,N_1305,N_1396);
or U1859 (N_1859,N_1227,N_1268);
nor U1860 (N_1860,N_1124,N_1114);
nand U1861 (N_1861,N_1410,N_1140);
nand U1862 (N_1862,N_1048,N_1196);
or U1863 (N_1863,N_1096,N_1323);
xnor U1864 (N_1864,N_1067,N_1337);
nor U1865 (N_1865,N_1351,N_1081);
xnor U1866 (N_1866,N_1377,N_1359);
or U1867 (N_1867,N_1066,N_1286);
nor U1868 (N_1868,N_1295,N_1357);
nand U1869 (N_1869,N_1494,N_1360);
nor U1870 (N_1870,N_1162,N_1499);
nand U1871 (N_1871,N_1346,N_1221);
nor U1872 (N_1872,N_1007,N_1383);
nand U1873 (N_1873,N_1404,N_1251);
and U1874 (N_1874,N_1262,N_1460);
nor U1875 (N_1875,N_1036,N_1487);
nor U1876 (N_1876,N_1388,N_1292);
and U1877 (N_1877,N_1465,N_1019);
or U1878 (N_1878,N_1286,N_1410);
or U1879 (N_1879,N_1219,N_1287);
nand U1880 (N_1880,N_1172,N_1303);
nor U1881 (N_1881,N_1129,N_1475);
nor U1882 (N_1882,N_1275,N_1110);
xor U1883 (N_1883,N_1292,N_1026);
or U1884 (N_1884,N_1003,N_1036);
or U1885 (N_1885,N_1066,N_1006);
and U1886 (N_1886,N_1320,N_1273);
and U1887 (N_1887,N_1230,N_1014);
nand U1888 (N_1888,N_1224,N_1129);
and U1889 (N_1889,N_1141,N_1019);
and U1890 (N_1890,N_1150,N_1054);
and U1891 (N_1891,N_1059,N_1400);
or U1892 (N_1892,N_1016,N_1441);
nor U1893 (N_1893,N_1081,N_1361);
nand U1894 (N_1894,N_1025,N_1242);
nor U1895 (N_1895,N_1209,N_1388);
nand U1896 (N_1896,N_1256,N_1048);
and U1897 (N_1897,N_1180,N_1095);
nor U1898 (N_1898,N_1478,N_1095);
or U1899 (N_1899,N_1484,N_1407);
nor U1900 (N_1900,N_1240,N_1095);
or U1901 (N_1901,N_1311,N_1238);
or U1902 (N_1902,N_1350,N_1468);
or U1903 (N_1903,N_1032,N_1180);
xnor U1904 (N_1904,N_1285,N_1052);
nor U1905 (N_1905,N_1085,N_1434);
or U1906 (N_1906,N_1100,N_1208);
nor U1907 (N_1907,N_1476,N_1461);
xor U1908 (N_1908,N_1364,N_1287);
nor U1909 (N_1909,N_1155,N_1062);
nand U1910 (N_1910,N_1028,N_1385);
or U1911 (N_1911,N_1143,N_1342);
nand U1912 (N_1912,N_1394,N_1364);
and U1913 (N_1913,N_1366,N_1154);
and U1914 (N_1914,N_1327,N_1183);
or U1915 (N_1915,N_1037,N_1223);
or U1916 (N_1916,N_1154,N_1064);
or U1917 (N_1917,N_1467,N_1157);
nand U1918 (N_1918,N_1464,N_1116);
and U1919 (N_1919,N_1359,N_1067);
and U1920 (N_1920,N_1041,N_1036);
xor U1921 (N_1921,N_1313,N_1451);
or U1922 (N_1922,N_1035,N_1410);
and U1923 (N_1923,N_1494,N_1368);
and U1924 (N_1924,N_1026,N_1190);
nand U1925 (N_1925,N_1099,N_1020);
and U1926 (N_1926,N_1426,N_1387);
nand U1927 (N_1927,N_1321,N_1136);
and U1928 (N_1928,N_1495,N_1267);
and U1929 (N_1929,N_1193,N_1423);
or U1930 (N_1930,N_1025,N_1263);
and U1931 (N_1931,N_1404,N_1129);
nand U1932 (N_1932,N_1360,N_1018);
or U1933 (N_1933,N_1305,N_1183);
or U1934 (N_1934,N_1491,N_1395);
and U1935 (N_1935,N_1311,N_1287);
nor U1936 (N_1936,N_1233,N_1392);
and U1937 (N_1937,N_1413,N_1048);
nor U1938 (N_1938,N_1048,N_1387);
nor U1939 (N_1939,N_1350,N_1277);
and U1940 (N_1940,N_1356,N_1186);
and U1941 (N_1941,N_1342,N_1177);
nand U1942 (N_1942,N_1267,N_1178);
and U1943 (N_1943,N_1492,N_1080);
nor U1944 (N_1944,N_1204,N_1451);
nand U1945 (N_1945,N_1429,N_1136);
nand U1946 (N_1946,N_1232,N_1084);
nor U1947 (N_1947,N_1051,N_1380);
nor U1948 (N_1948,N_1269,N_1410);
nand U1949 (N_1949,N_1464,N_1302);
and U1950 (N_1950,N_1465,N_1279);
and U1951 (N_1951,N_1180,N_1393);
and U1952 (N_1952,N_1025,N_1191);
and U1953 (N_1953,N_1217,N_1245);
or U1954 (N_1954,N_1403,N_1002);
nor U1955 (N_1955,N_1089,N_1004);
and U1956 (N_1956,N_1465,N_1448);
and U1957 (N_1957,N_1383,N_1133);
and U1958 (N_1958,N_1233,N_1488);
nor U1959 (N_1959,N_1369,N_1473);
nand U1960 (N_1960,N_1379,N_1355);
and U1961 (N_1961,N_1459,N_1462);
or U1962 (N_1962,N_1036,N_1390);
nand U1963 (N_1963,N_1150,N_1417);
nor U1964 (N_1964,N_1181,N_1196);
nand U1965 (N_1965,N_1061,N_1282);
nand U1966 (N_1966,N_1055,N_1233);
and U1967 (N_1967,N_1138,N_1447);
or U1968 (N_1968,N_1149,N_1217);
nor U1969 (N_1969,N_1197,N_1226);
and U1970 (N_1970,N_1118,N_1068);
and U1971 (N_1971,N_1258,N_1254);
nor U1972 (N_1972,N_1034,N_1076);
or U1973 (N_1973,N_1263,N_1125);
nand U1974 (N_1974,N_1042,N_1466);
nand U1975 (N_1975,N_1085,N_1234);
nand U1976 (N_1976,N_1175,N_1304);
and U1977 (N_1977,N_1072,N_1362);
nor U1978 (N_1978,N_1095,N_1028);
nand U1979 (N_1979,N_1066,N_1119);
and U1980 (N_1980,N_1182,N_1210);
or U1981 (N_1981,N_1402,N_1358);
nand U1982 (N_1982,N_1334,N_1150);
nand U1983 (N_1983,N_1109,N_1252);
and U1984 (N_1984,N_1442,N_1482);
nand U1985 (N_1985,N_1371,N_1130);
or U1986 (N_1986,N_1474,N_1009);
and U1987 (N_1987,N_1356,N_1406);
or U1988 (N_1988,N_1489,N_1052);
or U1989 (N_1989,N_1482,N_1224);
or U1990 (N_1990,N_1254,N_1352);
nor U1991 (N_1991,N_1171,N_1056);
xnor U1992 (N_1992,N_1086,N_1144);
or U1993 (N_1993,N_1046,N_1376);
nor U1994 (N_1994,N_1010,N_1177);
nor U1995 (N_1995,N_1316,N_1339);
nand U1996 (N_1996,N_1358,N_1021);
xnor U1997 (N_1997,N_1109,N_1375);
nor U1998 (N_1998,N_1189,N_1346);
or U1999 (N_1999,N_1212,N_1381);
nand U2000 (N_2000,N_1542,N_1692);
or U2001 (N_2001,N_1585,N_1893);
nor U2002 (N_2002,N_1822,N_1508);
nor U2003 (N_2003,N_1515,N_1629);
nand U2004 (N_2004,N_1906,N_1540);
xnor U2005 (N_2005,N_1850,N_1562);
nor U2006 (N_2006,N_1945,N_1755);
or U2007 (N_2007,N_1593,N_1733);
nor U2008 (N_2008,N_1897,N_1833);
nand U2009 (N_2009,N_1525,N_1617);
or U2010 (N_2010,N_1992,N_1716);
or U2011 (N_2011,N_1913,N_1884);
nand U2012 (N_2012,N_1886,N_1951);
nand U2013 (N_2013,N_1909,N_1854);
nand U2014 (N_2014,N_1547,N_1619);
nand U2015 (N_2015,N_1856,N_1753);
and U2016 (N_2016,N_1598,N_1848);
and U2017 (N_2017,N_1820,N_1663);
nand U2018 (N_2018,N_1538,N_1554);
nand U2019 (N_2019,N_1746,N_1703);
nor U2020 (N_2020,N_1930,N_1679);
and U2021 (N_2021,N_1650,N_1589);
or U2022 (N_2022,N_1803,N_1553);
or U2023 (N_2023,N_1699,N_1918);
or U2024 (N_2024,N_1682,N_1759);
and U2025 (N_2025,N_1828,N_1885);
and U2026 (N_2026,N_1980,N_1684);
nor U2027 (N_2027,N_1747,N_1727);
or U2028 (N_2028,N_1630,N_1997);
nand U2029 (N_2029,N_1739,N_1774);
or U2030 (N_2030,N_1528,N_1652);
nor U2031 (N_2031,N_1714,N_1974);
and U2032 (N_2032,N_1778,N_1505);
and U2033 (N_2033,N_1735,N_1901);
nor U2034 (N_2034,N_1624,N_1844);
or U2035 (N_2035,N_1726,N_1947);
or U2036 (N_2036,N_1892,N_1960);
nand U2037 (N_2037,N_1881,N_1504);
xor U2038 (N_2038,N_1923,N_1622);
nand U2039 (N_2039,N_1842,N_1794);
and U2040 (N_2040,N_1658,N_1745);
nand U2041 (N_2041,N_1738,N_1818);
nand U2042 (N_2042,N_1641,N_1957);
nor U2043 (N_2043,N_1758,N_1744);
and U2044 (N_2044,N_1985,N_1798);
nand U2045 (N_2045,N_1712,N_1823);
nor U2046 (N_2046,N_1648,N_1732);
and U2047 (N_2047,N_1864,N_1868);
nand U2048 (N_2048,N_1793,N_1602);
nand U2049 (N_2049,N_1862,N_1696);
or U2050 (N_2050,N_1565,N_1545);
or U2051 (N_2051,N_1940,N_1995);
nor U2052 (N_2052,N_1730,N_1668);
nand U2053 (N_2053,N_1685,N_1671);
nand U2054 (N_2054,N_1623,N_1888);
xor U2055 (N_2055,N_1950,N_1859);
or U2056 (N_2056,N_1559,N_1757);
nand U2057 (N_2057,N_1556,N_1713);
or U2058 (N_2058,N_1541,N_1601);
and U2059 (N_2059,N_1656,N_1972);
nand U2060 (N_2060,N_1989,N_1688);
and U2061 (N_2061,N_1973,N_1781);
and U2062 (N_2062,N_1825,N_1609);
xor U2063 (N_2063,N_1986,N_1569);
nor U2064 (N_2064,N_1644,N_1555);
or U2065 (N_2065,N_1719,N_1908);
and U2066 (N_2066,N_1795,N_1998);
or U2067 (N_2067,N_1966,N_1912);
and U2068 (N_2068,N_1572,N_1577);
nor U2069 (N_2069,N_1978,N_1865);
or U2070 (N_2070,N_1625,N_1670);
nand U2071 (N_2071,N_1519,N_1568);
and U2072 (N_2072,N_1734,N_1931);
and U2073 (N_2073,N_1988,N_1724);
or U2074 (N_2074,N_1874,N_1999);
and U2075 (N_2075,N_1655,N_1637);
nor U2076 (N_2076,N_1841,N_1900);
or U2077 (N_2077,N_1889,N_1858);
or U2078 (N_2078,N_1707,N_1697);
and U2079 (N_2079,N_1531,N_1829);
nor U2080 (N_2080,N_1635,N_1536);
nand U2081 (N_2081,N_1729,N_1691);
nand U2082 (N_2082,N_1996,N_1835);
or U2083 (N_2083,N_1802,N_1860);
nor U2084 (N_2084,N_1932,N_1706);
nor U2085 (N_2085,N_1870,N_1647);
nor U2086 (N_2086,N_1512,N_1840);
or U2087 (N_2087,N_1937,N_1915);
nand U2088 (N_2088,N_1956,N_1678);
nand U2089 (N_2089,N_1742,N_1968);
or U2090 (N_2090,N_1796,N_1883);
or U2091 (N_2091,N_1552,N_1718);
or U2092 (N_2092,N_1851,N_1632);
nor U2093 (N_2093,N_1643,N_1651);
or U2094 (N_2094,N_1831,N_1693);
nand U2095 (N_2095,N_1741,N_1961);
nor U2096 (N_2096,N_1701,N_1929);
or U2097 (N_2097,N_1958,N_1518);
nor U2098 (N_2098,N_1500,N_1627);
nor U2099 (N_2099,N_1946,N_1920);
nor U2100 (N_2100,N_1587,N_1936);
and U2101 (N_2101,N_1584,N_1959);
nand U2102 (N_2102,N_1836,N_1723);
nand U2103 (N_2103,N_1927,N_1938);
or U2104 (N_2104,N_1610,N_1580);
or U2105 (N_2105,N_1922,N_1673);
nand U2106 (N_2106,N_1866,N_1548);
nand U2107 (N_2107,N_1847,N_1967);
and U2108 (N_2108,N_1816,N_1677);
or U2109 (N_2109,N_1766,N_1586);
nor U2110 (N_2110,N_1775,N_1837);
nor U2111 (N_2111,N_1705,N_1722);
nor U2112 (N_2112,N_1815,N_1522);
nand U2113 (N_2113,N_1633,N_1964);
nand U2114 (N_2114,N_1575,N_1827);
nor U2115 (N_2115,N_1832,N_1567);
nor U2116 (N_2116,N_1771,N_1812);
or U2117 (N_2117,N_1549,N_1975);
or U2118 (N_2118,N_1579,N_1942);
or U2119 (N_2119,N_1516,N_1857);
nor U2120 (N_2120,N_1948,N_1954);
nand U2121 (N_2121,N_1869,N_1953);
and U2122 (N_2122,N_1955,N_1578);
nand U2123 (N_2123,N_1507,N_1910);
nand U2124 (N_2124,N_1702,N_1895);
and U2125 (N_2125,N_1700,N_1590);
nor U2126 (N_2126,N_1600,N_1506);
nand U2127 (N_2127,N_1916,N_1924);
nor U2128 (N_2128,N_1604,N_1620);
nor U2129 (N_2129,N_1941,N_1904);
or U2130 (N_2130,N_1736,N_1830);
nor U2131 (N_2131,N_1606,N_1596);
nand U2132 (N_2132,N_1546,N_1704);
or U2133 (N_2133,N_1800,N_1517);
or U2134 (N_2134,N_1560,N_1843);
and U2135 (N_2135,N_1898,N_1896);
nor U2136 (N_2136,N_1717,N_1939);
or U2137 (N_2137,N_1709,N_1510);
or U2138 (N_2138,N_1711,N_1534);
nor U2139 (N_2139,N_1708,N_1573);
nor U2140 (N_2140,N_1819,N_1981);
or U2141 (N_2141,N_1838,N_1676);
nor U2142 (N_2142,N_1595,N_1807);
nor U2143 (N_2143,N_1934,N_1698);
nor U2144 (N_2144,N_1666,N_1907);
nand U2145 (N_2145,N_1867,N_1921);
and U2146 (N_2146,N_1750,N_1839);
nand U2147 (N_2147,N_1943,N_1790);
nor U2148 (N_2148,N_1715,N_1965);
and U2149 (N_2149,N_1817,N_1571);
or U2150 (N_2150,N_1821,N_1765);
or U2151 (N_2151,N_1994,N_1982);
nand U2152 (N_2152,N_1944,N_1654);
nor U2153 (N_2153,N_1880,N_1680);
nand U2154 (N_2154,N_1566,N_1903);
nor U2155 (N_2155,N_1879,N_1513);
or U2156 (N_2156,N_1523,N_1877);
nand U2157 (N_2157,N_1532,N_1887);
or U2158 (N_2158,N_1582,N_1770);
nand U2159 (N_2159,N_1613,N_1768);
or U2160 (N_2160,N_1614,N_1626);
or U2161 (N_2161,N_1902,N_1791);
nor U2162 (N_2162,N_1890,N_1861);
nor U2163 (N_2163,N_1777,N_1977);
nand U2164 (N_2164,N_1645,N_1761);
or U2165 (N_2165,N_1675,N_1588);
and U2166 (N_2166,N_1792,N_1751);
nor U2167 (N_2167,N_1634,N_1526);
nor U2168 (N_2168,N_1611,N_1524);
nor U2169 (N_2169,N_1612,N_1826);
nor U2170 (N_2170,N_1756,N_1681);
or U2171 (N_2171,N_1592,N_1824);
nand U2172 (N_2172,N_1721,N_1871);
and U2173 (N_2173,N_1799,N_1882);
nand U2174 (N_2174,N_1917,N_1845);
nand U2175 (N_2175,N_1686,N_1811);
nor U2176 (N_2176,N_1689,N_1748);
nand U2177 (N_2177,N_1605,N_1878);
nand U2178 (N_2178,N_1984,N_1603);
or U2179 (N_2179,N_1749,N_1608);
nand U2180 (N_2180,N_1511,N_1661);
xor U2181 (N_2181,N_1616,N_1804);
nor U2182 (N_2182,N_1769,N_1963);
and U2183 (N_2183,N_1638,N_1783);
nor U2184 (N_2184,N_1782,N_1754);
or U2185 (N_2185,N_1779,N_1853);
and U2186 (N_2186,N_1894,N_1583);
nor U2187 (N_2187,N_1952,N_1971);
nor U2188 (N_2188,N_1914,N_1520);
and U2189 (N_2189,N_1657,N_1659);
nand U2190 (N_2190,N_1502,N_1615);
and U2191 (N_2191,N_1646,N_1808);
and U2192 (N_2192,N_1660,N_1695);
nand U2193 (N_2193,N_1551,N_1983);
or U2194 (N_2194,N_1899,N_1780);
nor U2195 (N_2195,N_1962,N_1872);
nor U2196 (N_2196,N_1762,N_1852);
or U2197 (N_2197,N_1797,N_1683);
and U2198 (N_2198,N_1905,N_1607);
and U2199 (N_2199,N_1876,N_1725);
nand U2200 (N_2200,N_1529,N_1537);
nand U2201 (N_2201,N_1558,N_1649);
and U2202 (N_2202,N_1667,N_1535);
nand U2203 (N_2203,N_1581,N_1662);
nor U2204 (N_2204,N_1576,N_1514);
and U2205 (N_2205,N_1891,N_1653);
nor U2206 (N_2206,N_1786,N_1849);
nor U2207 (N_2207,N_1533,N_1925);
and U2208 (N_2208,N_1669,N_1687);
nand U2209 (N_2209,N_1784,N_1846);
and U2210 (N_2210,N_1809,N_1911);
nand U2211 (N_2211,N_1501,N_1991);
xor U2212 (N_2212,N_1919,N_1789);
and U2213 (N_2213,N_1935,N_1564);
or U2214 (N_2214,N_1574,N_1767);
nand U2215 (N_2215,N_1949,N_1743);
nor U2216 (N_2216,N_1801,N_1806);
and U2217 (N_2217,N_1665,N_1970);
and U2218 (N_2218,N_1503,N_1550);
and U2219 (N_2219,N_1664,N_1763);
nor U2220 (N_2220,N_1530,N_1834);
nand U2221 (N_2221,N_1599,N_1672);
or U2222 (N_2222,N_1570,N_1776);
or U2223 (N_2223,N_1787,N_1591);
and U2224 (N_2224,N_1631,N_1764);
or U2225 (N_2225,N_1527,N_1788);
nor U2226 (N_2226,N_1594,N_1979);
and U2227 (N_2227,N_1543,N_1875);
and U2228 (N_2228,N_1928,N_1993);
and U2229 (N_2229,N_1731,N_1636);
or U2230 (N_2230,N_1728,N_1628);
nor U2231 (N_2231,N_1720,N_1752);
and U2232 (N_2232,N_1539,N_1813);
and U2233 (N_2233,N_1740,N_1814);
and U2234 (N_2234,N_1805,N_1737);
nor U2235 (N_2235,N_1557,N_1710);
nand U2236 (N_2236,N_1639,N_1561);
and U2237 (N_2237,N_1863,N_1810);
or U2238 (N_2238,N_1773,N_1674);
and U2239 (N_2239,N_1642,N_1873);
or U2240 (N_2240,N_1563,N_1509);
and U2241 (N_2241,N_1760,N_1621);
nand U2242 (N_2242,N_1521,N_1969);
and U2243 (N_2243,N_1926,N_1690);
nand U2244 (N_2244,N_1976,N_1785);
nor U2245 (N_2245,N_1544,N_1640);
nor U2246 (N_2246,N_1694,N_1990);
nor U2247 (N_2247,N_1597,N_1855);
and U2248 (N_2248,N_1772,N_1987);
nor U2249 (N_2249,N_1618,N_1933);
and U2250 (N_2250,N_1635,N_1657);
nor U2251 (N_2251,N_1963,N_1639);
and U2252 (N_2252,N_1610,N_1948);
or U2253 (N_2253,N_1622,N_1880);
nor U2254 (N_2254,N_1845,N_1872);
and U2255 (N_2255,N_1868,N_1878);
and U2256 (N_2256,N_1764,N_1758);
or U2257 (N_2257,N_1867,N_1854);
or U2258 (N_2258,N_1769,N_1971);
or U2259 (N_2259,N_1960,N_1835);
nor U2260 (N_2260,N_1669,N_1504);
and U2261 (N_2261,N_1657,N_1594);
or U2262 (N_2262,N_1765,N_1912);
and U2263 (N_2263,N_1563,N_1637);
and U2264 (N_2264,N_1513,N_1971);
or U2265 (N_2265,N_1852,N_1721);
nor U2266 (N_2266,N_1529,N_1508);
or U2267 (N_2267,N_1603,N_1907);
nand U2268 (N_2268,N_1942,N_1912);
nand U2269 (N_2269,N_1998,N_1617);
nor U2270 (N_2270,N_1899,N_1853);
or U2271 (N_2271,N_1627,N_1745);
and U2272 (N_2272,N_1726,N_1890);
and U2273 (N_2273,N_1684,N_1905);
nor U2274 (N_2274,N_1684,N_1896);
nand U2275 (N_2275,N_1686,N_1981);
and U2276 (N_2276,N_1706,N_1813);
nor U2277 (N_2277,N_1807,N_1814);
nand U2278 (N_2278,N_1514,N_1699);
nand U2279 (N_2279,N_1548,N_1948);
and U2280 (N_2280,N_1749,N_1801);
and U2281 (N_2281,N_1679,N_1632);
and U2282 (N_2282,N_1506,N_1548);
nand U2283 (N_2283,N_1775,N_1781);
or U2284 (N_2284,N_1890,N_1731);
and U2285 (N_2285,N_1723,N_1985);
or U2286 (N_2286,N_1684,N_1689);
or U2287 (N_2287,N_1931,N_1840);
nor U2288 (N_2288,N_1928,N_1979);
nor U2289 (N_2289,N_1667,N_1919);
or U2290 (N_2290,N_1592,N_1870);
or U2291 (N_2291,N_1824,N_1503);
or U2292 (N_2292,N_1777,N_1730);
or U2293 (N_2293,N_1989,N_1711);
xor U2294 (N_2294,N_1657,N_1620);
nor U2295 (N_2295,N_1881,N_1959);
and U2296 (N_2296,N_1841,N_1737);
nor U2297 (N_2297,N_1535,N_1556);
and U2298 (N_2298,N_1827,N_1626);
nor U2299 (N_2299,N_1580,N_1624);
nor U2300 (N_2300,N_1573,N_1848);
nand U2301 (N_2301,N_1524,N_1885);
and U2302 (N_2302,N_1993,N_1782);
nand U2303 (N_2303,N_1893,N_1672);
xnor U2304 (N_2304,N_1791,N_1965);
and U2305 (N_2305,N_1998,N_1941);
or U2306 (N_2306,N_1562,N_1930);
nor U2307 (N_2307,N_1607,N_1954);
and U2308 (N_2308,N_1677,N_1947);
nand U2309 (N_2309,N_1680,N_1809);
and U2310 (N_2310,N_1504,N_1574);
xnor U2311 (N_2311,N_1842,N_1697);
nand U2312 (N_2312,N_1571,N_1709);
or U2313 (N_2313,N_1955,N_1678);
and U2314 (N_2314,N_1928,N_1757);
nand U2315 (N_2315,N_1672,N_1882);
nor U2316 (N_2316,N_1729,N_1638);
nor U2317 (N_2317,N_1916,N_1547);
or U2318 (N_2318,N_1952,N_1640);
or U2319 (N_2319,N_1963,N_1710);
nand U2320 (N_2320,N_1897,N_1573);
nand U2321 (N_2321,N_1678,N_1886);
and U2322 (N_2322,N_1963,N_1753);
nand U2323 (N_2323,N_1521,N_1825);
nor U2324 (N_2324,N_1584,N_1512);
nor U2325 (N_2325,N_1940,N_1556);
nor U2326 (N_2326,N_1852,N_1573);
nand U2327 (N_2327,N_1886,N_1838);
or U2328 (N_2328,N_1870,N_1654);
or U2329 (N_2329,N_1846,N_1951);
and U2330 (N_2330,N_1963,N_1733);
nor U2331 (N_2331,N_1873,N_1684);
or U2332 (N_2332,N_1747,N_1721);
or U2333 (N_2333,N_1747,N_1537);
and U2334 (N_2334,N_1772,N_1829);
and U2335 (N_2335,N_1734,N_1949);
nand U2336 (N_2336,N_1787,N_1822);
and U2337 (N_2337,N_1659,N_1941);
and U2338 (N_2338,N_1974,N_1792);
or U2339 (N_2339,N_1525,N_1544);
or U2340 (N_2340,N_1566,N_1852);
and U2341 (N_2341,N_1906,N_1618);
xnor U2342 (N_2342,N_1990,N_1585);
and U2343 (N_2343,N_1719,N_1847);
and U2344 (N_2344,N_1750,N_1612);
and U2345 (N_2345,N_1917,N_1567);
xor U2346 (N_2346,N_1568,N_1872);
nor U2347 (N_2347,N_1519,N_1971);
nor U2348 (N_2348,N_1873,N_1756);
nor U2349 (N_2349,N_1787,N_1625);
nor U2350 (N_2350,N_1571,N_1664);
and U2351 (N_2351,N_1996,N_1566);
or U2352 (N_2352,N_1601,N_1887);
or U2353 (N_2353,N_1557,N_1583);
and U2354 (N_2354,N_1841,N_1870);
nor U2355 (N_2355,N_1551,N_1786);
nand U2356 (N_2356,N_1590,N_1731);
and U2357 (N_2357,N_1843,N_1680);
or U2358 (N_2358,N_1785,N_1886);
or U2359 (N_2359,N_1600,N_1585);
or U2360 (N_2360,N_1582,N_1850);
nor U2361 (N_2361,N_1597,N_1790);
or U2362 (N_2362,N_1702,N_1615);
nor U2363 (N_2363,N_1526,N_1755);
and U2364 (N_2364,N_1906,N_1576);
nor U2365 (N_2365,N_1500,N_1870);
nand U2366 (N_2366,N_1550,N_1885);
nor U2367 (N_2367,N_1563,N_1541);
and U2368 (N_2368,N_1725,N_1786);
nor U2369 (N_2369,N_1653,N_1936);
or U2370 (N_2370,N_1960,N_1519);
and U2371 (N_2371,N_1744,N_1799);
and U2372 (N_2372,N_1787,N_1885);
and U2373 (N_2373,N_1758,N_1625);
and U2374 (N_2374,N_1633,N_1939);
or U2375 (N_2375,N_1964,N_1800);
nand U2376 (N_2376,N_1636,N_1748);
nand U2377 (N_2377,N_1735,N_1654);
nor U2378 (N_2378,N_1909,N_1877);
or U2379 (N_2379,N_1650,N_1948);
nand U2380 (N_2380,N_1561,N_1563);
nor U2381 (N_2381,N_1981,N_1517);
nor U2382 (N_2382,N_1896,N_1659);
or U2383 (N_2383,N_1656,N_1996);
or U2384 (N_2384,N_1893,N_1645);
nor U2385 (N_2385,N_1870,N_1549);
nand U2386 (N_2386,N_1744,N_1807);
nand U2387 (N_2387,N_1925,N_1711);
nor U2388 (N_2388,N_1907,N_1875);
or U2389 (N_2389,N_1939,N_1953);
or U2390 (N_2390,N_1981,N_1612);
or U2391 (N_2391,N_1894,N_1764);
or U2392 (N_2392,N_1681,N_1838);
and U2393 (N_2393,N_1514,N_1550);
nor U2394 (N_2394,N_1709,N_1927);
nor U2395 (N_2395,N_1728,N_1686);
nor U2396 (N_2396,N_1799,N_1504);
or U2397 (N_2397,N_1869,N_1504);
or U2398 (N_2398,N_1894,N_1544);
and U2399 (N_2399,N_1673,N_1595);
nand U2400 (N_2400,N_1577,N_1961);
nor U2401 (N_2401,N_1710,N_1778);
and U2402 (N_2402,N_1807,N_1758);
nand U2403 (N_2403,N_1688,N_1752);
nand U2404 (N_2404,N_1645,N_1910);
and U2405 (N_2405,N_1986,N_1751);
nand U2406 (N_2406,N_1975,N_1984);
and U2407 (N_2407,N_1919,N_1830);
and U2408 (N_2408,N_1853,N_1638);
nor U2409 (N_2409,N_1906,N_1623);
or U2410 (N_2410,N_1817,N_1645);
and U2411 (N_2411,N_1600,N_1580);
or U2412 (N_2412,N_1865,N_1596);
nor U2413 (N_2413,N_1588,N_1785);
nand U2414 (N_2414,N_1723,N_1774);
nor U2415 (N_2415,N_1941,N_1969);
or U2416 (N_2416,N_1918,N_1645);
or U2417 (N_2417,N_1506,N_1707);
nand U2418 (N_2418,N_1926,N_1593);
nand U2419 (N_2419,N_1766,N_1755);
or U2420 (N_2420,N_1606,N_1947);
nand U2421 (N_2421,N_1557,N_1625);
or U2422 (N_2422,N_1790,N_1691);
and U2423 (N_2423,N_1588,N_1848);
and U2424 (N_2424,N_1792,N_1932);
or U2425 (N_2425,N_1792,N_1925);
and U2426 (N_2426,N_1632,N_1886);
nor U2427 (N_2427,N_1789,N_1879);
xnor U2428 (N_2428,N_1626,N_1671);
and U2429 (N_2429,N_1537,N_1954);
or U2430 (N_2430,N_1918,N_1737);
nand U2431 (N_2431,N_1537,N_1870);
nor U2432 (N_2432,N_1600,N_1708);
nand U2433 (N_2433,N_1756,N_1648);
and U2434 (N_2434,N_1804,N_1757);
or U2435 (N_2435,N_1781,N_1742);
or U2436 (N_2436,N_1822,N_1902);
xor U2437 (N_2437,N_1530,N_1934);
and U2438 (N_2438,N_1945,N_1672);
or U2439 (N_2439,N_1888,N_1713);
or U2440 (N_2440,N_1914,N_1856);
nor U2441 (N_2441,N_1628,N_1518);
or U2442 (N_2442,N_1561,N_1617);
nand U2443 (N_2443,N_1584,N_1865);
or U2444 (N_2444,N_1576,N_1969);
nand U2445 (N_2445,N_1771,N_1903);
nand U2446 (N_2446,N_1834,N_1870);
or U2447 (N_2447,N_1625,N_1937);
nand U2448 (N_2448,N_1555,N_1649);
nand U2449 (N_2449,N_1712,N_1930);
or U2450 (N_2450,N_1988,N_1868);
nand U2451 (N_2451,N_1674,N_1511);
nand U2452 (N_2452,N_1823,N_1587);
or U2453 (N_2453,N_1909,N_1918);
nor U2454 (N_2454,N_1806,N_1575);
or U2455 (N_2455,N_1652,N_1735);
and U2456 (N_2456,N_1510,N_1989);
or U2457 (N_2457,N_1530,N_1899);
nor U2458 (N_2458,N_1674,N_1527);
xnor U2459 (N_2459,N_1615,N_1598);
or U2460 (N_2460,N_1686,N_1848);
and U2461 (N_2461,N_1813,N_1867);
nor U2462 (N_2462,N_1557,N_1649);
nor U2463 (N_2463,N_1632,N_1557);
or U2464 (N_2464,N_1727,N_1761);
nor U2465 (N_2465,N_1865,N_1693);
nor U2466 (N_2466,N_1661,N_1568);
or U2467 (N_2467,N_1856,N_1797);
nor U2468 (N_2468,N_1588,N_1727);
nand U2469 (N_2469,N_1876,N_1755);
nor U2470 (N_2470,N_1825,N_1632);
and U2471 (N_2471,N_1713,N_1922);
and U2472 (N_2472,N_1543,N_1821);
nand U2473 (N_2473,N_1648,N_1849);
and U2474 (N_2474,N_1830,N_1857);
nand U2475 (N_2475,N_1555,N_1695);
and U2476 (N_2476,N_1653,N_1972);
nor U2477 (N_2477,N_1854,N_1774);
and U2478 (N_2478,N_1970,N_1792);
nor U2479 (N_2479,N_1960,N_1807);
nand U2480 (N_2480,N_1956,N_1776);
and U2481 (N_2481,N_1714,N_1600);
nand U2482 (N_2482,N_1508,N_1712);
xnor U2483 (N_2483,N_1615,N_1571);
nor U2484 (N_2484,N_1547,N_1545);
and U2485 (N_2485,N_1720,N_1524);
and U2486 (N_2486,N_1949,N_1887);
nor U2487 (N_2487,N_1585,N_1839);
and U2488 (N_2488,N_1598,N_1523);
nor U2489 (N_2489,N_1573,N_1687);
nand U2490 (N_2490,N_1987,N_1602);
nor U2491 (N_2491,N_1611,N_1676);
or U2492 (N_2492,N_1868,N_1950);
or U2493 (N_2493,N_1607,N_1648);
nand U2494 (N_2494,N_1835,N_1909);
and U2495 (N_2495,N_1634,N_1792);
or U2496 (N_2496,N_1750,N_1768);
nor U2497 (N_2497,N_1986,N_1992);
or U2498 (N_2498,N_1663,N_1536);
nand U2499 (N_2499,N_1959,N_1975);
and U2500 (N_2500,N_2464,N_2395);
nor U2501 (N_2501,N_2090,N_2081);
nor U2502 (N_2502,N_2293,N_2486);
nor U2503 (N_2503,N_2260,N_2118);
or U2504 (N_2504,N_2229,N_2275);
nand U2505 (N_2505,N_2431,N_2218);
or U2506 (N_2506,N_2310,N_2455);
or U2507 (N_2507,N_2454,N_2378);
or U2508 (N_2508,N_2141,N_2242);
nand U2509 (N_2509,N_2052,N_2091);
or U2510 (N_2510,N_2371,N_2366);
nand U2511 (N_2511,N_2369,N_2024);
nor U2512 (N_2512,N_2042,N_2194);
or U2513 (N_2513,N_2421,N_2397);
nand U2514 (N_2514,N_2410,N_2234);
and U2515 (N_2515,N_2450,N_2465);
or U2516 (N_2516,N_2349,N_2403);
and U2517 (N_2517,N_2282,N_2094);
and U2518 (N_2518,N_2105,N_2168);
or U2519 (N_2519,N_2128,N_2343);
nor U2520 (N_2520,N_2429,N_2083);
or U2521 (N_2521,N_2205,N_2364);
nor U2522 (N_2522,N_2393,N_2273);
or U2523 (N_2523,N_2233,N_2174);
nand U2524 (N_2524,N_2279,N_2276);
nand U2525 (N_2525,N_2108,N_2101);
or U2526 (N_2526,N_2157,N_2184);
and U2527 (N_2527,N_2250,N_2338);
nand U2528 (N_2528,N_2190,N_2207);
and U2529 (N_2529,N_2312,N_2341);
and U2530 (N_2530,N_2147,N_2002);
or U2531 (N_2531,N_2448,N_2295);
or U2532 (N_2532,N_2228,N_2358);
and U2533 (N_2533,N_2466,N_2380);
nand U2534 (N_2534,N_2309,N_2163);
and U2535 (N_2535,N_2236,N_2398);
and U2536 (N_2536,N_2331,N_2473);
nand U2537 (N_2537,N_2483,N_2495);
nand U2538 (N_2538,N_2212,N_2497);
or U2539 (N_2539,N_2107,N_2082);
nor U2540 (N_2540,N_2173,N_2475);
or U2541 (N_2541,N_2254,N_2478);
nor U2542 (N_2542,N_2326,N_2332);
or U2543 (N_2543,N_2158,N_2209);
or U2544 (N_2544,N_2425,N_2359);
and U2545 (N_2545,N_2400,N_2405);
nand U2546 (N_2546,N_2306,N_2285);
or U2547 (N_2547,N_2381,N_2015);
nand U2548 (N_2548,N_2409,N_2492);
nor U2549 (N_2549,N_2045,N_2166);
or U2550 (N_2550,N_2010,N_2489);
nor U2551 (N_2551,N_2152,N_2058);
and U2552 (N_2552,N_2027,N_2078);
nand U2553 (N_2553,N_2014,N_2135);
or U2554 (N_2554,N_2253,N_2076);
nand U2555 (N_2555,N_2440,N_2368);
nand U2556 (N_2556,N_2021,N_2385);
nor U2557 (N_2557,N_2424,N_2308);
xnor U2558 (N_2558,N_2204,N_2386);
nor U2559 (N_2559,N_2017,N_2472);
nor U2560 (N_2560,N_2235,N_2133);
and U2561 (N_2561,N_2456,N_2336);
or U2562 (N_2562,N_2469,N_2185);
nand U2563 (N_2563,N_2065,N_2446);
or U2564 (N_2564,N_2041,N_2323);
nand U2565 (N_2565,N_2384,N_2019);
nor U2566 (N_2566,N_2420,N_2264);
nor U2567 (N_2567,N_2334,N_2480);
nand U2568 (N_2568,N_2137,N_2297);
nor U2569 (N_2569,N_2004,N_2413);
nor U2570 (N_2570,N_2060,N_2084);
or U2571 (N_2571,N_2283,N_2307);
and U2572 (N_2572,N_2354,N_2022);
or U2573 (N_2573,N_2357,N_2311);
or U2574 (N_2574,N_2217,N_2088);
nor U2575 (N_2575,N_2415,N_2039);
or U2576 (N_2576,N_2374,N_2330);
nand U2577 (N_2577,N_2281,N_2302);
or U2578 (N_2578,N_2070,N_2224);
nand U2579 (N_2579,N_2248,N_2117);
xor U2580 (N_2580,N_2411,N_2116);
nor U2581 (N_2581,N_2051,N_2167);
or U2582 (N_2582,N_2121,N_2222);
and U2583 (N_2583,N_2300,N_2151);
nand U2584 (N_2584,N_2016,N_2267);
nor U2585 (N_2585,N_2046,N_2468);
and U2586 (N_2586,N_2054,N_2200);
and U2587 (N_2587,N_2098,N_2289);
and U2588 (N_2588,N_2050,N_2037);
and U2589 (N_2589,N_2073,N_2164);
and U2590 (N_2590,N_2048,N_2013);
nor U2591 (N_2591,N_2396,N_2035);
and U2592 (N_2592,N_2232,N_2442);
nand U2593 (N_2593,N_2294,N_2467);
or U2594 (N_2594,N_2443,N_2487);
nand U2595 (N_2595,N_2290,N_2485);
nor U2596 (N_2596,N_2372,N_2043);
nand U2597 (N_2597,N_2033,N_2159);
and U2598 (N_2598,N_2437,N_2100);
nand U2599 (N_2599,N_2303,N_2064);
and U2600 (N_2600,N_2461,N_2176);
nand U2601 (N_2601,N_2006,N_2053);
nand U2602 (N_2602,N_2191,N_2412);
nand U2603 (N_2603,N_2156,N_2320);
or U2604 (N_2604,N_2149,N_2179);
nor U2605 (N_2605,N_2195,N_2109);
nor U2606 (N_2606,N_2143,N_2382);
and U2607 (N_2607,N_2401,N_2139);
xor U2608 (N_2608,N_2251,N_2186);
nand U2609 (N_2609,N_2089,N_2047);
or U2610 (N_2610,N_2056,N_2460);
xnor U2611 (N_2611,N_2238,N_2085);
nand U2612 (N_2612,N_2278,N_2171);
or U2613 (N_2613,N_2146,N_2361);
nand U2614 (N_2614,N_2348,N_2444);
and U2615 (N_2615,N_2230,N_2243);
nor U2616 (N_2616,N_2430,N_2001);
or U2617 (N_2617,N_2114,N_2169);
nor U2618 (N_2618,N_2106,N_2129);
xor U2619 (N_2619,N_2202,N_2075);
nor U2620 (N_2620,N_2203,N_2291);
and U2621 (N_2621,N_2427,N_2000);
nand U2622 (N_2622,N_2339,N_2445);
nand U2623 (N_2623,N_2032,N_2245);
nor U2624 (N_2624,N_2170,N_2009);
nand U2625 (N_2625,N_2376,N_2426);
and U2626 (N_2626,N_2069,N_2287);
nand U2627 (N_2627,N_2189,N_2180);
and U2628 (N_2628,N_2482,N_2274);
and U2629 (N_2629,N_2178,N_2315);
and U2630 (N_2630,N_2417,N_2272);
or U2631 (N_2631,N_2347,N_2246);
and U2632 (N_2632,N_2219,N_2463);
or U2633 (N_2633,N_2447,N_2316);
or U2634 (N_2634,N_2402,N_2288);
xnor U2635 (N_2635,N_2277,N_2317);
nand U2636 (N_2636,N_2335,N_2220);
nand U2637 (N_2637,N_2110,N_2365);
nand U2638 (N_2638,N_2433,N_2130);
and U2639 (N_2639,N_2122,N_2057);
nor U2640 (N_2640,N_2153,N_2241);
nor U2641 (N_2641,N_2408,N_2353);
nand U2642 (N_2642,N_2007,N_2406);
nand U2643 (N_2643,N_2265,N_2329);
or U2644 (N_2644,N_2328,N_2011);
or U2645 (N_2645,N_2136,N_2025);
or U2646 (N_2646,N_2154,N_2177);
nand U2647 (N_2647,N_2257,N_2476);
nand U2648 (N_2648,N_2140,N_2499);
nand U2649 (N_2649,N_2240,N_2459);
and U2650 (N_2650,N_2390,N_2034);
nor U2651 (N_2651,N_2113,N_2115);
and U2652 (N_2652,N_2175,N_2252);
nor U2653 (N_2653,N_2367,N_2138);
nor U2654 (N_2654,N_2418,N_2271);
nor U2655 (N_2655,N_2355,N_2350);
and U2656 (N_2656,N_2301,N_2255);
or U2657 (N_2657,N_2484,N_2247);
nand U2658 (N_2658,N_2181,N_2155);
and U2659 (N_2659,N_2077,N_2481);
and U2660 (N_2660,N_2342,N_2352);
and U2661 (N_2661,N_2221,N_2008);
nand U2662 (N_2662,N_2457,N_2063);
nor U2663 (N_2663,N_2183,N_2362);
nand U2664 (N_2664,N_2262,N_2225);
and U2665 (N_2665,N_2313,N_2124);
nand U2666 (N_2666,N_2333,N_2496);
and U2667 (N_2667,N_2379,N_2451);
or U2668 (N_2668,N_2258,N_2102);
nand U2669 (N_2669,N_2095,N_2131);
nor U2670 (N_2670,N_2256,N_2375);
nor U2671 (N_2671,N_2389,N_2453);
nor U2672 (N_2672,N_2261,N_2227);
or U2673 (N_2673,N_2068,N_2345);
nor U2674 (N_2674,N_2193,N_2206);
and U2675 (N_2675,N_2211,N_2327);
nor U2676 (N_2676,N_2215,N_2145);
xor U2677 (N_2677,N_2123,N_2160);
nand U2678 (N_2678,N_2340,N_2298);
nand U2679 (N_2679,N_2321,N_2187);
and U2680 (N_2680,N_2391,N_2216);
nor U2681 (N_2681,N_2040,N_2226);
nand U2682 (N_2682,N_2162,N_2049);
nand U2683 (N_2683,N_2286,N_2249);
nor U2684 (N_2684,N_2337,N_2093);
nand U2685 (N_2685,N_2414,N_2432);
nor U2686 (N_2686,N_2055,N_2018);
nand U2687 (N_2687,N_2148,N_2325);
nor U2688 (N_2688,N_2005,N_2498);
and U2689 (N_2689,N_2493,N_2266);
or U2690 (N_2690,N_2299,N_2161);
nor U2691 (N_2691,N_2031,N_2351);
nand U2692 (N_2692,N_2491,N_2423);
nand U2693 (N_2693,N_2404,N_2092);
and U2694 (N_2694,N_2436,N_2003);
and U2695 (N_2695,N_2127,N_2182);
or U2696 (N_2696,N_2059,N_2314);
and U2697 (N_2697,N_2023,N_2012);
or U2698 (N_2698,N_2239,N_2201);
nand U2699 (N_2699,N_2097,N_2213);
nor U2700 (N_2700,N_2237,N_2080);
or U2701 (N_2701,N_2471,N_2479);
nand U2702 (N_2702,N_2086,N_2132);
nor U2703 (N_2703,N_2269,N_2125);
nand U2704 (N_2704,N_2144,N_2488);
nand U2705 (N_2705,N_2087,N_2126);
and U2706 (N_2706,N_2419,N_2304);
nand U2707 (N_2707,N_2120,N_2458);
and U2708 (N_2708,N_2270,N_2363);
or U2709 (N_2709,N_2387,N_2028);
or U2710 (N_2710,N_2020,N_2071);
and U2711 (N_2711,N_2346,N_2263);
nand U2712 (N_2712,N_2165,N_2231);
nor U2713 (N_2713,N_2029,N_2490);
and U2714 (N_2714,N_2038,N_2439);
nand U2715 (N_2715,N_2296,N_2111);
or U2716 (N_2716,N_2199,N_2066);
and U2717 (N_2717,N_2474,N_2356);
and U2718 (N_2718,N_2062,N_2026);
xor U2719 (N_2719,N_2284,N_2192);
nand U2720 (N_2720,N_2434,N_2197);
and U2721 (N_2721,N_2268,N_2305);
nor U2722 (N_2722,N_2388,N_2407);
xnor U2723 (N_2723,N_2099,N_2079);
or U2724 (N_2724,N_2318,N_2208);
or U2725 (N_2725,N_2449,N_2044);
xnor U2726 (N_2726,N_2292,N_2223);
nor U2727 (N_2727,N_2210,N_2074);
or U2728 (N_2728,N_2244,N_2422);
nor U2729 (N_2729,N_2394,N_2259);
and U2730 (N_2730,N_2370,N_2399);
xor U2731 (N_2731,N_2438,N_2462);
nor U2732 (N_2732,N_2119,N_2377);
nor U2733 (N_2733,N_2188,N_2104);
nand U2734 (N_2734,N_2214,N_2344);
nor U2735 (N_2735,N_2172,N_2280);
and U2736 (N_2736,N_2103,N_2067);
and U2737 (N_2737,N_2142,N_2373);
nor U2738 (N_2738,N_2150,N_2435);
nor U2739 (N_2739,N_2477,N_2324);
or U2740 (N_2740,N_2196,N_2416);
nand U2741 (N_2741,N_2061,N_2494);
nor U2742 (N_2742,N_2392,N_2112);
or U2743 (N_2743,N_2319,N_2072);
nand U2744 (N_2744,N_2428,N_2036);
nand U2745 (N_2745,N_2470,N_2030);
nand U2746 (N_2746,N_2360,N_2441);
or U2747 (N_2747,N_2134,N_2322);
or U2748 (N_2748,N_2198,N_2383);
nor U2749 (N_2749,N_2096,N_2452);
or U2750 (N_2750,N_2083,N_2200);
and U2751 (N_2751,N_2243,N_2489);
and U2752 (N_2752,N_2221,N_2276);
nand U2753 (N_2753,N_2256,N_2358);
and U2754 (N_2754,N_2122,N_2315);
nand U2755 (N_2755,N_2318,N_2072);
or U2756 (N_2756,N_2019,N_2169);
or U2757 (N_2757,N_2048,N_2272);
or U2758 (N_2758,N_2140,N_2356);
and U2759 (N_2759,N_2313,N_2304);
and U2760 (N_2760,N_2400,N_2252);
or U2761 (N_2761,N_2497,N_2136);
nand U2762 (N_2762,N_2130,N_2237);
nand U2763 (N_2763,N_2391,N_2318);
nor U2764 (N_2764,N_2182,N_2219);
and U2765 (N_2765,N_2411,N_2181);
xor U2766 (N_2766,N_2101,N_2261);
and U2767 (N_2767,N_2058,N_2299);
nand U2768 (N_2768,N_2120,N_2334);
nand U2769 (N_2769,N_2203,N_2266);
nor U2770 (N_2770,N_2284,N_2366);
nand U2771 (N_2771,N_2418,N_2116);
or U2772 (N_2772,N_2324,N_2240);
nand U2773 (N_2773,N_2233,N_2060);
and U2774 (N_2774,N_2380,N_2113);
nor U2775 (N_2775,N_2158,N_2078);
or U2776 (N_2776,N_2368,N_2377);
or U2777 (N_2777,N_2413,N_2163);
nand U2778 (N_2778,N_2333,N_2123);
nor U2779 (N_2779,N_2021,N_2329);
and U2780 (N_2780,N_2424,N_2047);
or U2781 (N_2781,N_2483,N_2041);
nor U2782 (N_2782,N_2052,N_2276);
and U2783 (N_2783,N_2358,N_2411);
nor U2784 (N_2784,N_2364,N_2186);
and U2785 (N_2785,N_2314,N_2230);
nor U2786 (N_2786,N_2021,N_2304);
nand U2787 (N_2787,N_2381,N_2458);
nor U2788 (N_2788,N_2264,N_2128);
nor U2789 (N_2789,N_2409,N_2456);
nor U2790 (N_2790,N_2204,N_2287);
and U2791 (N_2791,N_2071,N_2406);
nand U2792 (N_2792,N_2270,N_2411);
nand U2793 (N_2793,N_2298,N_2136);
and U2794 (N_2794,N_2362,N_2431);
nand U2795 (N_2795,N_2222,N_2174);
nor U2796 (N_2796,N_2146,N_2201);
nand U2797 (N_2797,N_2355,N_2210);
or U2798 (N_2798,N_2361,N_2007);
and U2799 (N_2799,N_2100,N_2056);
nor U2800 (N_2800,N_2367,N_2405);
and U2801 (N_2801,N_2088,N_2261);
or U2802 (N_2802,N_2295,N_2202);
or U2803 (N_2803,N_2384,N_2464);
nor U2804 (N_2804,N_2120,N_2136);
nor U2805 (N_2805,N_2150,N_2335);
or U2806 (N_2806,N_2021,N_2047);
and U2807 (N_2807,N_2298,N_2122);
nand U2808 (N_2808,N_2426,N_2022);
nand U2809 (N_2809,N_2037,N_2023);
or U2810 (N_2810,N_2129,N_2448);
nor U2811 (N_2811,N_2387,N_2029);
nor U2812 (N_2812,N_2401,N_2498);
or U2813 (N_2813,N_2012,N_2295);
nand U2814 (N_2814,N_2006,N_2169);
and U2815 (N_2815,N_2481,N_2095);
or U2816 (N_2816,N_2196,N_2293);
or U2817 (N_2817,N_2475,N_2176);
nor U2818 (N_2818,N_2496,N_2193);
nor U2819 (N_2819,N_2389,N_2446);
nor U2820 (N_2820,N_2298,N_2242);
nand U2821 (N_2821,N_2421,N_2390);
nor U2822 (N_2822,N_2262,N_2147);
or U2823 (N_2823,N_2045,N_2261);
or U2824 (N_2824,N_2363,N_2070);
nor U2825 (N_2825,N_2367,N_2374);
nand U2826 (N_2826,N_2459,N_2348);
and U2827 (N_2827,N_2302,N_2134);
nor U2828 (N_2828,N_2304,N_2109);
or U2829 (N_2829,N_2217,N_2348);
and U2830 (N_2830,N_2007,N_2017);
and U2831 (N_2831,N_2284,N_2169);
and U2832 (N_2832,N_2136,N_2010);
nor U2833 (N_2833,N_2017,N_2246);
nand U2834 (N_2834,N_2299,N_2383);
nor U2835 (N_2835,N_2148,N_2232);
nor U2836 (N_2836,N_2182,N_2471);
and U2837 (N_2837,N_2409,N_2149);
or U2838 (N_2838,N_2163,N_2014);
and U2839 (N_2839,N_2016,N_2494);
or U2840 (N_2840,N_2022,N_2351);
nor U2841 (N_2841,N_2041,N_2447);
or U2842 (N_2842,N_2398,N_2447);
nor U2843 (N_2843,N_2358,N_2055);
and U2844 (N_2844,N_2467,N_2105);
and U2845 (N_2845,N_2021,N_2228);
and U2846 (N_2846,N_2073,N_2017);
and U2847 (N_2847,N_2325,N_2038);
and U2848 (N_2848,N_2362,N_2248);
nor U2849 (N_2849,N_2307,N_2178);
xor U2850 (N_2850,N_2229,N_2385);
or U2851 (N_2851,N_2017,N_2434);
or U2852 (N_2852,N_2284,N_2091);
nor U2853 (N_2853,N_2391,N_2112);
or U2854 (N_2854,N_2235,N_2485);
or U2855 (N_2855,N_2410,N_2210);
and U2856 (N_2856,N_2210,N_2198);
nand U2857 (N_2857,N_2298,N_2094);
and U2858 (N_2858,N_2246,N_2061);
and U2859 (N_2859,N_2388,N_2341);
nor U2860 (N_2860,N_2047,N_2426);
and U2861 (N_2861,N_2055,N_2222);
nor U2862 (N_2862,N_2314,N_2130);
and U2863 (N_2863,N_2455,N_2201);
or U2864 (N_2864,N_2080,N_2457);
xnor U2865 (N_2865,N_2179,N_2486);
nor U2866 (N_2866,N_2028,N_2084);
and U2867 (N_2867,N_2017,N_2381);
nand U2868 (N_2868,N_2452,N_2406);
xnor U2869 (N_2869,N_2400,N_2364);
nand U2870 (N_2870,N_2467,N_2421);
xor U2871 (N_2871,N_2067,N_2309);
and U2872 (N_2872,N_2399,N_2214);
nor U2873 (N_2873,N_2490,N_2434);
or U2874 (N_2874,N_2094,N_2128);
nand U2875 (N_2875,N_2350,N_2120);
nor U2876 (N_2876,N_2333,N_2485);
and U2877 (N_2877,N_2435,N_2224);
nor U2878 (N_2878,N_2386,N_2079);
nor U2879 (N_2879,N_2046,N_2201);
or U2880 (N_2880,N_2225,N_2136);
nor U2881 (N_2881,N_2418,N_2020);
nor U2882 (N_2882,N_2101,N_2226);
nand U2883 (N_2883,N_2075,N_2072);
and U2884 (N_2884,N_2005,N_2053);
and U2885 (N_2885,N_2497,N_2151);
nor U2886 (N_2886,N_2421,N_2238);
or U2887 (N_2887,N_2458,N_2293);
or U2888 (N_2888,N_2152,N_2386);
and U2889 (N_2889,N_2066,N_2043);
or U2890 (N_2890,N_2461,N_2118);
nor U2891 (N_2891,N_2094,N_2181);
nor U2892 (N_2892,N_2019,N_2010);
and U2893 (N_2893,N_2192,N_2328);
nand U2894 (N_2894,N_2391,N_2215);
nand U2895 (N_2895,N_2296,N_2054);
or U2896 (N_2896,N_2248,N_2001);
nand U2897 (N_2897,N_2403,N_2020);
nand U2898 (N_2898,N_2369,N_2067);
and U2899 (N_2899,N_2139,N_2282);
and U2900 (N_2900,N_2153,N_2487);
or U2901 (N_2901,N_2261,N_2180);
nor U2902 (N_2902,N_2145,N_2325);
nand U2903 (N_2903,N_2412,N_2029);
or U2904 (N_2904,N_2396,N_2060);
xor U2905 (N_2905,N_2122,N_2357);
or U2906 (N_2906,N_2210,N_2334);
and U2907 (N_2907,N_2310,N_2437);
and U2908 (N_2908,N_2457,N_2403);
nor U2909 (N_2909,N_2325,N_2127);
and U2910 (N_2910,N_2199,N_2138);
and U2911 (N_2911,N_2311,N_2033);
and U2912 (N_2912,N_2106,N_2183);
nand U2913 (N_2913,N_2307,N_2076);
and U2914 (N_2914,N_2379,N_2013);
nand U2915 (N_2915,N_2463,N_2488);
or U2916 (N_2916,N_2483,N_2297);
nor U2917 (N_2917,N_2269,N_2097);
or U2918 (N_2918,N_2376,N_2432);
nand U2919 (N_2919,N_2205,N_2336);
xor U2920 (N_2920,N_2109,N_2072);
or U2921 (N_2921,N_2262,N_2066);
or U2922 (N_2922,N_2241,N_2092);
nor U2923 (N_2923,N_2302,N_2119);
and U2924 (N_2924,N_2120,N_2477);
nand U2925 (N_2925,N_2444,N_2431);
or U2926 (N_2926,N_2326,N_2342);
nand U2927 (N_2927,N_2450,N_2206);
or U2928 (N_2928,N_2204,N_2168);
nand U2929 (N_2929,N_2162,N_2337);
and U2930 (N_2930,N_2407,N_2154);
and U2931 (N_2931,N_2460,N_2150);
nor U2932 (N_2932,N_2208,N_2494);
nor U2933 (N_2933,N_2020,N_2121);
nor U2934 (N_2934,N_2260,N_2142);
nand U2935 (N_2935,N_2057,N_2323);
nand U2936 (N_2936,N_2108,N_2107);
or U2937 (N_2937,N_2074,N_2288);
nor U2938 (N_2938,N_2057,N_2498);
nor U2939 (N_2939,N_2363,N_2059);
nand U2940 (N_2940,N_2368,N_2424);
or U2941 (N_2941,N_2357,N_2203);
nor U2942 (N_2942,N_2467,N_2487);
and U2943 (N_2943,N_2297,N_2165);
or U2944 (N_2944,N_2406,N_2055);
nor U2945 (N_2945,N_2314,N_2347);
or U2946 (N_2946,N_2474,N_2461);
or U2947 (N_2947,N_2480,N_2216);
and U2948 (N_2948,N_2223,N_2175);
nor U2949 (N_2949,N_2050,N_2314);
or U2950 (N_2950,N_2369,N_2185);
xnor U2951 (N_2951,N_2236,N_2442);
and U2952 (N_2952,N_2498,N_2105);
and U2953 (N_2953,N_2394,N_2291);
and U2954 (N_2954,N_2195,N_2132);
nand U2955 (N_2955,N_2259,N_2196);
nand U2956 (N_2956,N_2297,N_2333);
nand U2957 (N_2957,N_2473,N_2433);
nand U2958 (N_2958,N_2346,N_2402);
nand U2959 (N_2959,N_2485,N_2202);
or U2960 (N_2960,N_2074,N_2361);
nand U2961 (N_2961,N_2352,N_2423);
and U2962 (N_2962,N_2485,N_2131);
nor U2963 (N_2963,N_2049,N_2438);
nor U2964 (N_2964,N_2373,N_2183);
nor U2965 (N_2965,N_2291,N_2110);
and U2966 (N_2966,N_2284,N_2209);
nand U2967 (N_2967,N_2062,N_2078);
nand U2968 (N_2968,N_2393,N_2478);
and U2969 (N_2969,N_2339,N_2326);
and U2970 (N_2970,N_2404,N_2459);
or U2971 (N_2971,N_2075,N_2081);
or U2972 (N_2972,N_2348,N_2384);
nand U2973 (N_2973,N_2109,N_2490);
or U2974 (N_2974,N_2447,N_2340);
nor U2975 (N_2975,N_2118,N_2355);
nor U2976 (N_2976,N_2250,N_2173);
and U2977 (N_2977,N_2356,N_2142);
nand U2978 (N_2978,N_2275,N_2353);
nand U2979 (N_2979,N_2221,N_2255);
nand U2980 (N_2980,N_2024,N_2164);
or U2981 (N_2981,N_2272,N_2308);
and U2982 (N_2982,N_2305,N_2491);
xor U2983 (N_2983,N_2351,N_2105);
and U2984 (N_2984,N_2406,N_2011);
or U2985 (N_2985,N_2258,N_2152);
nand U2986 (N_2986,N_2193,N_2240);
nor U2987 (N_2987,N_2081,N_2111);
nor U2988 (N_2988,N_2345,N_2108);
or U2989 (N_2989,N_2049,N_2011);
nand U2990 (N_2990,N_2328,N_2388);
xnor U2991 (N_2991,N_2326,N_2385);
or U2992 (N_2992,N_2078,N_2084);
nor U2993 (N_2993,N_2090,N_2470);
nand U2994 (N_2994,N_2306,N_2282);
xor U2995 (N_2995,N_2429,N_2468);
xor U2996 (N_2996,N_2352,N_2422);
or U2997 (N_2997,N_2187,N_2136);
or U2998 (N_2998,N_2130,N_2441);
nand U2999 (N_2999,N_2305,N_2497);
nor U3000 (N_3000,N_2925,N_2623);
nor U3001 (N_3001,N_2602,N_2700);
and U3002 (N_3002,N_2795,N_2807);
nor U3003 (N_3003,N_2546,N_2524);
nand U3004 (N_3004,N_2580,N_2798);
or U3005 (N_3005,N_2965,N_2573);
nand U3006 (N_3006,N_2797,N_2563);
nor U3007 (N_3007,N_2585,N_2599);
and U3008 (N_3008,N_2681,N_2938);
nor U3009 (N_3009,N_2567,N_2901);
nor U3010 (N_3010,N_2591,N_2637);
nand U3011 (N_3011,N_2900,N_2702);
nor U3012 (N_3012,N_2746,N_2613);
or U3013 (N_3013,N_2729,N_2656);
nand U3014 (N_3014,N_2978,N_2525);
nor U3015 (N_3015,N_2897,N_2832);
or U3016 (N_3016,N_2651,N_2849);
or U3017 (N_3017,N_2536,N_2636);
or U3018 (N_3018,N_2534,N_2590);
and U3019 (N_3019,N_2907,N_2606);
or U3020 (N_3020,N_2530,N_2587);
nor U3021 (N_3021,N_2894,N_2962);
or U3022 (N_3022,N_2548,N_2629);
and U3023 (N_3023,N_2604,N_2565);
and U3024 (N_3024,N_2779,N_2804);
or U3025 (N_3025,N_2516,N_2823);
xnor U3026 (N_3026,N_2595,N_2572);
and U3027 (N_3027,N_2691,N_2995);
nand U3028 (N_3028,N_2982,N_2500);
nand U3029 (N_3029,N_2951,N_2916);
or U3030 (N_3030,N_2910,N_2598);
nand U3031 (N_3031,N_2670,N_2762);
and U3032 (N_3032,N_2830,N_2844);
nand U3033 (N_3033,N_2686,N_2553);
nand U3034 (N_3034,N_2522,N_2557);
nor U3035 (N_3035,N_2754,N_2837);
xnor U3036 (N_3036,N_2724,N_2612);
or U3037 (N_3037,N_2772,N_2507);
and U3038 (N_3038,N_2955,N_2582);
nand U3039 (N_3039,N_2883,N_2794);
or U3040 (N_3040,N_2610,N_2699);
xor U3041 (N_3041,N_2682,N_2786);
nand U3042 (N_3042,N_2558,N_2842);
or U3043 (N_3043,N_2734,N_2966);
or U3044 (N_3044,N_2945,N_2929);
nor U3045 (N_3045,N_2722,N_2881);
nand U3046 (N_3046,N_2647,N_2969);
nand U3047 (N_3047,N_2993,N_2589);
and U3048 (N_3048,N_2757,N_2942);
nand U3049 (N_3049,N_2512,N_2954);
nor U3050 (N_3050,N_2728,N_2861);
nor U3051 (N_3051,N_2719,N_2800);
or U3052 (N_3052,N_2799,N_2669);
and U3053 (N_3053,N_2733,N_2555);
nor U3054 (N_3054,N_2609,N_2763);
or U3055 (N_3055,N_2840,N_2615);
nand U3056 (N_3056,N_2930,N_2860);
or U3057 (N_3057,N_2887,N_2931);
or U3058 (N_3058,N_2927,N_2863);
nor U3059 (N_3059,N_2759,N_2964);
nand U3060 (N_3060,N_2513,N_2544);
xnor U3061 (N_3061,N_2625,N_2663);
and U3062 (N_3062,N_2868,N_2811);
or U3063 (N_3063,N_2934,N_2908);
and U3064 (N_3064,N_2571,N_2685);
nor U3065 (N_3065,N_2603,N_2827);
and U3066 (N_3066,N_2627,N_2986);
nor U3067 (N_3067,N_2858,N_2828);
and U3068 (N_3068,N_2760,N_2698);
nor U3069 (N_3069,N_2706,N_2867);
nand U3070 (N_3070,N_2701,N_2696);
nor U3071 (N_3071,N_2501,N_2781);
or U3072 (N_3072,N_2869,N_2877);
and U3073 (N_3073,N_2674,N_2839);
or U3074 (N_3074,N_2574,N_2987);
nand U3075 (N_3075,N_2528,N_2535);
or U3076 (N_3076,N_2968,N_2853);
nand U3077 (N_3077,N_2825,N_2752);
and U3078 (N_3078,N_2977,N_2704);
and U3079 (N_3079,N_2758,N_2561);
or U3080 (N_3080,N_2905,N_2679);
nand U3081 (N_3081,N_2753,N_2694);
nand U3082 (N_3082,N_2914,N_2783);
nand U3083 (N_3083,N_2646,N_2997);
nor U3084 (N_3084,N_2873,N_2999);
and U3085 (N_3085,N_2747,N_2742);
nor U3086 (N_3086,N_2745,N_2741);
or U3087 (N_3087,N_2884,N_2521);
nand U3088 (N_3088,N_2956,N_2639);
nor U3089 (N_3089,N_2857,N_2633);
or U3090 (N_3090,N_2761,N_2855);
or U3091 (N_3091,N_2768,N_2851);
or U3092 (N_3092,N_2922,N_2791);
and U3093 (N_3093,N_2725,N_2766);
xor U3094 (N_3094,N_2985,N_2764);
nand U3095 (N_3095,N_2915,N_2551);
or U3096 (N_3096,N_2688,N_2990);
or U3097 (N_3097,N_2806,N_2892);
nand U3098 (N_3098,N_2787,N_2539);
and U3099 (N_3099,N_2785,N_2810);
or U3100 (N_3100,N_2972,N_2562);
and U3101 (N_3101,N_2805,N_2520);
nand U3102 (N_3102,N_2975,N_2709);
nor U3103 (N_3103,N_2852,N_2579);
or U3104 (N_3104,N_2967,N_2650);
and U3105 (N_3105,N_2959,N_2991);
nor U3106 (N_3106,N_2838,N_2826);
or U3107 (N_3107,N_2971,N_2621);
nor U3108 (N_3108,N_2952,N_2664);
xor U3109 (N_3109,N_2584,N_2617);
nor U3110 (N_3110,N_2820,N_2640);
or U3111 (N_3111,N_2891,N_2649);
nor U3112 (N_3112,N_2503,N_2726);
or U3113 (N_3113,N_2872,N_2953);
or U3114 (N_3114,N_2710,N_2665);
nand U3115 (N_3115,N_2963,N_2751);
nand U3116 (N_3116,N_2578,N_2831);
nand U3117 (N_3117,N_2773,N_2835);
nor U3118 (N_3118,N_2659,N_2635);
or U3119 (N_3119,N_2517,N_2943);
nor U3120 (N_3120,N_2708,N_2671);
and U3121 (N_3121,N_2755,N_2575);
nand U3122 (N_3122,N_2816,N_2846);
or U3123 (N_3123,N_2703,N_2833);
or U3124 (N_3124,N_2996,N_2850);
nor U3125 (N_3125,N_2560,N_2654);
nor U3126 (N_3126,N_2784,N_2712);
nand U3127 (N_3127,N_2677,N_2876);
or U3128 (N_3128,N_2903,N_2540);
nand U3129 (N_3129,N_2721,N_2845);
or U3130 (N_3130,N_2871,N_2814);
nor U3131 (N_3131,N_2879,N_2796);
nand U3132 (N_3132,N_2693,N_2949);
or U3133 (N_3133,N_2821,N_2776);
or U3134 (N_3134,N_2899,N_2643);
nor U3135 (N_3135,N_2933,N_2918);
and U3136 (N_3136,N_2994,N_2607);
nor U3137 (N_3137,N_2652,N_2778);
nor U3138 (N_3138,N_2818,N_2813);
or U3139 (N_3139,N_2655,N_2765);
nor U3140 (N_3140,N_2683,N_2672);
nor U3141 (N_3141,N_2614,N_2642);
or U3142 (N_3142,N_2676,N_2716);
nand U3143 (N_3143,N_2896,N_2526);
and U3144 (N_3144,N_2581,N_2774);
or U3145 (N_3145,N_2928,N_2543);
nor U3146 (N_3146,N_2577,N_2920);
nand U3147 (N_3147,N_2717,N_2793);
nand U3148 (N_3148,N_2932,N_2886);
nand U3149 (N_3149,N_2675,N_2618);
nor U3150 (N_3150,N_2554,N_2885);
and U3151 (N_3151,N_2748,N_2586);
or U3152 (N_3152,N_2707,N_2912);
nor U3153 (N_3153,N_2983,N_2518);
nand U3154 (N_3154,N_2780,N_2505);
nor U3155 (N_3155,N_2737,N_2510);
nand U3156 (N_3156,N_2600,N_2653);
and U3157 (N_3157,N_2735,N_2744);
nand U3158 (N_3158,N_2605,N_2570);
or U3159 (N_3159,N_2718,N_2750);
and U3160 (N_3160,N_2944,N_2988);
and U3161 (N_3161,N_2583,N_2859);
or U3162 (N_3162,N_2529,N_2819);
and U3163 (N_3163,N_2950,N_2713);
or U3164 (N_3164,N_2608,N_2559);
and U3165 (N_3165,N_2809,N_2504);
nor U3166 (N_3166,N_2947,N_2749);
or U3167 (N_3167,N_2801,N_2878);
nand U3168 (N_3168,N_2756,N_2616);
nand U3169 (N_3169,N_2715,N_2611);
and U3170 (N_3170,N_2593,N_2568);
nor U3171 (N_3171,N_2657,N_2630);
or U3172 (N_3172,N_2736,N_2533);
nor U3173 (N_3173,N_2870,N_2817);
nor U3174 (N_3174,N_2824,N_2957);
or U3175 (N_3175,N_2939,N_2815);
nand U3176 (N_3176,N_2508,N_2680);
or U3177 (N_3177,N_2898,N_2502);
nor U3178 (N_3178,N_2538,N_2547);
or U3179 (N_3179,N_2906,N_2509);
or U3180 (N_3180,N_2601,N_2666);
nor U3181 (N_3181,N_2732,N_2874);
nor U3182 (N_3182,N_2537,N_2727);
nand U3183 (N_3183,N_2668,N_2848);
nor U3184 (N_3184,N_2919,N_2979);
or U3185 (N_3185,N_2714,N_2658);
or U3186 (N_3186,N_2673,N_2803);
nor U3187 (N_3187,N_2523,N_2960);
and U3188 (N_3188,N_2739,N_2782);
nor U3189 (N_3189,N_2913,N_2738);
and U3190 (N_3190,N_2802,N_2948);
and U3191 (N_3191,N_2597,N_2767);
and U3192 (N_3192,N_2678,N_2632);
or U3193 (N_3193,N_2836,N_2909);
nor U3194 (N_3194,N_2695,N_2974);
or U3195 (N_3195,N_2847,N_2888);
and U3196 (N_3196,N_2923,N_2506);
or U3197 (N_3197,N_2973,N_2958);
nand U3198 (N_3198,N_2865,N_2550);
nand U3199 (N_3199,N_2532,N_2921);
nand U3200 (N_3200,N_2638,N_2684);
or U3201 (N_3201,N_2542,N_2989);
and U3202 (N_3202,N_2841,N_2961);
nand U3203 (N_3203,N_2941,N_2743);
and U3204 (N_3204,N_2875,N_2822);
nand U3205 (N_3205,N_2620,N_2984);
and U3206 (N_3206,N_2730,N_2864);
nor U3207 (N_3207,N_2622,N_2541);
and U3208 (N_3208,N_2917,N_2992);
nand U3209 (N_3209,N_2569,N_2940);
and U3210 (N_3210,N_2527,N_2619);
or U3211 (N_3211,N_2834,N_2723);
or U3212 (N_3212,N_2946,N_2777);
nand U3213 (N_3213,N_2662,N_2515);
and U3214 (N_3214,N_2660,N_2893);
nor U3215 (N_3215,N_2790,N_2624);
nand U3216 (N_3216,N_2545,N_2687);
nand U3217 (N_3217,N_2926,N_2829);
nor U3218 (N_3218,N_2970,N_2644);
nor U3219 (N_3219,N_2531,N_2519);
nor U3220 (N_3220,N_2566,N_2711);
nor U3221 (N_3221,N_2935,N_2588);
nand U3222 (N_3222,N_2690,N_2812);
nand U3223 (N_3223,N_2689,N_2882);
nor U3224 (N_3224,N_2731,N_2705);
nand U3225 (N_3225,N_2740,N_2936);
nand U3226 (N_3226,N_2895,N_2862);
xor U3227 (N_3227,N_2981,N_2880);
nand U3228 (N_3228,N_2770,N_2667);
nand U3229 (N_3229,N_2634,N_2980);
and U3230 (N_3230,N_2697,N_2808);
or U3231 (N_3231,N_2775,N_2924);
or U3232 (N_3232,N_2890,N_2645);
nor U3233 (N_3233,N_2789,N_2552);
nand U3234 (N_3234,N_2511,N_2631);
nor U3235 (N_3235,N_2792,N_2889);
and U3236 (N_3236,N_2564,N_2692);
nor U3237 (N_3237,N_2549,N_2594);
and U3238 (N_3238,N_2648,N_2854);
xnor U3239 (N_3239,N_2769,N_2788);
and U3240 (N_3240,N_2911,N_2576);
nor U3241 (N_3241,N_2592,N_2514);
nor U3242 (N_3242,N_2902,N_2628);
nor U3243 (N_3243,N_2904,N_2641);
or U3244 (N_3244,N_2556,N_2720);
or U3245 (N_3245,N_2866,N_2771);
nor U3246 (N_3246,N_2596,N_2843);
nor U3247 (N_3247,N_2856,N_2998);
and U3248 (N_3248,N_2626,N_2937);
or U3249 (N_3249,N_2661,N_2976);
xnor U3250 (N_3250,N_2875,N_2739);
nand U3251 (N_3251,N_2882,N_2594);
and U3252 (N_3252,N_2948,N_2923);
and U3253 (N_3253,N_2823,N_2758);
or U3254 (N_3254,N_2935,N_2504);
and U3255 (N_3255,N_2650,N_2679);
nor U3256 (N_3256,N_2791,N_2976);
nor U3257 (N_3257,N_2869,N_2603);
and U3258 (N_3258,N_2938,N_2525);
and U3259 (N_3259,N_2863,N_2578);
nand U3260 (N_3260,N_2867,N_2896);
or U3261 (N_3261,N_2579,N_2638);
nor U3262 (N_3262,N_2863,N_2598);
and U3263 (N_3263,N_2833,N_2851);
and U3264 (N_3264,N_2929,N_2742);
and U3265 (N_3265,N_2575,N_2625);
and U3266 (N_3266,N_2899,N_2836);
and U3267 (N_3267,N_2825,N_2937);
nor U3268 (N_3268,N_2842,N_2877);
nand U3269 (N_3269,N_2913,N_2640);
xor U3270 (N_3270,N_2842,N_2561);
and U3271 (N_3271,N_2521,N_2518);
and U3272 (N_3272,N_2617,N_2764);
or U3273 (N_3273,N_2848,N_2513);
nor U3274 (N_3274,N_2957,N_2622);
or U3275 (N_3275,N_2878,N_2676);
or U3276 (N_3276,N_2829,N_2671);
and U3277 (N_3277,N_2825,N_2527);
and U3278 (N_3278,N_2888,N_2993);
or U3279 (N_3279,N_2960,N_2874);
nor U3280 (N_3280,N_2542,N_2720);
nor U3281 (N_3281,N_2888,N_2669);
nand U3282 (N_3282,N_2571,N_2915);
nand U3283 (N_3283,N_2799,N_2986);
nor U3284 (N_3284,N_2936,N_2723);
nand U3285 (N_3285,N_2917,N_2775);
nor U3286 (N_3286,N_2966,N_2769);
and U3287 (N_3287,N_2568,N_2692);
and U3288 (N_3288,N_2807,N_2856);
nand U3289 (N_3289,N_2649,N_2579);
and U3290 (N_3290,N_2825,N_2823);
or U3291 (N_3291,N_2718,N_2864);
and U3292 (N_3292,N_2981,N_2858);
nand U3293 (N_3293,N_2955,N_2993);
and U3294 (N_3294,N_2667,N_2913);
or U3295 (N_3295,N_2651,N_2505);
and U3296 (N_3296,N_2761,N_2909);
nor U3297 (N_3297,N_2798,N_2771);
nor U3298 (N_3298,N_2911,N_2885);
and U3299 (N_3299,N_2882,N_2796);
nor U3300 (N_3300,N_2526,N_2566);
nor U3301 (N_3301,N_2635,N_2559);
and U3302 (N_3302,N_2532,N_2760);
nor U3303 (N_3303,N_2595,N_2529);
nor U3304 (N_3304,N_2719,N_2785);
nor U3305 (N_3305,N_2816,N_2512);
and U3306 (N_3306,N_2770,N_2910);
and U3307 (N_3307,N_2754,N_2786);
xnor U3308 (N_3308,N_2690,N_2950);
and U3309 (N_3309,N_2826,N_2527);
nand U3310 (N_3310,N_2711,N_2987);
and U3311 (N_3311,N_2793,N_2823);
nor U3312 (N_3312,N_2922,N_2533);
xor U3313 (N_3313,N_2831,N_2615);
nor U3314 (N_3314,N_2673,N_2689);
nand U3315 (N_3315,N_2644,N_2811);
and U3316 (N_3316,N_2904,N_2501);
or U3317 (N_3317,N_2602,N_2583);
and U3318 (N_3318,N_2764,N_2726);
xor U3319 (N_3319,N_2637,N_2506);
xnor U3320 (N_3320,N_2554,N_2716);
nor U3321 (N_3321,N_2802,N_2525);
nand U3322 (N_3322,N_2533,N_2984);
or U3323 (N_3323,N_2715,N_2516);
nand U3324 (N_3324,N_2627,N_2567);
and U3325 (N_3325,N_2687,N_2947);
or U3326 (N_3326,N_2720,N_2990);
or U3327 (N_3327,N_2554,N_2522);
and U3328 (N_3328,N_2605,N_2886);
and U3329 (N_3329,N_2545,N_2581);
and U3330 (N_3330,N_2782,N_2797);
or U3331 (N_3331,N_2915,N_2794);
and U3332 (N_3332,N_2936,N_2501);
and U3333 (N_3333,N_2507,N_2854);
and U3334 (N_3334,N_2897,N_2544);
or U3335 (N_3335,N_2763,N_2695);
nor U3336 (N_3336,N_2743,N_2536);
and U3337 (N_3337,N_2576,N_2775);
nor U3338 (N_3338,N_2627,N_2892);
nor U3339 (N_3339,N_2819,N_2736);
or U3340 (N_3340,N_2774,N_2932);
nor U3341 (N_3341,N_2912,N_2745);
nand U3342 (N_3342,N_2626,N_2612);
nand U3343 (N_3343,N_2579,N_2964);
and U3344 (N_3344,N_2682,N_2561);
and U3345 (N_3345,N_2923,N_2843);
nand U3346 (N_3346,N_2791,N_2544);
nor U3347 (N_3347,N_2517,N_2808);
and U3348 (N_3348,N_2970,N_2705);
or U3349 (N_3349,N_2520,N_2675);
nor U3350 (N_3350,N_2704,N_2577);
nor U3351 (N_3351,N_2783,N_2811);
nand U3352 (N_3352,N_2531,N_2976);
or U3353 (N_3353,N_2742,N_2611);
and U3354 (N_3354,N_2926,N_2831);
nor U3355 (N_3355,N_2641,N_2859);
or U3356 (N_3356,N_2936,N_2697);
nand U3357 (N_3357,N_2506,N_2522);
nor U3358 (N_3358,N_2643,N_2969);
nand U3359 (N_3359,N_2720,N_2535);
or U3360 (N_3360,N_2883,N_2930);
nand U3361 (N_3361,N_2951,N_2704);
nor U3362 (N_3362,N_2528,N_2663);
nand U3363 (N_3363,N_2542,N_2792);
and U3364 (N_3364,N_2797,N_2881);
and U3365 (N_3365,N_2706,N_2519);
and U3366 (N_3366,N_2918,N_2828);
nor U3367 (N_3367,N_2750,N_2555);
or U3368 (N_3368,N_2794,N_2613);
nand U3369 (N_3369,N_2736,N_2512);
nor U3370 (N_3370,N_2865,N_2819);
nor U3371 (N_3371,N_2963,N_2569);
or U3372 (N_3372,N_2513,N_2588);
and U3373 (N_3373,N_2794,N_2769);
or U3374 (N_3374,N_2679,N_2984);
nor U3375 (N_3375,N_2507,N_2769);
or U3376 (N_3376,N_2885,N_2558);
or U3377 (N_3377,N_2586,N_2876);
or U3378 (N_3378,N_2598,N_2645);
nor U3379 (N_3379,N_2911,N_2739);
and U3380 (N_3380,N_2826,N_2608);
and U3381 (N_3381,N_2889,N_2562);
nand U3382 (N_3382,N_2604,N_2760);
nor U3383 (N_3383,N_2732,N_2905);
and U3384 (N_3384,N_2974,N_2698);
or U3385 (N_3385,N_2954,N_2708);
nand U3386 (N_3386,N_2524,N_2976);
nor U3387 (N_3387,N_2705,N_2667);
nor U3388 (N_3388,N_2806,N_2953);
nand U3389 (N_3389,N_2924,N_2965);
or U3390 (N_3390,N_2704,N_2583);
xnor U3391 (N_3391,N_2542,N_2925);
nand U3392 (N_3392,N_2595,N_2979);
nand U3393 (N_3393,N_2569,N_2557);
nor U3394 (N_3394,N_2609,N_2627);
and U3395 (N_3395,N_2760,N_2745);
and U3396 (N_3396,N_2774,N_2570);
or U3397 (N_3397,N_2965,N_2960);
or U3398 (N_3398,N_2829,N_2963);
and U3399 (N_3399,N_2893,N_2997);
or U3400 (N_3400,N_2985,N_2577);
or U3401 (N_3401,N_2934,N_2594);
nor U3402 (N_3402,N_2893,N_2521);
nand U3403 (N_3403,N_2843,N_2837);
and U3404 (N_3404,N_2614,N_2704);
or U3405 (N_3405,N_2780,N_2874);
nand U3406 (N_3406,N_2945,N_2535);
nor U3407 (N_3407,N_2852,N_2867);
nor U3408 (N_3408,N_2505,N_2885);
and U3409 (N_3409,N_2959,N_2886);
nor U3410 (N_3410,N_2700,N_2810);
and U3411 (N_3411,N_2830,N_2942);
nand U3412 (N_3412,N_2719,N_2696);
nand U3413 (N_3413,N_2695,N_2648);
and U3414 (N_3414,N_2547,N_2796);
and U3415 (N_3415,N_2511,N_2555);
xor U3416 (N_3416,N_2550,N_2517);
and U3417 (N_3417,N_2918,N_2710);
nand U3418 (N_3418,N_2878,N_2713);
or U3419 (N_3419,N_2578,N_2891);
and U3420 (N_3420,N_2710,N_2608);
nand U3421 (N_3421,N_2538,N_2910);
and U3422 (N_3422,N_2839,N_2654);
or U3423 (N_3423,N_2972,N_2849);
and U3424 (N_3424,N_2807,N_2545);
nand U3425 (N_3425,N_2802,N_2996);
nand U3426 (N_3426,N_2564,N_2972);
or U3427 (N_3427,N_2626,N_2586);
nand U3428 (N_3428,N_2884,N_2876);
or U3429 (N_3429,N_2530,N_2863);
nor U3430 (N_3430,N_2684,N_2788);
nand U3431 (N_3431,N_2675,N_2534);
or U3432 (N_3432,N_2810,N_2935);
or U3433 (N_3433,N_2622,N_2559);
xor U3434 (N_3434,N_2805,N_2502);
nand U3435 (N_3435,N_2967,N_2617);
nor U3436 (N_3436,N_2586,N_2607);
or U3437 (N_3437,N_2932,N_2501);
and U3438 (N_3438,N_2758,N_2570);
and U3439 (N_3439,N_2959,N_2688);
and U3440 (N_3440,N_2650,N_2806);
nor U3441 (N_3441,N_2628,N_2687);
or U3442 (N_3442,N_2993,N_2717);
and U3443 (N_3443,N_2810,N_2679);
nand U3444 (N_3444,N_2721,N_2631);
nand U3445 (N_3445,N_2598,N_2932);
nand U3446 (N_3446,N_2647,N_2730);
and U3447 (N_3447,N_2715,N_2923);
nand U3448 (N_3448,N_2711,N_2937);
nor U3449 (N_3449,N_2758,N_2765);
and U3450 (N_3450,N_2683,N_2542);
and U3451 (N_3451,N_2781,N_2736);
nor U3452 (N_3452,N_2870,N_2785);
nand U3453 (N_3453,N_2656,N_2889);
xor U3454 (N_3454,N_2943,N_2555);
nor U3455 (N_3455,N_2948,N_2857);
nand U3456 (N_3456,N_2611,N_2526);
and U3457 (N_3457,N_2788,N_2752);
nand U3458 (N_3458,N_2950,N_2706);
nand U3459 (N_3459,N_2519,N_2775);
and U3460 (N_3460,N_2609,N_2680);
nor U3461 (N_3461,N_2729,N_2797);
or U3462 (N_3462,N_2788,N_2657);
nor U3463 (N_3463,N_2935,N_2743);
and U3464 (N_3464,N_2745,N_2979);
nor U3465 (N_3465,N_2827,N_2777);
nor U3466 (N_3466,N_2604,N_2746);
nand U3467 (N_3467,N_2738,N_2956);
or U3468 (N_3468,N_2575,N_2548);
or U3469 (N_3469,N_2813,N_2774);
and U3470 (N_3470,N_2783,N_2848);
nand U3471 (N_3471,N_2559,N_2612);
nor U3472 (N_3472,N_2753,N_2674);
nand U3473 (N_3473,N_2877,N_2556);
and U3474 (N_3474,N_2593,N_2564);
and U3475 (N_3475,N_2683,N_2878);
or U3476 (N_3476,N_2570,N_2880);
nor U3477 (N_3477,N_2704,N_2716);
or U3478 (N_3478,N_2705,N_2538);
and U3479 (N_3479,N_2875,N_2673);
nand U3480 (N_3480,N_2754,N_2828);
nor U3481 (N_3481,N_2881,N_2737);
nand U3482 (N_3482,N_2975,N_2745);
nor U3483 (N_3483,N_2847,N_2921);
nand U3484 (N_3484,N_2591,N_2789);
and U3485 (N_3485,N_2957,N_2547);
and U3486 (N_3486,N_2557,N_2521);
nand U3487 (N_3487,N_2544,N_2644);
xor U3488 (N_3488,N_2582,N_2781);
nor U3489 (N_3489,N_2849,N_2532);
or U3490 (N_3490,N_2602,N_2568);
nor U3491 (N_3491,N_2669,N_2638);
or U3492 (N_3492,N_2867,N_2647);
and U3493 (N_3493,N_2777,N_2759);
nand U3494 (N_3494,N_2676,N_2909);
nand U3495 (N_3495,N_2872,N_2572);
and U3496 (N_3496,N_2934,N_2720);
nor U3497 (N_3497,N_2621,N_2827);
or U3498 (N_3498,N_2704,N_2512);
nor U3499 (N_3499,N_2944,N_2795);
nor U3500 (N_3500,N_3453,N_3000);
and U3501 (N_3501,N_3450,N_3314);
nor U3502 (N_3502,N_3180,N_3308);
and U3503 (N_3503,N_3352,N_3261);
or U3504 (N_3504,N_3232,N_3489);
xnor U3505 (N_3505,N_3239,N_3138);
and U3506 (N_3506,N_3130,N_3062);
nor U3507 (N_3507,N_3167,N_3371);
or U3508 (N_3508,N_3250,N_3418);
or U3509 (N_3509,N_3330,N_3347);
or U3510 (N_3510,N_3054,N_3491);
nand U3511 (N_3511,N_3119,N_3118);
or U3512 (N_3512,N_3409,N_3073);
or U3513 (N_3513,N_3391,N_3066);
nor U3514 (N_3514,N_3077,N_3013);
or U3515 (N_3515,N_3154,N_3052);
nand U3516 (N_3516,N_3302,N_3482);
or U3517 (N_3517,N_3034,N_3063);
nor U3518 (N_3518,N_3114,N_3241);
and U3519 (N_3519,N_3475,N_3245);
and U3520 (N_3520,N_3351,N_3224);
and U3521 (N_3521,N_3354,N_3488);
xor U3522 (N_3522,N_3203,N_3191);
nand U3523 (N_3523,N_3202,N_3199);
or U3524 (N_3524,N_3356,N_3289);
and U3525 (N_3525,N_3246,N_3259);
nor U3526 (N_3526,N_3369,N_3374);
nor U3527 (N_3527,N_3218,N_3258);
and U3528 (N_3528,N_3108,N_3099);
and U3529 (N_3529,N_3042,N_3019);
xor U3530 (N_3530,N_3255,N_3431);
and U3531 (N_3531,N_3050,N_3048);
nand U3532 (N_3532,N_3164,N_3333);
nand U3533 (N_3533,N_3288,N_3003);
nor U3534 (N_3534,N_3210,N_3481);
and U3535 (N_3535,N_3280,N_3225);
or U3536 (N_3536,N_3343,N_3028);
and U3537 (N_3537,N_3070,N_3329);
nand U3538 (N_3538,N_3186,N_3367);
xnor U3539 (N_3539,N_3417,N_3365);
xnor U3540 (N_3540,N_3275,N_3057);
or U3541 (N_3541,N_3058,N_3012);
or U3542 (N_3542,N_3004,N_3484);
or U3543 (N_3543,N_3323,N_3140);
or U3544 (N_3544,N_3483,N_3421);
nand U3545 (N_3545,N_3122,N_3290);
nor U3546 (N_3546,N_3087,N_3277);
nand U3547 (N_3547,N_3105,N_3136);
and U3548 (N_3548,N_3016,N_3318);
nor U3549 (N_3549,N_3242,N_3303);
nand U3550 (N_3550,N_3056,N_3157);
or U3551 (N_3551,N_3260,N_3079);
nand U3552 (N_3552,N_3166,N_3233);
and U3553 (N_3553,N_3357,N_3030);
or U3554 (N_3554,N_3486,N_3425);
nand U3555 (N_3555,N_3040,N_3315);
and U3556 (N_3556,N_3036,N_3468);
nor U3557 (N_3557,N_3492,N_3403);
and U3558 (N_3558,N_3388,N_3123);
nor U3559 (N_3559,N_3359,N_3041);
nand U3560 (N_3560,N_3211,N_3452);
nor U3561 (N_3561,N_3080,N_3176);
nor U3562 (N_3562,N_3436,N_3462);
nor U3563 (N_3563,N_3212,N_3276);
and U3564 (N_3564,N_3010,N_3293);
xnor U3565 (N_3565,N_3069,N_3497);
and U3566 (N_3566,N_3410,N_3082);
nand U3567 (N_3567,N_3131,N_3072);
and U3568 (N_3568,N_3381,N_3071);
nand U3569 (N_3569,N_3256,N_3362);
and U3570 (N_3570,N_3132,N_3350);
and U3571 (N_3571,N_3023,N_3021);
and U3572 (N_3572,N_3401,N_3150);
nor U3573 (N_3573,N_3284,N_3393);
and U3574 (N_3574,N_3294,N_3395);
or U3575 (N_3575,N_3148,N_3430);
or U3576 (N_3576,N_3449,N_3229);
or U3577 (N_3577,N_3173,N_3024);
nor U3578 (N_3578,N_3018,N_3113);
nor U3579 (N_3579,N_3339,N_3262);
nand U3580 (N_3580,N_3363,N_3477);
nor U3581 (N_3581,N_3380,N_3423);
or U3582 (N_3582,N_3399,N_3473);
nand U3583 (N_3583,N_3149,N_3091);
nor U3584 (N_3584,N_3001,N_3181);
or U3585 (N_3585,N_3093,N_3207);
or U3586 (N_3586,N_3220,N_3402);
or U3587 (N_3587,N_3499,N_3404);
nor U3588 (N_3588,N_3397,N_3447);
nand U3589 (N_3589,N_3124,N_3291);
nand U3590 (N_3590,N_3109,N_3204);
or U3591 (N_3591,N_3265,N_3226);
nand U3592 (N_3592,N_3494,N_3183);
nor U3593 (N_3593,N_3243,N_3394);
or U3594 (N_3594,N_3353,N_3234);
nor U3595 (N_3595,N_3031,N_3435);
xnor U3596 (N_3596,N_3337,N_3014);
or U3597 (N_3597,N_3460,N_3219);
or U3598 (N_3598,N_3084,N_3295);
nand U3599 (N_3599,N_3469,N_3439);
or U3600 (N_3600,N_3228,N_3400);
or U3601 (N_3601,N_3476,N_3117);
and U3602 (N_3602,N_3376,N_3467);
and U3603 (N_3603,N_3116,N_3047);
or U3604 (N_3604,N_3478,N_3163);
and U3605 (N_3605,N_3089,N_3060);
and U3606 (N_3606,N_3195,N_3414);
nand U3607 (N_3607,N_3485,N_3463);
or U3608 (N_3608,N_3279,N_3107);
nand U3609 (N_3609,N_3461,N_3222);
nand U3610 (N_3610,N_3009,N_3364);
nor U3611 (N_3611,N_3197,N_3474);
and U3612 (N_3612,N_3493,N_3083);
or U3613 (N_3613,N_3322,N_3392);
or U3614 (N_3614,N_3102,N_3067);
nand U3615 (N_3615,N_3466,N_3035);
nor U3616 (N_3616,N_3086,N_3251);
or U3617 (N_3617,N_3214,N_3368);
nor U3618 (N_3618,N_3269,N_3139);
or U3619 (N_3619,N_3287,N_3045);
nor U3620 (N_3620,N_3487,N_3270);
nand U3621 (N_3621,N_3305,N_3076);
nand U3622 (N_3622,N_3465,N_3193);
and U3623 (N_3623,N_3049,N_3470);
or U3624 (N_3624,N_3115,N_3420);
nand U3625 (N_3625,N_3053,N_3064);
xnor U3626 (N_3626,N_3344,N_3104);
nand U3627 (N_3627,N_3128,N_3372);
nor U3628 (N_3628,N_3263,N_3398);
nor U3629 (N_3629,N_3142,N_3428);
nor U3630 (N_3630,N_3254,N_3038);
and U3631 (N_3631,N_3111,N_3006);
nor U3632 (N_3632,N_3094,N_3169);
xor U3633 (N_3633,N_3433,N_3160);
nand U3634 (N_3634,N_3216,N_3230);
or U3635 (N_3635,N_3286,N_3017);
and U3636 (N_3636,N_3144,N_3424);
and U3637 (N_3637,N_3349,N_3360);
and U3638 (N_3638,N_3422,N_3039);
nand U3639 (N_3639,N_3451,N_3158);
and U3640 (N_3640,N_3283,N_3358);
and U3641 (N_3641,N_3074,N_3426);
nor U3642 (N_3642,N_3065,N_3168);
nand U3643 (N_3643,N_3238,N_3007);
nor U3644 (N_3644,N_3137,N_3441);
nand U3645 (N_3645,N_3405,N_3313);
and U3646 (N_3646,N_3008,N_3172);
or U3647 (N_3647,N_3248,N_3464);
nor U3648 (N_3648,N_3103,N_3092);
nor U3649 (N_3649,N_3015,N_3434);
nor U3650 (N_3650,N_3236,N_3215);
and U3651 (N_3651,N_3386,N_3445);
nand U3652 (N_3652,N_3240,N_3145);
or U3653 (N_3653,N_3299,N_3440);
nand U3654 (N_3654,N_3155,N_3088);
and U3655 (N_3655,N_3162,N_3264);
nand U3656 (N_3656,N_3190,N_3253);
nor U3657 (N_3657,N_3427,N_3033);
nor U3658 (N_3658,N_3237,N_3200);
and U3659 (N_3659,N_3348,N_3319);
and U3660 (N_3660,N_3159,N_3194);
nor U3661 (N_3661,N_3061,N_3443);
and U3662 (N_3662,N_3387,N_3090);
or U3663 (N_3663,N_3298,N_3498);
nand U3664 (N_3664,N_3312,N_3437);
nand U3665 (N_3665,N_3025,N_3459);
nor U3666 (N_3666,N_3338,N_3340);
or U3667 (N_3667,N_3198,N_3309);
nor U3668 (N_3668,N_3438,N_3457);
and U3669 (N_3669,N_3133,N_3336);
or U3670 (N_3670,N_3141,N_3022);
and U3671 (N_3671,N_3310,N_3205);
or U3672 (N_3672,N_3324,N_3184);
nand U3673 (N_3673,N_3170,N_3495);
and U3674 (N_3674,N_3328,N_3382);
nand U3675 (N_3675,N_3292,N_3271);
or U3676 (N_3676,N_3296,N_3419);
nor U3677 (N_3677,N_3413,N_3126);
nand U3678 (N_3678,N_3385,N_3370);
and U3679 (N_3679,N_3335,N_3235);
and U3680 (N_3680,N_3496,N_3005);
or U3681 (N_3681,N_3444,N_3188);
nand U3682 (N_3682,N_3112,N_3120);
nor U3683 (N_3683,N_3231,N_3266);
nor U3684 (N_3684,N_3311,N_3378);
nor U3685 (N_3685,N_3026,N_3429);
nor U3686 (N_3686,N_3454,N_3249);
nor U3687 (N_3687,N_3455,N_3096);
nand U3688 (N_3688,N_3177,N_3274);
or U3689 (N_3689,N_3044,N_3285);
nand U3690 (N_3690,N_3411,N_3156);
nand U3691 (N_3691,N_3146,N_3227);
nand U3692 (N_3692,N_3272,N_3206);
or U3693 (N_3693,N_3377,N_3020);
nand U3694 (N_3694,N_3075,N_3389);
or U3695 (N_3695,N_3189,N_3165);
nor U3696 (N_3696,N_3110,N_3152);
or U3697 (N_3697,N_3366,N_3257);
and U3698 (N_3698,N_3479,N_3331);
nand U3699 (N_3699,N_3175,N_3247);
nor U3700 (N_3700,N_3316,N_3059);
nor U3701 (N_3701,N_3375,N_3281);
or U3702 (N_3702,N_3032,N_3027);
nor U3703 (N_3703,N_3297,N_3178);
nand U3704 (N_3704,N_3406,N_3321);
or U3705 (N_3705,N_3196,N_3304);
nor U3706 (N_3706,N_3320,N_3171);
and U3707 (N_3707,N_3472,N_3081);
nor U3708 (N_3708,N_3408,N_3301);
and U3709 (N_3709,N_3244,N_3208);
or U3710 (N_3710,N_3213,N_3278);
nor U3711 (N_3711,N_3327,N_3384);
nor U3712 (N_3712,N_3147,N_3458);
nand U3713 (N_3713,N_3490,N_3273);
nand U3714 (N_3714,N_3416,N_3355);
and U3715 (N_3715,N_3325,N_3095);
or U3716 (N_3716,N_3448,N_3043);
or U3717 (N_3717,N_3383,N_3101);
or U3718 (N_3718,N_3209,N_3252);
nor U3719 (N_3719,N_3129,N_3221);
and U3720 (N_3720,N_3051,N_3106);
nand U3721 (N_3721,N_3471,N_3097);
and U3722 (N_3722,N_3127,N_3134);
or U3723 (N_3723,N_3151,N_3268);
nand U3724 (N_3724,N_3346,N_3179);
or U3725 (N_3725,N_3161,N_3011);
and U3726 (N_3726,N_3185,N_3412);
or U3727 (N_3727,N_3379,N_3002);
nand U3728 (N_3728,N_3282,N_3037);
nand U3729 (N_3729,N_3174,N_3201);
and U3730 (N_3730,N_3143,N_3446);
or U3731 (N_3731,N_3456,N_3342);
nor U3732 (N_3732,N_3480,N_3415);
or U3733 (N_3733,N_3334,N_3345);
nand U3734 (N_3734,N_3267,N_3341);
or U3735 (N_3735,N_3100,N_3326);
nor U3736 (N_3736,N_3187,N_3317);
and U3737 (N_3737,N_3361,N_3192);
or U3738 (N_3738,N_3182,N_3332);
or U3739 (N_3739,N_3300,N_3085);
and U3740 (N_3740,N_3135,N_3121);
nand U3741 (N_3741,N_3432,N_3125);
and U3742 (N_3742,N_3153,N_3098);
xor U3743 (N_3743,N_3055,N_3029);
nand U3744 (N_3744,N_3217,N_3407);
nor U3745 (N_3745,N_3442,N_3223);
nor U3746 (N_3746,N_3078,N_3373);
and U3747 (N_3747,N_3307,N_3396);
nor U3748 (N_3748,N_3390,N_3046);
or U3749 (N_3749,N_3068,N_3306);
xor U3750 (N_3750,N_3013,N_3156);
nand U3751 (N_3751,N_3480,N_3478);
xnor U3752 (N_3752,N_3431,N_3420);
nor U3753 (N_3753,N_3227,N_3467);
or U3754 (N_3754,N_3378,N_3288);
nand U3755 (N_3755,N_3097,N_3151);
or U3756 (N_3756,N_3245,N_3448);
or U3757 (N_3757,N_3277,N_3009);
nor U3758 (N_3758,N_3384,N_3166);
and U3759 (N_3759,N_3488,N_3055);
nor U3760 (N_3760,N_3191,N_3394);
nand U3761 (N_3761,N_3305,N_3404);
nand U3762 (N_3762,N_3136,N_3096);
and U3763 (N_3763,N_3122,N_3038);
nand U3764 (N_3764,N_3253,N_3473);
nand U3765 (N_3765,N_3426,N_3466);
or U3766 (N_3766,N_3020,N_3183);
and U3767 (N_3767,N_3424,N_3057);
nand U3768 (N_3768,N_3267,N_3092);
nor U3769 (N_3769,N_3330,N_3111);
nand U3770 (N_3770,N_3085,N_3301);
or U3771 (N_3771,N_3375,N_3442);
nand U3772 (N_3772,N_3000,N_3156);
nand U3773 (N_3773,N_3252,N_3038);
nor U3774 (N_3774,N_3084,N_3185);
and U3775 (N_3775,N_3347,N_3174);
and U3776 (N_3776,N_3279,N_3349);
and U3777 (N_3777,N_3416,N_3206);
and U3778 (N_3778,N_3172,N_3287);
nor U3779 (N_3779,N_3059,N_3493);
and U3780 (N_3780,N_3312,N_3257);
nand U3781 (N_3781,N_3102,N_3240);
or U3782 (N_3782,N_3043,N_3032);
or U3783 (N_3783,N_3480,N_3115);
nor U3784 (N_3784,N_3170,N_3221);
or U3785 (N_3785,N_3162,N_3048);
or U3786 (N_3786,N_3348,N_3018);
nor U3787 (N_3787,N_3406,N_3499);
or U3788 (N_3788,N_3133,N_3352);
nor U3789 (N_3789,N_3101,N_3477);
or U3790 (N_3790,N_3067,N_3320);
nand U3791 (N_3791,N_3245,N_3246);
and U3792 (N_3792,N_3341,N_3104);
and U3793 (N_3793,N_3041,N_3100);
and U3794 (N_3794,N_3075,N_3456);
and U3795 (N_3795,N_3449,N_3126);
or U3796 (N_3796,N_3440,N_3483);
nor U3797 (N_3797,N_3119,N_3442);
or U3798 (N_3798,N_3246,N_3180);
and U3799 (N_3799,N_3374,N_3386);
xor U3800 (N_3800,N_3330,N_3231);
nand U3801 (N_3801,N_3098,N_3289);
nor U3802 (N_3802,N_3101,N_3040);
nand U3803 (N_3803,N_3078,N_3424);
or U3804 (N_3804,N_3358,N_3401);
or U3805 (N_3805,N_3345,N_3488);
or U3806 (N_3806,N_3012,N_3242);
nor U3807 (N_3807,N_3498,N_3012);
or U3808 (N_3808,N_3314,N_3440);
nand U3809 (N_3809,N_3110,N_3485);
nand U3810 (N_3810,N_3401,N_3293);
nand U3811 (N_3811,N_3454,N_3233);
and U3812 (N_3812,N_3209,N_3297);
nand U3813 (N_3813,N_3447,N_3399);
nand U3814 (N_3814,N_3281,N_3399);
nor U3815 (N_3815,N_3465,N_3116);
or U3816 (N_3816,N_3349,N_3063);
or U3817 (N_3817,N_3046,N_3408);
nand U3818 (N_3818,N_3477,N_3299);
or U3819 (N_3819,N_3320,N_3235);
and U3820 (N_3820,N_3143,N_3496);
and U3821 (N_3821,N_3355,N_3158);
nand U3822 (N_3822,N_3124,N_3419);
nor U3823 (N_3823,N_3027,N_3497);
nand U3824 (N_3824,N_3447,N_3155);
or U3825 (N_3825,N_3075,N_3144);
or U3826 (N_3826,N_3287,N_3192);
and U3827 (N_3827,N_3317,N_3493);
or U3828 (N_3828,N_3460,N_3325);
and U3829 (N_3829,N_3399,N_3373);
or U3830 (N_3830,N_3205,N_3000);
or U3831 (N_3831,N_3156,N_3029);
and U3832 (N_3832,N_3377,N_3222);
and U3833 (N_3833,N_3310,N_3036);
and U3834 (N_3834,N_3295,N_3039);
or U3835 (N_3835,N_3287,N_3001);
or U3836 (N_3836,N_3229,N_3355);
nand U3837 (N_3837,N_3492,N_3328);
nor U3838 (N_3838,N_3315,N_3266);
and U3839 (N_3839,N_3112,N_3432);
nor U3840 (N_3840,N_3370,N_3078);
nor U3841 (N_3841,N_3049,N_3129);
and U3842 (N_3842,N_3192,N_3132);
or U3843 (N_3843,N_3234,N_3383);
nor U3844 (N_3844,N_3007,N_3225);
nor U3845 (N_3845,N_3419,N_3020);
nor U3846 (N_3846,N_3059,N_3093);
nand U3847 (N_3847,N_3097,N_3154);
nand U3848 (N_3848,N_3295,N_3323);
and U3849 (N_3849,N_3319,N_3373);
or U3850 (N_3850,N_3200,N_3229);
nand U3851 (N_3851,N_3038,N_3417);
and U3852 (N_3852,N_3056,N_3387);
nand U3853 (N_3853,N_3086,N_3474);
or U3854 (N_3854,N_3035,N_3420);
nand U3855 (N_3855,N_3089,N_3376);
and U3856 (N_3856,N_3109,N_3003);
or U3857 (N_3857,N_3288,N_3165);
and U3858 (N_3858,N_3353,N_3465);
xnor U3859 (N_3859,N_3196,N_3387);
and U3860 (N_3860,N_3160,N_3300);
nand U3861 (N_3861,N_3322,N_3203);
or U3862 (N_3862,N_3210,N_3374);
or U3863 (N_3863,N_3386,N_3140);
and U3864 (N_3864,N_3434,N_3480);
and U3865 (N_3865,N_3282,N_3117);
nor U3866 (N_3866,N_3109,N_3030);
nor U3867 (N_3867,N_3118,N_3322);
nand U3868 (N_3868,N_3186,N_3078);
and U3869 (N_3869,N_3406,N_3299);
nand U3870 (N_3870,N_3209,N_3405);
and U3871 (N_3871,N_3091,N_3294);
or U3872 (N_3872,N_3328,N_3224);
or U3873 (N_3873,N_3203,N_3296);
nand U3874 (N_3874,N_3170,N_3135);
or U3875 (N_3875,N_3261,N_3467);
nand U3876 (N_3876,N_3112,N_3206);
and U3877 (N_3877,N_3323,N_3101);
and U3878 (N_3878,N_3499,N_3056);
nor U3879 (N_3879,N_3408,N_3017);
nand U3880 (N_3880,N_3092,N_3358);
nand U3881 (N_3881,N_3143,N_3055);
nand U3882 (N_3882,N_3393,N_3394);
nor U3883 (N_3883,N_3276,N_3451);
and U3884 (N_3884,N_3430,N_3130);
or U3885 (N_3885,N_3002,N_3095);
nor U3886 (N_3886,N_3249,N_3326);
nand U3887 (N_3887,N_3447,N_3132);
nand U3888 (N_3888,N_3443,N_3112);
or U3889 (N_3889,N_3285,N_3371);
nor U3890 (N_3890,N_3016,N_3444);
nand U3891 (N_3891,N_3033,N_3102);
nor U3892 (N_3892,N_3028,N_3154);
nor U3893 (N_3893,N_3278,N_3073);
or U3894 (N_3894,N_3090,N_3159);
nand U3895 (N_3895,N_3289,N_3385);
and U3896 (N_3896,N_3347,N_3013);
and U3897 (N_3897,N_3498,N_3313);
nor U3898 (N_3898,N_3490,N_3102);
nor U3899 (N_3899,N_3353,N_3076);
or U3900 (N_3900,N_3255,N_3278);
nor U3901 (N_3901,N_3325,N_3026);
nand U3902 (N_3902,N_3425,N_3458);
and U3903 (N_3903,N_3354,N_3021);
nor U3904 (N_3904,N_3233,N_3156);
xor U3905 (N_3905,N_3063,N_3449);
nand U3906 (N_3906,N_3455,N_3258);
or U3907 (N_3907,N_3455,N_3395);
or U3908 (N_3908,N_3346,N_3021);
and U3909 (N_3909,N_3374,N_3444);
nor U3910 (N_3910,N_3196,N_3202);
or U3911 (N_3911,N_3072,N_3170);
nor U3912 (N_3912,N_3016,N_3472);
nor U3913 (N_3913,N_3054,N_3034);
or U3914 (N_3914,N_3158,N_3096);
xnor U3915 (N_3915,N_3344,N_3264);
or U3916 (N_3916,N_3168,N_3063);
nand U3917 (N_3917,N_3498,N_3233);
xor U3918 (N_3918,N_3335,N_3070);
and U3919 (N_3919,N_3376,N_3103);
and U3920 (N_3920,N_3354,N_3365);
or U3921 (N_3921,N_3297,N_3470);
and U3922 (N_3922,N_3268,N_3393);
xnor U3923 (N_3923,N_3214,N_3341);
and U3924 (N_3924,N_3437,N_3150);
and U3925 (N_3925,N_3453,N_3372);
nand U3926 (N_3926,N_3058,N_3233);
nor U3927 (N_3927,N_3434,N_3280);
and U3928 (N_3928,N_3048,N_3205);
nand U3929 (N_3929,N_3003,N_3020);
nand U3930 (N_3930,N_3050,N_3116);
or U3931 (N_3931,N_3159,N_3454);
nor U3932 (N_3932,N_3419,N_3456);
nand U3933 (N_3933,N_3227,N_3255);
nor U3934 (N_3934,N_3448,N_3042);
and U3935 (N_3935,N_3333,N_3074);
nor U3936 (N_3936,N_3368,N_3315);
and U3937 (N_3937,N_3400,N_3226);
xnor U3938 (N_3938,N_3068,N_3007);
nand U3939 (N_3939,N_3343,N_3339);
nand U3940 (N_3940,N_3163,N_3054);
nor U3941 (N_3941,N_3068,N_3028);
nand U3942 (N_3942,N_3349,N_3213);
and U3943 (N_3943,N_3001,N_3157);
xnor U3944 (N_3944,N_3032,N_3421);
and U3945 (N_3945,N_3275,N_3335);
nand U3946 (N_3946,N_3473,N_3392);
nand U3947 (N_3947,N_3259,N_3328);
nor U3948 (N_3948,N_3495,N_3359);
or U3949 (N_3949,N_3237,N_3045);
nand U3950 (N_3950,N_3003,N_3124);
nor U3951 (N_3951,N_3466,N_3011);
and U3952 (N_3952,N_3473,N_3039);
nand U3953 (N_3953,N_3064,N_3293);
nor U3954 (N_3954,N_3004,N_3257);
nand U3955 (N_3955,N_3386,N_3025);
and U3956 (N_3956,N_3170,N_3345);
or U3957 (N_3957,N_3234,N_3222);
nor U3958 (N_3958,N_3138,N_3291);
nand U3959 (N_3959,N_3411,N_3367);
and U3960 (N_3960,N_3318,N_3488);
and U3961 (N_3961,N_3215,N_3383);
or U3962 (N_3962,N_3092,N_3075);
nor U3963 (N_3963,N_3366,N_3454);
or U3964 (N_3964,N_3050,N_3468);
nand U3965 (N_3965,N_3045,N_3023);
nand U3966 (N_3966,N_3152,N_3494);
and U3967 (N_3967,N_3289,N_3019);
nand U3968 (N_3968,N_3403,N_3373);
and U3969 (N_3969,N_3324,N_3497);
or U3970 (N_3970,N_3321,N_3417);
nand U3971 (N_3971,N_3213,N_3214);
nor U3972 (N_3972,N_3157,N_3106);
nor U3973 (N_3973,N_3343,N_3197);
nand U3974 (N_3974,N_3214,N_3307);
or U3975 (N_3975,N_3140,N_3275);
and U3976 (N_3976,N_3108,N_3032);
and U3977 (N_3977,N_3212,N_3013);
nand U3978 (N_3978,N_3481,N_3454);
and U3979 (N_3979,N_3206,N_3470);
nand U3980 (N_3980,N_3275,N_3387);
or U3981 (N_3981,N_3073,N_3288);
and U3982 (N_3982,N_3014,N_3109);
nor U3983 (N_3983,N_3289,N_3357);
nand U3984 (N_3984,N_3204,N_3126);
nand U3985 (N_3985,N_3238,N_3028);
or U3986 (N_3986,N_3426,N_3063);
nand U3987 (N_3987,N_3195,N_3311);
or U3988 (N_3988,N_3156,N_3152);
nor U3989 (N_3989,N_3437,N_3300);
or U3990 (N_3990,N_3060,N_3163);
nand U3991 (N_3991,N_3423,N_3449);
nand U3992 (N_3992,N_3492,N_3055);
or U3993 (N_3993,N_3293,N_3004);
nand U3994 (N_3994,N_3108,N_3024);
or U3995 (N_3995,N_3280,N_3468);
nor U3996 (N_3996,N_3012,N_3211);
or U3997 (N_3997,N_3417,N_3359);
nand U3998 (N_3998,N_3323,N_3009);
and U3999 (N_3999,N_3285,N_3038);
and U4000 (N_4000,N_3698,N_3763);
and U4001 (N_4001,N_3993,N_3783);
nor U4002 (N_4002,N_3603,N_3710);
nand U4003 (N_4003,N_3694,N_3661);
xnor U4004 (N_4004,N_3626,N_3722);
or U4005 (N_4005,N_3600,N_3664);
nor U4006 (N_4006,N_3965,N_3587);
or U4007 (N_4007,N_3572,N_3941);
nand U4008 (N_4008,N_3937,N_3911);
nor U4009 (N_4009,N_3645,N_3834);
or U4010 (N_4010,N_3795,N_3823);
xor U4011 (N_4011,N_3501,N_3735);
nand U4012 (N_4012,N_3923,N_3711);
and U4013 (N_4013,N_3932,N_3584);
and U4014 (N_4014,N_3537,N_3881);
nor U4015 (N_4015,N_3832,N_3833);
or U4016 (N_4016,N_3810,N_3819);
and U4017 (N_4017,N_3678,N_3560);
and U4018 (N_4018,N_3847,N_3982);
nor U4019 (N_4019,N_3590,N_3774);
nand U4020 (N_4020,N_3944,N_3918);
nand U4021 (N_4021,N_3970,N_3680);
and U4022 (N_4022,N_3503,N_3598);
nor U4023 (N_4023,N_3573,N_3951);
and U4024 (N_4024,N_3529,N_3548);
nor U4025 (N_4025,N_3748,N_3829);
nor U4026 (N_4026,N_3504,N_3788);
nand U4027 (N_4027,N_3618,N_3994);
nor U4028 (N_4028,N_3513,N_3632);
nand U4029 (N_4029,N_3903,N_3695);
or U4030 (N_4030,N_3507,N_3963);
nand U4031 (N_4031,N_3797,N_3804);
or U4032 (N_4032,N_3512,N_3790);
nand U4033 (N_4033,N_3607,N_3506);
nor U4034 (N_4034,N_3716,N_3822);
or U4035 (N_4035,N_3886,N_3756);
nor U4036 (N_4036,N_3967,N_3692);
nor U4037 (N_4037,N_3655,N_3690);
nor U4038 (N_4038,N_3636,N_3974);
nor U4039 (N_4039,N_3842,N_3902);
or U4040 (N_4040,N_3627,N_3516);
or U4041 (N_4041,N_3522,N_3563);
or U4042 (N_4042,N_3650,N_3651);
or U4043 (N_4043,N_3514,N_3633);
nor U4044 (N_4044,N_3968,N_3852);
nor U4045 (N_4045,N_3759,N_3525);
or U4046 (N_4046,N_3624,N_3988);
nor U4047 (N_4047,N_3879,N_3827);
nand U4048 (N_4048,N_3990,N_3532);
nor U4049 (N_4049,N_3976,N_3900);
nor U4050 (N_4050,N_3828,N_3565);
and U4051 (N_4051,N_3766,N_3571);
and U4052 (N_4052,N_3742,N_3700);
xnor U4053 (N_4053,N_3943,N_3746);
nand U4054 (N_4054,N_3801,N_3882);
nor U4055 (N_4055,N_3793,N_3569);
nand U4056 (N_4056,N_3595,N_3971);
nand U4057 (N_4057,N_3676,N_3719);
and U4058 (N_4058,N_3704,N_3892);
nand U4059 (N_4059,N_3551,N_3949);
and U4060 (N_4060,N_3684,N_3800);
nand U4061 (N_4061,N_3727,N_3677);
or U4062 (N_4062,N_3637,N_3764);
nand U4063 (N_4063,N_3740,N_3837);
nand U4064 (N_4064,N_3649,N_3653);
and U4065 (N_4065,N_3835,N_3814);
or U4066 (N_4066,N_3596,N_3745);
nor U4067 (N_4067,N_3582,N_3889);
or U4068 (N_4068,N_3796,N_3752);
nor U4069 (N_4069,N_3640,N_3726);
and U4070 (N_4070,N_3929,N_3562);
nor U4071 (N_4071,N_3777,N_3838);
or U4072 (N_4072,N_3639,N_3533);
or U4073 (N_4073,N_3861,N_3577);
nand U4074 (N_4074,N_3508,N_3914);
nand U4075 (N_4075,N_3916,N_3671);
nor U4076 (N_4076,N_3854,N_3975);
or U4077 (N_4077,N_3701,N_3579);
or U4078 (N_4078,N_3773,N_3973);
nor U4079 (N_4079,N_3939,N_3599);
nand U4080 (N_4080,N_3753,N_3897);
and U4081 (N_4081,N_3857,N_3705);
and U4082 (N_4082,N_3674,N_3905);
or U4083 (N_4083,N_3871,N_3799);
xor U4084 (N_4084,N_3948,N_3950);
nor U4085 (N_4085,N_3643,N_3991);
nor U4086 (N_4086,N_3917,N_3920);
nor U4087 (N_4087,N_3789,N_3818);
nor U4088 (N_4088,N_3635,N_3581);
or U4089 (N_4089,N_3915,N_3933);
nand U4090 (N_4090,N_3623,N_3865);
or U4091 (N_4091,N_3846,N_3862);
or U4092 (N_4092,N_3901,N_3841);
nand U4093 (N_4093,N_3502,N_3784);
nor U4094 (N_4094,N_3583,N_3665);
or U4095 (N_4095,N_3500,N_3884);
nor U4096 (N_4096,N_3863,N_3729);
or U4097 (N_4097,N_3675,N_3536);
nand U4098 (N_4098,N_3644,N_3732);
or U4099 (N_4099,N_3872,N_3605);
nor U4100 (N_4100,N_3638,N_3686);
nand U4101 (N_4101,N_3749,N_3725);
nand U4102 (N_4102,N_3682,N_3670);
nor U4103 (N_4103,N_3817,N_3712);
nor U4104 (N_4104,N_3647,N_3989);
and U4105 (N_4105,N_3807,N_3592);
nor U4106 (N_4106,N_3996,N_3805);
xnor U4107 (N_4107,N_3798,N_3806);
nor U4108 (N_4108,N_3617,N_3770);
nor U4109 (N_4109,N_3935,N_3885);
nor U4110 (N_4110,N_3921,N_3693);
or U4111 (N_4111,N_3812,N_3646);
or U4112 (N_4112,N_3708,N_3913);
nand U4113 (N_4113,N_3791,N_3767);
nand U4114 (N_4114,N_3622,N_3946);
nor U4115 (N_4115,N_3961,N_3864);
or U4116 (N_4116,N_3611,N_3699);
nand U4117 (N_4117,N_3808,N_3588);
or U4118 (N_4118,N_3540,N_3658);
xnor U4119 (N_4119,N_3831,N_3820);
nor U4120 (N_4120,N_3840,N_3762);
and U4121 (N_4121,N_3553,N_3743);
nand U4122 (N_4122,N_3535,N_3574);
nor U4123 (N_4123,N_3960,N_3985);
nand U4124 (N_4124,N_3778,N_3613);
and U4125 (N_4125,N_3546,N_3952);
or U4126 (N_4126,N_3668,N_3578);
nor U4127 (N_4127,N_3663,N_3620);
xor U4128 (N_4128,N_3981,N_3737);
and U4129 (N_4129,N_3866,N_3642);
and U4130 (N_4130,N_3550,N_3860);
and U4131 (N_4131,N_3717,N_3616);
and U4132 (N_4132,N_3926,N_3830);
nand U4133 (N_4133,N_3803,N_3849);
and U4134 (N_4134,N_3757,N_3679);
nor U4135 (N_4135,N_3602,N_3531);
or U4136 (N_4136,N_3591,N_3549);
nor U4137 (N_4137,N_3634,N_3555);
nand U4138 (N_4138,N_3844,N_3656);
xnor U4139 (N_4139,N_3815,N_3904);
and U4140 (N_4140,N_3713,N_3768);
nand U4141 (N_4141,N_3765,N_3594);
and U4142 (N_4142,N_3936,N_3621);
and U4143 (N_4143,N_3754,N_3606);
or U4144 (N_4144,N_3721,N_3541);
or U4145 (N_4145,N_3615,N_3683);
or U4146 (N_4146,N_3983,N_3586);
or U4147 (N_4147,N_3940,N_3659);
nand U4148 (N_4148,N_3505,N_3760);
or U4149 (N_4149,N_3517,N_3666);
and U4150 (N_4150,N_3922,N_3601);
nor U4151 (N_4151,N_3986,N_3906);
nand U4152 (N_4152,N_3999,N_3691);
nand U4153 (N_4153,N_3891,N_3570);
nand U4154 (N_4154,N_3912,N_3672);
nor U4155 (N_4155,N_3836,N_3959);
xor U4156 (N_4156,N_3776,N_3568);
nor U4157 (N_4157,N_3519,N_3567);
nor U4158 (N_4158,N_3995,N_3703);
nor U4159 (N_4159,N_3938,N_3954);
or U4160 (N_4160,N_3856,N_3772);
nor U4161 (N_4161,N_3564,N_3794);
nand U4162 (N_4162,N_3998,N_3654);
nand U4163 (N_4163,N_3530,N_3972);
nand U4164 (N_4164,N_3543,N_3887);
or U4165 (N_4165,N_3545,N_3552);
or U4166 (N_4166,N_3736,N_3909);
nor U4167 (N_4167,N_3955,N_3977);
xnor U4168 (N_4168,N_3589,N_3660);
nand U4169 (N_4169,N_3715,N_3855);
and U4170 (N_4170,N_3580,N_3612);
nor U4171 (N_4171,N_3811,N_3610);
nand U4172 (N_4172,N_3707,N_3681);
nor U4173 (N_4173,N_3769,N_3738);
or U4174 (N_4174,N_3641,N_3597);
and U4175 (N_4175,N_3724,N_3958);
or U4176 (N_4176,N_3741,N_3511);
and U4177 (N_4177,N_3910,N_3758);
nand U4178 (N_4178,N_3877,N_3771);
nor U4179 (N_4179,N_3896,N_3739);
and U4180 (N_4180,N_3809,N_3867);
and U4181 (N_4181,N_3880,N_3928);
nand U4182 (N_4182,N_3945,N_3883);
nor U4183 (N_4183,N_3907,N_3625);
and U4184 (N_4184,N_3874,N_3931);
nand U4185 (N_4185,N_3728,N_3539);
or U4186 (N_4186,N_3509,N_3924);
or U4187 (N_4187,N_3575,N_3526);
or U4188 (N_4188,N_3825,N_3802);
and U4189 (N_4189,N_3775,N_3566);
nor U4190 (N_4190,N_3687,N_3824);
nand U4191 (N_4191,N_3697,N_3576);
nand U4192 (N_4192,N_3609,N_3873);
or U4193 (N_4193,N_3528,N_3869);
nor U4194 (N_4194,N_3843,N_3761);
and U4195 (N_4195,N_3969,N_3934);
nand U4196 (N_4196,N_3731,N_3542);
nand U4197 (N_4197,N_3559,N_3527);
or U4198 (N_4198,N_3888,N_3667);
nand U4199 (N_4199,N_3899,N_3628);
nor U4200 (N_4200,N_3723,N_3781);
and U4201 (N_4201,N_3979,N_3547);
xor U4202 (N_4202,N_3755,N_3538);
nor U4203 (N_4203,N_3751,N_3953);
nor U4204 (N_4204,N_3558,N_3750);
or U4205 (N_4205,N_3930,N_3858);
nand U4206 (N_4206,N_3962,N_3696);
nand U4207 (N_4207,N_3652,N_3908);
or U4208 (N_4208,N_3813,N_3980);
and U4209 (N_4209,N_3848,N_3689);
and U4210 (N_4210,N_3688,N_3821);
nor U4211 (N_4211,N_3518,N_3964);
or U4212 (N_4212,N_3785,N_3956);
nand U4213 (N_4213,N_3997,N_3925);
nand U4214 (N_4214,N_3875,N_3685);
nand U4215 (N_4215,N_3714,N_3747);
nand U4216 (N_4216,N_3604,N_3608);
and U4217 (N_4217,N_3890,N_3870);
nand U4218 (N_4218,N_3554,N_3515);
nand U4219 (N_4219,N_3557,N_3845);
nor U4220 (N_4220,N_3733,N_3816);
or U4221 (N_4221,N_3893,N_3523);
and U4222 (N_4222,N_3629,N_3706);
and U4223 (N_4223,N_3630,N_3556);
nor U4224 (N_4224,N_3648,N_3966);
or U4225 (N_4225,N_3619,N_3510);
and U4226 (N_4226,N_3520,N_3521);
and U4227 (N_4227,N_3792,N_3895);
and U4228 (N_4228,N_3851,N_3782);
and U4229 (N_4229,N_3947,N_3984);
nor U4230 (N_4230,N_3898,N_3957);
nor U4231 (N_4231,N_3850,N_3779);
nand U4232 (N_4232,N_3780,N_3561);
nand U4233 (N_4233,N_3744,N_3669);
or U4234 (N_4234,N_3786,N_3730);
nand U4235 (N_4235,N_3868,N_3987);
xnor U4236 (N_4236,N_3593,N_3534);
nand U4237 (N_4237,N_3942,N_3978);
and U4238 (N_4238,N_3734,N_3878);
and U4239 (N_4239,N_3919,N_3544);
or U4240 (N_4240,N_3876,N_3720);
nand U4241 (N_4241,N_3787,N_3894);
or U4242 (N_4242,N_3853,N_3826);
and U4243 (N_4243,N_3673,N_3992);
and U4244 (N_4244,N_3839,N_3631);
nor U4245 (N_4245,N_3718,N_3614);
nor U4246 (N_4246,N_3709,N_3702);
nor U4247 (N_4247,N_3662,N_3524);
nor U4248 (N_4248,N_3927,N_3585);
or U4249 (N_4249,N_3859,N_3657);
nand U4250 (N_4250,N_3600,N_3807);
and U4251 (N_4251,N_3580,N_3562);
or U4252 (N_4252,N_3941,N_3792);
or U4253 (N_4253,N_3948,N_3799);
or U4254 (N_4254,N_3573,N_3581);
nand U4255 (N_4255,N_3923,N_3821);
nand U4256 (N_4256,N_3908,N_3912);
or U4257 (N_4257,N_3870,N_3677);
nand U4258 (N_4258,N_3674,N_3875);
nor U4259 (N_4259,N_3742,N_3876);
nand U4260 (N_4260,N_3890,N_3953);
or U4261 (N_4261,N_3834,N_3984);
and U4262 (N_4262,N_3735,N_3731);
nand U4263 (N_4263,N_3572,N_3535);
nor U4264 (N_4264,N_3558,N_3628);
or U4265 (N_4265,N_3679,N_3763);
nor U4266 (N_4266,N_3798,N_3504);
or U4267 (N_4267,N_3928,N_3788);
and U4268 (N_4268,N_3593,N_3884);
nand U4269 (N_4269,N_3930,N_3730);
and U4270 (N_4270,N_3821,N_3808);
nor U4271 (N_4271,N_3896,N_3812);
or U4272 (N_4272,N_3881,N_3558);
nand U4273 (N_4273,N_3913,N_3880);
or U4274 (N_4274,N_3956,N_3552);
or U4275 (N_4275,N_3943,N_3650);
or U4276 (N_4276,N_3889,N_3728);
nor U4277 (N_4277,N_3597,N_3537);
nor U4278 (N_4278,N_3693,N_3552);
or U4279 (N_4279,N_3869,N_3919);
or U4280 (N_4280,N_3646,N_3990);
nor U4281 (N_4281,N_3813,N_3990);
or U4282 (N_4282,N_3700,N_3528);
nor U4283 (N_4283,N_3864,N_3585);
nand U4284 (N_4284,N_3593,N_3507);
or U4285 (N_4285,N_3962,N_3761);
or U4286 (N_4286,N_3554,N_3884);
and U4287 (N_4287,N_3855,N_3554);
and U4288 (N_4288,N_3681,N_3984);
and U4289 (N_4289,N_3639,N_3976);
nor U4290 (N_4290,N_3930,N_3926);
or U4291 (N_4291,N_3617,N_3696);
nand U4292 (N_4292,N_3600,N_3554);
nand U4293 (N_4293,N_3848,N_3558);
nor U4294 (N_4294,N_3584,N_3805);
or U4295 (N_4295,N_3625,N_3830);
nand U4296 (N_4296,N_3561,N_3626);
nor U4297 (N_4297,N_3528,N_3612);
nor U4298 (N_4298,N_3602,N_3559);
nor U4299 (N_4299,N_3816,N_3895);
nand U4300 (N_4300,N_3596,N_3611);
nand U4301 (N_4301,N_3621,N_3573);
nand U4302 (N_4302,N_3701,N_3707);
nand U4303 (N_4303,N_3843,N_3685);
or U4304 (N_4304,N_3762,N_3864);
or U4305 (N_4305,N_3632,N_3654);
xor U4306 (N_4306,N_3947,N_3859);
nand U4307 (N_4307,N_3573,N_3871);
and U4308 (N_4308,N_3810,N_3614);
or U4309 (N_4309,N_3835,N_3512);
nand U4310 (N_4310,N_3932,N_3715);
nor U4311 (N_4311,N_3715,N_3599);
nand U4312 (N_4312,N_3542,N_3549);
xor U4313 (N_4313,N_3721,N_3978);
or U4314 (N_4314,N_3953,N_3960);
nand U4315 (N_4315,N_3582,N_3726);
nor U4316 (N_4316,N_3950,N_3980);
and U4317 (N_4317,N_3774,N_3522);
or U4318 (N_4318,N_3818,N_3657);
or U4319 (N_4319,N_3642,N_3592);
nor U4320 (N_4320,N_3689,N_3602);
or U4321 (N_4321,N_3917,N_3822);
nand U4322 (N_4322,N_3588,N_3861);
or U4323 (N_4323,N_3640,N_3785);
or U4324 (N_4324,N_3905,N_3569);
and U4325 (N_4325,N_3927,N_3588);
and U4326 (N_4326,N_3980,N_3854);
or U4327 (N_4327,N_3669,N_3536);
or U4328 (N_4328,N_3647,N_3637);
and U4329 (N_4329,N_3602,N_3841);
nand U4330 (N_4330,N_3825,N_3554);
or U4331 (N_4331,N_3837,N_3973);
nand U4332 (N_4332,N_3904,N_3759);
nor U4333 (N_4333,N_3545,N_3699);
nand U4334 (N_4334,N_3620,N_3881);
nand U4335 (N_4335,N_3754,N_3551);
xnor U4336 (N_4336,N_3851,N_3702);
nor U4337 (N_4337,N_3659,N_3898);
or U4338 (N_4338,N_3748,N_3904);
and U4339 (N_4339,N_3501,N_3592);
and U4340 (N_4340,N_3999,N_3778);
and U4341 (N_4341,N_3995,N_3601);
or U4342 (N_4342,N_3996,N_3727);
and U4343 (N_4343,N_3847,N_3976);
nand U4344 (N_4344,N_3817,N_3571);
and U4345 (N_4345,N_3578,N_3560);
or U4346 (N_4346,N_3842,N_3792);
and U4347 (N_4347,N_3787,N_3932);
or U4348 (N_4348,N_3535,N_3759);
and U4349 (N_4349,N_3880,N_3685);
or U4350 (N_4350,N_3871,N_3742);
nand U4351 (N_4351,N_3999,N_3912);
nor U4352 (N_4352,N_3852,N_3647);
and U4353 (N_4353,N_3821,N_3874);
or U4354 (N_4354,N_3875,N_3639);
and U4355 (N_4355,N_3897,N_3584);
nand U4356 (N_4356,N_3975,N_3596);
nor U4357 (N_4357,N_3757,N_3789);
nor U4358 (N_4358,N_3746,N_3803);
and U4359 (N_4359,N_3586,N_3750);
and U4360 (N_4360,N_3908,N_3581);
nand U4361 (N_4361,N_3815,N_3924);
or U4362 (N_4362,N_3698,N_3801);
nand U4363 (N_4363,N_3521,N_3535);
or U4364 (N_4364,N_3665,N_3620);
xnor U4365 (N_4365,N_3519,N_3978);
nor U4366 (N_4366,N_3586,N_3659);
nand U4367 (N_4367,N_3820,N_3629);
or U4368 (N_4368,N_3901,N_3880);
or U4369 (N_4369,N_3995,N_3955);
nor U4370 (N_4370,N_3845,N_3728);
nor U4371 (N_4371,N_3727,N_3758);
xor U4372 (N_4372,N_3524,N_3720);
nor U4373 (N_4373,N_3533,N_3701);
or U4374 (N_4374,N_3788,N_3712);
nor U4375 (N_4375,N_3569,N_3584);
nand U4376 (N_4376,N_3791,N_3906);
nor U4377 (N_4377,N_3788,N_3925);
nor U4378 (N_4378,N_3976,N_3505);
or U4379 (N_4379,N_3912,N_3748);
and U4380 (N_4380,N_3754,N_3593);
or U4381 (N_4381,N_3867,N_3905);
and U4382 (N_4382,N_3520,N_3701);
nand U4383 (N_4383,N_3814,N_3888);
or U4384 (N_4384,N_3753,N_3762);
and U4385 (N_4385,N_3682,N_3844);
nor U4386 (N_4386,N_3621,N_3947);
nand U4387 (N_4387,N_3766,N_3524);
nor U4388 (N_4388,N_3967,N_3510);
nor U4389 (N_4389,N_3503,N_3890);
nor U4390 (N_4390,N_3553,N_3995);
nor U4391 (N_4391,N_3723,N_3903);
or U4392 (N_4392,N_3925,N_3666);
or U4393 (N_4393,N_3904,N_3757);
and U4394 (N_4394,N_3715,N_3577);
and U4395 (N_4395,N_3957,N_3609);
nand U4396 (N_4396,N_3604,N_3550);
or U4397 (N_4397,N_3973,N_3525);
or U4398 (N_4398,N_3879,N_3614);
or U4399 (N_4399,N_3992,N_3891);
and U4400 (N_4400,N_3787,N_3937);
or U4401 (N_4401,N_3818,N_3543);
nand U4402 (N_4402,N_3676,N_3891);
or U4403 (N_4403,N_3554,N_3988);
nand U4404 (N_4404,N_3505,N_3751);
nand U4405 (N_4405,N_3624,N_3745);
and U4406 (N_4406,N_3518,N_3593);
and U4407 (N_4407,N_3549,N_3703);
or U4408 (N_4408,N_3705,N_3955);
xnor U4409 (N_4409,N_3622,N_3947);
nor U4410 (N_4410,N_3953,N_3989);
nand U4411 (N_4411,N_3732,N_3929);
nor U4412 (N_4412,N_3703,N_3690);
nand U4413 (N_4413,N_3726,N_3550);
and U4414 (N_4414,N_3872,N_3960);
and U4415 (N_4415,N_3592,N_3601);
or U4416 (N_4416,N_3534,N_3804);
nor U4417 (N_4417,N_3593,N_3620);
and U4418 (N_4418,N_3857,N_3762);
nand U4419 (N_4419,N_3783,N_3596);
and U4420 (N_4420,N_3766,N_3507);
and U4421 (N_4421,N_3658,N_3517);
or U4422 (N_4422,N_3810,N_3700);
nand U4423 (N_4423,N_3591,N_3778);
or U4424 (N_4424,N_3551,N_3842);
and U4425 (N_4425,N_3884,N_3980);
and U4426 (N_4426,N_3724,N_3950);
nor U4427 (N_4427,N_3977,N_3597);
or U4428 (N_4428,N_3717,N_3586);
nor U4429 (N_4429,N_3900,N_3702);
or U4430 (N_4430,N_3935,N_3609);
nand U4431 (N_4431,N_3727,N_3822);
or U4432 (N_4432,N_3822,N_3722);
and U4433 (N_4433,N_3827,N_3513);
nor U4434 (N_4434,N_3516,N_3615);
or U4435 (N_4435,N_3673,N_3661);
nor U4436 (N_4436,N_3540,N_3909);
or U4437 (N_4437,N_3666,N_3513);
nand U4438 (N_4438,N_3895,N_3964);
nor U4439 (N_4439,N_3739,N_3562);
nand U4440 (N_4440,N_3694,N_3845);
nor U4441 (N_4441,N_3721,N_3778);
nand U4442 (N_4442,N_3931,N_3951);
nor U4443 (N_4443,N_3633,N_3577);
nand U4444 (N_4444,N_3512,N_3840);
nor U4445 (N_4445,N_3953,N_3570);
and U4446 (N_4446,N_3932,N_3977);
and U4447 (N_4447,N_3633,N_3874);
nor U4448 (N_4448,N_3619,N_3987);
or U4449 (N_4449,N_3514,N_3994);
nor U4450 (N_4450,N_3855,N_3877);
nor U4451 (N_4451,N_3777,N_3596);
or U4452 (N_4452,N_3966,N_3820);
and U4453 (N_4453,N_3562,N_3555);
nand U4454 (N_4454,N_3976,N_3595);
nor U4455 (N_4455,N_3783,N_3646);
or U4456 (N_4456,N_3870,N_3833);
or U4457 (N_4457,N_3714,N_3531);
or U4458 (N_4458,N_3862,N_3880);
nor U4459 (N_4459,N_3862,N_3630);
or U4460 (N_4460,N_3589,N_3731);
or U4461 (N_4461,N_3512,N_3787);
nor U4462 (N_4462,N_3615,N_3750);
or U4463 (N_4463,N_3686,N_3674);
nand U4464 (N_4464,N_3744,N_3835);
nor U4465 (N_4465,N_3752,N_3851);
nand U4466 (N_4466,N_3575,N_3888);
and U4467 (N_4467,N_3748,N_3632);
nor U4468 (N_4468,N_3518,N_3945);
nor U4469 (N_4469,N_3696,N_3508);
nand U4470 (N_4470,N_3685,N_3986);
and U4471 (N_4471,N_3744,N_3819);
and U4472 (N_4472,N_3532,N_3692);
nand U4473 (N_4473,N_3584,N_3655);
nor U4474 (N_4474,N_3769,N_3686);
nand U4475 (N_4475,N_3778,N_3541);
or U4476 (N_4476,N_3749,N_3565);
nor U4477 (N_4477,N_3927,N_3986);
and U4478 (N_4478,N_3839,N_3714);
nor U4479 (N_4479,N_3694,N_3720);
xor U4480 (N_4480,N_3556,N_3824);
or U4481 (N_4481,N_3935,N_3668);
or U4482 (N_4482,N_3585,N_3721);
nor U4483 (N_4483,N_3831,N_3575);
and U4484 (N_4484,N_3614,N_3772);
and U4485 (N_4485,N_3811,N_3681);
nand U4486 (N_4486,N_3940,N_3508);
or U4487 (N_4487,N_3787,N_3608);
or U4488 (N_4488,N_3914,N_3813);
or U4489 (N_4489,N_3848,N_3998);
and U4490 (N_4490,N_3865,N_3798);
and U4491 (N_4491,N_3977,N_3642);
or U4492 (N_4492,N_3858,N_3827);
and U4493 (N_4493,N_3907,N_3584);
or U4494 (N_4494,N_3729,N_3635);
or U4495 (N_4495,N_3765,N_3662);
xnor U4496 (N_4496,N_3651,N_3926);
nor U4497 (N_4497,N_3754,N_3716);
nor U4498 (N_4498,N_3764,N_3996);
or U4499 (N_4499,N_3572,N_3943);
and U4500 (N_4500,N_4238,N_4399);
or U4501 (N_4501,N_4217,N_4301);
and U4502 (N_4502,N_4044,N_4009);
and U4503 (N_4503,N_4432,N_4237);
nor U4504 (N_4504,N_4265,N_4428);
and U4505 (N_4505,N_4156,N_4325);
or U4506 (N_4506,N_4283,N_4305);
nor U4507 (N_4507,N_4434,N_4048);
nor U4508 (N_4508,N_4057,N_4425);
nand U4509 (N_4509,N_4137,N_4060);
nor U4510 (N_4510,N_4133,N_4210);
and U4511 (N_4511,N_4069,N_4333);
or U4512 (N_4512,N_4151,N_4370);
and U4513 (N_4513,N_4066,N_4355);
or U4514 (N_4514,N_4036,N_4143);
nor U4515 (N_4515,N_4209,N_4000);
nand U4516 (N_4516,N_4170,N_4337);
or U4517 (N_4517,N_4465,N_4172);
nor U4518 (N_4518,N_4158,N_4216);
nor U4519 (N_4519,N_4456,N_4096);
and U4520 (N_4520,N_4250,N_4351);
or U4521 (N_4521,N_4336,N_4352);
nor U4522 (N_4522,N_4202,N_4068);
nor U4523 (N_4523,N_4065,N_4478);
nand U4524 (N_4524,N_4436,N_4472);
or U4525 (N_4525,N_4244,N_4341);
nand U4526 (N_4526,N_4225,N_4397);
and U4527 (N_4527,N_4037,N_4464);
nor U4528 (N_4528,N_4412,N_4014);
nor U4529 (N_4529,N_4086,N_4414);
xor U4530 (N_4530,N_4163,N_4299);
nand U4531 (N_4531,N_4422,N_4294);
nand U4532 (N_4532,N_4201,N_4362);
nor U4533 (N_4533,N_4282,N_4171);
xor U4534 (N_4534,N_4179,N_4120);
or U4535 (N_4535,N_4103,N_4295);
and U4536 (N_4536,N_4124,N_4175);
or U4537 (N_4537,N_4296,N_4186);
nor U4538 (N_4538,N_4426,N_4369);
nand U4539 (N_4539,N_4273,N_4184);
or U4540 (N_4540,N_4197,N_4485);
nand U4541 (N_4541,N_4483,N_4398);
nor U4542 (N_4542,N_4307,N_4098);
nand U4543 (N_4543,N_4257,N_4125);
nor U4544 (N_4544,N_4200,N_4415);
or U4545 (N_4545,N_4473,N_4017);
or U4546 (N_4546,N_4329,N_4354);
and U4547 (N_4547,N_4286,N_4361);
or U4548 (N_4548,N_4018,N_4338);
or U4549 (N_4549,N_4168,N_4013);
nand U4550 (N_4550,N_4330,N_4020);
or U4551 (N_4551,N_4302,N_4012);
and U4552 (N_4552,N_4052,N_4039);
or U4553 (N_4553,N_4107,N_4499);
nor U4554 (N_4554,N_4387,N_4240);
xnor U4555 (N_4555,N_4488,N_4291);
and U4556 (N_4556,N_4350,N_4061);
or U4557 (N_4557,N_4450,N_4167);
or U4558 (N_4558,N_4093,N_4384);
or U4559 (N_4559,N_4375,N_4342);
nand U4560 (N_4560,N_4034,N_4223);
or U4561 (N_4561,N_4391,N_4471);
or U4562 (N_4562,N_4259,N_4180);
and U4563 (N_4563,N_4188,N_4409);
and U4564 (N_4564,N_4251,N_4042);
or U4565 (N_4565,N_4453,N_4372);
and U4566 (N_4566,N_4208,N_4139);
nand U4567 (N_4567,N_4359,N_4314);
or U4568 (N_4568,N_4319,N_4152);
or U4569 (N_4569,N_4264,N_4493);
and U4570 (N_4570,N_4497,N_4262);
nand U4571 (N_4571,N_4451,N_4236);
and U4572 (N_4572,N_4082,N_4038);
or U4573 (N_4573,N_4430,N_4027);
nand U4574 (N_4574,N_4468,N_4281);
xnor U4575 (N_4575,N_4335,N_4444);
and U4576 (N_4576,N_4476,N_4081);
and U4577 (N_4577,N_4160,N_4449);
or U4578 (N_4578,N_4374,N_4150);
nand U4579 (N_4579,N_4418,N_4470);
or U4580 (N_4580,N_4356,N_4275);
or U4581 (N_4581,N_4187,N_4058);
and U4582 (N_4582,N_4241,N_4255);
or U4583 (N_4583,N_4317,N_4182);
nand U4584 (N_4584,N_4119,N_4343);
nand U4585 (N_4585,N_4407,N_4106);
or U4586 (N_4586,N_4159,N_4326);
or U4587 (N_4587,N_4490,N_4443);
nand U4588 (N_4588,N_4191,N_4452);
and U4589 (N_4589,N_4353,N_4248);
nor U4590 (N_4590,N_4463,N_4292);
nor U4591 (N_4591,N_4113,N_4222);
nand U4592 (N_4592,N_4141,N_4166);
and U4593 (N_4593,N_4123,N_4339);
nor U4594 (N_4594,N_4177,N_4029);
and U4595 (N_4595,N_4035,N_4135);
and U4596 (N_4596,N_4108,N_4489);
nand U4597 (N_4597,N_4131,N_4145);
nand U4598 (N_4598,N_4122,N_4173);
or U4599 (N_4599,N_4234,N_4115);
nand U4600 (N_4600,N_4388,N_4019);
nor U4601 (N_4601,N_4230,N_4393);
and U4602 (N_4602,N_4270,N_4461);
and U4603 (N_4603,N_4114,N_4348);
and U4604 (N_4604,N_4097,N_4022);
nor U4605 (N_4605,N_4192,N_4161);
nand U4606 (N_4606,N_4126,N_4015);
and U4607 (N_4607,N_4056,N_4381);
or U4608 (N_4608,N_4153,N_4303);
and U4609 (N_4609,N_4274,N_4331);
and U4610 (N_4610,N_4357,N_4079);
nor U4611 (N_4611,N_4261,N_4417);
and U4612 (N_4612,N_4363,N_4072);
or U4613 (N_4613,N_4232,N_4205);
nand U4614 (N_4614,N_4376,N_4423);
or U4615 (N_4615,N_4028,N_4030);
or U4616 (N_4616,N_4025,N_4204);
or U4617 (N_4617,N_4368,N_4413);
or U4618 (N_4618,N_4340,N_4227);
or U4619 (N_4619,N_4366,N_4117);
nor U4620 (N_4620,N_4406,N_4462);
and U4621 (N_4621,N_4053,N_4371);
nand U4622 (N_4622,N_4494,N_4040);
nand U4623 (N_4623,N_4466,N_4421);
nand U4624 (N_4624,N_4378,N_4334);
nor U4625 (N_4625,N_4440,N_4297);
and U4626 (N_4626,N_4380,N_4322);
xnor U4627 (N_4627,N_4190,N_4049);
nor U4628 (N_4628,N_4280,N_4147);
nor U4629 (N_4629,N_4112,N_4313);
or U4630 (N_4630,N_4311,N_4457);
xor U4631 (N_4631,N_4403,N_4401);
nand U4632 (N_4632,N_4074,N_4140);
nand U4633 (N_4633,N_4193,N_4320);
or U4634 (N_4634,N_4070,N_4142);
nand U4635 (N_4635,N_4385,N_4396);
and U4636 (N_4636,N_4071,N_4400);
nor U4637 (N_4637,N_4298,N_4454);
and U4638 (N_4638,N_4242,N_4001);
or U4639 (N_4639,N_4221,N_4395);
nand U4640 (N_4640,N_4149,N_4435);
nor U4641 (N_4641,N_4215,N_4101);
or U4642 (N_4642,N_4214,N_4116);
nor U4643 (N_4643,N_4469,N_4249);
nor U4644 (N_4644,N_4487,N_4185);
nand U4645 (N_4645,N_4136,N_4055);
or U4646 (N_4646,N_4031,N_4316);
or U4647 (N_4647,N_4105,N_4050);
nor U4648 (N_4648,N_4349,N_4008);
or U4649 (N_4649,N_4247,N_4196);
or U4650 (N_4650,N_4011,N_4383);
or U4651 (N_4651,N_4312,N_4392);
nor U4652 (N_4652,N_4382,N_4104);
and U4653 (N_4653,N_4345,N_4207);
or U4654 (N_4654,N_4373,N_4076);
nor U4655 (N_4655,N_4162,N_4344);
or U4656 (N_4656,N_4347,N_4279);
nor U4657 (N_4657,N_4441,N_4346);
nor U4658 (N_4658,N_4252,N_4007);
and U4659 (N_4659,N_4404,N_4367);
xnor U4660 (N_4660,N_4263,N_4491);
and U4661 (N_4661,N_4024,N_4364);
and U4662 (N_4662,N_4386,N_4220);
nor U4663 (N_4663,N_4181,N_4256);
or U4664 (N_4664,N_4475,N_4146);
nand U4665 (N_4665,N_4310,N_4431);
nor U4666 (N_4666,N_4455,N_4304);
nor U4667 (N_4667,N_4005,N_4051);
nor U4668 (N_4668,N_4445,N_4300);
nand U4669 (N_4669,N_4477,N_4138);
and U4670 (N_4670,N_4228,N_4067);
nor U4671 (N_4671,N_4258,N_4092);
or U4672 (N_4672,N_4267,N_4271);
nor U4673 (N_4673,N_4416,N_4004);
nor U4674 (N_4674,N_4481,N_4458);
or U4675 (N_4675,N_4046,N_4437);
nor U4676 (N_4676,N_4460,N_4266);
nor U4677 (N_4677,N_4144,N_4479);
or U4678 (N_4678,N_4110,N_4054);
nand U4679 (N_4679,N_4095,N_4402);
nand U4680 (N_4680,N_4023,N_4130);
and U4681 (N_4681,N_4287,N_4109);
nor U4682 (N_4682,N_4492,N_4411);
or U4683 (N_4683,N_4047,N_4010);
nand U4684 (N_4684,N_4498,N_4229);
nand U4685 (N_4685,N_4002,N_4219);
and U4686 (N_4686,N_4433,N_4148);
and U4687 (N_4687,N_4134,N_4064);
or U4688 (N_4688,N_4111,N_4006);
and U4689 (N_4689,N_4218,N_4100);
nand U4690 (N_4690,N_4429,N_4379);
nor U4691 (N_4691,N_4195,N_4077);
or U4692 (N_4692,N_4474,N_4089);
or U4693 (N_4693,N_4276,N_4408);
nand U4694 (N_4694,N_4360,N_4063);
and U4695 (N_4695,N_4269,N_4482);
nor U4696 (N_4696,N_4254,N_4278);
nand U4697 (N_4697,N_4243,N_4155);
or U4698 (N_4698,N_4327,N_4157);
nand U4699 (N_4699,N_4480,N_4021);
nand U4700 (N_4700,N_4448,N_4486);
and U4701 (N_4701,N_4211,N_4419);
nand U4702 (N_4702,N_4318,N_4164);
or U4703 (N_4703,N_4315,N_4099);
and U4704 (N_4704,N_4043,N_4003);
or U4705 (N_4705,N_4233,N_4213);
and U4706 (N_4706,N_4121,N_4459);
nand U4707 (N_4707,N_4041,N_4094);
and U4708 (N_4708,N_4189,N_4165);
and U4709 (N_4709,N_4442,N_4045);
nand U4710 (N_4710,N_4132,N_4154);
nand U4711 (N_4711,N_4088,N_4289);
and U4712 (N_4712,N_4212,N_4033);
or U4713 (N_4713,N_4206,N_4323);
nand U4714 (N_4714,N_4246,N_4328);
nand U4715 (N_4715,N_4467,N_4084);
and U4716 (N_4716,N_4394,N_4308);
nand U4717 (N_4717,N_4446,N_4389);
and U4718 (N_4718,N_4102,N_4231);
or U4719 (N_4719,N_4026,N_4427);
nand U4720 (N_4720,N_4176,N_4129);
nor U4721 (N_4721,N_4075,N_4226);
and U4722 (N_4722,N_4321,N_4253);
or U4723 (N_4723,N_4285,N_4324);
nand U4724 (N_4724,N_4484,N_4420);
nor U4725 (N_4725,N_4235,N_4016);
and U4726 (N_4726,N_4073,N_4224);
or U4727 (N_4727,N_4183,N_4090);
nand U4728 (N_4728,N_4080,N_4178);
or U4729 (N_4729,N_4174,N_4087);
nand U4730 (N_4730,N_4424,N_4260);
xnor U4731 (N_4731,N_4268,N_4239);
or U4732 (N_4732,N_4306,N_4377);
nor U4733 (N_4733,N_4083,N_4194);
nor U4734 (N_4734,N_4127,N_4390);
nand U4735 (N_4735,N_4078,N_4277);
or U4736 (N_4736,N_4438,N_4332);
and U4737 (N_4737,N_4059,N_4118);
and U4738 (N_4738,N_4309,N_4495);
nand U4739 (N_4739,N_4284,N_4410);
nor U4740 (N_4740,N_4439,N_4358);
and U4741 (N_4741,N_4365,N_4198);
nor U4742 (N_4742,N_4290,N_4128);
and U4743 (N_4743,N_4062,N_4272);
nor U4744 (N_4744,N_4203,N_4199);
or U4745 (N_4745,N_4245,N_4447);
nand U4746 (N_4746,N_4288,N_4032);
nor U4747 (N_4747,N_4169,N_4085);
or U4748 (N_4748,N_4405,N_4293);
and U4749 (N_4749,N_4496,N_4091);
or U4750 (N_4750,N_4335,N_4141);
nand U4751 (N_4751,N_4079,N_4027);
xnor U4752 (N_4752,N_4138,N_4316);
and U4753 (N_4753,N_4445,N_4456);
or U4754 (N_4754,N_4017,N_4089);
nor U4755 (N_4755,N_4309,N_4273);
nand U4756 (N_4756,N_4402,N_4074);
nand U4757 (N_4757,N_4165,N_4344);
nor U4758 (N_4758,N_4171,N_4312);
and U4759 (N_4759,N_4431,N_4358);
nand U4760 (N_4760,N_4213,N_4270);
nand U4761 (N_4761,N_4012,N_4470);
and U4762 (N_4762,N_4473,N_4135);
nand U4763 (N_4763,N_4099,N_4190);
nand U4764 (N_4764,N_4432,N_4369);
nand U4765 (N_4765,N_4182,N_4315);
nor U4766 (N_4766,N_4113,N_4279);
nor U4767 (N_4767,N_4254,N_4411);
and U4768 (N_4768,N_4487,N_4142);
nor U4769 (N_4769,N_4302,N_4269);
nand U4770 (N_4770,N_4416,N_4327);
or U4771 (N_4771,N_4144,N_4256);
nor U4772 (N_4772,N_4163,N_4087);
nand U4773 (N_4773,N_4402,N_4257);
and U4774 (N_4774,N_4208,N_4031);
or U4775 (N_4775,N_4005,N_4070);
nand U4776 (N_4776,N_4481,N_4346);
nand U4777 (N_4777,N_4318,N_4299);
or U4778 (N_4778,N_4085,N_4322);
nor U4779 (N_4779,N_4476,N_4117);
or U4780 (N_4780,N_4043,N_4097);
and U4781 (N_4781,N_4281,N_4030);
and U4782 (N_4782,N_4004,N_4260);
nor U4783 (N_4783,N_4408,N_4462);
nand U4784 (N_4784,N_4126,N_4289);
and U4785 (N_4785,N_4023,N_4024);
nor U4786 (N_4786,N_4026,N_4153);
or U4787 (N_4787,N_4067,N_4244);
and U4788 (N_4788,N_4169,N_4235);
nor U4789 (N_4789,N_4233,N_4345);
nand U4790 (N_4790,N_4078,N_4233);
nand U4791 (N_4791,N_4304,N_4044);
nand U4792 (N_4792,N_4478,N_4203);
nand U4793 (N_4793,N_4112,N_4404);
nor U4794 (N_4794,N_4167,N_4453);
nor U4795 (N_4795,N_4025,N_4356);
nor U4796 (N_4796,N_4358,N_4155);
nand U4797 (N_4797,N_4411,N_4021);
nor U4798 (N_4798,N_4477,N_4162);
or U4799 (N_4799,N_4441,N_4149);
or U4800 (N_4800,N_4064,N_4415);
nand U4801 (N_4801,N_4167,N_4108);
nor U4802 (N_4802,N_4171,N_4097);
or U4803 (N_4803,N_4483,N_4281);
nor U4804 (N_4804,N_4325,N_4093);
nand U4805 (N_4805,N_4204,N_4097);
nand U4806 (N_4806,N_4123,N_4037);
nor U4807 (N_4807,N_4234,N_4107);
nor U4808 (N_4808,N_4345,N_4461);
xnor U4809 (N_4809,N_4392,N_4288);
nand U4810 (N_4810,N_4483,N_4361);
nand U4811 (N_4811,N_4140,N_4375);
and U4812 (N_4812,N_4499,N_4323);
or U4813 (N_4813,N_4197,N_4091);
nand U4814 (N_4814,N_4367,N_4456);
nand U4815 (N_4815,N_4138,N_4366);
or U4816 (N_4816,N_4266,N_4030);
nor U4817 (N_4817,N_4129,N_4204);
or U4818 (N_4818,N_4474,N_4048);
or U4819 (N_4819,N_4340,N_4352);
or U4820 (N_4820,N_4205,N_4040);
or U4821 (N_4821,N_4145,N_4435);
and U4822 (N_4822,N_4178,N_4055);
nor U4823 (N_4823,N_4148,N_4120);
or U4824 (N_4824,N_4110,N_4412);
nand U4825 (N_4825,N_4331,N_4498);
and U4826 (N_4826,N_4212,N_4070);
and U4827 (N_4827,N_4178,N_4083);
nor U4828 (N_4828,N_4065,N_4372);
nor U4829 (N_4829,N_4433,N_4179);
and U4830 (N_4830,N_4203,N_4482);
nand U4831 (N_4831,N_4187,N_4134);
and U4832 (N_4832,N_4181,N_4073);
nor U4833 (N_4833,N_4075,N_4341);
or U4834 (N_4834,N_4111,N_4341);
nor U4835 (N_4835,N_4101,N_4485);
nand U4836 (N_4836,N_4453,N_4182);
and U4837 (N_4837,N_4080,N_4159);
nor U4838 (N_4838,N_4309,N_4161);
and U4839 (N_4839,N_4222,N_4283);
and U4840 (N_4840,N_4334,N_4166);
and U4841 (N_4841,N_4405,N_4245);
and U4842 (N_4842,N_4392,N_4448);
xor U4843 (N_4843,N_4166,N_4259);
nor U4844 (N_4844,N_4191,N_4348);
and U4845 (N_4845,N_4441,N_4181);
or U4846 (N_4846,N_4116,N_4482);
nor U4847 (N_4847,N_4176,N_4457);
nand U4848 (N_4848,N_4319,N_4269);
and U4849 (N_4849,N_4284,N_4374);
nor U4850 (N_4850,N_4067,N_4063);
and U4851 (N_4851,N_4283,N_4149);
xor U4852 (N_4852,N_4114,N_4197);
or U4853 (N_4853,N_4322,N_4395);
nand U4854 (N_4854,N_4352,N_4321);
nor U4855 (N_4855,N_4023,N_4403);
nor U4856 (N_4856,N_4270,N_4084);
nand U4857 (N_4857,N_4494,N_4340);
nor U4858 (N_4858,N_4202,N_4259);
nand U4859 (N_4859,N_4440,N_4087);
nand U4860 (N_4860,N_4297,N_4249);
nor U4861 (N_4861,N_4491,N_4155);
or U4862 (N_4862,N_4468,N_4119);
nor U4863 (N_4863,N_4204,N_4401);
nor U4864 (N_4864,N_4328,N_4445);
or U4865 (N_4865,N_4336,N_4232);
and U4866 (N_4866,N_4223,N_4126);
or U4867 (N_4867,N_4035,N_4238);
nand U4868 (N_4868,N_4420,N_4487);
nor U4869 (N_4869,N_4312,N_4172);
and U4870 (N_4870,N_4340,N_4388);
and U4871 (N_4871,N_4418,N_4380);
and U4872 (N_4872,N_4251,N_4275);
and U4873 (N_4873,N_4263,N_4115);
or U4874 (N_4874,N_4403,N_4235);
xor U4875 (N_4875,N_4071,N_4489);
nand U4876 (N_4876,N_4409,N_4195);
or U4877 (N_4877,N_4321,N_4460);
nor U4878 (N_4878,N_4412,N_4099);
nor U4879 (N_4879,N_4377,N_4441);
nand U4880 (N_4880,N_4374,N_4411);
nand U4881 (N_4881,N_4424,N_4134);
and U4882 (N_4882,N_4126,N_4333);
or U4883 (N_4883,N_4131,N_4492);
or U4884 (N_4884,N_4476,N_4268);
nor U4885 (N_4885,N_4188,N_4387);
and U4886 (N_4886,N_4194,N_4231);
nand U4887 (N_4887,N_4428,N_4053);
nor U4888 (N_4888,N_4061,N_4097);
xnor U4889 (N_4889,N_4063,N_4441);
or U4890 (N_4890,N_4007,N_4173);
nand U4891 (N_4891,N_4303,N_4077);
and U4892 (N_4892,N_4093,N_4414);
nand U4893 (N_4893,N_4352,N_4186);
nand U4894 (N_4894,N_4013,N_4262);
nand U4895 (N_4895,N_4008,N_4089);
nor U4896 (N_4896,N_4076,N_4228);
nand U4897 (N_4897,N_4022,N_4236);
and U4898 (N_4898,N_4239,N_4080);
nand U4899 (N_4899,N_4250,N_4255);
or U4900 (N_4900,N_4291,N_4052);
nand U4901 (N_4901,N_4074,N_4263);
or U4902 (N_4902,N_4159,N_4078);
nand U4903 (N_4903,N_4203,N_4368);
nor U4904 (N_4904,N_4152,N_4320);
nor U4905 (N_4905,N_4084,N_4097);
or U4906 (N_4906,N_4013,N_4375);
or U4907 (N_4907,N_4390,N_4418);
or U4908 (N_4908,N_4318,N_4265);
or U4909 (N_4909,N_4047,N_4323);
xnor U4910 (N_4910,N_4360,N_4104);
or U4911 (N_4911,N_4234,N_4213);
nor U4912 (N_4912,N_4082,N_4351);
nor U4913 (N_4913,N_4435,N_4282);
nor U4914 (N_4914,N_4347,N_4129);
nor U4915 (N_4915,N_4259,N_4255);
or U4916 (N_4916,N_4453,N_4407);
or U4917 (N_4917,N_4498,N_4435);
or U4918 (N_4918,N_4000,N_4394);
and U4919 (N_4919,N_4167,N_4267);
and U4920 (N_4920,N_4177,N_4160);
nor U4921 (N_4921,N_4068,N_4257);
or U4922 (N_4922,N_4126,N_4036);
or U4923 (N_4923,N_4231,N_4270);
xnor U4924 (N_4924,N_4263,N_4249);
and U4925 (N_4925,N_4093,N_4209);
nor U4926 (N_4926,N_4438,N_4288);
or U4927 (N_4927,N_4364,N_4313);
or U4928 (N_4928,N_4361,N_4166);
nand U4929 (N_4929,N_4179,N_4026);
or U4930 (N_4930,N_4305,N_4418);
or U4931 (N_4931,N_4120,N_4188);
nand U4932 (N_4932,N_4250,N_4383);
and U4933 (N_4933,N_4061,N_4096);
xor U4934 (N_4934,N_4402,N_4309);
nor U4935 (N_4935,N_4128,N_4035);
and U4936 (N_4936,N_4077,N_4322);
nand U4937 (N_4937,N_4190,N_4271);
nor U4938 (N_4938,N_4116,N_4240);
nand U4939 (N_4939,N_4337,N_4142);
nand U4940 (N_4940,N_4063,N_4012);
nor U4941 (N_4941,N_4089,N_4082);
nand U4942 (N_4942,N_4292,N_4020);
and U4943 (N_4943,N_4198,N_4469);
nand U4944 (N_4944,N_4236,N_4437);
nor U4945 (N_4945,N_4213,N_4126);
nor U4946 (N_4946,N_4459,N_4342);
and U4947 (N_4947,N_4167,N_4285);
and U4948 (N_4948,N_4173,N_4234);
or U4949 (N_4949,N_4149,N_4064);
or U4950 (N_4950,N_4422,N_4090);
nor U4951 (N_4951,N_4201,N_4471);
nor U4952 (N_4952,N_4070,N_4031);
nand U4953 (N_4953,N_4371,N_4376);
and U4954 (N_4954,N_4186,N_4372);
nor U4955 (N_4955,N_4483,N_4073);
nor U4956 (N_4956,N_4385,N_4050);
and U4957 (N_4957,N_4240,N_4437);
nor U4958 (N_4958,N_4199,N_4208);
or U4959 (N_4959,N_4113,N_4190);
or U4960 (N_4960,N_4275,N_4307);
nand U4961 (N_4961,N_4483,N_4358);
nor U4962 (N_4962,N_4467,N_4342);
nand U4963 (N_4963,N_4151,N_4085);
and U4964 (N_4964,N_4451,N_4135);
nand U4965 (N_4965,N_4496,N_4051);
or U4966 (N_4966,N_4132,N_4125);
and U4967 (N_4967,N_4070,N_4103);
or U4968 (N_4968,N_4051,N_4465);
nor U4969 (N_4969,N_4039,N_4258);
nand U4970 (N_4970,N_4017,N_4016);
nand U4971 (N_4971,N_4060,N_4094);
and U4972 (N_4972,N_4403,N_4212);
nand U4973 (N_4973,N_4105,N_4024);
nor U4974 (N_4974,N_4200,N_4467);
or U4975 (N_4975,N_4251,N_4329);
or U4976 (N_4976,N_4040,N_4118);
nor U4977 (N_4977,N_4330,N_4288);
and U4978 (N_4978,N_4403,N_4057);
and U4979 (N_4979,N_4217,N_4219);
nand U4980 (N_4980,N_4264,N_4027);
or U4981 (N_4981,N_4162,N_4370);
nand U4982 (N_4982,N_4160,N_4140);
and U4983 (N_4983,N_4196,N_4458);
nor U4984 (N_4984,N_4333,N_4287);
nor U4985 (N_4985,N_4257,N_4197);
nand U4986 (N_4986,N_4442,N_4096);
or U4987 (N_4987,N_4252,N_4397);
or U4988 (N_4988,N_4430,N_4168);
nand U4989 (N_4989,N_4161,N_4408);
nor U4990 (N_4990,N_4328,N_4007);
xor U4991 (N_4991,N_4050,N_4372);
or U4992 (N_4992,N_4492,N_4406);
or U4993 (N_4993,N_4064,N_4247);
and U4994 (N_4994,N_4332,N_4147);
and U4995 (N_4995,N_4344,N_4464);
nand U4996 (N_4996,N_4149,N_4418);
xor U4997 (N_4997,N_4260,N_4458);
and U4998 (N_4998,N_4285,N_4039);
nor U4999 (N_4999,N_4458,N_4152);
or UO_0 (O_0,N_4793,N_4872);
or UO_1 (O_1,N_4795,N_4950);
and UO_2 (O_2,N_4749,N_4623);
xnor UO_3 (O_3,N_4617,N_4952);
or UO_4 (O_4,N_4674,N_4896);
and UO_5 (O_5,N_4788,N_4994);
or UO_6 (O_6,N_4846,N_4669);
xnor UO_7 (O_7,N_4957,N_4739);
or UO_8 (O_8,N_4848,N_4721);
and UO_9 (O_9,N_4507,N_4620);
or UO_10 (O_10,N_4890,N_4999);
or UO_11 (O_11,N_4907,N_4947);
nor UO_12 (O_12,N_4933,N_4987);
nor UO_13 (O_13,N_4984,N_4975);
or UO_14 (O_14,N_4518,N_4819);
or UO_15 (O_15,N_4608,N_4966);
xor UO_16 (O_16,N_4857,N_4672);
and UO_17 (O_17,N_4718,N_4550);
nand UO_18 (O_18,N_4546,N_4508);
nor UO_19 (O_19,N_4610,N_4934);
and UO_20 (O_20,N_4666,N_4910);
nor UO_21 (O_21,N_4536,N_4554);
nand UO_22 (O_22,N_4866,N_4959);
nand UO_23 (O_23,N_4943,N_4563);
or UO_24 (O_24,N_4722,N_4501);
nand UO_25 (O_25,N_4525,N_4790);
nor UO_26 (O_26,N_4542,N_4825);
nor UO_27 (O_27,N_4515,N_4811);
and UO_28 (O_28,N_4626,N_4621);
and UO_29 (O_29,N_4551,N_4919);
nor UO_30 (O_30,N_4500,N_4644);
and UO_31 (O_31,N_4662,N_4660);
or UO_32 (O_32,N_4632,N_4742);
nand UO_33 (O_33,N_4821,N_4600);
or UO_34 (O_34,N_4572,N_4653);
xnor UO_35 (O_35,N_4937,N_4578);
or UO_36 (O_36,N_4614,N_4932);
nand UO_37 (O_37,N_4588,N_4510);
nand UO_38 (O_38,N_4897,N_4513);
nor UO_39 (O_39,N_4606,N_4983);
or UO_40 (O_40,N_4931,N_4687);
nor UO_41 (O_41,N_4949,N_4826);
and UO_42 (O_42,N_4690,N_4745);
nand UO_43 (O_43,N_4511,N_4831);
nor UO_44 (O_44,N_4695,N_4905);
nand UO_45 (O_45,N_4574,N_4523);
nor UO_46 (O_46,N_4991,N_4837);
or UO_47 (O_47,N_4516,N_4645);
nand UO_48 (O_48,N_4791,N_4858);
nor UO_49 (O_49,N_4961,N_4917);
or UO_50 (O_50,N_4703,N_4985);
nor UO_51 (O_51,N_4820,N_4719);
and UO_52 (O_52,N_4794,N_4878);
or UO_53 (O_53,N_4760,N_4899);
or UO_54 (O_54,N_4727,N_4571);
nand UO_55 (O_55,N_4834,N_4807);
nand UO_56 (O_56,N_4637,N_4861);
nand UO_57 (O_57,N_4816,N_4519);
and UO_58 (O_58,N_4928,N_4753);
nand UO_59 (O_59,N_4758,N_4969);
nand UO_60 (O_60,N_4589,N_4540);
or UO_61 (O_61,N_4971,N_4607);
or UO_62 (O_62,N_4895,N_4767);
nor UO_63 (O_63,N_4810,N_4775);
nor UO_64 (O_64,N_4527,N_4685);
and UO_65 (O_65,N_4786,N_4530);
and UO_66 (O_66,N_4988,N_4544);
nor UO_67 (O_67,N_4580,N_4534);
nand UO_68 (O_68,N_4676,N_4780);
nand UO_69 (O_69,N_4647,N_4938);
nor UO_70 (O_70,N_4747,N_4552);
or UO_71 (O_71,N_4770,N_4935);
or UO_72 (O_72,N_4888,N_4990);
and UO_73 (O_73,N_4643,N_4877);
nor UO_74 (O_74,N_4652,N_4512);
nand UO_75 (O_75,N_4893,N_4865);
nand UO_76 (O_76,N_4521,N_4976);
nor UO_77 (O_77,N_4989,N_4750);
nand UO_78 (O_78,N_4557,N_4978);
and UO_79 (O_79,N_4827,N_4867);
nand UO_80 (O_80,N_4651,N_4918);
or UO_81 (O_81,N_4913,N_4678);
nand UO_82 (O_82,N_4602,N_4879);
nand UO_83 (O_83,N_4716,N_4850);
nand UO_84 (O_84,N_4972,N_4680);
nand UO_85 (O_85,N_4843,N_4796);
xnor UO_86 (O_86,N_4828,N_4772);
nor UO_87 (O_87,N_4732,N_4693);
or UO_88 (O_88,N_4764,N_4956);
xor UO_89 (O_89,N_4936,N_4624);
or UO_90 (O_90,N_4586,N_4502);
nand UO_91 (O_91,N_4875,N_4777);
nand UO_92 (O_92,N_4691,N_4992);
nand UO_93 (O_93,N_4979,N_4964);
nor UO_94 (O_94,N_4616,N_4902);
nor UO_95 (O_95,N_4628,N_4668);
nand UO_96 (O_96,N_4731,N_4980);
and UO_97 (O_97,N_4582,N_4792);
or UO_98 (O_98,N_4892,N_4787);
or UO_99 (O_99,N_4562,N_4559);
nor UO_100 (O_100,N_4636,N_4667);
and UO_101 (O_101,N_4609,N_4532);
nand UO_102 (O_102,N_4684,N_4849);
nand UO_103 (O_103,N_4700,N_4830);
or UO_104 (O_104,N_4946,N_4520);
xnor UO_105 (O_105,N_4561,N_4973);
or UO_106 (O_106,N_4547,N_4661);
or UO_107 (O_107,N_4619,N_4939);
nor UO_108 (O_108,N_4744,N_4545);
or UO_109 (O_109,N_4748,N_4579);
or UO_110 (O_110,N_4640,N_4817);
nor UO_111 (O_111,N_4566,N_4771);
nand UO_112 (O_112,N_4577,N_4958);
and UO_113 (O_113,N_4862,N_4754);
nor UO_114 (O_114,N_4863,N_4555);
or UO_115 (O_115,N_4815,N_4945);
nor UO_116 (O_116,N_4798,N_4549);
nand UO_117 (O_117,N_4901,N_4675);
nand UO_118 (O_118,N_4911,N_4836);
nor UO_119 (O_119,N_4746,N_4997);
nand UO_120 (O_120,N_4597,N_4565);
nor UO_121 (O_121,N_4930,N_4738);
and UO_122 (O_122,N_4604,N_4853);
or UO_123 (O_123,N_4856,N_4755);
or UO_124 (O_124,N_4720,N_4974);
nor UO_125 (O_125,N_4648,N_4768);
nand UO_126 (O_126,N_4960,N_4942);
nor UO_127 (O_127,N_4638,N_4797);
or UO_128 (O_128,N_4735,N_4517);
nor UO_129 (O_129,N_4993,N_4649);
xnor UO_130 (O_130,N_4870,N_4965);
nand UO_131 (O_131,N_4708,N_4633);
nand UO_132 (O_132,N_4785,N_4977);
nand UO_133 (O_133,N_4522,N_4514);
nand UO_134 (O_134,N_4823,N_4524);
nor UO_135 (O_135,N_4528,N_4904);
nor UO_136 (O_136,N_4924,N_4809);
or UO_137 (O_137,N_4699,N_4506);
or UO_138 (O_138,N_4967,N_4963);
or UO_139 (O_139,N_4657,N_4835);
nand UO_140 (O_140,N_4541,N_4891);
nor UO_141 (O_141,N_4995,N_4576);
and UO_142 (O_142,N_4692,N_4779);
and UO_143 (O_143,N_4726,N_4923);
or UO_144 (O_144,N_4581,N_4646);
nand UO_145 (O_145,N_4629,N_4874);
nor UO_146 (O_146,N_4839,N_4740);
nor UO_147 (O_147,N_4951,N_4880);
xor UO_148 (O_148,N_4922,N_4886);
nor UO_149 (O_149,N_4812,N_4701);
and UO_150 (O_150,N_4885,N_4709);
nand UO_151 (O_151,N_4622,N_4635);
or UO_152 (O_152,N_4625,N_4808);
nor UO_153 (O_153,N_4603,N_4611);
or UO_154 (O_154,N_4766,N_4778);
or UO_155 (O_155,N_4906,N_4663);
or UO_156 (O_156,N_4587,N_4665);
and UO_157 (O_157,N_4583,N_4598);
xor UO_158 (O_158,N_4799,N_4761);
nor UO_159 (O_159,N_4654,N_4539);
and UO_160 (O_160,N_4682,N_4679);
and UO_161 (O_161,N_4671,N_4841);
xnor UO_162 (O_162,N_4864,N_4789);
nor UO_163 (O_163,N_4940,N_4915);
or UO_164 (O_164,N_4734,N_4529);
and UO_165 (O_165,N_4751,N_4822);
or UO_166 (O_166,N_4783,N_4929);
nand UO_167 (O_167,N_4650,N_4681);
or UO_168 (O_168,N_4504,N_4696);
or UO_169 (O_169,N_4655,N_4970);
and UO_170 (O_170,N_4543,N_4585);
nand UO_171 (O_171,N_4573,N_4535);
or UO_172 (O_172,N_4763,N_4509);
or UO_173 (O_173,N_4707,N_4714);
or UO_174 (O_174,N_4769,N_4756);
nor UO_175 (O_175,N_4531,N_4728);
and UO_176 (O_176,N_4968,N_4941);
nand UO_177 (O_177,N_4920,N_4833);
nor UO_178 (O_178,N_4800,N_4601);
and UO_179 (O_179,N_4774,N_4981);
nor UO_180 (O_180,N_4916,N_4677);
or UO_181 (O_181,N_4711,N_4802);
or UO_182 (O_182,N_4982,N_4723);
or UO_183 (O_183,N_4884,N_4715);
nand UO_184 (O_184,N_4845,N_4618);
and UO_185 (O_185,N_4824,N_4627);
or UO_186 (O_186,N_4847,N_4813);
nor UO_187 (O_187,N_4664,N_4526);
nor UO_188 (O_188,N_4832,N_4686);
nand UO_189 (O_189,N_4762,N_4962);
nand UO_190 (O_190,N_4613,N_4733);
nor UO_191 (O_191,N_4712,N_4925);
or UO_192 (O_192,N_4710,N_4590);
nand UO_193 (O_193,N_4752,N_4914);
and UO_194 (O_194,N_4605,N_4595);
or UO_195 (O_195,N_4683,N_4599);
nor UO_196 (O_196,N_4612,N_4903);
nor UO_197 (O_197,N_4986,N_4592);
and UO_198 (O_198,N_4730,N_4829);
or UO_199 (O_199,N_4656,N_4538);
or UO_200 (O_200,N_4805,N_4855);
or UO_201 (O_201,N_4505,N_4630);
or UO_202 (O_202,N_4954,N_4921);
nand UO_203 (O_203,N_4584,N_4537);
and UO_204 (O_204,N_4803,N_4871);
or UO_205 (O_205,N_4844,N_4804);
or UO_206 (O_206,N_4567,N_4704);
and UO_207 (O_207,N_4926,N_4729);
nor UO_208 (O_208,N_4898,N_4852);
nand UO_209 (O_209,N_4773,N_4670);
and UO_210 (O_210,N_4641,N_4909);
nand UO_211 (O_211,N_4781,N_4553);
nand UO_212 (O_212,N_4673,N_4503);
and UO_213 (O_213,N_4908,N_4876);
or UO_214 (O_214,N_4594,N_4998);
nor UO_215 (O_215,N_4570,N_4639);
xnor UO_216 (O_216,N_4694,N_4894);
or UO_217 (O_217,N_4806,N_4889);
and UO_218 (O_218,N_4702,N_4776);
nand UO_219 (O_219,N_4851,N_4569);
or UO_220 (O_220,N_4801,N_4568);
and UO_221 (O_221,N_4642,N_4873);
or UO_222 (O_222,N_4741,N_4996);
nor UO_223 (O_223,N_4944,N_4591);
or UO_224 (O_224,N_4658,N_4818);
or UO_225 (O_225,N_4759,N_4564);
nand UO_226 (O_226,N_4838,N_4724);
nor UO_227 (O_227,N_4688,N_4736);
or UO_228 (O_228,N_4713,N_4558);
xor UO_229 (O_229,N_4860,N_4782);
nand UO_230 (O_230,N_4955,N_4881);
xor UO_231 (O_231,N_4840,N_4927);
or UO_232 (O_232,N_4900,N_4757);
or UO_233 (O_233,N_4953,N_4883);
and UO_234 (O_234,N_4689,N_4548);
or UO_235 (O_235,N_4869,N_4887);
nor UO_236 (O_236,N_4615,N_4706);
nand UO_237 (O_237,N_4717,N_4705);
or UO_238 (O_238,N_4725,N_4634);
and UO_239 (O_239,N_4631,N_4743);
nand UO_240 (O_240,N_4859,N_4533);
and UO_241 (O_241,N_4560,N_4659);
and UO_242 (O_242,N_4765,N_4737);
nand UO_243 (O_243,N_4698,N_4882);
or UO_244 (O_244,N_4575,N_4784);
or UO_245 (O_245,N_4593,N_4842);
or UO_246 (O_246,N_4912,N_4596);
xnor UO_247 (O_247,N_4697,N_4948);
and UO_248 (O_248,N_4814,N_4868);
or UO_249 (O_249,N_4556,N_4854);
nor UO_250 (O_250,N_4841,N_4603);
nor UO_251 (O_251,N_4641,N_4752);
nor UO_252 (O_252,N_4806,N_4559);
and UO_253 (O_253,N_4519,N_4829);
nand UO_254 (O_254,N_4753,N_4675);
and UO_255 (O_255,N_4558,N_4572);
nand UO_256 (O_256,N_4565,N_4895);
or UO_257 (O_257,N_4834,N_4977);
nor UO_258 (O_258,N_4656,N_4672);
nor UO_259 (O_259,N_4872,N_4874);
and UO_260 (O_260,N_4555,N_4735);
nor UO_261 (O_261,N_4807,N_4723);
and UO_262 (O_262,N_4759,N_4936);
nor UO_263 (O_263,N_4696,N_4869);
or UO_264 (O_264,N_4747,N_4920);
nor UO_265 (O_265,N_4865,N_4559);
or UO_266 (O_266,N_4576,N_4937);
and UO_267 (O_267,N_4570,N_4664);
nand UO_268 (O_268,N_4620,N_4788);
nand UO_269 (O_269,N_4757,N_4749);
or UO_270 (O_270,N_4612,N_4527);
and UO_271 (O_271,N_4960,N_4607);
and UO_272 (O_272,N_4687,N_4885);
and UO_273 (O_273,N_4667,N_4503);
nor UO_274 (O_274,N_4908,N_4598);
and UO_275 (O_275,N_4677,N_4857);
and UO_276 (O_276,N_4730,N_4920);
nor UO_277 (O_277,N_4890,N_4577);
and UO_278 (O_278,N_4911,N_4979);
and UO_279 (O_279,N_4746,N_4741);
and UO_280 (O_280,N_4545,N_4515);
nand UO_281 (O_281,N_4662,N_4844);
and UO_282 (O_282,N_4774,N_4921);
and UO_283 (O_283,N_4874,N_4952);
and UO_284 (O_284,N_4687,N_4518);
and UO_285 (O_285,N_4861,N_4689);
nor UO_286 (O_286,N_4567,N_4811);
or UO_287 (O_287,N_4834,N_4696);
nor UO_288 (O_288,N_4522,N_4980);
nand UO_289 (O_289,N_4717,N_4710);
or UO_290 (O_290,N_4879,N_4778);
or UO_291 (O_291,N_4811,N_4954);
and UO_292 (O_292,N_4788,N_4690);
nor UO_293 (O_293,N_4586,N_4788);
and UO_294 (O_294,N_4672,N_4508);
nand UO_295 (O_295,N_4948,N_4621);
or UO_296 (O_296,N_4838,N_4701);
xor UO_297 (O_297,N_4927,N_4537);
nand UO_298 (O_298,N_4834,N_4636);
and UO_299 (O_299,N_4811,N_4652);
and UO_300 (O_300,N_4511,N_4525);
and UO_301 (O_301,N_4551,N_4580);
and UO_302 (O_302,N_4520,N_4986);
nand UO_303 (O_303,N_4668,N_4739);
nand UO_304 (O_304,N_4993,N_4714);
and UO_305 (O_305,N_4789,N_4778);
nor UO_306 (O_306,N_4632,N_4592);
or UO_307 (O_307,N_4539,N_4518);
nand UO_308 (O_308,N_4500,N_4538);
nor UO_309 (O_309,N_4642,N_4845);
nand UO_310 (O_310,N_4577,N_4532);
nand UO_311 (O_311,N_4556,N_4639);
or UO_312 (O_312,N_4902,N_4550);
and UO_313 (O_313,N_4545,N_4762);
nor UO_314 (O_314,N_4562,N_4769);
and UO_315 (O_315,N_4794,N_4810);
and UO_316 (O_316,N_4932,N_4586);
or UO_317 (O_317,N_4725,N_4611);
and UO_318 (O_318,N_4670,N_4678);
and UO_319 (O_319,N_4883,N_4641);
or UO_320 (O_320,N_4531,N_4691);
or UO_321 (O_321,N_4762,N_4621);
nor UO_322 (O_322,N_4693,N_4978);
or UO_323 (O_323,N_4751,N_4795);
or UO_324 (O_324,N_4939,N_4916);
or UO_325 (O_325,N_4886,N_4635);
nand UO_326 (O_326,N_4762,N_4759);
and UO_327 (O_327,N_4687,N_4667);
or UO_328 (O_328,N_4600,N_4609);
nand UO_329 (O_329,N_4854,N_4934);
nand UO_330 (O_330,N_4665,N_4824);
nor UO_331 (O_331,N_4540,N_4688);
or UO_332 (O_332,N_4669,N_4829);
or UO_333 (O_333,N_4836,N_4560);
and UO_334 (O_334,N_4658,N_4745);
nor UO_335 (O_335,N_4595,N_4885);
nor UO_336 (O_336,N_4610,N_4668);
nor UO_337 (O_337,N_4857,N_4745);
nor UO_338 (O_338,N_4737,N_4539);
or UO_339 (O_339,N_4922,N_4900);
nand UO_340 (O_340,N_4821,N_4618);
or UO_341 (O_341,N_4515,N_4948);
nand UO_342 (O_342,N_4911,N_4904);
nor UO_343 (O_343,N_4931,N_4533);
nor UO_344 (O_344,N_4738,N_4533);
nor UO_345 (O_345,N_4802,N_4529);
or UO_346 (O_346,N_4603,N_4724);
and UO_347 (O_347,N_4866,N_4998);
or UO_348 (O_348,N_4831,N_4515);
nor UO_349 (O_349,N_4566,N_4804);
nor UO_350 (O_350,N_4629,N_4549);
nor UO_351 (O_351,N_4931,N_4638);
and UO_352 (O_352,N_4635,N_4571);
nand UO_353 (O_353,N_4764,N_4699);
or UO_354 (O_354,N_4998,N_4584);
nor UO_355 (O_355,N_4832,N_4969);
nor UO_356 (O_356,N_4815,N_4708);
and UO_357 (O_357,N_4955,N_4658);
nand UO_358 (O_358,N_4804,N_4987);
xor UO_359 (O_359,N_4789,N_4803);
nand UO_360 (O_360,N_4661,N_4535);
nand UO_361 (O_361,N_4926,N_4975);
nor UO_362 (O_362,N_4520,N_4749);
nand UO_363 (O_363,N_4764,N_4915);
or UO_364 (O_364,N_4979,N_4954);
nor UO_365 (O_365,N_4955,N_4654);
and UO_366 (O_366,N_4640,N_4522);
nand UO_367 (O_367,N_4911,N_4578);
nand UO_368 (O_368,N_4766,N_4527);
and UO_369 (O_369,N_4957,N_4718);
nand UO_370 (O_370,N_4575,N_4632);
nor UO_371 (O_371,N_4911,N_4680);
or UO_372 (O_372,N_4812,N_4573);
and UO_373 (O_373,N_4996,N_4768);
or UO_374 (O_374,N_4556,N_4888);
nand UO_375 (O_375,N_4954,N_4540);
nand UO_376 (O_376,N_4764,N_4560);
nor UO_377 (O_377,N_4852,N_4821);
nor UO_378 (O_378,N_4746,N_4961);
or UO_379 (O_379,N_4602,N_4988);
nand UO_380 (O_380,N_4772,N_4871);
and UO_381 (O_381,N_4917,N_4719);
nor UO_382 (O_382,N_4841,N_4761);
nor UO_383 (O_383,N_4811,N_4757);
or UO_384 (O_384,N_4815,N_4946);
nand UO_385 (O_385,N_4853,N_4533);
or UO_386 (O_386,N_4832,N_4809);
nand UO_387 (O_387,N_4651,N_4963);
or UO_388 (O_388,N_4529,N_4682);
or UO_389 (O_389,N_4750,N_4951);
nor UO_390 (O_390,N_4732,N_4795);
nand UO_391 (O_391,N_4658,N_4813);
and UO_392 (O_392,N_4783,N_4511);
nand UO_393 (O_393,N_4631,N_4585);
nor UO_394 (O_394,N_4707,N_4692);
or UO_395 (O_395,N_4585,N_4919);
nor UO_396 (O_396,N_4552,N_4813);
or UO_397 (O_397,N_4693,N_4807);
nand UO_398 (O_398,N_4583,N_4775);
nor UO_399 (O_399,N_4674,N_4591);
nor UO_400 (O_400,N_4566,N_4984);
nor UO_401 (O_401,N_4602,N_4832);
and UO_402 (O_402,N_4866,N_4980);
or UO_403 (O_403,N_4810,N_4523);
or UO_404 (O_404,N_4628,N_4831);
and UO_405 (O_405,N_4877,N_4815);
or UO_406 (O_406,N_4514,N_4832);
and UO_407 (O_407,N_4996,N_4947);
nand UO_408 (O_408,N_4504,N_4899);
nand UO_409 (O_409,N_4716,N_4975);
and UO_410 (O_410,N_4590,N_4613);
nor UO_411 (O_411,N_4836,N_4680);
or UO_412 (O_412,N_4584,N_4800);
nor UO_413 (O_413,N_4639,N_4631);
and UO_414 (O_414,N_4940,N_4622);
or UO_415 (O_415,N_4578,N_4907);
nand UO_416 (O_416,N_4858,N_4512);
nor UO_417 (O_417,N_4749,N_4962);
nor UO_418 (O_418,N_4792,N_4701);
nand UO_419 (O_419,N_4926,N_4848);
and UO_420 (O_420,N_4889,N_4551);
or UO_421 (O_421,N_4945,N_4812);
and UO_422 (O_422,N_4506,N_4872);
and UO_423 (O_423,N_4644,N_4736);
nand UO_424 (O_424,N_4569,N_4929);
nor UO_425 (O_425,N_4932,N_4590);
nand UO_426 (O_426,N_4862,N_4709);
and UO_427 (O_427,N_4814,N_4752);
nand UO_428 (O_428,N_4694,N_4919);
and UO_429 (O_429,N_4821,N_4590);
nor UO_430 (O_430,N_4972,N_4571);
nor UO_431 (O_431,N_4824,N_4708);
nor UO_432 (O_432,N_4565,N_4807);
nand UO_433 (O_433,N_4803,N_4526);
and UO_434 (O_434,N_4730,N_4700);
nor UO_435 (O_435,N_4630,N_4753);
nor UO_436 (O_436,N_4870,N_4590);
nand UO_437 (O_437,N_4788,N_4635);
nor UO_438 (O_438,N_4568,N_4941);
and UO_439 (O_439,N_4766,N_4573);
and UO_440 (O_440,N_4617,N_4512);
or UO_441 (O_441,N_4876,N_4593);
nor UO_442 (O_442,N_4918,N_4877);
or UO_443 (O_443,N_4597,N_4930);
nor UO_444 (O_444,N_4828,N_4583);
nor UO_445 (O_445,N_4705,N_4838);
and UO_446 (O_446,N_4805,N_4776);
and UO_447 (O_447,N_4711,N_4695);
nand UO_448 (O_448,N_4725,N_4980);
or UO_449 (O_449,N_4755,N_4738);
nand UO_450 (O_450,N_4645,N_4566);
or UO_451 (O_451,N_4876,N_4836);
nand UO_452 (O_452,N_4963,N_4731);
and UO_453 (O_453,N_4503,N_4565);
or UO_454 (O_454,N_4548,N_4526);
and UO_455 (O_455,N_4725,N_4584);
nand UO_456 (O_456,N_4673,N_4763);
nor UO_457 (O_457,N_4962,N_4756);
xor UO_458 (O_458,N_4984,N_4638);
and UO_459 (O_459,N_4979,N_4645);
nor UO_460 (O_460,N_4988,N_4955);
or UO_461 (O_461,N_4872,N_4550);
or UO_462 (O_462,N_4896,N_4639);
or UO_463 (O_463,N_4554,N_4803);
or UO_464 (O_464,N_4791,N_4975);
nor UO_465 (O_465,N_4731,N_4782);
nand UO_466 (O_466,N_4860,N_4801);
nor UO_467 (O_467,N_4887,N_4864);
nand UO_468 (O_468,N_4997,N_4757);
nor UO_469 (O_469,N_4951,N_4990);
or UO_470 (O_470,N_4687,N_4626);
nand UO_471 (O_471,N_4815,N_4747);
and UO_472 (O_472,N_4625,N_4603);
and UO_473 (O_473,N_4608,N_4769);
nand UO_474 (O_474,N_4691,N_4589);
or UO_475 (O_475,N_4572,N_4555);
or UO_476 (O_476,N_4646,N_4544);
or UO_477 (O_477,N_4549,N_4507);
nand UO_478 (O_478,N_4694,N_4549);
and UO_479 (O_479,N_4917,N_4981);
or UO_480 (O_480,N_4565,N_4594);
or UO_481 (O_481,N_4768,N_4574);
nor UO_482 (O_482,N_4806,N_4711);
nor UO_483 (O_483,N_4648,N_4633);
or UO_484 (O_484,N_4958,N_4584);
nor UO_485 (O_485,N_4905,N_4904);
nor UO_486 (O_486,N_4767,N_4710);
nand UO_487 (O_487,N_4813,N_4719);
nor UO_488 (O_488,N_4870,N_4676);
or UO_489 (O_489,N_4806,N_4959);
nor UO_490 (O_490,N_4821,N_4868);
or UO_491 (O_491,N_4522,N_4604);
nand UO_492 (O_492,N_4880,N_4891);
nor UO_493 (O_493,N_4639,N_4739);
nor UO_494 (O_494,N_4867,N_4912);
and UO_495 (O_495,N_4918,N_4971);
nor UO_496 (O_496,N_4618,N_4942);
or UO_497 (O_497,N_4704,N_4603);
and UO_498 (O_498,N_4625,N_4939);
nor UO_499 (O_499,N_4959,N_4506);
or UO_500 (O_500,N_4925,N_4774);
or UO_501 (O_501,N_4681,N_4688);
or UO_502 (O_502,N_4923,N_4622);
nand UO_503 (O_503,N_4657,N_4622);
xnor UO_504 (O_504,N_4962,N_4687);
nand UO_505 (O_505,N_4621,N_4966);
nor UO_506 (O_506,N_4793,N_4699);
or UO_507 (O_507,N_4524,N_4652);
and UO_508 (O_508,N_4688,N_4518);
or UO_509 (O_509,N_4744,N_4572);
and UO_510 (O_510,N_4716,N_4713);
or UO_511 (O_511,N_4826,N_4668);
nor UO_512 (O_512,N_4742,N_4839);
and UO_513 (O_513,N_4961,N_4757);
nand UO_514 (O_514,N_4641,N_4992);
xnor UO_515 (O_515,N_4539,N_4846);
nand UO_516 (O_516,N_4640,N_4731);
nor UO_517 (O_517,N_4899,N_4923);
nor UO_518 (O_518,N_4769,N_4529);
nor UO_519 (O_519,N_4893,N_4578);
or UO_520 (O_520,N_4739,N_4547);
and UO_521 (O_521,N_4984,N_4753);
nor UO_522 (O_522,N_4798,N_4943);
xor UO_523 (O_523,N_4969,N_4672);
nor UO_524 (O_524,N_4919,N_4969);
nand UO_525 (O_525,N_4515,N_4754);
nor UO_526 (O_526,N_4960,N_4985);
nor UO_527 (O_527,N_4840,N_4579);
or UO_528 (O_528,N_4828,N_4739);
and UO_529 (O_529,N_4850,N_4953);
nor UO_530 (O_530,N_4807,N_4846);
nand UO_531 (O_531,N_4763,N_4979);
and UO_532 (O_532,N_4665,N_4658);
nor UO_533 (O_533,N_4605,N_4627);
nor UO_534 (O_534,N_4888,N_4708);
or UO_535 (O_535,N_4787,N_4500);
or UO_536 (O_536,N_4908,N_4889);
nor UO_537 (O_537,N_4915,N_4736);
or UO_538 (O_538,N_4612,N_4867);
nor UO_539 (O_539,N_4839,N_4953);
and UO_540 (O_540,N_4825,N_4819);
and UO_541 (O_541,N_4783,N_4607);
or UO_542 (O_542,N_4685,N_4667);
nand UO_543 (O_543,N_4926,N_4846);
nor UO_544 (O_544,N_4617,N_4812);
nor UO_545 (O_545,N_4946,N_4874);
or UO_546 (O_546,N_4707,N_4954);
and UO_547 (O_547,N_4960,N_4630);
and UO_548 (O_548,N_4600,N_4733);
or UO_549 (O_549,N_4753,N_4912);
and UO_550 (O_550,N_4692,N_4662);
nand UO_551 (O_551,N_4587,N_4670);
nand UO_552 (O_552,N_4935,N_4943);
or UO_553 (O_553,N_4922,N_4923);
and UO_554 (O_554,N_4764,N_4660);
nor UO_555 (O_555,N_4630,N_4936);
nand UO_556 (O_556,N_4940,N_4582);
and UO_557 (O_557,N_4781,N_4972);
and UO_558 (O_558,N_4689,N_4616);
and UO_559 (O_559,N_4878,N_4572);
nor UO_560 (O_560,N_4682,N_4822);
and UO_561 (O_561,N_4849,N_4575);
and UO_562 (O_562,N_4769,N_4572);
and UO_563 (O_563,N_4659,N_4664);
or UO_564 (O_564,N_4856,N_4736);
nor UO_565 (O_565,N_4704,N_4617);
nor UO_566 (O_566,N_4891,N_4532);
and UO_567 (O_567,N_4813,N_4735);
or UO_568 (O_568,N_4960,N_4969);
nor UO_569 (O_569,N_4956,N_4574);
nor UO_570 (O_570,N_4971,N_4523);
and UO_571 (O_571,N_4987,N_4762);
and UO_572 (O_572,N_4662,N_4727);
xnor UO_573 (O_573,N_4711,N_4702);
nand UO_574 (O_574,N_4732,N_4990);
or UO_575 (O_575,N_4814,N_4633);
and UO_576 (O_576,N_4948,N_4703);
and UO_577 (O_577,N_4666,N_4981);
and UO_578 (O_578,N_4557,N_4502);
nand UO_579 (O_579,N_4525,N_4933);
nor UO_580 (O_580,N_4638,N_4843);
nand UO_581 (O_581,N_4667,N_4878);
and UO_582 (O_582,N_4955,N_4799);
nor UO_583 (O_583,N_4617,N_4578);
nand UO_584 (O_584,N_4517,N_4577);
and UO_585 (O_585,N_4903,N_4582);
or UO_586 (O_586,N_4990,N_4694);
nor UO_587 (O_587,N_4961,N_4978);
nor UO_588 (O_588,N_4556,N_4719);
or UO_589 (O_589,N_4636,N_4886);
nand UO_590 (O_590,N_4882,N_4649);
or UO_591 (O_591,N_4783,N_4609);
and UO_592 (O_592,N_4651,N_4520);
nand UO_593 (O_593,N_4989,N_4608);
nor UO_594 (O_594,N_4975,N_4535);
nor UO_595 (O_595,N_4889,N_4547);
nor UO_596 (O_596,N_4869,N_4787);
or UO_597 (O_597,N_4950,N_4802);
xnor UO_598 (O_598,N_4803,N_4600);
nor UO_599 (O_599,N_4784,N_4827);
nand UO_600 (O_600,N_4841,N_4847);
xor UO_601 (O_601,N_4821,N_4804);
xnor UO_602 (O_602,N_4588,N_4612);
xor UO_603 (O_603,N_4540,N_4918);
nor UO_604 (O_604,N_4545,N_4747);
and UO_605 (O_605,N_4774,N_4887);
or UO_606 (O_606,N_4876,N_4943);
and UO_607 (O_607,N_4954,N_4953);
nor UO_608 (O_608,N_4633,N_4976);
and UO_609 (O_609,N_4938,N_4821);
and UO_610 (O_610,N_4575,N_4962);
nor UO_611 (O_611,N_4604,N_4956);
or UO_612 (O_612,N_4664,N_4837);
nand UO_613 (O_613,N_4648,N_4780);
and UO_614 (O_614,N_4637,N_4942);
or UO_615 (O_615,N_4971,N_4829);
and UO_616 (O_616,N_4690,N_4581);
nand UO_617 (O_617,N_4821,N_4784);
xor UO_618 (O_618,N_4676,N_4689);
and UO_619 (O_619,N_4708,N_4532);
nand UO_620 (O_620,N_4551,N_4755);
and UO_621 (O_621,N_4658,N_4787);
xor UO_622 (O_622,N_4584,N_4735);
or UO_623 (O_623,N_4937,N_4718);
and UO_624 (O_624,N_4621,N_4954);
nand UO_625 (O_625,N_4812,N_4748);
nor UO_626 (O_626,N_4667,N_4544);
nor UO_627 (O_627,N_4546,N_4592);
nor UO_628 (O_628,N_4593,N_4589);
and UO_629 (O_629,N_4627,N_4795);
nor UO_630 (O_630,N_4903,N_4895);
nor UO_631 (O_631,N_4550,N_4755);
xor UO_632 (O_632,N_4522,N_4932);
and UO_633 (O_633,N_4877,N_4813);
and UO_634 (O_634,N_4919,N_4957);
or UO_635 (O_635,N_4698,N_4899);
nor UO_636 (O_636,N_4793,N_4582);
nor UO_637 (O_637,N_4961,N_4970);
nand UO_638 (O_638,N_4964,N_4739);
or UO_639 (O_639,N_4846,N_4985);
nor UO_640 (O_640,N_4541,N_4659);
or UO_641 (O_641,N_4969,N_4653);
and UO_642 (O_642,N_4740,N_4755);
and UO_643 (O_643,N_4589,N_4601);
or UO_644 (O_644,N_4565,N_4544);
xnor UO_645 (O_645,N_4573,N_4966);
nor UO_646 (O_646,N_4950,N_4992);
or UO_647 (O_647,N_4841,N_4881);
and UO_648 (O_648,N_4861,N_4673);
or UO_649 (O_649,N_4988,N_4658);
or UO_650 (O_650,N_4993,N_4797);
nand UO_651 (O_651,N_4988,N_4540);
or UO_652 (O_652,N_4767,N_4961);
nor UO_653 (O_653,N_4626,N_4982);
and UO_654 (O_654,N_4598,N_4586);
and UO_655 (O_655,N_4786,N_4749);
nor UO_656 (O_656,N_4928,N_4919);
nand UO_657 (O_657,N_4585,N_4511);
or UO_658 (O_658,N_4894,N_4592);
nand UO_659 (O_659,N_4797,N_4759);
nand UO_660 (O_660,N_4512,N_4669);
or UO_661 (O_661,N_4668,N_4856);
or UO_662 (O_662,N_4946,N_4614);
or UO_663 (O_663,N_4605,N_4586);
nand UO_664 (O_664,N_4923,N_4576);
or UO_665 (O_665,N_4724,N_4800);
or UO_666 (O_666,N_4720,N_4574);
and UO_667 (O_667,N_4597,N_4545);
nor UO_668 (O_668,N_4506,N_4936);
nand UO_669 (O_669,N_4621,N_4823);
and UO_670 (O_670,N_4978,N_4722);
or UO_671 (O_671,N_4977,N_4738);
nand UO_672 (O_672,N_4839,N_4956);
or UO_673 (O_673,N_4707,N_4628);
or UO_674 (O_674,N_4662,N_4954);
or UO_675 (O_675,N_4596,N_4530);
nor UO_676 (O_676,N_4652,N_4563);
nand UO_677 (O_677,N_4604,N_4982);
or UO_678 (O_678,N_4616,N_4944);
nand UO_679 (O_679,N_4994,N_4811);
and UO_680 (O_680,N_4953,N_4917);
nand UO_681 (O_681,N_4642,N_4866);
or UO_682 (O_682,N_4824,N_4751);
and UO_683 (O_683,N_4958,N_4989);
and UO_684 (O_684,N_4937,N_4524);
nand UO_685 (O_685,N_4526,N_4758);
and UO_686 (O_686,N_4583,N_4809);
xnor UO_687 (O_687,N_4923,N_4893);
nor UO_688 (O_688,N_4693,N_4670);
and UO_689 (O_689,N_4947,N_4716);
or UO_690 (O_690,N_4714,N_4681);
nor UO_691 (O_691,N_4568,N_4892);
and UO_692 (O_692,N_4943,N_4545);
and UO_693 (O_693,N_4973,N_4599);
nand UO_694 (O_694,N_4990,N_4711);
or UO_695 (O_695,N_4513,N_4685);
nand UO_696 (O_696,N_4505,N_4554);
and UO_697 (O_697,N_4949,N_4519);
or UO_698 (O_698,N_4785,N_4955);
and UO_699 (O_699,N_4925,N_4585);
and UO_700 (O_700,N_4926,N_4845);
and UO_701 (O_701,N_4982,N_4612);
nand UO_702 (O_702,N_4649,N_4807);
xor UO_703 (O_703,N_4897,N_4930);
and UO_704 (O_704,N_4709,N_4523);
or UO_705 (O_705,N_4691,N_4915);
and UO_706 (O_706,N_4733,N_4571);
or UO_707 (O_707,N_4676,N_4835);
and UO_708 (O_708,N_4718,N_4880);
or UO_709 (O_709,N_4941,N_4799);
nor UO_710 (O_710,N_4502,N_4561);
nand UO_711 (O_711,N_4677,N_4705);
nor UO_712 (O_712,N_4908,N_4976);
and UO_713 (O_713,N_4676,N_4534);
nand UO_714 (O_714,N_4876,N_4865);
nor UO_715 (O_715,N_4745,N_4759);
nand UO_716 (O_716,N_4581,N_4714);
nor UO_717 (O_717,N_4561,N_4837);
nand UO_718 (O_718,N_4773,N_4693);
or UO_719 (O_719,N_4859,N_4651);
nor UO_720 (O_720,N_4755,N_4586);
and UO_721 (O_721,N_4947,N_4686);
and UO_722 (O_722,N_4844,N_4736);
and UO_723 (O_723,N_4879,N_4927);
and UO_724 (O_724,N_4700,N_4945);
and UO_725 (O_725,N_4915,N_4918);
nor UO_726 (O_726,N_4579,N_4908);
or UO_727 (O_727,N_4780,N_4501);
and UO_728 (O_728,N_4684,N_4699);
or UO_729 (O_729,N_4582,N_4539);
nor UO_730 (O_730,N_4647,N_4717);
nor UO_731 (O_731,N_4773,N_4896);
nand UO_732 (O_732,N_4997,N_4765);
nor UO_733 (O_733,N_4639,N_4679);
nand UO_734 (O_734,N_4610,N_4615);
nand UO_735 (O_735,N_4744,N_4726);
and UO_736 (O_736,N_4797,N_4730);
and UO_737 (O_737,N_4843,N_4565);
or UO_738 (O_738,N_4865,N_4617);
nor UO_739 (O_739,N_4986,N_4589);
or UO_740 (O_740,N_4836,N_4851);
nand UO_741 (O_741,N_4654,N_4879);
and UO_742 (O_742,N_4784,N_4605);
or UO_743 (O_743,N_4837,N_4879);
xor UO_744 (O_744,N_4656,N_4524);
nor UO_745 (O_745,N_4742,N_4613);
or UO_746 (O_746,N_4781,N_4730);
or UO_747 (O_747,N_4862,N_4611);
and UO_748 (O_748,N_4772,N_4558);
xor UO_749 (O_749,N_4748,N_4697);
or UO_750 (O_750,N_4776,N_4822);
nand UO_751 (O_751,N_4810,N_4620);
nor UO_752 (O_752,N_4986,N_4640);
nor UO_753 (O_753,N_4670,N_4561);
or UO_754 (O_754,N_4669,N_4508);
nor UO_755 (O_755,N_4640,N_4746);
nand UO_756 (O_756,N_4796,N_4885);
nand UO_757 (O_757,N_4737,N_4510);
or UO_758 (O_758,N_4917,N_4890);
and UO_759 (O_759,N_4859,N_4780);
and UO_760 (O_760,N_4893,N_4500);
nand UO_761 (O_761,N_4554,N_4606);
nand UO_762 (O_762,N_4712,N_4977);
nor UO_763 (O_763,N_4898,N_4571);
nor UO_764 (O_764,N_4698,N_4616);
nand UO_765 (O_765,N_4990,N_4724);
or UO_766 (O_766,N_4619,N_4813);
or UO_767 (O_767,N_4881,N_4711);
nor UO_768 (O_768,N_4527,N_4571);
nor UO_769 (O_769,N_4520,N_4689);
nor UO_770 (O_770,N_4586,N_4528);
or UO_771 (O_771,N_4757,N_4684);
and UO_772 (O_772,N_4736,N_4563);
or UO_773 (O_773,N_4529,N_4839);
and UO_774 (O_774,N_4754,N_4716);
and UO_775 (O_775,N_4941,N_4883);
nand UO_776 (O_776,N_4730,N_4836);
nand UO_777 (O_777,N_4890,N_4940);
nand UO_778 (O_778,N_4726,N_4979);
or UO_779 (O_779,N_4745,N_4829);
and UO_780 (O_780,N_4830,N_4668);
xnor UO_781 (O_781,N_4633,N_4912);
nor UO_782 (O_782,N_4855,N_4748);
nor UO_783 (O_783,N_4782,N_4905);
or UO_784 (O_784,N_4921,N_4627);
nand UO_785 (O_785,N_4733,N_4543);
nand UO_786 (O_786,N_4635,N_4512);
nand UO_787 (O_787,N_4504,N_4855);
and UO_788 (O_788,N_4987,N_4652);
or UO_789 (O_789,N_4691,N_4904);
and UO_790 (O_790,N_4919,N_4520);
or UO_791 (O_791,N_4653,N_4917);
nand UO_792 (O_792,N_4689,N_4589);
nand UO_793 (O_793,N_4591,N_4792);
and UO_794 (O_794,N_4857,N_4505);
and UO_795 (O_795,N_4789,N_4704);
and UO_796 (O_796,N_4917,N_4544);
nand UO_797 (O_797,N_4653,N_4771);
nor UO_798 (O_798,N_4533,N_4855);
and UO_799 (O_799,N_4810,N_4743);
or UO_800 (O_800,N_4565,N_4903);
nor UO_801 (O_801,N_4737,N_4557);
nand UO_802 (O_802,N_4576,N_4989);
nand UO_803 (O_803,N_4625,N_4770);
nor UO_804 (O_804,N_4747,N_4610);
and UO_805 (O_805,N_4605,N_4915);
nor UO_806 (O_806,N_4791,N_4758);
or UO_807 (O_807,N_4546,N_4794);
or UO_808 (O_808,N_4605,N_4869);
and UO_809 (O_809,N_4841,N_4579);
and UO_810 (O_810,N_4764,N_4690);
nor UO_811 (O_811,N_4727,N_4868);
or UO_812 (O_812,N_4813,N_4923);
nor UO_813 (O_813,N_4641,N_4507);
nor UO_814 (O_814,N_4941,N_4622);
nor UO_815 (O_815,N_4634,N_4601);
nand UO_816 (O_816,N_4829,N_4815);
nor UO_817 (O_817,N_4515,N_4943);
nor UO_818 (O_818,N_4844,N_4890);
and UO_819 (O_819,N_4572,N_4898);
and UO_820 (O_820,N_4926,N_4601);
nor UO_821 (O_821,N_4805,N_4536);
or UO_822 (O_822,N_4566,N_4598);
nor UO_823 (O_823,N_4778,N_4777);
and UO_824 (O_824,N_4854,N_4693);
and UO_825 (O_825,N_4725,N_4577);
or UO_826 (O_826,N_4900,N_4980);
nand UO_827 (O_827,N_4875,N_4678);
and UO_828 (O_828,N_4952,N_4575);
nand UO_829 (O_829,N_4935,N_4791);
xor UO_830 (O_830,N_4992,N_4704);
nand UO_831 (O_831,N_4856,N_4547);
nand UO_832 (O_832,N_4910,N_4604);
xnor UO_833 (O_833,N_4650,N_4785);
nand UO_834 (O_834,N_4586,N_4769);
nor UO_835 (O_835,N_4749,N_4880);
nand UO_836 (O_836,N_4822,N_4544);
nor UO_837 (O_837,N_4703,N_4578);
and UO_838 (O_838,N_4675,N_4810);
nor UO_839 (O_839,N_4891,N_4951);
nand UO_840 (O_840,N_4836,N_4733);
xnor UO_841 (O_841,N_4676,N_4577);
nor UO_842 (O_842,N_4507,N_4589);
nand UO_843 (O_843,N_4610,N_4538);
and UO_844 (O_844,N_4715,N_4819);
nor UO_845 (O_845,N_4620,N_4877);
nor UO_846 (O_846,N_4596,N_4994);
nor UO_847 (O_847,N_4726,N_4713);
nand UO_848 (O_848,N_4767,N_4545);
nand UO_849 (O_849,N_4583,N_4547);
nand UO_850 (O_850,N_4925,N_4858);
or UO_851 (O_851,N_4844,N_4550);
nand UO_852 (O_852,N_4987,N_4740);
nand UO_853 (O_853,N_4874,N_4884);
and UO_854 (O_854,N_4886,N_4880);
nand UO_855 (O_855,N_4531,N_4753);
or UO_856 (O_856,N_4929,N_4506);
nand UO_857 (O_857,N_4718,N_4762);
nor UO_858 (O_858,N_4860,N_4564);
nand UO_859 (O_859,N_4949,N_4743);
nor UO_860 (O_860,N_4638,N_4538);
and UO_861 (O_861,N_4828,N_4860);
or UO_862 (O_862,N_4746,N_4698);
nor UO_863 (O_863,N_4614,N_4935);
or UO_864 (O_864,N_4605,N_4530);
nor UO_865 (O_865,N_4812,N_4749);
nor UO_866 (O_866,N_4943,N_4857);
nor UO_867 (O_867,N_4585,N_4714);
or UO_868 (O_868,N_4722,N_4911);
nand UO_869 (O_869,N_4774,N_4915);
nor UO_870 (O_870,N_4675,N_4574);
and UO_871 (O_871,N_4930,N_4715);
nor UO_872 (O_872,N_4935,N_4525);
nand UO_873 (O_873,N_4710,N_4948);
and UO_874 (O_874,N_4630,N_4675);
nor UO_875 (O_875,N_4889,N_4534);
nand UO_876 (O_876,N_4947,N_4887);
and UO_877 (O_877,N_4897,N_4744);
nand UO_878 (O_878,N_4768,N_4978);
nor UO_879 (O_879,N_4681,N_4543);
nand UO_880 (O_880,N_4880,N_4712);
or UO_881 (O_881,N_4743,N_4883);
nor UO_882 (O_882,N_4753,N_4977);
nor UO_883 (O_883,N_4778,N_4584);
nand UO_884 (O_884,N_4623,N_4635);
and UO_885 (O_885,N_4613,N_4503);
and UO_886 (O_886,N_4738,N_4962);
or UO_887 (O_887,N_4552,N_4632);
or UO_888 (O_888,N_4879,N_4810);
nand UO_889 (O_889,N_4997,N_4840);
and UO_890 (O_890,N_4761,N_4517);
nand UO_891 (O_891,N_4739,N_4830);
nand UO_892 (O_892,N_4927,N_4961);
nor UO_893 (O_893,N_4703,N_4987);
nor UO_894 (O_894,N_4734,N_4706);
nand UO_895 (O_895,N_4509,N_4901);
and UO_896 (O_896,N_4686,N_4971);
and UO_897 (O_897,N_4612,N_4742);
nand UO_898 (O_898,N_4571,N_4584);
nor UO_899 (O_899,N_4593,N_4970);
and UO_900 (O_900,N_4989,N_4892);
nor UO_901 (O_901,N_4883,N_4643);
and UO_902 (O_902,N_4894,N_4617);
nand UO_903 (O_903,N_4853,N_4980);
nor UO_904 (O_904,N_4789,N_4538);
nor UO_905 (O_905,N_4938,N_4885);
nor UO_906 (O_906,N_4801,N_4586);
and UO_907 (O_907,N_4805,N_4804);
nor UO_908 (O_908,N_4689,N_4581);
and UO_909 (O_909,N_4762,N_4649);
xnor UO_910 (O_910,N_4579,N_4809);
and UO_911 (O_911,N_4915,N_4583);
and UO_912 (O_912,N_4937,N_4765);
nor UO_913 (O_913,N_4627,N_4597);
nor UO_914 (O_914,N_4960,N_4926);
or UO_915 (O_915,N_4704,N_4995);
or UO_916 (O_916,N_4864,N_4815);
nor UO_917 (O_917,N_4744,N_4753);
and UO_918 (O_918,N_4796,N_4988);
or UO_919 (O_919,N_4799,N_4986);
nand UO_920 (O_920,N_4776,N_4893);
nor UO_921 (O_921,N_4782,N_4981);
nand UO_922 (O_922,N_4698,N_4750);
nor UO_923 (O_923,N_4644,N_4898);
nand UO_924 (O_924,N_4605,N_4735);
or UO_925 (O_925,N_4819,N_4980);
nor UO_926 (O_926,N_4584,N_4835);
and UO_927 (O_927,N_4772,N_4795);
xor UO_928 (O_928,N_4878,N_4974);
nor UO_929 (O_929,N_4661,N_4651);
and UO_930 (O_930,N_4747,N_4687);
and UO_931 (O_931,N_4721,N_4776);
or UO_932 (O_932,N_4574,N_4912);
or UO_933 (O_933,N_4756,N_4537);
nand UO_934 (O_934,N_4750,N_4629);
nor UO_935 (O_935,N_4795,N_4944);
nor UO_936 (O_936,N_4653,N_4626);
or UO_937 (O_937,N_4505,N_4874);
and UO_938 (O_938,N_4660,N_4900);
nor UO_939 (O_939,N_4584,N_4908);
or UO_940 (O_940,N_4786,N_4537);
or UO_941 (O_941,N_4643,N_4510);
nor UO_942 (O_942,N_4895,N_4552);
and UO_943 (O_943,N_4702,N_4779);
nor UO_944 (O_944,N_4683,N_4515);
or UO_945 (O_945,N_4941,N_4519);
xnor UO_946 (O_946,N_4791,N_4552);
nor UO_947 (O_947,N_4812,N_4721);
nand UO_948 (O_948,N_4599,N_4758);
or UO_949 (O_949,N_4845,N_4548);
and UO_950 (O_950,N_4654,N_4614);
and UO_951 (O_951,N_4873,N_4997);
or UO_952 (O_952,N_4545,N_4578);
nor UO_953 (O_953,N_4634,N_4587);
nand UO_954 (O_954,N_4676,N_4604);
nand UO_955 (O_955,N_4543,N_4833);
nand UO_956 (O_956,N_4547,N_4717);
or UO_957 (O_957,N_4793,N_4567);
nand UO_958 (O_958,N_4630,N_4662);
nor UO_959 (O_959,N_4795,N_4635);
and UO_960 (O_960,N_4520,N_4803);
nand UO_961 (O_961,N_4518,N_4684);
and UO_962 (O_962,N_4594,N_4832);
nor UO_963 (O_963,N_4618,N_4860);
or UO_964 (O_964,N_4512,N_4587);
nand UO_965 (O_965,N_4977,N_4657);
nor UO_966 (O_966,N_4644,N_4771);
nor UO_967 (O_967,N_4624,N_4745);
and UO_968 (O_968,N_4748,N_4595);
nand UO_969 (O_969,N_4885,N_4509);
nor UO_970 (O_970,N_4795,N_4797);
or UO_971 (O_971,N_4773,N_4652);
nor UO_972 (O_972,N_4657,N_4818);
nand UO_973 (O_973,N_4958,N_4723);
nand UO_974 (O_974,N_4518,N_4605);
or UO_975 (O_975,N_4922,N_4859);
or UO_976 (O_976,N_4831,N_4909);
or UO_977 (O_977,N_4817,N_4871);
and UO_978 (O_978,N_4804,N_4616);
and UO_979 (O_979,N_4676,N_4763);
and UO_980 (O_980,N_4987,N_4926);
or UO_981 (O_981,N_4500,N_4646);
or UO_982 (O_982,N_4593,N_4639);
nor UO_983 (O_983,N_4692,N_4629);
xnor UO_984 (O_984,N_4989,N_4865);
nand UO_985 (O_985,N_4981,N_4767);
or UO_986 (O_986,N_4919,N_4896);
nand UO_987 (O_987,N_4777,N_4717);
or UO_988 (O_988,N_4542,N_4988);
nand UO_989 (O_989,N_4910,N_4696);
nor UO_990 (O_990,N_4815,N_4980);
or UO_991 (O_991,N_4921,N_4857);
nor UO_992 (O_992,N_4874,N_4657);
nor UO_993 (O_993,N_4618,N_4995);
or UO_994 (O_994,N_4866,N_4743);
nor UO_995 (O_995,N_4665,N_4620);
or UO_996 (O_996,N_4947,N_4671);
nor UO_997 (O_997,N_4638,N_4894);
or UO_998 (O_998,N_4882,N_4611);
nand UO_999 (O_999,N_4532,N_4778);
endmodule