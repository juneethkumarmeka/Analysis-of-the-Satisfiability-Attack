module basic_1500_15000_2000_120_levels_10xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
and U0 (N_0,In_1122,In_693);
nand U1 (N_1,In_49,In_612);
nand U2 (N_2,In_1253,In_391);
and U3 (N_3,In_665,In_1012);
xor U4 (N_4,In_491,In_268);
nor U5 (N_5,In_666,In_1164);
or U6 (N_6,In_1248,In_897);
nand U7 (N_7,In_976,In_1098);
or U8 (N_8,In_914,In_1343);
or U9 (N_9,In_54,In_427);
or U10 (N_10,In_1230,In_1147);
nor U11 (N_11,In_544,In_98);
xnor U12 (N_12,In_1282,In_1156);
nand U13 (N_13,In_842,In_15);
xnor U14 (N_14,In_219,In_63);
nand U15 (N_15,In_988,In_1371);
xor U16 (N_16,In_920,In_1200);
xnor U17 (N_17,In_1235,In_1417);
xnor U18 (N_18,In_1468,In_3);
xor U19 (N_19,In_406,In_1024);
nand U20 (N_20,In_404,In_849);
xnor U21 (N_21,In_1065,In_280);
nand U22 (N_22,In_1418,In_600);
or U23 (N_23,In_743,In_683);
or U24 (N_24,In_1390,In_1081);
xor U25 (N_25,In_763,In_933);
nor U26 (N_26,In_486,In_561);
or U27 (N_27,In_941,In_128);
xor U28 (N_28,In_399,In_1222);
and U29 (N_29,In_911,In_131);
nand U30 (N_30,In_862,In_791);
nand U31 (N_31,In_1313,In_354);
or U32 (N_32,In_1219,In_363);
nor U33 (N_33,In_374,In_783);
xnor U34 (N_34,In_906,In_333);
or U35 (N_35,In_292,In_1163);
and U36 (N_36,In_411,In_1119);
nand U37 (N_37,In_1168,In_325);
nor U38 (N_38,In_850,In_1158);
or U39 (N_39,In_1432,In_1456);
and U40 (N_40,In_1378,In_364);
nor U41 (N_41,In_702,In_787);
nor U42 (N_42,In_59,In_1057);
nand U43 (N_43,In_956,In_990);
or U44 (N_44,In_1427,In_921);
nand U45 (N_45,In_378,In_1127);
nand U46 (N_46,In_1047,In_690);
xnor U47 (N_47,In_1326,In_1197);
nand U48 (N_48,In_593,In_860);
or U49 (N_49,In_569,In_1305);
or U50 (N_50,In_422,In_242);
and U51 (N_51,In_64,In_963);
or U52 (N_52,In_197,In_403);
or U53 (N_53,In_440,In_1380);
xnor U54 (N_54,In_1388,In_1068);
xnor U55 (N_55,In_800,In_1079);
and U56 (N_56,In_28,In_603);
nor U57 (N_57,In_206,In_1279);
xnor U58 (N_58,In_24,In_839);
and U59 (N_59,In_201,In_540);
nor U60 (N_60,In_1171,In_939);
xor U61 (N_61,In_53,In_574);
nand U62 (N_62,In_589,In_821);
and U63 (N_63,In_742,In_1341);
nand U64 (N_64,In_151,In_177);
or U65 (N_65,In_519,In_913);
or U66 (N_66,In_1143,In_1294);
xor U67 (N_67,In_1394,In_298);
nand U68 (N_68,In_306,In_648);
and U69 (N_69,In_541,In_507);
nand U70 (N_70,In_459,In_892);
nand U71 (N_71,In_296,In_694);
xor U72 (N_72,In_1300,In_919);
or U73 (N_73,In_506,In_801);
nand U74 (N_74,In_426,In_1061);
xor U75 (N_75,In_522,In_577);
nor U76 (N_76,In_453,In_29);
xor U77 (N_77,In_408,In_863);
and U78 (N_78,In_543,In_464);
nand U79 (N_79,In_1392,In_996);
or U80 (N_80,In_969,In_1196);
or U81 (N_81,In_557,In_586);
nor U82 (N_82,In_1094,In_218);
nor U83 (N_83,In_657,In_444);
and U84 (N_84,In_1382,In_161);
nor U85 (N_85,In_931,In_164);
nor U86 (N_86,In_1285,In_1215);
nand U87 (N_87,In_527,In_1090);
and U88 (N_88,In_932,In_1130);
or U89 (N_89,In_181,In_594);
nor U90 (N_90,In_1223,In_212);
or U91 (N_91,In_1312,In_1302);
nand U92 (N_92,In_184,In_869);
or U93 (N_93,In_1157,In_1084);
xnor U94 (N_94,In_509,In_592);
xnor U95 (N_95,In_903,In_235);
xnor U96 (N_96,In_46,In_790);
nor U97 (N_97,In_33,In_1103);
nand U98 (N_98,In_1410,In_439);
or U99 (N_99,In_1177,In_741);
and U100 (N_100,In_1039,In_752);
xnor U101 (N_101,In_182,In_1421);
and U102 (N_102,In_595,In_767);
xor U103 (N_103,In_189,In_393);
nand U104 (N_104,In_895,In_409);
xnor U105 (N_105,In_872,In_588);
or U106 (N_106,In_667,In_1110);
xnor U107 (N_107,In_677,In_283);
nand U108 (N_108,In_1365,In_311);
nand U109 (N_109,In_1487,In_671);
or U110 (N_110,In_717,In_838);
xnor U111 (N_111,In_1311,In_203);
nand U112 (N_112,In_780,In_136);
and U113 (N_113,In_1250,In_1029);
or U114 (N_114,In_596,In_659);
xor U115 (N_115,In_301,In_120);
nor U116 (N_116,In_1465,In_1121);
and U117 (N_117,In_1320,In_13);
xnor U118 (N_118,In_277,In_1070);
nor U119 (N_119,In_97,In_599);
xnor U120 (N_120,In_273,In_315);
nand U121 (N_121,In_1287,In_836);
nand U122 (N_122,In_539,In_1357);
nor U123 (N_123,In_214,In_1035);
xor U124 (N_124,In_113,In_1236);
and U125 (N_125,In_1139,In_611);
and U126 (N_126,In_1495,In_972);
and U127 (N_127,In_178,In_725);
nand U128 (N_128,In_940,In_615);
nand U129 (N_129,In_997,In_629);
or U130 (N_130,In_468,In_951);
xor U131 (N_131,In_1149,In_443);
xor U132 (N_132,In_738,In_649);
nand U133 (N_133,N_23,In_1450);
and U134 (N_134,In_142,In_1071);
xnor U135 (N_135,In_815,In_67);
nand U136 (N_136,In_760,In_1315);
nor U137 (N_137,N_58,In_1292);
xor U138 (N_138,In_620,In_999);
nor U139 (N_139,In_331,In_1181);
or U140 (N_140,In_202,In_1009);
or U141 (N_141,In_882,In_1339);
xnor U142 (N_142,In_327,In_977);
or U143 (N_143,In_25,In_43);
and U144 (N_144,In_533,In_936);
nand U145 (N_145,In_32,In_1075);
or U146 (N_146,In_446,In_910);
or U147 (N_147,In_1144,In_180);
nand U148 (N_148,In_636,In_537);
and U149 (N_149,In_1281,In_1267);
nand U150 (N_150,In_187,In_697);
nor U151 (N_151,In_1490,In_482);
xor U152 (N_152,In_1379,In_476);
xor U153 (N_153,In_496,In_163);
nand U154 (N_154,In_449,In_153);
or U155 (N_155,N_31,In_1364);
or U156 (N_156,In_245,In_158);
xor U157 (N_157,In_748,In_9);
nor U158 (N_158,In_72,In_89);
xor U159 (N_159,In_1325,In_80);
xor U160 (N_160,In_822,In_835);
xor U161 (N_161,In_874,In_433);
or U162 (N_162,In_1272,In_1111);
nand U163 (N_163,In_1193,In_40);
nor U164 (N_164,In_204,In_1480);
nand U165 (N_165,N_24,In_704);
or U166 (N_166,In_118,In_719);
nand U167 (N_167,In_266,In_1097);
nor U168 (N_168,In_979,In_1474);
nor U169 (N_169,In_103,In_1);
or U170 (N_170,In_190,In_485);
and U171 (N_171,In_1423,In_547);
xnor U172 (N_172,In_891,In_851);
and U173 (N_173,In_1172,In_907);
nor U174 (N_174,N_101,In_101);
nor U175 (N_175,In_1195,In_339);
and U176 (N_176,In_1454,In_1360);
nor U177 (N_177,In_299,In_431);
nand U178 (N_178,In_176,In_241);
nor U179 (N_179,In_803,In_1316);
nand U180 (N_180,In_361,In_623);
nand U181 (N_181,In_1477,In_385);
xnor U182 (N_182,In_1232,In_768);
or U183 (N_183,In_844,In_1445);
and U184 (N_184,In_1411,In_1078);
or U185 (N_185,In_259,N_8);
or U186 (N_186,In_282,In_1214);
or U187 (N_187,In_1386,In_493);
xnor U188 (N_188,In_21,In_1413);
or U189 (N_189,In_428,In_148);
nor U190 (N_190,In_806,In_1132);
or U191 (N_191,In_162,In_1102);
and U192 (N_192,In_1161,In_384);
xnor U193 (N_193,N_18,In_645);
xnor U194 (N_194,In_814,In_929);
nor U195 (N_195,In_1488,In_1489);
or U196 (N_196,In_346,In_157);
nand U197 (N_197,In_832,N_107);
nand U198 (N_198,In_917,In_1082);
nand U199 (N_199,In_69,In_111);
nor U200 (N_200,In_669,In_55);
nand U201 (N_201,N_10,In_528);
nand U202 (N_202,In_542,In_1317);
and U203 (N_203,In_634,N_56);
and U204 (N_204,In_1131,In_194);
or U205 (N_205,In_1092,In_149);
nor U206 (N_206,In_451,In_232);
nor U207 (N_207,In_1249,N_118);
xnor U208 (N_208,In_878,In_662);
and U209 (N_209,In_966,In_968);
nand U210 (N_210,N_100,In_223);
and U211 (N_211,In_34,In_1055);
nor U212 (N_212,In_766,N_112);
and U213 (N_213,In_1023,In_1008);
xnor U214 (N_214,In_44,N_52);
xor U215 (N_215,In_978,N_86);
nand U216 (N_216,In_258,In_434);
xnor U217 (N_217,In_646,In_1472);
nand U218 (N_218,In_198,In_1176);
and U219 (N_219,In_174,In_837);
or U220 (N_220,In_711,In_1041);
nor U221 (N_221,In_126,In_856);
nor U222 (N_222,In_417,In_847);
and U223 (N_223,In_861,In_563);
xor U224 (N_224,In_1053,In_505);
xor U225 (N_225,In_362,In_678);
or U226 (N_226,In_351,In_744);
nand U227 (N_227,In_156,In_78);
or U228 (N_228,In_271,In_129);
and U229 (N_229,In_701,In_260);
xnor U230 (N_230,In_518,In_1153);
nor U231 (N_231,In_934,In_353);
nand U232 (N_232,In_1099,In_1431);
xor U233 (N_233,In_73,In_1414);
and U234 (N_234,In_448,N_105);
nand U235 (N_235,In_289,In_865);
nand U236 (N_236,In_1001,In_845);
and U237 (N_237,In_618,In_973);
nor U238 (N_238,In_224,In_713);
xnor U239 (N_239,In_281,In_1389);
or U240 (N_240,In_359,In_95);
xnor U241 (N_241,N_119,In_503);
xnor U242 (N_242,In_310,N_42);
or U243 (N_243,In_52,In_632);
and U244 (N_244,In_323,N_89);
or U245 (N_245,In_284,In_890);
xnor U246 (N_246,In_870,In_456);
xnor U247 (N_247,In_1396,In_820);
nor U248 (N_248,N_17,N_72);
or U249 (N_249,In_703,In_619);
or U250 (N_250,In_681,In_651);
or U251 (N_251,In_150,In_287);
xnor U252 (N_252,In_1322,In_338);
nor U253 (N_253,In_490,In_1146);
nand U254 (N_254,In_11,In_889);
or U255 (N_255,In_1058,In_984);
or U256 (N_256,In_390,In_1466);
or U257 (N_257,In_1464,In_1499);
or U258 (N_258,In_319,In_450);
or U259 (N_259,In_980,In_624);
and U260 (N_260,In_1353,In_1088);
xnor U261 (N_261,In_1104,N_106);
nand U262 (N_262,In_1331,In_279);
or U263 (N_263,N_14,N_7);
nand U264 (N_264,In_773,N_209);
nor U265 (N_265,In_81,In_721);
xnor U266 (N_266,N_225,In_366);
nor U267 (N_267,N_108,In_1178);
nor U268 (N_268,In_558,N_81);
or U269 (N_269,In_928,In_706);
and U270 (N_270,In_74,In_494);
nand U271 (N_271,N_174,N_232);
nor U272 (N_272,In_39,In_401);
xor U273 (N_273,N_19,In_179);
nand U274 (N_274,In_948,N_120);
and U275 (N_275,In_639,In_1227);
or U276 (N_276,N_140,N_45);
nor U277 (N_277,In_215,In_958);
nor U278 (N_278,In_1309,In_1013);
or U279 (N_279,In_601,In_286);
or U280 (N_280,N_151,In_70);
nand U281 (N_281,In_1204,N_197);
or U282 (N_282,In_1225,In_155);
nor U283 (N_283,In_342,In_954);
and U284 (N_284,In_240,N_88);
xnor U285 (N_285,N_43,In_8);
or U286 (N_286,In_1275,In_251);
xnor U287 (N_287,In_1005,In_949);
and U288 (N_288,N_183,In_943);
nor U289 (N_289,In_143,In_1314);
nor U290 (N_290,In_534,N_115);
nor U291 (N_291,In_1486,N_135);
and U292 (N_292,In_96,N_234);
or U293 (N_293,In_598,In_580);
or U294 (N_294,In_88,In_4);
nor U295 (N_295,In_1377,N_84);
nor U296 (N_296,In_789,In_894);
nand U297 (N_297,In_658,In_130);
nor U298 (N_298,In_1321,In_1000);
and U299 (N_299,N_4,In_421);
nor U300 (N_300,N_172,In_458);
nor U301 (N_301,In_133,In_425);
and U302 (N_302,N_176,N_242);
nor U303 (N_303,In_562,In_904);
nor U304 (N_304,In_1162,In_1351);
xor U305 (N_305,N_220,N_40);
nor U306 (N_306,In_275,In_530);
nand U307 (N_307,In_1406,In_345);
nand U308 (N_308,N_155,In_795);
and U309 (N_309,In_1120,In_524);
and U310 (N_310,N_186,In_689);
and U311 (N_311,In_734,In_22);
nor U312 (N_312,In_950,In_808);
nand U313 (N_313,N_147,In_1043);
nand U314 (N_314,In_1239,In_500);
or U315 (N_315,In_818,In_398);
and U316 (N_316,N_215,In_100);
nand U317 (N_317,In_722,In_747);
nor U318 (N_318,In_938,In_501);
xnor U319 (N_319,In_1247,In_437);
and U320 (N_320,In_1298,N_246);
nand U321 (N_321,In_170,N_201);
and U322 (N_322,In_777,In_858);
and U323 (N_323,In_412,In_640);
nor U324 (N_324,In_1405,In_23);
nor U325 (N_325,In_208,In_1073);
xor U326 (N_326,In_1352,N_149);
nand U327 (N_327,In_1165,In_1261);
nand U328 (N_328,In_852,In_447);
nand U329 (N_329,In_664,In_1060);
nor U330 (N_330,In_1115,In_316);
or U331 (N_331,In_1170,In_1221);
nand U332 (N_332,In_912,In_270);
nor U333 (N_333,In_848,In_631);
and U334 (N_334,In_883,In_309);
and U335 (N_335,In_1447,In_799);
or U336 (N_336,In_964,N_65);
and U337 (N_337,N_134,In_708);
nand U338 (N_338,In_840,In_1188);
nand U339 (N_339,In_1448,In_243);
and U340 (N_340,In_1350,N_231);
or U341 (N_341,In_635,N_238);
and U342 (N_342,In_402,In_1476);
nor U343 (N_343,In_1304,In_355);
or U344 (N_344,In_833,In_369);
xor U345 (N_345,In_1136,In_171);
nor U346 (N_346,In_614,N_241);
and U347 (N_347,In_1354,In_1198);
nand U348 (N_348,N_173,N_12);
nor U349 (N_349,In_1105,In_302);
xor U350 (N_350,In_492,In_1346);
nor U351 (N_351,In_712,In_602);
and U352 (N_352,In_1229,In_975);
and U353 (N_353,In_550,In_1367);
xor U354 (N_354,In_42,N_138);
nand U355 (N_355,In_1145,In_754);
nor U356 (N_356,In_498,In_613);
xor U357 (N_357,N_21,In_740);
or U358 (N_358,In_1277,In_1349);
nor U359 (N_359,In_764,N_129);
or U360 (N_360,In_326,In_735);
nor U361 (N_361,N_189,In_272);
or U362 (N_362,In_728,In_71);
or U363 (N_363,In_1191,In_1449);
nor U364 (N_364,N_85,N_153);
nand U365 (N_365,In_962,In_290);
xor U366 (N_366,In_675,In_942);
xnor U367 (N_367,N_50,In_857);
nor U368 (N_368,In_753,In_538);
xor U369 (N_369,N_27,In_1428);
nand U370 (N_370,In_1025,In_185);
nor U371 (N_371,N_51,N_90);
and U372 (N_372,In_261,In_731);
xnor U373 (N_373,In_955,In_626);
xor U374 (N_374,In_249,In_1015);
nand U375 (N_375,N_334,In_483);
and U376 (N_376,In_504,N_110);
and U377 (N_377,In_1407,In_520);
or U378 (N_378,In_1408,N_74);
nor U379 (N_379,In_57,In_1091);
or U380 (N_380,In_1056,N_210);
or U381 (N_381,N_168,N_75);
xor U382 (N_382,In_62,In_1199);
nand U383 (N_383,N_13,In_1338);
nor U384 (N_384,In_1451,In_442);
or U385 (N_385,N_182,In_1093);
and U386 (N_386,In_285,In_1205);
nor U387 (N_387,In_517,In_5);
nor U388 (N_388,In_582,N_353);
xnor U389 (N_389,In_680,In_465);
or U390 (N_390,In_1327,In_573);
and U391 (N_391,N_48,In_1213);
and U392 (N_392,In_1333,In_365);
nor U393 (N_393,N_167,In_405);
nor U394 (N_394,In_1242,N_226);
xnor U395 (N_395,N_55,In_140);
and U396 (N_396,In_535,N_330);
and U397 (N_397,N_1,In_477);
nand U398 (N_398,In_1034,In_854);
nand U399 (N_399,In_1062,In_1155);
or U400 (N_400,N_341,In_779);
xnor U401 (N_401,In_300,N_301);
xor U402 (N_402,N_156,N_273);
or U403 (N_403,In_1373,In_855);
nor U404 (N_404,N_69,In_682);
or U405 (N_405,In_1462,In_86);
nor U406 (N_406,In_1085,N_248);
nor U407 (N_407,In_516,In_1187);
nor U408 (N_408,In_262,In_1233);
and U409 (N_409,In_392,In_1318);
xnor U410 (N_410,In_222,N_53);
nand U411 (N_411,In_210,In_1208);
nor U412 (N_412,In_971,In_1049);
or U413 (N_413,N_202,In_893);
xor U414 (N_414,In_525,In_2);
nand U415 (N_415,In_1433,In_108);
xnor U416 (N_416,In_104,In_191);
or U417 (N_417,In_591,N_144);
or U418 (N_418,N_198,N_325);
nand U419 (N_419,N_308,In_565);
nand U420 (N_420,In_1175,N_304);
and U421 (N_421,In_736,N_247);
xor U422 (N_422,In_575,In_495);
and U423 (N_423,In_1393,In_1323);
or U424 (N_424,In_1276,In_51);
nor U425 (N_425,In_230,N_358);
nor U426 (N_426,In_568,N_97);
or U427 (N_427,In_644,In_107);
nand U428 (N_428,N_298,In_1135);
or U429 (N_429,N_39,In_1303);
or U430 (N_430,N_233,In_813);
nor U431 (N_431,In_888,In_816);
and U432 (N_432,In_205,N_166);
nand U433 (N_433,In_1470,In_159);
and U434 (N_434,In_276,In_1399);
nand U435 (N_435,In_1141,In_328);
xor U436 (N_436,In_1241,In_1166);
and U437 (N_437,In_1475,In_961);
or U438 (N_438,In_698,In_1209);
or U439 (N_439,N_141,In_622);
nand U440 (N_440,N_285,In_352);
and U441 (N_441,In_1036,In_145);
nand U442 (N_442,In_188,In_7);
nor U443 (N_443,In_370,N_57);
nor U444 (N_444,In_749,In_480);
or U445 (N_445,N_265,In_1290);
or U446 (N_446,N_114,N_165);
nor U447 (N_447,In_584,N_299);
nand U448 (N_448,In_1293,In_1436);
nor U449 (N_449,In_1366,N_154);
nand U450 (N_450,In_1273,In_183);
or U451 (N_451,In_922,In_512);
nor U452 (N_452,N_64,N_345);
nand U453 (N_453,N_184,In_511);
and U454 (N_454,In_19,In_781);
xor U455 (N_455,N_329,In_396);
or U456 (N_456,N_157,In_605);
xor U457 (N_457,N_250,In_1004);
xor U458 (N_458,N_288,N_208);
nor U459 (N_459,In_700,In_193);
or U460 (N_460,In_1017,In_400);
nand U461 (N_461,In_12,In_1169);
or U462 (N_462,In_556,N_46);
or U463 (N_463,N_70,N_229);
nand U464 (N_464,In_1059,N_98);
and U465 (N_465,In_220,In_1308);
or U466 (N_466,In_231,N_363);
nor U467 (N_467,N_222,In_386);
xor U468 (N_468,In_1374,In_1151);
nor U469 (N_469,In_1264,In_1332);
nand U470 (N_470,In_173,In_121);
and U471 (N_471,In_604,N_191);
nand U472 (N_472,In_381,N_196);
and U473 (N_473,In_812,N_26);
nor U474 (N_474,In_1429,In_1044);
xor U475 (N_475,In_1174,In_373);
nor U476 (N_476,In_937,In_1189);
nor U477 (N_477,In_1251,In_221);
nand U478 (N_478,N_36,In_898);
and U479 (N_479,In_1226,In_1479);
xnor U480 (N_480,In_1083,N_243);
and U481 (N_481,In_0,N_127);
nor U482 (N_482,N_190,In_707);
or U483 (N_483,In_1259,In_765);
nor U484 (N_484,In_1116,In_668);
nor U485 (N_485,N_123,N_158);
and U486 (N_486,N_252,In_1210);
nand U487 (N_487,In_83,In_1148);
and U488 (N_488,In_199,In_460);
nor U489 (N_489,In_1430,In_673);
nor U490 (N_490,In_901,In_225);
or U491 (N_491,In_1270,N_47);
nand U492 (N_492,In_983,N_181);
and U493 (N_493,In_826,In_1086);
nor U494 (N_494,In_521,In_687);
nor U495 (N_495,In_1458,N_82);
and U496 (N_496,N_77,In_1381);
xnor U497 (N_497,In_112,In_337);
or U498 (N_498,N_193,In_247);
and U499 (N_499,In_1179,In_782);
nand U500 (N_500,In_473,In_1076);
or U501 (N_501,In_125,In_1123);
or U502 (N_502,N_481,N_406);
and U503 (N_503,In_1180,In_474);
nor U504 (N_504,In_685,N_385);
nand U505 (N_505,In_367,In_982);
and U506 (N_506,In_1080,N_472);
nor U507 (N_507,In_1217,In_1415);
nand U508 (N_508,In_168,N_409);
or U509 (N_509,In_1211,N_20);
or U510 (N_510,In_864,N_432);
nor U511 (N_511,In_227,In_834);
nor U512 (N_512,N_442,In_1280);
or U513 (N_513,In_991,In_1118);
nand U514 (N_514,In_481,N_177);
nand U515 (N_515,N_274,N_67);
and U516 (N_516,N_326,N_347);
and U517 (N_517,In_819,N_336);
or U518 (N_518,N_271,N_54);
or U519 (N_519,In_567,In_435);
xnor U520 (N_520,N_436,In_165);
nor U521 (N_521,In_776,In_343);
nand U522 (N_522,In_770,In_946);
xnor U523 (N_523,In_1134,In_1301);
xor U524 (N_524,In_630,In_37);
nor U525 (N_525,N_381,In_371);
nand U526 (N_526,In_85,In_267);
and U527 (N_527,In_1329,N_403);
or U528 (N_528,In_726,In_1439);
nand U529 (N_529,N_324,N_438);
or U530 (N_530,N_456,N_462);
nand U531 (N_531,In_1434,In_256);
and U532 (N_532,In_1334,N_486);
xnor U533 (N_533,In_1461,In_960);
nor U534 (N_534,N_460,N_195);
nor U535 (N_535,N_83,In_1218);
and U536 (N_536,In_368,N_29);
and U537 (N_537,In_462,In_625);
and U538 (N_538,N_277,In_1038);
nand U539 (N_539,N_346,In_609);
xor U540 (N_540,In_1268,N_391);
nand U541 (N_541,In_228,N_465);
xor U542 (N_542,In_389,In_1419);
or U543 (N_543,In_47,In_686);
xor U544 (N_544,In_545,N_466);
or U545 (N_545,In_830,N_94);
nor U546 (N_546,N_498,In_115);
nand U547 (N_547,N_322,N_263);
or U548 (N_548,In_716,In_356);
xor U549 (N_549,In_1435,N_313);
or U550 (N_550,N_314,In_918);
xnor U551 (N_551,In_1066,In_1031);
nor U552 (N_552,In_297,In_1263);
nor U553 (N_553,N_464,N_41);
or U554 (N_554,In_597,N_192);
nor U555 (N_555,In_531,N_267);
and U556 (N_556,N_344,N_439);
nor U557 (N_557,N_453,In_1262);
or U558 (N_558,In_1019,N_440);
or U559 (N_559,In_1063,In_846);
nor U560 (N_560,In_1245,In_549);
nor U561 (N_561,In_691,In_590);
and U562 (N_562,N_398,N_188);
and U563 (N_563,N_73,In_1274);
nor U564 (N_564,In_471,In_1404);
nand U565 (N_565,In_654,N_170);
nor U566 (N_566,In_650,In_710);
xor U567 (N_567,N_386,N_200);
nand U568 (N_568,In_508,In_1256);
xnor U569 (N_569,In_798,In_407);
nor U570 (N_570,In_123,In_470);
nand U571 (N_571,N_476,In_759);
nand U572 (N_572,In_1173,In_278);
nand U573 (N_573,N_87,In_985);
or U574 (N_574,N_365,In_1459);
and U575 (N_575,N_493,In_1278);
and U576 (N_576,In_1359,N_62);
nand U577 (N_577,N_312,N_228);
nand U578 (N_578,N_289,In_478);
xnor U579 (N_579,In_109,N_293);
nor U580 (N_580,In_68,In_1074);
nor U581 (N_581,In_1159,In_119);
xnor U582 (N_582,In_876,N_292);
and U583 (N_583,In_312,N_337);
or U584 (N_584,In_566,N_359);
nor U585 (N_585,N_162,In_696);
and U586 (N_586,In_510,N_103);
xnor U587 (N_587,In_652,In_807);
and U588 (N_588,In_114,In_455);
xor U589 (N_589,In_745,N_467);
nand U590 (N_590,In_166,In_14);
nor U591 (N_591,In_264,In_295);
and U592 (N_592,In_186,N_113);
and U593 (N_593,In_413,In_233);
nor U594 (N_594,N_443,N_429);
and U595 (N_595,N_143,In_1228);
nand U596 (N_596,In_90,In_348);
nor U597 (N_597,In_952,In_758);
or U598 (N_598,In_1018,N_206);
and U599 (N_599,In_484,In_1006);
and U600 (N_600,N_327,In_461);
nor U601 (N_601,In_572,N_32);
or U602 (N_602,In_1257,N_416);
xor U603 (N_603,N_109,N_390);
nand U604 (N_604,In_925,In_82);
xor U605 (N_605,In_1069,In_1283);
nor U606 (N_606,In_1114,In_1375);
nand U607 (N_607,N_457,N_139);
and U608 (N_608,In_1342,In_1469);
nand U609 (N_609,N_33,N_321);
or U610 (N_610,In_947,In_674);
nor U611 (N_611,In_1296,In_1028);
and U612 (N_612,In_1109,In_660);
and U613 (N_613,In_6,In_576);
nand U614 (N_614,In_102,In_395);
nand U615 (N_615,N_131,In_347);
or U616 (N_616,N_133,In_321);
xnor U617 (N_617,In_1403,N_393);
nor U618 (N_618,N_489,In_1011);
or U619 (N_619,In_420,N_258);
xor U620 (N_620,In_92,In_778);
or U621 (N_621,N_378,In_853);
nand U622 (N_622,In_772,N_389);
or U623 (N_623,N_211,In_1491);
nand U624 (N_624,In_1160,N_305);
nand U625 (N_625,In_10,N_474);
xor U626 (N_626,N_379,N_503);
nand U627 (N_627,In_1306,In_237);
nor U628 (N_628,N_506,In_1284);
nand U629 (N_629,N_61,In_884);
xnor U630 (N_630,In_1416,N_34);
xor U631 (N_631,In_1471,In_1142);
and U632 (N_632,N_455,N_427);
or U633 (N_633,In_737,In_20);
and U634 (N_634,N_586,In_304);
nand U635 (N_635,In_900,N_566);
nor U636 (N_636,In_746,N_9);
nand U637 (N_637,In_607,N_490);
nor U638 (N_638,N_382,N_317);
xor U639 (N_639,In_1455,In_1224);
and U640 (N_640,N_610,N_412);
and U641 (N_641,In_1494,N_362);
and U642 (N_642,In_60,N_2);
or U643 (N_643,In_617,In_1420);
or U644 (N_644,In_91,In_134);
xnor U645 (N_645,In_229,N_264);
and U646 (N_646,In_135,In_110);
xor U647 (N_647,In_877,In_1391);
and U648 (N_648,N_116,In_1425);
nand U649 (N_649,In_987,In_375);
or U650 (N_650,N_377,N_600);
nand U651 (N_651,In_58,N_323);
nor U652 (N_652,In_303,N_392);
nand U653 (N_653,In_489,N_601);
nor U654 (N_654,In_344,N_614);
and U655 (N_655,In_793,N_256);
nor U656 (N_656,N_402,In_739);
and U657 (N_657,In_349,In_1484);
nor U658 (N_658,N_372,In_606);
and U659 (N_659,In_466,In_727);
nor U660 (N_660,In_695,In_688);
xor U661 (N_661,N_599,In_248);
xor U662 (N_662,In_330,In_265);
or U663 (N_663,N_212,In_1212);
and U664 (N_664,In_923,In_989);
nor U665 (N_665,In_610,N_619);
or U666 (N_666,In_583,In_560);
nand U667 (N_667,N_169,In_1295);
or U668 (N_668,N_249,N_618);
nand U669 (N_669,In_992,In_329);
xnor U670 (N_670,N_331,In_48);
or U671 (N_671,N_613,In_873);
xnor U672 (N_672,N_92,N_16);
nor U673 (N_673,N_617,In_1426);
xnor U674 (N_674,In_200,In_762);
nor U675 (N_675,N_418,In_1402);
or U676 (N_676,N_124,In_313);
nand U677 (N_677,In_31,In_1398);
nand U678 (N_678,N_370,In_1124);
and U679 (N_679,N_396,N_355);
nand U680 (N_680,N_606,N_538);
nand U681 (N_681,N_422,In_332);
nor U682 (N_682,N_354,In_786);
or U683 (N_683,In_30,In_970);
nand U684 (N_684,In_1202,N_413);
and U685 (N_685,In_1441,N_259);
nor U686 (N_686,In_207,In_41);
and U687 (N_687,In_529,N_482);
nor U688 (N_688,In_1032,In_1042);
or U689 (N_689,In_1258,In_1238);
nand U690 (N_690,In_885,In_641);
nor U691 (N_691,N_517,N_150);
and U692 (N_692,N_342,In_578);
or U693 (N_693,In_423,In_757);
nor U694 (N_694,In_679,In_1138);
and U695 (N_695,N_214,In_1330);
xnor U696 (N_696,N_117,In_1067);
nand U697 (N_697,In_1054,N_588);
xnor U698 (N_698,In_487,N_449);
nand U699 (N_699,In_709,N_473);
xnor U700 (N_700,In_305,N_203);
nor U701 (N_701,N_338,In_172);
or U702 (N_702,In_809,In_291);
nor U703 (N_703,N_171,In_216);
nor U704 (N_704,N_468,N_270);
nand U705 (N_705,N_510,In_515);
or U706 (N_706,In_1201,In_1291);
nor U707 (N_707,In_475,In_147);
and U708 (N_708,In_769,In_771);
nor U709 (N_709,N_559,In_383);
nand U710 (N_710,N_428,N_415);
or U711 (N_711,N_395,In_986);
nor U712 (N_712,In_76,In_841);
xnor U713 (N_713,In_1048,In_146);
or U714 (N_714,N_311,In_1246);
nor U715 (N_715,In_1007,In_238);
nand U716 (N_716,N_235,N_333);
and U717 (N_717,In_250,In_1243);
or U718 (N_718,In_1358,In_1473);
and U719 (N_719,N_479,In_902);
xor U720 (N_720,In_1021,In_1194);
xor U721 (N_721,In_1440,N_561);
xnor U722 (N_722,N_507,In_1022);
xnor U723 (N_723,In_959,N_574);
nand U724 (N_724,N_485,In_499);
nand U725 (N_725,In_579,In_122);
or U726 (N_726,N_194,N_602);
nor U727 (N_727,N_594,In_1095);
xor U728 (N_728,N_477,N_480);
xor U729 (N_729,N_269,In_1372);
nor U730 (N_730,In_467,In_1348);
nor U731 (N_731,In_723,N_224);
and U732 (N_732,In_154,In_1368);
xnor U733 (N_733,N_611,N_303);
nand U734 (N_734,N_445,N_533);
nand U735 (N_735,In_226,N_187);
xor U736 (N_736,N_549,In_438);
nor U737 (N_737,In_246,In_1237);
nand U738 (N_738,In_1087,N_282);
nor U739 (N_739,N_543,In_875);
nor U740 (N_740,In_1297,In_1252);
and U741 (N_741,In_653,N_78);
or U742 (N_742,N_60,N_261);
and U743 (N_743,In_16,In_1310);
xnor U744 (N_744,N_219,In_724);
and U745 (N_745,N_221,N_450);
and U746 (N_746,In_124,In_192);
or U747 (N_747,N_22,In_1183);
nor U748 (N_748,In_127,In_138);
xor U749 (N_749,N_504,N_268);
and U750 (N_750,In_36,N_641);
nor U751 (N_751,N_740,N_297);
nor U752 (N_752,N_548,N_478);
and U753 (N_753,N_281,N_496);
nor U754 (N_754,In_1137,N_744);
nand U755 (N_755,In_945,In_1269);
or U756 (N_756,N_520,In_523);
or U757 (N_757,N_578,N_148);
xnor U758 (N_758,N_25,In_797);
or U759 (N_759,In_144,N_560);
nand U760 (N_760,In_1203,N_146);
or U761 (N_761,N_714,In_926);
xnor U762 (N_762,In_1002,In_196);
nand U763 (N_763,N_539,In_441);
nand U764 (N_764,In_720,In_859);
xor U765 (N_765,In_1395,In_322);
and U766 (N_766,N_551,N_260);
nand U767 (N_767,N_707,N_49);
or U768 (N_768,In_419,In_1128);
or U769 (N_769,N_152,N_679);
nor U770 (N_770,N_747,In_234);
or U771 (N_771,N_505,In_294);
nor U772 (N_772,In_554,N_729);
and U773 (N_773,N_591,In_357);
and U774 (N_774,In_244,In_871);
nand U775 (N_775,N_724,In_175);
and U776 (N_776,N_589,In_1289);
and U777 (N_777,In_1443,N_502);
nand U778 (N_778,In_775,In_1271);
nand U779 (N_779,N_532,N_286);
nor U780 (N_780,In_616,N_604);
nor U781 (N_781,N_735,In_17);
nor U782 (N_782,N_556,N_137);
xor U783 (N_783,N_576,In_828);
and U784 (N_784,N_652,In_1385);
and U785 (N_785,N_484,N_689);
xnor U786 (N_786,N_446,N_410);
xor U787 (N_787,In_993,N_488);
nor U788 (N_788,N_66,In_967);
or U789 (N_789,N_681,In_77);
nor U790 (N_790,N_579,In_1106);
nor U791 (N_791,In_66,In_1400);
nor U792 (N_792,N_581,N_458);
and U793 (N_793,In_1016,N_470);
or U794 (N_794,N_128,N_435);
xor U795 (N_795,In_209,In_1307);
nand U796 (N_796,N_553,In_1113);
nand U797 (N_797,N_616,N_475);
xnor U798 (N_798,In_1260,In_1255);
nor U799 (N_799,N_701,N_694);
nand U800 (N_800,N_609,N_585);
or U801 (N_801,N_375,In_334);
nor U802 (N_802,N_732,N_28);
and U803 (N_803,N_111,N_628);
nand U804 (N_804,N_463,In_1167);
nand U805 (N_805,N_659,N_276);
and U806 (N_806,In_217,In_379);
nor U807 (N_807,N_245,In_1409);
nor U808 (N_808,In_335,In_879);
or U809 (N_809,In_905,N_667);
nand U810 (N_810,N_597,In_718);
or U811 (N_811,N_44,In_1424);
nand U812 (N_812,N_180,N_5);
and U813 (N_813,In_1340,N_163);
nand U814 (N_814,In_513,N_280);
and U815 (N_815,In_380,In_1254);
or U816 (N_816,In_1140,In_881);
xor U817 (N_817,In_526,In_944);
or U818 (N_818,N_96,In_479);
nor U819 (N_819,N_709,N_526);
nor U820 (N_820,In_805,N_237);
and U821 (N_821,N_290,In_637);
nand U822 (N_822,In_1496,In_320);
xnor U823 (N_823,In_314,N_63);
and U824 (N_824,In_792,N_657);
xnor U825 (N_825,N_572,N_535);
and U826 (N_826,In_1438,In_1444);
nor U827 (N_827,In_1089,N_651);
nand U828 (N_828,N_309,In_811);
or U829 (N_829,N_272,In_1453);
nor U830 (N_830,In_827,In_457);
nor U831 (N_831,N_430,In_1100);
or U832 (N_832,In_647,N_279);
xnor U833 (N_833,N_284,In_502);
or U834 (N_834,N_217,N_38);
or U835 (N_835,N_702,N_615);
or U836 (N_836,N_431,N_545);
xor U837 (N_837,N_207,N_302);
nand U838 (N_838,N_411,In_825);
nor U839 (N_839,N_291,In_169);
and U840 (N_840,N_204,In_452);
or U841 (N_841,N_487,N_319);
and U842 (N_842,In_585,N_524);
xor U843 (N_843,In_252,N_642);
xnor U844 (N_844,N_629,In_1077);
xnor U845 (N_845,In_1347,N_511);
xnor U846 (N_846,N_704,N_546);
nand U847 (N_847,N_491,In_255);
xnor U848 (N_848,N_699,N_587);
nand U849 (N_849,In_571,N_671);
xor U850 (N_850,In_1040,In_1355);
xnor U851 (N_851,N_91,N_633);
xor U852 (N_852,N_593,N_494);
or U853 (N_853,N_361,In_274);
or U854 (N_854,In_551,N_230);
nor U855 (N_855,In_1096,In_75);
nor U856 (N_856,In_488,N_649);
nand U857 (N_857,In_1324,N_437);
and U858 (N_858,N_716,N_380);
or U859 (N_859,N_352,In_866);
xnor U860 (N_860,N_145,N_595);
and U861 (N_861,N_662,In_382);
or U862 (N_862,N_332,N_35);
or U863 (N_863,N_731,In_1286);
nor U864 (N_864,N_541,In_497);
and U865 (N_865,N_567,N_254);
nand U866 (N_866,N_278,N_310);
nor U867 (N_867,In_643,N_682);
and U868 (N_868,N_441,N_497);
or U869 (N_869,N_397,In_627);
nor U870 (N_870,In_1101,N_557);
nor U871 (N_871,In_896,In_410);
and U872 (N_872,N_605,N_692);
and U873 (N_873,In_1492,In_1185);
and U874 (N_874,In_908,N_634);
and U875 (N_875,N_661,N_632);
nand U876 (N_876,In_804,N_672);
xnor U877 (N_877,N_399,N_349);
nor U878 (N_878,N_858,In_79);
and U879 (N_879,N_748,N_798);
nor U880 (N_880,In_1483,N_501);
xor U881 (N_881,N_813,N_575);
nand U882 (N_882,N_130,In_94);
and U883 (N_883,N_847,N_693);
and U884 (N_884,N_454,In_429);
and U885 (N_885,In_886,N_93);
nor U886 (N_886,In_1027,N_653);
or U887 (N_887,In_56,N_11);
nand U888 (N_888,N_550,In_105);
or U889 (N_889,N_255,N_637);
and U890 (N_890,In_638,N_296);
xnor U891 (N_891,N_287,In_1370);
nor U892 (N_892,In_957,N_540);
xnor U893 (N_893,In_106,N_712);
xor U894 (N_894,N_374,N_780);
nand U895 (N_895,In_84,In_909);
or U896 (N_896,N_726,N_320);
xor U897 (N_897,N_730,N_762);
xnor U898 (N_898,N_778,N_373);
xor U899 (N_899,N_817,In_254);
nor U900 (N_900,N_644,N_218);
and U901 (N_901,In_388,In_1482);
and U902 (N_902,In_116,In_998);
or U903 (N_903,In_788,N_741);
nand U904 (N_904,N_826,In_1045);
or U905 (N_905,In_672,N_519);
nand U906 (N_906,N_752,In_26);
nor U907 (N_907,In_924,In_514);
nand U908 (N_908,N_779,N_697);
xnor U909 (N_909,In_424,N_419);
nand U910 (N_910,In_995,N_737);
and U911 (N_911,N_71,N_627);
nor U912 (N_912,N_754,N_797);
nand U913 (N_913,In_552,N_216);
xor U914 (N_914,In_269,N_266);
nand U915 (N_915,In_195,N_125);
xnor U916 (N_916,N_227,N_185);
or U917 (N_917,N_364,In_823);
or U918 (N_918,In_705,N_59);
and U919 (N_919,In_1478,In_288);
or U920 (N_920,N_294,N_768);
nand U921 (N_921,N_580,In_432);
or U922 (N_922,In_1383,N_625);
or U923 (N_923,N_620,N_755);
nand U924 (N_924,N_315,N_573);
xnor U925 (N_925,In_341,In_1493);
nor U926 (N_926,N_867,N_95);
or U927 (N_927,In_360,N_544);
and U928 (N_928,In_1356,In_93);
nor U929 (N_929,N_806,N_824);
nor U930 (N_930,In_1336,N_663);
or U931 (N_931,In_213,In_1129);
nand U932 (N_932,N_700,In_1126);
nor U933 (N_933,N_792,In_802);
or U934 (N_934,In_454,In_965);
xor U935 (N_935,In_376,N_76);
nor U936 (N_936,In_1361,N_328);
nand U937 (N_937,N_306,N_795);
nor U938 (N_938,N_853,In_253);
xor U939 (N_939,In_548,N_542);
xnor U940 (N_940,In_1033,N_674);
and U941 (N_941,N_417,N_509);
and U942 (N_942,In_1003,N_626);
nand U943 (N_943,N_800,In_152);
and U944 (N_944,N_547,N_703);
nand U945 (N_945,N_240,N_750);
nand U946 (N_946,N_783,N_583);
and U947 (N_947,N_769,In_794);
and U948 (N_948,N_713,In_796);
nor U949 (N_949,N_676,N_360);
and U950 (N_950,N_828,N_534);
and U951 (N_951,N_469,In_18);
nand U952 (N_952,In_1014,In_761);
nor U953 (N_953,In_1125,N_102);
nand U954 (N_954,N_257,N_845);
nand U955 (N_955,N_199,N_854);
nor U956 (N_956,In_751,N_205);
and U957 (N_957,N_592,N_384);
nand U958 (N_958,In_1231,N_368);
and U959 (N_959,In_1345,In_1026);
nor U960 (N_960,N_760,N_864);
or U961 (N_961,N_805,N_774);
nand U962 (N_962,In_935,N_855);
and U963 (N_963,N_832,N_691);
nand U964 (N_964,N_723,N_809);
nor U965 (N_965,N_743,In_99);
nor U966 (N_966,In_45,In_132);
and U967 (N_967,In_1497,In_1401);
nand U968 (N_968,N_670,N_236);
or U969 (N_969,N_829,N_552);
nand U970 (N_970,In_167,In_581);
nor U971 (N_971,N_677,N_758);
or U972 (N_972,In_692,N_648);
xnor U973 (N_973,In_61,N_823);
xor U974 (N_974,In_35,In_784);
xnor U975 (N_975,In_1387,N_782);
and U976 (N_976,In_27,N_569);
nand U977 (N_977,N_696,In_714);
or U978 (N_978,N_787,N_733);
and U979 (N_979,N_664,In_141);
xor U980 (N_980,In_1010,In_1397);
xnor U981 (N_981,N_518,N_745);
or U982 (N_982,N_831,N_756);
nor U983 (N_983,In_1051,In_930);
xor U984 (N_984,N_655,In_394);
or U985 (N_985,In_472,N_536);
nand U986 (N_986,In_1192,In_1240);
nor U987 (N_987,N_495,N_376);
nor U988 (N_988,N_508,N_857);
or U989 (N_989,In_1234,N_444);
or U990 (N_990,N_673,In_756);
or U991 (N_991,N_631,N_827);
and U992 (N_992,N_523,N_424);
and U993 (N_993,In_1460,N_686);
nor U994 (N_994,N_819,N_821);
xor U995 (N_995,In_1337,In_1344);
and U996 (N_996,In_340,In_1467);
and U997 (N_997,In_559,N_262);
nand U998 (N_998,In_50,N_564);
nor U999 (N_999,In_994,N_788);
xor U1000 (N_1000,N_647,N_669);
and U1001 (N_1001,N_521,N_335);
or U1002 (N_1002,In_65,N_781);
nor U1003 (N_1003,N_932,N_923);
or U1004 (N_1004,N_807,N_295);
or U1005 (N_1005,In_1207,In_676);
and U1006 (N_1006,N_565,N_959);
or U1007 (N_1007,N_895,In_1154);
nor U1008 (N_1008,N_515,N_388);
nand U1009 (N_1009,N_80,N_964);
and U1010 (N_1010,N_837,In_1107);
xnor U1011 (N_1011,In_974,N_448);
xnor U1012 (N_1012,N_979,N_926);
and U1013 (N_1013,N_434,In_981);
nand U1014 (N_1014,N_537,In_308);
xor U1015 (N_1015,N_688,In_358);
or U1016 (N_1016,N_955,N_896);
nor U1017 (N_1017,N_394,N_164);
and U1018 (N_1018,N_654,N_811);
or U1019 (N_1019,N_367,N_514);
or U1020 (N_1020,N_859,N_851);
or U1021 (N_1021,N_865,In_887);
xor U1022 (N_1022,N_316,N_968);
xor U1023 (N_1023,N_757,In_1319);
nand U1024 (N_1024,N_638,N_999);
nor U1025 (N_1025,N_630,N_793);
or U1026 (N_1026,N_905,N_994);
or U1027 (N_1027,N_516,N_898);
and U1028 (N_1028,In_1376,N_965);
and U1029 (N_1029,In_532,N_767);
nand U1030 (N_1030,In_1046,In_257);
nand U1031 (N_1031,In_1328,N_658);
nand U1032 (N_1032,N_734,N_223);
xor U1033 (N_1033,N_947,In_899);
or U1034 (N_1034,N_300,N_251);
and U1035 (N_1035,N_350,In_293);
and U1036 (N_1036,N_283,In_546);
xor U1037 (N_1037,N_608,N_708);
xnor U1038 (N_1038,N_969,N_986);
and U1039 (N_1039,In_307,N_951);
or U1040 (N_1040,In_414,N_815);
nand U1041 (N_1041,N_684,N_351);
nor U1042 (N_1042,N_948,N_776);
xnor U1043 (N_1043,N_582,N_914);
nor U1044 (N_1044,N_977,N_887);
and U1045 (N_1045,N_791,In_137);
xnor U1046 (N_1046,N_933,N_126);
nand U1047 (N_1047,N_636,In_1412);
nand U1048 (N_1048,In_1299,N_356);
xor U1049 (N_1049,N_132,N_846);
xor U1050 (N_1050,N_830,N_839);
or U1051 (N_1051,N_906,N_911);
and U1052 (N_1052,N_159,N_571);
or U1053 (N_1053,N_30,In_608);
nor U1054 (N_1054,N_773,N_953);
or U1055 (N_1055,In_1265,N_623);
or U1056 (N_1056,In_1481,N_891);
nor U1057 (N_1057,N_820,N_975);
xor U1058 (N_1058,N_850,N_885);
or U1059 (N_1059,N_777,N_869);
xnor U1060 (N_1060,In_785,N_861);
or U1061 (N_1061,N_160,N_812);
and U1062 (N_1062,N_946,N_721);
nand U1063 (N_1063,N_698,N_993);
and U1064 (N_1064,N_890,N_68);
and U1065 (N_1065,In_1485,N_901);
nor U1066 (N_1066,N_997,In_1244);
nor U1067 (N_1067,N_404,N_3);
xnor U1068 (N_1068,N_622,N_920);
nand U1069 (N_1069,N_840,N_121);
xnor U1070 (N_1070,N_881,In_1182);
and U1071 (N_1071,In_1133,N_835);
and U1072 (N_1072,N_991,N_842);
nor U1073 (N_1073,N_717,N_531);
and U1074 (N_1074,N_889,N_984);
nand U1075 (N_1075,N_961,N_763);
or U1076 (N_1076,In_336,N_461);
xnor U1077 (N_1077,N_528,N_801);
xnor U1078 (N_1078,N_680,N_913);
nand U1079 (N_1079,N_142,In_1288);
xor U1080 (N_1080,N_998,In_733);
nand U1081 (N_1081,N_570,In_1186);
nor U1082 (N_1082,N_366,N_753);
or U1083 (N_1083,In_236,In_1362);
or U1084 (N_1084,N_876,N_941);
or U1085 (N_1085,N_957,N_383);
or U1086 (N_1086,In_621,N_856);
xnor U1087 (N_1087,N_872,N_175);
xnor U1088 (N_1088,In_824,N_990);
and U1089 (N_1089,In_139,N_775);
and U1090 (N_1090,N_790,N_451);
nand U1091 (N_1091,N_884,In_1052);
nand U1092 (N_1092,N_967,N_690);
xnor U1093 (N_1093,N_401,N_814);
and U1094 (N_1094,N_499,In_829);
or U1095 (N_1095,In_318,N_972);
nor U1096 (N_1096,N_900,In_750);
or U1097 (N_1097,In_555,N_433);
xnor U1098 (N_1098,N_940,In_1437);
or U1099 (N_1099,In_372,N_874);
nor U1100 (N_1100,In_927,N_339);
or U1101 (N_1101,In_774,N_0);
and U1102 (N_1102,N_759,In_656);
nand U1103 (N_1103,N_665,N_749);
xnor U1104 (N_1104,N_985,N_612);
and U1105 (N_1105,N_122,N_897);
and U1106 (N_1106,N_555,N_852);
nor U1107 (N_1107,N_136,In_670);
nor U1108 (N_1108,N_99,In_1446);
and U1109 (N_1109,N_942,N_725);
nor U1110 (N_1110,N_414,N_529);
and U1111 (N_1111,N_675,N_79);
nand U1112 (N_1112,In_730,N_640);
xnor U1113 (N_1113,N_275,N_907);
nand U1114 (N_1114,In_633,In_953);
and U1115 (N_1115,N_307,N_873);
or U1116 (N_1116,N_838,N_348);
nor U1117 (N_1117,In_843,N_6);
and U1118 (N_1118,N_843,N_908);
or U1119 (N_1119,N_584,N_849);
and U1120 (N_1120,N_844,N_666);
nand U1121 (N_1121,N_988,In_317);
xnor U1122 (N_1122,In_418,N_822);
xnor U1123 (N_1123,In_880,N_603);
nor U1124 (N_1124,In_1030,N_426);
xnor U1125 (N_1125,N_939,N_1015);
xor U1126 (N_1126,N_1039,N_816);
and U1127 (N_1127,N_1037,N_834);
or U1128 (N_1128,N_1012,N_1049);
nor U1129 (N_1129,In_436,N_179);
nand U1130 (N_1130,In_715,N_1071);
or U1131 (N_1131,N_950,N_1113);
nand U1132 (N_1132,N_1058,In_1216);
or U1133 (N_1133,N_1025,N_1086);
and U1134 (N_1134,N_492,N_645);
xor U1135 (N_1135,N_1032,N_1077);
or U1136 (N_1136,N_387,N_1094);
nor U1137 (N_1137,N_785,N_804);
and U1138 (N_1138,In_1220,In_915);
nor U1139 (N_1139,In_1190,N_1084);
nor U1140 (N_1140,N_1062,N_668);
nand U1141 (N_1141,In_755,N_980);
nand U1142 (N_1142,N_357,N_1034);
xor U1143 (N_1143,N_423,N_870);
or U1144 (N_1144,N_1035,N_970);
xnor U1145 (N_1145,N_833,N_1120);
nand U1146 (N_1146,N_400,N_922);
or U1147 (N_1147,N_1006,In_397);
xnor U1148 (N_1148,N_1101,In_684);
and U1149 (N_1149,In_642,In_1150);
nor U1150 (N_1150,N_678,N_405);
and U1151 (N_1151,N_650,N_902);
or U1152 (N_1152,In_1422,In_1498);
or U1153 (N_1153,N_1001,In_868);
nand U1154 (N_1154,N_527,N_746);
and U1155 (N_1155,N_1087,N_685);
and U1156 (N_1156,N_981,In_587);
and U1157 (N_1157,N_910,N_1054);
nand U1158 (N_1158,N_949,N_1081);
nor U1159 (N_1159,N_971,N_371);
and U1160 (N_1160,N_1085,N_764);
xnor U1161 (N_1161,In_160,In_732);
nor U1162 (N_1162,N_1105,N_1046);
xnor U1163 (N_1163,N_802,In_810);
or U1164 (N_1164,N_1114,N_1051);
nand U1165 (N_1165,N_1016,N_1100);
nor U1166 (N_1166,In_1184,N_1036);
nor U1167 (N_1167,N_452,N_1088);
nand U1168 (N_1168,In_699,N_1103);
or U1169 (N_1169,N_1000,N_929);
and U1170 (N_1170,N_808,In_430);
nor U1171 (N_1171,In_663,N_944);
xnor U1172 (N_1172,N_1031,N_1080);
and U1173 (N_1173,N_794,N_893);
and U1174 (N_1174,In_239,N_952);
and U1175 (N_1175,N_766,N_992);
xor U1176 (N_1176,In_117,N_935);
xor U1177 (N_1177,N_945,N_596);
nor U1178 (N_1178,N_1040,N_978);
xnor U1179 (N_1179,N_848,N_720);
and U1180 (N_1180,N_161,N_927);
and U1181 (N_1181,N_878,N_1061);
and U1182 (N_1182,N_738,N_892);
nor U1183 (N_1183,N_1026,N_882);
xnor U1184 (N_1184,N_899,N_1118);
xor U1185 (N_1185,N_868,N_562);
or U1186 (N_1186,N_1018,N_1047);
and U1187 (N_1187,N_1050,N_1115);
and U1188 (N_1188,In_415,N_607);
and U1189 (N_1189,N_639,In_1335);
nor U1190 (N_1190,N_369,N_739);
xnor U1191 (N_1191,N_1045,N_904);
nor U1192 (N_1192,N_1102,N_1029);
xnor U1193 (N_1193,N_863,N_960);
and U1194 (N_1194,N_866,N_803);
and U1195 (N_1195,N_1091,N_1090);
xnor U1196 (N_1196,In_1463,N_879);
and U1197 (N_1197,In_628,N_37);
nand U1198 (N_1198,N_1089,N_1056);
nand U1199 (N_1199,N_917,N_1043);
and U1200 (N_1200,N_983,N_253);
and U1201 (N_1201,In_324,N_343);
xnor U1202 (N_1202,N_982,N_996);
nand U1203 (N_1203,N_918,N_706);
and U1204 (N_1204,N_1097,N_931);
or U1205 (N_1205,N_530,N_727);
nor U1206 (N_1206,N_810,N_912);
nor U1207 (N_1207,N_1093,N_1067);
nor U1208 (N_1208,N_818,N_915);
nand U1209 (N_1209,In_916,N_1108);
nor U1210 (N_1210,N_1063,N_862);
or U1211 (N_1211,N_525,N_1076);
nand U1212 (N_1212,N_1008,N_925);
xnor U1213 (N_1213,N_1003,N_877);
and U1214 (N_1214,N_1066,In_416);
or U1215 (N_1215,N_1073,In_1206);
nand U1216 (N_1216,N_1022,N_1072);
nor U1217 (N_1217,N_1059,N_789);
and U1218 (N_1218,N_15,N_1123);
and U1219 (N_1219,N_894,N_1013);
nor U1220 (N_1220,N_1028,N_1021);
and U1221 (N_1221,N_718,N_425);
nand U1222 (N_1222,N_886,N_1041);
and U1223 (N_1223,N_1111,N_1011);
and U1224 (N_1224,N_1004,N_825);
nor U1225 (N_1225,N_178,N_213);
and U1226 (N_1226,In_211,In_1266);
nor U1227 (N_1227,N_1106,N_1014);
nand U1228 (N_1228,N_799,N_1070);
nand U1229 (N_1229,N_500,N_683);
nand U1230 (N_1230,N_736,In_387);
and U1231 (N_1231,N_624,N_646);
xnor U1232 (N_1232,N_958,N_784);
xor U1233 (N_1233,N_916,N_1009);
or U1234 (N_1234,In_1363,In_1112);
and U1235 (N_1235,In_350,N_1033);
nand U1236 (N_1236,N_796,N_1122);
xor U1237 (N_1237,In_564,N_1096);
and U1238 (N_1238,N_765,In_1072);
or U1239 (N_1239,N_1005,N_459);
xnor U1240 (N_1240,N_771,In_1452);
or U1241 (N_1241,N_936,N_1110);
xnor U1242 (N_1242,N_883,N_761);
or U1243 (N_1243,N_989,N_710);
nand U1244 (N_1244,N_1092,N_841);
or U1245 (N_1245,N_687,N_1027);
and U1246 (N_1246,N_1078,N_244);
xor U1247 (N_1247,N_1065,In_445);
nor U1248 (N_1248,In_729,N_937);
nand U1249 (N_1249,In_1020,N_563);
or U1250 (N_1250,In_817,N_512);
nand U1251 (N_1251,N_1146,N_987);
xnor U1252 (N_1252,N_318,N_1165);
and U1253 (N_1253,N_1196,N_1121);
and U1254 (N_1254,N_660,N_1167);
nor U1255 (N_1255,N_1148,N_1052);
xnor U1256 (N_1256,N_1181,N_1189);
and U1257 (N_1257,N_1116,N_1166);
xor U1258 (N_1258,In_1108,N_1185);
and U1259 (N_1259,N_635,N_1153);
xnor U1260 (N_1260,N_1098,N_1131);
nor U1261 (N_1261,N_1164,In_661);
or U1262 (N_1262,N_711,N_1221);
xnor U1263 (N_1263,N_1249,N_1203);
nand U1264 (N_1264,In_377,N_598);
xor U1265 (N_1265,In_38,N_1201);
or U1266 (N_1266,N_1010,N_1206);
nor U1267 (N_1267,N_1183,N_1209);
nand U1268 (N_1268,N_1202,N_558);
xor U1269 (N_1269,N_1133,N_919);
or U1270 (N_1270,N_447,N_1225);
nand U1271 (N_1271,N_1095,N_1007);
xor U1272 (N_1272,N_722,N_1195);
nand U1273 (N_1273,N_104,N_1223);
or U1274 (N_1274,N_1228,N_1219);
or U1275 (N_1275,N_408,N_973);
nand U1276 (N_1276,N_903,N_705);
or U1277 (N_1277,N_871,N_1140);
nand U1278 (N_1278,N_1171,N_1241);
nand U1279 (N_1279,N_772,N_1075);
nand U1280 (N_1280,N_1192,N_1242);
and U1281 (N_1281,In_570,N_1193);
nand U1282 (N_1282,N_1245,N_1176);
nor U1283 (N_1283,N_742,N_554);
or U1284 (N_1284,N_1162,N_995);
and U1285 (N_1285,N_1243,N_928);
or U1286 (N_1286,N_513,N_719);
or U1287 (N_1287,N_1002,N_1136);
or U1288 (N_1288,In_831,N_656);
nand U1289 (N_1289,In_469,N_1208);
and U1290 (N_1290,N_1128,N_1069);
or U1291 (N_1291,N_1112,N_1233);
xnor U1292 (N_1292,N_1099,In_867);
or U1293 (N_1293,N_909,N_1220);
nor U1294 (N_1294,N_728,N_956);
xnor U1295 (N_1295,N_1180,In_1442);
nand U1296 (N_1296,N_880,N_875);
and U1297 (N_1297,N_1044,N_1147);
or U1298 (N_1298,N_1210,N_1175);
xnor U1299 (N_1299,N_963,N_715);
nor U1300 (N_1300,N_1214,N_1229);
or U1301 (N_1301,In_1117,N_1151);
nand U1302 (N_1302,N_1191,N_1159);
nor U1303 (N_1303,N_1152,N_1205);
nor U1304 (N_1304,In_1384,N_1145);
xnor U1305 (N_1305,In_463,N_943);
xor U1306 (N_1306,N_1246,N_751);
and U1307 (N_1307,N_1182,N_1178);
nor U1308 (N_1308,N_1124,N_962);
or U1309 (N_1309,N_1042,N_1198);
or U1310 (N_1310,N_1134,N_836);
xnor U1311 (N_1311,N_1187,N_770);
nor U1312 (N_1312,N_1017,N_1248);
or U1313 (N_1313,N_1163,N_1212);
and U1314 (N_1314,N_1238,N_1200);
xor U1315 (N_1315,In_87,N_860);
nand U1316 (N_1316,N_1217,N_1155);
and U1317 (N_1317,N_1215,N_1057);
xnor U1318 (N_1318,N_1226,N_1053);
or U1319 (N_1319,N_1172,N_976);
and U1320 (N_1320,N_921,N_1038);
nor U1321 (N_1321,In_1369,N_974);
and U1322 (N_1322,N_924,N_1135);
xnor U1323 (N_1323,N_1247,N_1125);
nand U1324 (N_1324,N_1170,N_1230);
xor U1325 (N_1325,N_1104,N_1030);
or U1326 (N_1326,N_1169,N_1127);
nand U1327 (N_1327,N_577,N_1186);
or U1328 (N_1328,N_1023,N_1188);
xnor U1329 (N_1329,In_1457,N_1137);
or U1330 (N_1330,N_1199,N_621);
nor U1331 (N_1331,N_1150,N_1236);
and U1332 (N_1332,In_655,N_1244);
nand U1333 (N_1333,N_888,N_1179);
nand U1334 (N_1334,In_553,N_1138);
and U1335 (N_1335,In_1050,N_1126);
or U1336 (N_1336,N_1234,N_1168);
or U1337 (N_1337,N_1160,N_1239);
nor U1338 (N_1338,N_239,N_1107);
xor U1339 (N_1339,N_1082,N_1213);
and U1340 (N_1340,N_471,N_1149);
and U1341 (N_1341,N_421,N_1060);
nand U1342 (N_1342,N_938,N_1222);
nand U1343 (N_1343,N_1144,N_643);
or U1344 (N_1344,N_590,N_1156);
or U1345 (N_1345,N_1204,N_1232);
and U1346 (N_1346,N_1068,N_1141);
and U1347 (N_1347,N_1240,N_1161);
nand U1348 (N_1348,N_1197,N_1142);
or U1349 (N_1349,N_1083,N_1130);
nor U1350 (N_1350,N_568,In_536);
and U1351 (N_1351,N_695,N_1211);
nor U1352 (N_1352,N_786,N_420);
nor U1353 (N_1353,N_930,N_1079);
nand U1354 (N_1354,N_934,N_1224);
and U1355 (N_1355,N_1173,N_966);
and U1356 (N_1356,N_1231,N_1055);
xor U1357 (N_1357,N_1132,In_1064);
and U1358 (N_1358,N_1117,N_1119);
xor U1359 (N_1359,N_483,N_1129);
and U1360 (N_1360,N_1154,N_1194);
xor U1361 (N_1361,N_1158,N_1064);
nor U1362 (N_1362,N_1139,N_1237);
nand U1363 (N_1363,N_1048,N_954);
nand U1364 (N_1364,N_1020,N_1109);
and U1365 (N_1365,In_263,N_1074);
nand U1366 (N_1366,N_1019,N_1218);
nor U1367 (N_1367,N_1235,N_1143);
nand U1368 (N_1368,N_522,In_1152);
xor U1369 (N_1369,N_1227,N_1216);
nor U1370 (N_1370,N_1177,N_340);
nand U1371 (N_1371,N_407,N_1190);
nand U1372 (N_1372,In_1037,N_1207);
xnor U1373 (N_1373,N_1157,N_1174);
xnor U1374 (N_1374,N_1184,N_1024);
xnor U1375 (N_1375,N_1324,N_1319);
nor U1376 (N_1376,N_1276,N_1351);
nor U1377 (N_1377,N_1315,N_1290);
nand U1378 (N_1378,N_1298,N_1286);
and U1379 (N_1379,N_1312,N_1305);
or U1380 (N_1380,N_1355,N_1364);
and U1381 (N_1381,N_1283,N_1367);
nand U1382 (N_1382,N_1326,N_1264);
nor U1383 (N_1383,N_1320,N_1262);
nor U1384 (N_1384,N_1259,N_1346);
xnor U1385 (N_1385,N_1314,N_1357);
or U1386 (N_1386,N_1374,N_1363);
nand U1387 (N_1387,N_1253,N_1323);
and U1388 (N_1388,N_1352,N_1336);
xor U1389 (N_1389,N_1257,N_1269);
and U1390 (N_1390,N_1306,N_1339);
nor U1391 (N_1391,N_1282,N_1360);
nand U1392 (N_1392,N_1335,N_1349);
and U1393 (N_1393,N_1322,N_1293);
and U1394 (N_1394,N_1299,N_1288);
or U1395 (N_1395,N_1372,N_1342);
or U1396 (N_1396,N_1311,N_1278);
nand U1397 (N_1397,N_1369,N_1328);
nand U1398 (N_1398,N_1356,N_1341);
and U1399 (N_1399,N_1280,N_1317);
nand U1400 (N_1400,N_1272,N_1260);
and U1401 (N_1401,N_1258,N_1325);
or U1402 (N_1402,N_1294,N_1361);
nand U1403 (N_1403,N_1310,N_1337);
xor U1404 (N_1404,N_1295,N_1303);
or U1405 (N_1405,N_1291,N_1263);
nand U1406 (N_1406,N_1362,N_1365);
nand U1407 (N_1407,N_1345,N_1327);
or U1408 (N_1408,N_1251,N_1252);
and U1409 (N_1409,N_1302,N_1307);
and U1410 (N_1410,N_1309,N_1308);
or U1411 (N_1411,N_1340,N_1358);
or U1412 (N_1412,N_1347,N_1373);
and U1413 (N_1413,N_1370,N_1271);
xor U1414 (N_1414,N_1292,N_1332);
xnor U1415 (N_1415,N_1277,N_1256);
or U1416 (N_1416,N_1297,N_1343);
xor U1417 (N_1417,N_1254,N_1338);
nand U1418 (N_1418,N_1274,N_1250);
xor U1419 (N_1419,N_1348,N_1270);
nor U1420 (N_1420,N_1261,N_1279);
nor U1421 (N_1421,N_1366,N_1344);
xnor U1422 (N_1422,N_1316,N_1368);
nand U1423 (N_1423,N_1371,N_1359);
nor U1424 (N_1424,N_1273,N_1287);
nor U1425 (N_1425,N_1313,N_1284);
nor U1426 (N_1426,N_1329,N_1318);
or U1427 (N_1427,N_1289,N_1304);
nand U1428 (N_1428,N_1353,N_1255);
nand U1429 (N_1429,N_1266,N_1265);
or U1430 (N_1430,N_1354,N_1281);
and U1431 (N_1431,N_1296,N_1275);
nand U1432 (N_1432,N_1331,N_1268);
or U1433 (N_1433,N_1350,N_1267);
nand U1434 (N_1434,N_1330,N_1300);
or U1435 (N_1435,N_1285,N_1334);
or U1436 (N_1436,N_1333,N_1301);
nand U1437 (N_1437,N_1321,N_1259);
or U1438 (N_1438,N_1335,N_1267);
xor U1439 (N_1439,N_1253,N_1295);
and U1440 (N_1440,N_1320,N_1354);
nor U1441 (N_1441,N_1334,N_1255);
or U1442 (N_1442,N_1266,N_1282);
nand U1443 (N_1443,N_1341,N_1268);
or U1444 (N_1444,N_1302,N_1266);
xor U1445 (N_1445,N_1272,N_1340);
or U1446 (N_1446,N_1286,N_1267);
nor U1447 (N_1447,N_1319,N_1261);
and U1448 (N_1448,N_1291,N_1363);
nand U1449 (N_1449,N_1290,N_1285);
and U1450 (N_1450,N_1322,N_1330);
and U1451 (N_1451,N_1288,N_1262);
nor U1452 (N_1452,N_1301,N_1330);
and U1453 (N_1453,N_1300,N_1313);
or U1454 (N_1454,N_1269,N_1253);
and U1455 (N_1455,N_1358,N_1368);
xnor U1456 (N_1456,N_1306,N_1287);
and U1457 (N_1457,N_1374,N_1269);
or U1458 (N_1458,N_1253,N_1345);
and U1459 (N_1459,N_1252,N_1291);
nor U1460 (N_1460,N_1358,N_1300);
nand U1461 (N_1461,N_1335,N_1336);
nor U1462 (N_1462,N_1317,N_1372);
nand U1463 (N_1463,N_1284,N_1346);
nand U1464 (N_1464,N_1339,N_1368);
and U1465 (N_1465,N_1259,N_1341);
xor U1466 (N_1466,N_1270,N_1250);
nor U1467 (N_1467,N_1270,N_1321);
nand U1468 (N_1468,N_1257,N_1251);
xnor U1469 (N_1469,N_1273,N_1257);
nor U1470 (N_1470,N_1273,N_1349);
nor U1471 (N_1471,N_1324,N_1267);
or U1472 (N_1472,N_1256,N_1253);
nand U1473 (N_1473,N_1268,N_1288);
and U1474 (N_1474,N_1298,N_1301);
nor U1475 (N_1475,N_1332,N_1342);
or U1476 (N_1476,N_1275,N_1255);
and U1477 (N_1477,N_1255,N_1308);
nor U1478 (N_1478,N_1374,N_1304);
xor U1479 (N_1479,N_1256,N_1314);
and U1480 (N_1480,N_1276,N_1257);
nor U1481 (N_1481,N_1324,N_1269);
and U1482 (N_1482,N_1300,N_1362);
or U1483 (N_1483,N_1285,N_1336);
nor U1484 (N_1484,N_1349,N_1253);
xor U1485 (N_1485,N_1312,N_1358);
nand U1486 (N_1486,N_1298,N_1350);
xor U1487 (N_1487,N_1372,N_1297);
and U1488 (N_1488,N_1314,N_1293);
or U1489 (N_1489,N_1311,N_1331);
and U1490 (N_1490,N_1331,N_1271);
nor U1491 (N_1491,N_1256,N_1283);
nor U1492 (N_1492,N_1361,N_1254);
or U1493 (N_1493,N_1273,N_1295);
and U1494 (N_1494,N_1289,N_1309);
xnor U1495 (N_1495,N_1337,N_1360);
nand U1496 (N_1496,N_1308,N_1266);
xor U1497 (N_1497,N_1332,N_1254);
xor U1498 (N_1498,N_1267,N_1348);
or U1499 (N_1499,N_1336,N_1262);
nor U1500 (N_1500,N_1468,N_1404);
nand U1501 (N_1501,N_1463,N_1484);
and U1502 (N_1502,N_1453,N_1469);
xnor U1503 (N_1503,N_1486,N_1415);
or U1504 (N_1504,N_1487,N_1481);
or U1505 (N_1505,N_1428,N_1459);
or U1506 (N_1506,N_1457,N_1400);
and U1507 (N_1507,N_1375,N_1399);
or U1508 (N_1508,N_1498,N_1420);
nand U1509 (N_1509,N_1394,N_1437);
nor U1510 (N_1510,N_1402,N_1467);
nand U1511 (N_1511,N_1451,N_1376);
xor U1512 (N_1512,N_1377,N_1477);
xnor U1513 (N_1513,N_1378,N_1452);
xor U1514 (N_1514,N_1413,N_1390);
and U1515 (N_1515,N_1466,N_1393);
nand U1516 (N_1516,N_1429,N_1492);
xnor U1517 (N_1517,N_1499,N_1403);
nor U1518 (N_1518,N_1408,N_1462);
xor U1519 (N_1519,N_1485,N_1455);
nor U1520 (N_1520,N_1436,N_1406);
nor U1521 (N_1521,N_1454,N_1475);
nand U1522 (N_1522,N_1379,N_1401);
nand U1523 (N_1523,N_1411,N_1490);
xnor U1524 (N_1524,N_1471,N_1479);
nand U1525 (N_1525,N_1389,N_1495);
nor U1526 (N_1526,N_1494,N_1434);
nand U1527 (N_1527,N_1439,N_1419);
and U1528 (N_1528,N_1423,N_1438);
or U1529 (N_1529,N_1398,N_1470);
xor U1530 (N_1530,N_1396,N_1387);
xor U1531 (N_1531,N_1458,N_1473);
xnor U1532 (N_1532,N_1497,N_1493);
or U1533 (N_1533,N_1380,N_1480);
xnor U1534 (N_1534,N_1442,N_1407);
nor U1535 (N_1535,N_1465,N_1381);
xor U1536 (N_1536,N_1388,N_1446);
nand U1537 (N_1537,N_1405,N_1488);
nor U1538 (N_1538,N_1464,N_1392);
xnor U1539 (N_1539,N_1421,N_1412);
xnor U1540 (N_1540,N_1382,N_1426);
nand U1541 (N_1541,N_1417,N_1476);
nor U1542 (N_1542,N_1416,N_1409);
and U1543 (N_1543,N_1496,N_1425);
and U1544 (N_1544,N_1448,N_1424);
and U1545 (N_1545,N_1489,N_1483);
or U1546 (N_1546,N_1385,N_1456);
or U1547 (N_1547,N_1450,N_1478);
xor U1548 (N_1548,N_1443,N_1461);
xor U1549 (N_1549,N_1441,N_1386);
or U1550 (N_1550,N_1395,N_1491);
nand U1551 (N_1551,N_1384,N_1422);
nand U1552 (N_1552,N_1433,N_1472);
nor U1553 (N_1553,N_1430,N_1410);
or U1554 (N_1554,N_1440,N_1435);
nor U1555 (N_1555,N_1482,N_1427);
and U1556 (N_1556,N_1445,N_1432);
and U1557 (N_1557,N_1431,N_1418);
nor U1558 (N_1558,N_1397,N_1383);
nor U1559 (N_1559,N_1391,N_1460);
and U1560 (N_1560,N_1447,N_1414);
and U1561 (N_1561,N_1474,N_1449);
or U1562 (N_1562,N_1444,N_1382);
and U1563 (N_1563,N_1487,N_1477);
and U1564 (N_1564,N_1378,N_1464);
nor U1565 (N_1565,N_1461,N_1460);
nor U1566 (N_1566,N_1462,N_1459);
xnor U1567 (N_1567,N_1380,N_1436);
nor U1568 (N_1568,N_1377,N_1479);
or U1569 (N_1569,N_1437,N_1458);
or U1570 (N_1570,N_1411,N_1382);
nor U1571 (N_1571,N_1481,N_1405);
nor U1572 (N_1572,N_1375,N_1412);
nand U1573 (N_1573,N_1403,N_1446);
nor U1574 (N_1574,N_1440,N_1394);
xnor U1575 (N_1575,N_1433,N_1440);
and U1576 (N_1576,N_1394,N_1460);
xor U1577 (N_1577,N_1440,N_1432);
xnor U1578 (N_1578,N_1490,N_1409);
and U1579 (N_1579,N_1436,N_1473);
and U1580 (N_1580,N_1453,N_1496);
and U1581 (N_1581,N_1390,N_1445);
and U1582 (N_1582,N_1439,N_1474);
xor U1583 (N_1583,N_1413,N_1477);
or U1584 (N_1584,N_1425,N_1470);
nor U1585 (N_1585,N_1430,N_1415);
nand U1586 (N_1586,N_1385,N_1403);
nand U1587 (N_1587,N_1462,N_1456);
xnor U1588 (N_1588,N_1449,N_1466);
nand U1589 (N_1589,N_1387,N_1407);
xnor U1590 (N_1590,N_1442,N_1417);
xor U1591 (N_1591,N_1469,N_1379);
nor U1592 (N_1592,N_1470,N_1385);
nor U1593 (N_1593,N_1375,N_1426);
nand U1594 (N_1594,N_1462,N_1484);
or U1595 (N_1595,N_1462,N_1485);
nand U1596 (N_1596,N_1426,N_1433);
nor U1597 (N_1597,N_1377,N_1452);
nor U1598 (N_1598,N_1472,N_1488);
or U1599 (N_1599,N_1409,N_1394);
and U1600 (N_1600,N_1485,N_1380);
nand U1601 (N_1601,N_1420,N_1413);
nor U1602 (N_1602,N_1394,N_1475);
and U1603 (N_1603,N_1404,N_1477);
and U1604 (N_1604,N_1415,N_1409);
nand U1605 (N_1605,N_1432,N_1489);
xnor U1606 (N_1606,N_1391,N_1482);
nand U1607 (N_1607,N_1390,N_1397);
xnor U1608 (N_1608,N_1465,N_1456);
nor U1609 (N_1609,N_1469,N_1436);
xor U1610 (N_1610,N_1451,N_1379);
or U1611 (N_1611,N_1375,N_1387);
or U1612 (N_1612,N_1493,N_1402);
and U1613 (N_1613,N_1452,N_1420);
xnor U1614 (N_1614,N_1392,N_1440);
xor U1615 (N_1615,N_1482,N_1492);
nand U1616 (N_1616,N_1396,N_1386);
xor U1617 (N_1617,N_1481,N_1378);
xnor U1618 (N_1618,N_1389,N_1492);
nor U1619 (N_1619,N_1468,N_1459);
nand U1620 (N_1620,N_1387,N_1403);
or U1621 (N_1621,N_1386,N_1444);
nand U1622 (N_1622,N_1397,N_1382);
and U1623 (N_1623,N_1492,N_1441);
xnor U1624 (N_1624,N_1456,N_1495);
and U1625 (N_1625,N_1565,N_1510);
nand U1626 (N_1626,N_1582,N_1544);
xnor U1627 (N_1627,N_1614,N_1542);
nor U1628 (N_1628,N_1599,N_1509);
nor U1629 (N_1629,N_1535,N_1557);
and U1630 (N_1630,N_1527,N_1517);
nor U1631 (N_1631,N_1567,N_1585);
nand U1632 (N_1632,N_1613,N_1564);
nand U1633 (N_1633,N_1571,N_1578);
nand U1634 (N_1634,N_1529,N_1522);
and U1635 (N_1635,N_1577,N_1556);
nand U1636 (N_1636,N_1562,N_1568);
and U1637 (N_1637,N_1507,N_1570);
or U1638 (N_1638,N_1615,N_1597);
nor U1639 (N_1639,N_1587,N_1505);
xnor U1640 (N_1640,N_1551,N_1576);
xor U1641 (N_1641,N_1539,N_1596);
or U1642 (N_1642,N_1500,N_1612);
or U1643 (N_1643,N_1574,N_1524);
nand U1644 (N_1644,N_1501,N_1594);
xor U1645 (N_1645,N_1561,N_1607);
nor U1646 (N_1646,N_1516,N_1519);
nand U1647 (N_1647,N_1560,N_1555);
nor U1648 (N_1648,N_1604,N_1533);
nor U1649 (N_1649,N_1518,N_1502);
or U1650 (N_1650,N_1546,N_1595);
and U1651 (N_1651,N_1521,N_1549);
and U1652 (N_1652,N_1559,N_1558);
or U1653 (N_1653,N_1623,N_1508);
nor U1654 (N_1654,N_1554,N_1603);
nor U1655 (N_1655,N_1622,N_1563);
or U1656 (N_1656,N_1601,N_1515);
and U1657 (N_1657,N_1534,N_1608);
or U1658 (N_1658,N_1569,N_1616);
nor U1659 (N_1659,N_1620,N_1605);
or U1660 (N_1660,N_1621,N_1543);
nor U1661 (N_1661,N_1511,N_1504);
and U1662 (N_1662,N_1624,N_1579);
or U1663 (N_1663,N_1617,N_1586);
nand U1664 (N_1664,N_1580,N_1589);
nor U1665 (N_1665,N_1583,N_1618);
or U1666 (N_1666,N_1520,N_1592);
nand U1667 (N_1667,N_1513,N_1506);
or U1668 (N_1668,N_1610,N_1611);
nand U1669 (N_1669,N_1552,N_1591);
and U1670 (N_1670,N_1530,N_1600);
nor U1671 (N_1671,N_1526,N_1514);
xnor U1672 (N_1672,N_1523,N_1609);
nor U1673 (N_1673,N_1572,N_1619);
and U1674 (N_1674,N_1536,N_1538);
nand U1675 (N_1675,N_1553,N_1531);
nand U1676 (N_1676,N_1545,N_1540);
nor U1677 (N_1677,N_1503,N_1548);
xor U1678 (N_1678,N_1512,N_1532);
and U1679 (N_1679,N_1550,N_1528);
xor U1680 (N_1680,N_1573,N_1598);
xnor U1681 (N_1681,N_1602,N_1547);
xor U1682 (N_1682,N_1588,N_1590);
or U1683 (N_1683,N_1581,N_1606);
or U1684 (N_1684,N_1584,N_1575);
xor U1685 (N_1685,N_1537,N_1525);
or U1686 (N_1686,N_1593,N_1566);
xor U1687 (N_1687,N_1541,N_1570);
nand U1688 (N_1688,N_1622,N_1559);
and U1689 (N_1689,N_1524,N_1595);
and U1690 (N_1690,N_1562,N_1558);
and U1691 (N_1691,N_1547,N_1531);
nor U1692 (N_1692,N_1582,N_1511);
xnor U1693 (N_1693,N_1524,N_1577);
and U1694 (N_1694,N_1600,N_1521);
nor U1695 (N_1695,N_1541,N_1551);
nor U1696 (N_1696,N_1624,N_1559);
nor U1697 (N_1697,N_1515,N_1525);
or U1698 (N_1698,N_1582,N_1545);
and U1699 (N_1699,N_1574,N_1591);
or U1700 (N_1700,N_1549,N_1569);
and U1701 (N_1701,N_1588,N_1535);
nand U1702 (N_1702,N_1586,N_1578);
nand U1703 (N_1703,N_1573,N_1538);
nor U1704 (N_1704,N_1556,N_1553);
and U1705 (N_1705,N_1502,N_1572);
or U1706 (N_1706,N_1620,N_1618);
xor U1707 (N_1707,N_1516,N_1527);
nor U1708 (N_1708,N_1559,N_1540);
nor U1709 (N_1709,N_1553,N_1615);
or U1710 (N_1710,N_1576,N_1575);
and U1711 (N_1711,N_1537,N_1501);
nand U1712 (N_1712,N_1572,N_1570);
and U1713 (N_1713,N_1570,N_1566);
and U1714 (N_1714,N_1548,N_1541);
or U1715 (N_1715,N_1552,N_1539);
xnor U1716 (N_1716,N_1547,N_1612);
xor U1717 (N_1717,N_1613,N_1502);
nor U1718 (N_1718,N_1544,N_1548);
or U1719 (N_1719,N_1576,N_1605);
and U1720 (N_1720,N_1517,N_1604);
xnor U1721 (N_1721,N_1588,N_1598);
or U1722 (N_1722,N_1581,N_1505);
or U1723 (N_1723,N_1594,N_1623);
nor U1724 (N_1724,N_1542,N_1586);
or U1725 (N_1725,N_1619,N_1550);
and U1726 (N_1726,N_1520,N_1576);
xnor U1727 (N_1727,N_1556,N_1559);
and U1728 (N_1728,N_1547,N_1624);
nor U1729 (N_1729,N_1535,N_1517);
or U1730 (N_1730,N_1530,N_1540);
xnor U1731 (N_1731,N_1534,N_1612);
nor U1732 (N_1732,N_1530,N_1611);
nor U1733 (N_1733,N_1622,N_1570);
xnor U1734 (N_1734,N_1565,N_1574);
and U1735 (N_1735,N_1602,N_1601);
nor U1736 (N_1736,N_1605,N_1595);
nand U1737 (N_1737,N_1568,N_1597);
nand U1738 (N_1738,N_1610,N_1520);
or U1739 (N_1739,N_1562,N_1544);
or U1740 (N_1740,N_1536,N_1559);
nand U1741 (N_1741,N_1579,N_1576);
nor U1742 (N_1742,N_1580,N_1570);
xnor U1743 (N_1743,N_1589,N_1603);
or U1744 (N_1744,N_1575,N_1593);
or U1745 (N_1745,N_1609,N_1595);
xnor U1746 (N_1746,N_1623,N_1607);
xor U1747 (N_1747,N_1515,N_1534);
xor U1748 (N_1748,N_1581,N_1617);
and U1749 (N_1749,N_1539,N_1514);
and U1750 (N_1750,N_1743,N_1632);
and U1751 (N_1751,N_1711,N_1652);
or U1752 (N_1752,N_1641,N_1684);
xor U1753 (N_1753,N_1629,N_1631);
xnor U1754 (N_1754,N_1659,N_1681);
or U1755 (N_1755,N_1643,N_1680);
nor U1756 (N_1756,N_1710,N_1688);
and U1757 (N_1757,N_1661,N_1747);
or U1758 (N_1758,N_1731,N_1739);
and U1759 (N_1759,N_1742,N_1720);
and U1760 (N_1760,N_1634,N_1704);
nor U1761 (N_1761,N_1638,N_1705);
or U1762 (N_1762,N_1683,N_1734);
or U1763 (N_1763,N_1698,N_1708);
or U1764 (N_1764,N_1713,N_1662);
or U1765 (N_1765,N_1671,N_1678);
nor U1766 (N_1766,N_1650,N_1706);
nand U1767 (N_1767,N_1696,N_1700);
nand U1768 (N_1768,N_1729,N_1679);
and U1769 (N_1769,N_1635,N_1727);
or U1770 (N_1770,N_1689,N_1626);
xnor U1771 (N_1771,N_1745,N_1695);
xnor U1772 (N_1772,N_1721,N_1663);
nand U1773 (N_1773,N_1664,N_1633);
or U1774 (N_1774,N_1646,N_1716);
and U1775 (N_1775,N_1744,N_1674);
nor U1776 (N_1776,N_1737,N_1738);
and U1777 (N_1777,N_1670,N_1675);
nor U1778 (N_1778,N_1707,N_1717);
or U1779 (N_1779,N_1668,N_1697);
or U1780 (N_1780,N_1709,N_1636);
nor U1781 (N_1781,N_1667,N_1642);
and U1782 (N_1782,N_1677,N_1723);
nor U1783 (N_1783,N_1628,N_1669);
nor U1784 (N_1784,N_1736,N_1653);
nand U1785 (N_1785,N_1699,N_1749);
nand U1786 (N_1786,N_1733,N_1748);
or U1787 (N_1787,N_1637,N_1728);
and U1788 (N_1788,N_1644,N_1703);
xnor U1789 (N_1789,N_1645,N_1682);
xor U1790 (N_1790,N_1655,N_1724);
xor U1791 (N_1791,N_1686,N_1725);
nor U1792 (N_1792,N_1740,N_1693);
and U1793 (N_1793,N_1702,N_1647);
and U1794 (N_1794,N_1691,N_1657);
nor U1795 (N_1795,N_1654,N_1651);
nand U1796 (N_1796,N_1639,N_1715);
xor U1797 (N_1797,N_1719,N_1656);
nor U1798 (N_1798,N_1648,N_1625);
and U1799 (N_1799,N_1687,N_1627);
or U1800 (N_1800,N_1741,N_1735);
xor U1801 (N_1801,N_1673,N_1630);
or U1802 (N_1802,N_1694,N_1722);
or U1803 (N_1803,N_1692,N_1640);
or U1804 (N_1804,N_1718,N_1665);
nand U1805 (N_1805,N_1672,N_1666);
nand U1806 (N_1806,N_1746,N_1712);
nor U1807 (N_1807,N_1701,N_1658);
nor U1808 (N_1808,N_1690,N_1676);
xor U1809 (N_1809,N_1685,N_1649);
nand U1810 (N_1810,N_1660,N_1730);
xor U1811 (N_1811,N_1732,N_1714);
or U1812 (N_1812,N_1726,N_1708);
nand U1813 (N_1813,N_1693,N_1640);
nand U1814 (N_1814,N_1731,N_1651);
nand U1815 (N_1815,N_1651,N_1748);
and U1816 (N_1816,N_1672,N_1731);
nand U1817 (N_1817,N_1726,N_1738);
or U1818 (N_1818,N_1748,N_1740);
and U1819 (N_1819,N_1684,N_1656);
nor U1820 (N_1820,N_1719,N_1746);
xor U1821 (N_1821,N_1629,N_1637);
nor U1822 (N_1822,N_1724,N_1687);
or U1823 (N_1823,N_1688,N_1735);
nand U1824 (N_1824,N_1720,N_1680);
xor U1825 (N_1825,N_1714,N_1644);
xor U1826 (N_1826,N_1747,N_1705);
nand U1827 (N_1827,N_1641,N_1665);
or U1828 (N_1828,N_1712,N_1684);
nor U1829 (N_1829,N_1672,N_1746);
or U1830 (N_1830,N_1724,N_1740);
or U1831 (N_1831,N_1688,N_1641);
and U1832 (N_1832,N_1646,N_1730);
nand U1833 (N_1833,N_1652,N_1632);
xor U1834 (N_1834,N_1650,N_1698);
and U1835 (N_1835,N_1647,N_1691);
and U1836 (N_1836,N_1708,N_1713);
and U1837 (N_1837,N_1747,N_1691);
nor U1838 (N_1838,N_1725,N_1692);
nor U1839 (N_1839,N_1711,N_1715);
nor U1840 (N_1840,N_1714,N_1746);
and U1841 (N_1841,N_1749,N_1667);
nor U1842 (N_1842,N_1645,N_1725);
or U1843 (N_1843,N_1695,N_1699);
or U1844 (N_1844,N_1717,N_1670);
nand U1845 (N_1845,N_1724,N_1653);
and U1846 (N_1846,N_1657,N_1739);
and U1847 (N_1847,N_1729,N_1675);
or U1848 (N_1848,N_1733,N_1646);
nor U1849 (N_1849,N_1744,N_1714);
nand U1850 (N_1850,N_1744,N_1676);
or U1851 (N_1851,N_1727,N_1732);
nand U1852 (N_1852,N_1645,N_1742);
nor U1853 (N_1853,N_1643,N_1718);
nor U1854 (N_1854,N_1706,N_1626);
or U1855 (N_1855,N_1748,N_1743);
nor U1856 (N_1856,N_1704,N_1635);
nand U1857 (N_1857,N_1739,N_1649);
nand U1858 (N_1858,N_1719,N_1731);
and U1859 (N_1859,N_1629,N_1732);
xor U1860 (N_1860,N_1695,N_1689);
nand U1861 (N_1861,N_1684,N_1673);
xnor U1862 (N_1862,N_1631,N_1677);
or U1863 (N_1863,N_1732,N_1668);
xnor U1864 (N_1864,N_1746,N_1631);
and U1865 (N_1865,N_1721,N_1727);
xnor U1866 (N_1866,N_1711,N_1661);
xnor U1867 (N_1867,N_1692,N_1727);
and U1868 (N_1868,N_1749,N_1670);
xnor U1869 (N_1869,N_1749,N_1660);
or U1870 (N_1870,N_1670,N_1705);
and U1871 (N_1871,N_1663,N_1678);
and U1872 (N_1872,N_1712,N_1656);
nor U1873 (N_1873,N_1740,N_1734);
or U1874 (N_1874,N_1692,N_1746);
nand U1875 (N_1875,N_1764,N_1807);
nand U1876 (N_1876,N_1751,N_1799);
nor U1877 (N_1877,N_1857,N_1814);
and U1878 (N_1878,N_1833,N_1798);
or U1879 (N_1879,N_1817,N_1874);
and U1880 (N_1880,N_1841,N_1860);
or U1881 (N_1881,N_1856,N_1791);
nor U1882 (N_1882,N_1773,N_1818);
or U1883 (N_1883,N_1853,N_1835);
or U1884 (N_1884,N_1753,N_1840);
nor U1885 (N_1885,N_1863,N_1866);
nand U1886 (N_1886,N_1865,N_1846);
and U1887 (N_1887,N_1816,N_1766);
xor U1888 (N_1888,N_1768,N_1824);
nor U1889 (N_1889,N_1765,N_1858);
nand U1890 (N_1890,N_1792,N_1771);
nand U1891 (N_1891,N_1762,N_1830);
or U1892 (N_1892,N_1870,N_1794);
and U1893 (N_1893,N_1848,N_1843);
and U1894 (N_1894,N_1793,N_1781);
xor U1895 (N_1895,N_1810,N_1752);
or U1896 (N_1896,N_1850,N_1871);
or U1897 (N_1897,N_1769,N_1813);
nand U1898 (N_1898,N_1789,N_1786);
xor U1899 (N_1899,N_1782,N_1779);
and U1900 (N_1900,N_1855,N_1770);
xor U1901 (N_1901,N_1821,N_1826);
and U1902 (N_1902,N_1754,N_1800);
xnor U1903 (N_1903,N_1873,N_1758);
and U1904 (N_1904,N_1759,N_1805);
nand U1905 (N_1905,N_1829,N_1760);
nor U1906 (N_1906,N_1838,N_1811);
nand U1907 (N_1907,N_1862,N_1774);
nand U1908 (N_1908,N_1820,N_1859);
nand U1909 (N_1909,N_1822,N_1778);
or U1910 (N_1910,N_1797,N_1832);
nand U1911 (N_1911,N_1849,N_1834);
and U1912 (N_1912,N_1823,N_1819);
nor U1913 (N_1913,N_1802,N_1845);
and U1914 (N_1914,N_1790,N_1756);
xnor U1915 (N_1915,N_1825,N_1812);
or U1916 (N_1916,N_1868,N_1785);
nor U1917 (N_1917,N_1872,N_1796);
xor U1918 (N_1918,N_1803,N_1777);
nor U1919 (N_1919,N_1784,N_1767);
xor U1920 (N_1920,N_1763,N_1795);
xor U1921 (N_1921,N_1801,N_1755);
nor U1922 (N_1922,N_1827,N_1806);
and U1923 (N_1923,N_1772,N_1836);
nand U1924 (N_1924,N_1788,N_1847);
and U1925 (N_1925,N_1815,N_1828);
or U1926 (N_1926,N_1780,N_1809);
nor U1927 (N_1927,N_1831,N_1750);
xnor U1928 (N_1928,N_1854,N_1869);
xnor U1929 (N_1929,N_1839,N_1787);
xor U1930 (N_1930,N_1808,N_1852);
nand U1931 (N_1931,N_1861,N_1864);
or U1932 (N_1932,N_1844,N_1776);
nand U1933 (N_1933,N_1842,N_1837);
and U1934 (N_1934,N_1867,N_1851);
nand U1935 (N_1935,N_1804,N_1775);
nor U1936 (N_1936,N_1761,N_1783);
and U1937 (N_1937,N_1757,N_1855);
nor U1938 (N_1938,N_1867,N_1837);
nor U1939 (N_1939,N_1789,N_1858);
nand U1940 (N_1940,N_1871,N_1802);
nand U1941 (N_1941,N_1817,N_1831);
or U1942 (N_1942,N_1800,N_1815);
and U1943 (N_1943,N_1816,N_1821);
and U1944 (N_1944,N_1844,N_1771);
nand U1945 (N_1945,N_1814,N_1870);
and U1946 (N_1946,N_1800,N_1811);
xnor U1947 (N_1947,N_1792,N_1838);
or U1948 (N_1948,N_1757,N_1859);
nand U1949 (N_1949,N_1866,N_1760);
and U1950 (N_1950,N_1846,N_1870);
nor U1951 (N_1951,N_1824,N_1858);
nand U1952 (N_1952,N_1751,N_1845);
and U1953 (N_1953,N_1835,N_1845);
or U1954 (N_1954,N_1846,N_1763);
xnor U1955 (N_1955,N_1835,N_1866);
or U1956 (N_1956,N_1765,N_1805);
nor U1957 (N_1957,N_1756,N_1800);
xnor U1958 (N_1958,N_1814,N_1799);
nor U1959 (N_1959,N_1800,N_1804);
xor U1960 (N_1960,N_1821,N_1861);
and U1961 (N_1961,N_1785,N_1810);
nand U1962 (N_1962,N_1837,N_1831);
and U1963 (N_1963,N_1774,N_1752);
and U1964 (N_1964,N_1830,N_1759);
nand U1965 (N_1965,N_1822,N_1814);
and U1966 (N_1966,N_1783,N_1772);
and U1967 (N_1967,N_1871,N_1771);
and U1968 (N_1968,N_1863,N_1813);
or U1969 (N_1969,N_1803,N_1774);
or U1970 (N_1970,N_1794,N_1825);
and U1971 (N_1971,N_1821,N_1762);
xor U1972 (N_1972,N_1800,N_1870);
nor U1973 (N_1973,N_1851,N_1815);
xnor U1974 (N_1974,N_1845,N_1830);
and U1975 (N_1975,N_1767,N_1850);
or U1976 (N_1976,N_1786,N_1767);
and U1977 (N_1977,N_1786,N_1757);
nor U1978 (N_1978,N_1776,N_1797);
or U1979 (N_1979,N_1764,N_1862);
xor U1980 (N_1980,N_1797,N_1813);
nand U1981 (N_1981,N_1845,N_1783);
nor U1982 (N_1982,N_1770,N_1862);
xor U1983 (N_1983,N_1766,N_1837);
nand U1984 (N_1984,N_1795,N_1841);
and U1985 (N_1985,N_1844,N_1821);
nand U1986 (N_1986,N_1792,N_1837);
or U1987 (N_1987,N_1771,N_1828);
nor U1988 (N_1988,N_1844,N_1850);
and U1989 (N_1989,N_1768,N_1825);
and U1990 (N_1990,N_1872,N_1821);
nand U1991 (N_1991,N_1830,N_1809);
and U1992 (N_1992,N_1757,N_1762);
and U1993 (N_1993,N_1770,N_1824);
nand U1994 (N_1994,N_1813,N_1808);
or U1995 (N_1995,N_1791,N_1861);
and U1996 (N_1996,N_1806,N_1809);
and U1997 (N_1997,N_1850,N_1867);
or U1998 (N_1998,N_1854,N_1799);
xnor U1999 (N_1999,N_1800,N_1784);
xnor U2000 (N_2000,N_1987,N_1954);
nor U2001 (N_2001,N_1880,N_1990);
or U2002 (N_2002,N_1995,N_1994);
nand U2003 (N_2003,N_1879,N_1882);
and U2004 (N_2004,N_1993,N_1940);
nand U2005 (N_2005,N_1889,N_1921);
nor U2006 (N_2006,N_1976,N_1953);
nor U2007 (N_2007,N_1896,N_1970);
nand U2008 (N_2008,N_1933,N_1936);
nand U2009 (N_2009,N_1965,N_1895);
xor U2010 (N_2010,N_1939,N_1900);
or U2011 (N_2011,N_1905,N_1916);
or U2012 (N_2012,N_1887,N_1988);
nand U2013 (N_2013,N_1922,N_1893);
and U2014 (N_2014,N_1952,N_1923);
xor U2015 (N_2015,N_1911,N_1972);
xor U2016 (N_2016,N_1992,N_1986);
xor U2017 (N_2017,N_1958,N_1985);
nor U2018 (N_2018,N_1943,N_1980);
xnor U2019 (N_2019,N_1915,N_1981);
nor U2020 (N_2020,N_1960,N_1912);
or U2021 (N_2021,N_1964,N_1901);
and U2022 (N_2022,N_1991,N_1903);
xor U2023 (N_2023,N_1956,N_1883);
and U2024 (N_2024,N_1897,N_1907);
nand U2025 (N_2025,N_1969,N_1941);
nor U2026 (N_2026,N_1934,N_1978);
nor U2027 (N_2027,N_1910,N_1917);
nand U2028 (N_2028,N_1959,N_1931);
nor U2029 (N_2029,N_1949,N_1928);
and U2030 (N_2030,N_1971,N_1982);
xor U2031 (N_2031,N_1902,N_1975);
nand U2032 (N_2032,N_1926,N_1894);
nand U2033 (N_2033,N_1918,N_1898);
nor U2034 (N_2034,N_1989,N_1957);
nand U2035 (N_2035,N_1877,N_1996);
or U2036 (N_2036,N_1909,N_1892);
and U2037 (N_2037,N_1950,N_1932);
nor U2038 (N_2038,N_1963,N_1913);
or U2039 (N_2039,N_1884,N_1920);
nand U2040 (N_2040,N_1924,N_1955);
or U2041 (N_2041,N_1962,N_1944);
nor U2042 (N_2042,N_1935,N_1997);
nor U2043 (N_2043,N_1974,N_1878);
and U2044 (N_2044,N_1937,N_1881);
nor U2045 (N_2045,N_1891,N_1906);
or U2046 (N_2046,N_1998,N_1886);
and U2047 (N_2047,N_1888,N_1876);
and U2048 (N_2048,N_1914,N_1930);
nor U2049 (N_2049,N_1925,N_1973);
nor U2050 (N_2050,N_1967,N_1961);
xnor U2051 (N_2051,N_1999,N_1890);
and U2052 (N_2052,N_1908,N_1875);
nand U2053 (N_2053,N_1904,N_1899);
and U2054 (N_2054,N_1885,N_1929);
or U2055 (N_2055,N_1938,N_1945);
nand U2056 (N_2056,N_1927,N_1947);
or U2057 (N_2057,N_1946,N_1948);
and U2058 (N_2058,N_1979,N_1983);
xor U2059 (N_2059,N_1984,N_1966);
nor U2060 (N_2060,N_1942,N_1919);
or U2061 (N_2061,N_1968,N_1977);
or U2062 (N_2062,N_1951,N_1898);
xnor U2063 (N_2063,N_1893,N_1980);
nand U2064 (N_2064,N_1948,N_1898);
or U2065 (N_2065,N_1941,N_1992);
xnor U2066 (N_2066,N_1963,N_1998);
nand U2067 (N_2067,N_1956,N_1936);
or U2068 (N_2068,N_1933,N_1913);
and U2069 (N_2069,N_1994,N_1947);
nand U2070 (N_2070,N_1966,N_1911);
nand U2071 (N_2071,N_1941,N_1923);
and U2072 (N_2072,N_1977,N_1991);
xor U2073 (N_2073,N_1988,N_1886);
nand U2074 (N_2074,N_1879,N_1938);
and U2075 (N_2075,N_1921,N_1950);
nor U2076 (N_2076,N_1949,N_1978);
nor U2077 (N_2077,N_1950,N_1912);
xor U2078 (N_2078,N_1946,N_1966);
or U2079 (N_2079,N_1990,N_1936);
xnor U2080 (N_2080,N_1969,N_1898);
nor U2081 (N_2081,N_1906,N_1994);
xor U2082 (N_2082,N_1966,N_1888);
xor U2083 (N_2083,N_1997,N_1893);
nand U2084 (N_2084,N_1884,N_1891);
nor U2085 (N_2085,N_1922,N_1952);
and U2086 (N_2086,N_1981,N_1881);
and U2087 (N_2087,N_1937,N_1965);
and U2088 (N_2088,N_1991,N_1988);
nand U2089 (N_2089,N_1889,N_1926);
xor U2090 (N_2090,N_1896,N_1941);
and U2091 (N_2091,N_1995,N_1934);
or U2092 (N_2092,N_1974,N_1998);
nor U2093 (N_2093,N_1905,N_1915);
nor U2094 (N_2094,N_1921,N_1948);
and U2095 (N_2095,N_1915,N_1973);
xnor U2096 (N_2096,N_1932,N_1904);
nor U2097 (N_2097,N_1951,N_1969);
nand U2098 (N_2098,N_1886,N_1970);
or U2099 (N_2099,N_1977,N_1952);
xnor U2100 (N_2100,N_1998,N_1911);
and U2101 (N_2101,N_1995,N_1976);
nor U2102 (N_2102,N_1966,N_1875);
nor U2103 (N_2103,N_1882,N_1928);
and U2104 (N_2104,N_1927,N_1879);
and U2105 (N_2105,N_1965,N_1928);
or U2106 (N_2106,N_1935,N_1960);
nand U2107 (N_2107,N_1880,N_1935);
xor U2108 (N_2108,N_1984,N_1946);
and U2109 (N_2109,N_1892,N_1963);
or U2110 (N_2110,N_1989,N_1952);
nor U2111 (N_2111,N_1878,N_1947);
nor U2112 (N_2112,N_1921,N_1885);
and U2113 (N_2113,N_1944,N_1977);
xnor U2114 (N_2114,N_1904,N_1893);
xor U2115 (N_2115,N_1939,N_1943);
or U2116 (N_2116,N_1913,N_1924);
nand U2117 (N_2117,N_1925,N_1889);
nand U2118 (N_2118,N_1958,N_1983);
nand U2119 (N_2119,N_1988,N_1902);
nand U2120 (N_2120,N_1951,N_1882);
nand U2121 (N_2121,N_1977,N_1894);
and U2122 (N_2122,N_1876,N_1911);
nor U2123 (N_2123,N_1907,N_1972);
xor U2124 (N_2124,N_1988,N_1926);
and U2125 (N_2125,N_2077,N_2031);
nor U2126 (N_2126,N_2023,N_2052);
nor U2127 (N_2127,N_2054,N_2019);
nor U2128 (N_2128,N_2119,N_2041);
xnor U2129 (N_2129,N_2046,N_2027);
or U2130 (N_2130,N_2092,N_2030);
and U2131 (N_2131,N_2124,N_2107);
nor U2132 (N_2132,N_2014,N_2074);
xnor U2133 (N_2133,N_2058,N_2106);
nand U2134 (N_2134,N_2096,N_2038);
xnor U2135 (N_2135,N_2075,N_2013);
and U2136 (N_2136,N_2001,N_2010);
nor U2137 (N_2137,N_2007,N_2000);
nor U2138 (N_2138,N_2085,N_2061);
and U2139 (N_2139,N_2120,N_2012);
xnor U2140 (N_2140,N_2083,N_2048);
xor U2141 (N_2141,N_2004,N_2086);
nor U2142 (N_2142,N_2091,N_2084);
nand U2143 (N_2143,N_2088,N_2029);
and U2144 (N_2144,N_2051,N_2110);
and U2145 (N_2145,N_2042,N_2036);
nand U2146 (N_2146,N_2065,N_2006);
or U2147 (N_2147,N_2028,N_2109);
nor U2148 (N_2148,N_2011,N_2069);
nand U2149 (N_2149,N_2062,N_2111);
nor U2150 (N_2150,N_2089,N_2080);
nand U2151 (N_2151,N_2094,N_2108);
or U2152 (N_2152,N_2047,N_2097);
and U2153 (N_2153,N_2008,N_2101);
and U2154 (N_2154,N_2076,N_2103);
xor U2155 (N_2155,N_2068,N_2043);
and U2156 (N_2156,N_2040,N_2113);
and U2157 (N_2157,N_2104,N_2116);
xnor U2158 (N_2158,N_2037,N_2059);
and U2159 (N_2159,N_2064,N_2050);
or U2160 (N_2160,N_2115,N_2117);
xor U2161 (N_2161,N_2002,N_2102);
nor U2162 (N_2162,N_2122,N_2121);
nor U2163 (N_2163,N_2016,N_2005);
nand U2164 (N_2164,N_2044,N_2093);
xor U2165 (N_2165,N_2033,N_2045);
xor U2166 (N_2166,N_2017,N_2123);
or U2167 (N_2167,N_2060,N_2025);
nor U2168 (N_2168,N_2100,N_2020);
nand U2169 (N_2169,N_2118,N_2053);
nor U2170 (N_2170,N_2056,N_2039);
nand U2171 (N_2171,N_2034,N_2018);
nor U2172 (N_2172,N_2112,N_2035);
or U2173 (N_2173,N_2087,N_2049);
nor U2174 (N_2174,N_2024,N_2095);
or U2175 (N_2175,N_2082,N_2026);
or U2176 (N_2176,N_2078,N_2055);
or U2177 (N_2177,N_2021,N_2032);
xnor U2178 (N_2178,N_2079,N_2066);
nand U2179 (N_2179,N_2114,N_2071);
xnor U2180 (N_2180,N_2105,N_2003);
and U2181 (N_2181,N_2015,N_2063);
nand U2182 (N_2182,N_2098,N_2070);
and U2183 (N_2183,N_2009,N_2081);
and U2184 (N_2184,N_2022,N_2090);
and U2185 (N_2185,N_2067,N_2099);
or U2186 (N_2186,N_2057,N_2073);
nand U2187 (N_2187,N_2072,N_2026);
nand U2188 (N_2188,N_2042,N_2056);
nand U2189 (N_2189,N_2029,N_2078);
nor U2190 (N_2190,N_2063,N_2038);
nor U2191 (N_2191,N_2049,N_2070);
xor U2192 (N_2192,N_2107,N_2063);
or U2193 (N_2193,N_2074,N_2040);
xnor U2194 (N_2194,N_2096,N_2100);
nand U2195 (N_2195,N_2114,N_2120);
nand U2196 (N_2196,N_2036,N_2083);
nor U2197 (N_2197,N_2107,N_2038);
nand U2198 (N_2198,N_2114,N_2044);
xor U2199 (N_2199,N_2039,N_2055);
nand U2200 (N_2200,N_2029,N_2077);
nor U2201 (N_2201,N_2073,N_2032);
and U2202 (N_2202,N_2118,N_2055);
or U2203 (N_2203,N_2036,N_2068);
nor U2204 (N_2204,N_2032,N_2020);
and U2205 (N_2205,N_2102,N_2061);
or U2206 (N_2206,N_2080,N_2009);
nand U2207 (N_2207,N_2005,N_2119);
and U2208 (N_2208,N_2103,N_2108);
nor U2209 (N_2209,N_2008,N_2034);
xnor U2210 (N_2210,N_2110,N_2018);
or U2211 (N_2211,N_2044,N_2086);
or U2212 (N_2212,N_2088,N_2022);
and U2213 (N_2213,N_2105,N_2070);
nor U2214 (N_2214,N_2025,N_2086);
xor U2215 (N_2215,N_2109,N_2021);
nand U2216 (N_2216,N_2078,N_2000);
or U2217 (N_2217,N_2065,N_2042);
or U2218 (N_2218,N_2046,N_2088);
xor U2219 (N_2219,N_2076,N_2054);
nand U2220 (N_2220,N_2011,N_2043);
nand U2221 (N_2221,N_2060,N_2014);
nand U2222 (N_2222,N_2072,N_2018);
or U2223 (N_2223,N_2101,N_2085);
xor U2224 (N_2224,N_2087,N_2089);
nor U2225 (N_2225,N_2025,N_2047);
and U2226 (N_2226,N_2014,N_2077);
or U2227 (N_2227,N_2010,N_2061);
nand U2228 (N_2228,N_2016,N_2050);
and U2229 (N_2229,N_2096,N_2103);
nand U2230 (N_2230,N_2062,N_2033);
xor U2231 (N_2231,N_2100,N_2005);
xor U2232 (N_2232,N_2010,N_2101);
or U2233 (N_2233,N_2115,N_2025);
nor U2234 (N_2234,N_2004,N_2040);
or U2235 (N_2235,N_2034,N_2040);
or U2236 (N_2236,N_2000,N_2079);
xor U2237 (N_2237,N_2090,N_2063);
and U2238 (N_2238,N_2110,N_2032);
nor U2239 (N_2239,N_2017,N_2090);
xor U2240 (N_2240,N_2059,N_2013);
nor U2241 (N_2241,N_2043,N_2026);
nor U2242 (N_2242,N_2094,N_2029);
xnor U2243 (N_2243,N_2032,N_2066);
xnor U2244 (N_2244,N_2054,N_2105);
and U2245 (N_2245,N_2060,N_2075);
or U2246 (N_2246,N_2046,N_2095);
or U2247 (N_2247,N_2011,N_2034);
or U2248 (N_2248,N_2080,N_2008);
or U2249 (N_2249,N_2051,N_2067);
or U2250 (N_2250,N_2168,N_2156);
xnor U2251 (N_2251,N_2153,N_2131);
and U2252 (N_2252,N_2246,N_2155);
xor U2253 (N_2253,N_2195,N_2169);
nor U2254 (N_2254,N_2132,N_2180);
or U2255 (N_2255,N_2224,N_2201);
and U2256 (N_2256,N_2174,N_2235);
nand U2257 (N_2257,N_2144,N_2159);
nand U2258 (N_2258,N_2248,N_2221);
nor U2259 (N_2259,N_2223,N_2236);
xor U2260 (N_2260,N_2189,N_2196);
xnor U2261 (N_2261,N_2145,N_2143);
xor U2262 (N_2262,N_2154,N_2187);
xor U2263 (N_2263,N_2173,N_2214);
nor U2264 (N_2264,N_2230,N_2225);
nand U2265 (N_2265,N_2140,N_2164);
and U2266 (N_2266,N_2162,N_2146);
xor U2267 (N_2267,N_2185,N_2207);
and U2268 (N_2268,N_2138,N_2237);
xor U2269 (N_2269,N_2147,N_2217);
nand U2270 (N_2270,N_2166,N_2244);
or U2271 (N_2271,N_2175,N_2188);
or U2272 (N_2272,N_2249,N_2233);
nor U2273 (N_2273,N_2216,N_2234);
nand U2274 (N_2274,N_2184,N_2204);
nor U2275 (N_2275,N_2181,N_2206);
or U2276 (N_2276,N_2243,N_2192);
and U2277 (N_2277,N_2229,N_2199);
xnor U2278 (N_2278,N_2208,N_2213);
xnor U2279 (N_2279,N_2172,N_2127);
nand U2280 (N_2280,N_2218,N_2210);
xor U2281 (N_2281,N_2158,N_2232);
or U2282 (N_2282,N_2141,N_2163);
nand U2283 (N_2283,N_2129,N_2183);
or U2284 (N_2284,N_2179,N_2212);
nand U2285 (N_2285,N_2203,N_2190);
xor U2286 (N_2286,N_2125,N_2130);
or U2287 (N_2287,N_2151,N_2227);
and U2288 (N_2288,N_2171,N_2167);
nand U2289 (N_2289,N_2231,N_2202);
xnor U2290 (N_2290,N_2197,N_2142);
nor U2291 (N_2291,N_2239,N_2128);
nand U2292 (N_2292,N_2170,N_2219);
xor U2293 (N_2293,N_2228,N_2161);
nor U2294 (N_2294,N_2177,N_2226);
nand U2295 (N_2295,N_2133,N_2222);
nand U2296 (N_2296,N_2209,N_2150);
and U2297 (N_2297,N_2126,N_2157);
nand U2298 (N_2298,N_2198,N_2191);
or U2299 (N_2299,N_2139,N_2247);
xor U2300 (N_2300,N_2165,N_2215);
and U2301 (N_2301,N_2242,N_2211);
nor U2302 (N_2302,N_2148,N_2205);
and U2303 (N_2303,N_2240,N_2160);
nand U2304 (N_2304,N_2241,N_2194);
or U2305 (N_2305,N_2152,N_2135);
nor U2306 (N_2306,N_2193,N_2134);
nor U2307 (N_2307,N_2238,N_2245);
nor U2308 (N_2308,N_2182,N_2149);
xnor U2309 (N_2309,N_2186,N_2220);
and U2310 (N_2310,N_2178,N_2137);
xnor U2311 (N_2311,N_2136,N_2200);
nor U2312 (N_2312,N_2176,N_2164);
xor U2313 (N_2313,N_2157,N_2231);
or U2314 (N_2314,N_2155,N_2135);
xnor U2315 (N_2315,N_2198,N_2242);
xnor U2316 (N_2316,N_2142,N_2151);
nor U2317 (N_2317,N_2188,N_2183);
and U2318 (N_2318,N_2168,N_2249);
nand U2319 (N_2319,N_2129,N_2166);
xor U2320 (N_2320,N_2151,N_2153);
or U2321 (N_2321,N_2231,N_2129);
nor U2322 (N_2322,N_2220,N_2176);
xnor U2323 (N_2323,N_2140,N_2183);
xor U2324 (N_2324,N_2191,N_2183);
or U2325 (N_2325,N_2164,N_2154);
and U2326 (N_2326,N_2133,N_2130);
nand U2327 (N_2327,N_2186,N_2245);
and U2328 (N_2328,N_2135,N_2149);
xnor U2329 (N_2329,N_2244,N_2235);
or U2330 (N_2330,N_2127,N_2131);
or U2331 (N_2331,N_2139,N_2149);
xnor U2332 (N_2332,N_2135,N_2224);
and U2333 (N_2333,N_2209,N_2226);
nor U2334 (N_2334,N_2175,N_2164);
nand U2335 (N_2335,N_2168,N_2188);
xnor U2336 (N_2336,N_2156,N_2174);
nand U2337 (N_2337,N_2203,N_2154);
nor U2338 (N_2338,N_2242,N_2233);
or U2339 (N_2339,N_2249,N_2193);
or U2340 (N_2340,N_2227,N_2247);
nor U2341 (N_2341,N_2247,N_2199);
or U2342 (N_2342,N_2190,N_2217);
nor U2343 (N_2343,N_2174,N_2227);
nor U2344 (N_2344,N_2178,N_2218);
or U2345 (N_2345,N_2221,N_2151);
or U2346 (N_2346,N_2159,N_2232);
nor U2347 (N_2347,N_2140,N_2198);
and U2348 (N_2348,N_2218,N_2235);
nor U2349 (N_2349,N_2210,N_2232);
nand U2350 (N_2350,N_2196,N_2219);
nor U2351 (N_2351,N_2164,N_2139);
nand U2352 (N_2352,N_2151,N_2182);
xor U2353 (N_2353,N_2142,N_2233);
nor U2354 (N_2354,N_2197,N_2207);
xor U2355 (N_2355,N_2205,N_2159);
xor U2356 (N_2356,N_2150,N_2157);
xnor U2357 (N_2357,N_2242,N_2208);
and U2358 (N_2358,N_2182,N_2196);
nor U2359 (N_2359,N_2234,N_2197);
and U2360 (N_2360,N_2215,N_2201);
or U2361 (N_2361,N_2147,N_2190);
xor U2362 (N_2362,N_2217,N_2247);
nor U2363 (N_2363,N_2222,N_2203);
nor U2364 (N_2364,N_2126,N_2147);
and U2365 (N_2365,N_2242,N_2160);
nor U2366 (N_2366,N_2206,N_2169);
and U2367 (N_2367,N_2125,N_2207);
xor U2368 (N_2368,N_2176,N_2244);
nand U2369 (N_2369,N_2227,N_2199);
nor U2370 (N_2370,N_2129,N_2215);
or U2371 (N_2371,N_2132,N_2135);
and U2372 (N_2372,N_2176,N_2230);
xor U2373 (N_2373,N_2232,N_2141);
nor U2374 (N_2374,N_2169,N_2148);
xor U2375 (N_2375,N_2290,N_2310);
xnor U2376 (N_2376,N_2272,N_2297);
or U2377 (N_2377,N_2295,N_2269);
nor U2378 (N_2378,N_2323,N_2274);
nand U2379 (N_2379,N_2264,N_2354);
and U2380 (N_2380,N_2278,N_2282);
nand U2381 (N_2381,N_2324,N_2267);
or U2382 (N_2382,N_2280,N_2369);
and U2383 (N_2383,N_2338,N_2342);
nand U2384 (N_2384,N_2302,N_2270);
nor U2385 (N_2385,N_2330,N_2262);
nor U2386 (N_2386,N_2259,N_2303);
nor U2387 (N_2387,N_2289,N_2299);
or U2388 (N_2388,N_2350,N_2370);
and U2389 (N_2389,N_2333,N_2281);
nand U2390 (N_2390,N_2339,N_2288);
xor U2391 (N_2391,N_2358,N_2265);
xor U2392 (N_2392,N_2285,N_2291);
nand U2393 (N_2393,N_2361,N_2276);
nand U2394 (N_2394,N_2373,N_2301);
nand U2395 (N_2395,N_2341,N_2328);
and U2396 (N_2396,N_2293,N_2315);
and U2397 (N_2397,N_2296,N_2352);
nand U2398 (N_2398,N_2366,N_2307);
or U2399 (N_2399,N_2363,N_2322);
nor U2400 (N_2400,N_2359,N_2349);
xnor U2401 (N_2401,N_2263,N_2348);
nand U2402 (N_2402,N_2308,N_2316);
or U2403 (N_2403,N_2253,N_2258);
nand U2404 (N_2404,N_2372,N_2319);
xor U2405 (N_2405,N_2325,N_2306);
nand U2406 (N_2406,N_2317,N_2331);
nand U2407 (N_2407,N_2374,N_2273);
nor U2408 (N_2408,N_2309,N_2298);
and U2409 (N_2409,N_2329,N_2250);
nand U2410 (N_2410,N_2277,N_2335);
nor U2411 (N_2411,N_2304,N_2286);
and U2412 (N_2412,N_2300,N_2346);
nand U2413 (N_2413,N_2364,N_2334);
nor U2414 (N_2414,N_2368,N_2343);
xor U2415 (N_2415,N_2260,N_2326);
and U2416 (N_2416,N_2327,N_2271);
xor U2417 (N_2417,N_2283,N_2284);
nor U2418 (N_2418,N_2257,N_2371);
and U2419 (N_2419,N_2365,N_2312);
or U2420 (N_2420,N_2292,N_2254);
or U2421 (N_2421,N_2275,N_2356);
nor U2422 (N_2422,N_2340,N_2351);
nand U2423 (N_2423,N_2305,N_2287);
and U2424 (N_2424,N_2347,N_2320);
or U2425 (N_2425,N_2294,N_2332);
or U2426 (N_2426,N_2337,N_2266);
and U2427 (N_2427,N_2318,N_2336);
and U2428 (N_2428,N_2279,N_2362);
nand U2429 (N_2429,N_2353,N_2314);
nor U2430 (N_2430,N_2321,N_2345);
nand U2431 (N_2431,N_2367,N_2252);
nor U2432 (N_2432,N_2360,N_2261);
xnor U2433 (N_2433,N_2357,N_2344);
nand U2434 (N_2434,N_2268,N_2313);
xnor U2435 (N_2435,N_2256,N_2251);
xor U2436 (N_2436,N_2355,N_2255);
nand U2437 (N_2437,N_2311,N_2284);
xnor U2438 (N_2438,N_2257,N_2311);
and U2439 (N_2439,N_2372,N_2320);
and U2440 (N_2440,N_2327,N_2372);
nor U2441 (N_2441,N_2250,N_2335);
or U2442 (N_2442,N_2303,N_2340);
xor U2443 (N_2443,N_2365,N_2301);
and U2444 (N_2444,N_2335,N_2340);
xor U2445 (N_2445,N_2281,N_2309);
and U2446 (N_2446,N_2279,N_2303);
and U2447 (N_2447,N_2344,N_2349);
or U2448 (N_2448,N_2361,N_2319);
nand U2449 (N_2449,N_2342,N_2357);
and U2450 (N_2450,N_2372,N_2365);
and U2451 (N_2451,N_2278,N_2335);
or U2452 (N_2452,N_2256,N_2295);
nor U2453 (N_2453,N_2313,N_2357);
or U2454 (N_2454,N_2268,N_2281);
or U2455 (N_2455,N_2254,N_2372);
and U2456 (N_2456,N_2360,N_2319);
or U2457 (N_2457,N_2351,N_2267);
xor U2458 (N_2458,N_2302,N_2349);
nor U2459 (N_2459,N_2294,N_2312);
nand U2460 (N_2460,N_2293,N_2288);
or U2461 (N_2461,N_2347,N_2278);
nor U2462 (N_2462,N_2310,N_2279);
xnor U2463 (N_2463,N_2271,N_2269);
and U2464 (N_2464,N_2339,N_2369);
or U2465 (N_2465,N_2332,N_2315);
xor U2466 (N_2466,N_2267,N_2301);
and U2467 (N_2467,N_2306,N_2370);
nand U2468 (N_2468,N_2364,N_2264);
nor U2469 (N_2469,N_2290,N_2346);
and U2470 (N_2470,N_2328,N_2356);
and U2471 (N_2471,N_2356,N_2294);
nor U2472 (N_2472,N_2258,N_2339);
nor U2473 (N_2473,N_2356,N_2282);
and U2474 (N_2474,N_2252,N_2346);
xnor U2475 (N_2475,N_2259,N_2336);
and U2476 (N_2476,N_2266,N_2279);
nor U2477 (N_2477,N_2291,N_2286);
nor U2478 (N_2478,N_2313,N_2327);
or U2479 (N_2479,N_2301,N_2259);
nand U2480 (N_2480,N_2340,N_2353);
nor U2481 (N_2481,N_2328,N_2303);
nor U2482 (N_2482,N_2349,N_2271);
and U2483 (N_2483,N_2270,N_2269);
nand U2484 (N_2484,N_2262,N_2337);
or U2485 (N_2485,N_2338,N_2331);
xor U2486 (N_2486,N_2311,N_2365);
or U2487 (N_2487,N_2318,N_2372);
and U2488 (N_2488,N_2318,N_2357);
or U2489 (N_2489,N_2279,N_2366);
and U2490 (N_2490,N_2308,N_2283);
nor U2491 (N_2491,N_2345,N_2266);
nor U2492 (N_2492,N_2352,N_2311);
nor U2493 (N_2493,N_2305,N_2280);
and U2494 (N_2494,N_2342,N_2284);
and U2495 (N_2495,N_2368,N_2354);
and U2496 (N_2496,N_2310,N_2355);
xnor U2497 (N_2497,N_2292,N_2366);
nand U2498 (N_2498,N_2361,N_2260);
or U2499 (N_2499,N_2362,N_2295);
nor U2500 (N_2500,N_2396,N_2399);
xor U2501 (N_2501,N_2468,N_2379);
and U2502 (N_2502,N_2435,N_2417);
xor U2503 (N_2503,N_2451,N_2452);
or U2504 (N_2504,N_2450,N_2428);
or U2505 (N_2505,N_2423,N_2392);
and U2506 (N_2506,N_2397,N_2407);
nor U2507 (N_2507,N_2386,N_2471);
xor U2508 (N_2508,N_2491,N_2383);
nor U2509 (N_2509,N_2472,N_2456);
and U2510 (N_2510,N_2464,N_2400);
nand U2511 (N_2511,N_2421,N_2461);
or U2512 (N_2512,N_2387,N_2427);
or U2513 (N_2513,N_2391,N_2488);
nor U2514 (N_2514,N_2445,N_2486);
or U2515 (N_2515,N_2459,N_2495);
xor U2516 (N_2516,N_2385,N_2381);
and U2517 (N_2517,N_2376,N_2416);
and U2518 (N_2518,N_2414,N_2411);
nor U2519 (N_2519,N_2393,N_2475);
nor U2520 (N_2520,N_2430,N_2498);
xor U2521 (N_2521,N_2409,N_2478);
nor U2522 (N_2522,N_2462,N_2412);
and U2523 (N_2523,N_2403,N_2436);
xnor U2524 (N_2524,N_2454,N_2440);
xnor U2525 (N_2525,N_2453,N_2473);
or U2526 (N_2526,N_2493,N_2490);
or U2527 (N_2527,N_2434,N_2398);
or U2528 (N_2528,N_2460,N_2426);
nand U2529 (N_2529,N_2415,N_2429);
or U2530 (N_2530,N_2446,N_2389);
xnor U2531 (N_2531,N_2494,N_2476);
or U2532 (N_2532,N_2384,N_2404);
and U2533 (N_2533,N_2420,N_2441);
xnor U2534 (N_2534,N_2402,N_2449);
nor U2535 (N_2535,N_2419,N_2482);
xnor U2536 (N_2536,N_2443,N_2485);
and U2537 (N_2537,N_2487,N_2425);
or U2538 (N_2538,N_2448,N_2442);
nor U2539 (N_2539,N_2438,N_2496);
or U2540 (N_2540,N_2479,N_2394);
nand U2541 (N_2541,N_2432,N_2377);
or U2542 (N_2542,N_2424,N_2431);
xnor U2543 (N_2543,N_2390,N_2492);
xor U2544 (N_2544,N_2463,N_2474);
nand U2545 (N_2545,N_2418,N_2481);
nand U2546 (N_2546,N_2480,N_2401);
or U2547 (N_2547,N_2469,N_2380);
or U2548 (N_2548,N_2465,N_2477);
or U2549 (N_2549,N_2395,N_2437);
nand U2550 (N_2550,N_2408,N_2467);
nor U2551 (N_2551,N_2405,N_2489);
and U2552 (N_2552,N_2497,N_2413);
xnor U2553 (N_2553,N_2406,N_2433);
nand U2554 (N_2554,N_2484,N_2422);
or U2555 (N_2555,N_2444,N_2466);
and U2556 (N_2556,N_2410,N_2457);
nand U2557 (N_2557,N_2382,N_2447);
nand U2558 (N_2558,N_2439,N_2378);
or U2559 (N_2559,N_2470,N_2458);
nor U2560 (N_2560,N_2455,N_2483);
xnor U2561 (N_2561,N_2375,N_2499);
or U2562 (N_2562,N_2388,N_2406);
nor U2563 (N_2563,N_2379,N_2488);
or U2564 (N_2564,N_2471,N_2379);
and U2565 (N_2565,N_2449,N_2461);
xnor U2566 (N_2566,N_2462,N_2399);
nor U2567 (N_2567,N_2442,N_2496);
nor U2568 (N_2568,N_2435,N_2402);
nor U2569 (N_2569,N_2394,N_2384);
nand U2570 (N_2570,N_2457,N_2445);
nor U2571 (N_2571,N_2425,N_2377);
nor U2572 (N_2572,N_2418,N_2413);
nand U2573 (N_2573,N_2469,N_2423);
nor U2574 (N_2574,N_2393,N_2414);
nor U2575 (N_2575,N_2418,N_2444);
nand U2576 (N_2576,N_2404,N_2420);
xnor U2577 (N_2577,N_2398,N_2484);
xnor U2578 (N_2578,N_2485,N_2448);
nor U2579 (N_2579,N_2471,N_2468);
nor U2580 (N_2580,N_2492,N_2455);
nor U2581 (N_2581,N_2414,N_2446);
nand U2582 (N_2582,N_2453,N_2451);
nor U2583 (N_2583,N_2440,N_2413);
or U2584 (N_2584,N_2420,N_2468);
nand U2585 (N_2585,N_2411,N_2479);
nor U2586 (N_2586,N_2469,N_2399);
nor U2587 (N_2587,N_2485,N_2396);
xnor U2588 (N_2588,N_2428,N_2451);
and U2589 (N_2589,N_2392,N_2388);
and U2590 (N_2590,N_2406,N_2413);
xnor U2591 (N_2591,N_2481,N_2473);
nand U2592 (N_2592,N_2462,N_2485);
xor U2593 (N_2593,N_2389,N_2484);
or U2594 (N_2594,N_2470,N_2385);
or U2595 (N_2595,N_2407,N_2423);
nor U2596 (N_2596,N_2414,N_2441);
and U2597 (N_2597,N_2457,N_2498);
xnor U2598 (N_2598,N_2390,N_2473);
nor U2599 (N_2599,N_2487,N_2401);
nor U2600 (N_2600,N_2397,N_2409);
nor U2601 (N_2601,N_2411,N_2388);
xor U2602 (N_2602,N_2402,N_2376);
xnor U2603 (N_2603,N_2430,N_2447);
and U2604 (N_2604,N_2496,N_2420);
and U2605 (N_2605,N_2490,N_2464);
nand U2606 (N_2606,N_2497,N_2411);
and U2607 (N_2607,N_2411,N_2424);
nor U2608 (N_2608,N_2472,N_2414);
and U2609 (N_2609,N_2464,N_2475);
xor U2610 (N_2610,N_2458,N_2403);
nor U2611 (N_2611,N_2480,N_2470);
xor U2612 (N_2612,N_2375,N_2482);
or U2613 (N_2613,N_2499,N_2438);
xnor U2614 (N_2614,N_2479,N_2414);
nor U2615 (N_2615,N_2497,N_2426);
nor U2616 (N_2616,N_2469,N_2466);
or U2617 (N_2617,N_2375,N_2421);
or U2618 (N_2618,N_2450,N_2404);
and U2619 (N_2619,N_2482,N_2399);
or U2620 (N_2620,N_2452,N_2475);
nand U2621 (N_2621,N_2460,N_2443);
or U2622 (N_2622,N_2426,N_2388);
or U2623 (N_2623,N_2498,N_2471);
nand U2624 (N_2624,N_2383,N_2391);
or U2625 (N_2625,N_2583,N_2507);
nand U2626 (N_2626,N_2553,N_2557);
nand U2627 (N_2627,N_2615,N_2574);
and U2628 (N_2628,N_2504,N_2616);
xnor U2629 (N_2629,N_2579,N_2575);
or U2630 (N_2630,N_2587,N_2503);
or U2631 (N_2631,N_2617,N_2555);
nor U2632 (N_2632,N_2520,N_2543);
and U2633 (N_2633,N_2565,N_2576);
xnor U2634 (N_2634,N_2578,N_2526);
xnor U2635 (N_2635,N_2558,N_2609);
nand U2636 (N_2636,N_2593,N_2586);
nand U2637 (N_2637,N_2540,N_2514);
and U2638 (N_2638,N_2562,N_2500);
nand U2639 (N_2639,N_2550,N_2538);
and U2640 (N_2640,N_2539,N_2554);
xor U2641 (N_2641,N_2595,N_2512);
and U2642 (N_2642,N_2612,N_2572);
xor U2643 (N_2643,N_2551,N_2598);
or U2644 (N_2644,N_2618,N_2610);
nor U2645 (N_2645,N_2525,N_2620);
nand U2646 (N_2646,N_2501,N_2622);
nor U2647 (N_2647,N_2608,N_2519);
or U2648 (N_2648,N_2624,N_2528);
or U2649 (N_2649,N_2511,N_2573);
or U2650 (N_2650,N_2599,N_2596);
or U2651 (N_2651,N_2566,N_2602);
nor U2652 (N_2652,N_2548,N_2580);
or U2653 (N_2653,N_2571,N_2581);
nand U2654 (N_2654,N_2535,N_2614);
nor U2655 (N_2655,N_2600,N_2522);
xor U2656 (N_2656,N_2556,N_2567);
xnor U2657 (N_2657,N_2563,N_2516);
nor U2658 (N_2658,N_2537,N_2523);
nor U2659 (N_2659,N_2564,N_2584);
and U2660 (N_2660,N_2585,N_2592);
nor U2661 (N_2661,N_2588,N_2517);
xor U2662 (N_2662,N_2619,N_2510);
and U2663 (N_2663,N_2594,N_2623);
nand U2664 (N_2664,N_2569,N_2534);
or U2665 (N_2665,N_2590,N_2549);
nand U2666 (N_2666,N_2505,N_2552);
xnor U2667 (N_2667,N_2527,N_2582);
xor U2668 (N_2668,N_2597,N_2547);
or U2669 (N_2669,N_2502,N_2544);
and U2670 (N_2670,N_2542,N_2604);
nor U2671 (N_2671,N_2531,N_2508);
nand U2672 (N_2672,N_2515,N_2513);
xor U2673 (N_2673,N_2560,N_2545);
nor U2674 (N_2674,N_2568,N_2601);
and U2675 (N_2675,N_2561,N_2613);
xnor U2676 (N_2676,N_2506,N_2524);
xnor U2677 (N_2677,N_2606,N_2591);
nor U2678 (N_2678,N_2570,N_2532);
or U2679 (N_2679,N_2605,N_2530);
nand U2680 (N_2680,N_2541,N_2546);
nand U2681 (N_2681,N_2559,N_2533);
nor U2682 (N_2682,N_2509,N_2603);
and U2683 (N_2683,N_2607,N_2621);
nor U2684 (N_2684,N_2589,N_2536);
or U2685 (N_2685,N_2518,N_2521);
xnor U2686 (N_2686,N_2577,N_2529);
and U2687 (N_2687,N_2611,N_2587);
nor U2688 (N_2688,N_2506,N_2503);
nand U2689 (N_2689,N_2549,N_2532);
and U2690 (N_2690,N_2583,N_2521);
or U2691 (N_2691,N_2504,N_2557);
and U2692 (N_2692,N_2543,N_2500);
xor U2693 (N_2693,N_2500,N_2622);
xnor U2694 (N_2694,N_2549,N_2601);
or U2695 (N_2695,N_2563,N_2526);
xor U2696 (N_2696,N_2604,N_2500);
nand U2697 (N_2697,N_2530,N_2618);
or U2698 (N_2698,N_2548,N_2568);
or U2699 (N_2699,N_2550,N_2588);
nor U2700 (N_2700,N_2582,N_2548);
nand U2701 (N_2701,N_2522,N_2531);
or U2702 (N_2702,N_2507,N_2519);
xor U2703 (N_2703,N_2569,N_2550);
or U2704 (N_2704,N_2591,N_2573);
xor U2705 (N_2705,N_2595,N_2503);
nor U2706 (N_2706,N_2612,N_2552);
nor U2707 (N_2707,N_2521,N_2606);
or U2708 (N_2708,N_2551,N_2557);
or U2709 (N_2709,N_2564,N_2506);
nand U2710 (N_2710,N_2569,N_2577);
xnor U2711 (N_2711,N_2608,N_2547);
nor U2712 (N_2712,N_2542,N_2501);
nand U2713 (N_2713,N_2565,N_2591);
or U2714 (N_2714,N_2546,N_2516);
or U2715 (N_2715,N_2594,N_2550);
and U2716 (N_2716,N_2572,N_2611);
nor U2717 (N_2717,N_2559,N_2505);
xor U2718 (N_2718,N_2590,N_2613);
and U2719 (N_2719,N_2587,N_2618);
nor U2720 (N_2720,N_2521,N_2603);
xor U2721 (N_2721,N_2545,N_2605);
or U2722 (N_2722,N_2554,N_2519);
and U2723 (N_2723,N_2620,N_2541);
and U2724 (N_2724,N_2563,N_2591);
nor U2725 (N_2725,N_2530,N_2529);
xnor U2726 (N_2726,N_2535,N_2606);
nor U2727 (N_2727,N_2529,N_2510);
and U2728 (N_2728,N_2521,N_2595);
nor U2729 (N_2729,N_2505,N_2602);
nor U2730 (N_2730,N_2616,N_2605);
or U2731 (N_2731,N_2607,N_2543);
nor U2732 (N_2732,N_2614,N_2579);
and U2733 (N_2733,N_2570,N_2600);
nand U2734 (N_2734,N_2517,N_2502);
nor U2735 (N_2735,N_2508,N_2623);
and U2736 (N_2736,N_2547,N_2532);
or U2737 (N_2737,N_2582,N_2557);
xnor U2738 (N_2738,N_2523,N_2567);
or U2739 (N_2739,N_2581,N_2505);
and U2740 (N_2740,N_2608,N_2620);
and U2741 (N_2741,N_2576,N_2507);
nor U2742 (N_2742,N_2543,N_2562);
nand U2743 (N_2743,N_2517,N_2586);
and U2744 (N_2744,N_2566,N_2599);
xor U2745 (N_2745,N_2537,N_2585);
nor U2746 (N_2746,N_2520,N_2585);
nand U2747 (N_2747,N_2609,N_2547);
nand U2748 (N_2748,N_2534,N_2525);
nand U2749 (N_2749,N_2542,N_2504);
and U2750 (N_2750,N_2647,N_2707);
or U2751 (N_2751,N_2673,N_2712);
xor U2752 (N_2752,N_2636,N_2708);
nand U2753 (N_2753,N_2680,N_2739);
and U2754 (N_2754,N_2710,N_2679);
nand U2755 (N_2755,N_2703,N_2667);
or U2756 (N_2756,N_2684,N_2671);
xor U2757 (N_2757,N_2730,N_2657);
and U2758 (N_2758,N_2691,N_2714);
xnor U2759 (N_2759,N_2746,N_2699);
or U2760 (N_2760,N_2744,N_2737);
or U2761 (N_2761,N_2749,N_2745);
or U2762 (N_2762,N_2715,N_2687);
xor U2763 (N_2763,N_2627,N_2742);
nand U2764 (N_2764,N_2731,N_2669);
nand U2765 (N_2765,N_2666,N_2640);
and U2766 (N_2766,N_2692,N_2725);
nor U2767 (N_2767,N_2653,N_2706);
or U2768 (N_2768,N_2645,N_2656);
xnor U2769 (N_2769,N_2641,N_2676);
and U2770 (N_2770,N_2711,N_2690);
and U2771 (N_2771,N_2695,N_2697);
and U2772 (N_2772,N_2632,N_2705);
nand U2773 (N_2773,N_2748,N_2642);
nor U2774 (N_2774,N_2674,N_2654);
nor U2775 (N_2775,N_2722,N_2721);
nand U2776 (N_2776,N_2625,N_2670);
nand U2777 (N_2777,N_2688,N_2660);
and U2778 (N_2778,N_2644,N_2663);
or U2779 (N_2779,N_2727,N_2686);
nand U2780 (N_2780,N_2668,N_2633);
xor U2781 (N_2781,N_2701,N_2689);
xor U2782 (N_2782,N_2735,N_2719);
and U2783 (N_2783,N_2700,N_2681);
xor U2784 (N_2784,N_2677,N_2733);
nand U2785 (N_2785,N_2631,N_2635);
or U2786 (N_2786,N_2726,N_2639);
and U2787 (N_2787,N_2659,N_2728);
and U2788 (N_2788,N_2718,N_2723);
xnor U2789 (N_2789,N_2729,N_2655);
and U2790 (N_2790,N_2651,N_2661);
or U2791 (N_2791,N_2717,N_2720);
nor U2792 (N_2792,N_2683,N_2704);
nand U2793 (N_2793,N_2652,N_2743);
and U2794 (N_2794,N_2713,N_2648);
nor U2795 (N_2795,N_2740,N_2736);
and U2796 (N_2796,N_2685,N_2649);
nand U2797 (N_2797,N_2678,N_2650);
and U2798 (N_2798,N_2732,N_2747);
nor U2799 (N_2799,N_2626,N_2738);
nor U2800 (N_2800,N_2658,N_2630);
or U2801 (N_2801,N_2709,N_2682);
or U2802 (N_2802,N_2698,N_2646);
and U2803 (N_2803,N_2638,N_2643);
or U2804 (N_2804,N_2665,N_2716);
or U2805 (N_2805,N_2672,N_2662);
xor U2806 (N_2806,N_2741,N_2634);
and U2807 (N_2807,N_2664,N_2693);
nand U2808 (N_2808,N_2694,N_2734);
nand U2809 (N_2809,N_2724,N_2629);
and U2810 (N_2810,N_2702,N_2628);
or U2811 (N_2811,N_2637,N_2675);
nand U2812 (N_2812,N_2696,N_2687);
nand U2813 (N_2813,N_2656,N_2678);
nand U2814 (N_2814,N_2667,N_2653);
nand U2815 (N_2815,N_2656,N_2694);
nor U2816 (N_2816,N_2653,N_2675);
and U2817 (N_2817,N_2704,N_2710);
nor U2818 (N_2818,N_2738,N_2739);
xnor U2819 (N_2819,N_2653,N_2658);
and U2820 (N_2820,N_2744,N_2648);
or U2821 (N_2821,N_2627,N_2720);
xor U2822 (N_2822,N_2673,N_2721);
or U2823 (N_2823,N_2664,N_2657);
or U2824 (N_2824,N_2684,N_2628);
xor U2825 (N_2825,N_2666,N_2631);
nand U2826 (N_2826,N_2736,N_2693);
or U2827 (N_2827,N_2673,N_2665);
xnor U2828 (N_2828,N_2704,N_2722);
nand U2829 (N_2829,N_2680,N_2694);
or U2830 (N_2830,N_2647,N_2697);
nand U2831 (N_2831,N_2626,N_2702);
xor U2832 (N_2832,N_2658,N_2691);
or U2833 (N_2833,N_2737,N_2710);
nor U2834 (N_2834,N_2726,N_2748);
xor U2835 (N_2835,N_2648,N_2638);
xor U2836 (N_2836,N_2669,N_2712);
or U2837 (N_2837,N_2730,N_2725);
xnor U2838 (N_2838,N_2719,N_2653);
nand U2839 (N_2839,N_2698,N_2675);
nand U2840 (N_2840,N_2714,N_2710);
xor U2841 (N_2841,N_2713,N_2676);
nand U2842 (N_2842,N_2729,N_2625);
nor U2843 (N_2843,N_2699,N_2749);
nand U2844 (N_2844,N_2684,N_2709);
nor U2845 (N_2845,N_2688,N_2736);
or U2846 (N_2846,N_2631,N_2719);
nor U2847 (N_2847,N_2680,N_2693);
xor U2848 (N_2848,N_2651,N_2697);
xor U2849 (N_2849,N_2637,N_2710);
nor U2850 (N_2850,N_2702,N_2749);
xor U2851 (N_2851,N_2722,N_2681);
nor U2852 (N_2852,N_2719,N_2681);
and U2853 (N_2853,N_2735,N_2679);
and U2854 (N_2854,N_2658,N_2719);
nor U2855 (N_2855,N_2705,N_2665);
nor U2856 (N_2856,N_2731,N_2682);
xnor U2857 (N_2857,N_2701,N_2714);
and U2858 (N_2858,N_2625,N_2686);
nor U2859 (N_2859,N_2701,N_2705);
or U2860 (N_2860,N_2663,N_2638);
or U2861 (N_2861,N_2644,N_2726);
or U2862 (N_2862,N_2745,N_2704);
or U2863 (N_2863,N_2739,N_2713);
and U2864 (N_2864,N_2734,N_2661);
nor U2865 (N_2865,N_2700,N_2643);
nor U2866 (N_2866,N_2706,N_2725);
nand U2867 (N_2867,N_2732,N_2635);
xor U2868 (N_2868,N_2634,N_2635);
or U2869 (N_2869,N_2677,N_2718);
nor U2870 (N_2870,N_2635,N_2680);
or U2871 (N_2871,N_2648,N_2743);
xor U2872 (N_2872,N_2741,N_2694);
xnor U2873 (N_2873,N_2626,N_2639);
nand U2874 (N_2874,N_2748,N_2712);
and U2875 (N_2875,N_2846,N_2775);
xnor U2876 (N_2876,N_2791,N_2851);
or U2877 (N_2877,N_2816,N_2838);
xnor U2878 (N_2878,N_2815,N_2765);
and U2879 (N_2879,N_2849,N_2753);
nand U2880 (N_2880,N_2804,N_2793);
nor U2881 (N_2881,N_2780,N_2760);
nor U2882 (N_2882,N_2795,N_2784);
and U2883 (N_2883,N_2788,N_2763);
nand U2884 (N_2884,N_2840,N_2811);
nor U2885 (N_2885,N_2774,N_2865);
xnor U2886 (N_2886,N_2858,N_2808);
or U2887 (N_2887,N_2810,N_2752);
or U2888 (N_2888,N_2779,N_2862);
or U2889 (N_2889,N_2864,N_2839);
and U2890 (N_2890,N_2871,N_2819);
nand U2891 (N_2891,N_2859,N_2764);
nand U2892 (N_2892,N_2790,N_2826);
nor U2893 (N_2893,N_2854,N_2837);
nand U2894 (N_2894,N_2844,N_2809);
nor U2895 (N_2895,N_2757,N_2831);
xor U2896 (N_2896,N_2860,N_2853);
or U2897 (N_2897,N_2761,N_2800);
or U2898 (N_2898,N_2807,N_2767);
nand U2899 (N_2899,N_2855,N_2868);
nor U2900 (N_2900,N_2841,N_2817);
nor U2901 (N_2901,N_2798,N_2792);
nor U2902 (N_2902,N_2822,N_2867);
nor U2903 (N_2903,N_2812,N_2830);
xor U2904 (N_2904,N_2782,N_2869);
nand U2905 (N_2905,N_2751,N_2802);
nor U2906 (N_2906,N_2770,N_2772);
xor U2907 (N_2907,N_2756,N_2813);
nand U2908 (N_2908,N_2769,N_2785);
and U2909 (N_2909,N_2787,N_2856);
xor U2910 (N_2910,N_2776,N_2832);
nand U2911 (N_2911,N_2861,N_2872);
xnor U2912 (N_2912,N_2866,N_2870);
or U2913 (N_2913,N_2835,N_2824);
and U2914 (N_2914,N_2829,N_2762);
or U2915 (N_2915,N_2773,N_2755);
nor U2916 (N_2916,N_2771,N_2873);
nand U2917 (N_2917,N_2750,N_2778);
or U2918 (N_2918,N_2768,N_2857);
and U2919 (N_2919,N_2825,N_2754);
xor U2920 (N_2920,N_2801,N_2794);
and U2921 (N_2921,N_2847,N_2850);
or U2922 (N_2922,N_2852,N_2777);
and U2923 (N_2923,N_2827,N_2836);
xor U2924 (N_2924,N_2797,N_2766);
nand U2925 (N_2925,N_2783,N_2799);
and U2926 (N_2926,N_2759,N_2842);
and U2927 (N_2927,N_2818,N_2833);
and U2928 (N_2928,N_2786,N_2806);
xor U2929 (N_2929,N_2820,N_2874);
and U2930 (N_2930,N_2828,N_2758);
nand U2931 (N_2931,N_2796,N_2789);
or U2932 (N_2932,N_2781,N_2821);
and U2933 (N_2933,N_2848,N_2805);
nor U2934 (N_2934,N_2834,N_2843);
nor U2935 (N_2935,N_2823,N_2814);
and U2936 (N_2936,N_2803,N_2863);
or U2937 (N_2937,N_2845,N_2761);
and U2938 (N_2938,N_2814,N_2800);
xnor U2939 (N_2939,N_2788,N_2792);
or U2940 (N_2940,N_2774,N_2866);
nor U2941 (N_2941,N_2850,N_2843);
xor U2942 (N_2942,N_2827,N_2870);
or U2943 (N_2943,N_2827,N_2828);
or U2944 (N_2944,N_2750,N_2807);
or U2945 (N_2945,N_2828,N_2853);
xor U2946 (N_2946,N_2821,N_2797);
nand U2947 (N_2947,N_2831,N_2855);
nor U2948 (N_2948,N_2843,N_2790);
or U2949 (N_2949,N_2828,N_2851);
and U2950 (N_2950,N_2801,N_2815);
xnor U2951 (N_2951,N_2854,N_2824);
or U2952 (N_2952,N_2794,N_2829);
or U2953 (N_2953,N_2806,N_2782);
xor U2954 (N_2954,N_2859,N_2828);
and U2955 (N_2955,N_2760,N_2834);
xnor U2956 (N_2956,N_2754,N_2839);
nor U2957 (N_2957,N_2852,N_2871);
nor U2958 (N_2958,N_2814,N_2762);
nand U2959 (N_2959,N_2771,N_2758);
nor U2960 (N_2960,N_2832,N_2751);
nor U2961 (N_2961,N_2820,N_2786);
nor U2962 (N_2962,N_2840,N_2763);
xor U2963 (N_2963,N_2750,N_2794);
and U2964 (N_2964,N_2804,N_2780);
nor U2965 (N_2965,N_2803,N_2796);
or U2966 (N_2966,N_2853,N_2823);
nor U2967 (N_2967,N_2792,N_2847);
xnor U2968 (N_2968,N_2754,N_2774);
xnor U2969 (N_2969,N_2855,N_2838);
and U2970 (N_2970,N_2775,N_2758);
nor U2971 (N_2971,N_2797,N_2765);
xnor U2972 (N_2972,N_2845,N_2789);
and U2973 (N_2973,N_2859,N_2811);
nand U2974 (N_2974,N_2822,N_2827);
or U2975 (N_2975,N_2784,N_2850);
and U2976 (N_2976,N_2756,N_2873);
and U2977 (N_2977,N_2794,N_2847);
nor U2978 (N_2978,N_2757,N_2809);
nor U2979 (N_2979,N_2853,N_2838);
nand U2980 (N_2980,N_2790,N_2872);
xnor U2981 (N_2981,N_2781,N_2750);
and U2982 (N_2982,N_2774,N_2765);
nor U2983 (N_2983,N_2810,N_2869);
nand U2984 (N_2984,N_2804,N_2829);
and U2985 (N_2985,N_2753,N_2817);
or U2986 (N_2986,N_2774,N_2861);
nor U2987 (N_2987,N_2810,N_2759);
or U2988 (N_2988,N_2772,N_2844);
nand U2989 (N_2989,N_2776,N_2752);
and U2990 (N_2990,N_2826,N_2821);
nor U2991 (N_2991,N_2769,N_2845);
xor U2992 (N_2992,N_2800,N_2829);
and U2993 (N_2993,N_2765,N_2750);
and U2994 (N_2994,N_2853,N_2781);
nand U2995 (N_2995,N_2815,N_2764);
xor U2996 (N_2996,N_2761,N_2847);
nand U2997 (N_2997,N_2779,N_2772);
xnor U2998 (N_2998,N_2868,N_2835);
nand U2999 (N_2999,N_2842,N_2840);
nor U3000 (N_3000,N_2955,N_2929);
and U3001 (N_3001,N_2908,N_2966);
and U3002 (N_3002,N_2937,N_2896);
xnor U3003 (N_3003,N_2948,N_2935);
or U3004 (N_3004,N_2892,N_2918);
and U3005 (N_3005,N_2894,N_2979);
nor U3006 (N_3006,N_2989,N_2876);
or U3007 (N_3007,N_2893,N_2968);
nand U3008 (N_3008,N_2880,N_2921);
xnor U3009 (N_3009,N_2956,N_2925);
or U3010 (N_3010,N_2962,N_2971);
xnor U3011 (N_3011,N_2987,N_2899);
xnor U3012 (N_3012,N_2973,N_2957);
nand U3013 (N_3013,N_2952,N_2963);
nor U3014 (N_3014,N_2991,N_2949);
xnor U3015 (N_3015,N_2898,N_2917);
nand U3016 (N_3016,N_2912,N_2926);
and U3017 (N_3017,N_2878,N_2988);
nand U3018 (N_3018,N_2914,N_2886);
and U3019 (N_3019,N_2885,N_2950);
and U3020 (N_3020,N_2902,N_2923);
and U3021 (N_3021,N_2939,N_2986);
xor U3022 (N_3022,N_2932,N_2916);
or U3023 (N_3023,N_2901,N_2946);
nor U3024 (N_3024,N_2953,N_2961);
xnor U3025 (N_3025,N_2877,N_2959);
or U3026 (N_3026,N_2906,N_2910);
or U3027 (N_3027,N_2994,N_2982);
xnor U3028 (N_3028,N_2945,N_2990);
and U3029 (N_3029,N_2960,N_2911);
xor U3030 (N_3030,N_2889,N_2978);
nor U3031 (N_3031,N_2981,N_2922);
nand U3032 (N_3032,N_2931,N_2998);
xor U3033 (N_3033,N_2879,N_2930);
xnor U3034 (N_3034,N_2920,N_2881);
nand U3035 (N_3035,N_2924,N_2895);
and U3036 (N_3036,N_2938,N_2940);
nor U3037 (N_3037,N_2983,N_2958);
and U3038 (N_3038,N_2905,N_2954);
xnor U3039 (N_3039,N_2891,N_2997);
xnor U3040 (N_3040,N_2887,N_2969);
and U3041 (N_3041,N_2980,N_2951);
or U3042 (N_3042,N_2890,N_2999);
nand U3043 (N_3043,N_2919,N_2977);
nand U3044 (N_3044,N_2933,N_2884);
nor U3045 (N_3045,N_2903,N_2936);
xnor U3046 (N_3046,N_2996,N_2970);
or U3047 (N_3047,N_2942,N_2975);
nor U3048 (N_3048,N_2875,N_2915);
and U3049 (N_3049,N_2974,N_2888);
and U3050 (N_3050,N_2964,N_2992);
or U3051 (N_3051,N_2984,N_2909);
nor U3052 (N_3052,N_2965,N_2907);
xnor U3053 (N_3053,N_2967,N_2882);
xnor U3054 (N_3054,N_2993,N_2927);
nand U3055 (N_3055,N_2943,N_2947);
nand U3056 (N_3056,N_2976,N_2897);
nor U3057 (N_3057,N_2913,N_2900);
nor U3058 (N_3058,N_2941,N_2934);
xnor U3059 (N_3059,N_2928,N_2944);
nand U3060 (N_3060,N_2972,N_2985);
nor U3061 (N_3061,N_2904,N_2995);
xor U3062 (N_3062,N_2883,N_2903);
nor U3063 (N_3063,N_2895,N_2941);
or U3064 (N_3064,N_2903,N_2989);
and U3065 (N_3065,N_2947,N_2939);
xor U3066 (N_3066,N_2945,N_2934);
and U3067 (N_3067,N_2985,N_2957);
or U3068 (N_3068,N_2910,N_2896);
xnor U3069 (N_3069,N_2914,N_2882);
or U3070 (N_3070,N_2957,N_2980);
nand U3071 (N_3071,N_2910,N_2934);
nand U3072 (N_3072,N_2955,N_2878);
and U3073 (N_3073,N_2989,N_2928);
and U3074 (N_3074,N_2974,N_2911);
xnor U3075 (N_3075,N_2911,N_2954);
nor U3076 (N_3076,N_2980,N_2932);
and U3077 (N_3077,N_2886,N_2940);
nand U3078 (N_3078,N_2899,N_2954);
and U3079 (N_3079,N_2971,N_2904);
or U3080 (N_3080,N_2985,N_2999);
or U3081 (N_3081,N_2912,N_2883);
and U3082 (N_3082,N_2889,N_2916);
or U3083 (N_3083,N_2966,N_2951);
nor U3084 (N_3084,N_2965,N_2973);
and U3085 (N_3085,N_2958,N_2980);
or U3086 (N_3086,N_2876,N_2999);
nand U3087 (N_3087,N_2882,N_2947);
nor U3088 (N_3088,N_2908,N_2922);
and U3089 (N_3089,N_2968,N_2891);
xnor U3090 (N_3090,N_2983,N_2973);
nand U3091 (N_3091,N_2892,N_2929);
xor U3092 (N_3092,N_2875,N_2898);
and U3093 (N_3093,N_2895,N_2899);
and U3094 (N_3094,N_2890,N_2935);
or U3095 (N_3095,N_2923,N_2948);
and U3096 (N_3096,N_2920,N_2935);
nand U3097 (N_3097,N_2947,N_2942);
and U3098 (N_3098,N_2945,N_2950);
nor U3099 (N_3099,N_2896,N_2900);
nor U3100 (N_3100,N_2896,N_2959);
and U3101 (N_3101,N_2949,N_2875);
and U3102 (N_3102,N_2979,N_2876);
xnor U3103 (N_3103,N_2955,N_2924);
xor U3104 (N_3104,N_2897,N_2981);
or U3105 (N_3105,N_2926,N_2886);
nand U3106 (N_3106,N_2933,N_2934);
nor U3107 (N_3107,N_2960,N_2890);
nor U3108 (N_3108,N_2891,N_2972);
or U3109 (N_3109,N_2999,N_2893);
nand U3110 (N_3110,N_2878,N_2954);
nand U3111 (N_3111,N_2998,N_2944);
or U3112 (N_3112,N_2940,N_2914);
or U3113 (N_3113,N_2990,N_2956);
nand U3114 (N_3114,N_2882,N_2970);
xor U3115 (N_3115,N_2931,N_2951);
xor U3116 (N_3116,N_2993,N_2910);
and U3117 (N_3117,N_2912,N_2905);
or U3118 (N_3118,N_2965,N_2881);
nand U3119 (N_3119,N_2917,N_2932);
nand U3120 (N_3120,N_2980,N_2909);
nand U3121 (N_3121,N_2979,N_2999);
and U3122 (N_3122,N_2884,N_2958);
or U3123 (N_3123,N_2931,N_2976);
xnor U3124 (N_3124,N_2911,N_2900);
nor U3125 (N_3125,N_3056,N_3004);
nand U3126 (N_3126,N_3054,N_3052);
nand U3127 (N_3127,N_3062,N_3070);
or U3128 (N_3128,N_3082,N_3011);
nand U3129 (N_3129,N_3075,N_3058);
and U3130 (N_3130,N_3085,N_3023);
xor U3131 (N_3131,N_3022,N_3048);
nor U3132 (N_3132,N_3012,N_3064);
nor U3133 (N_3133,N_3107,N_3065);
nor U3134 (N_3134,N_3050,N_3018);
and U3135 (N_3135,N_3074,N_3110);
xor U3136 (N_3136,N_3120,N_3020);
nand U3137 (N_3137,N_3028,N_3097);
or U3138 (N_3138,N_3124,N_3057);
nor U3139 (N_3139,N_3067,N_3010);
nand U3140 (N_3140,N_3116,N_3027);
nand U3141 (N_3141,N_3014,N_3108);
or U3142 (N_3142,N_3095,N_3092);
nor U3143 (N_3143,N_3009,N_3040);
and U3144 (N_3144,N_3102,N_3080);
nand U3145 (N_3145,N_3066,N_3068);
nand U3146 (N_3146,N_3038,N_3113);
and U3147 (N_3147,N_3033,N_3060);
and U3148 (N_3148,N_3016,N_3007);
nand U3149 (N_3149,N_3101,N_3061);
nor U3150 (N_3150,N_3021,N_3087);
xnor U3151 (N_3151,N_3117,N_3094);
and U3152 (N_3152,N_3076,N_3079);
xor U3153 (N_3153,N_3069,N_3119);
nand U3154 (N_3154,N_3072,N_3041);
and U3155 (N_3155,N_3015,N_3077);
or U3156 (N_3156,N_3013,N_3000);
nor U3157 (N_3157,N_3121,N_3059);
nand U3158 (N_3158,N_3118,N_3051);
xnor U3159 (N_3159,N_3055,N_3029);
or U3160 (N_3160,N_3078,N_3123);
xnor U3161 (N_3161,N_3103,N_3106);
and U3162 (N_3162,N_3089,N_3017);
or U3163 (N_3163,N_3098,N_3036);
nand U3164 (N_3164,N_3037,N_3001);
and U3165 (N_3165,N_3086,N_3104);
nor U3166 (N_3166,N_3025,N_3096);
xor U3167 (N_3167,N_3008,N_3088);
or U3168 (N_3168,N_3035,N_3032);
nand U3169 (N_3169,N_3081,N_3044);
and U3170 (N_3170,N_3100,N_3024);
nor U3171 (N_3171,N_3046,N_3047);
xnor U3172 (N_3172,N_3114,N_3003);
or U3173 (N_3173,N_3105,N_3093);
nand U3174 (N_3174,N_3002,N_3122);
nor U3175 (N_3175,N_3030,N_3071);
xnor U3176 (N_3176,N_3073,N_3063);
or U3177 (N_3177,N_3111,N_3049);
or U3178 (N_3178,N_3043,N_3099);
and U3179 (N_3179,N_3034,N_3005);
and U3180 (N_3180,N_3090,N_3053);
nor U3181 (N_3181,N_3026,N_3042);
xor U3182 (N_3182,N_3045,N_3039);
or U3183 (N_3183,N_3006,N_3109);
nor U3184 (N_3184,N_3031,N_3083);
nand U3185 (N_3185,N_3019,N_3091);
and U3186 (N_3186,N_3112,N_3115);
xnor U3187 (N_3187,N_3084,N_3018);
nand U3188 (N_3188,N_3012,N_3071);
xor U3189 (N_3189,N_3082,N_3071);
and U3190 (N_3190,N_3089,N_3097);
nand U3191 (N_3191,N_3074,N_3124);
and U3192 (N_3192,N_3009,N_3083);
xor U3193 (N_3193,N_3071,N_3040);
or U3194 (N_3194,N_3113,N_3004);
nand U3195 (N_3195,N_3051,N_3004);
and U3196 (N_3196,N_3060,N_3117);
nor U3197 (N_3197,N_3077,N_3115);
nand U3198 (N_3198,N_3043,N_3115);
nor U3199 (N_3199,N_3075,N_3055);
and U3200 (N_3200,N_3003,N_3034);
xor U3201 (N_3201,N_3051,N_3017);
xnor U3202 (N_3202,N_3026,N_3047);
xnor U3203 (N_3203,N_3097,N_3091);
and U3204 (N_3204,N_3098,N_3118);
nor U3205 (N_3205,N_3082,N_3064);
nand U3206 (N_3206,N_3026,N_3093);
nand U3207 (N_3207,N_3033,N_3035);
or U3208 (N_3208,N_3022,N_3084);
or U3209 (N_3209,N_3072,N_3095);
xnor U3210 (N_3210,N_3042,N_3084);
and U3211 (N_3211,N_3040,N_3043);
and U3212 (N_3212,N_3008,N_3000);
nor U3213 (N_3213,N_3067,N_3077);
nand U3214 (N_3214,N_3074,N_3045);
xor U3215 (N_3215,N_3067,N_3083);
xnor U3216 (N_3216,N_3121,N_3030);
nand U3217 (N_3217,N_3119,N_3087);
and U3218 (N_3218,N_3119,N_3035);
nor U3219 (N_3219,N_3089,N_3108);
or U3220 (N_3220,N_3073,N_3062);
nor U3221 (N_3221,N_3085,N_3009);
nand U3222 (N_3222,N_3041,N_3032);
nand U3223 (N_3223,N_3110,N_3023);
xor U3224 (N_3224,N_3003,N_3026);
nand U3225 (N_3225,N_3054,N_3043);
xor U3226 (N_3226,N_3033,N_3123);
nor U3227 (N_3227,N_3111,N_3096);
nor U3228 (N_3228,N_3066,N_3009);
nor U3229 (N_3229,N_3043,N_3039);
xnor U3230 (N_3230,N_3086,N_3060);
or U3231 (N_3231,N_3017,N_3007);
or U3232 (N_3232,N_3122,N_3049);
xor U3233 (N_3233,N_3045,N_3094);
nand U3234 (N_3234,N_3078,N_3109);
and U3235 (N_3235,N_3070,N_3024);
nand U3236 (N_3236,N_3074,N_3014);
nor U3237 (N_3237,N_3023,N_3105);
xnor U3238 (N_3238,N_3100,N_3105);
nor U3239 (N_3239,N_3030,N_3120);
nand U3240 (N_3240,N_3067,N_3074);
and U3241 (N_3241,N_3009,N_3057);
or U3242 (N_3242,N_3000,N_3086);
or U3243 (N_3243,N_3117,N_3023);
nand U3244 (N_3244,N_3000,N_3122);
or U3245 (N_3245,N_3032,N_3022);
xnor U3246 (N_3246,N_3111,N_3015);
nor U3247 (N_3247,N_3023,N_3120);
nand U3248 (N_3248,N_3084,N_3049);
xor U3249 (N_3249,N_3115,N_3106);
nor U3250 (N_3250,N_3148,N_3185);
or U3251 (N_3251,N_3174,N_3193);
nor U3252 (N_3252,N_3223,N_3179);
xor U3253 (N_3253,N_3249,N_3141);
nor U3254 (N_3254,N_3143,N_3222);
nor U3255 (N_3255,N_3241,N_3172);
and U3256 (N_3256,N_3233,N_3162);
xnor U3257 (N_3257,N_3214,N_3215);
nand U3258 (N_3258,N_3213,N_3165);
or U3259 (N_3259,N_3189,N_3227);
xor U3260 (N_3260,N_3147,N_3180);
nand U3261 (N_3261,N_3211,N_3177);
and U3262 (N_3262,N_3125,N_3140);
and U3263 (N_3263,N_3191,N_3144);
and U3264 (N_3264,N_3134,N_3137);
and U3265 (N_3265,N_3200,N_3182);
xnor U3266 (N_3266,N_3132,N_3202);
and U3267 (N_3267,N_3168,N_3238);
nand U3268 (N_3268,N_3186,N_3230);
and U3269 (N_3269,N_3205,N_3212);
nor U3270 (N_3270,N_3234,N_3188);
and U3271 (N_3271,N_3232,N_3153);
and U3272 (N_3272,N_3128,N_3173);
nor U3273 (N_3273,N_3178,N_3151);
nand U3274 (N_3274,N_3210,N_3203);
and U3275 (N_3275,N_3246,N_3139);
and U3276 (N_3276,N_3175,N_3155);
nor U3277 (N_3277,N_3138,N_3240);
and U3278 (N_3278,N_3219,N_3208);
or U3279 (N_3279,N_3198,N_3192);
nand U3280 (N_3280,N_3183,N_3217);
xnor U3281 (N_3281,N_3184,N_3235);
xor U3282 (N_3282,N_3207,N_3156);
nor U3283 (N_3283,N_3194,N_3176);
and U3284 (N_3284,N_3169,N_3170);
and U3285 (N_3285,N_3161,N_3127);
nor U3286 (N_3286,N_3196,N_3149);
and U3287 (N_3287,N_3201,N_3181);
nand U3288 (N_3288,N_3199,N_3167);
xnor U3289 (N_3289,N_3160,N_3126);
nand U3290 (N_3290,N_3157,N_3142);
xor U3291 (N_3291,N_3236,N_3159);
nand U3292 (N_3292,N_3129,N_3218);
nand U3293 (N_3293,N_3231,N_3239);
nand U3294 (N_3294,N_3226,N_3237);
and U3295 (N_3295,N_3130,N_3243);
and U3296 (N_3296,N_3158,N_3146);
or U3297 (N_3297,N_3204,N_3244);
and U3298 (N_3298,N_3221,N_3229);
nor U3299 (N_3299,N_3164,N_3245);
nand U3300 (N_3300,N_3197,N_3216);
and U3301 (N_3301,N_3166,N_3145);
nor U3302 (N_3302,N_3171,N_3248);
or U3303 (N_3303,N_3195,N_3220);
xor U3304 (N_3304,N_3152,N_3131);
xnor U3305 (N_3305,N_3163,N_3206);
and U3306 (N_3306,N_3154,N_3133);
and U3307 (N_3307,N_3135,N_3224);
nand U3308 (N_3308,N_3150,N_3190);
nand U3309 (N_3309,N_3136,N_3187);
xnor U3310 (N_3310,N_3209,N_3242);
nand U3311 (N_3311,N_3228,N_3225);
and U3312 (N_3312,N_3247,N_3201);
nor U3313 (N_3313,N_3189,N_3207);
xor U3314 (N_3314,N_3133,N_3142);
and U3315 (N_3315,N_3204,N_3169);
nor U3316 (N_3316,N_3159,N_3170);
or U3317 (N_3317,N_3234,N_3127);
or U3318 (N_3318,N_3211,N_3237);
nand U3319 (N_3319,N_3227,N_3237);
xnor U3320 (N_3320,N_3224,N_3141);
or U3321 (N_3321,N_3192,N_3237);
nor U3322 (N_3322,N_3247,N_3181);
or U3323 (N_3323,N_3191,N_3246);
and U3324 (N_3324,N_3136,N_3191);
xnor U3325 (N_3325,N_3190,N_3217);
nor U3326 (N_3326,N_3227,N_3178);
and U3327 (N_3327,N_3169,N_3221);
and U3328 (N_3328,N_3161,N_3138);
nand U3329 (N_3329,N_3246,N_3184);
nor U3330 (N_3330,N_3147,N_3223);
xnor U3331 (N_3331,N_3231,N_3189);
xnor U3332 (N_3332,N_3159,N_3174);
xor U3333 (N_3333,N_3152,N_3155);
or U3334 (N_3334,N_3225,N_3227);
nand U3335 (N_3335,N_3227,N_3139);
nor U3336 (N_3336,N_3215,N_3228);
and U3337 (N_3337,N_3167,N_3237);
nand U3338 (N_3338,N_3181,N_3149);
nand U3339 (N_3339,N_3138,N_3131);
xor U3340 (N_3340,N_3211,N_3151);
nor U3341 (N_3341,N_3243,N_3181);
nand U3342 (N_3342,N_3135,N_3221);
xnor U3343 (N_3343,N_3188,N_3181);
nand U3344 (N_3344,N_3173,N_3230);
nand U3345 (N_3345,N_3134,N_3217);
nor U3346 (N_3346,N_3172,N_3188);
or U3347 (N_3347,N_3217,N_3193);
and U3348 (N_3348,N_3227,N_3233);
or U3349 (N_3349,N_3173,N_3224);
and U3350 (N_3350,N_3160,N_3225);
and U3351 (N_3351,N_3175,N_3203);
or U3352 (N_3352,N_3214,N_3243);
and U3353 (N_3353,N_3187,N_3199);
xnor U3354 (N_3354,N_3166,N_3226);
and U3355 (N_3355,N_3215,N_3133);
nand U3356 (N_3356,N_3181,N_3174);
or U3357 (N_3357,N_3231,N_3234);
nand U3358 (N_3358,N_3218,N_3196);
and U3359 (N_3359,N_3213,N_3192);
nand U3360 (N_3360,N_3234,N_3235);
nand U3361 (N_3361,N_3195,N_3214);
or U3362 (N_3362,N_3180,N_3171);
or U3363 (N_3363,N_3199,N_3154);
and U3364 (N_3364,N_3196,N_3158);
or U3365 (N_3365,N_3154,N_3153);
xnor U3366 (N_3366,N_3142,N_3128);
or U3367 (N_3367,N_3222,N_3242);
or U3368 (N_3368,N_3138,N_3126);
or U3369 (N_3369,N_3126,N_3185);
nor U3370 (N_3370,N_3155,N_3249);
nand U3371 (N_3371,N_3191,N_3227);
nor U3372 (N_3372,N_3226,N_3205);
nand U3373 (N_3373,N_3234,N_3183);
xnor U3374 (N_3374,N_3142,N_3148);
nor U3375 (N_3375,N_3338,N_3362);
or U3376 (N_3376,N_3351,N_3282);
or U3377 (N_3377,N_3353,N_3324);
or U3378 (N_3378,N_3330,N_3369);
nand U3379 (N_3379,N_3283,N_3310);
and U3380 (N_3380,N_3350,N_3254);
or U3381 (N_3381,N_3309,N_3257);
or U3382 (N_3382,N_3336,N_3298);
nor U3383 (N_3383,N_3302,N_3366);
nor U3384 (N_3384,N_3279,N_3270);
nor U3385 (N_3385,N_3335,N_3346);
or U3386 (N_3386,N_3323,N_3344);
and U3387 (N_3387,N_3370,N_3269);
and U3388 (N_3388,N_3267,N_3371);
nor U3389 (N_3389,N_3295,N_3343);
nor U3390 (N_3390,N_3311,N_3286);
or U3391 (N_3391,N_3329,N_3271);
nor U3392 (N_3392,N_3304,N_3345);
xor U3393 (N_3393,N_3327,N_3328);
nand U3394 (N_3394,N_3265,N_3352);
and U3395 (N_3395,N_3273,N_3252);
and U3396 (N_3396,N_3299,N_3320);
nand U3397 (N_3397,N_3349,N_3272);
nor U3398 (N_3398,N_3276,N_3290);
nand U3399 (N_3399,N_3359,N_3367);
and U3400 (N_3400,N_3300,N_3285);
or U3401 (N_3401,N_3342,N_3303);
nand U3402 (N_3402,N_3301,N_3315);
nor U3403 (N_3403,N_3284,N_3268);
nor U3404 (N_3404,N_3339,N_3374);
nor U3405 (N_3405,N_3275,N_3334);
xor U3406 (N_3406,N_3288,N_3280);
nand U3407 (N_3407,N_3251,N_3259);
xnor U3408 (N_3408,N_3314,N_3364);
nand U3409 (N_3409,N_3331,N_3337);
and U3410 (N_3410,N_3264,N_3358);
xnor U3411 (N_3411,N_3373,N_3355);
or U3412 (N_3412,N_3289,N_3363);
nand U3413 (N_3413,N_3360,N_3256);
and U3414 (N_3414,N_3317,N_3326);
or U3415 (N_3415,N_3263,N_3250);
nor U3416 (N_3416,N_3322,N_3294);
or U3417 (N_3417,N_3372,N_3340);
xnor U3418 (N_3418,N_3361,N_3316);
nor U3419 (N_3419,N_3356,N_3365);
nor U3420 (N_3420,N_3321,N_3306);
or U3421 (N_3421,N_3319,N_3368);
and U3422 (N_3422,N_3262,N_3347);
xor U3423 (N_3423,N_3325,N_3253);
and U3424 (N_3424,N_3287,N_3278);
xor U3425 (N_3425,N_3274,N_3260);
nor U3426 (N_3426,N_3266,N_3258);
and U3427 (N_3427,N_3305,N_3296);
nor U3428 (N_3428,N_3293,N_3261);
and U3429 (N_3429,N_3341,N_3354);
and U3430 (N_3430,N_3357,N_3308);
or U3431 (N_3431,N_3291,N_3277);
nand U3432 (N_3432,N_3333,N_3313);
or U3433 (N_3433,N_3255,N_3318);
nand U3434 (N_3434,N_3348,N_3281);
and U3435 (N_3435,N_3297,N_3312);
xnor U3436 (N_3436,N_3292,N_3307);
nand U3437 (N_3437,N_3332,N_3298);
nor U3438 (N_3438,N_3304,N_3306);
and U3439 (N_3439,N_3290,N_3263);
xnor U3440 (N_3440,N_3289,N_3264);
or U3441 (N_3441,N_3284,N_3303);
or U3442 (N_3442,N_3314,N_3341);
and U3443 (N_3443,N_3261,N_3297);
xnor U3444 (N_3444,N_3359,N_3358);
nand U3445 (N_3445,N_3252,N_3306);
xnor U3446 (N_3446,N_3299,N_3305);
xnor U3447 (N_3447,N_3350,N_3309);
or U3448 (N_3448,N_3290,N_3354);
nor U3449 (N_3449,N_3299,N_3294);
nand U3450 (N_3450,N_3293,N_3284);
nor U3451 (N_3451,N_3250,N_3296);
and U3452 (N_3452,N_3259,N_3374);
nand U3453 (N_3453,N_3276,N_3284);
nand U3454 (N_3454,N_3352,N_3326);
or U3455 (N_3455,N_3335,N_3268);
nand U3456 (N_3456,N_3276,N_3269);
nor U3457 (N_3457,N_3313,N_3374);
or U3458 (N_3458,N_3295,N_3340);
xor U3459 (N_3459,N_3313,N_3341);
and U3460 (N_3460,N_3307,N_3286);
or U3461 (N_3461,N_3277,N_3281);
and U3462 (N_3462,N_3297,N_3346);
nor U3463 (N_3463,N_3259,N_3339);
xnor U3464 (N_3464,N_3293,N_3325);
or U3465 (N_3465,N_3271,N_3292);
nand U3466 (N_3466,N_3350,N_3253);
and U3467 (N_3467,N_3367,N_3327);
or U3468 (N_3468,N_3348,N_3333);
nand U3469 (N_3469,N_3258,N_3263);
nor U3470 (N_3470,N_3347,N_3355);
or U3471 (N_3471,N_3358,N_3273);
or U3472 (N_3472,N_3351,N_3269);
and U3473 (N_3473,N_3369,N_3326);
and U3474 (N_3474,N_3295,N_3364);
xor U3475 (N_3475,N_3277,N_3295);
nor U3476 (N_3476,N_3306,N_3266);
xnor U3477 (N_3477,N_3293,N_3316);
and U3478 (N_3478,N_3335,N_3302);
or U3479 (N_3479,N_3347,N_3338);
xor U3480 (N_3480,N_3297,N_3257);
or U3481 (N_3481,N_3354,N_3312);
xor U3482 (N_3482,N_3284,N_3300);
nor U3483 (N_3483,N_3326,N_3351);
and U3484 (N_3484,N_3326,N_3346);
and U3485 (N_3485,N_3263,N_3320);
nand U3486 (N_3486,N_3318,N_3355);
nor U3487 (N_3487,N_3332,N_3259);
xor U3488 (N_3488,N_3335,N_3354);
nor U3489 (N_3489,N_3371,N_3333);
nor U3490 (N_3490,N_3271,N_3284);
or U3491 (N_3491,N_3288,N_3353);
or U3492 (N_3492,N_3362,N_3277);
xor U3493 (N_3493,N_3349,N_3255);
xnor U3494 (N_3494,N_3341,N_3273);
nand U3495 (N_3495,N_3348,N_3275);
and U3496 (N_3496,N_3286,N_3270);
and U3497 (N_3497,N_3293,N_3360);
and U3498 (N_3498,N_3348,N_3360);
or U3499 (N_3499,N_3280,N_3287);
nor U3500 (N_3500,N_3461,N_3378);
and U3501 (N_3501,N_3494,N_3493);
xnor U3502 (N_3502,N_3411,N_3467);
and U3503 (N_3503,N_3431,N_3426);
nor U3504 (N_3504,N_3403,N_3386);
nor U3505 (N_3505,N_3457,N_3414);
xnor U3506 (N_3506,N_3387,N_3384);
nor U3507 (N_3507,N_3498,N_3392);
nand U3508 (N_3508,N_3382,N_3441);
and U3509 (N_3509,N_3377,N_3473);
nand U3510 (N_3510,N_3479,N_3475);
nand U3511 (N_3511,N_3409,N_3385);
or U3512 (N_3512,N_3442,N_3471);
or U3513 (N_3513,N_3376,N_3396);
xor U3514 (N_3514,N_3481,N_3448);
xor U3515 (N_3515,N_3410,N_3460);
and U3516 (N_3516,N_3398,N_3435);
and U3517 (N_3517,N_3381,N_3499);
or U3518 (N_3518,N_3463,N_3459);
nand U3519 (N_3519,N_3452,N_3383);
nor U3520 (N_3520,N_3421,N_3379);
and U3521 (N_3521,N_3464,N_3486);
nand U3522 (N_3522,N_3478,N_3408);
xnor U3523 (N_3523,N_3497,N_3413);
or U3524 (N_3524,N_3492,N_3434);
or U3525 (N_3525,N_3454,N_3439);
or U3526 (N_3526,N_3405,N_3477);
xor U3527 (N_3527,N_3469,N_3428);
or U3528 (N_3528,N_3380,N_3404);
or U3529 (N_3529,N_3484,N_3445);
nor U3530 (N_3530,N_3406,N_3433);
and U3531 (N_3531,N_3446,N_3489);
nor U3532 (N_3532,N_3496,N_3491);
nand U3533 (N_3533,N_3468,N_3466);
xnor U3534 (N_3534,N_3447,N_3420);
xnor U3535 (N_3535,N_3375,N_3402);
and U3536 (N_3536,N_3470,N_3423);
nor U3537 (N_3537,N_3395,N_3417);
xnor U3538 (N_3538,N_3424,N_3440);
xnor U3539 (N_3539,N_3400,N_3432);
xor U3540 (N_3540,N_3399,N_3488);
nor U3541 (N_3541,N_3389,N_3436);
and U3542 (N_3542,N_3451,N_3485);
xor U3543 (N_3543,N_3425,N_3449);
nand U3544 (N_3544,N_3462,N_3437);
nor U3545 (N_3545,N_3495,N_3450);
nand U3546 (N_3546,N_3394,N_3474);
or U3547 (N_3547,N_3391,N_3444);
and U3548 (N_3548,N_3429,N_3388);
xnor U3549 (N_3549,N_3438,N_3482);
nor U3550 (N_3550,N_3393,N_3453);
and U3551 (N_3551,N_3458,N_3476);
xnor U3552 (N_3552,N_3415,N_3412);
nand U3553 (N_3553,N_3419,N_3472);
nor U3554 (N_3554,N_3397,N_3418);
or U3555 (N_3555,N_3465,N_3390);
nor U3556 (N_3556,N_3443,N_3480);
xnor U3557 (N_3557,N_3490,N_3456);
nand U3558 (N_3558,N_3487,N_3427);
nor U3559 (N_3559,N_3416,N_3430);
nand U3560 (N_3560,N_3483,N_3401);
and U3561 (N_3561,N_3455,N_3422);
or U3562 (N_3562,N_3407,N_3385);
or U3563 (N_3563,N_3499,N_3417);
nand U3564 (N_3564,N_3481,N_3442);
nand U3565 (N_3565,N_3434,N_3410);
or U3566 (N_3566,N_3406,N_3425);
nand U3567 (N_3567,N_3395,N_3378);
nand U3568 (N_3568,N_3432,N_3404);
nor U3569 (N_3569,N_3399,N_3436);
xor U3570 (N_3570,N_3407,N_3388);
nor U3571 (N_3571,N_3380,N_3453);
or U3572 (N_3572,N_3445,N_3462);
xnor U3573 (N_3573,N_3432,N_3384);
xnor U3574 (N_3574,N_3442,N_3455);
xnor U3575 (N_3575,N_3461,N_3498);
and U3576 (N_3576,N_3409,N_3382);
or U3577 (N_3577,N_3414,N_3396);
nand U3578 (N_3578,N_3457,N_3455);
xor U3579 (N_3579,N_3407,N_3465);
xnor U3580 (N_3580,N_3449,N_3397);
or U3581 (N_3581,N_3479,N_3494);
or U3582 (N_3582,N_3476,N_3448);
nand U3583 (N_3583,N_3445,N_3482);
nand U3584 (N_3584,N_3492,N_3497);
nand U3585 (N_3585,N_3468,N_3375);
and U3586 (N_3586,N_3478,N_3481);
xor U3587 (N_3587,N_3485,N_3442);
xor U3588 (N_3588,N_3428,N_3451);
and U3589 (N_3589,N_3418,N_3435);
and U3590 (N_3590,N_3393,N_3429);
nand U3591 (N_3591,N_3480,N_3429);
and U3592 (N_3592,N_3417,N_3473);
or U3593 (N_3593,N_3449,N_3435);
nand U3594 (N_3594,N_3386,N_3492);
or U3595 (N_3595,N_3406,N_3490);
xnor U3596 (N_3596,N_3460,N_3499);
xnor U3597 (N_3597,N_3471,N_3485);
xnor U3598 (N_3598,N_3478,N_3490);
and U3599 (N_3599,N_3414,N_3451);
nor U3600 (N_3600,N_3410,N_3489);
and U3601 (N_3601,N_3459,N_3456);
and U3602 (N_3602,N_3486,N_3483);
or U3603 (N_3603,N_3497,N_3475);
nor U3604 (N_3604,N_3382,N_3460);
and U3605 (N_3605,N_3383,N_3436);
and U3606 (N_3606,N_3487,N_3470);
or U3607 (N_3607,N_3381,N_3498);
or U3608 (N_3608,N_3473,N_3443);
nand U3609 (N_3609,N_3454,N_3463);
or U3610 (N_3610,N_3468,N_3478);
and U3611 (N_3611,N_3437,N_3432);
nand U3612 (N_3612,N_3494,N_3495);
or U3613 (N_3613,N_3493,N_3412);
or U3614 (N_3614,N_3379,N_3424);
or U3615 (N_3615,N_3386,N_3425);
nand U3616 (N_3616,N_3380,N_3479);
or U3617 (N_3617,N_3448,N_3423);
and U3618 (N_3618,N_3497,N_3416);
and U3619 (N_3619,N_3475,N_3444);
nand U3620 (N_3620,N_3426,N_3468);
nand U3621 (N_3621,N_3406,N_3485);
nand U3622 (N_3622,N_3415,N_3405);
or U3623 (N_3623,N_3457,N_3473);
nand U3624 (N_3624,N_3466,N_3381);
xnor U3625 (N_3625,N_3606,N_3605);
and U3626 (N_3626,N_3624,N_3560);
nor U3627 (N_3627,N_3591,N_3597);
or U3628 (N_3628,N_3505,N_3547);
nand U3629 (N_3629,N_3557,N_3564);
nand U3630 (N_3630,N_3534,N_3509);
nor U3631 (N_3631,N_3531,N_3510);
nor U3632 (N_3632,N_3555,N_3541);
or U3633 (N_3633,N_3553,N_3562);
and U3634 (N_3634,N_3586,N_3568);
or U3635 (N_3635,N_3528,N_3575);
and U3636 (N_3636,N_3599,N_3603);
or U3637 (N_3637,N_3621,N_3592);
and U3638 (N_3638,N_3532,N_3590);
nand U3639 (N_3639,N_3604,N_3596);
nor U3640 (N_3640,N_3556,N_3537);
or U3641 (N_3641,N_3538,N_3561);
or U3642 (N_3642,N_3558,N_3578);
and U3643 (N_3643,N_3623,N_3530);
or U3644 (N_3644,N_3551,N_3559);
or U3645 (N_3645,N_3580,N_3594);
nor U3646 (N_3646,N_3513,N_3588);
nand U3647 (N_3647,N_3540,N_3506);
and U3648 (N_3648,N_3573,N_3529);
or U3649 (N_3649,N_3614,N_3527);
or U3650 (N_3650,N_3546,N_3579);
or U3651 (N_3651,N_3502,N_3549);
nor U3652 (N_3652,N_3593,N_3598);
xor U3653 (N_3653,N_3507,N_3525);
nand U3654 (N_3654,N_3620,N_3601);
nand U3655 (N_3655,N_3571,N_3518);
or U3656 (N_3656,N_3581,N_3539);
nand U3657 (N_3657,N_3608,N_3609);
xor U3658 (N_3658,N_3512,N_3610);
and U3659 (N_3659,N_3521,N_3611);
xor U3660 (N_3660,N_3566,N_3607);
xor U3661 (N_3661,N_3511,N_3504);
xor U3662 (N_3662,N_3552,N_3517);
or U3663 (N_3663,N_3570,N_3577);
xor U3664 (N_3664,N_3500,N_3584);
nand U3665 (N_3665,N_3548,N_3613);
and U3666 (N_3666,N_3543,N_3522);
and U3667 (N_3667,N_3563,N_3526);
nor U3668 (N_3668,N_3612,N_3545);
nor U3669 (N_3669,N_3516,N_3501);
and U3670 (N_3670,N_3542,N_3508);
nand U3671 (N_3671,N_3617,N_3587);
or U3672 (N_3672,N_3589,N_3536);
nand U3673 (N_3673,N_3583,N_3515);
xnor U3674 (N_3674,N_3544,N_3618);
and U3675 (N_3675,N_3582,N_3533);
xor U3676 (N_3676,N_3554,N_3569);
or U3677 (N_3677,N_3520,N_3600);
nand U3678 (N_3678,N_3585,N_3524);
and U3679 (N_3679,N_3567,N_3619);
and U3680 (N_3680,N_3565,N_3535);
nand U3681 (N_3681,N_3519,N_3572);
and U3682 (N_3682,N_3595,N_3622);
or U3683 (N_3683,N_3503,N_3602);
or U3684 (N_3684,N_3514,N_3574);
xor U3685 (N_3685,N_3615,N_3616);
nor U3686 (N_3686,N_3523,N_3550);
nor U3687 (N_3687,N_3576,N_3543);
nand U3688 (N_3688,N_3531,N_3596);
nand U3689 (N_3689,N_3525,N_3558);
nand U3690 (N_3690,N_3509,N_3546);
nand U3691 (N_3691,N_3592,N_3619);
or U3692 (N_3692,N_3518,N_3612);
xor U3693 (N_3693,N_3523,N_3575);
or U3694 (N_3694,N_3604,N_3584);
nand U3695 (N_3695,N_3582,N_3591);
and U3696 (N_3696,N_3511,N_3608);
or U3697 (N_3697,N_3521,N_3590);
nor U3698 (N_3698,N_3623,N_3621);
nor U3699 (N_3699,N_3511,N_3619);
nand U3700 (N_3700,N_3589,N_3586);
and U3701 (N_3701,N_3573,N_3616);
nor U3702 (N_3702,N_3573,N_3567);
nand U3703 (N_3703,N_3538,N_3542);
and U3704 (N_3704,N_3621,N_3588);
nand U3705 (N_3705,N_3502,N_3517);
nand U3706 (N_3706,N_3537,N_3515);
nor U3707 (N_3707,N_3587,N_3591);
nand U3708 (N_3708,N_3515,N_3539);
xnor U3709 (N_3709,N_3538,N_3599);
xor U3710 (N_3710,N_3612,N_3582);
or U3711 (N_3711,N_3593,N_3610);
and U3712 (N_3712,N_3622,N_3562);
and U3713 (N_3713,N_3607,N_3576);
nand U3714 (N_3714,N_3527,N_3559);
xor U3715 (N_3715,N_3533,N_3546);
xnor U3716 (N_3716,N_3619,N_3503);
nand U3717 (N_3717,N_3559,N_3599);
or U3718 (N_3718,N_3584,N_3547);
and U3719 (N_3719,N_3549,N_3575);
nand U3720 (N_3720,N_3618,N_3583);
or U3721 (N_3721,N_3518,N_3528);
nand U3722 (N_3722,N_3623,N_3555);
nor U3723 (N_3723,N_3517,N_3545);
xnor U3724 (N_3724,N_3520,N_3621);
xnor U3725 (N_3725,N_3525,N_3503);
xor U3726 (N_3726,N_3542,N_3621);
xor U3727 (N_3727,N_3537,N_3598);
nand U3728 (N_3728,N_3522,N_3621);
and U3729 (N_3729,N_3584,N_3513);
nand U3730 (N_3730,N_3542,N_3548);
xnor U3731 (N_3731,N_3547,N_3575);
and U3732 (N_3732,N_3524,N_3596);
xor U3733 (N_3733,N_3590,N_3608);
nor U3734 (N_3734,N_3552,N_3524);
nand U3735 (N_3735,N_3529,N_3606);
nor U3736 (N_3736,N_3513,N_3561);
and U3737 (N_3737,N_3612,N_3530);
and U3738 (N_3738,N_3624,N_3576);
nor U3739 (N_3739,N_3592,N_3571);
nand U3740 (N_3740,N_3539,N_3612);
or U3741 (N_3741,N_3549,N_3584);
nand U3742 (N_3742,N_3618,N_3615);
nor U3743 (N_3743,N_3620,N_3554);
xnor U3744 (N_3744,N_3539,N_3563);
nand U3745 (N_3745,N_3607,N_3512);
nand U3746 (N_3746,N_3582,N_3550);
or U3747 (N_3747,N_3598,N_3599);
xor U3748 (N_3748,N_3533,N_3504);
nand U3749 (N_3749,N_3512,N_3563);
xor U3750 (N_3750,N_3742,N_3684);
xnor U3751 (N_3751,N_3645,N_3749);
nor U3752 (N_3752,N_3693,N_3648);
xnor U3753 (N_3753,N_3679,N_3660);
xnor U3754 (N_3754,N_3722,N_3686);
nand U3755 (N_3755,N_3746,N_3747);
or U3756 (N_3756,N_3731,N_3650);
or U3757 (N_3757,N_3631,N_3717);
and U3758 (N_3758,N_3720,N_3744);
nor U3759 (N_3759,N_3732,N_3688);
nor U3760 (N_3760,N_3735,N_3740);
and U3761 (N_3761,N_3713,N_3625);
and U3762 (N_3762,N_3656,N_3672);
nor U3763 (N_3763,N_3670,N_3711);
xnor U3764 (N_3764,N_3638,N_3729);
nor U3765 (N_3765,N_3632,N_3727);
xor U3766 (N_3766,N_3745,N_3704);
xor U3767 (N_3767,N_3642,N_3741);
nand U3768 (N_3768,N_3689,N_3721);
or U3769 (N_3769,N_3698,N_3634);
xnor U3770 (N_3770,N_3659,N_3702);
nand U3771 (N_3771,N_3666,N_3633);
or U3772 (N_3772,N_3635,N_3730);
xor U3773 (N_3773,N_3664,N_3676);
nor U3774 (N_3774,N_3671,N_3738);
or U3775 (N_3775,N_3630,N_3691);
xnor U3776 (N_3776,N_3748,N_3674);
or U3777 (N_3777,N_3651,N_3627);
nor U3778 (N_3778,N_3685,N_3724);
nor U3779 (N_3779,N_3703,N_3667);
nand U3780 (N_3780,N_3718,N_3716);
nand U3781 (N_3781,N_3626,N_3681);
and U3782 (N_3782,N_3641,N_3663);
and U3783 (N_3783,N_3700,N_3669);
and U3784 (N_3784,N_3643,N_3712);
nand U3785 (N_3785,N_3726,N_3675);
nand U3786 (N_3786,N_3714,N_3706);
and U3787 (N_3787,N_3723,N_3636);
xor U3788 (N_3788,N_3637,N_3709);
and U3789 (N_3789,N_3707,N_3639);
or U3790 (N_3790,N_3739,N_3658);
or U3791 (N_3791,N_3733,N_3710);
nor U3792 (N_3792,N_3647,N_3743);
nor U3793 (N_3793,N_3653,N_3725);
or U3794 (N_3794,N_3661,N_3673);
and U3795 (N_3795,N_3690,N_3646);
and U3796 (N_3796,N_3655,N_3644);
or U3797 (N_3797,N_3680,N_3677);
or U3798 (N_3798,N_3695,N_3701);
nor U3799 (N_3799,N_3736,N_3652);
or U3800 (N_3800,N_3697,N_3629);
or U3801 (N_3801,N_3728,N_3682);
nor U3802 (N_3802,N_3662,N_3654);
nand U3803 (N_3803,N_3715,N_3640);
nand U3804 (N_3804,N_3665,N_3719);
and U3805 (N_3805,N_3668,N_3734);
or U3806 (N_3806,N_3699,N_3708);
nand U3807 (N_3807,N_3687,N_3678);
or U3808 (N_3808,N_3657,N_3694);
and U3809 (N_3809,N_3692,N_3683);
nand U3810 (N_3810,N_3737,N_3649);
and U3811 (N_3811,N_3696,N_3705);
nor U3812 (N_3812,N_3628,N_3730);
or U3813 (N_3813,N_3646,N_3689);
and U3814 (N_3814,N_3664,N_3626);
xnor U3815 (N_3815,N_3725,N_3626);
nor U3816 (N_3816,N_3660,N_3630);
nor U3817 (N_3817,N_3642,N_3654);
nor U3818 (N_3818,N_3736,N_3648);
and U3819 (N_3819,N_3682,N_3699);
nor U3820 (N_3820,N_3701,N_3726);
xnor U3821 (N_3821,N_3633,N_3715);
nand U3822 (N_3822,N_3702,N_3673);
or U3823 (N_3823,N_3699,N_3684);
and U3824 (N_3824,N_3629,N_3726);
nand U3825 (N_3825,N_3662,N_3678);
nor U3826 (N_3826,N_3631,N_3730);
nor U3827 (N_3827,N_3728,N_3648);
nor U3828 (N_3828,N_3649,N_3661);
and U3829 (N_3829,N_3679,N_3749);
xor U3830 (N_3830,N_3740,N_3666);
nand U3831 (N_3831,N_3662,N_3642);
nand U3832 (N_3832,N_3681,N_3627);
or U3833 (N_3833,N_3675,N_3693);
and U3834 (N_3834,N_3672,N_3738);
or U3835 (N_3835,N_3699,N_3691);
or U3836 (N_3836,N_3625,N_3632);
or U3837 (N_3837,N_3692,N_3748);
or U3838 (N_3838,N_3656,N_3699);
nor U3839 (N_3839,N_3713,N_3685);
or U3840 (N_3840,N_3639,N_3636);
and U3841 (N_3841,N_3722,N_3632);
or U3842 (N_3842,N_3722,N_3626);
nor U3843 (N_3843,N_3742,N_3749);
nand U3844 (N_3844,N_3706,N_3699);
or U3845 (N_3845,N_3700,N_3659);
or U3846 (N_3846,N_3633,N_3724);
and U3847 (N_3847,N_3674,N_3721);
and U3848 (N_3848,N_3643,N_3743);
nor U3849 (N_3849,N_3730,N_3746);
or U3850 (N_3850,N_3676,N_3646);
and U3851 (N_3851,N_3650,N_3665);
or U3852 (N_3852,N_3747,N_3708);
or U3853 (N_3853,N_3679,N_3721);
nor U3854 (N_3854,N_3649,N_3646);
or U3855 (N_3855,N_3725,N_3701);
nor U3856 (N_3856,N_3717,N_3719);
xor U3857 (N_3857,N_3688,N_3679);
nand U3858 (N_3858,N_3747,N_3716);
xnor U3859 (N_3859,N_3742,N_3678);
or U3860 (N_3860,N_3744,N_3705);
nor U3861 (N_3861,N_3710,N_3672);
and U3862 (N_3862,N_3685,N_3714);
nand U3863 (N_3863,N_3656,N_3690);
or U3864 (N_3864,N_3655,N_3653);
xor U3865 (N_3865,N_3687,N_3701);
nand U3866 (N_3866,N_3657,N_3727);
xor U3867 (N_3867,N_3657,N_3704);
and U3868 (N_3868,N_3725,N_3727);
and U3869 (N_3869,N_3703,N_3687);
and U3870 (N_3870,N_3746,N_3686);
nor U3871 (N_3871,N_3684,N_3741);
nor U3872 (N_3872,N_3704,N_3655);
nand U3873 (N_3873,N_3744,N_3696);
nor U3874 (N_3874,N_3743,N_3630);
and U3875 (N_3875,N_3867,N_3836);
nand U3876 (N_3876,N_3837,N_3775);
and U3877 (N_3877,N_3797,N_3794);
and U3878 (N_3878,N_3862,N_3824);
nor U3879 (N_3879,N_3785,N_3786);
or U3880 (N_3880,N_3851,N_3872);
xnor U3881 (N_3881,N_3802,N_3774);
nor U3882 (N_3882,N_3776,N_3842);
xor U3883 (N_3883,N_3798,N_3750);
and U3884 (N_3884,N_3827,N_3765);
xnor U3885 (N_3885,N_3820,N_3865);
or U3886 (N_3886,N_3783,N_3792);
xor U3887 (N_3887,N_3815,N_3859);
or U3888 (N_3888,N_3873,N_3844);
and U3889 (N_3889,N_3796,N_3809);
or U3890 (N_3890,N_3808,N_3868);
or U3891 (N_3891,N_3766,N_3850);
xnor U3892 (N_3892,N_3759,N_3816);
nor U3893 (N_3893,N_3830,N_3860);
or U3894 (N_3894,N_3769,N_3763);
and U3895 (N_3895,N_3854,N_3788);
nor U3896 (N_3896,N_3861,N_3782);
and U3897 (N_3897,N_3840,N_3807);
xnor U3898 (N_3898,N_3857,N_3787);
nor U3899 (N_3899,N_3781,N_3849);
and U3900 (N_3900,N_3864,N_3777);
and U3901 (N_3901,N_3845,N_3767);
and U3902 (N_3902,N_3812,N_3773);
nor U3903 (N_3903,N_3858,N_3762);
xor U3904 (N_3904,N_3805,N_3871);
and U3905 (N_3905,N_3795,N_3822);
nor U3906 (N_3906,N_3778,N_3801);
nor U3907 (N_3907,N_3770,N_3853);
or U3908 (N_3908,N_3791,N_3757);
and U3909 (N_3909,N_3847,N_3814);
and U3910 (N_3910,N_3768,N_3833);
xnor U3911 (N_3911,N_3841,N_3838);
xor U3912 (N_3912,N_3752,N_3826);
nor U3913 (N_3913,N_3761,N_3772);
xnor U3914 (N_3914,N_3751,N_3832);
and U3915 (N_3915,N_3758,N_3821);
nand U3916 (N_3916,N_3779,N_3793);
and U3917 (N_3917,N_3754,N_3784);
and U3918 (N_3918,N_3818,N_3771);
and U3919 (N_3919,N_3848,N_3804);
and U3920 (N_3920,N_3831,N_3823);
xnor U3921 (N_3921,N_3817,N_3839);
and U3922 (N_3922,N_3790,N_3800);
nand U3923 (N_3923,N_3852,N_3870);
xnor U3924 (N_3924,N_3813,N_3835);
and U3925 (N_3925,N_3764,N_3825);
or U3926 (N_3926,N_3856,N_3756);
and U3927 (N_3927,N_3869,N_3806);
nand U3928 (N_3928,N_3855,N_3874);
or U3929 (N_3929,N_3760,N_3811);
or U3930 (N_3930,N_3803,N_3866);
xor U3931 (N_3931,N_3789,N_3810);
nand U3932 (N_3932,N_3829,N_3755);
xor U3933 (N_3933,N_3819,N_3846);
nor U3934 (N_3934,N_3828,N_3834);
or U3935 (N_3935,N_3843,N_3799);
nor U3936 (N_3936,N_3863,N_3780);
xor U3937 (N_3937,N_3753,N_3857);
or U3938 (N_3938,N_3867,N_3800);
xor U3939 (N_3939,N_3823,N_3817);
xor U3940 (N_3940,N_3822,N_3792);
nor U3941 (N_3941,N_3827,N_3754);
xor U3942 (N_3942,N_3825,N_3873);
and U3943 (N_3943,N_3779,N_3845);
xor U3944 (N_3944,N_3849,N_3872);
nor U3945 (N_3945,N_3797,N_3857);
xnor U3946 (N_3946,N_3798,N_3818);
nor U3947 (N_3947,N_3855,N_3840);
or U3948 (N_3948,N_3751,N_3846);
or U3949 (N_3949,N_3795,N_3873);
nor U3950 (N_3950,N_3840,N_3837);
nor U3951 (N_3951,N_3814,N_3851);
xor U3952 (N_3952,N_3832,N_3817);
xor U3953 (N_3953,N_3817,N_3774);
xor U3954 (N_3954,N_3847,N_3807);
or U3955 (N_3955,N_3824,N_3818);
nand U3956 (N_3956,N_3759,N_3855);
nand U3957 (N_3957,N_3769,N_3797);
and U3958 (N_3958,N_3791,N_3776);
or U3959 (N_3959,N_3760,N_3755);
or U3960 (N_3960,N_3753,N_3803);
nand U3961 (N_3961,N_3763,N_3787);
and U3962 (N_3962,N_3786,N_3788);
or U3963 (N_3963,N_3862,N_3783);
xnor U3964 (N_3964,N_3758,N_3818);
xor U3965 (N_3965,N_3854,N_3858);
nor U3966 (N_3966,N_3802,N_3820);
xnor U3967 (N_3967,N_3874,N_3775);
nand U3968 (N_3968,N_3781,N_3777);
or U3969 (N_3969,N_3793,N_3801);
nand U3970 (N_3970,N_3834,N_3827);
nor U3971 (N_3971,N_3828,N_3820);
nor U3972 (N_3972,N_3784,N_3766);
xor U3973 (N_3973,N_3789,N_3867);
nor U3974 (N_3974,N_3776,N_3802);
nor U3975 (N_3975,N_3761,N_3804);
xnor U3976 (N_3976,N_3751,N_3755);
and U3977 (N_3977,N_3837,N_3843);
and U3978 (N_3978,N_3827,N_3802);
nand U3979 (N_3979,N_3761,N_3780);
nand U3980 (N_3980,N_3871,N_3790);
nor U3981 (N_3981,N_3796,N_3869);
and U3982 (N_3982,N_3785,N_3853);
and U3983 (N_3983,N_3776,N_3833);
xnor U3984 (N_3984,N_3827,N_3848);
xor U3985 (N_3985,N_3766,N_3820);
nand U3986 (N_3986,N_3788,N_3763);
or U3987 (N_3987,N_3761,N_3806);
or U3988 (N_3988,N_3815,N_3789);
nor U3989 (N_3989,N_3846,N_3789);
or U3990 (N_3990,N_3754,N_3842);
and U3991 (N_3991,N_3835,N_3821);
nor U3992 (N_3992,N_3846,N_3824);
nor U3993 (N_3993,N_3829,N_3832);
nor U3994 (N_3994,N_3780,N_3812);
or U3995 (N_3995,N_3785,N_3784);
and U3996 (N_3996,N_3783,N_3855);
xnor U3997 (N_3997,N_3826,N_3873);
and U3998 (N_3998,N_3834,N_3759);
and U3999 (N_3999,N_3856,N_3844);
xor U4000 (N_4000,N_3986,N_3877);
and U4001 (N_4001,N_3991,N_3969);
and U4002 (N_4002,N_3972,N_3994);
or U4003 (N_4003,N_3882,N_3927);
and U4004 (N_4004,N_3962,N_3906);
and U4005 (N_4005,N_3967,N_3913);
nand U4006 (N_4006,N_3903,N_3957);
nand U4007 (N_4007,N_3895,N_3911);
or U4008 (N_4008,N_3908,N_3975);
xnor U4009 (N_4009,N_3883,N_3936);
nor U4010 (N_4010,N_3892,N_3881);
and U4011 (N_4011,N_3964,N_3995);
and U4012 (N_4012,N_3978,N_3880);
nor U4013 (N_4013,N_3989,N_3944);
nor U4014 (N_4014,N_3938,N_3947);
xnor U4015 (N_4015,N_3876,N_3940);
xor U4016 (N_4016,N_3909,N_3937);
and U4017 (N_4017,N_3985,N_3907);
xor U4018 (N_4018,N_3951,N_3891);
nor U4019 (N_4019,N_3902,N_3992);
or U4020 (N_4020,N_3982,N_3916);
xnor U4021 (N_4021,N_3959,N_3878);
xor U4022 (N_4022,N_3875,N_3996);
nor U4023 (N_4023,N_3950,N_3946);
nand U4024 (N_4024,N_3900,N_3948);
nand U4025 (N_4025,N_3918,N_3983);
xnor U4026 (N_4026,N_3912,N_3988);
or U4027 (N_4027,N_3889,N_3954);
nand U4028 (N_4028,N_3921,N_3981);
nand U4029 (N_4029,N_3939,N_3887);
nand U4030 (N_4030,N_3901,N_3941);
or U4031 (N_4031,N_3897,N_3929);
nor U4032 (N_4032,N_3885,N_3976);
xor U4033 (N_4033,N_3935,N_3953);
and U4034 (N_4034,N_3990,N_3993);
nand U4035 (N_4035,N_3893,N_3915);
and U4036 (N_4036,N_3958,N_3949);
and U4037 (N_4037,N_3890,N_3961);
nor U4038 (N_4038,N_3971,N_3917);
and U4039 (N_4039,N_3919,N_3888);
nand U4040 (N_4040,N_3930,N_3984);
nand U4041 (N_4041,N_3965,N_3898);
nand U4042 (N_4042,N_3960,N_3955);
nor U4043 (N_4043,N_3970,N_3977);
xor U4044 (N_4044,N_3896,N_3905);
or U4045 (N_4045,N_3968,N_3928);
or U4046 (N_4046,N_3943,N_3923);
and U4047 (N_4047,N_3920,N_3974);
or U4048 (N_4048,N_3924,N_3933);
or U4049 (N_4049,N_3966,N_3925);
and U4050 (N_4050,N_3945,N_3914);
nand U4051 (N_4051,N_3952,N_3932);
xor U4052 (N_4052,N_3934,N_3980);
nor U4053 (N_4053,N_3998,N_3956);
nor U4054 (N_4054,N_3904,N_3926);
and U4055 (N_4055,N_3997,N_3910);
or U4056 (N_4056,N_3942,N_3999);
xor U4057 (N_4057,N_3922,N_3979);
xnor U4058 (N_4058,N_3987,N_3884);
nand U4059 (N_4059,N_3973,N_3899);
nand U4060 (N_4060,N_3894,N_3879);
and U4061 (N_4061,N_3931,N_3963);
nand U4062 (N_4062,N_3886,N_3901);
nand U4063 (N_4063,N_3940,N_3962);
nand U4064 (N_4064,N_3898,N_3925);
xnor U4065 (N_4065,N_3971,N_3892);
nor U4066 (N_4066,N_3918,N_3915);
and U4067 (N_4067,N_3958,N_3930);
and U4068 (N_4068,N_3991,N_3912);
and U4069 (N_4069,N_3879,N_3889);
nor U4070 (N_4070,N_3934,N_3979);
and U4071 (N_4071,N_3892,N_3958);
xnor U4072 (N_4072,N_3994,N_3921);
or U4073 (N_4073,N_3927,N_3954);
xor U4074 (N_4074,N_3915,N_3930);
nor U4075 (N_4075,N_3983,N_3964);
nor U4076 (N_4076,N_3919,N_3985);
xnor U4077 (N_4077,N_3901,N_3953);
nor U4078 (N_4078,N_3880,N_3939);
xor U4079 (N_4079,N_3911,N_3985);
and U4080 (N_4080,N_3987,N_3891);
or U4081 (N_4081,N_3952,N_3878);
nand U4082 (N_4082,N_3972,N_3927);
nand U4083 (N_4083,N_3981,N_3951);
nor U4084 (N_4084,N_3907,N_3992);
or U4085 (N_4085,N_3928,N_3919);
or U4086 (N_4086,N_3908,N_3877);
and U4087 (N_4087,N_3878,N_3977);
nand U4088 (N_4088,N_3947,N_3953);
or U4089 (N_4089,N_3885,N_3942);
and U4090 (N_4090,N_3961,N_3962);
xor U4091 (N_4091,N_3927,N_3899);
and U4092 (N_4092,N_3889,N_3918);
xnor U4093 (N_4093,N_3881,N_3893);
nand U4094 (N_4094,N_3900,N_3881);
xnor U4095 (N_4095,N_3959,N_3918);
or U4096 (N_4096,N_3912,N_3913);
nand U4097 (N_4097,N_3891,N_3888);
nor U4098 (N_4098,N_3908,N_3978);
and U4099 (N_4099,N_3971,N_3885);
nor U4100 (N_4100,N_3889,N_3899);
and U4101 (N_4101,N_3915,N_3982);
and U4102 (N_4102,N_3951,N_3893);
nor U4103 (N_4103,N_3947,N_3900);
nor U4104 (N_4104,N_3968,N_3939);
nor U4105 (N_4105,N_3967,N_3882);
nor U4106 (N_4106,N_3917,N_3925);
or U4107 (N_4107,N_3897,N_3983);
nor U4108 (N_4108,N_3963,N_3913);
and U4109 (N_4109,N_3918,N_3974);
nand U4110 (N_4110,N_3911,N_3899);
or U4111 (N_4111,N_3984,N_3998);
nor U4112 (N_4112,N_3896,N_3909);
or U4113 (N_4113,N_3949,N_3918);
or U4114 (N_4114,N_3965,N_3922);
and U4115 (N_4115,N_3997,N_3912);
and U4116 (N_4116,N_3982,N_3986);
or U4117 (N_4117,N_3966,N_3922);
nor U4118 (N_4118,N_3928,N_3946);
nor U4119 (N_4119,N_3968,N_3993);
nand U4120 (N_4120,N_3920,N_3972);
nor U4121 (N_4121,N_3956,N_3911);
and U4122 (N_4122,N_3962,N_3986);
nor U4123 (N_4123,N_3936,N_3931);
or U4124 (N_4124,N_3914,N_3996);
nand U4125 (N_4125,N_4113,N_4009);
xor U4126 (N_4126,N_4093,N_4072);
nand U4127 (N_4127,N_4084,N_4092);
nor U4128 (N_4128,N_4078,N_4089);
nand U4129 (N_4129,N_4006,N_4051);
nand U4130 (N_4130,N_4081,N_4109);
nand U4131 (N_4131,N_4067,N_4003);
and U4132 (N_4132,N_4087,N_4117);
and U4133 (N_4133,N_4119,N_4040);
or U4134 (N_4134,N_4052,N_4121);
xor U4135 (N_4135,N_4039,N_4035);
and U4136 (N_4136,N_4090,N_4049);
nand U4137 (N_4137,N_4055,N_4008);
nor U4138 (N_4138,N_4069,N_4043);
xor U4139 (N_4139,N_4059,N_4034);
nor U4140 (N_4140,N_4115,N_4036);
nor U4141 (N_4141,N_4100,N_4062);
nor U4142 (N_4142,N_4022,N_4077);
nand U4143 (N_4143,N_4083,N_4076);
or U4144 (N_4144,N_4038,N_4098);
nand U4145 (N_4145,N_4031,N_4068);
nand U4146 (N_4146,N_4026,N_4120);
or U4147 (N_4147,N_4048,N_4088);
and U4148 (N_4148,N_4001,N_4046);
xor U4149 (N_4149,N_4041,N_4095);
and U4150 (N_4150,N_4091,N_4020);
nand U4151 (N_4151,N_4082,N_4027);
nor U4152 (N_4152,N_4101,N_4075);
and U4153 (N_4153,N_4071,N_4070);
nor U4154 (N_4154,N_4086,N_4114);
nand U4155 (N_4155,N_4102,N_4042);
xor U4156 (N_4156,N_4057,N_4029);
xnor U4157 (N_4157,N_4002,N_4116);
and U4158 (N_4158,N_4018,N_4108);
or U4159 (N_4159,N_4104,N_4021);
or U4160 (N_4160,N_4105,N_4096);
nor U4161 (N_4161,N_4045,N_4053);
or U4162 (N_4162,N_4024,N_4015);
or U4163 (N_4163,N_4013,N_4094);
nand U4164 (N_4164,N_4047,N_4032);
nand U4165 (N_4165,N_4014,N_4060);
nand U4166 (N_4166,N_4061,N_4064);
xnor U4167 (N_4167,N_4066,N_4056);
xor U4168 (N_4168,N_4124,N_4044);
xnor U4169 (N_4169,N_4103,N_4111);
xnor U4170 (N_4170,N_4005,N_4050);
and U4171 (N_4171,N_4028,N_4054);
and U4172 (N_4172,N_4079,N_4118);
or U4173 (N_4173,N_4033,N_4000);
or U4174 (N_4174,N_4010,N_4030);
and U4175 (N_4175,N_4073,N_4017);
and U4176 (N_4176,N_4110,N_4007);
and U4177 (N_4177,N_4063,N_4011);
and U4178 (N_4178,N_4037,N_4085);
xor U4179 (N_4179,N_4058,N_4107);
nand U4180 (N_4180,N_4065,N_4112);
nor U4181 (N_4181,N_4004,N_4097);
nand U4182 (N_4182,N_4016,N_4012);
nand U4183 (N_4183,N_4122,N_4123);
nand U4184 (N_4184,N_4080,N_4106);
or U4185 (N_4185,N_4023,N_4019);
nand U4186 (N_4186,N_4099,N_4025);
nor U4187 (N_4187,N_4074,N_4048);
xnor U4188 (N_4188,N_4012,N_4119);
nand U4189 (N_4189,N_4048,N_4079);
and U4190 (N_4190,N_4034,N_4046);
or U4191 (N_4191,N_4040,N_4124);
and U4192 (N_4192,N_4101,N_4034);
or U4193 (N_4193,N_4059,N_4063);
nand U4194 (N_4194,N_4061,N_4015);
nand U4195 (N_4195,N_4052,N_4117);
xnor U4196 (N_4196,N_4046,N_4068);
nand U4197 (N_4197,N_4078,N_4020);
or U4198 (N_4198,N_4114,N_4017);
or U4199 (N_4199,N_4115,N_4024);
nand U4200 (N_4200,N_4078,N_4091);
and U4201 (N_4201,N_4099,N_4052);
or U4202 (N_4202,N_4070,N_4023);
or U4203 (N_4203,N_4007,N_4050);
and U4204 (N_4204,N_4082,N_4006);
nor U4205 (N_4205,N_4105,N_4111);
or U4206 (N_4206,N_4070,N_4093);
xor U4207 (N_4207,N_4002,N_4122);
nor U4208 (N_4208,N_4048,N_4005);
nor U4209 (N_4209,N_4038,N_4119);
nor U4210 (N_4210,N_4090,N_4003);
or U4211 (N_4211,N_4053,N_4055);
xor U4212 (N_4212,N_4083,N_4012);
nand U4213 (N_4213,N_4054,N_4103);
nor U4214 (N_4214,N_4026,N_4001);
and U4215 (N_4215,N_4017,N_4029);
nor U4216 (N_4216,N_4072,N_4083);
or U4217 (N_4217,N_4061,N_4111);
nand U4218 (N_4218,N_4119,N_4113);
xor U4219 (N_4219,N_4034,N_4123);
xnor U4220 (N_4220,N_4007,N_4065);
nor U4221 (N_4221,N_4035,N_4036);
nor U4222 (N_4222,N_4105,N_4031);
nand U4223 (N_4223,N_4019,N_4030);
nor U4224 (N_4224,N_4088,N_4067);
or U4225 (N_4225,N_4106,N_4101);
nand U4226 (N_4226,N_4083,N_4051);
xor U4227 (N_4227,N_4110,N_4113);
xor U4228 (N_4228,N_4016,N_4053);
or U4229 (N_4229,N_4025,N_4065);
or U4230 (N_4230,N_4075,N_4072);
and U4231 (N_4231,N_4116,N_4012);
nand U4232 (N_4232,N_4017,N_4097);
and U4233 (N_4233,N_4090,N_4019);
and U4234 (N_4234,N_4037,N_4101);
and U4235 (N_4235,N_4046,N_4119);
nand U4236 (N_4236,N_4080,N_4005);
nand U4237 (N_4237,N_4045,N_4088);
nor U4238 (N_4238,N_4016,N_4119);
or U4239 (N_4239,N_4029,N_4085);
nor U4240 (N_4240,N_4076,N_4074);
and U4241 (N_4241,N_4123,N_4020);
xnor U4242 (N_4242,N_4103,N_4116);
or U4243 (N_4243,N_4008,N_4051);
nor U4244 (N_4244,N_4026,N_4095);
nor U4245 (N_4245,N_4030,N_4091);
nor U4246 (N_4246,N_4110,N_4005);
nor U4247 (N_4247,N_4089,N_4103);
and U4248 (N_4248,N_4024,N_4091);
or U4249 (N_4249,N_4044,N_4108);
nor U4250 (N_4250,N_4170,N_4208);
nand U4251 (N_4251,N_4146,N_4211);
or U4252 (N_4252,N_4189,N_4244);
and U4253 (N_4253,N_4157,N_4241);
xor U4254 (N_4254,N_4190,N_4182);
nand U4255 (N_4255,N_4137,N_4153);
or U4256 (N_4256,N_4239,N_4169);
or U4257 (N_4257,N_4200,N_4249);
xnor U4258 (N_4258,N_4145,N_4181);
and U4259 (N_4259,N_4159,N_4209);
xnor U4260 (N_4260,N_4140,N_4150);
xnor U4261 (N_4261,N_4219,N_4185);
xor U4262 (N_4262,N_4168,N_4127);
nand U4263 (N_4263,N_4151,N_4186);
nand U4264 (N_4264,N_4248,N_4213);
nand U4265 (N_4265,N_4128,N_4135);
xor U4266 (N_4266,N_4187,N_4160);
nor U4267 (N_4267,N_4217,N_4230);
or U4268 (N_4268,N_4223,N_4233);
or U4269 (N_4269,N_4156,N_4215);
xor U4270 (N_4270,N_4167,N_4221);
nor U4271 (N_4271,N_4192,N_4161);
xor U4272 (N_4272,N_4232,N_4173);
nand U4273 (N_4273,N_4228,N_4227);
and U4274 (N_4274,N_4149,N_4216);
nand U4275 (N_4275,N_4155,N_4143);
and U4276 (N_4276,N_4238,N_4158);
and U4277 (N_4277,N_4152,N_4197);
nand U4278 (N_4278,N_4133,N_4172);
xnor U4279 (N_4279,N_4247,N_4130);
and U4280 (N_4280,N_4226,N_4125);
and U4281 (N_4281,N_4203,N_4236);
or U4282 (N_4282,N_4163,N_4184);
nand U4283 (N_4283,N_4176,N_4148);
and U4284 (N_4284,N_4202,N_4162);
and U4285 (N_4285,N_4191,N_4242);
nand U4286 (N_4286,N_4246,N_4165);
nor U4287 (N_4287,N_4234,N_4243);
or U4288 (N_4288,N_4204,N_4164);
nand U4289 (N_4289,N_4179,N_4206);
nand U4290 (N_4290,N_4240,N_4205);
nor U4291 (N_4291,N_4225,N_4171);
or U4292 (N_4292,N_4144,N_4195);
xnor U4293 (N_4293,N_4207,N_4174);
nor U4294 (N_4294,N_4147,N_4141);
and U4295 (N_4295,N_4235,N_4212);
nand U4296 (N_4296,N_4198,N_4196);
or U4297 (N_4297,N_4142,N_4199);
or U4298 (N_4298,N_4139,N_4166);
and U4299 (N_4299,N_4188,N_4220);
nor U4300 (N_4300,N_4193,N_4194);
xor U4301 (N_4301,N_4201,N_4136);
xor U4302 (N_4302,N_4138,N_4132);
nand U4303 (N_4303,N_4218,N_4222);
nor U4304 (N_4304,N_4177,N_4134);
nand U4305 (N_4305,N_4237,N_4175);
xor U4306 (N_4306,N_4224,N_4154);
nand U4307 (N_4307,N_4231,N_4229);
and U4308 (N_4308,N_4126,N_4245);
or U4309 (N_4309,N_4180,N_4178);
or U4310 (N_4310,N_4214,N_4210);
and U4311 (N_4311,N_4183,N_4131);
and U4312 (N_4312,N_4129,N_4167);
or U4313 (N_4313,N_4221,N_4232);
nor U4314 (N_4314,N_4165,N_4240);
or U4315 (N_4315,N_4190,N_4212);
and U4316 (N_4316,N_4166,N_4180);
xor U4317 (N_4317,N_4231,N_4140);
or U4318 (N_4318,N_4142,N_4145);
or U4319 (N_4319,N_4214,N_4221);
nand U4320 (N_4320,N_4126,N_4224);
or U4321 (N_4321,N_4184,N_4221);
nor U4322 (N_4322,N_4241,N_4221);
and U4323 (N_4323,N_4169,N_4194);
nor U4324 (N_4324,N_4220,N_4128);
or U4325 (N_4325,N_4162,N_4188);
nand U4326 (N_4326,N_4184,N_4205);
and U4327 (N_4327,N_4180,N_4153);
and U4328 (N_4328,N_4196,N_4241);
and U4329 (N_4329,N_4247,N_4166);
and U4330 (N_4330,N_4236,N_4132);
and U4331 (N_4331,N_4237,N_4131);
nor U4332 (N_4332,N_4187,N_4130);
nor U4333 (N_4333,N_4202,N_4149);
and U4334 (N_4334,N_4170,N_4154);
nor U4335 (N_4335,N_4249,N_4134);
or U4336 (N_4336,N_4144,N_4201);
or U4337 (N_4337,N_4215,N_4177);
and U4338 (N_4338,N_4130,N_4219);
xor U4339 (N_4339,N_4219,N_4142);
and U4340 (N_4340,N_4209,N_4219);
xnor U4341 (N_4341,N_4196,N_4134);
or U4342 (N_4342,N_4244,N_4161);
nand U4343 (N_4343,N_4193,N_4200);
xor U4344 (N_4344,N_4129,N_4229);
nor U4345 (N_4345,N_4147,N_4188);
nor U4346 (N_4346,N_4143,N_4216);
and U4347 (N_4347,N_4208,N_4135);
nor U4348 (N_4348,N_4244,N_4228);
nor U4349 (N_4349,N_4219,N_4180);
nand U4350 (N_4350,N_4142,N_4205);
and U4351 (N_4351,N_4207,N_4222);
nand U4352 (N_4352,N_4171,N_4224);
or U4353 (N_4353,N_4165,N_4229);
and U4354 (N_4354,N_4232,N_4214);
and U4355 (N_4355,N_4193,N_4212);
or U4356 (N_4356,N_4204,N_4160);
nor U4357 (N_4357,N_4126,N_4169);
or U4358 (N_4358,N_4183,N_4155);
nor U4359 (N_4359,N_4225,N_4194);
or U4360 (N_4360,N_4157,N_4133);
xnor U4361 (N_4361,N_4239,N_4219);
and U4362 (N_4362,N_4156,N_4209);
nor U4363 (N_4363,N_4125,N_4196);
and U4364 (N_4364,N_4212,N_4215);
xor U4365 (N_4365,N_4177,N_4198);
nor U4366 (N_4366,N_4197,N_4127);
xor U4367 (N_4367,N_4245,N_4200);
nand U4368 (N_4368,N_4133,N_4246);
nand U4369 (N_4369,N_4212,N_4228);
nand U4370 (N_4370,N_4128,N_4230);
nand U4371 (N_4371,N_4179,N_4232);
xnor U4372 (N_4372,N_4165,N_4178);
and U4373 (N_4373,N_4202,N_4175);
nand U4374 (N_4374,N_4230,N_4238);
xor U4375 (N_4375,N_4259,N_4362);
xnor U4376 (N_4376,N_4360,N_4366);
xor U4377 (N_4377,N_4276,N_4361);
nor U4378 (N_4378,N_4352,N_4255);
nor U4379 (N_4379,N_4261,N_4283);
or U4380 (N_4380,N_4309,N_4299);
or U4381 (N_4381,N_4293,N_4373);
nor U4382 (N_4382,N_4305,N_4271);
and U4383 (N_4383,N_4348,N_4265);
and U4384 (N_4384,N_4278,N_4272);
xor U4385 (N_4385,N_4301,N_4339);
or U4386 (N_4386,N_4357,N_4304);
or U4387 (N_4387,N_4329,N_4338);
or U4388 (N_4388,N_4317,N_4279);
or U4389 (N_4389,N_4280,N_4258);
and U4390 (N_4390,N_4253,N_4297);
or U4391 (N_4391,N_4295,N_4359);
and U4392 (N_4392,N_4343,N_4328);
or U4393 (N_4393,N_4346,N_4356);
or U4394 (N_4394,N_4353,N_4256);
or U4395 (N_4395,N_4333,N_4316);
or U4396 (N_4396,N_4302,N_4288);
and U4397 (N_4397,N_4370,N_4312);
xor U4398 (N_4398,N_4367,N_4296);
and U4399 (N_4399,N_4264,N_4341);
xor U4400 (N_4400,N_4326,N_4314);
xor U4401 (N_4401,N_4277,N_4351);
nor U4402 (N_4402,N_4350,N_4325);
or U4403 (N_4403,N_4298,N_4267);
nor U4404 (N_4404,N_4303,N_4273);
and U4405 (N_4405,N_4251,N_4374);
or U4406 (N_4406,N_4363,N_4372);
nor U4407 (N_4407,N_4365,N_4263);
nor U4408 (N_4408,N_4252,N_4324);
nor U4409 (N_4409,N_4250,N_4355);
nor U4410 (N_4410,N_4331,N_4307);
xnor U4411 (N_4411,N_4270,N_4371);
xor U4412 (N_4412,N_4281,N_4347);
xor U4413 (N_4413,N_4257,N_4260);
xnor U4414 (N_4414,N_4368,N_4315);
xnor U4415 (N_4415,N_4340,N_4349);
and U4416 (N_4416,N_4292,N_4318);
nand U4417 (N_4417,N_4354,N_4335);
nor U4418 (N_4418,N_4306,N_4310);
nor U4419 (N_4419,N_4269,N_4311);
or U4420 (N_4420,N_4290,N_4358);
or U4421 (N_4421,N_4274,N_4289);
xor U4422 (N_4422,N_4284,N_4285);
xor U4423 (N_4423,N_4262,N_4300);
xor U4424 (N_4424,N_4342,N_4327);
nor U4425 (N_4425,N_4330,N_4323);
and U4426 (N_4426,N_4322,N_4254);
or U4427 (N_4427,N_4291,N_4364);
xnor U4428 (N_4428,N_4334,N_4294);
and U4429 (N_4429,N_4319,N_4308);
nor U4430 (N_4430,N_4282,N_4268);
nand U4431 (N_4431,N_4313,N_4287);
and U4432 (N_4432,N_4336,N_4345);
nor U4433 (N_4433,N_4344,N_4275);
xor U4434 (N_4434,N_4320,N_4286);
xnor U4435 (N_4435,N_4266,N_4332);
or U4436 (N_4436,N_4321,N_4369);
nand U4437 (N_4437,N_4337,N_4290);
nand U4438 (N_4438,N_4322,N_4259);
xor U4439 (N_4439,N_4360,N_4299);
nand U4440 (N_4440,N_4303,N_4260);
or U4441 (N_4441,N_4282,N_4311);
or U4442 (N_4442,N_4259,N_4328);
nand U4443 (N_4443,N_4352,N_4251);
nand U4444 (N_4444,N_4313,N_4325);
nor U4445 (N_4445,N_4360,N_4307);
and U4446 (N_4446,N_4267,N_4349);
nor U4447 (N_4447,N_4303,N_4276);
and U4448 (N_4448,N_4348,N_4367);
nor U4449 (N_4449,N_4313,N_4338);
and U4450 (N_4450,N_4337,N_4288);
and U4451 (N_4451,N_4343,N_4299);
nor U4452 (N_4452,N_4287,N_4253);
nor U4453 (N_4453,N_4369,N_4255);
nor U4454 (N_4454,N_4316,N_4353);
nand U4455 (N_4455,N_4262,N_4362);
nand U4456 (N_4456,N_4265,N_4299);
nand U4457 (N_4457,N_4304,N_4332);
and U4458 (N_4458,N_4261,N_4344);
nand U4459 (N_4459,N_4286,N_4268);
or U4460 (N_4460,N_4311,N_4325);
nor U4461 (N_4461,N_4288,N_4255);
and U4462 (N_4462,N_4336,N_4309);
nor U4463 (N_4463,N_4318,N_4304);
or U4464 (N_4464,N_4294,N_4315);
nand U4465 (N_4465,N_4274,N_4352);
nand U4466 (N_4466,N_4340,N_4364);
nand U4467 (N_4467,N_4346,N_4270);
or U4468 (N_4468,N_4303,N_4278);
xor U4469 (N_4469,N_4321,N_4324);
and U4470 (N_4470,N_4341,N_4360);
xnor U4471 (N_4471,N_4306,N_4304);
nor U4472 (N_4472,N_4285,N_4352);
xor U4473 (N_4473,N_4323,N_4332);
nor U4474 (N_4474,N_4294,N_4359);
nor U4475 (N_4475,N_4258,N_4302);
and U4476 (N_4476,N_4334,N_4368);
xor U4477 (N_4477,N_4295,N_4371);
xnor U4478 (N_4478,N_4363,N_4250);
nand U4479 (N_4479,N_4355,N_4273);
and U4480 (N_4480,N_4365,N_4255);
xnor U4481 (N_4481,N_4308,N_4337);
or U4482 (N_4482,N_4252,N_4315);
and U4483 (N_4483,N_4347,N_4302);
xor U4484 (N_4484,N_4259,N_4344);
xor U4485 (N_4485,N_4328,N_4348);
nand U4486 (N_4486,N_4349,N_4361);
and U4487 (N_4487,N_4374,N_4255);
nor U4488 (N_4488,N_4356,N_4299);
nor U4489 (N_4489,N_4262,N_4291);
nor U4490 (N_4490,N_4353,N_4321);
or U4491 (N_4491,N_4328,N_4287);
or U4492 (N_4492,N_4360,N_4294);
and U4493 (N_4493,N_4341,N_4261);
nand U4494 (N_4494,N_4256,N_4311);
or U4495 (N_4495,N_4320,N_4361);
nand U4496 (N_4496,N_4265,N_4333);
or U4497 (N_4497,N_4269,N_4369);
or U4498 (N_4498,N_4319,N_4345);
or U4499 (N_4499,N_4311,N_4338);
xnor U4500 (N_4500,N_4497,N_4404);
xnor U4501 (N_4501,N_4384,N_4402);
and U4502 (N_4502,N_4405,N_4407);
nor U4503 (N_4503,N_4399,N_4483);
or U4504 (N_4504,N_4416,N_4456);
and U4505 (N_4505,N_4458,N_4478);
nor U4506 (N_4506,N_4390,N_4495);
xor U4507 (N_4507,N_4398,N_4425);
and U4508 (N_4508,N_4385,N_4392);
or U4509 (N_4509,N_4417,N_4418);
xor U4510 (N_4510,N_4415,N_4480);
nor U4511 (N_4511,N_4432,N_4381);
and U4512 (N_4512,N_4394,N_4410);
and U4513 (N_4513,N_4378,N_4421);
xnor U4514 (N_4514,N_4489,N_4482);
or U4515 (N_4515,N_4444,N_4414);
nor U4516 (N_4516,N_4455,N_4470);
nand U4517 (N_4517,N_4427,N_4488);
nand U4518 (N_4518,N_4436,N_4428);
and U4519 (N_4519,N_4412,N_4377);
nand U4520 (N_4520,N_4469,N_4491);
nand U4521 (N_4521,N_4431,N_4481);
nor U4522 (N_4522,N_4383,N_4492);
and U4523 (N_4523,N_4499,N_4494);
or U4524 (N_4524,N_4433,N_4490);
nand U4525 (N_4525,N_4382,N_4453);
or U4526 (N_4526,N_4380,N_4464);
nand U4527 (N_4527,N_4387,N_4375);
or U4528 (N_4528,N_4391,N_4400);
or U4529 (N_4529,N_4413,N_4420);
xor U4530 (N_4530,N_4439,N_4376);
and U4531 (N_4531,N_4449,N_4406);
or U4532 (N_4532,N_4445,N_4487);
and U4533 (N_4533,N_4459,N_4477);
xor U4534 (N_4534,N_4467,N_4498);
xor U4535 (N_4535,N_4461,N_4452);
and U4536 (N_4536,N_4484,N_4437);
and U4537 (N_4537,N_4396,N_4448);
nor U4538 (N_4538,N_4451,N_4457);
or U4539 (N_4539,N_4438,N_4468);
nor U4540 (N_4540,N_4430,N_4403);
or U4541 (N_4541,N_4386,N_4493);
nor U4542 (N_4542,N_4409,N_4397);
or U4543 (N_4543,N_4471,N_4443);
nand U4544 (N_4544,N_4446,N_4434);
xnor U4545 (N_4545,N_4447,N_4476);
or U4546 (N_4546,N_4411,N_4423);
or U4547 (N_4547,N_4440,N_4473);
xor U4548 (N_4548,N_4486,N_4463);
nor U4549 (N_4549,N_4408,N_4393);
or U4550 (N_4550,N_4479,N_4474);
or U4551 (N_4551,N_4462,N_4466);
xnor U4552 (N_4552,N_4496,N_4379);
xor U4553 (N_4553,N_4388,N_4419);
or U4554 (N_4554,N_4422,N_4435);
xor U4555 (N_4555,N_4429,N_4426);
nand U4556 (N_4556,N_4424,N_4465);
and U4557 (N_4557,N_4450,N_4485);
and U4558 (N_4558,N_4442,N_4460);
nand U4559 (N_4559,N_4441,N_4401);
nor U4560 (N_4560,N_4472,N_4389);
xor U4561 (N_4561,N_4454,N_4475);
nand U4562 (N_4562,N_4395,N_4498);
and U4563 (N_4563,N_4380,N_4499);
and U4564 (N_4564,N_4404,N_4499);
or U4565 (N_4565,N_4443,N_4387);
or U4566 (N_4566,N_4469,N_4436);
xnor U4567 (N_4567,N_4392,N_4400);
nor U4568 (N_4568,N_4449,N_4404);
nand U4569 (N_4569,N_4477,N_4481);
and U4570 (N_4570,N_4406,N_4482);
and U4571 (N_4571,N_4448,N_4390);
and U4572 (N_4572,N_4394,N_4404);
xnor U4573 (N_4573,N_4449,N_4492);
nand U4574 (N_4574,N_4376,N_4428);
nand U4575 (N_4575,N_4436,N_4433);
nor U4576 (N_4576,N_4484,N_4470);
nand U4577 (N_4577,N_4377,N_4481);
nor U4578 (N_4578,N_4462,N_4403);
xnor U4579 (N_4579,N_4464,N_4463);
xor U4580 (N_4580,N_4469,N_4488);
nand U4581 (N_4581,N_4441,N_4380);
nor U4582 (N_4582,N_4456,N_4488);
nor U4583 (N_4583,N_4492,N_4463);
nor U4584 (N_4584,N_4397,N_4460);
nand U4585 (N_4585,N_4394,N_4478);
nand U4586 (N_4586,N_4429,N_4379);
nand U4587 (N_4587,N_4437,N_4398);
or U4588 (N_4588,N_4481,N_4443);
and U4589 (N_4589,N_4408,N_4418);
and U4590 (N_4590,N_4378,N_4483);
xor U4591 (N_4591,N_4451,N_4390);
nand U4592 (N_4592,N_4406,N_4458);
xnor U4593 (N_4593,N_4450,N_4429);
nand U4594 (N_4594,N_4411,N_4393);
nand U4595 (N_4595,N_4401,N_4419);
nand U4596 (N_4596,N_4470,N_4439);
xnor U4597 (N_4597,N_4416,N_4428);
nor U4598 (N_4598,N_4425,N_4411);
nor U4599 (N_4599,N_4422,N_4479);
nor U4600 (N_4600,N_4482,N_4474);
xor U4601 (N_4601,N_4429,N_4439);
and U4602 (N_4602,N_4412,N_4493);
and U4603 (N_4603,N_4447,N_4481);
nand U4604 (N_4604,N_4440,N_4429);
xnor U4605 (N_4605,N_4377,N_4415);
nand U4606 (N_4606,N_4496,N_4498);
nand U4607 (N_4607,N_4468,N_4399);
xnor U4608 (N_4608,N_4451,N_4463);
or U4609 (N_4609,N_4476,N_4409);
xnor U4610 (N_4610,N_4493,N_4487);
xor U4611 (N_4611,N_4389,N_4400);
and U4612 (N_4612,N_4424,N_4487);
xnor U4613 (N_4613,N_4392,N_4425);
or U4614 (N_4614,N_4404,N_4490);
and U4615 (N_4615,N_4429,N_4400);
nand U4616 (N_4616,N_4429,N_4468);
and U4617 (N_4617,N_4460,N_4492);
nor U4618 (N_4618,N_4408,N_4422);
xnor U4619 (N_4619,N_4382,N_4499);
nand U4620 (N_4620,N_4448,N_4429);
nor U4621 (N_4621,N_4457,N_4484);
and U4622 (N_4622,N_4491,N_4382);
nor U4623 (N_4623,N_4407,N_4396);
or U4624 (N_4624,N_4392,N_4475);
nor U4625 (N_4625,N_4531,N_4613);
or U4626 (N_4626,N_4500,N_4513);
or U4627 (N_4627,N_4509,N_4576);
nand U4628 (N_4628,N_4602,N_4599);
xnor U4629 (N_4629,N_4591,N_4600);
nand U4630 (N_4630,N_4561,N_4567);
xnor U4631 (N_4631,N_4551,N_4589);
nor U4632 (N_4632,N_4533,N_4565);
or U4633 (N_4633,N_4583,N_4549);
nand U4634 (N_4634,N_4596,N_4536);
xor U4635 (N_4635,N_4504,N_4547);
xor U4636 (N_4636,N_4528,N_4605);
or U4637 (N_4637,N_4594,N_4524);
nand U4638 (N_4638,N_4570,N_4568);
nand U4639 (N_4639,N_4537,N_4609);
nand U4640 (N_4640,N_4523,N_4514);
xnor U4641 (N_4641,N_4520,N_4557);
nor U4642 (N_4642,N_4562,N_4580);
xor U4643 (N_4643,N_4542,N_4622);
or U4644 (N_4644,N_4588,N_4606);
nand U4645 (N_4645,N_4538,N_4621);
nor U4646 (N_4646,N_4521,N_4539);
nand U4647 (N_4647,N_4604,N_4593);
xor U4648 (N_4648,N_4552,N_4595);
nor U4649 (N_4649,N_4526,N_4546);
nand U4650 (N_4650,N_4584,N_4607);
or U4651 (N_4651,N_4555,N_4571);
and U4652 (N_4652,N_4519,N_4507);
and U4653 (N_4653,N_4534,N_4573);
or U4654 (N_4654,N_4510,N_4578);
nor U4655 (N_4655,N_4582,N_4543);
nand U4656 (N_4656,N_4619,N_4517);
and U4657 (N_4657,N_4585,N_4529);
nor U4658 (N_4658,N_4512,N_4564);
and U4659 (N_4659,N_4615,N_4590);
xnor U4660 (N_4660,N_4511,N_4566);
xor U4661 (N_4661,N_4612,N_4581);
nand U4662 (N_4662,N_4614,N_4532);
and U4663 (N_4663,N_4522,N_4544);
or U4664 (N_4664,N_4554,N_4563);
and U4665 (N_4665,N_4506,N_4587);
nand U4666 (N_4666,N_4508,N_4597);
and U4667 (N_4667,N_4618,N_4530);
xor U4668 (N_4668,N_4586,N_4556);
and U4669 (N_4669,N_4515,N_4577);
nand U4670 (N_4670,N_4569,N_4550);
nor U4671 (N_4671,N_4502,N_4601);
xnor U4672 (N_4672,N_4623,N_4501);
or U4673 (N_4673,N_4592,N_4610);
nor U4674 (N_4674,N_4535,N_4575);
xnor U4675 (N_4675,N_4541,N_4598);
and U4676 (N_4676,N_4553,N_4558);
nor U4677 (N_4677,N_4624,N_4548);
nand U4678 (N_4678,N_4617,N_4559);
xnor U4679 (N_4679,N_4574,N_4616);
and U4680 (N_4680,N_4505,N_4603);
nand U4681 (N_4681,N_4516,N_4560);
or U4682 (N_4682,N_4525,N_4545);
nand U4683 (N_4683,N_4540,N_4527);
nor U4684 (N_4684,N_4518,N_4620);
and U4685 (N_4685,N_4611,N_4572);
or U4686 (N_4686,N_4608,N_4579);
or U4687 (N_4687,N_4503,N_4542);
nor U4688 (N_4688,N_4526,N_4520);
nand U4689 (N_4689,N_4501,N_4512);
nand U4690 (N_4690,N_4593,N_4529);
or U4691 (N_4691,N_4524,N_4564);
nand U4692 (N_4692,N_4589,N_4582);
nor U4693 (N_4693,N_4601,N_4572);
and U4694 (N_4694,N_4548,N_4533);
or U4695 (N_4695,N_4529,N_4569);
xor U4696 (N_4696,N_4617,N_4543);
nor U4697 (N_4697,N_4624,N_4527);
or U4698 (N_4698,N_4506,N_4519);
nor U4699 (N_4699,N_4531,N_4546);
xor U4700 (N_4700,N_4607,N_4556);
xnor U4701 (N_4701,N_4528,N_4505);
nand U4702 (N_4702,N_4547,N_4526);
xnor U4703 (N_4703,N_4516,N_4535);
nor U4704 (N_4704,N_4507,N_4621);
xnor U4705 (N_4705,N_4607,N_4567);
xor U4706 (N_4706,N_4549,N_4527);
or U4707 (N_4707,N_4523,N_4623);
and U4708 (N_4708,N_4607,N_4612);
xnor U4709 (N_4709,N_4571,N_4540);
or U4710 (N_4710,N_4576,N_4527);
nor U4711 (N_4711,N_4525,N_4553);
nand U4712 (N_4712,N_4586,N_4618);
nor U4713 (N_4713,N_4504,N_4548);
nand U4714 (N_4714,N_4618,N_4595);
nor U4715 (N_4715,N_4550,N_4575);
nand U4716 (N_4716,N_4534,N_4516);
nor U4717 (N_4717,N_4503,N_4585);
nor U4718 (N_4718,N_4552,N_4622);
and U4719 (N_4719,N_4559,N_4532);
or U4720 (N_4720,N_4542,N_4605);
and U4721 (N_4721,N_4619,N_4576);
and U4722 (N_4722,N_4526,N_4540);
and U4723 (N_4723,N_4583,N_4526);
nand U4724 (N_4724,N_4604,N_4520);
nand U4725 (N_4725,N_4512,N_4537);
or U4726 (N_4726,N_4596,N_4543);
nand U4727 (N_4727,N_4554,N_4558);
or U4728 (N_4728,N_4525,N_4527);
nand U4729 (N_4729,N_4566,N_4545);
nor U4730 (N_4730,N_4594,N_4555);
and U4731 (N_4731,N_4594,N_4542);
or U4732 (N_4732,N_4614,N_4546);
xnor U4733 (N_4733,N_4566,N_4577);
nand U4734 (N_4734,N_4568,N_4574);
or U4735 (N_4735,N_4558,N_4613);
or U4736 (N_4736,N_4575,N_4543);
and U4737 (N_4737,N_4610,N_4601);
nor U4738 (N_4738,N_4572,N_4596);
and U4739 (N_4739,N_4541,N_4560);
and U4740 (N_4740,N_4574,N_4520);
nand U4741 (N_4741,N_4570,N_4530);
xor U4742 (N_4742,N_4594,N_4553);
nand U4743 (N_4743,N_4616,N_4514);
or U4744 (N_4744,N_4501,N_4601);
or U4745 (N_4745,N_4609,N_4519);
and U4746 (N_4746,N_4529,N_4549);
nand U4747 (N_4747,N_4605,N_4536);
nor U4748 (N_4748,N_4594,N_4519);
nor U4749 (N_4749,N_4556,N_4618);
and U4750 (N_4750,N_4698,N_4661);
and U4751 (N_4751,N_4743,N_4634);
xnor U4752 (N_4752,N_4647,N_4709);
nand U4753 (N_4753,N_4729,N_4684);
xor U4754 (N_4754,N_4732,N_4719);
and U4755 (N_4755,N_4688,N_4740);
nand U4756 (N_4756,N_4701,N_4715);
nand U4757 (N_4757,N_4640,N_4703);
or U4758 (N_4758,N_4636,N_4731);
and U4759 (N_4759,N_4638,N_4723);
or U4760 (N_4760,N_4694,N_4635);
xnor U4761 (N_4761,N_4749,N_4669);
nand U4762 (N_4762,N_4683,N_4662);
nor U4763 (N_4763,N_4744,N_4639);
and U4764 (N_4764,N_4716,N_4642);
nor U4765 (N_4765,N_4734,N_4670);
or U4766 (N_4766,N_4663,N_4682);
and U4767 (N_4767,N_4727,N_4726);
nand U4768 (N_4768,N_4676,N_4686);
and U4769 (N_4769,N_4697,N_4700);
and U4770 (N_4770,N_4745,N_4718);
nand U4771 (N_4771,N_4707,N_4728);
or U4772 (N_4772,N_4691,N_4742);
nor U4773 (N_4773,N_4748,N_4651);
and U4774 (N_4774,N_4650,N_4643);
nand U4775 (N_4775,N_4648,N_4702);
nor U4776 (N_4776,N_4660,N_4721);
nor U4777 (N_4777,N_4704,N_4730);
nand U4778 (N_4778,N_4738,N_4664);
xnor U4779 (N_4779,N_4652,N_4722);
or U4780 (N_4780,N_4712,N_4708);
or U4781 (N_4781,N_4667,N_4720);
xor U4782 (N_4782,N_4678,N_4711);
and U4783 (N_4783,N_4673,N_4675);
xnor U4784 (N_4784,N_4689,N_4654);
xnor U4785 (N_4785,N_4666,N_4695);
xnor U4786 (N_4786,N_4674,N_4677);
nor U4787 (N_4787,N_4630,N_4627);
and U4788 (N_4788,N_4625,N_4696);
nor U4789 (N_4789,N_4665,N_4736);
nor U4790 (N_4790,N_4645,N_4706);
xnor U4791 (N_4791,N_4649,N_4739);
xnor U4792 (N_4792,N_4687,N_4655);
xnor U4793 (N_4793,N_4685,N_4657);
nand U4794 (N_4794,N_4637,N_4671);
and U4795 (N_4795,N_4746,N_4626);
and U4796 (N_4796,N_4633,N_4672);
nor U4797 (N_4797,N_4705,N_4733);
nor U4798 (N_4798,N_4741,N_4628);
and U4799 (N_4799,N_4659,N_4714);
or U4800 (N_4800,N_4641,N_4699);
nor U4801 (N_4801,N_4724,N_4692);
or U4802 (N_4802,N_4713,N_4679);
and U4803 (N_4803,N_4681,N_4680);
nand U4804 (N_4804,N_4725,N_4717);
xnor U4805 (N_4805,N_4735,N_4747);
nor U4806 (N_4806,N_4646,N_4693);
or U4807 (N_4807,N_4690,N_4629);
xor U4808 (N_4808,N_4656,N_4710);
nand U4809 (N_4809,N_4632,N_4668);
xnor U4810 (N_4810,N_4644,N_4737);
xnor U4811 (N_4811,N_4631,N_4653);
or U4812 (N_4812,N_4658,N_4739);
and U4813 (N_4813,N_4704,N_4673);
xor U4814 (N_4814,N_4710,N_4633);
nor U4815 (N_4815,N_4646,N_4716);
nand U4816 (N_4816,N_4727,N_4669);
nand U4817 (N_4817,N_4699,N_4626);
and U4818 (N_4818,N_4723,N_4631);
nand U4819 (N_4819,N_4685,N_4662);
nor U4820 (N_4820,N_4689,N_4644);
and U4821 (N_4821,N_4679,N_4746);
and U4822 (N_4822,N_4643,N_4678);
and U4823 (N_4823,N_4685,N_4709);
xnor U4824 (N_4824,N_4677,N_4668);
and U4825 (N_4825,N_4706,N_4656);
and U4826 (N_4826,N_4670,N_4689);
nand U4827 (N_4827,N_4678,N_4721);
nand U4828 (N_4828,N_4643,N_4743);
or U4829 (N_4829,N_4672,N_4696);
or U4830 (N_4830,N_4724,N_4709);
nor U4831 (N_4831,N_4706,N_4679);
xor U4832 (N_4832,N_4746,N_4692);
nand U4833 (N_4833,N_4723,N_4708);
nand U4834 (N_4834,N_4729,N_4746);
nor U4835 (N_4835,N_4712,N_4666);
and U4836 (N_4836,N_4747,N_4720);
nand U4837 (N_4837,N_4710,N_4744);
and U4838 (N_4838,N_4740,N_4735);
xnor U4839 (N_4839,N_4626,N_4734);
or U4840 (N_4840,N_4746,N_4633);
and U4841 (N_4841,N_4647,N_4731);
nor U4842 (N_4842,N_4695,N_4716);
nand U4843 (N_4843,N_4732,N_4666);
nor U4844 (N_4844,N_4734,N_4660);
nand U4845 (N_4845,N_4683,N_4695);
and U4846 (N_4846,N_4647,N_4698);
nor U4847 (N_4847,N_4634,N_4710);
nand U4848 (N_4848,N_4726,N_4695);
xnor U4849 (N_4849,N_4683,N_4637);
and U4850 (N_4850,N_4676,N_4725);
and U4851 (N_4851,N_4644,N_4640);
xnor U4852 (N_4852,N_4733,N_4726);
nor U4853 (N_4853,N_4730,N_4665);
nand U4854 (N_4854,N_4678,N_4645);
nor U4855 (N_4855,N_4625,N_4702);
nand U4856 (N_4856,N_4632,N_4740);
nand U4857 (N_4857,N_4657,N_4725);
xor U4858 (N_4858,N_4731,N_4653);
and U4859 (N_4859,N_4642,N_4675);
nor U4860 (N_4860,N_4705,N_4749);
nor U4861 (N_4861,N_4654,N_4646);
or U4862 (N_4862,N_4679,N_4701);
nor U4863 (N_4863,N_4738,N_4649);
nand U4864 (N_4864,N_4703,N_4744);
and U4865 (N_4865,N_4631,N_4646);
and U4866 (N_4866,N_4697,N_4662);
and U4867 (N_4867,N_4727,N_4687);
nor U4868 (N_4868,N_4661,N_4737);
xor U4869 (N_4869,N_4689,N_4720);
nand U4870 (N_4870,N_4691,N_4627);
or U4871 (N_4871,N_4701,N_4722);
nor U4872 (N_4872,N_4702,N_4693);
and U4873 (N_4873,N_4695,N_4703);
and U4874 (N_4874,N_4670,N_4680);
nand U4875 (N_4875,N_4813,N_4759);
nor U4876 (N_4876,N_4825,N_4820);
xnor U4877 (N_4877,N_4753,N_4804);
or U4878 (N_4878,N_4790,N_4866);
nand U4879 (N_4879,N_4830,N_4835);
nand U4880 (N_4880,N_4803,N_4750);
nor U4881 (N_4881,N_4786,N_4773);
nor U4882 (N_4882,N_4756,N_4807);
and U4883 (N_4883,N_4772,N_4839);
xor U4884 (N_4884,N_4853,N_4789);
xor U4885 (N_4885,N_4785,N_4868);
xor U4886 (N_4886,N_4826,N_4808);
or U4887 (N_4887,N_4817,N_4847);
nand U4888 (N_4888,N_4796,N_4770);
nor U4889 (N_4889,N_4794,N_4771);
nand U4890 (N_4890,N_4840,N_4872);
nand U4891 (N_4891,N_4752,N_4871);
nand U4892 (N_4892,N_4762,N_4812);
nor U4893 (N_4893,N_4834,N_4865);
and U4894 (N_4894,N_4819,N_4763);
or U4895 (N_4895,N_4761,N_4795);
nand U4896 (N_4896,N_4860,N_4767);
or U4897 (N_4897,N_4855,N_4791);
nand U4898 (N_4898,N_4846,N_4861);
xor U4899 (N_4899,N_4776,N_4798);
nor U4900 (N_4900,N_4870,N_4851);
or U4901 (N_4901,N_4842,N_4782);
xnor U4902 (N_4902,N_4751,N_4765);
nand U4903 (N_4903,N_4768,N_4754);
nand U4904 (N_4904,N_4780,N_4764);
and U4905 (N_4905,N_4774,N_4850);
and U4906 (N_4906,N_4836,N_4845);
xnor U4907 (N_4907,N_4769,N_4856);
and U4908 (N_4908,N_4869,N_4805);
or U4909 (N_4909,N_4787,N_4858);
nor U4910 (N_4910,N_4793,N_4854);
xnor U4911 (N_4911,N_4802,N_4755);
nand U4912 (N_4912,N_4779,N_4781);
xnor U4913 (N_4913,N_4783,N_4800);
or U4914 (N_4914,N_4824,N_4760);
xnor U4915 (N_4915,N_4823,N_4801);
nor U4916 (N_4916,N_4775,N_4837);
or U4917 (N_4917,N_4799,N_4867);
and U4918 (N_4918,N_4848,N_4832);
xor U4919 (N_4919,N_4797,N_4841);
and U4920 (N_4920,N_4833,N_4815);
nor U4921 (N_4921,N_4852,N_4873);
or U4922 (N_4922,N_4816,N_4821);
and U4923 (N_4923,N_4831,N_4844);
and U4924 (N_4924,N_4838,N_4864);
nand U4925 (N_4925,N_4857,N_4766);
nor U4926 (N_4926,N_4828,N_4862);
xnor U4927 (N_4927,N_4806,N_4822);
or U4928 (N_4928,N_4792,N_4811);
and U4929 (N_4929,N_4849,N_4843);
xnor U4930 (N_4930,N_4818,N_4809);
or U4931 (N_4931,N_4758,N_4810);
and U4932 (N_4932,N_4829,N_4827);
nand U4933 (N_4933,N_4784,N_4788);
or U4934 (N_4934,N_4778,N_4814);
xnor U4935 (N_4935,N_4777,N_4874);
or U4936 (N_4936,N_4859,N_4757);
nand U4937 (N_4937,N_4863,N_4755);
and U4938 (N_4938,N_4865,N_4824);
nand U4939 (N_4939,N_4774,N_4831);
xnor U4940 (N_4940,N_4811,N_4763);
xor U4941 (N_4941,N_4805,N_4816);
xnor U4942 (N_4942,N_4870,N_4854);
and U4943 (N_4943,N_4831,N_4843);
xnor U4944 (N_4944,N_4871,N_4837);
nor U4945 (N_4945,N_4794,N_4767);
xnor U4946 (N_4946,N_4776,N_4782);
xnor U4947 (N_4947,N_4821,N_4751);
and U4948 (N_4948,N_4766,N_4833);
xnor U4949 (N_4949,N_4765,N_4760);
or U4950 (N_4950,N_4758,N_4856);
nand U4951 (N_4951,N_4851,N_4854);
and U4952 (N_4952,N_4852,N_4811);
or U4953 (N_4953,N_4849,N_4850);
xor U4954 (N_4954,N_4760,N_4828);
and U4955 (N_4955,N_4761,N_4756);
xnor U4956 (N_4956,N_4779,N_4844);
nand U4957 (N_4957,N_4840,N_4808);
xor U4958 (N_4958,N_4837,N_4828);
nand U4959 (N_4959,N_4858,N_4867);
nor U4960 (N_4960,N_4762,N_4835);
nor U4961 (N_4961,N_4761,N_4835);
xor U4962 (N_4962,N_4862,N_4754);
nor U4963 (N_4963,N_4783,N_4865);
or U4964 (N_4964,N_4825,N_4853);
xor U4965 (N_4965,N_4799,N_4844);
xor U4966 (N_4966,N_4814,N_4859);
and U4967 (N_4967,N_4784,N_4792);
nand U4968 (N_4968,N_4804,N_4820);
or U4969 (N_4969,N_4832,N_4847);
and U4970 (N_4970,N_4823,N_4755);
xnor U4971 (N_4971,N_4809,N_4769);
nand U4972 (N_4972,N_4851,N_4791);
or U4973 (N_4973,N_4816,N_4848);
nand U4974 (N_4974,N_4862,N_4871);
and U4975 (N_4975,N_4837,N_4763);
xor U4976 (N_4976,N_4813,N_4795);
and U4977 (N_4977,N_4869,N_4757);
xnor U4978 (N_4978,N_4842,N_4816);
and U4979 (N_4979,N_4750,N_4843);
or U4980 (N_4980,N_4819,N_4758);
and U4981 (N_4981,N_4833,N_4873);
nor U4982 (N_4982,N_4816,N_4854);
nand U4983 (N_4983,N_4756,N_4831);
nor U4984 (N_4984,N_4757,N_4844);
or U4985 (N_4985,N_4774,N_4814);
nor U4986 (N_4986,N_4871,N_4778);
xnor U4987 (N_4987,N_4759,N_4828);
nor U4988 (N_4988,N_4752,N_4824);
and U4989 (N_4989,N_4862,N_4801);
xnor U4990 (N_4990,N_4826,N_4827);
and U4991 (N_4991,N_4766,N_4807);
and U4992 (N_4992,N_4821,N_4795);
and U4993 (N_4993,N_4777,N_4856);
xnor U4994 (N_4994,N_4792,N_4850);
nand U4995 (N_4995,N_4771,N_4789);
and U4996 (N_4996,N_4805,N_4841);
xor U4997 (N_4997,N_4772,N_4841);
or U4998 (N_4998,N_4827,N_4848);
or U4999 (N_4999,N_4833,N_4849);
and U5000 (N_5000,N_4968,N_4961);
or U5001 (N_5001,N_4933,N_4997);
and U5002 (N_5002,N_4994,N_4908);
nor U5003 (N_5003,N_4901,N_4934);
and U5004 (N_5004,N_4927,N_4878);
xnor U5005 (N_5005,N_4979,N_4941);
xnor U5006 (N_5006,N_4935,N_4949);
nor U5007 (N_5007,N_4971,N_4930);
nor U5008 (N_5008,N_4890,N_4911);
nand U5009 (N_5009,N_4959,N_4940);
or U5010 (N_5010,N_4889,N_4923);
nor U5011 (N_5011,N_4974,N_4989);
nand U5012 (N_5012,N_4945,N_4980);
xnor U5013 (N_5013,N_4899,N_4972);
and U5014 (N_5014,N_4884,N_4999);
xor U5015 (N_5015,N_4882,N_4932);
xor U5016 (N_5016,N_4938,N_4877);
nand U5017 (N_5017,N_4982,N_4996);
xnor U5018 (N_5018,N_4895,N_4929);
nand U5019 (N_5019,N_4903,N_4969);
and U5020 (N_5020,N_4993,N_4909);
or U5021 (N_5021,N_4954,N_4998);
and U5022 (N_5022,N_4926,N_4946);
and U5023 (N_5023,N_4956,N_4985);
nor U5024 (N_5024,N_4912,N_4944);
or U5025 (N_5025,N_4928,N_4916);
or U5026 (N_5026,N_4883,N_4896);
or U5027 (N_5027,N_4963,N_4966);
or U5028 (N_5028,N_4951,N_4891);
nand U5029 (N_5029,N_4886,N_4914);
nand U5030 (N_5030,N_4892,N_4953);
and U5031 (N_5031,N_4950,N_4981);
nand U5032 (N_5032,N_4918,N_4879);
nor U5033 (N_5033,N_4978,N_4960);
nand U5034 (N_5034,N_4984,N_4900);
nor U5035 (N_5035,N_4965,N_4905);
xor U5036 (N_5036,N_4976,N_4990);
nor U5037 (N_5037,N_4988,N_4983);
nand U5038 (N_5038,N_4977,N_4875);
nand U5039 (N_5039,N_4973,N_4937);
nor U5040 (N_5040,N_4907,N_4902);
nand U5041 (N_5041,N_4995,N_4962);
and U5042 (N_5042,N_4881,N_4936);
or U5043 (N_5043,N_4986,N_4925);
and U5044 (N_5044,N_4948,N_4970);
nor U5045 (N_5045,N_4876,N_4921);
nor U5046 (N_5046,N_4924,N_4922);
or U5047 (N_5047,N_4987,N_4958);
nor U5048 (N_5048,N_4898,N_4919);
and U5049 (N_5049,N_4880,N_4885);
and U5050 (N_5050,N_4888,N_4887);
xnor U5051 (N_5051,N_4952,N_4975);
xnor U5052 (N_5052,N_4910,N_4947);
xnor U5053 (N_5053,N_4964,N_4942);
or U5054 (N_5054,N_4931,N_4991);
xor U5055 (N_5055,N_4893,N_4967);
nand U5056 (N_5056,N_4913,N_4897);
and U5057 (N_5057,N_4955,N_4906);
nand U5058 (N_5058,N_4894,N_4904);
nor U5059 (N_5059,N_4917,N_4992);
nor U5060 (N_5060,N_4915,N_4939);
and U5061 (N_5061,N_4957,N_4943);
or U5062 (N_5062,N_4920,N_4954);
nand U5063 (N_5063,N_4968,N_4952);
xor U5064 (N_5064,N_4932,N_4999);
or U5065 (N_5065,N_4949,N_4901);
and U5066 (N_5066,N_4924,N_4892);
or U5067 (N_5067,N_4961,N_4937);
xnor U5068 (N_5068,N_4913,N_4934);
xnor U5069 (N_5069,N_4967,N_4905);
nand U5070 (N_5070,N_4904,N_4885);
nor U5071 (N_5071,N_4894,N_4925);
nor U5072 (N_5072,N_4947,N_4981);
and U5073 (N_5073,N_4973,N_4955);
xor U5074 (N_5074,N_4898,N_4894);
or U5075 (N_5075,N_4997,N_4976);
nand U5076 (N_5076,N_4998,N_4983);
nand U5077 (N_5077,N_4914,N_4919);
xor U5078 (N_5078,N_4932,N_4917);
xnor U5079 (N_5079,N_4958,N_4925);
xnor U5080 (N_5080,N_4959,N_4998);
or U5081 (N_5081,N_4959,N_4878);
nor U5082 (N_5082,N_4913,N_4997);
and U5083 (N_5083,N_4919,N_4971);
and U5084 (N_5084,N_4983,N_4982);
and U5085 (N_5085,N_4947,N_4965);
and U5086 (N_5086,N_4949,N_4957);
xnor U5087 (N_5087,N_4942,N_4986);
nor U5088 (N_5088,N_4945,N_4902);
nand U5089 (N_5089,N_4999,N_4958);
or U5090 (N_5090,N_4928,N_4988);
nor U5091 (N_5091,N_4877,N_4908);
nand U5092 (N_5092,N_4891,N_4884);
nor U5093 (N_5093,N_4956,N_4971);
or U5094 (N_5094,N_4889,N_4971);
nand U5095 (N_5095,N_4878,N_4962);
and U5096 (N_5096,N_4918,N_4901);
nand U5097 (N_5097,N_4881,N_4939);
xor U5098 (N_5098,N_4930,N_4992);
or U5099 (N_5099,N_4941,N_4982);
xnor U5100 (N_5100,N_4971,N_4942);
or U5101 (N_5101,N_4925,N_4969);
and U5102 (N_5102,N_4897,N_4904);
xor U5103 (N_5103,N_4928,N_4958);
or U5104 (N_5104,N_4924,N_4992);
nand U5105 (N_5105,N_4946,N_4950);
nand U5106 (N_5106,N_4909,N_4963);
and U5107 (N_5107,N_4939,N_4957);
nand U5108 (N_5108,N_4942,N_4953);
nor U5109 (N_5109,N_4909,N_4954);
nand U5110 (N_5110,N_4880,N_4979);
nor U5111 (N_5111,N_4942,N_4998);
nor U5112 (N_5112,N_4933,N_4913);
and U5113 (N_5113,N_4950,N_4884);
and U5114 (N_5114,N_4963,N_4935);
or U5115 (N_5115,N_4981,N_4909);
nor U5116 (N_5116,N_4893,N_4920);
xnor U5117 (N_5117,N_4886,N_4887);
xnor U5118 (N_5118,N_4958,N_4906);
nand U5119 (N_5119,N_4953,N_4998);
and U5120 (N_5120,N_4899,N_4900);
nand U5121 (N_5121,N_4882,N_4945);
nand U5122 (N_5122,N_4940,N_4932);
xnor U5123 (N_5123,N_4924,N_4962);
nand U5124 (N_5124,N_4953,N_4988);
nand U5125 (N_5125,N_5047,N_5009);
or U5126 (N_5126,N_5112,N_5103);
nor U5127 (N_5127,N_5018,N_5066);
nor U5128 (N_5128,N_5013,N_5005);
or U5129 (N_5129,N_5087,N_5029);
nor U5130 (N_5130,N_5043,N_5023);
xor U5131 (N_5131,N_5022,N_5093);
nor U5132 (N_5132,N_5036,N_5086);
or U5133 (N_5133,N_5000,N_5020);
and U5134 (N_5134,N_5069,N_5083);
nand U5135 (N_5135,N_5025,N_5094);
nor U5136 (N_5136,N_5057,N_5031);
nand U5137 (N_5137,N_5104,N_5032);
and U5138 (N_5138,N_5028,N_5105);
nand U5139 (N_5139,N_5120,N_5067);
or U5140 (N_5140,N_5113,N_5001);
nand U5141 (N_5141,N_5034,N_5007);
and U5142 (N_5142,N_5045,N_5004);
nand U5143 (N_5143,N_5095,N_5121);
nand U5144 (N_5144,N_5014,N_5111);
and U5145 (N_5145,N_5116,N_5012);
nor U5146 (N_5146,N_5101,N_5077);
or U5147 (N_5147,N_5107,N_5040);
nand U5148 (N_5148,N_5092,N_5048);
or U5149 (N_5149,N_5085,N_5115);
or U5150 (N_5150,N_5076,N_5065);
and U5151 (N_5151,N_5060,N_5122);
xor U5152 (N_5152,N_5061,N_5068);
and U5153 (N_5153,N_5117,N_5070);
nor U5154 (N_5154,N_5055,N_5044);
nand U5155 (N_5155,N_5006,N_5063);
nand U5156 (N_5156,N_5100,N_5064);
nand U5157 (N_5157,N_5041,N_5072);
or U5158 (N_5158,N_5033,N_5119);
nor U5159 (N_5159,N_5082,N_5016);
nor U5160 (N_5160,N_5114,N_5015);
or U5161 (N_5161,N_5011,N_5075);
or U5162 (N_5162,N_5106,N_5081);
xor U5163 (N_5163,N_5003,N_5054);
nor U5164 (N_5164,N_5089,N_5037);
nor U5165 (N_5165,N_5088,N_5056);
xor U5166 (N_5166,N_5027,N_5039);
or U5167 (N_5167,N_5071,N_5042);
or U5168 (N_5168,N_5035,N_5058);
and U5169 (N_5169,N_5049,N_5024);
nor U5170 (N_5170,N_5051,N_5108);
and U5171 (N_5171,N_5079,N_5099);
nor U5172 (N_5172,N_5059,N_5017);
or U5173 (N_5173,N_5074,N_5124);
nand U5174 (N_5174,N_5038,N_5109);
and U5175 (N_5175,N_5021,N_5050);
nand U5176 (N_5176,N_5110,N_5010);
or U5177 (N_5177,N_5052,N_5097);
and U5178 (N_5178,N_5084,N_5030);
and U5179 (N_5179,N_5090,N_5096);
nor U5180 (N_5180,N_5091,N_5102);
xnor U5181 (N_5181,N_5008,N_5053);
nand U5182 (N_5182,N_5073,N_5026);
nand U5183 (N_5183,N_5046,N_5019);
or U5184 (N_5184,N_5118,N_5078);
xnor U5185 (N_5185,N_5098,N_5080);
xor U5186 (N_5186,N_5062,N_5002);
or U5187 (N_5187,N_5123,N_5111);
nand U5188 (N_5188,N_5020,N_5122);
and U5189 (N_5189,N_5007,N_5102);
and U5190 (N_5190,N_5056,N_5016);
and U5191 (N_5191,N_5063,N_5103);
nand U5192 (N_5192,N_5044,N_5004);
or U5193 (N_5193,N_5028,N_5046);
or U5194 (N_5194,N_5074,N_5103);
or U5195 (N_5195,N_5025,N_5069);
xor U5196 (N_5196,N_5110,N_5063);
nand U5197 (N_5197,N_5001,N_5045);
or U5198 (N_5198,N_5044,N_5086);
nand U5199 (N_5199,N_5076,N_5033);
and U5200 (N_5200,N_5088,N_5028);
or U5201 (N_5201,N_5100,N_5106);
or U5202 (N_5202,N_5026,N_5000);
nand U5203 (N_5203,N_5045,N_5056);
xnor U5204 (N_5204,N_5096,N_5099);
xor U5205 (N_5205,N_5000,N_5101);
nor U5206 (N_5206,N_5112,N_5015);
xnor U5207 (N_5207,N_5023,N_5057);
nand U5208 (N_5208,N_5123,N_5120);
nand U5209 (N_5209,N_5031,N_5116);
or U5210 (N_5210,N_5055,N_5083);
xor U5211 (N_5211,N_5086,N_5006);
nand U5212 (N_5212,N_5089,N_5033);
or U5213 (N_5213,N_5103,N_5056);
or U5214 (N_5214,N_5090,N_5115);
or U5215 (N_5215,N_5101,N_5109);
nor U5216 (N_5216,N_5113,N_5027);
or U5217 (N_5217,N_5016,N_5104);
or U5218 (N_5218,N_5004,N_5042);
xor U5219 (N_5219,N_5017,N_5073);
nor U5220 (N_5220,N_5097,N_5103);
xor U5221 (N_5221,N_5098,N_5033);
and U5222 (N_5222,N_5087,N_5102);
xnor U5223 (N_5223,N_5050,N_5123);
nor U5224 (N_5224,N_5098,N_5056);
and U5225 (N_5225,N_5108,N_5098);
and U5226 (N_5226,N_5073,N_5054);
and U5227 (N_5227,N_5072,N_5039);
or U5228 (N_5228,N_5054,N_5036);
or U5229 (N_5229,N_5072,N_5005);
or U5230 (N_5230,N_5054,N_5041);
xor U5231 (N_5231,N_5092,N_5112);
nor U5232 (N_5232,N_5100,N_5049);
nand U5233 (N_5233,N_5120,N_5046);
xnor U5234 (N_5234,N_5022,N_5040);
and U5235 (N_5235,N_5075,N_5050);
nand U5236 (N_5236,N_5031,N_5021);
or U5237 (N_5237,N_5101,N_5057);
xnor U5238 (N_5238,N_5054,N_5075);
nor U5239 (N_5239,N_5062,N_5084);
nand U5240 (N_5240,N_5106,N_5029);
nor U5241 (N_5241,N_5115,N_5096);
and U5242 (N_5242,N_5103,N_5094);
xnor U5243 (N_5243,N_5002,N_5003);
xor U5244 (N_5244,N_5065,N_5095);
nor U5245 (N_5245,N_5102,N_5078);
or U5246 (N_5246,N_5032,N_5099);
and U5247 (N_5247,N_5070,N_5037);
and U5248 (N_5248,N_5042,N_5073);
nor U5249 (N_5249,N_5036,N_5055);
nor U5250 (N_5250,N_5157,N_5194);
nand U5251 (N_5251,N_5183,N_5181);
nor U5252 (N_5252,N_5148,N_5207);
or U5253 (N_5253,N_5140,N_5163);
and U5254 (N_5254,N_5169,N_5177);
nor U5255 (N_5255,N_5240,N_5125);
xnor U5256 (N_5256,N_5135,N_5137);
and U5257 (N_5257,N_5246,N_5191);
and U5258 (N_5258,N_5198,N_5206);
and U5259 (N_5259,N_5159,N_5220);
and U5260 (N_5260,N_5205,N_5180);
nand U5261 (N_5261,N_5235,N_5166);
or U5262 (N_5262,N_5171,N_5182);
nor U5263 (N_5263,N_5197,N_5192);
nand U5264 (N_5264,N_5151,N_5241);
and U5265 (N_5265,N_5212,N_5215);
and U5266 (N_5266,N_5228,N_5225);
nor U5267 (N_5267,N_5167,N_5203);
nor U5268 (N_5268,N_5146,N_5222);
xor U5269 (N_5269,N_5179,N_5132);
and U5270 (N_5270,N_5243,N_5244);
nand U5271 (N_5271,N_5216,N_5136);
and U5272 (N_5272,N_5161,N_5230);
nor U5273 (N_5273,N_5134,N_5229);
and U5274 (N_5274,N_5144,N_5141);
and U5275 (N_5275,N_5162,N_5208);
and U5276 (N_5276,N_5202,N_5138);
nor U5277 (N_5277,N_5233,N_5178);
or U5278 (N_5278,N_5147,N_5131);
xor U5279 (N_5279,N_5188,N_5145);
xor U5280 (N_5280,N_5217,N_5173);
nor U5281 (N_5281,N_5153,N_5236);
or U5282 (N_5282,N_5195,N_5214);
and U5283 (N_5283,N_5128,N_5142);
nor U5284 (N_5284,N_5237,N_5143);
nor U5285 (N_5285,N_5172,N_5149);
xnor U5286 (N_5286,N_5155,N_5209);
nor U5287 (N_5287,N_5213,N_5218);
nor U5288 (N_5288,N_5187,N_5158);
and U5289 (N_5289,N_5150,N_5126);
nand U5290 (N_5290,N_5224,N_5133);
nand U5291 (N_5291,N_5160,N_5168);
nand U5292 (N_5292,N_5247,N_5219);
or U5293 (N_5293,N_5201,N_5130);
xnor U5294 (N_5294,N_5129,N_5165);
nor U5295 (N_5295,N_5127,N_5184);
nand U5296 (N_5296,N_5175,N_5245);
xor U5297 (N_5297,N_5238,N_5154);
xnor U5298 (N_5298,N_5210,N_5186);
xnor U5299 (N_5299,N_5190,N_5139);
nor U5300 (N_5300,N_5248,N_5232);
nor U5301 (N_5301,N_5164,N_5174);
nor U5302 (N_5302,N_5193,N_5204);
nand U5303 (N_5303,N_5242,N_5239);
and U5304 (N_5304,N_5234,N_5199);
nand U5305 (N_5305,N_5189,N_5170);
nand U5306 (N_5306,N_5211,N_5249);
nor U5307 (N_5307,N_5221,N_5196);
xnor U5308 (N_5308,N_5176,N_5152);
and U5309 (N_5309,N_5226,N_5200);
xor U5310 (N_5310,N_5156,N_5227);
or U5311 (N_5311,N_5223,N_5231);
and U5312 (N_5312,N_5185,N_5219);
nor U5313 (N_5313,N_5142,N_5161);
xnor U5314 (N_5314,N_5208,N_5155);
nor U5315 (N_5315,N_5245,N_5200);
and U5316 (N_5316,N_5174,N_5176);
nand U5317 (N_5317,N_5193,N_5185);
and U5318 (N_5318,N_5154,N_5181);
nor U5319 (N_5319,N_5168,N_5136);
nor U5320 (N_5320,N_5194,N_5141);
xor U5321 (N_5321,N_5127,N_5201);
or U5322 (N_5322,N_5224,N_5188);
and U5323 (N_5323,N_5181,N_5160);
or U5324 (N_5324,N_5170,N_5166);
nor U5325 (N_5325,N_5203,N_5127);
nand U5326 (N_5326,N_5214,N_5222);
nor U5327 (N_5327,N_5171,N_5229);
or U5328 (N_5328,N_5135,N_5206);
nand U5329 (N_5329,N_5126,N_5180);
and U5330 (N_5330,N_5153,N_5226);
and U5331 (N_5331,N_5177,N_5171);
nand U5332 (N_5332,N_5220,N_5246);
nor U5333 (N_5333,N_5149,N_5177);
xnor U5334 (N_5334,N_5222,N_5129);
nand U5335 (N_5335,N_5136,N_5182);
or U5336 (N_5336,N_5154,N_5158);
nor U5337 (N_5337,N_5186,N_5196);
nand U5338 (N_5338,N_5201,N_5185);
nand U5339 (N_5339,N_5185,N_5154);
nand U5340 (N_5340,N_5171,N_5240);
and U5341 (N_5341,N_5217,N_5180);
or U5342 (N_5342,N_5236,N_5224);
nand U5343 (N_5343,N_5132,N_5218);
nand U5344 (N_5344,N_5231,N_5209);
nor U5345 (N_5345,N_5181,N_5193);
and U5346 (N_5346,N_5125,N_5176);
xor U5347 (N_5347,N_5135,N_5185);
nand U5348 (N_5348,N_5233,N_5229);
or U5349 (N_5349,N_5177,N_5220);
or U5350 (N_5350,N_5233,N_5198);
nor U5351 (N_5351,N_5136,N_5221);
nand U5352 (N_5352,N_5144,N_5167);
or U5353 (N_5353,N_5144,N_5226);
nand U5354 (N_5354,N_5169,N_5220);
nand U5355 (N_5355,N_5178,N_5177);
nor U5356 (N_5356,N_5246,N_5239);
nor U5357 (N_5357,N_5220,N_5179);
xor U5358 (N_5358,N_5193,N_5147);
and U5359 (N_5359,N_5126,N_5177);
xnor U5360 (N_5360,N_5222,N_5174);
nor U5361 (N_5361,N_5184,N_5214);
or U5362 (N_5362,N_5215,N_5196);
nand U5363 (N_5363,N_5243,N_5242);
xor U5364 (N_5364,N_5150,N_5140);
and U5365 (N_5365,N_5125,N_5214);
nand U5366 (N_5366,N_5163,N_5214);
nand U5367 (N_5367,N_5193,N_5249);
xor U5368 (N_5368,N_5208,N_5247);
xnor U5369 (N_5369,N_5196,N_5199);
xor U5370 (N_5370,N_5164,N_5234);
or U5371 (N_5371,N_5215,N_5198);
nand U5372 (N_5372,N_5183,N_5173);
nor U5373 (N_5373,N_5204,N_5238);
and U5374 (N_5374,N_5242,N_5223);
xnor U5375 (N_5375,N_5283,N_5313);
or U5376 (N_5376,N_5362,N_5308);
or U5377 (N_5377,N_5258,N_5274);
or U5378 (N_5378,N_5350,N_5312);
and U5379 (N_5379,N_5348,N_5262);
xnor U5380 (N_5380,N_5342,N_5271);
nand U5381 (N_5381,N_5259,N_5358);
nand U5382 (N_5382,N_5336,N_5306);
and U5383 (N_5383,N_5324,N_5325);
and U5384 (N_5384,N_5261,N_5351);
nor U5385 (N_5385,N_5335,N_5367);
xnor U5386 (N_5386,N_5291,N_5373);
and U5387 (N_5387,N_5269,N_5363);
xnor U5388 (N_5388,N_5328,N_5270);
nand U5389 (N_5389,N_5349,N_5294);
nor U5390 (N_5390,N_5332,N_5266);
xnor U5391 (N_5391,N_5366,N_5317);
and U5392 (N_5392,N_5315,N_5357);
nand U5393 (N_5393,N_5343,N_5368);
xor U5394 (N_5394,N_5288,N_5302);
nor U5395 (N_5395,N_5305,N_5278);
nor U5396 (N_5396,N_5322,N_5303);
and U5397 (N_5397,N_5264,N_5285);
nand U5398 (N_5398,N_5293,N_5361);
nand U5399 (N_5399,N_5333,N_5279);
xnor U5400 (N_5400,N_5316,N_5319);
and U5401 (N_5401,N_5296,N_5355);
and U5402 (N_5402,N_5321,N_5370);
and U5403 (N_5403,N_5281,N_5272);
xnor U5404 (N_5404,N_5365,N_5330);
nand U5405 (N_5405,N_5304,N_5356);
nand U5406 (N_5406,N_5299,N_5263);
or U5407 (N_5407,N_5301,N_5295);
or U5408 (N_5408,N_5300,N_5298);
nand U5409 (N_5409,N_5337,N_5275);
or U5410 (N_5410,N_5251,N_5250);
nand U5411 (N_5411,N_5267,N_5360);
and U5412 (N_5412,N_5286,N_5268);
xnor U5413 (N_5413,N_5289,N_5353);
xnor U5414 (N_5414,N_5341,N_5292);
and U5415 (N_5415,N_5329,N_5290);
xnor U5416 (N_5416,N_5372,N_5280);
xnor U5417 (N_5417,N_5257,N_5276);
nand U5418 (N_5418,N_5369,N_5326);
and U5419 (N_5419,N_5297,N_5327);
and U5420 (N_5420,N_5309,N_5273);
or U5421 (N_5421,N_5347,N_5359);
nor U5422 (N_5422,N_5346,N_5345);
or U5423 (N_5423,N_5311,N_5352);
xnor U5424 (N_5424,N_5334,N_5371);
or U5425 (N_5425,N_5339,N_5253);
nand U5426 (N_5426,N_5277,N_5282);
and U5427 (N_5427,N_5340,N_5254);
xor U5428 (N_5428,N_5252,N_5364);
nor U5429 (N_5429,N_5260,N_5265);
nor U5430 (N_5430,N_5314,N_5287);
nand U5431 (N_5431,N_5310,N_5354);
nor U5432 (N_5432,N_5338,N_5255);
xnor U5433 (N_5433,N_5320,N_5256);
or U5434 (N_5434,N_5374,N_5307);
and U5435 (N_5435,N_5318,N_5331);
or U5436 (N_5436,N_5284,N_5344);
nand U5437 (N_5437,N_5323,N_5360);
xnor U5438 (N_5438,N_5271,N_5366);
nor U5439 (N_5439,N_5361,N_5297);
nor U5440 (N_5440,N_5294,N_5363);
nor U5441 (N_5441,N_5253,N_5257);
nor U5442 (N_5442,N_5311,N_5310);
or U5443 (N_5443,N_5315,N_5258);
nor U5444 (N_5444,N_5294,N_5315);
or U5445 (N_5445,N_5314,N_5269);
xnor U5446 (N_5446,N_5359,N_5341);
nand U5447 (N_5447,N_5338,N_5334);
nand U5448 (N_5448,N_5341,N_5271);
nor U5449 (N_5449,N_5367,N_5310);
and U5450 (N_5450,N_5278,N_5357);
nand U5451 (N_5451,N_5352,N_5342);
and U5452 (N_5452,N_5277,N_5342);
or U5453 (N_5453,N_5296,N_5276);
and U5454 (N_5454,N_5315,N_5251);
nand U5455 (N_5455,N_5335,N_5353);
and U5456 (N_5456,N_5285,N_5255);
xnor U5457 (N_5457,N_5310,N_5293);
and U5458 (N_5458,N_5356,N_5267);
nor U5459 (N_5459,N_5329,N_5345);
or U5460 (N_5460,N_5295,N_5320);
or U5461 (N_5461,N_5364,N_5288);
nor U5462 (N_5462,N_5302,N_5282);
and U5463 (N_5463,N_5297,N_5259);
or U5464 (N_5464,N_5356,N_5318);
nor U5465 (N_5465,N_5333,N_5360);
and U5466 (N_5466,N_5340,N_5280);
xor U5467 (N_5467,N_5343,N_5254);
xnor U5468 (N_5468,N_5372,N_5310);
nor U5469 (N_5469,N_5364,N_5320);
or U5470 (N_5470,N_5274,N_5286);
xor U5471 (N_5471,N_5297,N_5276);
nor U5472 (N_5472,N_5338,N_5347);
nor U5473 (N_5473,N_5332,N_5346);
xnor U5474 (N_5474,N_5319,N_5310);
nand U5475 (N_5475,N_5343,N_5373);
or U5476 (N_5476,N_5329,N_5304);
nor U5477 (N_5477,N_5355,N_5316);
and U5478 (N_5478,N_5276,N_5306);
nor U5479 (N_5479,N_5253,N_5346);
and U5480 (N_5480,N_5327,N_5350);
or U5481 (N_5481,N_5292,N_5301);
and U5482 (N_5482,N_5319,N_5293);
nand U5483 (N_5483,N_5343,N_5258);
or U5484 (N_5484,N_5347,N_5252);
nor U5485 (N_5485,N_5252,N_5250);
xnor U5486 (N_5486,N_5352,N_5335);
or U5487 (N_5487,N_5331,N_5329);
nor U5488 (N_5488,N_5254,N_5288);
or U5489 (N_5489,N_5295,N_5319);
nor U5490 (N_5490,N_5309,N_5351);
and U5491 (N_5491,N_5274,N_5339);
or U5492 (N_5492,N_5254,N_5325);
xnor U5493 (N_5493,N_5276,N_5304);
and U5494 (N_5494,N_5293,N_5273);
xor U5495 (N_5495,N_5275,N_5347);
nand U5496 (N_5496,N_5366,N_5373);
nor U5497 (N_5497,N_5300,N_5296);
xnor U5498 (N_5498,N_5339,N_5293);
and U5499 (N_5499,N_5328,N_5304);
nor U5500 (N_5500,N_5478,N_5483);
and U5501 (N_5501,N_5435,N_5484);
xnor U5502 (N_5502,N_5486,N_5445);
and U5503 (N_5503,N_5479,N_5410);
and U5504 (N_5504,N_5381,N_5399);
or U5505 (N_5505,N_5475,N_5403);
and U5506 (N_5506,N_5434,N_5394);
nand U5507 (N_5507,N_5413,N_5468);
and U5508 (N_5508,N_5444,N_5458);
nand U5509 (N_5509,N_5460,N_5491);
nor U5510 (N_5510,N_5455,N_5380);
xor U5511 (N_5511,N_5432,N_5462);
or U5512 (N_5512,N_5390,N_5467);
nand U5513 (N_5513,N_5499,N_5459);
and U5514 (N_5514,N_5383,N_5490);
xor U5515 (N_5515,N_5477,N_5427);
nand U5516 (N_5516,N_5485,N_5431);
xnor U5517 (N_5517,N_5482,N_5471);
or U5518 (N_5518,N_5401,N_5408);
and U5519 (N_5519,N_5418,N_5416);
xor U5520 (N_5520,N_5470,N_5495);
nand U5521 (N_5521,N_5426,N_5451);
and U5522 (N_5522,N_5405,N_5457);
and U5523 (N_5523,N_5385,N_5448);
nand U5524 (N_5524,N_5409,N_5442);
nand U5525 (N_5525,N_5496,N_5430);
or U5526 (N_5526,N_5480,N_5406);
nand U5527 (N_5527,N_5397,N_5447);
nand U5528 (N_5528,N_5481,N_5425);
or U5529 (N_5529,N_5452,N_5454);
xor U5530 (N_5530,N_5439,N_5465);
xor U5531 (N_5531,N_5494,N_5433);
and U5532 (N_5532,N_5396,N_5407);
nor U5533 (N_5533,N_5469,N_5461);
or U5534 (N_5534,N_5423,N_5466);
nor U5535 (N_5535,N_5404,N_5376);
nor U5536 (N_5536,N_5414,N_5489);
nand U5537 (N_5537,N_5443,N_5453);
nand U5538 (N_5538,N_5474,N_5378);
and U5539 (N_5539,N_5386,N_5412);
or U5540 (N_5540,N_5392,N_5382);
and U5541 (N_5541,N_5437,N_5384);
nor U5542 (N_5542,N_5428,N_5456);
nand U5543 (N_5543,N_5436,N_5464);
nor U5544 (N_5544,N_5449,N_5488);
nand U5545 (N_5545,N_5441,N_5417);
and U5546 (N_5546,N_5493,N_5398);
and U5547 (N_5547,N_5377,N_5438);
or U5548 (N_5548,N_5450,N_5487);
nor U5549 (N_5549,N_5422,N_5393);
and U5550 (N_5550,N_5440,N_5389);
and U5551 (N_5551,N_5472,N_5476);
or U5552 (N_5552,N_5492,N_5419);
nand U5553 (N_5553,N_5473,N_5411);
nor U5554 (N_5554,N_5387,N_5388);
nor U5555 (N_5555,N_5395,N_5446);
and U5556 (N_5556,N_5498,N_5429);
nor U5557 (N_5557,N_5421,N_5391);
xnor U5558 (N_5558,N_5497,N_5420);
xnor U5559 (N_5559,N_5463,N_5402);
nand U5560 (N_5560,N_5379,N_5415);
nand U5561 (N_5561,N_5400,N_5424);
or U5562 (N_5562,N_5375,N_5396);
and U5563 (N_5563,N_5408,N_5445);
and U5564 (N_5564,N_5412,N_5483);
and U5565 (N_5565,N_5426,N_5474);
and U5566 (N_5566,N_5407,N_5394);
or U5567 (N_5567,N_5378,N_5456);
nand U5568 (N_5568,N_5398,N_5473);
xnor U5569 (N_5569,N_5413,N_5419);
nand U5570 (N_5570,N_5497,N_5379);
nor U5571 (N_5571,N_5493,N_5443);
xnor U5572 (N_5572,N_5402,N_5437);
nand U5573 (N_5573,N_5472,N_5437);
nor U5574 (N_5574,N_5454,N_5403);
nor U5575 (N_5575,N_5436,N_5382);
and U5576 (N_5576,N_5423,N_5412);
and U5577 (N_5577,N_5438,N_5490);
or U5578 (N_5578,N_5414,N_5444);
and U5579 (N_5579,N_5388,N_5391);
nand U5580 (N_5580,N_5377,N_5447);
nor U5581 (N_5581,N_5491,N_5471);
nand U5582 (N_5582,N_5379,N_5488);
nand U5583 (N_5583,N_5449,N_5413);
nand U5584 (N_5584,N_5439,N_5422);
or U5585 (N_5585,N_5379,N_5417);
xor U5586 (N_5586,N_5446,N_5420);
and U5587 (N_5587,N_5378,N_5479);
nand U5588 (N_5588,N_5428,N_5397);
nand U5589 (N_5589,N_5416,N_5403);
and U5590 (N_5590,N_5442,N_5419);
nor U5591 (N_5591,N_5492,N_5471);
xor U5592 (N_5592,N_5395,N_5418);
nand U5593 (N_5593,N_5488,N_5375);
nor U5594 (N_5594,N_5494,N_5480);
xnor U5595 (N_5595,N_5451,N_5429);
xor U5596 (N_5596,N_5387,N_5496);
or U5597 (N_5597,N_5394,N_5473);
nor U5598 (N_5598,N_5435,N_5421);
xor U5599 (N_5599,N_5429,N_5410);
nor U5600 (N_5600,N_5425,N_5381);
or U5601 (N_5601,N_5389,N_5477);
nor U5602 (N_5602,N_5406,N_5427);
xnor U5603 (N_5603,N_5419,N_5386);
and U5604 (N_5604,N_5379,N_5445);
xnor U5605 (N_5605,N_5425,N_5403);
or U5606 (N_5606,N_5481,N_5410);
nand U5607 (N_5607,N_5429,N_5430);
nor U5608 (N_5608,N_5419,N_5440);
nand U5609 (N_5609,N_5484,N_5378);
nor U5610 (N_5610,N_5397,N_5418);
nor U5611 (N_5611,N_5471,N_5385);
or U5612 (N_5612,N_5479,N_5476);
xor U5613 (N_5613,N_5392,N_5468);
or U5614 (N_5614,N_5464,N_5411);
or U5615 (N_5615,N_5417,N_5462);
nor U5616 (N_5616,N_5403,N_5375);
or U5617 (N_5617,N_5385,N_5427);
nand U5618 (N_5618,N_5376,N_5456);
nor U5619 (N_5619,N_5377,N_5385);
and U5620 (N_5620,N_5381,N_5428);
nor U5621 (N_5621,N_5413,N_5406);
and U5622 (N_5622,N_5495,N_5477);
and U5623 (N_5623,N_5449,N_5387);
xnor U5624 (N_5624,N_5428,N_5451);
nor U5625 (N_5625,N_5591,N_5580);
or U5626 (N_5626,N_5547,N_5574);
and U5627 (N_5627,N_5603,N_5508);
and U5628 (N_5628,N_5548,N_5618);
and U5629 (N_5629,N_5620,N_5537);
xnor U5630 (N_5630,N_5573,N_5583);
and U5631 (N_5631,N_5585,N_5578);
xor U5632 (N_5632,N_5598,N_5563);
nor U5633 (N_5633,N_5516,N_5588);
and U5634 (N_5634,N_5560,N_5557);
nand U5635 (N_5635,N_5538,N_5503);
nand U5636 (N_5636,N_5599,N_5522);
nand U5637 (N_5637,N_5619,N_5505);
nand U5638 (N_5638,N_5621,N_5512);
nor U5639 (N_5639,N_5504,N_5587);
xor U5640 (N_5640,N_5514,N_5553);
and U5641 (N_5641,N_5612,N_5622);
xnor U5642 (N_5642,N_5554,N_5546);
nor U5643 (N_5643,N_5534,N_5523);
nand U5644 (N_5644,N_5525,N_5519);
nor U5645 (N_5645,N_5543,N_5624);
nand U5646 (N_5646,N_5582,N_5604);
nand U5647 (N_5647,N_5536,N_5524);
xor U5648 (N_5648,N_5531,N_5507);
or U5649 (N_5649,N_5510,N_5608);
xor U5650 (N_5650,N_5500,N_5579);
nor U5651 (N_5651,N_5567,N_5530);
or U5652 (N_5652,N_5575,N_5571);
nor U5653 (N_5653,N_5518,N_5556);
and U5654 (N_5654,N_5517,N_5590);
xnor U5655 (N_5655,N_5610,N_5542);
xnor U5656 (N_5656,N_5589,N_5607);
nor U5657 (N_5657,N_5555,N_5562);
or U5658 (N_5658,N_5602,N_5515);
xnor U5659 (N_5659,N_5564,N_5606);
or U5660 (N_5660,N_5509,N_5558);
nor U5661 (N_5661,N_5511,N_5595);
nor U5662 (N_5662,N_5615,N_5529);
or U5663 (N_5663,N_5513,N_5594);
and U5664 (N_5664,N_5541,N_5597);
xor U5665 (N_5665,N_5539,N_5570);
or U5666 (N_5666,N_5623,N_5600);
or U5667 (N_5667,N_5586,N_5501);
nor U5668 (N_5668,N_5527,N_5616);
nor U5669 (N_5669,N_5532,N_5561);
nand U5670 (N_5670,N_5601,N_5568);
and U5671 (N_5671,N_5569,N_5520);
or U5672 (N_5672,N_5540,N_5550);
nand U5673 (N_5673,N_5581,N_5614);
nand U5674 (N_5674,N_5605,N_5609);
xnor U5675 (N_5675,N_5528,N_5545);
nor U5676 (N_5676,N_5576,N_5566);
or U5677 (N_5677,N_5535,N_5617);
xnor U5678 (N_5678,N_5533,N_5544);
and U5679 (N_5679,N_5592,N_5502);
and U5680 (N_5680,N_5577,N_5506);
nand U5681 (N_5681,N_5593,N_5596);
nor U5682 (N_5682,N_5613,N_5549);
or U5683 (N_5683,N_5559,N_5526);
xor U5684 (N_5684,N_5521,N_5565);
nor U5685 (N_5685,N_5611,N_5552);
or U5686 (N_5686,N_5572,N_5551);
or U5687 (N_5687,N_5584,N_5569);
or U5688 (N_5688,N_5513,N_5600);
nand U5689 (N_5689,N_5600,N_5586);
nand U5690 (N_5690,N_5551,N_5594);
nor U5691 (N_5691,N_5507,N_5506);
xor U5692 (N_5692,N_5577,N_5601);
or U5693 (N_5693,N_5612,N_5595);
nor U5694 (N_5694,N_5504,N_5600);
xnor U5695 (N_5695,N_5583,N_5523);
and U5696 (N_5696,N_5543,N_5607);
or U5697 (N_5697,N_5619,N_5581);
and U5698 (N_5698,N_5534,N_5581);
nor U5699 (N_5699,N_5551,N_5586);
and U5700 (N_5700,N_5609,N_5525);
xor U5701 (N_5701,N_5501,N_5599);
xnor U5702 (N_5702,N_5584,N_5573);
nor U5703 (N_5703,N_5517,N_5501);
nand U5704 (N_5704,N_5539,N_5522);
nand U5705 (N_5705,N_5508,N_5589);
or U5706 (N_5706,N_5617,N_5612);
or U5707 (N_5707,N_5540,N_5572);
nand U5708 (N_5708,N_5546,N_5571);
nor U5709 (N_5709,N_5618,N_5586);
or U5710 (N_5710,N_5534,N_5570);
nand U5711 (N_5711,N_5521,N_5605);
nor U5712 (N_5712,N_5581,N_5516);
nor U5713 (N_5713,N_5560,N_5502);
nand U5714 (N_5714,N_5513,N_5537);
and U5715 (N_5715,N_5516,N_5546);
xor U5716 (N_5716,N_5571,N_5617);
and U5717 (N_5717,N_5571,N_5605);
nor U5718 (N_5718,N_5617,N_5555);
nand U5719 (N_5719,N_5502,N_5574);
and U5720 (N_5720,N_5559,N_5567);
xor U5721 (N_5721,N_5617,N_5505);
or U5722 (N_5722,N_5501,N_5597);
or U5723 (N_5723,N_5518,N_5589);
or U5724 (N_5724,N_5585,N_5604);
and U5725 (N_5725,N_5542,N_5526);
and U5726 (N_5726,N_5544,N_5585);
and U5727 (N_5727,N_5584,N_5577);
or U5728 (N_5728,N_5621,N_5502);
xnor U5729 (N_5729,N_5614,N_5525);
or U5730 (N_5730,N_5503,N_5520);
nand U5731 (N_5731,N_5616,N_5523);
and U5732 (N_5732,N_5556,N_5603);
nand U5733 (N_5733,N_5611,N_5576);
and U5734 (N_5734,N_5578,N_5576);
or U5735 (N_5735,N_5574,N_5508);
and U5736 (N_5736,N_5602,N_5573);
xor U5737 (N_5737,N_5515,N_5618);
nand U5738 (N_5738,N_5556,N_5559);
and U5739 (N_5739,N_5608,N_5505);
nor U5740 (N_5740,N_5547,N_5582);
nor U5741 (N_5741,N_5598,N_5613);
or U5742 (N_5742,N_5556,N_5502);
nand U5743 (N_5743,N_5508,N_5576);
or U5744 (N_5744,N_5527,N_5548);
or U5745 (N_5745,N_5550,N_5553);
and U5746 (N_5746,N_5546,N_5579);
nor U5747 (N_5747,N_5507,N_5613);
xor U5748 (N_5748,N_5528,N_5510);
and U5749 (N_5749,N_5594,N_5555);
nand U5750 (N_5750,N_5709,N_5651);
and U5751 (N_5751,N_5675,N_5710);
nor U5752 (N_5752,N_5741,N_5670);
xor U5753 (N_5753,N_5706,N_5717);
xor U5754 (N_5754,N_5668,N_5657);
nand U5755 (N_5755,N_5679,N_5639);
nand U5756 (N_5756,N_5676,N_5723);
nand U5757 (N_5757,N_5678,N_5677);
or U5758 (N_5758,N_5733,N_5705);
and U5759 (N_5759,N_5626,N_5748);
xnor U5760 (N_5760,N_5652,N_5707);
and U5761 (N_5761,N_5701,N_5711);
or U5762 (N_5762,N_5745,N_5735);
xor U5763 (N_5763,N_5704,N_5728);
xor U5764 (N_5764,N_5700,N_5642);
nor U5765 (N_5765,N_5649,N_5714);
nand U5766 (N_5766,N_5713,N_5637);
nand U5767 (N_5767,N_5742,N_5662);
or U5768 (N_5768,N_5654,N_5731);
or U5769 (N_5769,N_5665,N_5724);
nor U5770 (N_5770,N_5743,N_5659);
and U5771 (N_5771,N_5722,N_5632);
nor U5772 (N_5772,N_5739,N_5736);
or U5773 (N_5773,N_5744,N_5640);
or U5774 (N_5774,N_5631,N_5727);
xor U5775 (N_5775,N_5645,N_5650);
xnor U5776 (N_5776,N_5692,N_5697);
or U5777 (N_5777,N_5694,N_5720);
xnor U5778 (N_5778,N_5680,N_5635);
or U5779 (N_5779,N_5691,N_5708);
nand U5780 (N_5780,N_5684,N_5730);
nor U5781 (N_5781,N_5702,N_5669);
nor U5782 (N_5782,N_5667,N_5629);
nor U5783 (N_5783,N_5740,N_5673);
nand U5784 (N_5784,N_5718,N_5746);
nand U5785 (N_5785,N_5647,N_5627);
and U5786 (N_5786,N_5671,N_5695);
or U5787 (N_5787,N_5686,N_5698);
nand U5788 (N_5788,N_5658,N_5726);
and U5789 (N_5789,N_5656,N_5699);
and U5790 (N_5790,N_5719,N_5625);
nand U5791 (N_5791,N_5663,N_5747);
and U5792 (N_5792,N_5683,N_5688);
nor U5793 (N_5793,N_5634,N_5636);
and U5794 (N_5794,N_5738,N_5655);
nor U5795 (N_5795,N_5661,N_5690);
or U5796 (N_5796,N_5696,N_5681);
and U5797 (N_5797,N_5712,N_5630);
or U5798 (N_5798,N_5725,N_5664);
or U5799 (N_5799,N_5672,N_5653);
or U5800 (N_5800,N_5732,N_5703);
xor U5801 (N_5801,N_5721,N_5628);
and U5802 (N_5802,N_5643,N_5644);
or U5803 (N_5803,N_5749,N_5666);
xor U5804 (N_5804,N_5715,N_5734);
nor U5805 (N_5805,N_5689,N_5674);
nand U5806 (N_5806,N_5729,N_5737);
xnor U5807 (N_5807,N_5682,N_5633);
xnor U5808 (N_5808,N_5646,N_5641);
xor U5809 (N_5809,N_5687,N_5685);
xor U5810 (N_5810,N_5648,N_5693);
and U5811 (N_5811,N_5660,N_5716);
and U5812 (N_5812,N_5638,N_5692);
nor U5813 (N_5813,N_5729,N_5657);
or U5814 (N_5814,N_5722,N_5678);
nand U5815 (N_5815,N_5688,N_5686);
nor U5816 (N_5816,N_5676,N_5657);
and U5817 (N_5817,N_5635,N_5746);
nor U5818 (N_5818,N_5682,N_5629);
and U5819 (N_5819,N_5706,N_5684);
or U5820 (N_5820,N_5634,N_5737);
or U5821 (N_5821,N_5632,N_5744);
and U5822 (N_5822,N_5692,N_5698);
or U5823 (N_5823,N_5726,N_5732);
xnor U5824 (N_5824,N_5696,N_5629);
xor U5825 (N_5825,N_5716,N_5651);
nand U5826 (N_5826,N_5716,N_5672);
xnor U5827 (N_5827,N_5735,N_5724);
nand U5828 (N_5828,N_5633,N_5726);
nor U5829 (N_5829,N_5744,N_5724);
nand U5830 (N_5830,N_5646,N_5642);
xnor U5831 (N_5831,N_5637,N_5634);
and U5832 (N_5832,N_5670,N_5633);
and U5833 (N_5833,N_5648,N_5714);
nand U5834 (N_5834,N_5670,N_5650);
and U5835 (N_5835,N_5718,N_5650);
and U5836 (N_5836,N_5745,N_5733);
nor U5837 (N_5837,N_5739,N_5695);
nand U5838 (N_5838,N_5657,N_5672);
or U5839 (N_5839,N_5648,N_5727);
xor U5840 (N_5840,N_5695,N_5639);
xor U5841 (N_5841,N_5746,N_5645);
or U5842 (N_5842,N_5641,N_5711);
and U5843 (N_5843,N_5655,N_5668);
and U5844 (N_5844,N_5679,N_5685);
nand U5845 (N_5845,N_5640,N_5698);
xnor U5846 (N_5846,N_5667,N_5648);
nor U5847 (N_5847,N_5683,N_5743);
nor U5848 (N_5848,N_5628,N_5656);
nand U5849 (N_5849,N_5713,N_5645);
and U5850 (N_5850,N_5742,N_5628);
and U5851 (N_5851,N_5747,N_5739);
nor U5852 (N_5852,N_5685,N_5671);
xor U5853 (N_5853,N_5652,N_5676);
xnor U5854 (N_5854,N_5704,N_5651);
and U5855 (N_5855,N_5672,N_5631);
xor U5856 (N_5856,N_5664,N_5737);
xnor U5857 (N_5857,N_5639,N_5668);
nor U5858 (N_5858,N_5651,N_5638);
nand U5859 (N_5859,N_5683,N_5681);
nand U5860 (N_5860,N_5668,N_5650);
and U5861 (N_5861,N_5732,N_5632);
nand U5862 (N_5862,N_5699,N_5660);
nor U5863 (N_5863,N_5639,N_5739);
nor U5864 (N_5864,N_5706,N_5645);
and U5865 (N_5865,N_5717,N_5674);
and U5866 (N_5866,N_5691,N_5683);
nand U5867 (N_5867,N_5663,N_5689);
and U5868 (N_5868,N_5664,N_5738);
and U5869 (N_5869,N_5717,N_5748);
or U5870 (N_5870,N_5696,N_5705);
nor U5871 (N_5871,N_5630,N_5637);
and U5872 (N_5872,N_5634,N_5643);
nand U5873 (N_5873,N_5740,N_5715);
xnor U5874 (N_5874,N_5749,N_5687);
nand U5875 (N_5875,N_5772,N_5811);
or U5876 (N_5876,N_5789,N_5756);
xnor U5877 (N_5877,N_5774,N_5841);
xor U5878 (N_5878,N_5752,N_5804);
xor U5879 (N_5879,N_5819,N_5853);
and U5880 (N_5880,N_5805,N_5848);
nor U5881 (N_5881,N_5767,N_5806);
or U5882 (N_5882,N_5765,N_5801);
nand U5883 (N_5883,N_5840,N_5854);
nand U5884 (N_5884,N_5809,N_5778);
nor U5885 (N_5885,N_5834,N_5863);
and U5886 (N_5886,N_5861,N_5779);
nor U5887 (N_5887,N_5781,N_5783);
xnor U5888 (N_5888,N_5808,N_5855);
or U5889 (N_5889,N_5803,N_5828);
nand U5890 (N_5890,N_5835,N_5792);
or U5891 (N_5891,N_5817,N_5825);
nand U5892 (N_5892,N_5826,N_5844);
or U5893 (N_5893,N_5857,N_5800);
nand U5894 (N_5894,N_5799,N_5754);
and U5895 (N_5895,N_5793,N_5874);
and U5896 (N_5896,N_5818,N_5852);
nand U5897 (N_5897,N_5813,N_5823);
xnor U5898 (N_5898,N_5764,N_5788);
or U5899 (N_5899,N_5870,N_5768);
nand U5900 (N_5900,N_5777,N_5751);
nor U5901 (N_5901,N_5784,N_5860);
and U5902 (N_5902,N_5866,N_5833);
or U5903 (N_5903,N_5830,N_5821);
nor U5904 (N_5904,N_5786,N_5760);
xnor U5905 (N_5905,N_5865,N_5753);
nand U5906 (N_5906,N_5859,N_5780);
xor U5907 (N_5907,N_5815,N_5842);
nor U5908 (N_5908,N_5869,N_5790);
or U5909 (N_5909,N_5814,N_5795);
or U5910 (N_5910,N_5824,N_5791);
nor U5911 (N_5911,N_5755,N_5766);
xor U5912 (N_5912,N_5782,N_5812);
and U5913 (N_5913,N_5871,N_5836);
and U5914 (N_5914,N_5831,N_5757);
nor U5915 (N_5915,N_5838,N_5750);
and U5916 (N_5916,N_5763,N_5820);
or U5917 (N_5917,N_5851,N_5873);
nor U5918 (N_5918,N_5797,N_5775);
nand U5919 (N_5919,N_5794,N_5769);
and U5920 (N_5920,N_5802,N_5868);
or U5921 (N_5921,N_5807,N_5856);
and U5922 (N_5922,N_5845,N_5771);
xnor U5923 (N_5923,N_5770,N_5864);
nor U5924 (N_5924,N_5867,N_5858);
or U5925 (N_5925,N_5785,N_5787);
xnor U5926 (N_5926,N_5839,N_5759);
or U5927 (N_5927,N_5816,N_5837);
nand U5928 (N_5928,N_5829,N_5810);
xor U5929 (N_5929,N_5832,N_5827);
or U5930 (N_5930,N_5798,N_5846);
or U5931 (N_5931,N_5862,N_5847);
xnor U5932 (N_5932,N_5849,N_5822);
nor U5933 (N_5933,N_5762,N_5776);
xnor U5934 (N_5934,N_5843,N_5773);
or U5935 (N_5935,N_5796,N_5758);
nor U5936 (N_5936,N_5872,N_5761);
xor U5937 (N_5937,N_5850,N_5798);
and U5938 (N_5938,N_5826,N_5847);
nand U5939 (N_5939,N_5860,N_5851);
nor U5940 (N_5940,N_5847,N_5756);
or U5941 (N_5941,N_5801,N_5836);
nand U5942 (N_5942,N_5774,N_5751);
nand U5943 (N_5943,N_5844,N_5840);
and U5944 (N_5944,N_5843,N_5755);
and U5945 (N_5945,N_5805,N_5833);
or U5946 (N_5946,N_5772,N_5764);
nor U5947 (N_5947,N_5813,N_5833);
nand U5948 (N_5948,N_5838,N_5806);
nor U5949 (N_5949,N_5784,N_5812);
nand U5950 (N_5950,N_5786,N_5752);
and U5951 (N_5951,N_5818,N_5830);
nand U5952 (N_5952,N_5824,N_5750);
nand U5953 (N_5953,N_5839,N_5751);
or U5954 (N_5954,N_5868,N_5796);
or U5955 (N_5955,N_5874,N_5777);
or U5956 (N_5956,N_5820,N_5808);
xor U5957 (N_5957,N_5863,N_5754);
xnor U5958 (N_5958,N_5840,N_5782);
and U5959 (N_5959,N_5750,N_5835);
xnor U5960 (N_5960,N_5818,N_5772);
nand U5961 (N_5961,N_5820,N_5865);
or U5962 (N_5962,N_5863,N_5824);
nand U5963 (N_5963,N_5836,N_5775);
xnor U5964 (N_5964,N_5790,N_5825);
xnor U5965 (N_5965,N_5777,N_5783);
or U5966 (N_5966,N_5754,N_5858);
and U5967 (N_5967,N_5840,N_5816);
nor U5968 (N_5968,N_5869,N_5843);
and U5969 (N_5969,N_5764,N_5820);
or U5970 (N_5970,N_5801,N_5759);
and U5971 (N_5971,N_5807,N_5784);
nand U5972 (N_5972,N_5872,N_5856);
nor U5973 (N_5973,N_5839,N_5802);
or U5974 (N_5974,N_5813,N_5816);
or U5975 (N_5975,N_5844,N_5813);
nor U5976 (N_5976,N_5779,N_5808);
nand U5977 (N_5977,N_5777,N_5794);
and U5978 (N_5978,N_5842,N_5824);
nand U5979 (N_5979,N_5786,N_5865);
nand U5980 (N_5980,N_5809,N_5870);
xor U5981 (N_5981,N_5868,N_5811);
nor U5982 (N_5982,N_5787,N_5783);
nand U5983 (N_5983,N_5806,N_5853);
or U5984 (N_5984,N_5803,N_5863);
and U5985 (N_5985,N_5754,N_5752);
or U5986 (N_5986,N_5776,N_5766);
nand U5987 (N_5987,N_5783,N_5775);
nand U5988 (N_5988,N_5827,N_5788);
nand U5989 (N_5989,N_5821,N_5779);
nand U5990 (N_5990,N_5834,N_5807);
nor U5991 (N_5991,N_5816,N_5750);
nor U5992 (N_5992,N_5807,N_5824);
nand U5993 (N_5993,N_5794,N_5776);
nand U5994 (N_5994,N_5816,N_5800);
and U5995 (N_5995,N_5856,N_5811);
or U5996 (N_5996,N_5857,N_5852);
and U5997 (N_5997,N_5823,N_5787);
xnor U5998 (N_5998,N_5813,N_5766);
or U5999 (N_5999,N_5780,N_5788);
nand U6000 (N_6000,N_5920,N_5956);
or U6001 (N_6001,N_5935,N_5985);
nand U6002 (N_6002,N_5960,N_5962);
or U6003 (N_6003,N_5999,N_5988);
or U6004 (N_6004,N_5877,N_5959);
xor U6005 (N_6005,N_5885,N_5943);
and U6006 (N_6006,N_5970,N_5924);
or U6007 (N_6007,N_5986,N_5979);
nand U6008 (N_6008,N_5977,N_5890);
nor U6009 (N_6009,N_5881,N_5949);
and U6010 (N_6010,N_5934,N_5968);
or U6011 (N_6011,N_5973,N_5906);
nand U6012 (N_6012,N_5895,N_5992);
and U6013 (N_6013,N_5897,N_5940);
nand U6014 (N_6014,N_5904,N_5997);
and U6015 (N_6015,N_5909,N_5886);
and U6016 (N_6016,N_5899,N_5880);
and U6017 (N_6017,N_5954,N_5927);
and U6018 (N_6018,N_5916,N_5894);
or U6019 (N_6019,N_5896,N_5878);
and U6020 (N_6020,N_5946,N_5998);
nand U6021 (N_6021,N_5942,N_5939);
nand U6022 (N_6022,N_5995,N_5963);
nor U6023 (N_6023,N_5913,N_5883);
nand U6024 (N_6024,N_5975,N_5993);
nor U6025 (N_6025,N_5907,N_5961);
nor U6026 (N_6026,N_5965,N_5969);
nor U6027 (N_6027,N_5987,N_5966);
and U6028 (N_6028,N_5978,N_5936);
nor U6029 (N_6029,N_5951,N_5955);
nand U6030 (N_6030,N_5910,N_5923);
xnor U6031 (N_6031,N_5928,N_5991);
or U6032 (N_6032,N_5914,N_5911);
or U6033 (N_6033,N_5900,N_5938);
xnor U6034 (N_6034,N_5989,N_5950);
nand U6035 (N_6035,N_5958,N_5994);
xnor U6036 (N_6036,N_5887,N_5903);
nand U6037 (N_6037,N_5980,N_5929);
and U6038 (N_6038,N_5957,N_5931);
xnor U6039 (N_6039,N_5884,N_5937);
or U6040 (N_6040,N_5948,N_5901);
nor U6041 (N_6041,N_5932,N_5976);
or U6042 (N_6042,N_5889,N_5945);
or U6043 (N_6043,N_5982,N_5930);
and U6044 (N_6044,N_5990,N_5882);
or U6045 (N_6045,N_5875,N_5926);
or U6046 (N_6046,N_5891,N_5971);
xor U6047 (N_6047,N_5933,N_5876);
or U6048 (N_6048,N_5925,N_5905);
nor U6049 (N_6049,N_5908,N_5893);
nand U6050 (N_6050,N_5898,N_5947);
and U6051 (N_6051,N_5879,N_5892);
nor U6052 (N_6052,N_5983,N_5941);
nor U6053 (N_6053,N_5953,N_5921);
xor U6054 (N_6054,N_5888,N_5917);
or U6055 (N_6055,N_5974,N_5919);
or U6056 (N_6056,N_5964,N_5984);
xor U6057 (N_6057,N_5915,N_5967);
nand U6058 (N_6058,N_5944,N_5918);
or U6059 (N_6059,N_5972,N_5912);
xor U6060 (N_6060,N_5981,N_5922);
xor U6061 (N_6061,N_5996,N_5952);
nand U6062 (N_6062,N_5902,N_5885);
and U6063 (N_6063,N_5930,N_5895);
or U6064 (N_6064,N_5888,N_5947);
or U6065 (N_6065,N_5875,N_5986);
nor U6066 (N_6066,N_5961,N_5945);
nand U6067 (N_6067,N_5891,N_5882);
and U6068 (N_6068,N_5929,N_5949);
nand U6069 (N_6069,N_5980,N_5911);
nor U6070 (N_6070,N_5975,N_5904);
nor U6071 (N_6071,N_5968,N_5925);
nor U6072 (N_6072,N_5982,N_5971);
nor U6073 (N_6073,N_5884,N_5878);
xnor U6074 (N_6074,N_5917,N_5985);
nand U6075 (N_6075,N_5881,N_5979);
xnor U6076 (N_6076,N_5936,N_5933);
and U6077 (N_6077,N_5920,N_5951);
and U6078 (N_6078,N_5897,N_5911);
or U6079 (N_6079,N_5966,N_5897);
nor U6080 (N_6080,N_5976,N_5894);
nand U6081 (N_6081,N_5891,N_5975);
nor U6082 (N_6082,N_5971,N_5905);
nand U6083 (N_6083,N_5905,N_5956);
and U6084 (N_6084,N_5877,N_5997);
or U6085 (N_6085,N_5906,N_5945);
or U6086 (N_6086,N_5927,N_5937);
xnor U6087 (N_6087,N_5886,N_5878);
nand U6088 (N_6088,N_5989,N_5891);
xnor U6089 (N_6089,N_5921,N_5942);
xnor U6090 (N_6090,N_5988,N_5889);
xor U6091 (N_6091,N_5896,N_5938);
nor U6092 (N_6092,N_5956,N_5972);
or U6093 (N_6093,N_5949,N_5986);
or U6094 (N_6094,N_5898,N_5961);
and U6095 (N_6095,N_5895,N_5886);
or U6096 (N_6096,N_5907,N_5973);
xnor U6097 (N_6097,N_5891,N_5982);
nand U6098 (N_6098,N_5916,N_5891);
and U6099 (N_6099,N_5882,N_5935);
nand U6100 (N_6100,N_5976,N_5921);
xor U6101 (N_6101,N_5879,N_5991);
xor U6102 (N_6102,N_5969,N_5954);
nor U6103 (N_6103,N_5967,N_5882);
and U6104 (N_6104,N_5962,N_5957);
xor U6105 (N_6105,N_5912,N_5880);
and U6106 (N_6106,N_5991,N_5997);
xnor U6107 (N_6107,N_5906,N_5921);
xnor U6108 (N_6108,N_5973,N_5966);
xnor U6109 (N_6109,N_5905,N_5994);
and U6110 (N_6110,N_5951,N_5943);
or U6111 (N_6111,N_5977,N_5973);
nand U6112 (N_6112,N_5992,N_5909);
and U6113 (N_6113,N_5933,N_5961);
or U6114 (N_6114,N_5884,N_5899);
nand U6115 (N_6115,N_5944,N_5989);
or U6116 (N_6116,N_5938,N_5943);
nor U6117 (N_6117,N_5916,N_5885);
nand U6118 (N_6118,N_5921,N_5933);
or U6119 (N_6119,N_5943,N_5877);
or U6120 (N_6120,N_5925,N_5994);
xnor U6121 (N_6121,N_5935,N_5977);
and U6122 (N_6122,N_5951,N_5892);
or U6123 (N_6123,N_5993,N_5977);
xor U6124 (N_6124,N_5899,N_5910);
xor U6125 (N_6125,N_6108,N_6069);
nor U6126 (N_6126,N_6085,N_6019);
nand U6127 (N_6127,N_6083,N_6098);
and U6128 (N_6128,N_6096,N_6119);
and U6129 (N_6129,N_6052,N_6065);
xnor U6130 (N_6130,N_6056,N_6023);
or U6131 (N_6131,N_6020,N_6018);
nand U6132 (N_6132,N_6113,N_6072);
nor U6133 (N_6133,N_6058,N_6022);
nand U6134 (N_6134,N_6059,N_6114);
or U6135 (N_6135,N_6051,N_6097);
or U6136 (N_6136,N_6042,N_6102);
xnor U6137 (N_6137,N_6062,N_6036);
xor U6138 (N_6138,N_6079,N_6037);
xnor U6139 (N_6139,N_6112,N_6034);
xnor U6140 (N_6140,N_6060,N_6015);
or U6141 (N_6141,N_6088,N_6117);
xnor U6142 (N_6142,N_6009,N_6092);
nor U6143 (N_6143,N_6045,N_6087);
nor U6144 (N_6144,N_6067,N_6103);
xor U6145 (N_6145,N_6082,N_6038);
nand U6146 (N_6146,N_6120,N_6109);
nand U6147 (N_6147,N_6106,N_6002);
and U6148 (N_6148,N_6055,N_6046);
nand U6149 (N_6149,N_6063,N_6021);
nand U6150 (N_6150,N_6100,N_6124);
nand U6151 (N_6151,N_6074,N_6010);
nor U6152 (N_6152,N_6025,N_6066);
and U6153 (N_6153,N_6013,N_6064);
or U6154 (N_6154,N_6110,N_6073);
nor U6155 (N_6155,N_6090,N_6123);
or U6156 (N_6156,N_6027,N_6057);
or U6157 (N_6157,N_6047,N_6000);
or U6158 (N_6158,N_6026,N_6029);
or U6159 (N_6159,N_6121,N_6054);
nand U6160 (N_6160,N_6122,N_6031);
xor U6161 (N_6161,N_6091,N_6099);
nor U6162 (N_6162,N_6017,N_6086);
or U6163 (N_6163,N_6115,N_6118);
and U6164 (N_6164,N_6101,N_6039);
xnor U6165 (N_6165,N_6070,N_6048);
and U6166 (N_6166,N_6077,N_6075);
and U6167 (N_6167,N_6068,N_6016);
nand U6168 (N_6168,N_6094,N_6005);
xor U6169 (N_6169,N_6105,N_6071);
nor U6170 (N_6170,N_6028,N_6111);
nor U6171 (N_6171,N_6012,N_6004);
or U6172 (N_6172,N_6050,N_6024);
or U6173 (N_6173,N_6053,N_6089);
nor U6174 (N_6174,N_6006,N_6080);
nor U6175 (N_6175,N_6044,N_6107);
and U6176 (N_6176,N_6095,N_6003);
and U6177 (N_6177,N_6104,N_6040);
nor U6178 (N_6178,N_6084,N_6035);
or U6179 (N_6179,N_6061,N_6081);
xor U6180 (N_6180,N_6078,N_6116);
and U6181 (N_6181,N_6076,N_6030);
xnor U6182 (N_6182,N_6014,N_6043);
xnor U6183 (N_6183,N_6041,N_6093);
nand U6184 (N_6184,N_6011,N_6008);
nor U6185 (N_6185,N_6033,N_6032);
nor U6186 (N_6186,N_6007,N_6001);
xor U6187 (N_6187,N_6049,N_6113);
and U6188 (N_6188,N_6053,N_6013);
or U6189 (N_6189,N_6096,N_6078);
or U6190 (N_6190,N_6108,N_6079);
and U6191 (N_6191,N_6014,N_6030);
nor U6192 (N_6192,N_6094,N_6111);
nand U6193 (N_6193,N_6087,N_6093);
nand U6194 (N_6194,N_6114,N_6042);
and U6195 (N_6195,N_6060,N_6003);
nor U6196 (N_6196,N_6035,N_6061);
or U6197 (N_6197,N_6028,N_6117);
nor U6198 (N_6198,N_6076,N_6091);
and U6199 (N_6199,N_6111,N_6108);
nor U6200 (N_6200,N_6073,N_6028);
xor U6201 (N_6201,N_6099,N_6065);
or U6202 (N_6202,N_6092,N_6000);
xor U6203 (N_6203,N_6063,N_6073);
or U6204 (N_6204,N_6008,N_6053);
nand U6205 (N_6205,N_6034,N_6060);
or U6206 (N_6206,N_6124,N_6122);
nand U6207 (N_6207,N_6090,N_6074);
nand U6208 (N_6208,N_6062,N_6050);
nand U6209 (N_6209,N_6090,N_6054);
nor U6210 (N_6210,N_6088,N_6116);
nand U6211 (N_6211,N_6069,N_6086);
nor U6212 (N_6212,N_6042,N_6098);
and U6213 (N_6213,N_6086,N_6038);
and U6214 (N_6214,N_6108,N_6039);
and U6215 (N_6215,N_6089,N_6056);
xor U6216 (N_6216,N_6013,N_6113);
and U6217 (N_6217,N_6084,N_6104);
or U6218 (N_6218,N_6035,N_6086);
xor U6219 (N_6219,N_6015,N_6065);
xnor U6220 (N_6220,N_6061,N_6010);
xor U6221 (N_6221,N_6014,N_6054);
nor U6222 (N_6222,N_6024,N_6010);
nand U6223 (N_6223,N_6082,N_6024);
or U6224 (N_6224,N_6025,N_6080);
xnor U6225 (N_6225,N_6104,N_6116);
xnor U6226 (N_6226,N_6074,N_6063);
or U6227 (N_6227,N_6112,N_6056);
nand U6228 (N_6228,N_6003,N_6098);
nor U6229 (N_6229,N_6023,N_6011);
nor U6230 (N_6230,N_6063,N_6025);
xnor U6231 (N_6231,N_6019,N_6120);
nor U6232 (N_6232,N_6013,N_6060);
nand U6233 (N_6233,N_6104,N_6067);
nor U6234 (N_6234,N_6059,N_6086);
and U6235 (N_6235,N_6016,N_6048);
or U6236 (N_6236,N_6057,N_6025);
nand U6237 (N_6237,N_6102,N_6123);
or U6238 (N_6238,N_6019,N_6005);
nand U6239 (N_6239,N_6088,N_6065);
and U6240 (N_6240,N_6014,N_6007);
nor U6241 (N_6241,N_6116,N_6081);
and U6242 (N_6242,N_6121,N_6109);
xor U6243 (N_6243,N_6090,N_6102);
nor U6244 (N_6244,N_6055,N_6043);
xnor U6245 (N_6245,N_6100,N_6115);
nor U6246 (N_6246,N_6048,N_6066);
nand U6247 (N_6247,N_6025,N_6102);
and U6248 (N_6248,N_6074,N_6050);
xnor U6249 (N_6249,N_6042,N_6101);
nand U6250 (N_6250,N_6225,N_6143);
nand U6251 (N_6251,N_6141,N_6163);
xnor U6252 (N_6252,N_6155,N_6179);
and U6253 (N_6253,N_6127,N_6247);
nand U6254 (N_6254,N_6140,N_6165);
nor U6255 (N_6255,N_6215,N_6133);
nor U6256 (N_6256,N_6187,N_6193);
nand U6257 (N_6257,N_6139,N_6241);
or U6258 (N_6258,N_6181,N_6232);
nand U6259 (N_6259,N_6239,N_6176);
nand U6260 (N_6260,N_6168,N_6147);
nand U6261 (N_6261,N_6214,N_6200);
nand U6262 (N_6262,N_6229,N_6244);
or U6263 (N_6263,N_6189,N_6138);
and U6264 (N_6264,N_6210,N_6228);
nand U6265 (N_6265,N_6175,N_6135);
xor U6266 (N_6266,N_6172,N_6167);
nand U6267 (N_6267,N_6243,N_6185);
nor U6268 (N_6268,N_6131,N_6171);
xnor U6269 (N_6269,N_6240,N_6150);
or U6270 (N_6270,N_6157,N_6158);
and U6271 (N_6271,N_6156,N_6197);
xnor U6272 (N_6272,N_6132,N_6195);
or U6273 (N_6273,N_6216,N_6169);
xor U6274 (N_6274,N_6130,N_6166);
nor U6275 (N_6275,N_6242,N_6209);
nand U6276 (N_6276,N_6170,N_6180);
nor U6277 (N_6277,N_6148,N_6173);
xnor U6278 (N_6278,N_6192,N_6217);
and U6279 (N_6279,N_6161,N_6142);
and U6280 (N_6280,N_6178,N_6211);
xnor U6281 (N_6281,N_6224,N_6238);
xor U6282 (N_6282,N_6134,N_6198);
nand U6283 (N_6283,N_6226,N_6154);
xor U6284 (N_6284,N_6153,N_6246);
and U6285 (N_6285,N_6223,N_6159);
nor U6286 (N_6286,N_6212,N_6191);
nand U6287 (N_6287,N_6236,N_6233);
and U6288 (N_6288,N_6206,N_6162);
or U6289 (N_6289,N_6151,N_6207);
nor U6290 (N_6290,N_6199,N_6136);
xnor U6291 (N_6291,N_6203,N_6227);
or U6292 (N_6292,N_6230,N_6164);
and U6293 (N_6293,N_6248,N_6202);
and U6294 (N_6294,N_6222,N_6218);
xnor U6295 (N_6295,N_6149,N_6186);
xor U6296 (N_6296,N_6144,N_6213);
or U6297 (N_6297,N_6125,N_6188);
nor U6298 (N_6298,N_6177,N_6249);
nor U6299 (N_6299,N_6201,N_6146);
or U6300 (N_6300,N_6219,N_6182);
nand U6301 (N_6301,N_6208,N_6129);
nand U6302 (N_6302,N_6174,N_6235);
nand U6303 (N_6303,N_6137,N_6184);
or U6304 (N_6304,N_6190,N_6221);
and U6305 (N_6305,N_6128,N_6145);
nand U6306 (N_6306,N_6220,N_6205);
nor U6307 (N_6307,N_6204,N_6152);
and U6308 (N_6308,N_6234,N_6245);
and U6309 (N_6309,N_6237,N_6160);
and U6310 (N_6310,N_6183,N_6126);
nand U6311 (N_6311,N_6231,N_6194);
nor U6312 (N_6312,N_6196,N_6137);
nand U6313 (N_6313,N_6233,N_6129);
and U6314 (N_6314,N_6141,N_6240);
nand U6315 (N_6315,N_6191,N_6160);
or U6316 (N_6316,N_6227,N_6220);
nand U6317 (N_6317,N_6190,N_6173);
nand U6318 (N_6318,N_6185,N_6249);
or U6319 (N_6319,N_6137,N_6201);
nand U6320 (N_6320,N_6196,N_6248);
or U6321 (N_6321,N_6156,N_6192);
nor U6322 (N_6322,N_6159,N_6188);
nand U6323 (N_6323,N_6128,N_6190);
nand U6324 (N_6324,N_6215,N_6210);
or U6325 (N_6325,N_6167,N_6128);
nand U6326 (N_6326,N_6243,N_6154);
nand U6327 (N_6327,N_6154,N_6248);
nor U6328 (N_6328,N_6220,N_6184);
nor U6329 (N_6329,N_6193,N_6157);
xnor U6330 (N_6330,N_6191,N_6151);
nor U6331 (N_6331,N_6226,N_6143);
xor U6332 (N_6332,N_6143,N_6243);
xor U6333 (N_6333,N_6240,N_6225);
nand U6334 (N_6334,N_6154,N_6138);
nand U6335 (N_6335,N_6249,N_6243);
nand U6336 (N_6336,N_6204,N_6161);
nor U6337 (N_6337,N_6182,N_6165);
nand U6338 (N_6338,N_6193,N_6191);
and U6339 (N_6339,N_6222,N_6166);
nand U6340 (N_6340,N_6131,N_6183);
and U6341 (N_6341,N_6162,N_6177);
nor U6342 (N_6342,N_6157,N_6218);
nand U6343 (N_6343,N_6244,N_6228);
or U6344 (N_6344,N_6223,N_6200);
xor U6345 (N_6345,N_6153,N_6179);
nor U6346 (N_6346,N_6202,N_6145);
nor U6347 (N_6347,N_6206,N_6239);
nand U6348 (N_6348,N_6223,N_6144);
nand U6349 (N_6349,N_6154,N_6237);
nor U6350 (N_6350,N_6196,N_6174);
and U6351 (N_6351,N_6244,N_6152);
and U6352 (N_6352,N_6180,N_6165);
nand U6353 (N_6353,N_6139,N_6205);
and U6354 (N_6354,N_6164,N_6183);
xnor U6355 (N_6355,N_6173,N_6229);
xor U6356 (N_6356,N_6206,N_6225);
nor U6357 (N_6357,N_6163,N_6204);
xor U6358 (N_6358,N_6233,N_6143);
xor U6359 (N_6359,N_6206,N_6172);
and U6360 (N_6360,N_6218,N_6155);
nor U6361 (N_6361,N_6145,N_6191);
xnor U6362 (N_6362,N_6201,N_6162);
xnor U6363 (N_6363,N_6179,N_6207);
nor U6364 (N_6364,N_6240,N_6189);
or U6365 (N_6365,N_6208,N_6179);
and U6366 (N_6366,N_6172,N_6179);
and U6367 (N_6367,N_6131,N_6166);
or U6368 (N_6368,N_6236,N_6141);
and U6369 (N_6369,N_6182,N_6210);
nor U6370 (N_6370,N_6219,N_6130);
and U6371 (N_6371,N_6210,N_6185);
or U6372 (N_6372,N_6141,N_6213);
or U6373 (N_6373,N_6170,N_6155);
nand U6374 (N_6374,N_6133,N_6227);
or U6375 (N_6375,N_6324,N_6274);
nand U6376 (N_6376,N_6347,N_6306);
and U6377 (N_6377,N_6320,N_6361);
or U6378 (N_6378,N_6261,N_6270);
xnor U6379 (N_6379,N_6354,N_6372);
or U6380 (N_6380,N_6289,N_6342);
nand U6381 (N_6381,N_6327,N_6281);
or U6382 (N_6382,N_6262,N_6346);
and U6383 (N_6383,N_6283,N_6338);
xor U6384 (N_6384,N_6254,N_6301);
nand U6385 (N_6385,N_6318,N_6370);
and U6386 (N_6386,N_6334,N_6287);
and U6387 (N_6387,N_6250,N_6294);
and U6388 (N_6388,N_6272,N_6276);
xnor U6389 (N_6389,N_6308,N_6331);
or U6390 (N_6390,N_6352,N_6312);
nand U6391 (N_6391,N_6298,N_6268);
nand U6392 (N_6392,N_6323,N_6357);
or U6393 (N_6393,N_6315,N_6310);
or U6394 (N_6394,N_6348,N_6297);
or U6395 (N_6395,N_6269,N_6366);
nor U6396 (N_6396,N_6286,N_6260);
nor U6397 (N_6397,N_6311,N_6358);
and U6398 (N_6398,N_6314,N_6282);
xor U6399 (N_6399,N_6295,N_6267);
nor U6400 (N_6400,N_6316,N_6374);
and U6401 (N_6401,N_6319,N_6359);
or U6402 (N_6402,N_6309,N_6371);
and U6403 (N_6403,N_6362,N_6292);
nand U6404 (N_6404,N_6252,N_6322);
nor U6405 (N_6405,N_6367,N_6266);
or U6406 (N_6406,N_6313,N_6326);
nand U6407 (N_6407,N_6344,N_6263);
or U6408 (N_6408,N_6332,N_6337);
or U6409 (N_6409,N_6328,N_6304);
nand U6410 (N_6410,N_6363,N_6345);
or U6411 (N_6411,N_6341,N_6339);
xnor U6412 (N_6412,N_6356,N_6273);
nor U6413 (N_6413,N_6299,N_6291);
and U6414 (N_6414,N_6307,N_6271);
and U6415 (N_6415,N_6296,N_6277);
and U6416 (N_6416,N_6373,N_6364);
xor U6417 (N_6417,N_6259,N_6251);
and U6418 (N_6418,N_6349,N_6253);
or U6419 (N_6419,N_6293,N_6335);
nand U6420 (N_6420,N_6265,N_6284);
or U6421 (N_6421,N_6350,N_6290);
or U6422 (N_6422,N_6336,N_6280);
or U6423 (N_6423,N_6275,N_6255);
nor U6424 (N_6424,N_6325,N_6351);
and U6425 (N_6425,N_6355,N_6258);
and U6426 (N_6426,N_6369,N_6329);
and U6427 (N_6427,N_6256,N_6368);
xnor U6428 (N_6428,N_6365,N_6303);
nor U6429 (N_6429,N_6279,N_6343);
xor U6430 (N_6430,N_6264,N_6257);
xor U6431 (N_6431,N_6340,N_6300);
and U6432 (N_6432,N_6330,N_6285);
and U6433 (N_6433,N_6321,N_6360);
and U6434 (N_6434,N_6305,N_6302);
xor U6435 (N_6435,N_6333,N_6353);
nand U6436 (N_6436,N_6278,N_6317);
and U6437 (N_6437,N_6288,N_6291);
nor U6438 (N_6438,N_6327,N_6311);
or U6439 (N_6439,N_6360,N_6277);
nor U6440 (N_6440,N_6257,N_6374);
nand U6441 (N_6441,N_6287,N_6322);
nor U6442 (N_6442,N_6342,N_6261);
nand U6443 (N_6443,N_6371,N_6290);
and U6444 (N_6444,N_6302,N_6277);
and U6445 (N_6445,N_6303,N_6351);
nand U6446 (N_6446,N_6260,N_6280);
and U6447 (N_6447,N_6250,N_6374);
nand U6448 (N_6448,N_6326,N_6303);
nand U6449 (N_6449,N_6294,N_6307);
nor U6450 (N_6450,N_6340,N_6272);
or U6451 (N_6451,N_6364,N_6257);
nor U6452 (N_6452,N_6290,N_6352);
and U6453 (N_6453,N_6353,N_6346);
nor U6454 (N_6454,N_6253,N_6286);
or U6455 (N_6455,N_6310,N_6304);
nand U6456 (N_6456,N_6263,N_6328);
or U6457 (N_6457,N_6342,N_6254);
xnor U6458 (N_6458,N_6324,N_6251);
or U6459 (N_6459,N_6330,N_6367);
or U6460 (N_6460,N_6337,N_6366);
or U6461 (N_6461,N_6326,N_6366);
nand U6462 (N_6462,N_6318,N_6369);
nor U6463 (N_6463,N_6299,N_6256);
or U6464 (N_6464,N_6347,N_6297);
nor U6465 (N_6465,N_6289,N_6307);
nand U6466 (N_6466,N_6349,N_6266);
nor U6467 (N_6467,N_6289,N_6374);
nor U6468 (N_6468,N_6291,N_6358);
or U6469 (N_6469,N_6322,N_6298);
and U6470 (N_6470,N_6359,N_6276);
and U6471 (N_6471,N_6281,N_6286);
nor U6472 (N_6472,N_6288,N_6332);
nand U6473 (N_6473,N_6289,N_6265);
and U6474 (N_6474,N_6322,N_6374);
nand U6475 (N_6475,N_6317,N_6289);
and U6476 (N_6476,N_6271,N_6322);
and U6477 (N_6477,N_6291,N_6374);
and U6478 (N_6478,N_6350,N_6314);
or U6479 (N_6479,N_6292,N_6274);
or U6480 (N_6480,N_6312,N_6251);
nand U6481 (N_6481,N_6292,N_6349);
or U6482 (N_6482,N_6282,N_6340);
xor U6483 (N_6483,N_6347,N_6317);
or U6484 (N_6484,N_6272,N_6307);
or U6485 (N_6485,N_6329,N_6348);
or U6486 (N_6486,N_6270,N_6285);
or U6487 (N_6487,N_6363,N_6357);
xnor U6488 (N_6488,N_6299,N_6307);
nor U6489 (N_6489,N_6372,N_6346);
nand U6490 (N_6490,N_6350,N_6331);
or U6491 (N_6491,N_6334,N_6360);
and U6492 (N_6492,N_6254,N_6359);
nand U6493 (N_6493,N_6355,N_6300);
nor U6494 (N_6494,N_6284,N_6293);
and U6495 (N_6495,N_6309,N_6351);
and U6496 (N_6496,N_6308,N_6299);
xor U6497 (N_6497,N_6328,N_6365);
and U6498 (N_6498,N_6266,N_6373);
nor U6499 (N_6499,N_6351,N_6354);
or U6500 (N_6500,N_6455,N_6464);
or U6501 (N_6501,N_6487,N_6486);
nand U6502 (N_6502,N_6476,N_6461);
and U6503 (N_6503,N_6438,N_6459);
xor U6504 (N_6504,N_6386,N_6403);
nand U6505 (N_6505,N_6389,N_6467);
and U6506 (N_6506,N_6397,N_6456);
xor U6507 (N_6507,N_6430,N_6451);
xnor U6508 (N_6508,N_6423,N_6485);
xnor U6509 (N_6509,N_6379,N_6382);
and U6510 (N_6510,N_6463,N_6499);
and U6511 (N_6511,N_6484,N_6473);
nand U6512 (N_6512,N_6458,N_6385);
nand U6513 (N_6513,N_6471,N_6483);
nand U6514 (N_6514,N_6401,N_6470);
xor U6515 (N_6515,N_6462,N_6425);
and U6516 (N_6516,N_6394,N_6468);
nand U6517 (N_6517,N_6497,N_6406);
nor U6518 (N_6518,N_6413,N_6465);
and U6519 (N_6519,N_6410,N_6436);
xor U6520 (N_6520,N_6432,N_6404);
or U6521 (N_6521,N_6439,N_6444);
and U6522 (N_6522,N_6417,N_6431);
nor U6523 (N_6523,N_6492,N_6447);
and U6524 (N_6524,N_6489,N_6445);
nor U6525 (N_6525,N_6493,N_6494);
or U6526 (N_6526,N_6449,N_6435);
xnor U6527 (N_6527,N_6388,N_6478);
nor U6528 (N_6528,N_6407,N_6405);
nand U6529 (N_6529,N_6391,N_6384);
and U6530 (N_6530,N_6427,N_6452);
and U6531 (N_6531,N_6383,N_6433);
and U6532 (N_6532,N_6390,N_6420);
xnor U6533 (N_6533,N_6426,N_6479);
nand U6534 (N_6534,N_6442,N_6443);
nand U6535 (N_6535,N_6375,N_6472);
nand U6536 (N_6536,N_6460,N_6491);
nor U6537 (N_6537,N_6482,N_6378);
and U6538 (N_6538,N_6408,N_6469);
xnor U6539 (N_6539,N_6419,N_6399);
and U6540 (N_6540,N_6429,N_6498);
xnor U6541 (N_6541,N_6488,N_6396);
and U6542 (N_6542,N_6412,N_6414);
nand U6543 (N_6543,N_6400,N_6422);
nand U6544 (N_6544,N_6437,N_6450);
and U6545 (N_6545,N_6377,N_6474);
or U6546 (N_6546,N_6424,N_6380);
or U6547 (N_6547,N_6392,N_6466);
xnor U6548 (N_6548,N_6454,N_6415);
and U6549 (N_6549,N_6490,N_6428);
and U6550 (N_6550,N_6440,N_6448);
nor U6551 (N_6551,N_6411,N_6477);
nor U6552 (N_6552,N_6446,N_6496);
nand U6553 (N_6553,N_6421,N_6480);
xor U6554 (N_6554,N_6434,N_6398);
and U6555 (N_6555,N_6381,N_6376);
xor U6556 (N_6556,N_6402,N_6481);
or U6557 (N_6557,N_6457,N_6395);
or U6558 (N_6558,N_6393,N_6453);
nor U6559 (N_6559,N_6441,N_6409);
xor U6560 (N_6560,N_6475,N_6418);
nor U6561 (N_6561,N_6495,N_6416);
nor U6562 (N_6562,N_6387,N_6403);
nor U6563 (N_6563,N_6426,N_6437);
nand U6564 (N_6564,N_6492,N_6385);
nand U6565 (N_6565,N_6411,N_6440);
or U6566 (N_6566,N_6428,N_6454);
xor U6567 (N_6567,N_6440,N_6423);
and U6568 (N_6568,N_6461,N_6441);
and U6569 (N_6569,N_6473,N_6476);
and U6570 (N_6570,N_6429,N_6378);
nand U6571 (N_6571,N_6417,N_6390);
xnor U6572 (N_6572,N_6467,N_6440);
nor U6573 (N_6573,N_6419,N_6499);
and U6574 (N_6574,N_6402,N_6386);
and U6575 (N_6575,N_6455,N_6378);
or U6576 (N_6576,N_6494,N_6491);
xnor U6577 (N_6577,N_6435,N_6436);
nand U6578 (N_6578,N_6427,N_6472);
or U6579 (N_6579,N_6440,N_6408);
and U6580 (N_6580,N_6424,N_6461);
xor U6581 (N_6581,N_6491,N_6487);
nor U6582 (N_6582,N_6448,N_6496);
or U6583 (N_6583,N_6444,N_6420);
nor U6584 (N_6584,N_6433,N_6446);
and U6585 (N_6585,N_6382,N_6474);
and U6586 (N_6586,N_6392,N_6445);
nor U6587 (N_6587,N_6390,N_6401);
or U6588 (N_6588,N_6459,N_6436);
and U6589 (N_6589,N_6429,N_6404);
nand U6590 (N_6590,N_6438,N_6492);
or U6591 (N_6591,N_6497,N_6426);
nand U6592 (N_6592,N_6463,N_6474);
xor U6593 (N_6593,N_6439,N_6450);
xor U6594 (N_6594,N_6456,N_6495);
nand U6595 (N_6595,N_6388,N_6441);
xor U6596 (N_6596,N_6455,N_6462);
nor U6597 (N_6597,N_6459,N_6401);
nor U6598 (N_6598,N_6400,N_6383);
nand U6599 (N_6599,N_6376,N_6423);
xnor U6600 (N_6600,N_6433,N_6418);
nor U6601 (N_6601,N_6433,N_6377);
and U6602 (N_6602,N_6412,N_6432);
nand U6603 (N_6603,N_6419,N_6436);
nand U6604 (N_6604,N_6378,N_6452);
or U6605 (N_6605,N_6487,N_6453);
and U6606 (N_6606,N_6447,N_6464);
nor U6607 (N_6607,N_6412,N_6461);
and U6608 (N_6608,N_6409,N_6474);
or U6609 (N_6609,N_6409,N_6458);
and U6610 (N_6610,N_6427,N_6419);
nor U6611 (N_6611,N_6444,N_6401);
nand U6612 (N_6612,N_6423,N_6412);
xnor U6613 (N_6613,N_6452,N_6494);
nand U6614 (N_6614,N_6439,N_6479);
nand U6615 (N_6615,N_6385,N_6461);
xor U6616 (N_6616,N_6497,N_6392);
xnor U6617 (N_6617,N_6379,N_6473);
xnor U6618 (N_6618,N_6478,N_6437);
xnor U6619 (N_6619,N_6459,N_6481);
nand U6620 (N_6620,N_6397,N_6380);
or U6621 (N_6621,N_6467,N_6424);
nand U6622 (N_6622,N_6465,N_6445);
xnor U6623 (N_6623,N_6401,N_6462);
nand U6624 (N_6624,N_6465,N_6475);
or U6625 (N_6625,N_6543,N_6513);
xor U6626 (N_6626,N_6528,N_6618);
nand U6627 (N_6627,N_6590,N_6538);
or U6628 (N_6628,N_6612,N_6525);
and U6629 (N_6629,N_6584,N_6502);
nor U6630 (N_6630,N_6539,N_6515);
and U6631 (N_6631,N_6597,N_6517);
xnor U6632 (N_6632,N_6586,N_6554);
nor U6633 (N_6633,N_6556,N_6519);
nand U6634 (N_6634,N_6552,N_6545);
nand U6635 (N_6635,N_6593,N_6582);
or U6636 (N_6636,N_6544,N_6533);
and U6637 (N_6637,N_6537,N_6621);
or U6638 (N_6638,N_6588,N_6561);
nand U6639 (N_6639,N_6574,N_6548);
nand U6640 (N_6640,N_6595,N_6576);
and U6641 (N_6641,N_6564,N_6572);
nand U6642 (N_6642,N_6523,N_6606);
or U6643 (N_6643,N_6547,N_6542);
nor U6644 (N_6644,N_6617,N_6506);
or U6645 (N_6645,N_6596,N_6592);
or U6646 (N_6646,N_6504,N_6550);
or U6647 (N_6647,N_6591,N_6585);
nor U6648 (N_6648,N_6553,N_6580);
and U6649 (N_6649,N_6579,N_6536);
nand U6650 (N_6650,N_6503,N_6534);
nor U6651 (N_6651,N_6581,N_6594);
or U6652 (N_6652,N_6583,N_6609);
nor U6653 (N_6653,N_6568,N_6524);
nor U6654 (N_6654,N_6604,N_6551);
nand U6655 (N_6655,N_6616,N_6600);
nand U6656 (N_6656,N_6510,N_6611);
xnor U6657 (N_6657,N_6546,N_6516);
and U6658 (N_6658,N_6535,N_6615);
and U6659 (N_6659,N_6607,N_6602);
nand U6660 (N_6660,N_6549,N_6622);
or U6661 (N_6661,N_6613,N_6540);
and U6662 (N_6662,N_6587,N_6575);
and U6663 (N_6663,N_6507,N_6577);
nor U6664 (N_6664,N_6619,N_6541);
and U6665 (N_6665,N_6505,N_6555);
or U6666 (N_6666,N_6514,N_6559);
nor U6667 (N_6667,N_6501,N_6601);
nor U6668 (N_6668,N_6521,N_6500);
nand U6669 (N_6669,N_6624,N_6511);
xor U6670 (N_6670,N_6532,N_6557);
or U6671 (N_6671,N_6569,N_6623);
or U6672 (N_6672,N_6560,N_6527);
nand U6673 (N_6673,N_6526,N_6598);
and U6674 (N_6674,N_6620,N_6599);
or U6675 (N_6675,N_6520,N_6566);
xor U6676 (N_6676,N_6570,N_6562);
xor U6677 (N_6677,N_6522,N_6605);
xor U6678 (N_6678,N_6509,N_6531);
or U6679 (N_6679,N_6589,N_6518);
nor U6680 (N_6680,N_6565,N_6578);
or U6681 (N_6681,N_6608,N_6563);
and U6682 (N_6682,N_6603,N_6573);
and U6683 (N_6683,N_6530,N_6614);
nand U6684 (N_6684,N_6610,N_6571);
and U6685 (N_6685,N_6558,N_6512);
or U6686 (N_6686,N_6529,N_6567);
xor U6687 (N_6687,N_6508,N_6506);
nand U6688 (N_6688,N_6512,N_6522);
nor U6689 (N_6689,N_6591,N_6572);
or U6690 (N_6690,N_6508,N_6568);
or U6691 (N_6691,N_6591,N_6623);
or U6692 (N_6692,N_6619,N_6602);
and U6693 (N_6693,N_6535,N_6504);
nand U6694 (N_6694,N_6603,N_6563);
or U6695 (N_6695,N_6556,N_6538);
xor U6696 (N_6696,N_6576,N_6617);
nand U6697 (N_6697,N_6538,N_6543);
xor U6698 (N_6698,N_6540,N_6623);
and U6699 (N_6699,N_6580,N_6545);
nor U6700 (N_6700,N_6556,N_6508);
xor U6701 (N_6701,N_6580,N_6563);
nor U6702 (N_6702,N_6525,N_6538);
or U6703 (N_6703,N_6619,N_6600);
xor U6704 (N_6704,N_6577,N_6516);
or U6705 (N_6705,N_6540,N_6562);
and U6706 (N_6706,N_6580,N_6538);
and U6707 (N_6707,N_6523,N_6601);
nor U6708 (N_6708,N_6608,N_6555);
and U6709 (N_6709,N_6592,N_6606);
nand U6710 (N_6710,N_6549,N_6566);
or U6711 (N_6711,N_6614,N_6572);
nand U6712 (N_6712,N_6619,N_6507);
nor U6713 (N_6713,N_6603,N_6538);
or U6714 (N_6714,N_6520,N_6522);
xor U6715 (N_6715,N_6515,N_6581);
and U6716 (N_6716,N_6503,N_6605);
xnor U6717 (N_6717,N_6524,N_6603);
and U6718 (N_6718,N_6572,N_6524);
and U6719 (N_6719,N_6570,N_6621);
xor U6720 (N_6720,N_6623,N_6624);
nor U6721 (N_6721,N_6575,N_6608);
or U6722 (N_6722,N_6554,N_6601);
xnor U6723 (N_6723,N_6533,N_6585);
xor U6724 (N_6724,N_6547,N_6562);
xor U6725 (N_6725,N_6533,N_6569);
nor U6726 (N_6726,N_6578,N_6510);
or U6727 (N_6727,N_6557,N_6608);
or U6728 (N_6728,N_6597,N_6576);
nor U6729 (N_6729,N_6535,N_6521);
xnor U6730 (N_6730,N_6608,N_6584);
nor U6731 (N_6731,N_6554,N_6506);
nor U6732 (N_6732,N_6527,N_6559);
nor U6733 (N_6733,N_6574,N_6591);
and U6734 (N_6734,N_6505,N_6582);
or U6735 (N_6735,N_6594,N_6513);
nor U6736 (N_6736,N_6567,N_6615);
xnor U6737 (N_6737,N_6533,N_6546);
nor U6738 (N_6738,N_6525,N_6545);
nand U6739 (N_6739,N_6536,N_6537);
and U6740 (N_6740,N_6507,N_6532);
nor U6741 (N_6741,N_6532,N_6503);
and U6742 (N_6742,N_6502,N_6528);
xor U6743 (N_6743,N_6521,N_6511);
nor U6744 (N_6744,N_6578,N_6539);
nor U6745 (N_6745,N_6614,N_6521);
xor U6746 (N_6746,N_6522,N_6518);
nor U6747 (N_6747,N_6621,N_6573);
nor U6748 (N_6748,N_6608,N_6538);
nor U6749 (N_6749,N_6605,N_6589);
or U6750 (N_6750,N_6711,N_6632);
nand U6751 (N_6751,N_6707,N_6696);
or U6752 (N_6752,N_6689,N_6662);
nand U6753 (N_6753,N_6686,N_6684);
and U6754 (N_6754,N_6736,N_6641);
or U6755 (N_6755,N_6625,N_6636);
or U6756 (N_6756,N_6743,N_6635);
nor U6757 (N_6757,N_6650,N_6727);
nor U6758 (N_6758,N_6681,N_6687);
and U6759 (N_6759,N_6638,N_6725);
xnor U6760 (N_6760,N_6730,N_6648);
xor U6761 (N_6761,N_6649,N_6693);
or U6762 (N_6762,N_6735,N_6633);
and U6763 (N_6763,N_6685,N_6690);
xnor U6764 (N_6764,N_6669,N_6676);
nand U6765 (N_6765,N_6717,N_6700);
and U6766 (N_6766,N_6733,N_6668);
or U6767 (N_6767,N_6708,N_6691);
nand U6768 (N_6768,N_6709,N_6723);
or U6769 (N_6769,N_6626,N_6722);
and U6770 (N_6770,N_6739,N_6705);
and U6771 (N_6771,N_6653,N_6639);
and U6772 (N_6772,N_6721,N_6694);
or U6773 (N_6773,N_6679,N_6629);
nor U6774 (N_6774,N_6628,N_6703);
nand U6775 (N_6775,N_6719,N_6695);
nand U6776 (N_6776,N_6664,N_6715);
xnor U6777 (N_6777,N_6637,N_6688);
nor U6778 (N_6778,N_6665,N_6652);
or U6779 (N_6779,N_6671,N_6682);
nor U6780 (N_6780,N_6673,N_6646);
nor U6781 (N_6781,N_6718,N_6670);
or U6782 (N_6782,N_6713,N_6701);
nand U6783 (N_6783,N_6658,N_6657);
xor U6784 (N_6784,N_6698,N_6627);
nor U6785 (N_6785,N_6643,N_6748);
nor U6786 (N_6786,N_6738,N_6675);
nor U6787 (N_6787,N_6645,N_6660);
nor U6788 (N_6788,N_6654,N_6702);
and U6789 (N_6789,N_6745,N_6699);
and U6790 (N_6790,N_6631,N_6729);
nand U6791 (N_6791,N_6644,N_6661);
nand U6792 (N_6792,N_6720,N_6744);
nor U6793 (N_6793,N_6732,N_6642);
xnor U6794 (N_6794,N_6749,N_6674);
or U6795 (N_6795,N_6634,N_6647);
nor U6796 (N_6796,N_6737,N_6666);
xnor U6797 (N_6797,N_6710,N_6734);
and U6798 (N_6798,N_6640,N_6692);
nor U6799 (N_6799,N_6747,N_6740);
or U6800 (N_6800,N_6697,N_6672);
xor U6801 (N_6801,N_6704,N_6741);
nor U6802 (N_6802,N_6716,N_6728);
and U6803 (N_6803,N_6630,N_6655);
nand U6804 (N_6804,N_6659,N_6714);
xnor U6805 (N_6805,N_6680,N_6706);
xnor U6806 (N_6806,N_6667,N_6746);
nand U6807 (N_6807,N_6656,N_6683);
nand U6808 (N_6808,N_6726,N_6712);
nand U6809 (N_6809,N_6677,N_6663);
and U6810 (N_6810,N_6724,N_6731);
nand U6811 (N_6811,N_6651,N_6678);
nand U6812 (N_6812,N_6742,N_6722);
xnor U6813 (N_6813,N_6740,N_6691);
nor U6814 (N_6814,N_6719,N_6650);
nor U6815 (N_6815,N_6700,N_6741);
nand U6816 (N_6816,N_6637,N_6744);
or U6817 (N_6817,N_6646,N_6700);
xnor U6818 (N_6818,N_6737,N_6698);
nand U6819 (N_6819,N_6694,N_6625);
nand U6820 (N_6820,N_6740,N_6720);
or U6821 (N_6821,N_6725,N_6728);
xnor U6822 (N_6822,N_6747,N_6653);
nor U6823 (N_6823,N_6708,N_6643);
nor U6824 (N_6824,N_6692,N_6689);
nor U6825 (N_6825,N_6732,N_6640);
nand U6826 (N_6826,N_6739,N_6700);
and U6827 (N_6827,N_6746,N_6642);
nor U6828 (N_6828,N_6639,N_6732);
nor U6829 (N_6829,N_6627,N_6701);
and U6830 (N_6830,N_6705,N_6662);
or U6831 (N_6831,N_6627,N_6649);
xnor U6832 (N_6832,N_6647,N_6644);
nand U6833 (N_6833,N_6669,N_6684);
nand U6834 (N_6834,N_6731,N_6665);
nor U6835 (N_6835,N_6715,N_6662);
or U6836 (N_6836,N_6691,N_6667);
xnor U6837 (N_6837,N_6710,N_6735);
xnor U6838 (N_6838,N_6669,N_6647);
xor U6839 (N_6839,N_6669,N_6672);
nor U6840 (N_6840,N_6727,N_6733);
and U6841 (N_6841,N_6644,N_6668);
or U6842 (N_6842,N_6632,N_6724);
xor U6843 (N_6843,N_6728,N_6713);
xnor U6844 (N_6844,N_6692,N_6740);
xor U6845 (N_6845,N_6635,N_6645);
nor U6846 (N_6846,N_6731,N_6734);
and U6847 (N_6847,N_6652,N_6724);
and U6848 (N_6848,N_6668,N_6736);
nand U6849 (N_6849,N_6728,N_6712);
xnor U6850 (N_6850,N_6730,N_6636);
or U6851 (N_6851,N_6685,N_6651);
nand U6852 (N_6852,N_6640,N_6659);
xor U6853 (N_6853,N_6672,N_6749);
nand U6854 (N_6854,N_6626,N_6698);
nor U6855 (N_6855,N_6739,N_6749);
nor U6856 (N_6856,N_6682,N_6742);
xnor U6857 (N_6857,N_6673,N_6660);
or U6858 (N_6858,N_6654,N_6680);
and U6859 (N_6859,N_6632,N_6735);
and U6860 (N_6860,N_6725,N_6689);
xor U6861 (N_6861,N_6633,N_6746);
nor U6862 (N_6862,N_6658,N_6653);
nor U6863 (N_6863,N_6688,N_6686);
nand U6864 (N_6864,N_6747,N_6652);
or U6865 (N_6865,N_6673,N_6743);
and U6866 (N_6866,N_6703,N_6679);
nand U6867 (N_6867,N_6677,N_6745);
and U6868 (N_6868,N_6699,N_6640);
nor U6869 (N_6869,N_6696,N_6705);
nand U6870 (N_6870,N_6700,N_6715);
and U6871 (N_6871,N_6631,N_6670);
xor U6872 (N_6872,N_6687,N_6703);
xor U6873 (N_6873,N_6748,N_6647);
or U6874 (N_6874,N_6706,N_6686);
or U6875 (N_6875,N_6780,N_6862);
nand U6876 (N_6876,N_6819,N_6849);
nor U6877 (N_6877,N_6798,N_6855);
and U6878 (N_6878,N_6799,N_6757);
nand U6879 (N_6879,N_6775,N_6806);
nand U6880 (N_6880,N_6751,N_6812);
and U6881 (N_6881,N_6835,N_6865);
nand U6882 (N_6882,N_6826,N_6857);
or U6883 (N_6883,N_6801,N_6829);
nand U6884 (N_6884,N_6800,N_6773);
and U6885 (N_6885,N_6866,N_6863);
and U6886 (N_6886,N_6831,N_6785);
nor U6887 (N_6887,N_6816,N_6752);
nand U6888 (N_6888,N_6838,N_6789);
xor U6889 (N_6889,N_6864,N_6815);
xnor U6890 (N_6890,N_6804,N_6759);
and U6891 (N_6891,N_6823,N_6779);
xor U6892 (N_6892,N_6784,N_6843);
and U6893 (N_6893,N_6807,N_6818);
nor U6894 (N_6894,N_6754,N_6874);
nor U6895 (N_6895,N_6782,N_6770);
and U6896 (N_6896,N_6766,N_6822);
and U6897 (N_6897,N_6837,N_6841);
nand U6898 (N_6898,N_6794,N_6796);
or U6899 (N_6899,N_6861,N_6762);
and U6900 (N_6900,N_6786,N_6845);
nor U6901 (N_6901,N_6870,N_6834);
nand U6902 (N_6902,N_6795,N_6783);
nand U6903 (N_6903,N_6790,N_6768);
and U6904 (N_6904,N_6791,N_6788);
nand U6905 (N_6905,N_6828,N_6760);
or U6906 (N_6906,N_6774,N_6776);
nor U6907 (N_6907,N_6753,N_6847);
and U6908 (N_6908,N_6873,N_6765);
and U6909 (N_6909,N_6839,N_6850);
xnor U6910 (N_6910,N_6810,N_6860);
nand U6911 (N_6911,N_6756,N_6808);
xor U6912 (N_6912,N_6858,N_6755);
and U6913 (N_6913,N_6769,N_6821);
or U6914 (N_6914,N_6761,N_6777);
xor U6915 (N_6915,N_6787,N_6851);
xor U6916 (N_6916,N_6830,N_6797);
or U6917 (N_6917,N_6805,N_6781);
and U6918 (N_6918,N_6868,N_6767);
nand U6919 (N_6919,N_6811,N_6763);
or U6920 (N_6920,N_6872,N_6871);
or U6921 (N_6921,N_6848,N_6758);
or U6922 (N_6922,N_6809,N_6844);
or U6923 (N_6923,N_6853,N_6824);
and U6924 (N_6924,N_6840,N_6836);
or U6925 (N_6925,N_6846,N_6778);
xor U6926 (N_6926,N_6750,N_6820);
xor U6927 (N_6927,N_6856,N_6817);
nand U6928 (N_6928,N_6792,N_6803);
or U6929 (N_6929,N_6814,N_6854);
and U6930 (N_6930,N_6869,N_6802);
nor U6931 (N_6931,N_6833,N_6771);
xnor U6932 (N_6932,N_6859,N_6764);
or U6933 (N_6933,N_6825,N_6827);
nor U6934 (N_6934,N_6842,N_6793);
nand U6935 (N_6935,N_6867,N_6852);
xnor U6936 (N_6936,N_6832,N_6772);
nor U6937 (N_6937,N_6813,N_6804);
and U6938 (N_6938,N_6832,N_6873);
xnor U6939 (N_6939,N_6776,N_6780);
nor U6940 (N_6940,N_6788,N_6809);
xor U6941 (N_6941,N_6809,N_6817);
and U6942 (N_6942,N_6781,N_6872);
and U6943 (N_6943,N_6829,N_6782);
or U6944 (N_6944,N_6863,N_6869);
or U6945 (N_6945,N_6867,N_6836);
or U6946 (N_6946,N_6873,N_6793);
xnor U6947 (N_6947,N_6764,N_6871);
nor U6948 (N_6948,N_6835,N_6825);
and U6949 (N_6949,N_6828,N_6761);
xnor U6950 (N_6950,N_6811,N_6769);
nand U6951 (N_6951,N_6763,N_6828);
and U6952 (N_6952,N_6856,N_6794);
nand U6953 (N_6953,N_6794,N_6844);
nor U6954 (N_6954,N_6807,N_6820);
and U6955 (N_6955,N_6870,N_6871);
or U6956 (N_6956,N_6761,N_6818);
and U6957 (N_6957,N_6751,N_6843);
and U6958 (N_6958,N_6791,N_6779);
and U6959 (N_6959,N_6800,N_6760);
xor U6960 (N_6960,N_6807,N_6829);
xnor U6961 (N_6961,N_6760,N_6789);
or U6962 (N_6962,N_6753,N_6808);
nor U6963 (N_6963,N_6844,N_6861);
and U6964 (N_6964,N_6799,N_6837);
and U6965 (N_6965,N_6840,N_6779);
xor U6966 (N_6966,N_6834,N_6821);
and U6967 (N_6967,N_6827,N_6754);
xor U6968 (N_6968,N_6808,N_6863);
xnor U6969 (N_6969,N_6810,N_6813);
and U6970 (N_6970,N_6797,N_6769);
and U6971 (N_6971,N_6784,N_6838);
nand U6972 (N_6972,N_6787,N_6828);
nand U6973 (N_6973,N_6783,N_6848);
nor U6974 (N_6974,N_6759,N_6852);
xor U6975 (N_6975,N_6764,N_6869);
xor U6976 (N_6976,N_6810,N_6807);
or U6977 (N_6977,N_6759,N_6863);
nor U6978 (N_6978,N_6798,N_6772);
nor U6979 (N_6979,N_6863,N_6799);
xor U6980 (N_6980,N_6811,N_6835);
or U6981 (N_6981,N_6867,N_6809);
and U6982 (N_6982,N_6770,N_6804);
and U6983 (N_6983,N_6778,N_6844);
xor U6984 (N_6984,N_6786,N_6789);
xnor U6985 (N_6985,N_6824,N_6863);
and U6986 (N_6986,N_6751,N_6766);
nor U6987 (N_6987,N_6786,N_6825);
xnor U6988 (N_6988,N_6815,N_6832);
nand U6989 (N_6989,N_6858,N_6850);
nor U6990 (N_6990,N_6812,N_6787);
xnor U6991 (N_6991,N_6783,N_6799);
xor U6992 (N_6992,N_6794,N_6870);
or U6993 (N_6993,N_6819,N_6769);
nand U6994 (N_6994,N_6863,N_6845);
and U6995 (N_6995,N_6787,N_6869);
or U6996 (N_6996,N_6794,N_6779);
xor U6997 (N_6997,N_6784,N_6844);
and U6998 (N_6998,N_6824,N_6770);
xnor U6999 (N_6999,N_6759,N_6822);
or U7000 (N_7000,N_6964,N_6905);
nor U7001 (N_7001,N_6919,N_6934);
nor U7002 (N_7002,N_6909,N_6961);
nand U7003 (N_7003,N_6898,N_6953);
nand U7004 (N_7004,N_6970,N_6986);
and U7005 (N_7005,N_6944,N_6904);
nand U7006 (N_7006,N_6889,N_6929);
and U7007 (N_7007,N_6960,N_6892);
nor U7008 (N_7008,N_6890,N_6937);
xor U7009 (N_7009,N_6918,N_6975);
nand U7010 (N_7010,N_6948,N_6922);
nor U7011 (N_7011,N_6875,N_6933);
xnor U7012 (N_7012,N_6893,N_6981);
or U7013 (N_7013,N_6880,N_6977);
or U7014 (N_7014,N_6997,N_6942);
nand U7015 (N_7015,N_6965,N_6967);
xnor U7016 (N_7016,N_6938,N_6923);
or U7017 (N_7017,N_6976,N_6951);
and U7018 (N_7018,N_6991,N_6989);
nor U7019 (N_7019,N_6887,N_6972);
or U7020 (N_7020,N_6932,N_6903);
nor U7021 (N_7021,N_6966,N_6882);
and U7022 (N_7022,N_6883,N_6911);
xor U7023 (N_7023,N_6982,N_6950);
xor U7024 (N_7024,N_6987,N_6902);
and U7025 (N_7025,N_6900,N_6959);
or U7026 (N_7026,N_6984,N_6928);
or U7027 (N_7027,N_6896,N_6886);
and U7028 (N_7028,N_6974,N_6962);
nor U7029 (N_7029,N_6956,N_6957);
or U7030 (N_7030,N_6978,N_6908);
and U7031 (N_7031,N_6910,N_6885);
nand U7032 (N_7032,N_6927,N_6985);
nor U7033 (N_7033,N_6931,N_6925);
and U7034 (N_7034,N_6949,N_6954);
nand U7035 (N_7035,N_6915,N_6945);
nor U7036 (N_7036,N_6879,N_6926);
xor U7037 (N_7037,N_6941,N_6878);
nand U7038 (N_7038,N_6920,N_6901);
nor U7039 (N_7039,N_6940,N_6971);
or U7040 (N_7040,N_6983,N_6958);
nor U7041 (N_7041,N_6969,N_6921);
nand U7042 (N_7042,N_6947,N_6998);
and U7043 (N_7043,N_6906,N_6877);
xor U7044 (N_7044,N_6876,N_6936);
nor U7045 (N_7045,N_6935,N_6946);
or U7046 (N_7046,N_6993,N_6907);
nand U7047 (N_7047,N_6899,N_6952);
or U7048 (N_7048,N_6930,N_6979);
or U7049 (N_7049,N_6968,N_6999);
xor U7050 (N_7050,N_6994,N_6895);
or U7051 (N_7051,N_6897,N_6939);
or U7052 (N_7052,N_6894,N_6995);
nor U7053 (N_7053,N_6881,N_6917);
or U7054 (N_7054,N_6973,N_6996);
nand U7055 (N_7055,N_6912,N_6891);
nand U7056 (N_7056,N_6884,N_6990);
or U7057 (N_7057,N_6992,N_6924);
and U7058 (N_7058,N_6963,N_6988);
and U7059 (N_7059,N_6888,N_6913);
xor U7060 (N_7060,N_6914,N_6916);
and U7061 (N_7061,N_6955,N_6980);
and U7062 (N_7062,N_6943,N_6971);
and U7063 (N_7063,N_6909,N_6988);
xor U7064 (N_7064,N_6921,N_6888);
and U7065 (N_7065,N_6875,N_6935);
nand U7066 (N_7066,N_6980,N_6938);
nor U7067 (N_7067,N_6920,N_6932);
nand U7068 (N_7068,N_6943,N_6883);
and U7069 (N_7069,N_6933,N_6894);
nand U7070 (N_7070,N_6877,N_6958);
xnor U7071 (N_7071,N_6941,N_6932);
nor U7072 (N_7072,N_6889,N_6962);
or U7073 (N_7073,N_6954,N_6948);
nand U7074 (N_7074,N_6920,N_6960);
nor U7075 (N_7075,N_6881,N_6946);
nor U7076 (N_7076,N_6938,N_6975);
or U7077 (N_7077,N_6995,N_6893);
and U7078 (N_7078,N_6972,N_6878);
nor U7079 (N_7079,N_6912,N_6928);
or U7080 (N_7080,N_6987,N_6981);
nor U7081 (N_7081,N_6956,N_6937);
and U7082 (N_7082,N_6968,N_6894);
xnor U7083 (N_7083,N_6891,N_6971);
nor U7084 (N_7084,N_6919,N_6968);
and U7085 (N_7085,N_6947,N_6914);
xnor U7086 (N_7086,N_6956,N_6877);
nor U7087 (N_7087,N_6892,N_6954);
nand U7088 (N_7088,N_6951,N_6877);
and U7089 (N_7089,N_6881,N_6936);
xnor U7090 (N_7090,N_6939,N_6983);
or U7091 (N_7091,N_6992,N_6895);
or U7092 (N_7092,N_6882,N_6970);
nor U7093 (N_7093,N_6960,N_6925);
and U7094 (N_7094,N_6931,N_6895);
and U7095 (N_7095,N_6913,N_6980);
and U7096 (N_7096,N_6924,N_6919);
nand U7097 (N_7097,N_6953,N_6934);
or U7098 (N_7098,N_6965,N_6897);
and U7099 (N_7099,N_6960,N_6957);
and U7100 (N_7100,N_6978,N_6957);
nor U7101 (N_7101,N_6911,N_6986);
and U7102 (N_7102,N_6976,N_6888);
nand U7103 (N_7103,N_6983,N_6954);
nor U7104 (N_7104,N_6966,N_6881);
nor U7105 (N_7105,N_6944,N_6999);
nor U7106 (N_7106,N_6996,N_6941);
and U7107 (N_7107,N_6880,N_6922);
and U7108 (N_7108,N_6995,N_6957);
xnor U7109 (N_7109,N_6981,N_6886);
xnor U7110 (N_7110,N_6971,N_6875);
and U7111 (N_7111,N_6909,N_6962);
nor U7112 (N_7112,N_6919,N_6935);
nand U7113 (N_7113,N_6946,N_6904);
or U7114 (N_7114,N_6955,N_6964);
nand U7115 (N_7115,N_6916,N_6907);
nand U7116 (N_7116,N_6977,N_6961);
nor U7117 (N_7117,N_6932,N_6969);
and U7118 (N_7118,N_6989,N_6930);
nor U7119 (N_7119,N_6927,N_6914);
xor U7120 (N_7120,N_6875,N_6892);
nand U7121 (N_7121,N_6984,N_6951);
xor U7122 (N_7122,N_6989,N_6920);
nand U7123 (N_7123,N_6973,N_6910);
nor U7124 (N_7124,N_6960,N_6947);
xor U7125 (N_7125,N_7096,N_7119);
nor U7126 (N_7126,N_7006,N_7076);
or U7127 (N_7127,N_7104,N_7013);
nand U7128 (N_7128,N_7075,N_7063);
or U7129 (N_7129,N_7022,N_7087);
nor U7130 (N_7130,N_7037,N_7035);
and U7131 (N_7131,N_7109,N_7027);
nor U7132 (N_7132,N_7054,N_7030);
or U7133 (N_7133,N_7080,N_7114);
or U7134 (N_7134,N_7017,N_7029);
xnor U7135 (N_7135,N_7001,N_7045);
nand U7136 (N_7136,N_7051,N_7020);
nor U7137 (N_7137,N_7118,N_7071);
nand U7138 (N_7138,N_7101,N_7012);
nor U7139 (N_7139,N_7002,N_7003);
or U7140 (N_7140,N_7000,N_7064);
nor U7141 (N_7141,N_7015,N_7117);
or U7142 (N_7142,N_7116,N_7073);
nor U7143 (N_7143,N_7018,N_7039);
nand U7144 (N_7144,N_7090,N_7122);
xnor U7145 (N_7145,N_7004,N_7112);
or U7146 (N_7146,N_7011,N_7049);
and U7147 (N_7147,N_7010,N_7047);
or U7148 (N_7148,N_7016,N_7069);
nand U7149 (N_7149,N_7083,N_7121);
nand U7150 (N_7150,N_7065,N_7105);
nor U7151 (N_7151,N_7024,N_7048);
nand U7152 (N_7152,N_7021,N_7056);
and U7153 (N_7153,N_7032,N_7058);
and U7154 (N_7154,N_7115,N_7052);
nor U7155 (N_7155,N_7113,N_7097);
or U7156 (N_7156,N_7060,N_7120);
nor U7157 (N_7157,N_7086,N_7055);
and U7158 (N_7158,N_7005,N_7103);
nand U7159 (N_7159,N_7079,N_7014);
nor U7160 (N_7160,N_7007,N_7100);
xnor U7161 (N_7161,N_7070,N_7106);
xnor U7162 (N_7162,N_7094,N_7053);
nor U7163 (N_7163,N_7091,N_7046);
and U7164 (N_7164,N_7059,N_7062);
nand U7165 (N_7165,N_7043,N_7033);
nand U7166 (N_7166,N_7088,N_7040);
or U7167 (N_7167,N_7031,N_7057);
nand U7168 (N_7168,N_7082,N_7107);
and U7169 (N_7169,N_7068,N_7095);
xnor U7170 (N_7170,N_7028,N_7081);
nor U7171 (N_7171,N_7077,N_7041);
and U7172 (N_7172,N_7023,N_7061);
xnor U7173 (N_7173,N_7072,N_7124);
nand U7174 (N_7174,N_7050,N_7110);
xnor U7175 (N_7175,N_7019,N_7098);
nand U7176 (N_7176,N_7008,N_7042);
or U7177 (N_7177,N_7026,N_7102);
nand U7178 (N_7178,N_7111,N_7074);
nand U7179 (N_7179,N_7085,N_7066);
or U7180 (N_7180,N_7099,N_7089);
and U7181 (N_7181,N_7067,N_7038);
nor U7182 (N_7182,N_7009,N_7084);
nor U7183 (N_7183,N_7036,N_7034);
or U7184 (N_7184,N_7044,N_7123);
nand U7185 (N_7185,N_7093,N_7078);
or U7186 (N_7186,N_7092,N_7025);
nor U7187 (N_7187,N_7108,N_7102);
nor U7188 (N_7188,N_7079,N_7076);
nor U7189 (N_7189,N_7111,N_7058);
xor U7190 (N_7190,N_7082,N_7015);
nand U7191 (N_7191,N_7115,N_7062);
xnor U7192 (N_7192,N_7050,N_7053);
or U7193 (N_7193,N_7077,N_7092);
and U7194 (N_7194,N_7015,N_7088);
nor U7195 (N_7195,N_7082,N_7030);
nand U7196 (N_7196,N_7038,N_7044);
xor U7197 (N_7197,N_7055,N_7068);
nand U7198 (N_7198,N_7086,N_7064);
or U7199 (N_7199,N_7030,N_7046);
or U7200 (N_7200,N_7043,N_7026);
nor U7201 (N_7201,N_7110,N_7025);
nor U7202 (N_7202,N_7119,N_7020);
and U7203 (N_7203,N_7099,N_7025);
nor U7204 (N_7204,N_7051,N_7032);
or U7205 (N_7205,N_7104,N_7040);
or U7206 (N_7206,N_7119,N_7077);
or U7207 (N_7207,N_7072,N_7019);
and U7208 (N_7208,N_7113,N_7047);
xor U7209 (N_7209,N_7075,N_7034);
nand U7210 (N_7210,N_7040,N_7046);
or U7211 (N_7211,N_7116,N_7076);
nand U7212 (N_7212,N_7105,N_7044);
and U7213 (N_7213,N_7024,N_7098);
nor U7214 (N_7214,N_7042,N_7106);
xnor U7215 (N_7215,N_7016,N_7032);
xnor U7216 (N_7216,N_7045,N_7069);
xnor U7217 (N_7217,N_7051,N_7101);
and U7218 (N_7218,N_7076,N_7070);
xnor U7219 (N_7219,N_7007,N_7099);
nand U7220 (N_7220,N_7052,N_7117);
xor U7221 (N_7221,N_7049,N_7090);
nand U7222 (N_7222,N_7108,N_7035);
xnor U7223 (N_7223,N_7115,N_7031);
nand U7224 (N_7224,N_7017,N_7063);
nand U7225 (N_7225,N_7038,N_7028);
nor U7226 (N_7226,N_7039,N_7001);
nand U7227 (N_7227,N_7056,N_7009);
nand U7228 (N_7228,N_7024,N_7114);
nand U7229 (N_7229,N_7081,N_7005);
or U7230 (N_7230,N_7103,N_7030);
nand U7231 (N_7231,N_7000,N_7047);
nand U7232 (N_7232,N_7043,N_7118);
and U7233 (N_7233,N_7050,N_7124);
xnor U7234 (N_7234,N_7073,N_7113);
nand U7235 (N_7235,N_7016,N_7065);
and U7236 (N_7236,N_7115,N_7036);
nand U7237 (N_7237,N_7025,N_7087);
nand U7238 (N_7238,N_7035,N_7014);
or U7239 (N_7239,N_7094,N_7047);
or U7240 (N_7240,N_7042,N_7082);
nand U7241 (N_7241,N_7083,N_7118);
nor U7242 (N_7242,N_7106,N_7047);
or U7243 (N_7243,N_7006,N_7111);
or U7244 (N_7244,N_7061,N_7063);
or U7245 (N_7245,N_7079,N_7098);
xnor U7246 (N_7246,N_7055,N_7045);
nand U7247 (N_7247,N_7015,N_7116);
or U7248 (N_7248,N_7092,N_7039);
xor U7249 (N_7249,N_7012,N_7039);
and U7250 (N_7250,N_7223,N_7202);
or U7251 (N_7251,N_7172,N_7249);
nor U7252 (N_7252,N_7136,N_7160);
and U7253 (N_7253,N_7187,N_7192);
or U7254 (N_7254,N_7178,N_7216);
xnor U7255 (N_7255,N_7218,N_7132);
nor U7256 (N_7256,N_7135,N_7139);
xnor U7257 (N_7257,N_7155,N_7185);
nor U7258 (N_7258,N_7222,N_7213);
or U7259 (N_7259,N_7149,N_7151);
nand U7260 (N_7260,N_7201,N_7181);
or U7261 (N_7261,N_7145,N_7128);
nand U7262 (N_7262,N_7130,N_7236);
nor U7263 (N_7263,N_7174,N_7229);
nor U7264 (N_7264,N_7239,N_7150);
nand U7265 (N_7265,N_7211,N_7180);
and U7266 (N_7266,N_7241,N_7183);
nor U7267 (N_7267,N_7126,N_7228);
nor U7268 (N_7268,N_7246,N_7153);
or U7269 (N_7269,N_7129,N_7200);
and U7270 (N_7270,N_7157,N_7203);
nor U7271 (N_7271,N_7186,N_7167);
or U7272 (N_7272,N_7163,N_7170);
or U7273 (N_7273,N_7152,N_7169);
nand U7274 (N_7274,N_7162,N_7217);
xnor U7275 (N_7275,N_7147,N_7137);
or U7276 (N_7276,N_7207,N_7194);
or U7277 (N_7277,N_7168,N_7204);
or U7278 (N_7278,N_7134,N_7219);
nand U7279 (N_7279,N_7237,N_7148);
or U7280 (N_7280,N_7189,N_7238);
nand U7281 (N_7281,N_7154,N_7247);
xnor U7282 (N_7282,N_7221,N_7208);
xor U7283 (N_7283,N_7240,N_7242);
nor U7284 (N_7284,N_7171,N_7220);
or U7285 (N_7285,N_7215,N_7214);
nand U7286 (N_7286,N_7175,N_7212);
nand U7287 (N_7287,N_7165,N_7144);
nand U7288 (N_7288,N_7210,N_7156);
nor U7289 (N_7289,N_7190,N_7182);
xor U7290 (N_7290,N_7232,N_7188);
and U7291 (N_7291,N_7177,N_7140);
nand U7292 (N_7292,N_7191,N_7127);
xnor U7293 (N_7293,N_7225,N_7231);
xor U7294 (N_7294,N_7196,N_7206);
or U7295 (N_7295,N_7227,N_7209);
xor U7296 (N_7296,N_7248,N_7234);
and U7297 (N_7297,N_7176,N_7141);
xor U7298 (N_7298,N_7244,N_7138);
nand U7299 (N_7299,N_7158,N_7131);
and U7300 (N_7300,N_7193,N_7226);
nor U7301 (N_7301,N_7166,N_7146);
and U7302 (N_7302,N_7224,N_7161);
nor U7303 (N_7303,N_7184,N_7133);
nor U7304 (N_7304,N_7230,N_7179);
nor U7305 (N_7305,N_7125,N_7199);
xor U7306 (N_7306,N_7195,N_7205);
and U7307 (N_7307,N_7243,N_7233);
or U7308 (N_7308,N_7235,N_7142);
or U7309 (N_7309,N_7159,N_7173);
nand U7310 (N_7310,N_7245,N_7164);
nand U7311 (N_7311,N_7198,N_7143);
nand U7312 (N_7312,N_7197,N_7181);
nand U7313 (N_7313,N_7148,N_7192);
nand U7314 (N_7314,N_7167,N_7129);
nand U7315 (N_7315,N_7218,N_7213);
and U7316 (N_7316,N_7211,N_7154);
or U7317 (N_7317,N_7181,N_7174);
nor U7318 (N_7318,N_7241,N_7167);
nor U7319 (N_7319,N_7168,N_7213);
nand U7320 (N_7320,N_7152,N_7173);
and U7321 (N_7321,N_7138,N_7140);
xor U7322 (N_7322,N_7140,N_7246);
or U7323 (N_7323,N_7213,N_7151);
nand U7324 (N_7324,N_7125,N_7161);
xnor U7325 (N_7325,N_7218,N_7136);
xor U7326 (N_7326,N_7159,N_7186);
xor U7327 (N_7327,N_7238,N_7185);
nand U7328 (N_7328,N_7224,N_7180);
or U7329 (N_7329,N_7207,N_7225);
or U7330 (N_7330,N_7128,N_7211);
nor U7331 (N_7331,N_7233,N_7191);
xor U7332 (N_7332,N_7164,N_7210);
and U7333 (N_7333,N_7167,N_7222);
xor U7334 (N_7334,N_7174,N_7140);
xnor U7335 (N_7335,N_7157,N_7168);
and U7336 (N_7336,N_7191,N_7135);
and U7337 (N_7337,N_7205,N_7137);
xnor U7338 (N_7338,N_7167,N_7220);
nor U7339 (N_7339,N_7195,N_7222);
or U7340 (N_7340,N_7175,N_7226);
nand U7341 (N_7341,N_7176,N_7130);
or U7342 (N_7342,N_7191,N_7164);
or U7343 (N_7343,N_7177,N_7184);
or U7344 (N_7344,N_7169,N_7175);
nand U7345 (N_7345,N_7131,N_7227);
or U7346 (N_7346,N_7236,N_7235);
and U7347 (N_7347,N_7168,N_7165);
nor U7348 (N_7348,N_7150,N_7173);
and U7349 (N_7349,N_7229,N_7128);
or U7350 (N_7350,N_7173,N_7180);
nand U7351 (N_7351,N_7219,N_7152);
nand U7352 (N_7352,N_7159,N_7217);
or U7353 (N_7353,N_7134,N_7236);
xor U7354 (N_7354,N_7149,N_7190);
or U7355 (N_7355,N_7215,N_7176);
nand U7356 (N_7356,N_7146,N_7232);
nor U7357 (N_7357,N_7213,N_7237);
nand U7358 (N_7358,N_7146,N_7141);
and U7359 (N_7359,N_7242,N_7221);
nor U7360 (N_7360,N_7175,N_7216);
and U7361 (N_7361,N_7163,N_7187);
nand U7362 (N_7362,N_7243,N_7159);
and U7363 (N_7363,N_7234,N_7219);
nand U7364 (N_7364,N_7218,N_7179);
nand U7365 (N_7365,N_7244,N_7127);
nor U7366 (N_7366,N_7143,N_7189);
nor U7367 (N_7367,N_7149,N_7247);
or U7368 (N_7368,N_7225,N_7203);
nand U7369 (N_7369,N_7165,N_7206);
and U7370 (N_7370,N_7198,N_7185);
nand U7371 (N_7371,N_7246,N_7160);
nand U7372 (N_7372,N_7191,N_7210);
and U7373 (N_7373,N_7244,N_7165);
and U7374 (N_7374,N_7196,N_7242);
nand U7375 (N_7375,N_7317,N_7316);
nand U7376 (N_7376,N_7330,N_7318);
nand U7377 (N_7377,N_7351,N_7344);
nand U7378 (N_7378,N_7296,N_7367);
and U7379 (N_7379,N_7372,N_7329);
or U7380 (N_7380,N_7328,N_7341);
and U7381 (N_7381,N_7289,N_7324);
xnor U7382 (N_7382,N_7280,N_7307);
xnor U7383 (N_7383,N_7274,N_7327);
xor U7384 (N_7384,N_7253,N_7331);
nor U7385 (N_7385,N_7265,N_7254);
and U7386 (N_7386,N_7276,N_7271);
nor U7387 (N_7387,N_7360,N_7359);
and U7388 (N_7388,N_7295,N_7298);
nor U7389 (N_7389,N_7277,N_7332);
xnor U7390 (N_7390,N_7285,N_7251);
and U7391 (N_7391,N_7353,N_7349);
or U7392 (N_7392,N_7370,N_7270);
and U7393 (N_7393,N_7363,N_7259);
nor U7394 (N_7394,N_7357,N_7369);
nor U7395 (N_7395,N_7304,N_7262);
nand U7396 (N_7396,N_7313,N_7288);
or U7397 (N_7397,N_7373,N_7263);
nand U7398 (N_7398,N_7279,N_7340);
or U7399 (N_7399,N_7286,N_7252);
or U7400 (N_7400,N_7362,N_7343);
or U7401 (N_7401,N_7365,N_7339);
nand U7402 (N_7402,N_7358,N_7314);
or U7403 (N_7403,N_7257,N_7334);
nor U7404 (N_7404,N_7333,N_7258);
nand U7405 (N_7405,N_7354,N_7311);
nand U7406 (N_7406,N_7306,N_7335);
nor U7407 (N_7407,N_7320,N_7275);
nand U7408 (N_7408,N_7267,N_7273);
nor U7409 (N_7409,N_7347,N_7303);
and U7410 (N_7410,N_7282,N_7250);
xnor U7411 (N_7411,N_7325,N_7348);
xnor U7412 (N_7412,N_7301,N_7299);
and U7413 (N_7413,N_7319,N_7350);
or U7414 (N_7414,N_7266,N_7291);
nor U7415 (N_7415,N_7256,N_7315);
or U7416 (N_7416,N_7310,N_7290);
nor U7417 (N_7417,N_7326,N_7366);
nand U7418 (N_7418,N_7305,N_7268);
and U7419 (N_7419,N_7281,N_7352);
and U7420 (N_7420,N_7355,N_7342);
xnor U7421 (N_7421,N_7361,N_7338);
nand U7422 (N_7422,N_7272,N_7374);
and U7423 (N_7423,N_7297,N_7278);
nand U7424 (N_7424,N_7309,N_7364);
xor U7425 (N_7425,N_7323,N_7302);
nor U7426 (N_7426,N_7321,N_7346);
nand U7427 (N_7427,N_7264,N_7261);
nor U7428 (N_7428,N_7287,N_7292);
or U7429 (N_7429,N_7293,N_7337);
nor U7430 (N_7430,N_7284,N_7260);
or U7431 (N_7431,N_7322,N_7308);
nand U7432 (N_7432,N_7356,N_7283);
nor U7433 (N_7433,N_7294,N_7312);
nor U7434 (N_7434,N_7368,N_7371);
nor U7435 (N_7435,N_7336,N_7269);
and U7436 (N_7436,N_7345,N_7255);
and U7437 (N_7437,N_7300,N_7362);
or U7438 (N_7438,N_7257,N_7330);
nand U7439 (N_7439,N_7319,N_7293);
xor U7440 (N_7440,N_7321,N_7261);
nor U7441 (N_7441,N_7261,N_7257);
or U7442 (N_7442,N_7289,N_7341);
or U7443 (N_7443,N_7318,N_7273);
xor U7444 (N_7444,N_7250,N_7325);
and U7445 (N_7445,N_7314,N_7287);
nand U7446 (N_7446,N_7324,N_7348);
xnor U7447 (N_7447,N_7337,N_7330);
nand U7448 (N_7448,N_7317,N_7299);
xnor U7449 (N_7449,N_7303,N_7371);
nor U7450 (N_7450,N_7285,N_7318);
nor U7451 (N_7451,N_7267,N_7285);
and U7452 (N_7452,N_7252,N_7354);
nand U7453 (N_7453,N_7262,N_7299);
or U7454 (N_7454,N_7299,N_7370);
nor U7455 (N_7455,N_7348,N_7309);
nand U7456 (N_7456,N_7373,N_7303);
nor U7457 (N_7457,N_7359,N_7365);
nor U7458 (N_7458,N_7298,N_7310);
and U7459 (N_7459,N_7285,N_7337);
xor U7460 (N_7460,N_7261,N_7295);
xnor U7461 (N_7461,N_7317,N_7351);
xor U7462 (N_7462,N_7365,N_7355);
and U7463 (N_7463,N_7373,N_7340);
or U7464 (N_7464,N_7307,N_7330);
and U7465 (N_7465,N_7340,N_7339);
nor U7466 (N_7466,N_7274,N_7278);
nand U7467 (N_7467,N_7373,N_7356);
xor U7468 (N_7468,N_7294,N_7360);
xor U7469 (N_7469,N_7258,N_7358);
nor U7470 (N_7470,N_7374,N_7305);
nor U7471 (N_7471,N_7257,N_7269);
or U7472 (N_7472,N_7309,N_7363);
or U7473 (N_7473,N_7277,N_7266);
and U7474 (N_7474,N_7280,N_7332);
nor U7475 (N_7475,N_7332,N_7369);
and U7476 (N_7476,N_7339,N_7271);
or U7477 (N_7477,N_7327,N_7363);
and U7478 (N_7478,N_7363,N_7293);
xnor U7479 (N_7479,N_7331,N_7260);
or U7480 (N_7480,N_7306,N_7330);
xnor U7481 (N_7481,N_7273,N_7337);
xnor U7482 (N_7482,N_7348,N_7296);
nor U7483 (N_7483,N_7332,N_7325);
nor U7484 (N_7484,N_7280,N_7283);
or U7485 (N_7485,N_7337,N_7290);
nand U7486 (N_7486,N_7354,N_7277);
nor U7487 (N_7487,N_7313,N_7251);
xnor U7488 (N_7488,N_7270,N_7291);
and U7489 (N_7489,N_7356,N_7269);
and U7490 (N_7490,N_7344,N_7273);
xnor U7491 (N_7491,N_7299,N_7374);
xnor U7492 (N_7492,N_7293,N_7334);
nor U7493 (N_7493,N_7298,N_7313);
nor U7494 (N_7494,N_7351,N_7361);
and U7495 (N_7495,N_7359,N_7295);
and U7496 (N_7496,N_7314,N_7300);
or U7497 (N_7497,N_7325,N_7290);
nor U7498 (N_7498,N_7312,N_7326);
or U7499 (N_7499,N_7303,N_7336);
or U7500 (N_7500,N_7392,N_7427);
nand U7501 (N_7501,N_7485,N_7375);
xor U7502 (N_7502,N_7439,N_7428);
nor U7503 (N_7503,N_7406,N_7400);
nand U7504 (N_7504,N_7432,N_7426);
nand U7505 (N_7505,N_7493,N_7407);
and U7506 (N_7506,N_7433,N_7408);
and U7507 (N_7507,N_7453,N_7489);
nor U7508 (N_7508,N_7378,N_7390);
and U7509 (N_7509,N_7402,N_7454);
xnor U7510 (N_7510,N_7481,N_7435);
and U7511 (N_7511,N_7380,N_7470);
or U7512 (N_7512,N_7465,N_7376);
nand U7513 (N_7513,N_7383,N_7421);
nand U7514 (N_7514,N_7456,N_7498);
nand U7515 (N_7515,N_7450,N_7420);
and U7516 (N_7516,N_7473,N_7377);
and U7517 (N_7517,N_7394,N_7417);
and U7518 (N_7518,N_7446,N_7438);
and U7519 (N_7519,N_7440,N_7466);
and U7520 (N_7520,N_7412,N_7452);
and U7521 (N_7521,N_7411,N_7398);
and U7522 (N_7522,N_7449,N_7445);
or U7523 (N_7523,N_7483,N_7499);
or U7524 (N_7524,N_7419,N_7387);
xnor U7525 (N_7525,N_7399,N_7415);
xnor U7526 (N_7526,N_7441,N_7388);
nor U7527 (N_7527,N_7429,N_7469);
or U7528 (N_7528,N_7424,N_7444);
nor U7529 (N_7529,N_7389,N_7397);
or U7530 (N_7530,N_7448,N_7474);
nand U7531 (N_7531,N_7443,N_7395);
xnor U7532 (N_7532,N_7478,N_7488);
or U7533 (N_7533,N_7492,N_7468);
nor U7534 (N_7534,N_7487,N_7458);
nor U7535 (N_7535,N_7455,N_7416);
nor U7536 (N_7536,N_7471,N_7437);
nor U7537 (N_7537,N_7490,N_7430);
nand U7538 (N_7538,N_7436,N_7496);
nand U7539 (N_7539,N_7425,N_7404);
and U7540 (N_7540,N_7393,N_7447);
nand U7541 (N_7541,N_7401,N_7482);
or U7542 (N_7542,N_7476,N_7477);
nand U7543 (N_7543,N_7391,N_7413);
nor U7544 (N_7544,N_7414,N_7472);
nor U7545 (N_7545,N_7451,N_7434);
nand U7546 (N_7546,N_7463,N_7467);
or U7547 (N_7547,N_7418,N_7480);
and U7548 (N_7548,N_7459,N_7486);
and U7549 (N_7549,N_7382,N_7461);
xnor U7550 (N_7550,N_7384,N_7405);
xnor U7551 (N_7551,N_7423,N_7379);
nor U7552 (N_7552,N_7460,N_7484);
nand U7553 (N_7553,N_7409,N_7457);
or U7554 (N_7554,N_7497,N_7464);
xor U7555 (N_7555,N_7386,N_7381);
nand U7556 (N_7556,N_7475,N_7396);
or U7557 (N_7557,N_7495,N_7385);
and U7558 (N_7558,N_7479,N_7422);
xnor U7559 (N_7559,N_7431,N_7491);
nand U7560 (N_7560,N_7410,N_7403);
nand U7561 (N_7561,N_7462,N_7494);
and U7562 (N_7562,N_7442,N_7376);
or U7563 (N_7563,N_7383,N_7442);
nor U7564 (N_7564,N_7496,N_7415);
nand U7565 (N_7565,N_7488,N_7467);
and U7566 (N_7566,N_7412,N_7386);
xnor U7567 (N_7567,N_7393,N_7376);
nand U7568 (N_7568,N_7485,N_7426);
nor U7569 (N_7569,N_7404,N_7388);
nand U7570 (N_7570,N_7388,N_7482);
or U7571 (N_7571,N_7427,N_7486);
and U7572 (N_7572,N_7402,N_7420);
xor U7573 (N_7573,N_7380,N_7442);
nand U7574 (N_7574,N_7462,N_7382);
or U7575 (N_7575,N_7484,N_7393);
nand U7576 (N_7576,N_7425,N_7445);
xor U7577 (N_7577,N_7402,N_7452);
xnor U7578 (N_7578,N_7427,N_7462);
nand U7579 (N_7579,N_7496,N_7421);
and U7580 (N_7580,N_7452,N_7464);
or U7581 (N_7581,N_7423,N_7450);
xnor U7582 (N_7582,N_7401,N_7408);
nand U7583 (N_7583,N_7388,N_7432);
and U7584 (N_7584,N_7499,N_7380);
and U7585 (N_7585,N_7425,N_7417);
nor U7586 (N_7586,N_7381,N_7485);
and U7587 (N_7587,N_7466,N_7452);
and U7588 (N_7588,N_7438,N_7426);
or U7589 (N_7589,N_7453,N_7397);
and U7590 (N_7590,N_7401,N_7497);
nand U7591 (N_7591,N_7435,N_7476);
nand U7592 (N_7592,N_7400,N_7393);
nor U7593 (N_7593,N_7382,N_7442);
xor U7594 (N_7594,N_7426,N_7428);
and U7595 (N_7595,N_7455,N_7476);
nor U7596 (N_7596,N_7459,N_7494);
xnor U7597 (N_7597,N_7436,N_7429);
and U7598 (N_7598,N_7381,N_7429);
nand U7599 (N_7599,N_7429,N_7437);
and U7600 (N_7600,N_7405,N_7421);
xnor U7601 (N_7601,N_7463,N_7461);
nand U7602 (N_7602,N_7493,N_7395);
and U7603 (N_7603,N_7429,N_7391);
nand U7604 (N_7604,N_7432,N_7419);
or U7605 (N_7605,N_7442,N_7390);
nor U7606 (N_7606,N_7376,N_7463);
nor U7607 (N_7607,N_7460,N_7445);
nand U7608 (N_7608,N_7404,N_7417);
or U7609 (N_7609,N_7408,N_7452);
and U7610 (N_7610,N_7472,N_7408);
and U7611 (N_7611,N_7390,N_7414);
or U7612 (N_7612,N_7446,N_7403);
nand U7613 (N_7613,N_7467,N_7399);
or U7614 (N_7614,N_7470,N_7403);
or U7615 (N_7615,N_7475,N_7423);
xor U7616 (N_7616,N_7479,N_7443);
xor U7617 (N_7617,N_7407,N_7389);
nor U7618 (N_7618,N_7482,N_7419);
nor U7619 (N_7619,N_7440,N_7378);
nor U7620 (N_7620,N_7458,N_7399);
nand U7621 (N_7621,N_7420,N_7380);
and U7622 (N_7622,N_7397,N_7494);
nand U7623 (N_7623,N_7449,N_7497);
nand U7624 (N_7624,N_7469,N_7440);
and U7625 (N_7625,N_7506,N_7511);
nand U7626 (N_7626,N_7566,N_7526);
nand U7627 (N_7627,N_7572,N_7603);
nand U7628 (N_7628,N_7597,N_7606);
nand U7629 (N_7629,N_7589,N_7599);
xor U7630 (N_7630,N_7580,N_7620);
nor U7631 (N_7631,N_7544,N_7536);
nor U7632 (N_7632,N_7554,N_7604);
nor U7633 (N_7633,N_7613,N_7583);
nor U7634 (N_7634,N_7516,N_7518);
xnor U7635 (N_7635,N_7533,N_7517);
or U7636 (N_7636,N_7507,N_7615);
nor U7637 (N_7637,N_7548,N_7556);
or U7638 (N_7638,N_7553,N_7596);
nor U7639 (N_7639,N_7546,N_7577);
nor U7640 (N_7640,N_7579,N_7564);
and U7641 (N_7641,N_7514,N_7528);
xnor U7642 (N_7642,N_7614,N_7617);
and U7643 (N_7643,N_7503,N_7542);
and U7644 (N_7644,N_7622,N_7581);
nor U7645 (N_7645,N_7539,N_7505);
nand U7646 (N_7646,N_7521,N_7569);
or U7647 (N_7647,N_7594,N_7537);
xor U7648 (N_7648,N_7508,N_7515);
nand U7649 (N_7649,N_7501,N_7570);
and U7650 (N_7650,N_7559,N_7519);
xnor U7651 (N_7651,N_7523,N_7562);
nand U7652 (N_7652,N_7587,N_7551);
nand U7653 (N_7653,N_7522,N_7592);
and U7654 (N_7654,N_7605,N_7561);
xor U7655 (N_7655,N_7575,N_7545);
or U7656 (N_7656,N_7567,N_7621);
nand U7657 (N_7657,N_7563,N_7565);
and U7658 (N_7658,N_7568,N_7532);
and U7659 (N_7659,N_7550,N_7549);
xnor U7660 (N_7660,N_7531,N_7552);
and U7661 (N_7661,N_7590,N_7608);
xnor U7662 (N_7662,N_7601,N_7595);
nand U7663 (N_7663,N_7512,N_7607);
nand U7664 (N_7664,N_7525,N_7540);
xor U7665 (N_7665,N_7612,N_7547);
xor U7666 (N_7666,N_7513,N_7591);
xnor U7667 (N_7667,N_7611,N_7585);
nor U7668 (N_7668,N_7593,N_7527);
xor U7669 (N_7669,N_7584,N_7610);
nor U7670 (N_7670,N_7578,N_7520);
nor U7671 (N_7671,N_7588,N_7602);
and U7672 (N_7672,N_7609,N_7598);
nand U7673 (N_7673,N_7619,N_7616);
or U7674 (N_7674,N_7538,N_7557);
and U7675 (N_7675,N_7573,N_7504);
or U7676 (N_7676,N_7534,N_7535);
nand U7677 (N_7677,N_7574,N_7586);
nand U7678 (N_7678,N_7560,N_7582);
nor U7679 (N_7679,N_7600,N_7543);
or U7680 (N_7680,N_7500,N_7502);
and U7681 (N_7681,N_7624,N_7618);
and U7682 (N_7682,N_7558,N_7576);
and U7683 (N_7683,N_7571,N_7541);
or U7684 (N_7684,N_7529,N_7510);
nor U7685 (N_7685,N_7530,N_7623);
or U7686 (N_7686,N_7524,N_7555);
and U7687 (N_7687,N_7509,N_7614);
and U7688 (N_7688,N_7592,N_7535);
and U7689 (N_7689,N_7523,N_7587);
xnor U7690 (N_7690,N_7572,N_7511);
or U7691 (N_7691,N_7504,N_7574);
or U7692 (N_7692,N_7613,N_7615);
xor U7693 (N_7693,N_7517,N_7570);
nor U7694 (N_7694,N_7599,N_7556);
nand U7695 (N_7695,N_7549,N_7506);
xor U7696 (N_7696,N_7565,N_7501);
or U7697 (N_7697,N_7538,N_7544);
and U7698 (N_7698,N_7558,N_7573);
or U7699 (N_7699,N_7551,N_7603);
nor U7700 (N_7700,N_7576,N_7589);
nor U7701 (N_7701,N_7573,N_7545);
xor U7702 (N_7702,N_7525,N_7516);
nand U7703 (N_7703,N_7503,N_7521);
nand U7704 (N_7704,N_7532,N_7541);
xor U7705 (N_7705,N_7521,N_7528);
nand U7706 (N_7706,N_7594,N_7565);
and U7707 (N_7707,N_7503,N_7507);
xor U7708 (N_7708,N_7580,N_7589);
or U7709 (N_7709,N_7576,N_7546);
and U7710 (N_7710,N_7575,N_7548);
nand U7711 (N_7711,N_7557,N_7572);
xnor U7712 (N_7712,N_7535,N_7516);
nor U7713 (N_7713,N_7527,N_7575);
nor U7714 (N_7714,N_7532,N_7593);
and U7715 (N_7715,N_7578,N_7613);
and U7716 (N_7716,N_7508,N_7537);
and U7717 (N_7717,N_7556,N_7613);
or U7718 (N_7718,N_7519,N_7523);
nand U7719 (N_7719,N_7621,N_7569);
or U7720 (N_7720,N_7608,N_7588);
nor U7721 (N_7721,N_7521,N_7561);
nand U7722 (N_7722,N_7501,N_7574);
xor U7723 (N_7723,N_7622,N_7568);
nand U7724 (N_7724,N_7577,N_7616);
or U7725 (N_7725,N_7613,N_7589);
nor U7726 (N_7726,N_7546,N_7561);
nand U7727 (N_7727,N_7620,N_7548);
nand U7728 (N_7728,N_7609,N_7516);
and U7729 (N_7729,N_7607,N_7613);
or U7730 (N_7730,N_7597,N_7574);
or U7731 (N_7731,N_7534,N_7608);
or U7732 (N_7732,N_7616,N_7557);
xor U7733 (N_7733,N_7525,N_7583);
nor U7734 (N_7734,N_7501,N_7606);
nor U7735 (N_7735,N_7601,N_7532);
nor U7736 (N_7736,N_7552,N_7506);
nor U7737 (N_7737,N_7541,N_7511);
nor U7738 (N_7738,N_7529,N_7623);
nor U7739 (N_7739,N_7534,N_7553);
xor U7740 (N_7740,N_7576,N_7531);
or U7741 (N_7741,N_7552,N_7585);
nor U7742 (N_7742,N_7507,N_7623);
nand U7743 (N_7743,N_7618,N_7507);
or U7744 (N_7744,N_7534,N_7549);
nand U7745 (N_7745,N_7503,N_7608);
and U7746 (N_7746,N_7623,N_7506);
xor U7747 (N_7747,N_7604,N_7545);
nand U7748 (N_7748,N_7609,N_7617);
nand U7749 (N_7749,N_7525,N_7504);
and U7750 (N_7750,N_7647,N_7733);
nor U7751 (N_7751,N_7717,N_7683);
xor U7752 (N_7752,N_7703,N_7666);
nor U7753 (N_7753,N_7704,N_7698);
xor U7754 (N_7754,N_7634,N_7650);
nand U7755 (N_7755,N_7652,N_7741);
or U7756 (N_7756,N_7715,N_7731);
nand U7757 (N_7757,N_7735,N_7665);
or U7758 (N_7758,N_7658,N_7630);
or U7759 (N_7759,N_7719,N_7727);
or U7760 (N_7760,N_7669,N_7638);
nand U7761 (N_7761,N_7695,N_7685);
nand U7762 (N_7762,N_7716,N_7680);
or U7763 (N_7763,N_7691,N_7649);
and U7764 (N_7764,N_7625,N_7681);
and U7765 (N_7765,N_7674,N_7646);
or U7766 (N_7766,N_7642,N_7654);
and U7767 (N_7767,N_7739,N_7742);
nand U7768 (N_7768,N_7690,N_7656);
xnor U7769 (N_7769,N_7626,N_7648);
or U7770 (N_7770,N_7740,N_7701);
nor U7771 (N_7771,N_7662,N_7706);
or U7772 (N_7772,N_7664,N_7633);
nand U7773 (N_7773,N_7641,N_7708);
xnor U7774 (N_7774,N_7718,N_7678);
and U7775 (N_7775,N_7628,N_7744);
xnor U7776 (N_7776,N_7747,N_7677);
nor U7777 (N_7777,N_7702,N_7645);
and U7778 (N_7778,N_7700,N_7692);
nor U7779 (N_7779,N_7668,N_7639);
xor U7780 (N_7780,N_7725,N_7672);
nor U7781 (N_7781,N_7714,N_7660);
and U7782 (N_7782,N_7670,N_7729);
nand U7783 (N_7783,N_7712,N_7689);
xnor U7784 (N_7784,N_7732,N_7673);
and U7785 (N_7785,N_7743,N_7724);
or U7786 (N_7786,N_7675,N_7657);
xor U7787 (N_7787,N_7655,N_7707);
and U7788 (N_7788,N_7699,N_7682);
or U7789 (N_7789,N_7722,N_7694);
xor U7790 (N_7790,N_7644,N_7710);
nor U7791 (N_7791,N_7738,N_7697);
and U7792 (N_7792,N_7679,N_7734);
and U7793 (N_7793,N_7746,N_7728);
or U7794 (N_7794,N_7637,N_7663);
nor U7795 (N_7795,N_7737,N_7684);
nor U7796 (N_7796,N_7736,N_7636);
or U7797 (N_7797,N_7627,N_7730);
xnor U7798 (N_7798,N_7651,N_7661);
nand U7799 (N_7799,N_7671,N_7635);
nand U7800 (N_7800,N_7688,N_7693);
and U7801 (N_7801,N_7686,N_7749);
xnor U7802 (N_7802,N_7721,N_7653);
and U7803 (N_7803,N_7709,N_7629);
nor U7804 (N_7804,N_7745,N_7713);
xor U7805 (N_7805,N_7676,N_7696);
xnor U7806 (N_7806,N_7705,N_7726);
xnor U7807 (N_7807,N_7632,N_7631);
nor U7808 (N_7808,N_7748,N_7640);
nand U7809 (N_7809,N_7711,N_7720);
nor U7810 (N_7810,N_7667,N_7687);
xnor U7811 (N_7811,N_7723,N_7659);
or U7812 (N_7812,N_7643,N_7677);
or U7813 (N_7813,N_7679,N_7726);
nand U7814 (N_7814,N_7676,N_7626);
nor U7815 (N_7815,N_7699,N_7627);
nand U7816 (N_7816,N_7732,N_7668);
nor U7817 (N_7817,N_7651,N_7659);
or U7818 (N_7818,N_7694,N_7669);
nand U7819 (N_7819,N_7683,N_7741);
nand U7820 (N_7820,N_7651,N_7688);
and U7821 (N_7821,N_7721,N_7681);
xnor U7822 (N_7822,N_7689,N_7694);
nor U7823 (N_7823,N_7630,N_7700);
or U7824 (N_7824,N_7672,N_7662);
or U7825 (N_7825,N_7698,N_7747);
or U7826 (N_7826,N_7704,N_7715);
or U7827 (N_7827,N_7745,N_7690);
xnor U7828 (N_7828,N_7651,N_7655);
nand U7829 (N_7829,N_7634,N_7638);
and U7830 (N_7830,N_7699,N_7629);
xnor U7831 (N_7831,N_7641,N_7671);
and U7832 (N_7832,N_7702,N_7685);
xor U7833 (N_7833,N_7685,N_7637);
nor U7834 (N_7834,N_7670,N_7699);
nor U7835 (N_7835,N_7636,N_7641);
nand U7836 (N_7836,N_7685,N_7745);
and U7837 (N_7837,N_7675,N_7636);
and U7838 (N_7838,N_7714,N_7647);
nand U7839 (N_7839,N_7657,N_7669);
nor U7840 (N_7840,N_7715,N_7638);
xor U7841 (N_7841,N_7666,N_7658);
or U7842 (N_7842,N_7629,N_7663);
nor U7843 (N_7843,N_7652,N_7709);
nand U7844 (N_7844,N_7632,N_7705);
or U7845 (N_7845,N_7689,N_7746);
xor U7846 (N_7846,N_7697,N_7670);
nand U7847 (N_7847,N_7675,N_7728);
nand U7848 (N_7848,N_7707,N_7689);
xor U7849 (N_7849,N_7681,N_7748);
and U7850 (N_7850,N_7634,N_7707);
and U7851 (N_7851,N_7696,N_7724);
nor U7852 (N_7852,N_7695,N_7744);
nand U7853 (N_7853,N_7693,N_7697);
and U7854 (N_7854,N_7723,N_7685);
nor U7855 (N_7855,N_7702,N_7643);
or U7856 (N_7856,N_7656,N_7731);
xnor U7857 (N_7857,N_7660,N_7670);
nand U7858 (N_7858,N_7724,N_7627);
and U7859 (N_7859,N_7719,N_7659);
or U7860 (N_7860,N_7666,N_7739);
or U7861 (N_7861,N_7644,N_7694);
nand U7862 (N_7862,N_7661,N_7653);
and U7863 (N_7863,N_7675,N_7627);
nand U7864 (N_7864,N_7695,N_7660);
xor U7865 (N_7865,N_7725,N_7668);
or U7866 (N_7866,N_7658,N_7632);
or U7867 (N_7867,N_7676,N_7627);
and U7868 (N_7868,N_7719,N_7725);
nand U7869 (N_7869,N_7700,N_7741);
nor U7870 (N_7870,N_7673,N_7685);
or U7871 (N_7871,N_7699,N_7677);
or U7872 (N_7872,N_7625,N_7655);
or U7873 (N_7873,N_7639,N_7663);
nand U7874 (N_7874,N_7697,N_7653);
nand U7875 (N_7875,N_7777,N_7835);
nand U7876 (N_7876,N_7802,N_7752);
nor U7877 (N_7877,N_7778,N_7789);
nor U7878 (N_7878,N_7786,N_7787);
and U7879 (N_7879,N_7838,N_7849);
nand U7880 (N_7880,N_7819,N_7825);
and U7881 (N_7881,N_7845,N_7826);
nor U7882 (N_7882,N_7824,N_7860);
nand U7883 (N_7883,N_7841,N_7776);
or U7884 (N_7884,N_7812,N_7830);
xor U7885 (N_7885,N_7754,N_7794);
nor U7886 (N_7886,N_7863,N_7839);
and U7887 (N_7887,N_7864,N_7766);
nand U7888 (N_7888,N_7798,N_7837);
nand U7889 (N_7889,N_7805,N_7840);
or U7890 (N_7890,N_7809,N_7851);
and U7891 (N_7891,N_7871,N_7764);
nor U7892 (N_7892,N_7829,N_7753);
xnor U7893 (N_7893,N_7822,N_7866);
xor U7894 (N_7894,N_7751,N_7765);
nor U7895 (N_7895,N_7813,N_7846);
and U7896 (N_7896,N_7795,N_7788);
or U7897 (N_7897,N_7781,N_7862);
or U7898 (N_7898,N_7821,N_7854);
nor U7899 (N_7899,N_7850,N_7779);
or U7900 (N_7900,N_7807,N_7796);
xnor U7901 (N_7901,N_7816,N_7803);
nand U7902 (N_7902,N_7844,N_7792);
nand U7903 (N_7903,N_7832,N_7793);
nand U7904 (N_7904,N_7769,N_7772);
and U7905 (N_7905,N_7759,N_7815);
and U7906 (N_7906,N_7833,N_7799);
or U7907 (N_7907,N_7783,N_7870);
and U7908 (N_7908,N_7827,N_7797);
nor U7909 (N_7909,N_7810,N_7872);
and U7910 (N_7910,N_7861,N_7828);
nor U7911 (N_7911,N_7859,N_7853);
nand U7912 (N_7912,N_7867,N_7852);
or U7913 (N_7913,N_7855,N_7820);
nand U7914 (N_7914,N_7873,N_7831);
and U7915 (N_7915,N_7808,N_7811);
xor U7916 (N_7916,N_7762,N_7814);
or U7917 (N_7917,N_7784,N_7757);
or U7918 (N_7918,N_7800,N_7823);
xor U7919 (N_7919,N_7770,N_7847);
or U7920 (N_7920,N_7750,N_7801);
and U7921 (N_7921,N_7768,N_7818);
and U7922 (N_7922,N_7804,N_7834);
or U7923 (N_7923,N_7865,N_7763);
nor U7924 (N_7924,N_7843,N_7858);
xnor U7925 (N_7925,N_7775,N_7791);
and U7926 (N_7926,N_7773,N_7760);
or U7927 (N_7927,N_7755,N_7785);
xor U7928 (N_7928,N_7774,N_7806);
and U7929 (N_7929,N_7756,N_7817);
and U7930 (N_7930,N_7842,N_7780);
or U7931 (N_7931,N_7874,N_7848);
xnor U7932 (N_7932,N_7868,N_7758);
or U7933 (N_7933,N_7790,N_7771);
and U7934 (N_7934,N_7761,N_7857);
nand U7935 (N_7935,N_7767,N_7856);
nor U7936 (N_7936,N_7836,N_7869);
nand U7937 (N_7937,N_7782,N_7862);
xnor U7938 (N_7938,N_7864,N_7806);
or U7939 (N_7939,N_7805,N_7778);
and U7940 (N_7940,N_7766,N_7795);
nand U7941 (N_7941,N_7778,N_7869);
nand U7942 (N_7942,N_7869,N_7849);
nor U7943 (N_7943,N_7854,N_7832);
nor U7944 (N_7944,N_7801,N_7834);
nand U7945 (N_7945,N_7839,N_7803);
nor U7946 (N_7946,N_7834,N_7864);
or U7947 (N_7947,N_7753,N_7833);
nand U7948 (N_7948,N_7763,N_7862);
xnor U7949 (N_7949,N_7769,N_7821);
nand U7950 (N_7950,N_7848,N_7854);
or U7951 (N_7951,N_7782,N_7776);
xor U7952 (N_7952,N_7792,N_7831);
nor U7953 (N_7953,N_7791,N_7836);
nand U7954 (N_7954,N_7763,N_7755);
xor U7955 (N_7955,N_7828,N_7805);
and U7956 (N_7956,N_7863,N_7840);
xor U7957 (N_7957,N_7865,N_7812);
nand U7958 (N_7958,N_7790,N_7874);
xor U7959 (N_7959,N_7852,N_7808);
nand U7960 (N_7960,N_7760,N_7790);
nor U7961 (N_7961,N_7754,N_7824);
or U7962 (N_7962,N_7829,N_7751);
nand U7963 (N_7963,N_7814,N_7841);
nor U7964 (N_7964,N_7780,N_7789);
nor U7965 (N_7965,N_7850,N_7801);
or U7966 (N_7966,N_7836,N_7830);
and U7967 (N_7967,N_7797,N_7809);
or U7968 (N_7968,N_7857,N_7864);
nor U7969 (N_7969,N_7820,N_7760);
nor U7970 (N_7970,N_7755,N_7874);
and U7971 (N_7971,N_7828,N_7855);
nor U7972 (N_7972,N_7853,N_7820);
nand U7973 (N_7973,N_7834,N_7781);
nand U7974 (N_7974,N_7822,N_7807);
nor U7975 (N_7975,N_7771,N_7750);
nor U7976 (N_7976,N_7804,N_7874);
nand U7977 (N_7977,N_7812,N_7759);
and U7978 (N_7978,N_7795,N_7765);
or U7979 (N_7979,N_7804,N_7812);
nor U7980 (N_7980,N_7843,N_7758);
nand U7981 (N_7981,N_7811,N_7845);
nand U7982 (N_7982,N_7781,N_7845);
or U7983 (N_7983,N_7816,N_7798);
and U7984 (N_7984,N_7814,N_7857);
or U7985 (N_7985,N_7753,N_7800);
and U7986 (N_7986,N_7776,N_7811);
xor U7987 (N_7987,N_7761,N_7805);
nand U7988 (N_7988,N_7844,N_7863);
or U7989 (N_7989,N_7815,N_7807);
xor U7990 (N_7990,N_7790,N_7843);
or U7991 (N_7991,N_7850,N_7849);
nor U7992 (N_7992,N_7780,N_7776);
and U7993 (N_7993,N_7783,N_7867);
xor U7994 (N_7994,N_7778,N_7861);
or U7995 (N_7995,N_7870,N_7799);
nand U7996 (N_7996,N_7864,N_7772);
xor U7997 (N_7997,N_7830,N_7794);
and U7998 (N_7998,N_7849,N_7783);
nand U7999 (N_7999,N_7754,N_7809);
nand U8000 (N_8000,N_7912,N_7911);
or U8001 (N_8001,N_7910,N_7905);
or U8002 (N_8002,N_7875,N_7962);
nand U8003 (N_8003,N_7983,N_7935);
nor U8004 (N_8004,N_7880,N_7895);
nor U8005 (N_8005,N_7918,N_7921);
nand U8006 (N_8006,N_7967,N_7960);
or U8007 (N_8007,N_7986,N_7941);
and U8008 (N_8008,N_7946,N_7975);
or U8009 (N_8009,N_7897,N_7878);
and U8010 (N_8010,N_7898,N_7973);
and U8011 (N_8011,N_7926,N_7953);
and U8012 (N_8012,N_7977,N_7970);
nor U8013 (N_8013,N_7996,N_7879);
nand U8014 (N_8014,N_7890,N_7995);
nand U8015 (N_8015,N_7952,N_7957);
nor U8016 (N_8016,N_7954,N_7903);
or U8017 (N_8017,N_7914,N_7981);
nor U8018 (N_8018,N_7915,N_7951);
nor U8019 (N_8019,N_7959,N_7929);
and U8020 (N_8020,N_7998,N_7987);
or U8021 (N_8021,N_7876,N_7945);
nor U8022 (N_8022,N_7931,N_7938);
and U8023 (N_8023,N_7949,N_7989);
and U8024 (N_8024,N_7950,N_7992);
xor U8025 (N_8025,N_7932,N_7974);
nor U8026 (N_8026,N_7881,N_7899);
xor U8027 (N_8027,N_7990,N_7980);
xnor U8028 (N_8028,N_7947,N_7939);
xor U8029 (N_8029,N_7877,N_7901);
nand U8030 (N_8030,N_7942,N_7985);
or U8031 (N_8031,N_7891,N_7893);
xnor U8032 (N_8032,N_7979,N_7968);
or U8033 (N_8033,N_7982,N_7896);
nand U8034 (N_8034,N_7991,N_7955);
nor U8035 (N_8035,N_7940,N_7923);
nor U8036 (N_8036,N_7965,N_7925);
nor U8037 (N_8037,N_7907,N_7964);
nand U8038 (N_8038,N_7885,N_7930);
nor U8039 (N_8039,N_7976,N_7971);
xnor U8040 (N_8040,N_7944,N_7943);
nand U8041 (N_8041,N_7963,N_7994);
nand U8042 (N_8042,N_7958,N_7886);
nor U8043 (N_8043,N_7894,N_7920);
xor U8044 (N_8044,N_7908,N_7999);
and U8045 (N_8045,N_7969,N_7936);
or U8046 (N_8046,N_7972,N_7889);
nand U8047 (N_8047,N_7892,N_7937);
nand U8048 (N_8048,N_7913,N_7906);
xnor U8049 (N_8049,N_7927,N_7924);
nor U8050 (N_8050,N_7956,N_7919);
nor U8051 (N_8051,N_7993,N_7966);
xor U8052 (N_8052,N_7978,N_7909);
nand U8053 (N_8053,N_7884,N_7883);
xor U8054 (N_8054,N_7997,N_7887);
and U8055 (N_8055,N_7961,N_7917);
and U8056 (N_8056,N_7904,N_7922);
xnor U8057 (N_8057,N_7902,N_7888);
and U8058 (N_8058,N_7882,N_7948);
nor U8059 (N_8059,N_7928,N_7916);
and U8060 (N_8060,N_7933,N_7934);
or U8061 (N_8061,N_7984,N_7988);
nand U8062 (N_8062,N_7900,N_7971);
or U8063 (N_8063,N_7988,N_7946);
and U8064 (N_8064,N_7973,N_7894);
nor U8065 (N_8065,N_7878,N_7967);
and U8066 (N_8066,N_7882,N_7990);
and U8067 (N_8067,N_7881,N_7884);
and U8068 (N_8068,N_7907,N_7940);
or U8069 (N_8069,N_7996,N_7898);
xor U8070 (N_8070,N_7952,N_7897);
and U8071 (N_8071,N_7985,N_7962);
nand U8072 (N_8072,N_7945,N_7931);
and U8073 (N_8073,N_7930,N_7984);
or U8074 (N_8074,N_7969,N_7948);
nor U8075 (N_8075,N_7995,N_7917);
xnor U8076 (N_8076,N_7919,N_7954);
or U8077 (N_8077,N_7937,N_7983);
nand U8078 (N_8078,N_7881,N_7955);
nand U8079 (N_8079,N_7893,N_7897);
xnor U8080 (N_8080,N_7880,N_7943);
or U8081 (N_8081,N_7926,N_7879);
xor U8082 (N_8082,N_7924,N_7970);
xnor U8083 (N_8083,N_7946,N_7942);
xnor U8084 (N_8084,N_7904,N_7926);
nor U8085 (N_8085,N_7888,N_7950);
nor U8086 (N_8086,N_7993,N_7988);
xor U8087 (N_8087,N_7926,N_7983);
nor U8088 (N_8088,N_7905,N_7899);
and U8089 (N_8089,N_7884,N_7949);
xor U8090 (N_8090,N_7944,N_7930);
xnor U8091 (N_8091,N_7892,N_7963);
or U8092 (N_8092,N_7924,N_7912);
nor U8093 (N_8093,N_7974,N_7968);
nand U8094 (N_8094,N_7971,N_7972);
nand U8095 (N_8095,N_7963,N_7894);
xnor U8096 (N_8096,N_7965,N_7949);
xor U8097 (N_8097,N_7937,N_7969);
and U8098 (N_8098,N_7879,N_7976);
and U8099 (N_8099,N_7897,N_7982);
nor U8100 (N_8100,N_7941,N_7915);
xnor U8101 (N_8101,N_7974,N_7975);
or U8102 (N_8102,N_7878,N_7921);
or U8103 (N_8103,N_7980,N_7974);
and U8104 (N_8104,N_7884,N_7990);
nor U8105 (N_8105,N_7982,N_7952);
and U8106 (N_8106,N_7883,N_7966);
nand U8107 (N_8107,N_7923,N_7969);
nor U8108 (N_8108,N_7964,N_7880);
or U8109 (N_8109,N_7920,N_7903);
xnor U8110 (N_8110,N_7944,N_7965);
nand U8111 (N_8111,N_7961,N_7978);
or U8112 (N_8112,N_7952,N_7901);
or U8113 (N_8113,N_7880,N_7916);
nand U8114 (N_8114,N_7969,N_7961);
xnor U8115 (N_8115,N_7968,N_7930);
nand U8116 (N_8116,N_7881,N_7989);
and U8117 (N_8117,N_7896,N_7994);
nor U8118 (N_8118,N_7932,N_7904);
nand U8119 (N_8119,N_7882,N_7881);
or U8120 (N_8120,N_7970,N_7933);
nand U8121 (N_8121,N_7954,N_7967);
nand U8122 (N_8122,N_7932,N_7887);
nor U8123 (N_8123,N_7948,N_7958);
nand U8124 (N_8124,N_7906,N_7942);
xnor U8125 (N_8125,N_8121,N_8057);
nand U8126 (N_8126,N_8117,N_8072);
xor U8127 (N_8127,N_8116,N_8065);
xor U8128 (N_8128,N_8005,N_8031);
xnor U8129 (N_8129,N_8046,N_8011);
nor U8130 (N_8130,N_8026,N_8093);
and U8131 (N_8131,N_8100,N_8099);
and U8132 (N_8132,N_8052,N_8067);
or U8133 (N_8133,N_8101,N_8069);
xnor U8134 (N_8134,N_8013,N_8114);
nand U8135 (N_8135,N_8029,N_8064);
nor U8136 (N_8136,N_8016,N_8086);
xnor U8137 (N_8137,N_8043,N_8090);
nor U8138 (N_8138,N_8014,N_8058);
and U8139 (N_8139,N_8035,N_8103);
and U8140 (N_8140,N_8083,N_8006);
nor U8141 (N_8141,N_8056,N_8060);
nand U8142 (N_8142,N_8082,N_8107);
xor U8143 (N_8143,N_8028,N_8092);
xnor U8144 (N_8144,N_8078,N_8094);
or U8145 (N_8145,N_8084,N_8113);
or U8146 (N_8146,N_8124,N_8112);
or U8147 (N_8147,N_8027,N_8024);
and U8148 (N_8148,N_8081,N_8044);
xnor U8149 (N_8149,N_8012,N_8076);
or U8150 (N_8150,N_8106,N_8021);
nand U8151 (N_8151,N_8001,N_8095);
nor U8152 (N_8152,N_8073,N_8119);
nor U8153 (N_8153,N_8080,N_8025);
and U8154 (N_8154,N_8087,N_8111);
and U8155 (N_8155,N_8068,N_8074);
nand U8156 (N_8156,N_8037,N_8048);
and U8157 (N_8157,N_8091,N_8017);
nand U8158 (N_8158,N_8104,N_8059);
and U8159 (N_8159,N_8015,N_8075);
nor U8160 (N_8160,N_8034,N_8007);
nand U8161 (N_8161,N_8110,N_8105);
nand U8162 (N_8162,N_8030,N_8000);
nand U8163 (N_8163,N_8122,N_8045);
or U8164 (N_8164,N_8061,N_8102);
xnor U8165 (N_8165,N_8018,N_8120);
and U8166 (N_8166,N_8108,N_8062);
or U8167 (N_8167,N_8042,N_8050);
xor U8168 (N_8168,N_8097,N_8070);
nand U8169 (N_8169,N_8010,N_8079);
nand U8170 (N_8170,N_8019,N_8123);
xor U8171 (N_8171,N_8055,N_8009);
and U8172 (N_8172,N_8040,N_8003);
nand U8173 (N_8173,N_8051,N_8023);
xnor U8174 (N_8174,N_8002,N_8004);
or U8175 (N_8175,N_8036,N_8088);
nor U8176 (N_8176,N_8032,N_8039);
and U8177 (N_8177,N_8115,N_8008);
or U8178 (N_8178,N_8022,N_8033);
xnor U8179 (N_8179,N_8066,N_8089);
or U8180 (N_8180,N_8098,N_8049);
and U8181 (N_8181,N_8053,N_8047);
or U8182 (N_8182,N_8096,N_8071);
or U8183 (N_8183,N_8085,N_8020);
nand U8184 (N_8184,N_8054,N_8109);
and U8185 (N_8185,N_8063,N_8041);
or U8186 (N_8186,N_8118,N_8077);
nor U8187 (N_8187,N_8038,N_8077);
and U8188 (N_8188,N_8117,N_8040);
nand U8189 (N_8189,N_8067,N_8015);
xnor U8190 (N_8190,N_8035,N_8087);
nor U8191 (N_8191,N_8003,N_8069);
or U8192 (N_8192,N_8073,N_8108);
nor U8193 (N_8193,N_8025,N_8116);
nand U8194 (N_8194,N_8049,N_8009);
or U8195 (N_8195,N_8034,N_8083);
nor U8196 (N_8196,N_8110,N_8081);
or U8197 (N_8197,N_8110,N_8077);
and U8198 (N_8198,N_8035,N_8054);
xnor U8199 (N_8199,N_8013,N_8124);
nor U8200 (N_8200,N_8099,N_8024);
nand U8201 (N_8201,N_8015,N_8060);
nand U8202 (N_8202,N_8113,N_8025);
or U8203 (N_8203,N_8069,N_8050);
nand U8204 (N_8204,N_8024,N_8015);
nor U8205 (N_8205,N_8011,N_8081);
nor U8206 (N_8206,N_8088,N_8075);
xnor U8207 (N_8207,N_8076,N_8123);
or U8208 (N_8208,N_8032,N_8003);
xor U8209 (N_8209,N_8066,N_8014);
or U8210 (N_8210,N_8054,N_8029);
nor U8211 (N_8211,N_8123,N_8097);
or U8212 (N_8212,N_8028,N_8048);
nor U8213 (N_8213,N_8009,N_8002);
nand U8214 (N_8214,N_8054,N_8011);
nor U8215 (N_8215,N_8058,N_8097);
xor U8216 (N_8216,N_8090,N_8050);
xnor U8217 (N_8217,N_8116,N_8015);
nand U8218 (N_8218,N_8020,N_8065);
and U8219 (N_8219,N_8068,N_8100);
xnor U8220 (N_8220,N_8113,N_8075);
and U8221 (N_8221,N_8052,N_8064);
or U8222 (N_8222,N_8034,N_8060);
or U8223 (N_8223,N_8065,N_8106);
and U8224 (N_8224,N_8107,N_8087);
or U8225 (N_8225,N_8100,N_8102);
xnor U8226 (N_8226,N_8118,N_8023);
xnor U8227 (N_8227,N_8031,N_8105);
nor U8228 (N_8228,N_8048,N_8095);
xor U8229 (N_8229,N_8037,N_8087);
and U8230 (N_8230,N_8095,N_8058);
nor U8231 (N_8231,N_8020,N_8099);
nand U8232 (N_8232,N_8062,N_8105);
or U8233 (N_8233,N_8104,N_8035);
nand U8234 (N_8234,N_8089,N_8014);
xnor U8235 (N_8235,N_8083,N_8002);
nor U8236 (N_8236,N_8058,N_8002);
nor U8237 (N_8237,N_8074,N_8056);
xnor U8238 (N_8238,N_8071,N_8008);
nor U8239 (N_8239,N_8071,N_8040);
nor U8240 (N_8240,N_8075,N_8098);
nand U8241 (N_8241,N_8033,N_8042);
or U8242 (N_8242,N_8024,N_8039);
nor U8243 (N_8243,N_8042,N_8115);
or U8244 (N_8244,N_8120,N_8068);
nand U8245 (N_8245,N_8009,N_8111);
nor U8246 (N_8246,N_8118,N_8088);
nor U8247 (N_8247,N_8083,N_8081);
nor U8248 (N_8248,N_8116,N_8018);
xnor U8249 (N_8249,N_8082,N_8073);
or U8250 (N_8250,N_8208,N_8151);
nor U8251 (N_8251,N_8238,N_8247);
or U8252 (N_8252,N_8148,N_8199);
or U8253 (N_8253,N_8156,N_8154);
or U8254 (N_8254,N_8188,N_8183);
nor U8255 (N_8255,N_8157,N_8165);
nand U8256 (N_8256,N_8173,N_8219);
nor U8257 (N_8257,N_8245,N_8166);
nand U8258 (N_8258,N_8131,N_8137);
nand U8259 (N_8259,N_8187,N_8202);
nor U8260 (N_8260,N_8223,N_8220);
or U8261 (N_8261,N_8175,N_8159);
nand U8262 (N_8262,N_8239,N_8136);
xor U8263 (N_8263,N_8170,N_8143);
and U8264 (N_8264,N_8232,N_8164);
or U8265 (N_8265,N_8204,N_8162);
nor U8266 (N_8266,N_8152,N_8182);
nor U8267 (N_8267,N_8218,N_8216);
nand U8268 (N_8268,N_8209,N_8194);
and U8269 (N_8269,N_8190,N_8210);
xor U8270 (N_8270,N_8142,N_8177);
or U8271 (N_8271,N_8158,N_8144);
or U8272 (N_8272,N_8172,N_8125);
nor U8273 (N_8273,N_8217,N_8180);
and U8274 (N_8274,N_8244,N_8129);
nor U8275 (N_8275,N_8213,N_8127);
xor U8276 (N_8276,N_8193,N_8168);
or U8277 (N_8277,N_8149,N_8160);
xnor U8278 (N_8278,N_8207,N_8241);
xnor U8279 (N_8279,N_8249,N_8132);
xor U8280 (N_8280,N_8184,N_8248);
nor U8281 (N_8281,N_8196,N_8153);
or U8282 (N_8282,N_8133,N_8169);
nand U8283 (N_8283,N_8135,N_8211);
and U8284 (N_8284,N_8130,N_8195);
nor U8285 (N_8285,N_8226,N_8222);
nand U8286 (N_8286,N_8230,N_8240);
or U8287 (N_8287,N_8215,N_8201);
or U8288 (N_8288,N_8139,N_8192);
nor U8289 (N_8289,N_8246,N_8147);
xor U8290 (N_8290,N_8214,N_8212);
nor U8291 (N_8291,N_8186,N_8237);
xor U8292 (N_8292,N_8181,N_8243);
xnor U8293 (N_8293,N_8163,N_8242);
nand U8294 (N_8294,N_8145,N_8171);
nor U8295 (N_8295,N_8178,N_8134);
nor U8296 (N_8296,N_8234,N_8200);
or U8297 (N_8297,N_8221,N_8126);
nand U8298 (N_8298,N_8224,N_8197);
xor U8299 (N_8299,N_8176,N_8174);
nor U8300 (N_8300,N_8198,N_8225);
nor U8301 (N_8301,N_8141,N_8146);
xor U8302 (N_8302,N_8229,N_8155);
xnor U8303 (N_8303,N_8203,N_8227);
xor U8304 (N_8304,N_8140,N_8231);
nand U8305 (N_8305,N_8233,N_8236);
nand U8306 (N_8306,N_8167,N_8138);
xor U8307 (N_8307,N_8185,N_8189);
and U8308 (N_8308,N_8191,N_8206);
nor U8309 (N_8309,N_8235,N_8128);
nand U8310 (N_8310,N_8179,N_8161);
or U8311 (N_8311,N_8228,N_8205);
nor U8312 (N_8312,N_8150,N_8174);
nand U8313 (N_8313,N_8206,N_8214);
xor U8314 (N_8314,N_8156,N_8132);
xnor U8315 (N_8315,N_8132,N_8232);
xor U8316 (N_8316,N_8181,N_8220);
or U8317 (N_8317,N_8134,N_8227);
or U8318 (N_8318,N_8154,N_8147);
xor U8319 (N_8319,N_8149,N_8161);
xnor U8320 (N_8320,N_8230,N_8227);
xor U8321 (N_8321,N_8175,N_8236);
nand U8322 (N_8322,N_8144,N_8179);
and U8323 (N_8323,N_8145,N_8141);
xor U8324 (N_8324,N_8218,N_8179);
xor U8325 (N_8325,N_8248,N_8221);
xor U8326 (N_8326,N_8186,N_8187);
nor U8327 (N_8327,N_8134,N_8128);
nand U8328 (N_8328,N_8168,N_8192);
or U8329 (N_8329,N_8188,N_8181);
or U8330 (N_8330,N_8155,N_8186);
or U8331 (N_8331,N_8214,N_8211);
nand U8332 (N_8332,N_8148,N_8223);
and U8333 (N_8333,N_8134,N_8237);
and U8334 (N_8334,N_8229,N_8214);
nor U8335 (N_8335,N_8140,N_8248);
nor U8336 (N_8336,N_8132,N_8167);
or U8337 (N_8337,N_8247,N_8158);
or U8338 (N_8338,N_8163,N_8143);
nand U8339 (N_8339,N_8226,N_8144);
and U8340 (N_8340,N_8136,N_8203);
nand U8341 (N_8341,N_8206,N_8219);
xor U8342 (N_8342,N_8141,N_8167);
xor U8343 (N_8343,N_8188,N_8197);
xor U8344 (N_8344,N_8150,N_8194);
nand U8345 (N_8345,N_8206,N_8159);
nor U8346 (N_8346,N_8187,N_8158);
and U8347 (N_8347,N_8244,N_8169);
nand U8348 (N_8348,N_8163,N_8144);
xor U8349 (N_8349,N_8195,N_8127);
xor U8350 (N_8350,N_8189,N_8179);
xor U8351 (N_8351,N_8208,N_8167);
nand U8352 (N_8352,N_8147,N_8204);
or U8353 (N_8353,N_8216,N_8245);
nand U8354 (N_8354,N_8177,N_8217);
or U8355 (N_8355,N_8197,N_8158);
xnor U8356 (N_8356,N_8170,N_8169);
or U8357 (N_8357,N_8199,N_8149);
and U8358 (N_8358,N_8155,N_8242);
and U8359 (N_8359,N_8239,N_8244);
nor U8360 (N_8360,N_8205,N_8239);
and U8361 (N_8361,N_8209,N_8224);
and U8362 (N_8362,N_8226,N_8177);
and U8363 (N_8363,N_8165,N_8243);
nand U8364 (N_8364,N_8133,N_8209);
nand U8365 (N_8365,N_8170,N_8180);
nand U8366 (N_8366,N_8126,N_8133);
nor U8367 (N_8367,N_8169,N_8129);
or U8368 (N_8368,N_8225,N_8235);
nor U8369 (N_8369,N_8179,N_8225);
or U8370 (N_8370,N_8173,N_8222);
xnor U8371 (N_8371,N_8245,N_8159);
and U8372 (N_8372,N_8238,N_8195);
or U8373 (N_8373,N_8214,N_8138);
nor U8374 (N_8374,N_8147,N_8161);
nand U8375 (N_8375,N_8259,N_8306);
nor U8376 (N_8376,N_8294,N_8369);
and U8377 (N_8377,N_8253,N_8335);
or U8378 (N_8378,N_8317,N_8302);
nor U8379 (N_8379,N_8373,N_8305);
nor U8380 (N_8380,N_8359,N_8268);
and U8381 (N_8381,N_8279,N_8320);
and U8382 (N_8382,N_8338,N_8367);
nor U8383 (N_8383,N_8311,N_8276);
and U8384 (N_8384,N_8301,N_8258);
and U8385 (N_8385,N_8303,N_8362);
xor U8386 (N_8386,N_8281,N_8256);
xor U8387 (N_8387,N_8345,N_8331);
nand U8388 (N_8388,N_8283,N_8348);
nand U8389 (N_8389,N_8290,N_8364);
nand U8390 (N_8390,N_8336,N_8263);
or U8391 (N_8391,N_8261,N_8368);
and U8392 (N_8392,N_8324,N_8333);
xnor U8393 (N_8393,N_8295,N_8291);
or U8394 (N_8394,N_8366,N_8262);
and U8395 (N_8395,N_8329,N_8354);
xor U8396 (N_8396,N_8323,N_8342);
nand U8397 (N_8397,N_8314,N_8327);
nor U8398 (N_8398,N_8353,N_8287);
xnor U8399 (N_8399,N_8312,N_8266);
nor U8400 (N_8400,N_8357,N_8271);
nand U8401 (N_8401,N_8264,N_8332);
and U8402 (N_8402,N_8289,N_8308);
xor U8403 (N_8403,N_8299,N_8252);
and U8404 (N_8404,N_8349,N_8278);
nor U8405 (N_8405,N_8282,N_8360);
or U8406 (N_8406,N_8292,N_8285);
xor U8407 (N_8407,N_8269,N_8339);
and U8408 (N_8408,N_8310,N_8255);
nor U8409 (N_8409,N_8374,N_8363);
nor U8410 (N_8410,N_8267,N_8273);
nand U8411 (N_8411,N_8326,N_8280);
nand U8412 (N_8412,N_8355,N_8260);
nor U8413 (N_8413,N_8270,N_8254);
and U8414 (N_8414,N_8344,N_8351);
or U8415 (N_8415,N_8288,N_8319);
and U8416 (N_8416,N_8325,N_8272);
or U8417 (N_8417,N_8361,N_8250);
and U8418 (N_8418,N_8265,N_8257);
nor U8419 (N_8419,N_8274,N_8341);
and U8420 (N_8420,N_8346,N_8275);
nand U8421 (N_8421,N_8352,N_8330);
xnor U8422 (N_8422,N_8315,N_8284);
xnor U8423 (N_8423,N_8337,N_8372);
or U8424 (N_8424,N_8334,N_8328);
and U8425 (N_8425,N_8340,N_8296);
and U8426 (N_8426,N_8293,N_8286);
xor U8427 (N_8427,N_8356,N_8370);
or U8428 (N_8428,N_8365,N_8316);
nor U8429 (N_8429,N_8251,N_8309);
nand U8430 (N_8430,N_8371,N_8358);
or U8431 (N_8431,N_8313,N_8350);
nand U8432 (N_8432,N_8343,N_8322);
xor U8433 (N_8433,N_8307,N_8298);
or U8434 (N_8434,N_8277,N_8347);
or U8435 (N_8435,N_8321,N_8318);
nor U8436 (N_8436,N_8300,N_8297);
nor U8437 (N_8437,N_8304,N_8362);
nand U8438 (N_8438,N_8336,N_8250);
nor U8439 (N_8439,N_8301,N_8360);
and U8440 (N_8440,N_8309,N_8311);
nor U8441 (N_8441,N_8286,N_8347);
and U8442 (N_8442,N_8372,N_8274);
or U8443 (N_8443,N_8372,N_8315);
nand U8444 (N_8444,N_8318,N_8259);
xor U8445 (N_8445,N_8291,N_8334);
nand U8446 (N_8446,N_8356,N_8290);
nand U8447 (N_8447,N_8317,N_8316);
and U8448 (N_8448,N_8262,N_8295);
nor U8449 (N_8449,N_8251,N_8322);
or U8450 (N_8450,N_8286,N_8261);
nand U8451 (N_8451,N_8298,N_8305);
or U8452 (N_8452,N_8357,N_8255);
nand U8453 (N_8453,N_8328,N_8314);
xnor U8454 (N_8454,N_8301,N_8321);
and U8455 (N_8455,N_8299,N_8262);
xnor U8456 (N_8456,N_8287,N_8308);
xor U8457 (N_8457,N_8306,N_8360);
or U8458 (N_8458,N_8298,N_8290);
nand U8459 (N_8459,N_8366,N_8301);
nor U8460 (N_8460,N_8362,N_8305);
and U8461 (N_8461,N_8299,N_8289);
xnor U8462 (N_8462,N_8361,N_8315);
nor U8463 (N_8463,N_8330,N_8344);
nor U8464 (N_8464,N_8252,N_8341);
nand U8465 (N_8465,N_8311,N_8345);
nor U8466 (N_8466,N_8263,N_8291);
and U8467 (N_8467,N_8357,N_8317);
xnor U8468 (N_8468,N_8348,N_8345);
xnor U8469 (N_8469,N_8319,N_8273);
and U8470 (N_8470,N_8314,N_8363);
nor U8471 (N_8471,N_8322,N_8317);
xor U8472 (N_8472,N_8331,N_8365);
xor U8473 (N_8473,N_8330,N_8276);
nand U8474 (N_8474,N_8334,N_8350);
nor U8475 (N_8475,N_8264,N_8343);
or U8476 (N_8476,N_8336,N_8268);
xor U8477 (N_8477,N_8295,N_8264);
nor U8478 (N_8478,N_8312,N_8259);
and U8479 (N_8479,N_8366,N_8349);
or U8480 (N_8480,N_8302,N_8285);
or U8481 (N_8481,N_8273,N_8358);
xor U8482 (N_8482,N_8289,N_8278);
nor U8483 (N_8483,N_8275,N_8300);
nand U8484 (N_8484,N_8314,N_8338);
nor U8485 (N_8485,N_8359,N_8341);
nor U8486 (N_8486,N_8301,N_8295);
or U8487 (N_8487,N_8303,N_8262);
nor U8488 (N_8488,N_8373,N_8257);
xor U8489 (N_8489,N_8312,N_8362);
nor U8490 (N_8490,N_8267,N_8264);
nor U8491 (N_8491,N_8305,N_8344);
nand U8492 (N_8492,N_8304,N_8332);
nor U8493 (N_8493,N_8365,N_8362);
nand U8494 (N_8494,N_8255,N_8331);
xor U8495 (N_8495,N_8332,N_8333);
and U8496 (N_8496,N_8357,N_8354);
and U8497 (N_8497,N_8329,N_8263);
xnor U8498 (N_8498,N_8282,N_8333);
nand U8499 (N_8499,N_8336,N_8275);
nor U8500 (N_8500,N_8491,N_8478);
nor U8501 (N_8501,N_8420,N_8452);
xnor U8502 (N_8502,N_8406,N_8460);
and U8503 (N_8503,N_8459,N_8484);
nand U8504 (N_8504,N_8441,N_8380);
nand U8505 (N_8505,N_8475,N_8450);
xnor U8506 (N_8506,N_8423,N_8432);
and U8507 (N_8507,N_8447,N_8403);
nor U8508 (N_8508,N_8477,N_8474);
nor U8509 (N_8509,N_8488,N_8487);
or U8510 (N_8510,N_8396,N_8387);
and U8511 (N_8511,N_8411,N_8449);
or U8512 (N_8512,N_8457,N_8443);
or U8513 (N_8513,N_8461,N_8481);
or U8514 (N_8514,N_8456,N_8498);
nand U8515 (N_8515,N_8472,N_8405);
or U8516 (N_8516,N_8421,N_8383);
nand U8517 (N_8517,N_8410,N_8479);
or U8518 (N_8518,N_8429,N_8390);
xnor U8519 (N_8519,N_8399,N_8400);
and U8520 (N_8520,N_8430,N_8480);
xnor U8521 (N_8521,N_8376,N_8385);
and U8522 (N_8522,N_8473,N_8428);
xnor U8523 (N_8523,N_8397,N_8495);
and U8524 (N_8524,N_8407,N_8448);
or U8525 (N_8525,N_8416,N_8438);
or U8526 (N_8526,N_8377,N_8389);
nand U8527 (N_8527,N_8466,N_8493);
or U8528 (N_8528,N_8388,N_8497);
xor U8529 (N_8529,N_8436,N_8465);
nand U8530 (N_8530,N_8482,N_8454);
nand U8531 (N_8531,N_8492,N_8418);
nand U8532 (N_8532,N_8409,N_8381);
or U8533 (N_8533,N_8453,N_8468);
or U8534 (N_8534,N_8490,N_8485);
xnor U8535 (N_8535,N_8417,N_8398);
xor U8536 (N_8536,N_8375,N_8499);
nor U8537 (N_8537,N_8408,N_8455);
or U8538 (N_8538,N_8433,N_8422);
or U8539 (N_8539,N_8404,N_8412);
or U8540 (N_8540,N_8469,N_8445);
and U8541 (N_8541,N_8467,N_8431);
nor U8542 (N_8542,N_8391,N_8442);
nor U8543 (N_8543,N_8496,N_8419);
and U8544 (N_8544,N_8427,N_8462);
or U8545 (N_8545,N_8463,N_8470);
xor U8546 (N_8546,N_8425,N_8437);
nand U8547 (N_8547,N_8444,N_8384);
xnor U8548 (N_8548,N_8489,N_8401);
or U8549 (N_8549,N_8439,N_8434);
nor U8550 (N_8550,N_8435,N_8471);
nor U8551 (N_8551,N_8464,N_8483);
or U8552 (N_8552,N_8486,N_8446);
nor U8553 (N_8553,N_8402,N_8393);
nor U8554 (N_8554,N_8392,N_8378);
nor U8555 (N_8555,N_8382,N_8379);
xor U8556 (N_8556,N_8395,N_8394);
xor U8557 (N_8557,N_8413,N_8414);
or U8558 (N_8558,N_8386,N_8440);
and U8559 (N_8559,N_8458,N_8415);
or U8560 (N_8560,N_8494,N_8426);
or U8561 (N_8561,N_8424,N_8476);
nand U8562 (N_8562,N_8451,N_8463);
xor U8563 (N_8563,N_8448,N_8395);
or U8564 (N_8564,N_8481,N_8402);
or U8565 (N_8565,N_8398,N_8426);
nor U8566 (N_8566,N_8412,N_8489);
xor U8567 (N_8567,N_8383,N_8382);
and U8568 (N_8568,N_8461,N_8471);
or U8569 (N_8569,N_8452,N_8397);
nand U8570 (N_8570,N_8497,N_8492);
and U8571 (N_8571,N_8401,N_8469);
nand U8572 (N_8572,N_8494,N_8432);
xor U8573 (N_8573,N_8499,N_8484);
nand U8574 (N_8574,N_8437,N_8408);
nor U8575 (N_8575,N_8471,N_8412);
nand U8576 (N_8576,N_8497,N_8491);
and U8577 (N_8577,N_8460,N_8411);
nand U8578 (N_8578,N_8455,N_8388);
nand U8579 (N_8579,N_8475,N_8448);
and U8580 (N_8580,N_8486,N_8471);
nor U8581 (N_8581,N_8400,N_8459);
or U8582 (N_8582,N_8468,N_8479);
xnor U8583 (N_8583,N_8388,N_8422);
and U8584 (N_8584,N_8457,N_8438);
nand U8585 (N_8585,N_8472,N_8457);
xor U8586 (N_8586,N_8395,N_8446);
nor U8587 (N_8587,N_8449,N_8455);
nor U8588 (N_8588,N_8401,N_8493);
nand U8589 (N_8589,N_8435,N_8459);
and U8590 (N_8590,N_8491,N_8486);
and U8591 (N_8591,N_8458,N_8449);
xnor U8592 (N_8592,N_8431,N_8466);
nor U8593 (N_8593,N_8462,N_8392);
and U8594 (N_8594,N_8379,N_8392);
and U8595 (N_8595,N_8440,N_8493);
xnor U8596 (N_8596,N_8400,N_8412);
xnor U8597 (N_8597,N_8426,N_8464);
xnor U8598 (N_8598,N_8427,N_8423);
nand U8599 (N_8599,N_8388,N_8396);
xnor U8600 (N_8600,N_8495,N_8432);
xor U8601 (N_8601,N_8402,N_8429);
nand U8602 (N_8602,N_8466,N_8391);
nor U8603 (N_8603,N_8380,N_8384);
and U8604 (N_8604,N_8464,N_8406);
or U8605 (N_8605,N_8388,N_8434);
or U8606 (N_8606,N_8466,N_8394);
nor U8607 (N_8607,N_8412,N_8379);
nand U8608 (N_8608,N_8492,N_8453);
nand U8609 (N_8609,N_8467,N_8447);
nand U8610 (N_8610,N_8437,N_8469);
xnor U8611 (N_8611,N_8452,N_8400);
or U8612 (N_8612,N_8469,N_8456);
xor U8613 (N_8613,N_8493,N_8467);
nor U8614 (N_8614,N_8453,N_8476);
nor U8615 (N_8615,N_8408,N_8391);
xnor U8616 (N_8616,N_8459,N_8438);
or U8617 (N_8617,N_8427,N_8403);
xnor U8618 (N_8618,N_8392,N_8439);
nor U8619 (N_8619,N_8482,N_8453);
nand U8620 (N_8620,N_8412,N_8402);
xnor U8621 (N_8621,N_8378,N_8415);
nand U8622 (N_8622,N_8499,N_8400);
and U8623 (N_8623,N_8450,N_8426);
or U8624 (N_8624,N_8429,N_8424);
or U8625 (N_8625,N_8582,N_8547);
xor U8626 (N_8626,N_8518,N_8536);
or U8627 (N_8627,N_8604,N_8539);
or U8628 (N_8628,N_8602,N_8526);
nand U8629 (N_8629,N_8529,N_8623);
nand U8630 (N_8630,N_8624,N_8599);
nand U8631 (N_8631,N_8595,N_8504);
or U8632 (N_8632,N_8607,N_8580);
nor U8633 (N_8633,N_8519,N_8577);
xor U8634 (N_8634,N_8612,N_8611);
xnor U8635 (N_8635,N_8610,N_8520);
nor U8636 (N_8636,N_8578,N_8618);
xnor U8637 (N_8637,N_8558,N_8543);
or U8638 (N_8638,N_8613,N_8506);
or U8639 (N_8639,N_8572,N_8508);
xnor U8640 (N_8640,N_8592,N_8554);
or U8641 (N_8641,N_8565,N_8606);
or U8642 (N_8642,N_8524,N_8615);
and U8643 (N_8643,N_8523,N_8589);
and U8644 (N_8644,N_8574,N_8597);
and U8645 (N_8645,N_8593,N_8531);
xnor U8646 (N_8646,N_8511,N_8583);
nand U8647 (N_8647,N_8567,N_8517);
or U8648 (N_8648,N_8588,N_8616);
and U8649 (N_8649,N_8619,N_8561);
xor U8650 (N_8650,N_8548,N_8538);
nand U8651 (N_8651,N_8621,N_8552);
nor U8652 (N_8652,N_8515,N_8541);
xor U8653 (N_8653,N_8514,N_8591);
xnor U8654 (N_8654,N_8500,N_8581);
nand U8655 (N_8655,N_8601,N_8560);
nor U8656 (N_8656,N_8528,N_8614);
and U8657 (N_8657,N_8503,N_8537);
nand U8658 (N_8658,N_8509,N_8571);
or U8659 (N_8659,N_8516,N_8608);
nor U8660 (N_8660,N_8533,N_8603);
nor U8661 (N_8661,N_8521,N_8510);
or U8662 (N_8662,N_8596,N_8532);
xor U8663 (N_8663,N_8620,N_8598);
or U8664 (N_8664,N_8535,N_8556);
and U8665 (N_8665,N_8501,N_8566);
nor U8666 (N_8666,N_8573,N_8586);
or U8667 (N_8667,N_8512,N_8505);
nor U8668 (N_8668,N_8502,N_8594);
nand U8669 (N_8669,N_8590,N_8555);
or U8670 (N_8670,N_8600,N_8585);
nor U8671 (N_8671,N_8576,N_8534);
xor U8672 (N_8672,N_8564,N_8559);
or U8673 (N_8673,N_8605,N_8513);
or U8674 (N_8674,N_8622,N_8551);
nand U8675 (N_8675,N_8584,N_8579);
nor U8676 (N_8676,N_8525,N_8522);
and U8677 (N_8677,N_8609,N_8562);
or U8678 (N_8678,N_8550,N_8570);
nand U8679 (N_8679,N_8557,N_8544);
and U8680 (N_8680,N_8527,N_8553);
and U8681 (N_8681,N_8617,N_8540);
or U8682 (N_8682,N_8563,N_8568);
nor U8683 (N_8683,N_8569,N_8507);
nand U8684 (N_8684,N_8549,N_8587);
nor U8685 (N_8685,N_8575,N_8545);
nor U8686 (N_8686,N_8542,N_8530);
nor U8687 (N_8687,N_8546,N_8613);
nor U8688 (N_8688,N_8528,N_8566);
and U8689 (N_8689,N_8593,N_8571);
nor U8690 (N_8690,N_8532,N_8501);
and U8691 (N_8691,N_8623,N_8544);
or U8692 (N_8692,N_8509,N_8576);
and U8693 (N_8693,N_8530,N_8565);
and U8694 (N_8694,N_8614,N_8510);
xor U8695 (N_8695,N_8622,N_8539);
and U8696 (N_8696,N_8618,N_8588);
xnor U8697 (N_8697,N_8535,N_8521);
xor U8698 (N_8698,N_8532,N_8524);
nand U8699 (N_8699,N_8579,N_8539);
xnor U8700 (N_8700,N_8544,N_8601);
nor U8701 (N_8701,N_8597,N_8550);
nor U8702 (N_8702,N_8601,N_8562);
and U8703 (N_8703,N_8595,N_8522);
and U8704 (N_8704,N_8584,N_8567);
nand U8705 (N_8705,N_8571,N_8597);
nand U8706 (N_8706,N_8501,N_8616);
or U8707 (N_8707,N_8518,N_8516);
xnor U8708 (N_8708,N_8526,N_8597);
nor U8709 (N_8709,N_8572,N_8545);
or U8710 (N_8710,N_8544,N_8515);
or U8711 (N_8711,N_8542,N_8551);
xnor U8712 (N_8712,N_8515,N_8519);
xnor U8713 (N_8713,N_8531,N_8544);
xnor U8714 (N_8714,N_8592,N_8533);
or U8715 (N_8715,N_8502,N_8566);
xnor U8716 (N_8716,N_8523,N_8527);
and U8717 (N_8717,N_8517,N_8551);
nand U8718 (N_8718,N_8577,N_8516);
xnor U8719 (N_8719,N_8621,N_8519);
nand U8720 (N_8720,N_8537,N_8520);
nor U8721 (N_8721,N_8606,N_8563);
nand U8722 (N_8722,N_8500,N_8559);
nor U8723 (N_8723,N_8535,N_8623);
nand U8724 (N_8724,N_8538,N_8540);
and U8725 (N_8725,N_8513,N_8561);
nor U8726 (N_8726,N_8575,N_8542);
and U8727 (N_8727,N_8581,N_8619);
or U8728 (N_8728,N_8618,N_8616);
xnor U8729 (N_8729,N_8529,N_8589);
nor U8730 (N_8730,N_8576,N_8586);
and U8731 (N_8731,N_8623,N_8571);
and U8732 (N_8732,N_8556,N_8596);
xnor U8733 (N_8733,N_8567,N_8553);
or U8734 (N_8734,N_8558,N_8582);
xor U8735 (N_8735,N_8536,N_8583);
and U8736 (N_8736,N_8601,N_8609);
and U8737 (N_8737,N_8574,N_8581);
nor U8738 (N_8738,N_8528,N_8556);
and U8739 (N_8739,N_8595,N_8553);
and U8740 (N_8740,N_8561,N_8557);
xor U8741 (N_8741,N_8567,N_8543);
and U8742 (N_8742,N_8582,N_8529);
nand U8743 (N_8743,N_8589,N_8606);
nor U8744 (N_8744,N_8586,N_8610);
nor U8745 (N_8745,N_8584,N_8582);
nand U8746 (N_8746,N_8559,N_8515);
or U8747 (N_8747,N_8508,N_8518);
or U8748 (N_8748,N_8589,N_8583);
nand U8749 (N_8749,N_8588,N_8601);
xor U8750 (N_8750,N_8736,N_8661);
xor U8751 (N_8751,N_8677,N_8678);
or U8752 (N_8752,N_8628,N_8701);
or U8753 (N_8753,N_8702,N_8669);
or U8754 (N_8754,N_8627,N_8687);
nand U8755 (N_8755,N_8728,N_8690);
nand U8756 (N_8756,N_8682,N_8668);
nor U8757 (N_8757,N_8693,N_8703);
nand U8758 (N_8758,N_8667,N_8743);
nor U8759 (N_8759,N_8729,N_8663);
nor U8760 (N_8760,N_8730,N_8719);
xnor U8761 (N_8761,N_8652,N_8691);
nor U8762 (N_8762,N_8681,N_8686);
and U8763 (N_8763,N_8721,N_8657);
nor U8764 (N_8764,N_8699,N_8746);
or U8765 (N_8765,N_8723,N_8718);
and U8766 (N_8766,N_8732,N_8725);
nor U8767 (N_8767,N_8700,N_8670);
nor U8768 (N_8768,N_8696,N_8632);
or U8769 (N_8769,N_8711,N_8685);
xor U8770 (N_8770,N_8724,N_8655);
nand U8771 (N_8771,N_8708,N_8648);
and U8772 (N_8772,N_8705,N_8658);
nor U8773 (N_8773,N_8674,N_8650);
nand U8774 (N_8774,N_8709,N_8712);
xor U8775 (N_8775,N_8694,N_8731);
nand U8776 (N_8776,N_8737,N_8676);
or U8777 (N_8777,N_8643,N_8749);
nor U8778 (N_8778,N_8715,N_8664);
or U8779 (N_8779,N_8747,N_8706);
nand U8780 (N_8780,N_8722,N_8683);
nand U8781 (N_8781,N_8636,N_8653);
xor U8782 (N_8782,N_8645,N_8739);
or U8783 (N_8783,N_8727,N_8662);
nor U8784 (N_8784,N_8734,N_8741);
and U8785 (N_8785,N_8720,N_8704);
nor U8786 (N_8786,N_8630,N_8659);
nor U8787 (N_8787,N_8666,N_8697);
nand U8788 (N_8788,N_8633,N_8692);
or U8789 (N_8789,N_8646,N_8726);
nor U8790 (N_8790,N_8689,N_8626);
and U8791 (N_8791,N_8654,N_8625);
xor U8792 (N_8792,N_8640,N_8671);
nand U8793 (N_8793,N_8744,N_8688);
xnor U8794 (N_8794,N_8634,N_8707);
and U8795 (N_8795,N_8631,N_8713);
and U8796 (N_8796,N_8745,N_8695);
xnor U8797 (N_8797,N_8735,N_8638);
nor U8798 (N_8798,N_8651,N_8716);
nand U8799 (N_8799,N_8679,N_8684);
and U8800 (N_8800,N_8710,N_8675);
or U8801 (N_8801,N_8733,N_8717);
xor U8802 (N_8802,N_8672,N_8698);
nor U8803 (N_8803,N_8660,N_8642);
xor U8804 (N_8804,N_8738,N_8629);
nor U8805 (N_8805,N_8656,N_8742);
and U8806 (N_8806,N_8647,N_8649);
or U8807 (N_8807,N_8680,N_8635);
xnor U8808 (N_8808,N_8714,N_8673);
xnor U8809 (N_8809,N_8644,N_8748);
and U8810 (N_8810,N_8637,N_8641);
and U8811 (N_8811,N_8665,N_8639);
nor U8812 (N_8812,N_8740,N_8717);
nor U8813 (N_8813,N_8695,N_8730);
xnor U8814 (N_8814,N_8666,N_8663);
and U8815 (N_8815,N_8742,N_8698);
xnor U8816 (N_8816,N_8653,N_8648);
or U8817 (N_8817,N_8646,N_8714);
or U8818 (N_8818,N_8695,N_8686);
nor U8819 (N_8819,N_8704,N_8675);
and U8820 (N_8820,N_8690,N_8697);
nor U8821 (N_8821,N_8706,N_8678);
or U8822 (N_8822,N_8686,N_8739);
xor U8823 (N_8823,N_8667,N_8748);
xor U8824 (N_8824,N_8747,N_8705);
nand U8825 (N_8825,N_8724,N_8742);
or U8826 (N_8826,N_8650,N_8649);
or U8827 (N_8827,N_8665,N_8694);
nor U8828 (N_8828,N_8747,N_8734);
and U8829 (N_8829,N_8687,N_8671);
or U8830 (N_8830,N_8739,N_8653);
nor U8831 (N_8831,N_8638,N_8748);
nor U8832 (N_8832,N_8696,N_8743);
xnor U8833 (N_8833,N_8679,N_8740);
and U8834 (N_8834,N_8687,N_8678);
xor U8835 (N_8835,N_8659,N_8664);
nand U8836 (N_8836,N_8638,N_8652);
xor U8837 (N_8837,N_8686,N_8723);
or U8838 (N_8838,N_8636,N_8692);
and U8839 (N_8839,N_8737,N_8748);
nor U8840 (N_8840,N_8690,N_8669);
nand U8841 (N_8841,N_8636,N_8709);
xor U8842 (N_8842,N_8641,N_8710);
and U8843 (N_8843,N_8678,N_8705);
and U8844 (N_8844,N_8708,N_8721);
xnor U8845 (N_8845,N_8636,N_8651);
or U8846 (N_8846,N_8705,N_8659);
nor U8847 (N_8847,N_8680,N_8654);
nand U8848 (N_8848,N_8735,N_8705);
or U8849 (N_8849,N_8662,N_8663);
nand U8850 (N_8850,N_8627,N_8694);
nor U8851 (N_8851,N_8630,N_8714);
nand U8852 (N_8852,N_8741,N_8715);
nor U8853 (N_8853,N_8641,N_8645);
nor U8854 (N_8854,N_8731,N_8680);
xor U8855 (N_8855,N_8640,N_8635);
or U8856 (N_8856,N_8652,N_8747);
nor U8857 (N_8857,N_8697,N_8728);
and U8858 (N_8858,N_8687,N_8643);
nor U8859 (N_8859,N_8656,N_8699);
nor U8860 (N_8860,N_8654,N_8735);
xnor U8861 (N_8861,N_8723,N_8629);
and U8862 (N_8862,N_8699,N_8652);
xor U8863 (N_8863,N_8688,N_8661);
and U8864 (N_8864,N_8685,N_8735);
and U8865 (N_8865,N_8661,N_8742);
nor U8866 (N_8866,N_8746,N_8636);
nor U8867 (N_8867,N_8685,N_8746);
nor U8868 (N_8868,N_8710,N_8683);
nand U8869 (N_8869,N_8625,N_8720);
and U8870 (N_8870,N_8719,N_8646);
or U8871 (N_8871,N_8711,N_8733);
or U8872 (N_8872,N_8671,N_8713);
nor U8873 (N_8873,N_8724,N_8714);
nor U8874 (N_8874,N_8696,N_8633);
nand U8875 (N_8875,N_8854,N_8820);
nor U8876 (N_8876,N_8833,N_8819);
and U8877 (N_8877,N_8858,N_8774);
or U8878 (N_8878,N_8861,N_8825);
or U8879 (N_8879,N_8776,N_8766);
nor U8880 (N_8880,N_8836,N_8811);
nand U8881 (N_8881,N_8801,N_8756);
nand U8882 (N_8882,N_8871,N_8830);
xor U8883 (N_8883,N_8837,N_8794);
nor U8884 (N_8884,N_8761,N_8868);
nor U8885 (N_8885,N_8764,N_8855);
nand U8886 (N_8886,N_8831,N_8865);
or U8887 (N_8887,N_8818,N_8769);
nand U8888 (N_8888,N_8824,N_8823);
or U8889 (N_8889,N_8797,N_8753);
nor U8890 (N_8890,N_8847,N_8853);
and U8891 (N_8891,N_8852,N_8792);
or U8892 (N_8892,N_8846,N_8767);
xnor U8893 (N_8893,N_8803,N_8808);
xnor U8894 (N_8894,N_8786,N_8829);
and U8895 (N_8895,N_8799,N_8869);
nand U8896 (N_8896,N_8859,N_8780);
nand U8897 (N_8897,N_8812,N_8793);
nor U8898 (N_8898,N_8775,N_8750);
and U8899 (N_8899,N_8843,N_8784);
and U8900 (N_8900,N_8773,N_8874);
and U8901 (N_8901,N_8782,N_8813);
nor U8902 (N_8902,N_8788,N_8768);
or U8903 (N_8903,N_8867,N_8839);
nor U8904 (N_8904,N_8851,N_8844);
or U8905 (N_8905,N_8751,N_8815);
and U8906 (N_8906,N_8821,N_8850);
or U8907 (N_8907,N_8848,N_8762);
or U8908 (N_8908,N_8845,N_8770);
nor U8909 (N_8909,N_8835,N_8771);
and U8910 (N_8910,N_8787,N_8863);
nor U8911 (N_8911,N_8814,N_8834);
nor U8912 (N_8912,N_8760,N_8800);
or U8913 (N_8913,N_8870,N_8826);
xor U8914 (N_8914,N_8802,N_8790);
and U8915 (N_8915,N_8857,N_8804);
xor U8916 (N_8916,N_8841,N_8789);
nor U8917 (N_8917,N_8872,N_8755);
or U8918 (N_8918,N_8828,N_8758);
xor U8919 (N_8919,N_8783,N_8840);
xor U8920 (N_8920,N_8752,N_8860);
and U8921 (N_8921,N_8798,N_8765);
xor U8922 (N_8922,N_8759,N_8791);
nand U8923 (N_8923,N_8754,N_8849);
nor U8924 (N_8924,N_8805,N_8807);
xor U8925 (N_8925,N_8763,N_8866);
nor U8926 (N_8926,N_8778,N_8856);
nand U8927 (N_8927,N_8806,N_8842);
nand U8928 (N_8928,N_8795,N_8864);
or U8929 (N_8929,N_8827,N_8873);
xor U8930 (N_8930,N_8832,N_8816);
nand U8931 (N_8931,N_8810,N_8777);
or U8932 (N_8932,N_8809,N_8772);
or U8933 (N_8933,N_8817,N_8757);
and U8934 (N_8934,N_8796,N_8781);
and U8935 (N_8935,N_8862,N_8779);
or U8936 (N_8936,N_8822,N_8785);
nor U8937 (N_8937,N_8838,N_8863);
and U8938 (N_8938,N_8801,N_8828);
xnor U8939 (N_8939,N_8825,N_8866);
xnor U8940 (N_8940,N_8868,N_8844);
and U8941 (N_8941,N_8860,N_8788);
nand U8942 (N_8942,N_8851,N_8818);
or U8943 (N_8943,N_8769,N_8792);
xnor U8944 (N_8944,N_8797,N_8789);
nor U8945 (N_8945,N_8836,N_8787);
and U8946 (N_8946,N_8850,N_8762);
xor U8947 (N_8947,N_8851,N_8874);
or U8948 (N_8948,N_8804,N_8849);
and U8949 (N_8949,N_8782,N_8819);
xor U8950 (N_8950,N_8783,N_8761);
nand U8951 (N_8951,N_8784,N_8758);
or U8952 (N_8952,N_8805,N_8768);
or U8953 (N_8953,N_8856,N_8800);
or U8954 (N_8954,N_8872,N_8779);
nand U8955 (N_8955,N_8855,N_8844);
xnor U8956 (N_8956,N_8802,N_8858);
xor U8957 (N_8957,N_8808,N_8784);
or U8958 (N_8958,N_8856,N_8872);
and U8959 (N_8959,N_8757,N_8783);
or U8960 (N_8960,N_8872,N_8842);
and U8961 (N_8961,N_8807,N_8873);
and U8962 (N_8962,N_8797,N_8823);
xnor U8963 (N_8963,N_8874,N_8769);
nor U8964 (N_8964,N_8806,N_8820);
nand U8965 (N_8965,N_8799,N_8760);
nand U8966 (N_8966,N_8777,N_8869);
or U8967 (N_8967,N_8842,N_8759);
nand U8968 (N_8968,N_8825,N_8841);
xnor U8969 (N_8969,N_8840,N_8791);
nand U8970 (N_8970,N_8855,N_8797);
or U8971 (N_8971,N_8782,N_8779);
nor U8972 (N_8972,N_8754,N_8790);
xnor U8973 (N_8973,N_8866,N_8796);
or U8974 (N_8974,N_8754,N_8837);
and U8975 (N_8975,N_8869,N_8763);
xor U8976 (N_8976,N_8833,N_8811);
nor U8977 (N_8977,N_8753,N_8868);
and U8978 (N_8978,N_8790,N_8820);
nand U8979 (N_8979,N_8831,N_8810);
or U8980 (N_8980,N_8812,N_8816);
or U8981 (N_8981,N_8838,N_8804);
xnor U8982 (N_8982,N_8838,N_8854);
xor U8983 (N_8983,N_8821,N_8785);
or U8984 (N_8984,N_8841,N_8754);
or U8985 (N_8985,N_8872,N_8772);
and U8986 (N_8986,N_8871,N_8803);
nand U8987 (N_8987,N_8819,N_8866);
or U8988 (N_8988,N_8783,N_8763);
xnor U8989 (N_8989,N_8821,N_8801);
nor U8990 (N_8990,N_8791,N_8794);
or U8991 (N_8991,N_8778,N_8770);
or U8992 (N_8992,N_8855,N_8840);
xor U8993 (N_8993,N_8831,N_8811);
nand U8994 (N_8994,N_8761,N_8781);
nor U8995 (N_8995,N_8818,N_8845);
and U8996 (N_8996,N_8802,N_8856);
and U8997 (N_8997,N_8871,N_8850);
or U8998 (N_8998,N_8779,N_8771);
and U8999 (N_8999,N_8873,N_8782);
and U9000 (N_9000,N_8983,N_8946);
nor U9001 (N_9001,N_8933,N_8926);
nand U9002 (N_9002,N_8950,N_8968);
nand U9003 (N_9003,N_8884,N_8994);
nor U9004 (N_9004,N_8931,N_8959);
nor U9005 (N_9005,N_8932,N_8928);
or U9006 (N_9006,N_8992,N_8981);
and U9007 (N_9007,N_8986,N_8875);
or U9008 (N_9008,N_8925,N_8987);
xnor U9009 (N_9009,N_8969,N_8880);
and U9010 (N_9010,N_8977,N_8912);
nand U9011 (N_9011,N_8882,N_8938);
xor U9012 (N_9012,N_8951,N_8988);
and U9013 (N_9013,N_8909,N_8878);
nor U9014 (N_9014,N_8897,N_8887);
nor U9015 (N_9015,N_8900,N_8889);
nand U9016 (N_9016,N_8908,N_8916);
and U9017 (N_9017,N_8965,N_8996);
xor U9018 (N_9018,N_8947,N_8975);
or U9019 (N_9019,N_8901,N_8972);
or U9020 (N_9020,N_8895,N_8924);
or U9021 (N_9021,N_8999,N_8935);
xnor U9022 (N_9022,N_8930,N_8953);
and U9023 (N_9023,N_8963,N_8910);
xor U9024 (N_9024,N_8896,N_8922);
nand U9025 (N_9025,N_8903,N_8890);
and U9026 (N_9026,N_8995,N_8891);
nor U9027 (N_9027,N_8949,N_8905);
xnor U9028 (N_9028,N_8907,N_8985);
nor U9029 (N_9029,N_8979,N_8990);
and U9030 (N_9030,N_8894,N_8964);
nor U9031 (N_9031,N_8940,N_8962);
or U9032 (N_9032,N_8982,N_8956);
and U9033 (N_9033,N_8998,N_8917);
or U9034 (N_9034,N_8958,N_8942);
and U9035 (N_9035,N_8902,N_8923);
and U9036 (N_9036,N_8976,N_8914);
nand U9037 (N_9037,N_8943,N_8920);
and U9038 (N_9038,N_8904,N_8893);
nand U9039 (N_9039,N_8934,N_8973);
and U9040 (N_9040,N_8919,N_8881);
nand U9041 (N_9041,N_8945,N_8974);
or U9042 (N_9042,N_8876,N_8885);
nand U9043 (N_9043,N_8888,N_8921);
and U9044 (N_9044,N_8879,N_8993);
and U9045 (N_9045,N_8948,N_8883);
and U9046 (N_9046,N_8970,N_8997);
nand U9047 (N_9047,N_8991,N_8906);
nand U9048 (N_9048,N_8966,N_8899);
and U9049 (N_9049,N_8941,N_8967);
xor U9050 (N_9050,N_8961,N_8937);
xnor U9051 (N_9051,N_8978,N_8944);
xnor U9052 (N_9052,N_8911,N_8955);
and U9053 (N_9053,N_8952,N_8989);
nor U9054 (N_9054,N_8898,N_8980);
nand U9055 (N_9055,N_8913,N_8971);
xnor U9056 (N_9056,N_8886,N_8927);
nor U9057 (N_9057,N_8936,N_8954);
or U9058 (N_9058,N_8918,N_8877);
or U9059 (N_9059,N_8957,N_8984);
or U9060 (N_9060,N_8960,N_8929);
xor U9061 (N_9061,N_8892,N_8915);
nor U9062 (N_9062,N_8939,N_8913);
nand U9063 (N_9063,N_8943,N_8919);
xnor U9064 (N_9064,N_8986,N_8927);
xnor U9065 (N_9065,N_8984,N_8926);
nor U9066 (N_9066,N_8889,N_8962);
nor U9067 (N_9067,N_8981,N_8963);
nand U9068 (N_9068,N_8958,N_8970);
xor U9069 (N_9069,N_8984,N_8928);
and U9070 (N_9070,N_8990,N_8948);
or U9071 (N_9071,N_8935,N_8957);
xor U9072 (N_9072,N_8980,N_8951);
nor U9073 (N_9073,N_8972,N_8903);
xor U9074 (N_9074,N_8988,N_8912);
nand U9075 (N_9075,N_8997,N_8950);
nor U9076 (N_9076,N_8925,N_8927);
nor U9077 (N_9077,N_8945,N_8910);
nand U9078 (N_9078,N_8998,N_8883);
nand U9079 (N_9079,N_8974,N_8994);
nor U9080 (N_9080,N_8943,N_8964);
and U9081 (N_9081,N_8968,N_8913);
nand U9082 (N_9082,N_8892,N_8980);
and U9083 (N_9083,N_8902,N_8907);
or U9084 (N_9084,N_8940,N_8967);
or U9085 (N_9085,N_8998,N_8905);
xor U9086 (N_9086,N_8951,N_8981);
and U9087 (N_9087,N_8980,N_8903);
nand U9088 (N_9088,N_8878,N_8939);
nor U9089 (N_9089,N_8945,N_8952);
and U9090 (N_9090,N_8895,N_8920);
and U9091 (N_9091,N_8962,N_8935);
nand U9092 (N_9092,N_8940,N_8928);
xor U9093 (N_9093,N_8889,N_8953);
nor U9094 (N_9094,N_8936,N_8956);
nor U9095 (N_9095,N_8929,N_8943);
and U9096 (N_9096,N_8944,N_8888);
nor U9097 (N_9097,N_8947,N_8991);
nand U9098 (N_9098,N_8927,N_8939);
and U9099 (N_9099,N_8896,N_8888);
xor U9100 (N_9100,N_8943,N_8991);
and U9101 (N_9101,N_8955,N_8977);
or U9102 (N_9102,N_8946,N_8922);
nor U9103 (N_9103,N_8943,N_8899);
nor U9104 (N_9104,N_8881,N_8928);
nor U9105 (N_9105,N_8930,N_8983);
or U9106 (N_9106,N_8910,N_8958);
xnor U9107 (N_9107,N_8961,N_8900);
and U9108 (N_9108,N_8956,N_8893);
or U9109 (N_9109,N_8889,N_8880);
or U9110 (N_9110,N_8907,N_8893);
nor U9111 (N_9111,N_8977,N_8922);
nand U9112 (N_9112,N_8972,N_8919);
or U9113 (N_9113,N_8929,N_8996);
nand U9114 (N_9114,N_8900,N_8875);
nand U9115 (N_9115,N_8922,N_8945);
and U9116 (N_9116,N_8897,N_8963);
and U9117 (N_9117,N_8949,N_8895);
or U9118 (N_9118,N_8989,N_8906);
or U9119 (N_9119,N_8919,N_8975);
nand U9120 (N_9120,N_8936,N_8879);
xor U9121 (N_9121,N_8886,N_8976);
nand U9122 (N_9122,N_8961,N_8943);
nand U9123 (N_9123,N_8929,N_8877);
nor U9124 (N_9124,N_8987,N_8956);
nor U9125 (N_9125,N_9020,N_9082);
or U9126 (N_9126,N_9030,N_9045);
or U9127 (N_9127,N_9034,N_9063);
nand U9128 (N_9128,N_9021,N_9038);
or U9129 (N_9129,N_9015,N_9031);
xnor U9130 (N_9130,N_9016,N_9035);
nand U9131 (N_9131,N_9053,N_9047);
xor U9132 (N_9132,N_9105,N_9056);
nand U9133 (N_9133,N_9076,N_9033);
xor U9134 (N_9134,N_9075,N_9026);
nand U9135 (N_9135,N_9064,N_9072);
and U9136 (N_9136,N_9012,N_9050);
xnor U9137 (N_9137,N_9115,N_9058);
or U9138 (N_9138,N_9117,N_9089);
and U9139 (N_9139,N_9057,N_9087);
xnor U9140 (N_9140,N_9044,N_9084);
and U9141 (N_9141,N_9039,N_9046);
and U9142 (N_9142,N_9043,N_9060);
or U9143 (N_9143,N_9019,N_9013);
nand U9144 (N_9144,N_9002,N_9065);
or U9145 (N_9145,N_9118,N_9003);
or U9146 (N_9146,N_9023,N_9024);
xor U9147 (N_9147,N_9018,N_9054);
xor U9148 (N_9148,N_9109,N_9107);
or U9149 (N_9149,N_9102,N_9069);
nor U9150 (N_9150,N_9055,N_9011);
nand U9151 (N_9151,N_9093,N_9124);
nor U9152 (N_9152,N_9088,N_9108);
nor U9153 (N_9153,N_9014,N_9000);
and U9154 (N_9154,N_9008,N_9101);
nor U9155 (N_9155,N_9032,N_9073);
xnor U9156 (N_9156,N_9027,N_9001);
xor U9157 (N_9157,N_9048,N_9009);
nor U9158 (N_9158,N_9096,N_9120);
and U9159 (N_9159,N_9114,N_9071);
and U9160 (N_9160,N_9099,N_9067);
xnor U9161 (N_9161,N_9110,N_9095);
or U9162 (N_9162,N_9051,N_9037);
nand U9163 (N_9163,N_9116,N_9103);
xor U9164 (N_9164,N_9061,N_9070);
or U9165 (N_9165,N_9074,N_9104);
nand U9166 (N_9166,N_9005,N_9052);
nand U9167 (N_9167,N_9007,N_9017);
or U9168 (N_9168,N_9097,N_9111);
xnor U9169 (N_9169,N_9041,N_9029);
nand U9170 (N_9170,N_9022,N_9006);
nand U9171 (N_9171,N_9123,N_9004);
nand U9172 (N_9172,N_9085,N_9025);
or U9173 (N_9173,N_9091,N_9113);
xnor U9174 (N_9174,N_9079,N_9121);
nor U9175 (N_9175,N_9078,N_9098);
xor U9176 (N_9176,N_9010,N_9092);
nor U9177 (N_9177,N_9059,N_9106);
xor U9178 (N_9178,N_9062,N_9112);
xor U9179 (N_9179,N_9081,N_9094);
or U9180 (N_9180,N_9040,N_9049);
or U9181 (N_9181,N_9036,N_9090);
nand U9182 (N_9182,N_9042,N_9100);
nand U9183 (N_9183,N_9122,N_9066);
or U9184 (N_9184,N_9080,N_9083);
or U9185 (N_9185,N_9086,N_9028);
and U9186 (N_9186,N_9068,N_9119);
and U9187 (N_9187,N_9077,N_9085);
xor U9188 (N_9188,N_9068,N_9093);
or U9189 (N_9189,N_9011,N_9087);
and U9190 (N_9190,N_9123,N_9083);
xnor U9191 (N_9191,N_9062,N_9048);
and U9192 (N_9192,N_9010,N_9038);
and U9193 (N_9193,N_9061,N_9096);
or U9194 (N_9194,N_9114,N_9110);
and U9195 (N_9195,N_9091,N_9061);
nand U9196 (N_9196,N_9014,N_9068);
and U9197 (N_9197,N_9073,N_9065);
nand U9198 (N_9198,N_9002,N_9067);
nor U9199 (N_9199,N_9003,N_9082);
and U9200 (N_9200,N_9021,N_9041);
or U9201 (N_9201,N_9087,N_9020);
nand U9202 (N_9202,N_9108,N_9052);
nand U9203 (N_9203,N_9053,N_9064);
xor U9204 (N_9204,N_9087,N_9016);
nor U9205 (N_9205,N_9102,N_9055);
nor U9206 (N_9206,N_9114,N_9056);
nand U9207 (N_9207,N_9104,N_9025);
or U9208 (N_9208,N_9090,N_9050);
and U9209 (N_9209,N_9120,N_9097);
nand U9210 (N_9210,N_9119,N_9115);
nor U9211 (N_9211,N_9082,N_9113);
or U9212 (N_9212,N_9102,N_9043);
nor U9213 (N_9213,N_9089,N_9096);
nor U9214 (N_9214,N_9044,N_9011);
nor U9215 (N_9215,N_9110,N_9046);
nand U9216 (N_9216,N_9091,N_9079);
nand U9217 (N_9217,N_9094,N_9031);
nor U9218 (N_9218,N_9078,N_9103);
or U9219 (N_9219,N_9018,N_9067);
and U9220 (N_9220,N_9073,N_9066);
or U9221 (N_9221,N_9074,N_9032);
and U9222 (N_9222,N_9024,N_9100);
xnor U9223 (N_9223,N_9020,N_9073);
and U9224 (N_9224,N_9114,N_9018);
or U9225 (N_9225,N_9020,N_9055);
nand U9226 (N_9226,N_9068,N_9017);
and U9227 (N_9227,N_9089,N_9056);
and U9228 (N_9228,N_9107,N_9073);
nand U9229 (N_9229,N_9039,N_9111);
or U9230 (N_9230,N_9000,N_9019);
nand U9231 (N_9231,N_9082,N_9083);
nor U9232 (N_9232,N_9068,N_9079);
nand U9233 (N_9233,N_9027,N_9051);
or U9234 (N_9234,N_9053,N_9049);
nor U9235 (N_9235,N_9032,N_9028);
nand U9236 (N_9236,N_9070,N_9000);
nor U9237 (N_9237,N_9082,N_9061);
nand U9238 (N_9238,N_9084,N_9015);
or U9239 (N_9239,N_9083,N_9113);
or U9240 (N_9240,N_9022,N_9038);
or U9241 (N_9241,N_9119,N_9071);
xnor U9242 (N_9242,N_9075,N_9046);
and U9243 (N_9243,N_9049,N_9026);
nor U9244 (N_9244,N_9064,N_9108);
nor U9245 (N_9245,N_9099,N_9022);
and U9246 (N_9246,N_9045,N_9041);
nor U9247 (N_9247,N_9061,N_9102);
xor U9248 (N_9248,N_9060,N_9109);
nor U9249 (N_9249,N_9066,N_9008);
and U9250 (N_9250,N_9240,N_9164);
nand U9251 (N_9251,N_9184,N_9125);
or U9252 (N_9252,N_9201,N_9220);
and U9253 (N_9253,N_9152,N_9185);
or U9254 (N_9254,N_9157,N_9215);
nor U9255 (N_9255,N_9190,N_9237);
nor U9256 (N_9256,N_9169,N_9198);
nor U9257 (N_9257,N_9158,N_9143);
and U9258 (N_9258,N_9219,N_9228);
or U9259 (N_9259,N_9170,N_9168);
nor U9260 (N_9260,N_9167,N_9239);
nor U9261 (N_9261,N_9178,N_9223);
nand U9262 (N_9262,N_9249,N_9133);
nand U9263 (N_9263,N_9221,N_9243);
nand U9264 (N_9264,N_9236,N_9216);
xor U9265 (N_9265,N_9138,N_9166);
nor U9266 (N_9266,N_9230,N_9224);
xnor U9267 (N_9267,N_9132,N_9245);
xor U9268 (N_9268,N_9146,N_9229);
xor U9269 (N_9269,N_9244,N_9179);
and U9270 (N_9270,N_9202,N_9234);
xor U9271 (N_9271,N_9214,N_9130);
nand U9272 (N_9272,N_9218,N_9210);
xnor U9273 (N_9273,N_9145,N_9144);
or U9274 (N_9274,N_9128,N_9196);
nor U9275 (N_9275,N_9209,N_9232);
or U9276 (N_9276,N_9174,N_9187);
xnor U9277 (N_9277,N_9242,N_9199);
nand U9278 (N_9278,N_9137,N_9127);
and U9279 (N_9279,N_9172,N_9197);
nor U9280 (N_9280,N_9177,N_9246);
nor U9281 (N_9281,N_9212,N_9171);
xnor U9282 (N_9282,N_9183,N_9135);
xnor U9283 (N_9283,N_9182,N_9142);
nand U9284 (N_9284,N_9238,N_9227);
nand U9285 (N_9285,N_9225,N_9141);
xor U9286 (N_9286,N_9213,N_9233);
and U9287 (N_9287,N_9247,N_9159);
or U9288 (N_9288,N_9206,N_9153);
nand U9289 (N_9289,N_9139,N_9150);
or U9290 (N_9290,N_9160,N_9189);
nand U9291 (N_9291,N_9226,N_9200);
nand U9292 (N_9292,N_9241,N_9235);
xor U9293 (N_9293,N_9165,N_9186);
nor U9294 (N_9294,N_9175,N_9161);
nand U9295 (N_9295,N_9149,N_9194);
or U9296 (N_9296,N_9148,N_9173);
nor U9297 (N_9297,N_9231,N_9151);
xor U9298 (N_9298,N_9195,N_9140);
nand U9299 (N_9299,N_9188,N_9136);
or U9300 (N_9300,N_9131,N_9181);
and U9301 (N_9301,N_9207,N_9162);
or U9302 (N_9302,N_9193,N_9147);
or U9303 (N_9303,N_9203,N_9156);
or U9304 (N_9304,N_9208,N_9126);
or U9305 (N_9305,N_9129,N_9180);
or U9306 (N_9306,N_9211,N_9222);
nand U9307 (N_9307,N_9154,N_9217);
or U9308 (N_9308,N_9205,N_9163);
and U9309 (N_9309,N_9248,N_9155);
nor U9310 (N_9310,N_9192,N_9134);
nand U9311 (N_9311,N_9204,N_9191);
nand U9312 (N_9312,N_9176,N_9159);
xnor U9313 (N_9313,N_9157,N_9176);
nand U9314 (N_9314,N_9201,N_9133);
xnor U9315 (N_9315,N_9166,N_9211);
nor U9316 (N_9316,N_9212,N_9135);
xnor U9317 (N_9317,N_9191,N_9240);
nor U9318 (N_9318,N_9232,N_9162);
or U9319 (N_9319,N_9249,N_9199);
and U9320 (N_9320,N_9238,N_9249);
and U9321 (N_9321,N_9186,N_9227);
or U9322 (N_9322,N_9194,N_9180);
and U9323 (N_9323,N_9200,N_9153);
or U9324 (N_9324,N_9162,N_9150);
nor U9325 (N_9325,N_9219,N_9216);
xnor U9326 (N_9326,N_9181,N_9177);
or U9327 (N_9327,N_9210,N_9242);
or U9328 (N_9328,N_9199,N_9243);
nor U9329 (N_9329,N_9244,N_9191);
xnor U9330 (N_9330,N_9226,N_9180);
nor U9331 (N_9331,N_9232,N_9140);
or U9332 (N_9332,N_9176,N_9132);
nor U9333 (N_9333,N_9177,N_9210);
nor U9334 (N_9334,N_9239,N_9205);
xnor U9335 (N_9335,N_9149,N_9135);
and U9336 (N_9336,N_9246,N_9143);
and U9337 (N_9337,N_9232,N_9188);
xnor U9338 (N_9338,N_9249,N_9134);
or U9339 (N_9339,N_9139,N_9221);
nor U9340 (N_9340,N_9160,N_9134);
or U9341 (N_9341,N_9165,N_9143);
nor U9342 (N_9342,N_9226,N_9199);
or U9343 (N_9343,N_9126,N_9147);
or U9344 (N_9344,N_9192,N_9129);
and U9345 (N_9345,N_9210,N_9205);
nand U9346 (N_9346,N_9233,N_9189);
nand U9347 (N_9347,N_9159,N_9131);
or U9348 (N_9348,N_9147,N_9196);
nand U9349 (N_9349,N_9216,N_9201);
and U9350 (N_9350,N_9141,N_9240);
nand U9351 (N_9351,N_9202,N_9228);
nor U9352 (N_9352,N_9202,N_9127);
nand U9353 (N_9353,N_9171,N_9188);
and U9354 (N_9354,N_9245,N_9229);
or U9355 (N_9355,N_9248,N_9138);
nor U9356 (N_9356,N_9187,N_9217);
and U9357 (N_9357,N_9241,N_9168);
and U9358 (N_9358,N_9232,N_9230);
xnor U9359 (N_9359,N_9201,N_9129);
or U9360 (N_9360,N_9185,N_9199);
or U9361 (N_9361,N_9236,N_9228);
xnor U9362 (N_9362,N_9230,N_9211);
nor U9363 (N_9363,N_9174,N_9235);
nand U9364 (N_9364,N_9173,N_9198);
xnor U9365 (N_9365,N_9233,N_9156);
nand U9366 (N_9366,N_9173,N_9177);
or U9367 (N_9367,N_9167,N_9166);
or U9368 (N_9368,N_9210,N_9195);
or U9369 (N_9369,N_9214,N_9180);
nand U9370 (N_9370,N_9157,N_9128);
nand U9371 (N_9371,N_9161,N_9184);
nor U9372 (N_9372,N_9185,N_9184);
nand U9373 (N_9373,N_9185,N_9131);
nand U9374 (N_9374,N_9241,N_9195);
and U9375 (N_9375,N_9330,N_9307);
nor U9376 (N_9376,N_9251,N_9349);
or U9377 (N_9377,N_9355,N_9354);
nor U9378 (N_9378,N_9259,N_9341);
nor U9379 (N_9379,N_9266,N_9369);
nand U9380 (N_9380,N_9284,N_9345);
nor U9381 (N_9381,N_9253,N_9320);
xor U9382 (N_9382,N_9256,N_9250);
or U9383 (N_9383,N_9263,N_9276);
nor U9384 (N_9384,N_9267,N_9321);
nor U9385 (N_9385,N_9370,N_9372);
and U9386 (N_9386,N_9337,N_9306);
xnor U9387 (N_9387,N_9353,N_9310);
or U9388 (N_9388,N_9347,N_9314);
xnor U9389 (N_9389,N_9297,N_9368);
nand U9390 (N_9390,N_9287,N_9364);
and U9391 (N_9391,N_9277,N_9329);
or U9392 (N_9392,N_9301,N_9346);
or U9393 (N_9393,N_9294,N_9374);
or U9394 (N_9394,N_9289,N_9336);
and U9395 (N_9395,N_9325,N_9268);
and U9396 (N_9396,N_9254,N_9296);
nor U9397 (N_9397,N_9282,N_9285);
or U9398 (N_9398,N_9357,N_9308);
and U9399 (N_9399,N_9290,N_9270);
or U9400 (N_9400,N_9313,N_9316);
nand U9401 (N_9401,N_9309,N_9324);
nor U9402 (N_9402,N_9286,N_9359);
xor U9403 (N_9403,N_9302,N_9255);
nand U9404 (N_9404,N_9257,N_9319);
xor U9405 (N_9405,N_9366,N_9252);
nand U9406 (N_9406,N_9315,N_9305);
nand U9407 (N_9407,N_9356,N_9279);
nand U9408 (N_9408,N_9258,N_9326);
xor U9409 (N_9409,N_9274,N_9333);
xor U9410 (N_9410,N_9339,N_9318);
xor U9411 (N_9411,N_9265,N_9311);
or U9412 (N_9412,N_9292,N_9362);
and U9413 (N_9413,N_9343,N_9262);
and U9414 (N_9414,N_9360,N_9334);
and U9415 (N_9415,N_9298,N_9338);
nand U9416 (N_9416,N_9342,N_9352);
nand U9417 (N_9417,N_9280,N_9300);
and U9418 (N_9418,N_9273,N_9335);
xor U9419 (N_9419,N_9312,N_9281);
xnor U9420 (N_9420,N_9348,N_9367);
nand U9421 (N_9421,N_9328,N_9295);
xnor U9422 (N_9422,N_9340,N_9304);
nor U9423 (N_9423,N_9269,N_9291);
and U9424 (N_9424,N_9371,N_9283);
and U9425 (N_9425,N_9288,N_9327);
or U9426 (N_9426,N_9299,N_9363);
or U9427 (N_9427,N_9261,N_9260);
and U9428 (N_9428,N_9365,N_9358);
nor U9429 (N_9429,N_9293,N_9332);
xnor U9430 (N_9430,N_9272,N_9271);
nand U9431 (N_9431,N_9322,N_9323);
and U9432 (N_9432,N_9317,N_9373);
nand U9433 (N_9433,N_9275,N_9303);
nor U9434 (N_9434,N_9264,N_9344);
xnor U9435 (N_9435,N_9361,N_9351);
xnor U9436 (N_9436,N_9350,N_9278);
and U9437 (N_9437,N_9331,N_9314);
or U9438 (N_9438,N_9269,N_9363);
or U9439 (N_9439,N_9276,N_9301);
nand U9440 (N_9440,N_9346,N_9335);
or U9441 (N_9441,N_9290,N_9338);
nor U9442 (N_9442,N_9302,N_9298);
xor U9443 (N_9443,N_9286,N_9318);
nor U9444 (N_9444,N_9269,N_9271);
nor U9445 (N_9445,N_9297,N_9283);
or U9446 (N_9446,N_9251,N_9282);
xor U9447 (N_9447,N_9352,N_9346);
or U9448 (N_9448,N_9311,N_9328);
nand U9449 (N_9449,N_9273,N_9272);
and U9450 (N_9450,N_9361,N_9330);
nand U9451 (N_9451,N_9372,N_9371);
xnor U9452 (N_9452,N_9311,N_9363);
or U9453 (N_9453,N_9335,N_9325);
and U9454 (N_9454,N_9314,N_9272);
or U9455 (N_9455,N_9303,N_9326);
nor U9456 (N_9456,N_9352,N_9298);
and U9457 (N_9457,N_9326,N_9264);
and U9458 (N_9458,N_9355,N_9258);
xnor U9459 (N_9459,N_9336,N_9293);
nor U9460 (N_9460,N_9342,N_9274);
and U9461 (N_9461,N_9303,N_9355);
nand U9462 (N_9462,N_9360,N_9259);
nand U9463 (N_9463,N_9366,N_9362);
nand U9464 (N_9464,N_9274,N_9358);
or U9465 (N_9465,N_9357,N_9342);
xnor U9466 (N_9466,N_9328,N_9286);
xor U9467 (N_9467,N_9317,N_9294);
xnor U9468 (N_9468,N_9370,N_9274);
nor U9469 (N_9469,N_9305,N_9369);
nor U9470 (N_9470,N_9283,N_9337);
nand U9471 (N_9471,N_9318,N_9366);
nor U9472 (N_9472,N_9350,N_9253);
nor U9473 (N_9473,N_9341,N_9263);
nand U9474 (N_9474,N_9362,N_9348);
xnor U9475 (N_9475,N_9285,N_9362);
and U9476 (N_9476,N_9273,N_9365);
xnor U9477 (N_9477,N_9288,N_9351);
nand U9478 (N_9478,N_9343,N_9307);
or U9479 (N_9479,N_9297,N_9360);
and U9480 (N_9480,N_9359,N_9351);
and U9481 (N_9481,N_9287,N_9358);
xor U9482 (N_9482,N_9325,N_9259);
nand U9483 (N_9483,N_9354,N_9282);
nand U9484 (N_9484,N_9326,N_9351);
or U9485 (N_9485,N_9260,N_9299);
nand U9486 (N_9486,N_9260,N_9300);
nand U9487 (N_9487,N_9300,N_9262);
xnor U9488 (N_9488,N_9297,N_9319);
nand U9489 (N_9489,N_9285,N_9365);
nand U9490 (N_9490,N_9286,N_9270);
xor U9491 (N_9491,N_9298,N_9324);
nand U9492 (N_9492,N_9369,N_9278);
nor U9493 (N_9493,N_9296,N_9337);
xor U9494 (N_9494,N_9272,N_9323);
or U9495 (N_9495,N_9343,N_9269);
nor U9496 (N_9496,N_9263,N_9261);
or U9497 (N_9497,N_9315,N_9304);
nor U9498 (N_9498,N_9278,N_9308);
nor U9499 (N_9499,N_9306,N_9286);
nor U9500 (N_9500,N_9422,N_9397);
or U9501 (N_9501,N_9448,N_9403);
and U9502 (N_9502,N_9474,N_9480);
nand U9503 (N_9503,N_9426,N_9447);
nor U9504 (N_9504,N_9491,N_9445);
nand U9505 (N_9505,N_9468,N_9453);
xnor U9506 (N_9506,N_9395,N_9462);
xor U9507 (N_9507,N_9377,N_9458);
and U9508 (N_9508,N_9467,N_9452);
and U9509 (N_9509,N_9443,N_9384);
or U9510 (N_9510,N_9483,N_9425);
nand U9511 (N_9511,N_9407,N_9489);
nand U9512 (N_9512,N_9406,N_9411);
or U9513 (N_9513,N_9488,N_9424);
nand U9514 (N_9514,N_9444,N_9461);
nand U9515 (N_9515,N_9439,N_9446);
nand U9516 (N_9516,N_9393,N_9460);
nor U9517 (N_9517,N_9434,N_9451);
nand U9518 (N_9518,N_9404,N_9482);
xnor U9519 (N_9519,N_9497,N_9389);
or U9520 (N_9520,N_9398,N_9490);
or U9521 (N_9521,N_9429,N_9402);
nand U9522 (N_9522,N_9382,N_9401);
and U9523 (N_9523,N_9437,N_9400);
xor U9524 (N_9524,N_9463,N_9486);
xnor U9525 (N_9525,N_9477,N_9387);
or U9526 (N_9526,N_9427,N_9469);
xnor U9527 (N_9527,N_9376,N_9423);
nor U9528 (N_9528,N_9476,N_9432);
xor U9529 (N_9529,N_9433,N_9388);
or U9530 (N_9530,N_9380,N_9484);
or U9531 (N_9531,N_9485,N_9405);
nand U9532 (N_9532,N_9464,N_9492);
nor U9533 (N_9533,N_9396,N_9441);
nand U9534 (N_9534,N_9494,N_9392);
nor U9535 (N_9535,N_9410,N_9412);
and U9536 (N_9536,N_9436,N_9449);
nor U9537 (N_9537,N_9440,N_9379);
or U9538 (N_9538,N_9390,N_9457);
xnor U9539 (N_9539,N_9495,N_9438);
and U9540 (N_9540,N_9481,N_9408);
and U9541 (N_9541,N_9414,N_9409);
nor U9542 (N_9542,N_9418,N_9416);
xnor U9543 (N_9543,N_9394,N_9435);
or U9544 (N_9544,N_9378,N_9470);
nor U9545 (N_9545,N_9466,N_9442);
nand U9546 (N_9546,N_9385,N_9454);
and U9547 (N_9547,N_9456,N_9383);
xnor U9548 (N_9548,N_9493,N_9498);
or U9549 (N_9549,N_9421,N_9450);
and U9550 (N_9550,N_9487,N_9399);
nand U9551 (N_9551,N_9428,N_9459);
or U9552 (N_9552,N_9472,N_9465);
nand U9553 (N_9553,N_9413,N_9417);
and U9554 (N_9554,N_9381,N_9386);
or U9555 (N_9555,N_9471,N_9473);
nor U9556 (N_9556,N_9431,N_9496);
nand U9557 (N_9557,N_9419,N_9455);
xnor U9558 (N_9558,N_9499,N_9479);
nand U9559 (N_9559,N_9430,N_9475);
nand U9560 (N_9560,N_9375,N_9478);
nor U9561 (N_9561,N_9391,N_9415);
xnor U9562 (N_9562,N_9420,N_9381);
xor U9563 (N_9563,N_9425,N_9479);
nor U9564 (N_9564,N_9491,N_9401);
xnor U9565 (N_9565,N_9376,N_9389);
nand U9566 (N_9566,N_9431,N_9421);
xor U9567 (N_9567,N_9387,N_9447);
and U9568 (N_9568,N_9460,N_9411);
nand U9569 (N_9569,N_9430,N_9480);
and U9570 (N_9570,N_9408,N_9412);
nor U9571 (N_9571,N_9427,N_9390);
and U9572 (N_9572,N_9395,N_9447);
xor U9573 (N_9573,N_9427,N_9400);
and U9574 (N_9574,N_9461,N_9471);
and U9575 (N_9575,N_9440,N_9452);
and U9576 (N_9576,N_9480,N_9389);
nand U9577 (N_9577,N_9400,N_9472);
or U9578 (N_9578,N_9388,N_9427);
xor U9579 (N_9579,N_9430,N_9443);
or U9580 (N_9580,N_9467,N_9458);
and U9581 (N_9581,N_9467,N_9498);
nor U9582 (N_9582,N_9401,N_9438);
nand U9583 (N_9583,N_9474,N_9499);
or U9584 (N_9584,N_9415,N_9426);
xnor U9585 (N_9585,N_9405,N_9491);
nand U9586 (N_9586,N_9428,N_9470);
or U9587 (N_9587,N_9405,N_9447);
xnor U9588 (N_9588,N_9428,N_9437);
and U9589 (N_9589,N_9451,N_9408);
xnor U9590 (N_9590,N_9452,N_9455);
nor U9591 (N_9591,N_9400,N_9446);
nand U9592 (N_9592,N_9460,N_9492);
nand U9593 (N_9593,N_9471,N_9397);
xor U9594 (N_9594,N_9493,N_9390);
xor U9595 (N_9595,N_9395,N_9446);
and U9596 (N_9596,N_9477,N_9407);
and U9597 (N_9597,N_9413,N_9390);
nor U9598 (N_9598,N_9423,N_9451);
nand U9599 (N_9599,N_9423,N_9396);
xor U9600 (N_9600,N_9468,N_9490);
nand U9601 (N_9601,N_9481,N_9485);
xor U9602 (N_9602,N_9403,N_9493);
nand U9603 (N_9603,N_9489,N_9404);
nand U9604 (N_9604,N_9461,N_9460);
nor U9605 (N_9605,N_9454,N_9457);
nor U9606 (N_9606,N_9475,N_9482);
and U9607 (N_9607,N_9390,N_9417);
xor U9608 (N_9608,N_9405,N_9444);
and U9609 (N_9609,N_9498,N_9457);
xnor U9610 (N_9610,N_9423,N_9433);
or U9611 (N_9611,N_9442,N_9389);
or U9612 (N_9612,N_9388,N_9496);
xnor U9613 (N_9613,N_9382,N_9395);
and U9614 (N_9614,N_9481,N_9439);
or U9615 (N_9615,N_9489,N_9434);
or U9616 (N_9616,N_9396,N_9424);
and U9617 (N_9617,N_9428,N_9406);
and U9618 (N_9618,N_9389,N_9434);
and U9619 (N_9619,N_9384,N_9387);
nor U9620 (N_9620,N_9456,N_9422);
xor U9621 (N_9621,N_9459,N_9427);
xnor U9622 (N_9622,N_9457,N_9389);
or U9623 (N_9623,N_9414,N_9441);
nand U9624 (N_9624,N_9483,N_9487);
nor U9625 (N_9625,N_9559,N_9603);
nor U9626 (N_9626,N_9565,N_9579);
xnor U9627 (N_9627,N_9550,N_9518);
or U9628 (N_9628,N_9569,N_9501);
nand U9629 (N_9629,N_9529,N_9584);
nand U9630 (N_9630,N_9548,N_9554);
nand U9631 (N_9631,N_9562,N_9618);
nand U9632 (N_9632,N_9553,N_9524);
or U9633 (N_9633,N_9564,N_9536);
xnor U9634 (N_9634,N_9511,N_9571);
nor U9635 (N_9635,N_9600,N_9598);
xnor U9636 (N_9636,N_9523,N_9602);
nor U9637 (N_9637,N_9522,N_9599);
nor U9638 (N_9638,N_9560,N_9503);
or U9639 (N_9639,N_9541,N_9509);
xor U9640 (N_9640,N_9581,N_9596);
nor U9641 (N_9641,N_9537,N_9516);
and U9642 (N_9642,N_9556,N_9543);
and U9643 (N_9643,N_9594,N_9587);
nand U9644 (N_9644,N_9610,N_9577);
nand U9645 (N_9645,N_9613,N_9586);
xnor U9646 (N_9646,N_9542,N_9604);
and U9647 (N_9647,N_9614,N_9580);
nand U9648 (N_9648,N_9526,N_9510);
and U9649 (N_9649,N_9558,N_9615);
or U9650 (N_9650,N_9578,N_9551);
and U9651 (N_9651,N_9525,N_9534);
nor U9652 (N_9652,N_9530,N_9532);
and U9653 (N_9653,N_9607,N_9561);
and U9654 (N_9654,N_9620,N_9505);
nor U9655 (N_9655,N_9549,N_9521);
nand U9656 (N_9656,N_9612,N_9591);
nor U9657 (N_9657,N_9616,N_9544);
and U9658 (N_9658,N_9570,N_9504);
and U9659 (N_9659,N_9506,N_9502);
and U9660 (N_9660,N_9514,N_9508);
nand U9661 (N_9661,N_9590,N_9546);
nand U9662 (N_9662,N_9621,N_9573);
nor U9663 (N_9663,N_9585,N_9545);
xnor U9664 (N_9664,N_9531,N_9513);
nor U9665 (N_9665,N_9609,N_9608);
xnor U9666 (N_9666,N_9540,N_9572);
and U9667 (N_9667,N_9617,N_9528);
nor U9668 (N_9668,N_9619,N_9563);
and U9669 (N_9669,N_9500,N_9533);
nand U9670 (N_9670,N_9595,N_9519);
nor U9671 (N_9671,N_9539,N_9605);
or U9672 (N_9672,N_9538,N_9622);
nor U9673 (N_9673,N_9606,N_9588);
xor U9674 (N_9674,N_9515,N_9583);
nand U9675 (N_9675,N_9623,N_9566);
xnor U9676 (N_9676,N_9517,N_9557);
xnor U9677 (N_9677,N_9611,N_9597);
and U9678 (N_9678,N_9527,N_9574);
nand U9679 (N_9679,N_9601,N_9576);
or U9680 (N_9680,N_9592,N_9555);
or U9681 (N_9681,N_9575,N_9624);
nand U9682 (N_9682,N_9582,N_9520);
and U9683 (N_9683,N_9567,N_9568);
nand U9684 (N_9684,N_9547,N_9535);
and U9685 (N_9685,N_9512,N_9589);
nand U9686 (N_9686,N_9552,N_9507);
nand U9687 (N_9687,N_9593,N_9602);
nor U9688 (N_9688,N_9502,N_9513);
nor U9689 (N_9689,N_9614,N_9567);
nor U9690 (N_9690,N_9500,N_9514);
nand U9691 (N_9691,N_9574,N_9544);
nor U9692 (N_9692,N_9623,N_9621);
and U9693 (N_9693,N_9571,N_9594);
or U9694 (N_9694,N_9537,N_9551);
nor U9695 (N_9695,N_9523,N_9541);
xor U9696 (N_9696,N_9589,N_9581);
nand U9697 (N_9697,N_9561,N_9580);
nor U9698 (N_9698,N_9569,N_9601);
xor U9699 (N_9699,N_9609,N_9597);
xor U9700 (N_9700,N_9624,N_9508);
or U9701 (N_9701,N_9567,N_9584);
nor U9702 (N_9702,N_9510,N_9580);
nand U9703 (N_9703,N_9507,N_9564);
nor U9704 (N_9704,N_9517,N_9511);
xor U9705 (N_9705,N_9534,N_9502);
and U9706 (N_9706,N_9589,N_9502);
and U9707 (N_9707,N_9578,N_9544);
and U9708 (N_9708,N_9558,N_9574);
or U9709 (N_9709,N_9622,N_9558);
nand U9710 (N_9710,N_9570,N_9513);
xnor U9711 (N_9711,N_9613,N_9587);
nand U9712 (N_9712,N_9545,N_9509);
nor U9713 (N_9713,N_9527,N_9618);
or U9714 (N_9714,N_9532,N_9515);
xor U9715 (N_9715,N_9579,N_9548);
xnor U9716 (N_9716,N_9502,N_9501);
and U9717 (N_9717,N_9591,N_9596);
and U9718 (N_9718,N_9598,N_9623);
xor U9719 (N_9719,N_9548,N_9591);
xor U9720 (N_9720,N_9595,N_9508);
nand U9721 (N_9721,N_9576,N_9532);
nand U9722 (N_9722,N_9504,N_9538);
nand U9723 (N_9723,N_9504,N_9605);
or U9724 (N_9724,N_9620,N_9603);
xnor U9725 (N_9725,N_9617,N_9592);
and U9726 (N_9726,N_9578,N_9533);
xor U9727 (N_9727,N_9602,N_9539);
and U9728 (N_9728,N_9612,N_9555);
nand U9729 (N_9729,N_9593,N_9575);
nor U9730 (N_9730,N_9617,N_9500);
nand U9731 (N_9731,N_9547,N_9575);
and U9732 (N_9732,N_9555,N_9533);
nor U9733 (N_9733,N_9543,N_9523);
or U9734 (N_9734,N_9596,N_9576);
and U9735 (N_9735,N_9620,N_9590);
xnor U9736 (N_9736,N_9575,N_9576);
and U9737 (N_9737,N_9593,N_9508);
or U9738 (N_9738,N_9595,N_9613);
nand U9739 (N_9739,N_9506,N_9539);
nand U9740 (N_9740,N_9555,N_9622);
nand U9741 (N_9741,N_9535,N_9601);
nand U9742 (N_9742,N_9587,N_9567);
xor U9743 (N_9743,N_9556,N_9533);
nand U9744 (N_9744,N_9622,N_9613);
nor U9745 (N_9745,N_9527,N_9512);
and U9746 (N_9746,N_9577,N_9509);
or U9747 (N_9747,N_9557,N_9535);
xor U9748 (N_9748,N_9525,N_9603);
xor U9749 (N_9749,N_9598,N_9556);
or U9750 (N_9750,N_9707,N_9635);
nor U9751 (N_9751,N_9680,N_9712);
nand U9752 (N_9752,N_9702,N_9718);
nor U9753 (N_9753,N_9634,N_9628);
xor U9754 (N_9754,N_9721,N_9661);
nand U9755 (N_9755,N_9650,N_9703);
nor U9756 (N_9756,N_9639,N_9709);
and U9757 (N_9757,N_9663,N_9696);
nand U9758 (N_9758,N_9659,N_9726);
nand U9759 (N_9759,N_9738,N_9694);
or U9760 (N_9760,N_9644,N_9670);
xnor U9761 (N_9761,N_9739,N_9743);
nor U9762 (N_9762,N_9675,N_9677);
or U9763 (N_9763,N_9679,N_9638);
xor U9764 (N_9764,N_9745,N_9686);
xor U9765 (N_9765,N_9626,N_9643);
xnor U9766 (N_9766,N_9632,N_9719);
xnor U9767 (N_9767,N_9735,N_9693);
or U9768 (N_9768,N_9710,N_9630);
nor U9769 (N_9769,N_9681,N_9691);
nand U9770 (N_9770,N_9734,N_9746);
xor U9771 (N_9771,N_9706,N_9683);
or U9772 (N_9772,N_9698,N_9688);
xor U9773 (N_9773,N_9649,N_9676);
and U9774 (N_9774,N_9692,N_9652);
nor U9775 (N_9775,N_9657,N_9722);
or U9776 (N_9776,N_9700,N_9687);
and U9777 (N_9777,N_9662,N_9653);
or U9778 (N_9778,N_9671,N_9715);
or U9779 (N_9779,N_9629,N_9697);
nor U9780 (N_9780,N_9724,N_9747);
or U9781 (N_9781,N_9631,N_9672);
or U9782 (N_9782,N_9725,N_9749);
or U9783 (N_9783,N_9633,N_9723);
xor U9784 (N_9784,N_9741,N_9682);
nand U9785 (N_9785,N_9705,N_9658);
xnor U9786 (N_9786,N_9665,N_9674);
nor U9787 (N_9787,N_9699,N_9711);
or U9788 (N_9788,N_9690,N_9627);
nor U9789 (N_9789,N_9730,N_9654);
or U9790 (N_9790,N_9636,N_9642);
xnor U9791 (N_9791,N_9714,N_9728);
and U9792 (N_9792,N_9742,N_9744);
nor U9793 (N_9793,N_9668,N_9648);
nor U9794 (N_9794,N_9646,N_9736);
nand U9795 (N_9795,N_9647,N_9645);
and U9796 (N_9796,N_9667,N_9732);
or U9797 (N_9797,N_9720,N_9713);
xor U9798 (N_9798,N_9666,N_9717);
nor U9799 (N_9799,N_9673,N_9708);
nand U9800 (N_9800,N_9701,N_9684);
nor U9801 (N_9801,N_9716,N_9641);
and U9802 (N_9802,N_9727,N_9669);
nor U9803 (N_9803,N_9704,N_9655);
or U9804 (N_9804,N_9685,N_9731);
or U9805 (N_9805,N_9656,N_9695);
xnor U9806 (N_9806,N_9729,N_9748);
or U9807 (N_9807,N_9640,N_9740);
nor U9808 (N_9808,N_9660,N_9637);
nor U9809 (N_9809,N_9737,N_9678);
and U9810 (N_9810,N_9651,N_9664);
nor U9811 (N_9811,N_9733,N_9689);
or U9812 (N_9812,N_9625,N_9696);
nor U9813 (N_9813,N_9664,N_9705);
and U9814 (N_9814,N_9668,N_9660);
nor U9815 (N_9815,N_9629,N_9738);
or U9816 (N_9816,N_9743,N_9738);
xor U9817 (N_9817,N_9658,N_9706);
or U9818 (N_9818,N_9728,N_9627);
and U9819 (N_9819,N_9720,N_9642);
xor U9820 (N_9820,N_9748,N_9643);
and U9821 (N_9821,N_9653,N_9698);
or U9822 (N_9822,N_9682,N_9654);
and U9823 (N_9823,N_9643,N_9641);
or U9824 (N_9824,N_9661,N_9714);
xnor U9825 (N_9825,N_9732,N_9656);
and U9826 (N_9826,N_9654,N_9679);
and U9827 (N_9827,N_9662,N_9681);
xor U9828 (N_9828,N_9685,N_9737);
or U9829 (N_9829,N_9636,N_9681);
or U9830 (N_9830,N_9651,N_9643);
xor U9831 (N_9831,N_9666,N_9702);
and U9832 (N_9832,N_9692,N_9658);
xor U9833 (N_9833,N_9749,N_9682);
xor U9834 (N_9834,N_9634,N_9737);
and U9835 (N_9835,N_9658,N_9710);
or U9836 (N_9836,N_9722,N_9645);
nand U9837 (N_9837,N_9748,N_9641);
and U9838 (N_9838,N_9675,N_9740);
nor U9839 (N_9839,N_9652,N_9645);
nand U9840 (N_9840,N_9732,N_9639);
nor U9841 (N_9841,N_9669,N_9728);
nand U9842 (N_9842,N_9740,N_9669);
nor U9843 (N_9843,N_9702,N_9626);
xor U9844 (N_9844,N_9717,N_9706);
and U9845 (N_9845,N_9691,N_9729);
nor U9846 (N_9846,N_9716,N_9628);
or U9847 (N_9847,N_9718,N_9676);
and U9848 (N_9848,N_9741,N_9711);
xnor U9849 (N_9849,N_9660,N_9738);
nor U9850 (N_9850,N_9696,N_9649);
nor U9851 (N_9851,N_9694,N_9720);
nand U9852 (N_9852,N_9707,N_9657);
and U9853 (N_9853,N_9720,N_9626);
and U9854 (N_9854,N_9720,N_9688);
xor U9855 (N_9855,N_9633,N_9630);
xnor U9856 (N_9856,N_9636,N_9643);
and U9857 (N_9857,N_9667,N_9721);
xnor U9858 (N_9858,N_9730,N_9701);
xnor U9859 (N_9859,N_9663,N_9743);
or U9860 (N_9860,N_9705,N_9699);
or U9861 (N_9861,N_9726,N_9708);
or U9862 (N_9862,N_9655,N_9669);
and U9863 (N_9863,N_9695,N_9641);
nand U9864 (N_9864,N_9652,N_9740);
nand U9865 (N_9865,N_9685,N_9702);
and U9866 (N_9866,N_9631,N_9708);
xnor U9867 (N_9867,N_9721,N_9700);
or U9868 (N_9868,N_9713,N_9731);
xor U9869 (N_9869,N_9723,N_9675);
xor U9870 (N_9870,N_9714,N_9700);
nand U9871 (N_9871,N_9726,N_9724);
and U9872 (N_9872,N_9680,N_9637);
or U9873 (N_9873,N_9684,N_9680);
or U9874 (N_9874,N_9737,N_9727);
nor U9875 (N_9875,N_9827,N_9779);
and U9876 (N_9876,N_9801,N_9826);
or U9877 (N_9877,N_9820,N_9770);
xor U9878 (N_9878,N_9864,N_9851);
or U9879 (N_9879,N_9805,N_9856);
xor U9880 (N_9880,N_9857,N_9841);
xor U9881 (N_9881,N_9843,N_9873);
xnor U9882 (N_9882,N_9837,N_9824);
and U9883 (N_9883,N_9798,N_9758);
nor U9884 (N_9884,N_9791,N_9814);
xor U9885 (N_9885,N_9750,N_9800);
and U9886 (N_9886,N_9807,N_9764);
nand U9887 (N_9887,N_9834,N_9753);
and U9888 (N_9888,N_9808,N_9833);
nand U9889 (N_9889,N_9777,N_9810);
xor U9890 (N_9890,N_9793,N_9829);
nor U9891 (N_9891,N_9862,N_9761);
xor U9892 (N_9892,N_9784,N_9803);
nor U9893 (N_9893,N_9760,N_9858);
and U9894 (N_9894,N_9815,N_9774);
or U9895 (N_9895,N_9769,N_9868);
nor U9896 (N_9896,N_9809,N_9786);
nor U9897 (N_9897,N_9783,N_9812);
or U9898 (N_9898,N_9790,N_9804);
nand U9899 (N_9899,N_9766,N_9811);
and U9900 (N_9900,N_9835,N_9861);
nor U9901 (N_9901,N_9840,N_9752);
xnor U9902 (N_9902,N_9765,N_9838);
nand U9903 (N_9903,N_9792,N_9757);
and U9904 (N_9904,N_9782,N_9756);
or U9905 (N_9905,N_9780,N_9855);
nor U9906 (N_9906,N_9859,N_9759);
xor U9907 (N_9907,N_9796,N_9822);
or U9908 (N_9908,N_9788,N_9754);
nor U9909 (N_9909,N_9848,N_9853);
nand U9910 (N_9910,N_9768,N_9842);
and U9911 (N_9911,N_9863,N_9865);
nand U9912 (N_9912,N_9755,N_9776);
and U9913 (N_9913,N_9806,N_9771);
xnor U9914 (N_9914,N_9773,N_9821);
nand U9915 (N_9915,N_9799,N_9871);
nand U9916 (N_9916,N_9869,N_9802);
nand U9917 (N_9917,N_9823,N_9797);
and U9918 (N_9918,N_9866,N_9854);
nand U9919 (N_9919,N_9763,N_9860);
or U9920 (N_9920,N_9849,N_9867);
nand U9921 (N_9921,N_9874,N_9775);
nand U9922 (N_9922,N_9825,N_9839);
nor U9923 (N_9923,N_9785,N_9787);
xnor U9924 (N_9924,N_9830,N_9817);
and U9925 (N_9925,N_9778,N_9852);
nor U9926 (N_9926,N_9813,N_9846);
nand U9927 (N_9927,N_9818,N_9872);
nand U9928 (N_9928,N_9762,N_9847);
nor U9929 (N_9929,N_9772,N_9794);
nand U9930 (N_9930,N_9819,N_9844);
or U9931 (N_9931,N_9751,N_9789);
nor U9932 (N_9932,N_9850,N_9845);
or U9933 (N_9933,N_9828,N_9831);
or U9934 (N_9934,N_9781,N_9832);
xnor U9935 (N_9935,N_9836,N_9795);
xnor U9936 (N_9936,N_9870,N_9816);
nand U9937 (N_9937,N_9767,N_9789);
nand U9938 (N_9938,N_9760,N_9811);
or U9939 (N_9939,N_9841,N_9834);
xnor U9940 (N_9940,N_9820,N_9813);
and U9941 (N_9941,N_9768,N_9828);
xor U9942 (N_9942,N_9810,N_9813);
or U9943 (N_9943,N_9753,N_9856);
or U9944 (N_9944,N_9823,N_9769);
xor U9945 (N_9945,N_9788,N_9853);
or U9946 (N_9946,N_9815,N_9785);
nor U9947 (N_9947,N_9825,N_9809);
nor U9948 (N_9948,N_9858,N_9786);
or U9949 (N_9949,N_9851,N_9762);
or U9950 (N_9950,N_9791,N_9808);
and U9951 (N_9951,N_9775,N_9809);
nor U9952 (N_9952,N_9770,N_9809);
xnor U9953 (N_9953,N_9754,N_9769);
nor U9954 (N_9954,N_9840,N_9825);
nor U9955 (N_9955,N_9768,N_9775);
nand U9956 (N_9956,N_9772,N_9796);
or U9957 (N_9957,N_9825,N_9790);
xnor U9958 (N_9958,N_9874,N_9789);
nor U9959 (N_9959,N_9813,N_9861);
and U9960 (N_9960,N_9819,N_9770);
xnor U9961 (N_9961,N_9758,N_9762);
or U9962 (N_9962,N_9836,N_9874);
nor U9963 (N_9963,N_9867,N_9859);
and U9964 (N_9964,N_9798,N_9834);
nor U9965 (N_9965,N_9800,N_9853);
or U9966 (N_9966,N_9841,N_9822);
or U9967 (N_9967,N_9874,N_9858);
nor U9968 (N_9968,N_9850,N_9828);
and U9969 (N_9969,N_9790,N_9843);
xnor U9970 (N_9970,N_9874,N_9871);
nand U9971 (N_9971,N_9847,N_9789);
or U9972 (N_9972,N_9760,N_9808);
xnor U9973 (N_9973,N_9770,N_9843);
xnor U9974 (N_9974,N_9763,N_9842);
or U9975 (N_9975,N_9829,N_9765);
nor U9976 (N_9976,N_9832,N_9864);
nor U9977 (N_9977,N_9793,N_9768);
nand U9978 (N_9978,N_9856,N_9784);
nand U9979 (N_9979,N_9817,N_9848);
nor U9980 (N_9980,N_9871,N_9770);
nand U9981 (N_9981,N_9772,N_9775);
nand U9982 (N_9982,N_9801,N_9787);
nor U9983 (N_9983,N_9864,N_9827);
or U9984 (N_9984,N_9781,N_9760);
and U9985 (N_9985,N_9784,N_9830);
or U9986 (N_9986,N_9798,N_9778);
and U9987 (N_9987,N_9853,N_9854);
and U9988 (N_9988,N_9783,N_9805);
and U9989 (N_9989,N_9751,N_9835);
and U9990 (N_9990,N_9798,N_9791);
xor U9991 (N_9991,N_9838,N_9806);
nand U9992 (N_9992,N_9816,N_9828);
xnor U9993 (N_9993,N_9787,N_9756);
or U9994 (N_9994,N_9830,N_9787);
nand U9995 (N_9995,N_9854,N_9757);
nor U9996 (N_9996,N_9860,N_9788);
xor U9997 (N_9997,N_9820,N_9860);
xnor U9998 (N_9998,N_9808,N_9829);
xnor U9999 (N_9999,N_9780,N_9785);
xor U10000 (N_10000,N_9976,N_9905);
and U10001 (N_10001,N_9883,N_9966);
nand U10002 (N_10002,N_9887,N_9971);
nand U10003 (N_10003,N_9948,N_9891);
and U10004 (N_10004,N_9918,N_9978);
and U10005 (N_10005,N_9890,N_9888);
and U10006 (N_10006,N_9906,N_9878);
nand U10007 (N_10007,N_9896,N_9907);
and U10008 (N_10008,N_9898,N_9877);
or U10009 (N_10009,N_9929,N_9988);
xor U10010 (N_10010,N_9920,N_9982);
and U10011 (N_10011,N_9919,N_9892);
nand U10012 (N_10012,N_9952,N_9980);
nor U10013 (N_10013,N_9926,N_9880);
or U10014 (N_10014,N_9881,N_9957);
xor U10015 (N_10015,N_9884,N_9947);
nand U10016 (N_10016,N_9902,N_9916);
nor U10017 (N_10017,N_9979,N_9917);
or U10018 (N_10018,N_9989,N_9944);
and U10019 (N_10019,N_9908,N_9893);
and U10020 (N_10020,N_9960,N_9993);
and U10021 (N_10021,N_9974,N_9885);
nor U10022 (N_10022,N_9981,N_9934);
nor U10023 (N_10023,N_9897,N_9939);
nor U10024 (N_10024,N_9899,N_9994);
nor U10025 (N_10025,N_9953,N_9889);
or U10026 (N_10026,N_9901,N_9962);
and U10027 (N_10027,N_9875,N_9932);
or U10028 (N_10028,N_9963,N_9911);
xnor U10029 (N_10029,N_9922,N_9910);
xnor U10030 (N_10030,N_9914,N_9925);
and U10031 (N_10031,N_9999,N_9965);
or U10032 (N_10032,N_9956,N_9923);
or U10033 (N_10033,N_9968,N_9894);
or U10034 (N_10034,N_9938,N_9970);
nor U10035 (N_10035,N_9969,N_9998);
or U10036 (N_10036,N_9972,N_9927);
nand U10037 (N_10037,N_9886,N_9983);
and U10038 (N_10038,N_9996,N_9943);
nor U10039 (N_10039,N_9900,N_9931);
nor U10040 (N_10040,N_9895,N_9903);
nor U10041 (N_10041,N_9990,N_9955);
nor U10042 (N_10042,N_9995,N_9967);
or U10043 (N_10043,N_9909,N_9959);
nor U10044 (N_10044,N_9958,N_9985);
xnor U10045 (N_10045,N_9946,N_9949);
xnor U10046 (N_10046,N_9986,N_9924);
nand U10047 (N_10047,N_9942,N_9987);
xnor U10048 (N_10048,N_9945,N_9997);
nor U10049 (N_10049,N_9950,N_9879);
and U10050 (N_10050,N_9915,N_9936);
or U10051 (N_10051,N_9975,N_9912);
nor U10052 (N_10052,N_9921,N_9991);
nor U10053 (N_10053,N_9882,N_9913);
nor U10054 (N_10054,N_9876,N_9954);
and U10055 (N_10055,N_9977,N_9984);
and U10056 (N_10056,N_9951,N_9904);
xnor U10057 (N_10057,N_9941,N_9940);
and U10058 (N_10058,N_9930,N_9937);
nand U10059 (N_10059,N_9935,N_9973);
or U10060 (N_10060,N_9928,N_9933);
xnor U10061 (N_10061,N_9992,N_9961);
and U10062 (N_10062,N_9964,N_9977);
or U10063 (N_10063,N_9944,N_9997);
or U10064 (N_10064,N_9912,N_9934);
or U10065 (N_10065,N_9950,N_9956);
and U10066 (N_10066,N_9964,N_9925);
xor U10067 (N_10067,N_9947,N_9961);
or U10068 (N_10068,N_9924,N_9889);
or U10069 (N_10069,N_9957,N_9943);
nor U10070 (N_10070,N_9963,N_9969);
and U10071 (N_10071,N_9937,N_9895);
nand U10072 (N_10072,N_9933,N_9908);
and U10073 (N_10073,N_9920,N_9990);
nand U10074 (N_10074,N_9897,N_9998);
nand U10075 (N_10075,N_9906,N_9876);
or U10076 (N_10076,N_9919,N_9912);
and U10077 (N_10077,N_9884,N_9894);
xnor U10078 (N_10078,N_9919,N_9968);
nand U10079 (N_10079,N_9884,N_9881);
or U10080 (N_10080,N_9912,N_9923);
nand U10081 (N_10081,N_9940,N_9875);
xor U10082 (N_10082,N_9967,N_9951);
xor U10083 (N_10083,N_9971,N_9942);
nand U10084 (N_10084,N_9950,N_9997);
and U10085 (N_10085,N_9979,N_9927);
nor U10086 (N_10086,N_9984,N_9976);
xnor U10087 (N_10087,N_9912,N_9946);
nor U10088 (N_10088,N_9978,N_9909);
nand U10089 (N_10089,N_9897,N_9997);
or U10090 (N_10090,N_9980,N_9909);
xnor U10091 (N_10091,N_9904,N_9990);
xor U10092 (N_10092,N_9972,N_9940);
and U10093 (N_10093,N_9890,N_9975);
nand U10094 (N_10094,N_9879,N_9981);
nand U10095 (N_10095,N_9997,N_9980);
and U10096 (N_10096,N_9985,N_9925);
nor U10097 (N_10097,N_9991,N_9990);
nor U10098 (N_10098,N_9947,N_9944);
and U10099 (N_10099,N_9945,N_9974);
or U10100 (N_10100,N_9955,N_9895);
xnor U10101 (N_10101,N_9981,N_9978);
xnor U10102 (N_10102,N_9902,N_9957);
nand U10103 (N_10103,N_9972,N_9974);
nand U10104 (N_10104,N_9907,N_9986);
nor U10105 (N_10105,N_9986,N_9899);
nor U10106 (N_10106,N_9947,N_9994);
or U10107 (N_10107,N_9888,N_9891);
nor U10108 (N_10108,N_9986,N_9977);
xor U10109 (N_10109,N_9916,N_9887);
nor U10110 (N_10110,N_9900,N_9976);
nor U10111 (N_10111,N_9978,N_9931);
and U10112 (N_10112,N_9940,N_9897);
xnor U10113 (N_10113,N_9995,N_9933);
nor U10114 (N_10114,N_9971,N_9950);
and U10115 (N_10115,N_9917,N_9997);
nand U10116 (N_10116,N_9909,N_9927);
nor U10117 (N_10117,N_9972,N_9914);
nor U10118 (N_10118,N_9887,N_9898);
and U10119 (N_10119,N_9935,N_9930);
nor U10120 (N_10120,N_9994,N_9886);
xor U10121 (N_10121,N_9964,N_9922);
or U10122 (N_10122,N_9896,N_9899);
nor U10123 (N_10123,N_9942,N_9973);
and U10124 (N_10124,N_9900,N_9892);
nand U10125 (N_10125,N_10011,N_10116);
xor U10126 (N_10126,N_10028,N_10103);
or U10127 (N_10127,N_10007,N_10000);
and U10128 (N_10128,N_10076,N_10115);
and U10129 (N_10129,N_10060,N_10001);
and U10130 (N_10130,N_10113,N_10021);
or U10131 (N_10131,N_10071,N_10012);
nand U10132 (N_10132,N_10009,N_10063);
xor U10133 (N_10133,N_10014,N_10057);
or U10134 (N_10134,N_10002,N_10122);
or U10135 (N_10135,N_10008,N_10020);
nand U10136 (N_10136,N_10083,N_10069);
nor U10137 (N_10137,N_10098,N_10029);
nor U10138 (N_10138,N_10036,N_10065);
or U10139 (N_10139,N_10033,N_10110);
xnor U10140 (N_10140,N_10015,N_10093);
or U10141 (N_10141,N_10042,N_10017);
nand U10142 (N_10142,N_10034,N_10104);
or U10143 (N_10143,N_10059,N_10114);
nand U10144 (N_10144,N_10091,N_10051);
nand U10145 (N_10145,N_10074,N_10038);
xnor U10146 (N_10146,N_10101,N_10022);
and U10147 (N_10147,N_10124,N_10062);
nand U10148 (N_10148,N_10018,N_10092);
nor U10149 (N_10149,N_10089,N_10067);
and U10150 (N_10150,N_10095,N_10005);
or U10151 (N_10151,N_10047,N_10117);
or U10152 (N_10152,N_10026,N_10121);
nand U10153 (N_10153,N_10044,N_10081);
nor U10154 (N_10154,N_10019,N_10032);
nand U10155 (N_10155,N_10072,N_10077);
or U10156 (N_10156,N_10107,N_10056);
nor U10157 (N_10157,N_10037,N_10054);
xor U10158 (N_10158,N_10004,N_10090);
or U10159 (N_10159,N_10084,N_10087);
nor U10160 (N_10160,N_10013,N_10119);
and U10161 (N_10161,N_10064,N_10023);
nor U10162 (N_10162,N_10118,N_10043);
nand U10163 (N_10163,N_10053,N_10111);
and U10164 (N_10164,N_10061,N_10070);
xor U10165 (N_10165,N_10045,N_10106);
and U10166 (N_10166,N_10082,N_10025);
nor U10167 (N_10167,N_10108,N_10010);
and U10168 (N_10168,N_10040,N_10055);
and U10169 (N_10169,N_10003,N_10024);
or U10170 (N_10170,N_10112,N_10046);
nor U10171 (N_10171,N_10123,N_10120);
nand U10172 (N_10172,N_10039,N_10050);
nor U10173 (N_10173,N_10105,N_10048);
or U10174 (N_10174,N_10030,N_10049);
and U10175 (N_10175,N_10006,N_10096);
and U10176 (N_10176,N_10079,N_10080);
or U10177 (N_10177,N_10085,N_10088);
nor U10178 (N_10178,N_10052,N_10097);
nand U10179 (N_10179,N_10075,N_10102);
xor U10180 (N_10180,N_10086,N_10078);
or U10181 (N_10181,N_10041,N_10094);
and U10182 (N_10182,N_10109,N_10058);
nand U10183 (N_10183,N_10068,N_10027);
xor U10184 (N_10184,N_10066,N_10031);
nor U10185 (N_10185,N_10016,N_10099);
nand U10186 (N_10186,N_10073,N_10035);
and U10187 (N_10187,N_10100,N_10062);
and U10188 (N_10188,N_10120,N_10114);
xor U10189 (N_10189,N_10122,N_10063);
xnor U10190 (N_10190,N_10106,N_10061);
or U10191 (N_10191,N_10078,N_10051);
or U10192 (N_10192,N_10046,N_10017);
nor U10193 (N_10193,N_10123,N_10048);
or U10194 (N_10194,N_10047,N_10017);
nor U10195 (N_10195,N_10025,N_10064);
nor U10196 (N_10196,N_10007,N_10062);
or U10197 (N_10197,N_10031,N_10052);
xnor U10198 (N_10198,N_10079,N_10090);
and U10199 (N_10199,N_10066,N_10045);
nand U10200 (N_10200,N_10082,N_10065);
nand U10201 (N_10201,N_10101,N_10077);
nand U10202 (N_10202,N_10066,N_10103);
nand U10203 (N_10203,N_10006,N_10022);
or U10204 (N_10204,N_10032,N_10033);
xor U10205 (N_10205,N_10043,N_10040);
xnor U10206 (N_10206,N_10114,N_10049);
and U10207 (N_10207,N_10011,N_10096);
nand U10208 (N_10208,N_10069,N_10036);
nor U10209 (N_10209,N_10053,N_10056);
and U10210 (N_10210,N_10060,N_10098);
and U10211 (N_10211,N_10046,N_10035);
and U10212 (N_10212,N_10061,N_10105);
nand U10213 (N_10213,N_10059,N_10089);
or U10214 (N_10214,N_10027,N_10066);
xnor U10215 (N_10215,N_10109,N_10004);
nor U10216 (N_10216,N_10090,N_10022);
nor U10217 (N_10217,N_10078,N_10012);
or U10218 (N_10218,N_10058,N_10114);
nor U10219 (N_10219,N_10072,N_10085);
nor U10220 (N_10220,N_10010,N_10088);
or U10221 (N_10221,N_10078,N_10041);
nor U10222 (N_10222,N_10053,N_10027);
nand U10223 (N_10223,N_10003,N_10118);
xnor U10224 (N_10224,N_10068,N_10093);
or U10225 (N_10225,N_10055,N_10019);
and U10226 (N_10226,N_10095,N_10027);
or U10227 (N_10227,N_10025,N_10030);
nand U10228 (N_10228,N_10114,N_10068);
xnor U10229 (N_10229,N_10078,N_10117);
nor U10230 (N_10230,N_10068,N_10119);
and U10231 (N_10231,N_10002,N_10110);
nand U10232 (N_10232,N_10121,N_10069);
nor U10233 (N_10233,N_10009,N_10113);
xnor U10234 (N_10234,N_10022,N_10076);
nand U10235 (N_10235,N_10089,N_10086);
or U10236 (N_10236,N_10085,N_10053);
and U10237 (N_10237,N_10113,N_10078);
xor U10238 (N_10238,N_10051,N_10033);
or U10239 (N_10239,N_10014,N_10041);
nor U10240 (N_10240,N_10066,N_10096);
nand U10241 (N_10241,N_10066,N_10036);
xor U10242 (N_10242,N_10037,N_10007);
xnor U10243 (N_10243,N_10083,N_10116);
nor U10244 (N_10244,N_10065,N_10109);
or U10245 (N_10245,N_10009,N_10029);
nor U10246 (N_10246,N_10118,N_10081);
and U10247 (N_10247,N_10073,N_10009);
xor U10248 (N_10248,N_10047,N_10058);
xor U10249 (N_10249,N_10019,N_10028);
nor U10250 (N_10250,N_10211,N_10162);
or U10251 (N_10251,N_10227,N_10130);
nand U10252 (N_10252,N_10248,N_10163);
nand U10253 (N_10253,N_10128,N_10176);
xor U10254 (N_10254,N_10177,N_10238);
xor U10255 (N_10255,N_10125,N_10155);
and U10256 (N_10256,N_10213,N_10190);
and U10257 (N_10257,N_10224,N_10178);
nor U10258 (N_10258,N_10133,N_10167);
and U10259 (N_10259,N_10191,N_10172);
nor U10260 (N_10260,N_10135,N_10146);
xor U10261 (N_10261,N_10221,N_10240);
nand U10262 (N_10262,N_10182,N_10225);
and U10263 (N_10263,N_10171,N_10193);
or U10264 (N_10264,N_10205,N_10144);
nand U10265 (N_10265,N_10247,N_10242);
nand U10266 (N_10266,N_10218,N_10134);
and U10267 (N_10267,N_10245,N_10129);
xor U10268 (N_10268,N_10132,N_10142);
or U10269 (N_10269,N_10180,N_10157);
nand U10270 (N_10270,N_10217,N_10241);
xnor U10271 (N_10271,N_10209,N_10152);
nand U10272 (N_10272,N_10232,N_10199);
nor U10273 (N_10273,N_10215,N_10138);
or U10274 (N_10274,N_10197,N_10235);
xor U10275 (N_10275,N_10194,N_10181);
nor U10276 (N_10276,N_10228,N_10233);
xor U10277 (N_10277,N_10184,N_10196);
nor U10278 (N_10278,N_10139,N_10203);
xnor U10279 (N_10279,N_10222,N_10143);
and U10280 (N_10280,N_10174,N_10186);
nor U10281 (N_10281,N_10187,N_10185);
xnor U10282 (N_10282,N_10136,N_10151);
nand U10283 (N_10283,N_10214,N_10137);
xor U10284 (N_10284,N_10179,N_10150);
xnor U10285 (N_10285,N_10223,N_10127);
or U10286 (N_10286,N_10244,N_10208);
nor U10287 (N_10287,N_10220,N_10234);
nor U10288 (N_10288,N_10212,N_10154);
or U10289 (N_10289,N_10148,N_10149);
nand U10290 (N_10290,N_10145,N_10192);
and U10291 (N_10291,N_10141,N_10165);
nor U10292 (N_10292,N_10207,N_10158);
nor U10293 (N_10293,N_10219,N_10126);
xnor U10294 (N_10294,N_10166,N_10147);
or U10295 (N_10295,N_10206,N_10140);
or U10296 (N_10296,N_10153,N_10243);
nor U10297 (N_10297,N_10216,N_10188);
nor U10298 (N_10298,N_10237,N_10168);
or U10299 (N_10299,N_10156,N_10204);
nand U10300 (N_10300,N_10231,N_10229);
xnor U10301 (N_10301,N_10160,N_10198);
or U10302 (N_10302,N_10170,N_10249);
nor U10303 (N_10303,N_10195,N_10210);
nor U10304 (N_10304,N_10189,N_10131);
xnor U10305 (N_10305,N_10202,N_10183);
nand U10306 (N_10306,N_10230,N_10246);
xor U10307 (N_10307,N_10239,N_10159);
or U10308 (N_10308,N_10226,N_10175);
and U10309 (N_10309,N_10164,N_10236);
nand U10310 (N_10310,N_10169,N_10201);
or U10311 (N_10311,N_10161,N_10200);
xnor U10312 (N_10312,N_10173,N_10183);
xnor U10313 (N_10313,N_10140,N_10147);
nand U10314 (N_10314,N_10235,N_10134);
or U10315 (N_10315,N_10214,N_10220);
nand U10316 (N_10316,N_10134,N_10175);
nor U10317 (N_10317,N_10143,N_10188);
nor U10318 (N_10318,N_10133,N_10175);
xnor U10319 (N_10319,N_10179,N_10211);
nand U10320 (N_10320,N_10143,N_10200);
nor U10321 (N_10321,N_10223,N_10239);
and U10322 (N_10322,N_10167,N_10185);
xnor U10323 (N_10323,N_10147,N_10180);
nor U10324 (N_10324,N_10175,N_10244);
and U10325 (N_10325,N_10211,N_10130);
nand U10326 (N_10326,N_10202,N_10205);
nor U10327 (N_10327,N_10236,N_10166);
and U10328 (N_10328,N_10183,N_10140);
or U10329 (N_10329,N_10218,N_10188);
or U10330 (N_10330,N_10219,N_10217);
or U10331 (N_10331,N_10239,N_10181);
nand U10332 (N_10332,N_10189,N_10201);
nor U10333 (N_10333,N_10242,N_10166);
xnor U10334 (N_10334,N_10198,N_10241);
xnor U10335 (N_10335,N_10137,N_10219);
or U10336 (N_10336,N_10218,N_10235);
or U10337 (N_10337,N_10240,N_10158);
and U10338 (N_10338,N_10143,N_10211);
or U10339 (N_10339,N_10133,N_10173);
nand U10340 (N_10340,N_10152,N_10190);
and U10341 (N_10341,N_10134,N_10167);
nand U10342 (N_10342,N_10175,N_10222);
or U10343 (N_10343,N_10158,N_10236);
nand U10344 (N_10344,N_10169,N_10133);
and U10345 (N_10345,N_10173,N_10135);
nand U10346 (N_10346,N_10225,N_10235);
nand U10347 (N_10347,N_10211,N_10227);
xnor U10348 (N_10348,N_10170,N_10165);
nor U10349 (N_10349,N_10207,N_10155);
or U10350 (N_10350,N_10175,N_10146);
nand U10351 (N_10351,N_10195,N_10242);
nor U10352 (N_10352,N_10177,N_10141);
or U10353 (N_10353,N_10181,N_10161);
xor U10354 (N_10354,N_10144,N_10147);
nand U10355 (N_10355,N_10173,N_10126);
nand U10356 (N_10356,N_10201,N_10249);
xor U10357 (N_10357,N_10239,N_10161);
nand U10358 (N_10358,N_10178,N_10127);
and U10359 (N_10359,N_10244,N_10220);
and U10360 (N_10360,N_10192,N_10218);
nor U10361 (N_10361,N_10149,N_10152);
nor U10362 (N_10362,N_10192,N_10211);
or U10363 (N_10363,N_10146,N_10196);
nor U10364 (N_10364,N_10213,N_10206);
nor U10365 (N_10365,N_10248,N_10214);
nor U10366 (N_10366,N_10240,N_10175);
and U10367 (N_10367,N_10146,N_10160);
xor U10368 (N_10368,N_10185,N_10142);
nor U10369 (N_10369,N_10143,N_10227);
nor U10370 (N_10370,N_10210,N_10138);
nand U10371 (N_10371,N_10175,N_10161);
xnor U10372 (N_10372,N_10244,N_10127);
nor U10373 (N_10373,N_10211,N_10166);
nand U10374 (N_10374,N_10193,N_10204);
nor U10375 (N_10375,N_10302,N_10343);
xor U10376 (N_10376,N_10318,N_10373);
nor U10377 (N_10377,N_10297,N_10308);
nor U10378 (N_10378,N_10340,N_10354);
xnor U10379 (N_10379,N_10298,N_10251);
and U10380 (N_10380,N_10273,N_10327);
nor U10381 (N_10381,N_10293,N_10339);
xnor U10382 (N_10382,N_10270,N_10271);
or U10383 (N_10383,N_10320,N_10277);
nor U10384 (N_10384,N_10304,N_10371);
xnor U10385 (N_10385,N_10261,N_10284);
or U10386 (N_10386,N_10265,N_10316);
nand U10387 (N_10387,N_10328,N_10250);
and U10388 (N_10388,N_10263,N_10370);
nor U10389 (N_10389,N_10367,N_10355);
xor U10390 (N_10390,N_10357,N_10366);
or U10391 (N_10391,N_10260,N_10358);
or U10392 (N_10392,N_10344,N_10295);
xnor U10393 (N_10393,N_10359,N_10317);
nor U10394 (N_10394,N_10319,N_10351);
nor U10395 (N_10395,N_10296,N_10347);
nor U10396 (N_10396,N_10360,N_10356);
or U10397 (N_10397,N_10274,N_10300);
xor U10398 (N_10398,N_10303,N_10278);
nor U10399 (N_10399,N_10348,N_10337);
xor U10400 (N_10400,N_10290,N_10372);
or U10401 (N_10401,N_10330,N_10353);
nand U10402 (N_10402,N_10311,N_10306);
and U10403 (N_10403,N_10291,N_10324);
or U10404 (N_10404,N_10350,N_10364);
xnor U10405 (N_10405,N_10352,N_10333);
or U10406 (N_10406,N_10282,N_10331);
nand U10407 (N_10407,N_10279,N_10338);
nor U10408 (N_10408,N_10254,N_10287);
xnor U10409 (N_10409,N_10259,N_10256);
and U10410 (N_10410,N_10289,N_10361);
xnor U10411 (N_10411,N_10341,N_10365);
nand U10412 (N_10412,N_10255,N_10286);
nor U10413 (N_10413,N_10362,N_10309);
or U10414 (N_10414,N_10285,N_10281);
or U10415 (N_10415,N_10258,N_10283);
nand U10416 (N_10416,N_10257,N_10276);
xnor U10417 (N_10417,N_10335,N_10321);
nand U10418 (N_10418,N_10305,N_10368);
xnor U10419 (N_10419,N_10369,N_10329);
and U10420 (N_10420,N_10294,N_10374);
nor U10421 (N_10421,N_10272,N_10292);
or U10422 (N_10422,N_10301,N_10252);
xnor U10423 (N_10423,N_10332,N_10345);
nand U10424 (N_10424,N_10314,N_10322);
xor U10425 (N_10425,N_10312,N_10275);
nand U10426 (N_10426,N_10307,N_10349);
nand U10427 (N_10427,N_10310,N_10299);
and U10428 (N_10428,N_10269,N_10253);
or U10429 (N_10429,N_10326,N_10323);
nand U10430 (N_10430,N_10264,N_10288);
xnor U10431 (N_10431,N_10346,N_10268);
xnor U10432 (N_10432,N_10315,N_10280);
nand U10433 (N_10433,N_10363,N_10262);
nand U10434 (N_10434,N_10325,N_10334);
xnor U10435 (N_10435,N_10267,N_10342);
nand U10436 (N_10436,N_10313,N_10336);
and U10437 (N_10437,N_10266,N_10253);
nand U10438 (N_10438,N_10251,N_10297);
nand U10439 (N_10439,N_10330,N_10268);
nor U10440 (N_10440,N_10343,N_10278);
or U10441 (N_10441,N_10302,N_10358);
or U10442 (N_10442,N_10308,N_10268);
and U10443 (N_10443,N_10360,N_10364);
xnor U10444 (N_10444,N_10261,N_10298);
nor U10445 (N_10445,N_10351,N_10283);
xnor U10446 (N_10446,N_10286,N_10302);
nand U10447 (N_10447,N_10277,N_10275);
xor U10448 (N_10448,N_10281,N_10274);
and U10449 (N_10449,N_10320,N_10307);
and U10450 (N_10450,N_10274,N_10343);
xor U10451 (N_10451,N_10347,N_10277);
nor U10452 (N_10452,N_10321,N_10342);
or U10453 (N_10453,N_10311,N_10281);
and U10454 (N_10454,N_10337,N_10340);
nor U10455 (N_10455,N_10338,N_10355);
or U10456 (N_10456,N_10370,N_10347);
xor U10457 (N_10457,N_10344,N_10302);
or U10458 (N_10458,N_10268,N_10252);
xnor U10459 (N_10459,N_10250,N_10314);
xnor U10460 (N_10460,N_10345,N_10338);
and U10461 (N_10461,N_10275,N_10287);
and U10462 (N_10462,N_10325,N_10268);
xnor U10463 (N_10463,N_10293,N_10370);
nor U10464 (N_10464,N_10268,N_10363);
or U10465 (N_10465,N_10287,N_10284);
xnor U10466 (N_10466,N_10295,N_10339);
nor U10467 (N_10467,N_10331,N_10344);
nor U10468 (N_10468,N_10279,N_10250);
or U10469 (N_10469,N_10362,N_10301);
xnor U10470 (N_10470,N_10358,N_10322);
and U10471 (N_10471,N_10327,N_10348);
or U10472 (N_10472,N_10320,N_10286);
or U10473 (N_10473,N_10370,N_10334);
and U10474 (N_10474,N_10363,N_10336);
or U10475 (N_10475,N_10306,N_10360);
or U10476 (N_10476,N_10360,N_10265);
nor U10477 (N_10477,N_10370,N_10373);
and U10478 (N_10478,N_10368,N_10311);
nor U10479 (N_10479,N_10313,N_10367);
and U10480 (N_10480,N_10289,N_10252);
and U10481 (N_10481,N_10280,N_10347);
nor U10482 (N_10482,N_10311,N_10344);
xnor U10483 (N_10483,N_10322,N_10266);
and U10484 (N_10484,N_10272,N_10301);
nor U10485 (N_10485,N_10275,N_10363);
xnor U10486 (N_10486,N_10357,N_10362);
or U10487 (N_10487,N_10347,N_10353);
nor U10488 (N_10488,N_10267,N_10270);
xnor U10489 (N_10489,N_10278,N_10356);
nand U10490 (N_10490,N_10332,N_10258);
nor U10491 (N_10491,N_10293,N_10305);
or U10492 (N_10492,N_10258,N_10367);
xor U10493 (N_10493,N_10279,N_10285);
nand U10494 (N_10494,N_10370,N_10274);
nor U10495 (N_10495,N_10268,N_10263);
xnor U10496 (N_10496,N_10277,N_10374);
and U10497 (N_10497,N_10283,N_10255);
xor U10498 (N_10498,N_10296,N_10278);
or U10499 (N_10499,N_10363,N_10255);
nor U10500 (N_10500,N_10450,N_10425);
nand U10501 (N_10501,N_10397,N_10404);
nor U10502 (N_10502,N_10491,N_10439);
xor U10503 (N_10503,N_10451,N_10376);
or U10504 (N_10504,N_10430,N_10488);
xnor U10505 (N_10505,N_10419,N_10498);
nor U10506 (N_10506,N_10481,N_10384);
nor U10507 (N_10507,N_10445,N_10442);
or U10508 (N_10508,N_10471,N_10473);
xnor U10509 (N_10509,N_10475,N_10433);
nor U10510 (N_10510,N_10455,N_10416);
nor U10511 (N_10511,N_10423,N_10453);
and U10512 (N_10512,N_10493,N_10467);
or U10513 (N_10513,N_10414,N_10420);
or U10514 (N_10514,N_10474,N_10496);
or U10515 (N_10515,N_10378,N_10470);
xor U10516 (N_10516,N_10459,N_10438);
and U10517 (N_10517,N_10380,N_10476);
nand U10518 (N_10518,N_10457,N_10490);
or U10519 (N_10519,N_10417,N_10452);
xnor U10520 (N_10520,N_10408,N_10413);
xnor U10521 (N_10521,N_10392,N_10401);
nor U10522 (N_10522,N_10407,N_10432);
and U10523 (N_10523,N_10441,N_10446);
xor U10524 (N_10524,N_10447,N_10434);
nand U10525 (N_10525,N_10383,N_10497);
nor U10526 (N_10526,N_10465,N_10431);
nor U10527 (N_10527,N_10482,N_10400);
xnor U10528 (N_10528,N_10387,N_10484);
and U10529 (N_10529,N_10485,N_10435);
nand U10530 (N_10530,N_10396,N_10479);
or U10531 (N_10531,N_10478,N_10440);
nor U10532 (N_10532,N_10437,N_10444);
nor U10533 (N_10533,N_10461,N_10487);
xor U10534 (N_10534,N_10426,N_10464);
xor U10535 (N_10535,N_10499,N_10456);
xnor U10536 (N_10536,N_10421,N_10489);
xnor U10537 (N_10537,N_10466,N_10428);
or U10538 (N_10538,N_10449,N_10395);
or U10539 (N_10539,N_10443,N_10427);
nand U10540 (N_10540,N_10480,N_10405);
or U10541 (N_10541,N_10469,N_10393);
and U10542 (N_10542,N_10429,N_10409);
xnor U10543 (N_10543,N_10381,N_10410);
nand U10544 (N_10544,N_10377,N_10412);
nand U10545 (N_10545,N_10388,N_10495);
nor U10546 (N_10546,N_10458,N_10382);
and U10547 (N_10547,N_10389,N_10398);
xor U10548 (N_10548,N_10486,N_10379);
and U10549 (N_10549,N_10477,N_10386);
and U10550 (N_10550,N_10424,N_10418);
nand U10551 (N_10551,N_10436,N_10406);
or U10552 (N_10552,N_10448,N_10399);
nor U10553 (N_10553,N_10462,N_10391);
nand U10554 (N_10554,N_10403,N_10415);
nor U10555 (N_10555,N_10385,N_10483);
xnor U10556 (N_10556,N_10390,N_10472);
nor U10557 (N_10557,N_10402,N_10375);
or U10558 (N_10558,N_10492,N_10460);
and U10559 (N_10559,N_10468,N_10494);
nor U10560 (N_10560,N_10394,N_10454);
xnor U10561 (N_10561,N_10422,N_10411);
xnor U10562 (N_10562,N_10463,N_10378);
or U10563 (N_10563,N_10383,N_10387);
xor U10564 (N_10564,N_10380,N_10399);
nor U10565 (N_10565,N_10375,N_10422);
xor U10566 (N_10566,N_10384,N_10467);
and U10567 (N_10567,N_10457,N_10447);
nor U10568 (N_10568,N_10435,N_10471);
nand U10569 (N_10569,N_10498,N_10450);
xor U10570 (N_10570,N_10390,N_10379);
and U10571 (N_10571,N_10498,N_10476);
and U10572 (N_10572,N_10381,N_10412);
or U10573 (N_10573,N_10412,N_10407);
or U10574 (N_10574,N_10393,N_10457);
and U10575 (N_10575,N_10456,N_10395);
and U10576 (N_10576,N_10420,N_10450);
nor U10577 (N_10577,N_10378,N_10441);
and U10578 (N_10578,N_10492,N_10431);
nor U10579 (N_10579,N_10465,N_10481);
or U10580 (N_10580,N_10475,N_10409);
xnor U10581 (N_10581,N_10425,N_10385);
and U10582 (N_10582,N_10423,N_10392);
nor U10583 (N_10583,N_10412,N_10473);
or U10584 (N_10584,N_10387,N_10399);
xor U10585 (N_10585,N_10403,N_10399);
and U10586 (N_10586,N_10488,N_10409);
and U10587 (N_10587,N_10432,N_10461);
or U10588 (N_10588,N_10407,N_10395);
and U10589 (N_10589,N_10498,N_10377);
or U10590 (N_10590,N_10475,N_10458);
xnor U10591 (N_10591,N_10463,N_10454);
nor U10592 (N_10592,N_10416,N_10423);
or U10593 (N_10593,N_10382,N_10426);
or U10594 (N_10594,N_10432,N_10448);
or U10595 (N_10595,N_10453,N_10471);
and U10596 (N_10596,N_10471,N_10464);
nor U10597 (N_10597,N_10385,N_10451);
and U10598 (N_10598,N_10409,N_10454);
or U10599 (N_10599,N_10404,N_10476);
nand U10600 (N_10600,N_10445,N_10433);
nand U10601 (N_10601,N_10474,N_10424);
or U10602 (N_10602,N_10456,N_10444);
xnor U10603 (N_10603,N_10395,N_10402);
xor U10604 (N_10604,N_10393,N_10422);
xor U10605 (N_10605,N_10496,N_10407);
nor U10606 (N_10606,N_10428,N_10495);
nand U10607 (N_10607,N_10460,N_10443);
or U10608 (N_10608,N_10405,N_10454);
nor U10609 (N_10609,N_10483,N_10388);
or U10610 (N_10610,N_10463,N_10496);
or U10611 (N_10611,N_10496,N_10395);
xor U10612 (N_10612,N_10423,N_10406);
nand U10613 (N_10613,N_10468,N_10382);
xnor U10614 (N_10614,N_10462,N_10439);
nand U10615 (N_10615,N_10408,N_10457);
xor U10616 (N_10616,N_10484,N_10464);
or U10617 (N_10617,N_10405,N_10461);
or U10618 (N_10618,N_10429,N_10474);
xnor U10619 (N_10619,N_10493,N_10425);
xor U10620 (N_10620,N_10454,N_10395);
and U10621 (N_10621,N_10392,N_10408);
nand U10622 (N_10622,N_10440,N_10382);
xor U10623 (N_10623,N_10470,N_10495);
and U10624 (N_10624,N_10456,N_10440);
nor U10625 (N_10625,N_10505,N_10533);
or U10626 (N_10626,N_10508,N_10510);
and U10627 (N_10627,N_10569,N_10580);
nor U10628 (N_10628,N_10567,N_10516);
and U10629 (N_10629,N_10554,N_10602);
nor U10630 (N_10630,N_10520,N_10603);
or U10631 (N_10631,N_10503,N_10566);
nor U10632 (N_10632,N_10541,N_10622);
or U10633 (N_10633,N_10517,N_10585);
nand U10634 (N_10634,N_10624,N_10500);
nor U10635 (N_10635,N_10548,N_10591);
xor U10636 (N_10636,N_10515,N_10575);
nand U10637 (N_10637,N_10506,N_10538);
nor U10638 (N_10638,N_10527,N_10536);
xor U10639 (N_10639,N_10576,N_10599);
and U10640 (N_10640,N_10558,N_10590);
xnor U10641 (N_10641,N_10513,N_10557);
or U10642 (N_10642,N_10561,N_10525);
or U10643 (N_10643,N_10615,N_10560);
or U10644 (N_10644,N_10540,N_10523);
or U10645 (N_10645,N_10552,N_10612);
nand U10646 (N_10646,N_10530,N_10543);
nand U10647 (N_10647,N_10584,N_10619);
xnor U10648 (N_10648,N_10596,N_10617);
or U10649 (N_10649,N_10563,N_10572);
nand U10650 (N_10650,N_10532,N_10609);
or U10651 (N_10651,N_10608,N_10511);
nand U10652 (N_10652,N_10549,N_10597);
nand U10653 (N_10653,N_10577,N_10581);
or U10654 (N_10654,N_10507,N_10586);
xor U10655 (N_10655,N_10553,N_10588);
and U10656 (N_10656,N_10504,N_10528);
or U10657 (N_10657,N_10551,N_10601);
or U10658 (N_10658,N_10582,N_10565);
or U10659 (N_10659,N_10531,N_10521);
nand U10660 (N_10660,N_10562,N_10544);
xnor U10661 (N_10661,N_10539,N_10547);
nor U10662 (N_10662,N_10589,N_10579);
xor U10663 (N_10663,N_10550,N_10600);
nand U10664 (N_10664,N_10570,N_10556);
nor U10665 (N_10665,N_10545,N_10514);
and U10666 (N_10666,N_10592,N_10518);
and U10667 (N_10667,N_10509,N_10604);
and U10668 (N_10668,N_10611,N_10546);
nand U10669 (N_10669,N_10623,N_10542);
xnor U10670 (N_10670,N_10573,N_10512);
and U10671 (N_10671,N_10610,N_10613);
nor U10672 (N_10672,N_10559,N_10519);
xnor U10673 (N_10673,N_10595,N_10524);
nor U10674 (N_10674,N_10555,N_10574);
nand U10675 (N_10675,N_10534,N_10526);
and U10676 (N_10676,N_10620,N_10501);
nor U10677 (N_10677,N_10607,N_10621);
nand U10678 (N_10678,N_10571,N_10583);
nor U10679 (N_10679,N_10614,N_10568);
or U10680 (N_10680,N_10616,N_10593);
and U10681 (N_10681,N_10522,N_10537);
nand U10682 (N_10682,N_10598,N_10587);
nor U10683 (N_10683,N_10578,N_10605);
nand U10684 (N_10684,N_10502,N_10535);
xor U10685 (N_10685,N_10564,N_10606);
nand U10686 (N_10686,N_10529,N_10594);
nor U10687 (N_10687,N_10618,N_10551);
nor U10688 (N_10688,N_10593,N_10557);
and U10689 (N_10689,N_10610,N_10505);
nor U10690 (N_10690,N_10521,N_10504);
nor U10691 (N_10691,N_10607,N_10560);
nand U10692 (N_10692,N_10586,N_10582);
nor U10693 (N_10693,N_10602,N_10614);
and U10694 (N_10694,N_10555,N_10603);
and U10695 (N_10695,N_10504,N_10505);
or U10696 (N_10696,N_10589,N_10522);
nor U10697 (N_10697,N_10562,N_10610);
nor U10698 (N_10698,N_10614,N_10557);
xnor U10699 (N_10699,N_10593,N_10552);
or U10700 (N_10700,N_10580,N_10558);
nor U10701 (N_10701,N_10619,N_10507);
or U10702 (N_10702,N_10602,N_10561);
xnor U10703 (N_10703,N_10612,N_10618);
or U10704 (N_10704,N_10589,N_10595);
nand U10705 (N_10705,N_10513,N_10516);
xor U10706 (N_10706,N_10589,N_10610);
xor U10707 (N_10707,N_10554,N_10534);
xnor U10708 (N_10708,N_10572,N_10524);
nor U10709 (N_10709,N_10592,N_10575);
or U10710 (N_10710,N_10621,N_10585);
nor U10711 (N_10711,N_10609,N_10533);
nor U10712 (N_10712,N_10622,N_10505);
and U10713 (N_10713,N_10504,N_10611);
and U10714 (N_10714,N_10543,N_10605);
nand U10715 (N_10715,N_10556,N_10541);
and U10716 (N_10716,N_10502,N_10612);
and U10717 (N_10717,N_10619,N_10591);
xnor U10718 (N_10718,N_10519,N_10580);
xnor U10719 (N_10719,N_10589,N_10545);
nor U10720 (N_10720,N_10549,N_10569);
nor U10721 (N_10721,N_10528,N_10616);
or U10722 (N_10722,N_10582,N_10510);
nor U10723 (N_10723,N_10614,N_10539);
nor U10724 (N_10724,N_10603,N_10610);
and U10725 (N_10725,N_10618,N_10527);
nand U10726 (N_10726,N_10531,N_10500);
and U10727 (N_10727,N_10615,N_10570);
or U10728 (N_10728,N_10619,N_10508);
or U10729 (N_10729,N_10605,N_10604);
or U10730 (N_10730,N_10534,N_10577);
nand U10731 (N_10731,N_10582,N_10596);
or U10732 (N_10732,N_10514,N_10585);
nor U10733 (N_10733,N_10540,N_10545);
and U10734 (N_10734,N_10525,N_10543);
nand U10735 (N_10735,N_10598,N_10612);
xor U10736 (N_10736,N_10544,N_10598);
nor U10737 (N_10737,N_10536,N_10555);
nor U10738 (N_10738,N_10513,N_10533);
or U10739 (N_10739,N_10540,N_10574);
or U10740 (N_10740,N_10567,N_10598);
nor U10741 (N_10741,N_10506,N_10520);
nand U10742 (N_10742,N_10539,N_10561);
and U10743 (N_10743,N_10624,N_10591);
xnor U10744 (N_10744,N_10624,N_10613);
nor U10745 (N_10745,N_10544,N_10535);
and U10746 (N_10746,N_10547,N_10585);
or U10747 (N_10747,N_10521,N_10617);
nand U10748 (N_10748,N_10609,N_10585);
or U10749 (N_10749,N_10515,N_10546);
nor U10750 (N_10750,N_10631,N_10694);
and U10751 (N_10751,N_10630,N_10691);
xnor U10752 (N_10752,N_10693,N_10746);
xor U10753 (N_10753,N_10706,N_10696);
xnor U10754 (N_10754,N_10689,N_10731);
or U10755 (N_10755,N_10718,N_10687);
or U10756 (N_10756,N_10659,N_10692);
nor U10757 (N_10757,N_10721,N_10724);
nand U10758 (N_10758,N_10677,N_10716);
xor U10759 (N_10759,N_10629,N_10652);
nand U10760 (N_10760,N_10744,N_10699);
or U10761 (N_10761,N_10661,N_10668);
and U10762 (N_10762,N_10664,N_10737);
or U10763 (N_10763,N_10723,N_10714);
or U10764 (N_10764,N_10732,N_10636);
xnor U10765 (N_10765,N_10719,N_10634);
nand U10766 (N_10766,N_10669,N_10642);
and U10767 (N_10767,N_10701,N_10640);
or U10768 (N_10768,N_10660,N_10740);
and U10769 (N_10769,N_10729,N_10678);
nand U10770 (N_10770,N_10626,N_10681);
nor U10771 (N_10771,N_10698,N_10707);
or U10772 (N_10772,N_10730,N_10666);
or U10773 (N_10773,N_10748,N_10702);
xor U10774 (N_10774,N_10734,N_10651);
and U10775 (N_10775,N_10641,N_10720);
xnor U10776 (N_10776,N_10713,N_10646);
nor U10777 (N_10777,N_10662,N_10654);
nor U10778 (N_10778,N_10682,N_10717);
nor U10779 (N_10779,N_10627,N_10728);
nor U10780 (N_10780,N_10658,N_10633);
nand U10781 (N_10781,N_10738,N_10733);
or U10782 (N_10782,N_10684,N_10710);
xor U10783 (N_10783,N_10670,N_10690);
nand U10784 (N_10784,N_10650,N_10709);
or U10785 (N_10785,N_10643,N_10686);
nor U10786 (N_10786,N_10703,N_10679);
nor U10787 (N_10787,N_10739,N_10632);
xnor U10788 (N_10788,N_10674,N_10647);
nor U10789 (N_10789,N_10625,N_10656);
nor U10790 (N_10790,N_10742,N_10671);
nand U10791 (N_10791,N_10683,N_10675);
or U10792 (N_10792,N_10715,N_10708);
nor U10793 (N_10793,N_10705,N_10657);
nor U10794 (N_10794,N_10644,N_10704);
or U10795 (N_10795,N_10743,N_10722);
xor U10796 (N_10796,N_10712,N_10711);
nand U10797 (N_10797,N_10700,N_10672);
or U10798 (N_10798,N_10653,N_10726);
or U10799 (N_10799,N_10725,N_10735);
nand U10800 (N_10800,N_10685,N_10741);
or U10801 (N_10801,N_10663,N_10676);
nand U10802 (N_10802,N_10655,N_10649);
nor U10803 (N_10803,N_10680,N_10745);
xor U10804 (N_10804,N_10628,N_10688);
nor U10805 (N_10805,N_10747,N_10637);
or U10806 (N_10806,N_10638,N_10697);
and U10807 (N_10807,N_10645,N_10695);
xnor U10808 (N_10808,N_10639,N_10736);
nor U10809 (N_10809,N_10727,N_10665);
or U10810 (N_10810,N_10673,N_10667);
xnor U10811 (N_10811,N_10749,N_10648);
or U10812 (N_10812,N_10635,N_10726);
nand U10813 (N_10813,N_10662,N_10735);
or U10814 (N_10814,N_10730,N_10743);
nor U10815 (N_10815,N_10659,N_10711);
nand U10816 (N_10816,N_10734,N_10720);
and U10817 (N_10817,N_10678,N_10645);
nor U10818 (N_10818,N_10676,N_10718);
or U10819 (N_10819,N_10665,N_10671);
xor U10820 (N_10820,N_10688,N_10738);
or U10821 (N_10821,N_10726,N_10666);
or U10822 (N_10822,N_10703,N_10646);
nor U10823 (N_10823,N_10656,N_10734);
or U10824 (N_10824,N_10661,N_10677);
or U10825 (N_10825,N_10658,N_10727);
or U10826 (N_10826,N_10681,N_10738);
nor U10827 (N_10827,N_10716,N_10724);
or U10828 (N_10828,N_10732,N_10683);
nor U10829 (N_10829,N_10635,N_10701);
and U10830 (N_10830,N_10707,N_10727);
nor U10831 (N_10831,N_10683,N_10730);
xor U10832 (N_10832,N_10724,N_10677);
xnor U10833 (N_10833,N_10749,N_10745);
nand U10834 (N_10834,N_10727,N_10737);
and U10835 (N_10835,N_10703,N_10746);
and U10836 (N_10836,N_10635,N_10641);
or U10837 (N_10837,N_10685,N_10715);
and U10838 (N_10838,N_10686,N_10660);
nor U10839 (N_10839,N_10731,N_10642);
and U10840 (N_10840,N_10715,N_10719);
nand U10841 (N_10841,N_10714,N_10687);
nand U10842 (N_10842,N_10633,N_10682);
nand U10843 (N_10843,N_10741,N_10648);
xnor U10844 (N_10844,N_10733,N_10736);
nor U10845 (N_10845,N_10718,N_10632);
xnor U10846 (N_10846,N_10667,N_10650);
nor U10847 (N_10847,N_10748,N_10715);
and U10848 (N_10848,N_10724,N_10744);
xnor U10849 (N_10849,N_10679,N_10738);
or U10850 (N_10850,N_10625,N_10695);
nor U10851 (N_10851,N_10686,N_10668);
nand U10852 (N_10852,N_10712,N_10635);
nand U10853 (N_10853,N_10668,N_10685);
nand U10854 (N_10854,N_10734,N_10718);
xor U10855 (N_10855,N_10735,N_10709);
nand U10856 (N_10856,N_10648,N_10739);
xor U10857 (N_10857,N_10667,N_10672);
xnor U10858 (N_10858,N_10662,N_10676);
xnor U10859 (N_10859,N_10693,N_10665);
nor U10860 (N_10860,N_10708,N_10680);
or U10861 (N_10861,N_10678,N_10661);
and U10862 (N_10862,N_10722,N_10708);
nand U10863 (N_10863,N_10717,N_10671);
or U10864 (N_10864,N_10643,N_10705);
nand U10865 (N_10865,N_10681,N_10697);
xor U10866 (N_10866,N_10722,N_10680);
nor U10867 (N_10867,N_10658,N_10670);
and U10868 (N_10868,N_10647,N_10733);
and U10869 (N_10869,N_10728,N_10694);
and U10870 (N_10870,N_10691,N_10695);
nand U10871 (N_10871,N_10728,N_10690);
xor U10872 (N_10872,N_10662,N_10644);
and U10873 (N_10873,N_10641,N_10677);
or U10874 (N_10874,N_10647,N_10732);
nand U10875 (N_10875,N_10827,N_10768);
or U10876 (N_10876,N_10817,N_10838);
nor U10877 (N_10877,N_10757,N_10848);
nand U10878 (N_10878,N_10861,N_10826);
or U10879 (N_10879,N_10829,N_10816);
nor U10880 (N_10880,N_10799,N_10845);
nand U10881 (N_10881,N_10855,N_10831);
or U10882 (N_10882,N_10794,N_10793);
or U10883 (N_10883,N_10869,N_10830);
or U10884 (N_10884,N_10772,N_10778);
or U10885 (N_10885,N_10786,N_10860);
xnor U10886 (N_10886,N_10850,N_10767);
or U10887 (N_10887,N_10873,N_10763);
nor U10888 (N_10888,N_10854,N_10821);
xnor U10889 (N_10889,N_10849,N_10784);
nand U10890 (N_10890,N_10865,N_10753);
and U10891 (N_10891,N_10758,N_10800);
nand U10892 (N_10892,N_10787,N_10864);
or U10893 (N_10893,N_10777,N_10774);
or U10894 (N_10894,N_10859,N_10790);
nor U10895 (N_10895,N_10792,N_10762);
nand U10896 (N_10896,N_10773,N_10871);
nand U10897 (N_10897,N_10853,N_10847);
nand U10898 (N_10898,N_10818,N_10771);
or U10899 (N_10899,N_10825,N_10781);
and U10900 (N_10900,N_10857,N_10805);
nor U10901 (N_10901,N_10775,N_10810);
or U10902 (N_10902,N_10841,N_10863);
or U10903 (N_10903,N_10776,N_10755);
and U10904 (N_10904,N_10851,N_10788);
or U10905 (N_10905,N_10812,N_10785);
nor U10906 (N_10906,N_10796,N_10837);
and U10907 (N_10907,N_10872,N_10867);
nand U10908 (N_10908,N_10836,N_10823);
or U10909 (N_10909,N_10766,N_10783);
nor U10910 (N_10910,N_10822,N_10807);
xor U10911 (N_10911,N_10751,N_10874);
nor U10912 (N_10912,N_10820,N_10814);
nand U10913 (N_10913,N_10804,N_10824);
nor U10914 (N_10914,N_10782,N_10819);
nor U10915 (N_10915,N_10770,N_10866);
nand U10916 (N_10916,N_10808,N_10862);
nor U10917 (N_10917,N_10843,N_10809);
nor U10918 (N_10918,N_10846,N_10835);
nand U10919 (N_10919,N_10828,N_10858);
and U10920 (N_10920,N_10833,N_10815);
and U10921 (N_10921,N_10842,N_10780);
and U10922 (N_10922,N_10868,N_10765);
or U10923 (N_10923,N_10761,N_10752);
nor U10924 (N_10924,N_10795,N_10839);
nor U10925 (N_10925,N_10813,N_10803);
xnor U10926 (N_10926,N_10779,N_10797);
nand U10927 (N_10927,N_10806,N_10759);
or U10928 (N_10928,N_10791,N_10789);
and U10929 (N_10929,N_10754,N_10811);
xor U10930 (N_10930,N_10834,N_10852);
nor U10931 (N_10931,N_10844,N_10856);
nor U10932 (N_10932,N_10769,N_10798);
or U10933 (N_10933,N_10832,N_10750);
nor U10934 (N_10934,N_10802,N_10760);
or U10935 (N_10935,N_10764,N_10870);
xor U10936 (N_10936,N_10840,N_10756);
nand U10937 (N_10937,N_10801,N_10862);
nor U10938 (N_10938,N_10787,N_10869);
nand U10939 (N_10939,N_10855,N_10846);
or U10940 (N_10940,N_10799,N_10798);
nor U10941 (N_10941,N_10855,N_10809);
or U10942 (N_10942,N_10832,N_10840);
nand U10943 (N_10943,N_10797,N_10842);
xnor U10944 (N_10944,N_10827,N_10799);
nand U10945 (N_10945,N_10867,N_10834);
nor U10946 (N_10946,N_10807,N_10801);
nor U10947 (N_10947,N_10772,N_10766);
nand U10948 (N_10948,N_10776,N_10835);
xor U10949 (N_10949,N_10782,N_10812);
or U10950 (N_10950,N_10793,N_10858);
nand U10951 (N_10951,N_10829,N_10856);
and U10952 (N_10952,N_10825,N_10759);
nor U10953 (N_10953,N_10758,N_10812);
nor U10954 (N_10954,N_10786,N_10792);
or U10955 (N_10955,N_10861,N_10834);
nor U10956 (N_10956,N_10806,N_10834);
nand U10957 (N_10957,N_10817,N_10782);
nor U10958 (N_10958,N_10752,N_10765);
nor U10959 (N_10959,N_10868,N_10756);
and U10960 (N_10960,N_10767,N_10774);
xor U10961 (N_10961,N_10825,N_10789);
nand U10962 (N_10962,N_10867,N_10791);
nor U10963 (N_10963,N_10832,N_10837);
xnor U10964 (N_10964,N_10788,N_10756);
nor U10965 (N_10965,N_10873,N_10844);
and U10966 (N_10966,N_10849,N_10844);
nor U10967 (N_10967,N_10837,N_10755);
or U10968 (N_10968,N_10792,N_10870);
or U10969 (N_10969,N_10797,N_10753);
xnor U10970 (N_10970,N_10787,N_10865);
xnor U10971 (N_10971,N_10856,N_10755);
nor U10972 (N_10972,N_10835,N_10778);
nand U10973 (N_10973,N_10750,N_10873);
nor U10974 (N_10974,N_10849,N_10766);
nor U10975 (N_10975,N_10800,N_10785);
nand U10976 (N_10976,N_10799,N_10802);
xnor U10977 (N_10977,N_10807,N_10769);
and U10978 (N_10978,N_10796,N_10819);
nand U10979 (N_10979,N_10794,N_10805);
or U10980 (N_10980,N_10844,N_10826);
xor U10981 (N_10981,N_10819,N_10804);
nor U10982 (N_10982,N_10850,N_10759);
or U10983 (N_10983,N_10783,N_10853);
or U10984 (N_10984,N_10820,N_10811);
nor U10985 (N_10985,N_10763,N_10836);
nor U10986 (N_10986,N_10774,N_10803);
and U10987 (N_10987,N_10848,N_10861);
xor U10988 (N_10988,N_10781,N_10816);
xnor U10989 (N_10989,N_10750,N_10776);
xnor U10990 (N_10990,N_10753,N_10764);
nand U10991 (N_10991,N_10847,N_10830);
and U10992 (N_10992,N_10836,N_10778);
and U10993 (N_10993,N_10857,N_10752);
or U10994 (N_10994,N_10792,N_10832);
nor U10995 (N_10995,N_10838,N_10787);
xor U10996 (N_10996,N_10798,N_10871);
or U10997 (N_10997,N_10803,N_10753);
xor U10998 (N_10998,N_10831,N_10795);
nand U10999 (N_10999,N_10794,N_10763);
or U11000 (N_11000,N_10910,N_10929);
xnor U11001 (N_11001,N_10912,N_10939);
nor U11002 (N_11002,N_10914,N_10889);
or U11003 (N_11003,N_10954,N_10883);
and U11004 (N_11004,N_10989,N_10995);
nor U11005 (N_11005,N_10934,N_10900);
nor U11006 (N_11006,N_10973,N_10955);
nand U11007 (N_11007,N_10878,N_10977);
or U11008 (N_11008,N_10880,N_10935);
nor U11009 (N_11009,N_10923,N_10894);
or U11010 (N_11010,N_10930,N_10927);
or U11011 (N_11011,N_10957,N_10907);
and U11012 (N_11012,N_10921,N_10959);
nor U11013 (N_11013,N_10985,N_10932);
nand U11014 (N_11014,N_10950,N_10975);
or U11015 (N_11015,N_10951,N_10982);
nand U11016 (N_11016,N_10958,N_10956);
xnor U11017 (N_11017,N_10941,N_10903);
nand U11018 (N_11018,N_10965,N_10897);
or U11019 (N_11019,N_10997,N_10986);
nor U11020 (N_11020,N_10901,N_10919);
xor U11021 (N_11021,N_10996,N_10931);
nor U11022 (N_11022,N_10972,N_10981);
xnor U11023 (N_11023,N_10928,N_10979);
nand U11024 (N_11024,N_10940,N_10902);
xnor U11025 (N_11025,N_10879,N_10938);
nand U11026 (N_11026,N_10968,N_10875);
and U11027 (N_11027,N_10966,N_10963);
nand U11028 (N_11028,N_10876,N_10918);
xor U11029 (N_11029,N_10882,N_10961);
nor U11030 (N_11030,N_10917,N_10906);
or U11031 (N_11031,N_10896,N_10885);
nand U11032 (N_11032,N_10887,N_10913);
or U11033 (N_11033,N_10933,N_10908);
xor U11034 (N_11034,N_10904,N_10969);
and U11035 (N_11035,N_10971,N_10953);
nand U11036 (N_11036,N_10984,N_10895);
and U11037 (N_11037,N_10967,N_10987);
and U11038 (N_11038,N_10909,N_10893);
and U11039 (N_11039,N_10952,N_10964);
nand U11040 (N_11040,N_10920,N_10945);
or U11041 (N_11041,N_10942,N_10947);
nand U11042 (N_11042,N_10898,N_10978);
xnor U11043 (N_11043,N_10992,N_10892);
nor U11044 (N_11044,N_10962,N_10976);
and U11045 (N_11045,N_10974,N_10916);
xnor U11046 (N_11046,N_10946,N_10949);
nor U11047 (N_11047,N_10948,N_10994);
nor U11048 (N_11048,N_10998,N_10915);
nor U11049 (N_11049,N_10911,N_10980);
nor U11050 (N_11050,N_10937,N_10891);
xnor U11051 (N_11051,N_10922,N_10925);
xor U11052 (N_11052,N_10970,N_10936);
nand U11053 (N_11053,N_10899,N_10993);
nor U11054 (N_11054,N_10890,N_10960);
or U11055 (N_11055,N_10999,N_10905);
and U11056 (N_11056,N_10943,N_10884);
nor U11057 (N_11057,N_10990,N_10926);
nand U11058 (N_11058,N_10888,N_10881);
nor U11059 (N_11059,N_10886,N_10924);
nor U11060 (N_11060,N_10991,N_10983);
nor U11061 (N_11061,N_10877,N_10988);
nand U11062 (N_11062,N_10944,N_10979);
and U11063 (N_11063,N_10885,N_10964);
nor U11064 (N_11064,N_10888,N_10926);
and U11065 (N_11065,N_10918,N_10898);
nor U11066 (N_11066,N_10937,N_10941);
or U11067 (N_11067,N_10975,N_10983);
and U11068 (N_11068,N_10997,N_10944);
xor U11069 (N_11069,N_10950,N_10890);
nor U11070 (N_11070,N_10884,N_10921);
or U11071 (N_11071,N_10974,N_10895);
xnor U11072 (N_11072,N_10962,N_10910);
or U11073 (N_11073,N_10918,N_10940);
nor U11074 (N_11074,N_10982,N_10944);
or U11075 (N_11075,N_10979,N_10912);
or U11076 (N_11076,N_10992,N_10900);
nand U11077 (N_11077,N_10991,N_10971);
or U11078 (N_11078,N_10875,N_10918);
nand U11079 (N_11079,N_10964,N_10934);
nor U11080 (N_11080,N_10990,N_10989);
and U11081 (N_11081,N_10915,N_10934);
and U11082 (N_11082,N_10967,N_10902);
and U11083 (N_11083,N_10885,N_10914);
nor U11084 (N_11084,N_10917,N_10955);
and U11085 (N_11085,N_10945,N_10968);
and U11086 (N_11086,N_10924,N_10936);
and U11087 (N_11087,N_10912,N_10984);
xor U11088 (N_11088,N_10995,N_10973);
and U11089 (N_11089,N_10946,N_10888);
xnor U11090 (N_11090,N_10893,N_10964);
xor U11091 (N_11091,N_10908,N_10913);
nor U11092 (N_11092,N_10927,N_10917);
nor U11093 (N_11093,N_10898,N_10963);
nor U11094 (N_11094,N_10919,N_10946);
nor U11095 (N_11095,N_10993,N_10967);
nor U11096 (N_11096,N_10988,N_10900);
xnor U11097 (N_11097,N_10917,N_10911);
nor U11098 (N_11098,N_10998,N_10971);
or U11099 (N_11099,N_10953,N_10877);
and U11100 (N_11100,N_10914,N_10901);
and U11101 (N_11101,N_10880,N_10958);
and U11102 (N_11102,N_10901,N_10965);
and U11103 (N_11103,N_10894,N_10882);
nand U11104 (N_11104,N_10986,N_10951);
xnor U11105 (N_11105,N_10906,N_10879);
xnor U11106 (N_11106,N_10887,N_10990);
nand U11107 (N_11107,N_10965,N_10939);
nand U11108 (N_11108,N_10966,N_10893);
xor U11109 (N_11109,N_10973,N_10992);
xnor U11110 (N_11110,N_10960,N_10891);
xor U11111 (N_11111,N_10879,N_10885);
xor U11112 (N_11112,N_10936,N_10942);
or U11113 (N_11113,N_10990,N_10890);
nand U11114 (N_11114,N_10959,N_10881);
nor U11115 (N_11115,N_10946,N_10951);
or U11116 (N_11116,N_10942,N_10933);
xor U11117 (N_11117,N_10944,N_10991);
and U11118 (N_11118,N_10968,N_10926);
nor U11119 (N_11119,N_10887,N_10916);
or U11120 (N_11120,N_10953,N_10887);
and U11121 (N_11121,N_10932,N_10882);
or U11122 (N_11122,N_10940,N_10986);
nand U11123 (N_11123,N_10931,N_10913);
or U11124 (N_11124,N_10967,N_10935);
and U11125 (N_11125,N_11048,N_11098);
xor U11126 (N_11126,N_11063,N_11100);
and U11127 (N_11127,N_11122,N_11019);
nor U11128 (N_11128,N_11031,N_11023);
xor U11129 (N_11129,N_11039,N_11104);
and U11130 (N_11130,N_11083,N_11054);
xnor U11131 (N_11131,N_11041,N_11058);
and U11132 (N_11132,N_11084,N_11050);
xor U11133 (N_11133,N_11094,N_11116);
nor U11134 (N_11134,N_11038,N_11096);
or U11135 (N_11135,N_11042,N_11012);
nor U11136 (N_11136,N_11073,N_11061);
nor U11137 (N_11137,N_11005,N_11066);
xnor U11138 (N_11138,N_11027,N_11106);
nor U11139 (N_11139,N_11044,N_11006);
xnor U11140 (N_11140,N_11060,N_11033);
xor U11141 (N_11141,N_11117,N_11085);
nor U11142 (N_11142,N_11046,N_11010);
and U11143 (N_11143,N_11053,N_11108);
or U11144 (N_11144,N_11065,N_11112);
nand U11145 (N_11145,N_11037,N_11043);
or U11146 (N_11146,N_11072,N_11062);
or U11147 (N_11147,N_11001,N_11086);
or U11148 (N_11148,N_11013,N_11034);
or U11149 (N_11149,N_11091,N_11078);
nor U11150 (N_11150,N_11089,N_11113);
nand U11151 (N_11151,N_11035,N_11057);
and U11152 (N_11152,N_11118,N_11022);
xor U11153 (N_11153,N_11103,N_11014);
or U11154 (N_11154,N_11095,N_11101);
and U11155 (N_11155,N_11105,N_11099);
or U11156 (N_11156,N_11087,N_11024);
nor U11157 (N_11157,N_11121,N_11088);
or U11158 (N_11158,N_11081,N_11120);
nor U11159 (N_11159,N_11097,N_11002);
xor U11160 (N_11160,N_11090,N_11026);
xor U11161 (N_11161,N_11052,N_11047);
xor U11162 (N_11162,N_11068,N_11036);
nand U11163 (N_11163,N_11076,N_11055);
nor U11164 (N_11164,N_11075,N_11074);
or U11165 (N_11165,N_11124,N_11000);
and U11166 (N_11166,N_11114,N_11107);
xor U11167 (N_11167,N_11071,N_11069);
nand U11168 (N_11168,N_11020,N_11092);
xor U11169 (N_11169,N_11059,N_11018);
xor U11170 (N_11170,N_11030,N_11003);
nand U11171 (N_11171,N_11007,N_11040);
nand U11172 (N_11172,N_11110,N_11045);
xor U11173 (N_11173,N_11025,N_11017);
xor U11174 (N_11174,N_11082,N_11021);
nand U11175 (N_11175,N_11016,N_11067);
or U11176 (N_11176,N_11079,N_11111);
xor U11177 (N_11177,N_11009,N_11008);
or U11178 (N_11178,N_11032,N_11011);
or U11179 (N_11179,N_11056,N_11049);
nand U11180 (N_11180,N_11119,N_11070);
nand U11181 (N_11181,N_11080,N_11109);
and U11182 (N_11182,N_11029,N_11077);
nor U11183 (N_11183,N_11028,N_11051);
nand U11184 (N_11184,N_11115,N_11093);
nor U11185 (N_11185,N_11004,N_11123);
nor U11186 (N_11186,N_11102,N_11015);
or U11187 (N_11187,N_11064,N_11098);
nand U11188 (N_11188,N_11047,N_11070);
xnor U11189 (N_11189,N_11110,N_11084);
xnor U11190 (N_11190,N_11051,N_11035);
nor U11191 (N_11191,N_11103,N_11018);
xor U11192 (N_11192,N_11087,N_11070);
or U11193 (N_11193,N_11031,N_11025);
and U11194 (N_11194,N_11008,N_11053);
nor U11195 (N_11195,N_11103,N_11072);
nand U11196 (N_11196,N_11022,N_11078);
nand U11197 (N_11197,N_11056,N_11120);
xnor U11198 (N_11198,N_11089,N_11052);
or U11199 (N_11199,N_11062,N_11058);
nand U11200 (N_11200,N_11051,N_11067);
and U11201 (N_11201,N_11081,N_11055);
xnor U11202 (N_11202,N_11107,N_11039);
and U11203 (N_11203,N_11045,N_11044);
nand U11204 (N_11204,N_11005,N_11000);
and U11205 (N_11205,N_11076,N_11047);
xor U11206 (N_11206,N_11076,N_11108);
and U11207 (N_11207,N_11029,N_11045);
and U11208 (N_11208,N_11103,N_11050);
xor U11209 (N_11209,N_11022,N_11069);
or U11210 (N_11210,N_11108,N_11043);
or U11211 (N_11211,N_11027,N_11080);
and U11212 (N_11212,N_11001,N_11078);
and U11213 (N_11213,N_11070,N_11062);
nand U11214 (N_11214,N_11092,N_11094);
xnor U11215 (N_11215,N_11065,N_11100);
or U11216 (N_11216,N_11106,N_11119);
nand U11217 (N_11217,N_11013,N_11062);
xnor U11218 (N_11218,N_11042,N_11077);
xor U11219 (N_11219,N_11077,N_11112);
nor U11220 (N_11220,N_11085,N_11020);
xnor U11221 (N_11221,N_11100,N_11033);
or U11222 (N_11222,N_11094,N_11046);
xor U11223 (N_11223,N_11099,N_11070);
nand U11224 (N_11224,N_11118,N_11105);
and U11225 (N_11225,N_11010,N_11009);
and U11226 (N_11226,N_11051,N_11054);
nor U11227 (N_11227,N_11038,N_11052);
xor U11228 (N_11228,N_11071,N_11047);
nand U11229 (N_11229,N_11043,N_11045);
or U11230 (N_11230,N_11017,N_11061);
and U11231 (N_11231,N_11068,N_11013);
xor U11232 (N_11232,N_11113,N_11025);
nand U11233 (N_11233,N_11006,N_11032);
or U11234 (N_11234,N_11059,N_11048);
nand U11235 (N_11235,N_11018,N_11108);
nor U11236 (N_11236,N_11020,N_11051);
or U11237 (N_11237,N_11104,N_11119);
xor U11238 (N_11238,N_11076,N_11015);
nand U11239 (N_11239,N_11077,N_11035);
and U11240 (N_11240,N_11096,N_11056);
nand U11241 (N_11241,N_11111,N_11098);
nand U11242 (N_11242,N_11077,N_11054);
xor U11243 (N_11243,N_11071,N_11043);
nand U11244 (N_11244,N_11077,N_11107);
and U11245 (N_11245,N_11076,N_11007);
xnor U11246 (N_11246,N_11045,N_11054);
and U11247 (N_11247,N_11120,N_11030);
nand U11248 (N_11248,N_11098,N_11091);
nand U11249 (N_11249,N_11031,N_11077);
nand U11250 (N_11250,N_11189,N_11224);
nand U11251 (N_11251,N_11202,N_11213);
and U11252 (N_11252,N_11248,N_11196);
xor U11253 (N_11253,N_11186,N_11172);
xnor U11254 (N_11254,N_11241,N_11203);
or U11255 (N_11255,N_11180,N_11205);
nor U11256 (N_11256,N_11201,N_11144);
nand U11257 (N_11257,N_11212,N_11195);
xnor U11258 (N_11258,N_11245,N_11228);
and U11259 (N_11259,N_11183,N_11239);
and U11260 (N_11260,N_11139,N_11171);
and U11261 (N_11261,N_11226,N_11176);
or U11262 (N_11262,N_11188,N_11135);
xnor U11263 (N_11263,N_11147,N_11193);
nand U11264 (N_11264,N_11198,N_11225);
or U11265 (N_11265,N_11136,N_11143);
nand U11266 (N_11266,N_11128,N_11243);
nor U11267 (N_11267,N_11204,N_11238);
nor U11268 (N_11268,N_11210,N_11170);
or U11269 (N_11269,N_11217,N_11154);
xor U11270 (N_11270,N_11129,N_11133);
nor U11271 (N_11271,N_11234,N_11148);
and U11272 (N_11272,N_11216,N_11167);
and U11273 (N_11273,N_11126,N_11207);
and U11274 (N_11274,N_11229,N_11182);
and U11275 (N_11275,N_11232,N_11165);
xnor U11276 (N_11276,N_11208,N_11191);
and U11277 (N_11277,N_11231,N_11247);
or U11278 (N_11278,N_11141,N_11174);
nand U11279 (N_11279,N_11240,N_11192);
nor U11280 (N_11280,N_11199,N_11236);
nand U11281 (N_11281,N_11160,N_11184);
or U11282 (N_11282,N_11146,N_11233);
or U11283 (N_11283,N_11162,N_11220);
or U11284 (N_11284,N_11166,N_11175);
xor U11285 (N_11285,N_11221,N_11214);
and U11286 (N_11286,N_11242,N_11177);
or U11287 (N_11287,N_11159,N_11249);
nand U11288 (N_11288,N_11169,N_11125);
and U11289 (N_11289,N_11246,N_11215);
or U11290 (N_11290,N_11211,N_11209);
xnor U11291 (N_11291,N_11137,N_11244);
xor U11292 (N_11292,N_11150,N_11230);
nand U11293 (N_11293,N_11142,N_11219);
nor U11294 (N_11294,N_11161,N_11178);
nand U11295 (N_11295,N_11235,N_11156);
nand U11296 (N_11296,N_11153,N_11151);
or U11297 (N_11297,N_11163,N_11206);
nor U11298 (N_11298,N_11185,N_11181);
or U11299 (N_11299,N_11130,N_11179);
xnor U11300 (N_11300,N_11227,N_11223);
nand U11301 (N_11301,N_11200,N_11173);
nor U11302 (N_11302,N_11149,N_11157);
nand U11303 (N_11303,N_11140,N_11197);
and U11304 (N_11304,N_11218,N_11158);
nand U11305 (N_11305,N_11138,N_11190);
nor U11306 (N_11306,N_11237,N_11134);
nor U11307 (N_11307,N_11131,N_11155);
nand U11308 (N_11308,N_11222,N_11132);
nand U11309 (N_11309,N_11168,N_11194);
or U11310 (N_11310,N_11187,N_11145);
nand U11311 (N_11311,N_11164,N_11127);
or U11312 (N_11312,N_11152,N_11198);
or U11313 (N_11313,N_11145,N_11180);
xor U11314 (N_11314,N_11234,N_11196);
or U11315 (N_11315,N_11137,N_11185);
nor U11316 (N_11316,N_11205,N_11219);
xnor U11317 (N_11317,N_11226,N_11221);
and U11318 (N_11318,N_11210,N_11219);
or U11319 (N_11319,N_11245,N_11157);
and U11320 (N_11320,N_11126,N_11228);
and U11321 (N_11321,N_11145,N_11144);
or U11322 (N_11322,N_11236,N_11227);
xnor U11323 (N_11323,N_11126,N_11143);
nor U11324 (N_11324,N_11130,N_11199);
nand U11325 (N_11325,N_11220,N_11204);
nor U11326 (N_11326,N_11163,N_11155);
nor U11327 (N_11327,N_11219,N_11206);
nor U11328 (N_11328,N_11168,N_11127);
nand U11329 (N_11329,N_11168,N_11202);
nor U11330 (N_11330,N_11143,N_11189);
nand U11331 (N_11331,N_11155,N_11232);
or U11332 (N_11332,N_11136,N_11213);
nand U11333 (N_11333,N_11151,N_11243);
or U11334 (N_11334,N_11149,N_11133);
or U11335 (N_11335,N_11125,N_11208);
and U11336 (N_11336,N_11226,N_11162);
xnor U11337 (N_11337,N_11159,N_11133);
or U11338 (N_11338,N_11127,N_11209);
xnor U11339 (N_11339,N_11210,N_11156);
or U11340 (N_11340,N_11237,N_11222);
xnor U11341 (N_11341,N_11247,N_11178);
nor U11342 (N_11342,N_11145,N_11211);
and U11343 (N_11343,N_11185,N_11239);
xnor U11344 (N_11344,N_11150,N_11219);
nor U11345 (N_11345,N_11165,N_11193);
and U11346 (N_11346,N_11165,N_11133);
nand U11347 (N_11347,N_11217,N_11197);
nand U11348 (N_11348,N_11245,N_11206);
xor U11349 (N_11349,N_11192,N_11158);
and U11350 (N_11350,N_11125,N_11211);
xnor U11351 (N_11351,N_11219,N_11237);
nor U11352 (N_11352,N_11225,N_11180);
nor U11353 (N_11353,N_11151,N_11247);
nand U11354 (N_11354,N_11128,N_11201);
nor U11355 (N_11355,N_11248,N_11165);
or U11356 (N_11356,N_11133,N_11138);
or U11357 (N_11357,N_11135,N_11241);
xnor U11358 (N_11358,N_11246,N_11247);
nor U11359 (N_11359,N_11224,N_11223);
nor U11360 (N_11360,N_11131,N_11195);
nand U11361 (N_11361,N_11220,N_11154);
and U11362 (N_11362,N_11234,N_11147);
nand U11363 (N_11363,N_11212,N_11196);
nand U11364 (N_11364,N_11237,N_11175);
nor U11365 (N_11365,N_11189,N_11163);
or U11366 (N_11366,N_11131,N_11192);
xor U11367 (N_11367,N_11206,N_11215);
nand U11368 (N_11368,N_11212,N_11186);
or U11369 (N_11369,N_11171,N_11161);
and U11370 (N_11370,N_11134,N_11226);
xnor U11371 (N_11371,N_11205,N_11238);
and U11372 (N_11372,N_11172,N_11184);
and U11373 (N_11373,N_11127,N_11228);
or U11374 (N_11374,N_11203,N_11132);
xor U11375 (N_11375,N_11332,N_11352);
nand U11376 (N_11376,N_11364,N_11368);
and U11377 (N_11377,N_11330,N_11314);
xor U11378 (N_11378,N_11305,N_11286);
nand U11379 (N_11379,N_11353,N_11300);
xnor U11380 (N_11380,N_11251,N_11267);
or U11381 (N_11381,N_11309,N_11284);
xor U11382 (N_11382,N_11321,N_11256);
and U11383 (N_11383,N_11301,N_11273);
xor U11384 (N_11384,N_11366,N_11354);
or U11385 (N_11385,N_11289,N_11265);
or U11386 (N_11386,N_11329,N_11262);
nor U11387 (N_11387,N_11250,N_11363);
nor U11388 (N_11388,N_11374,N_11313);
and U11389 (N_11389,N_11281,N_11346);
xnor U11390 (N_11390,N_11343,N_11272);
xor U11391 (N_11391,N_11299,N_11358);
and U11392 (N_11392,N_11258,N_11295);
and U11393 (N_11393,N_11342,N_11348);
nand U11394 (N_11394,N_11335,N_11319);
nand U11395 (N_11395,N_11345,N_11277);
xnor U11396 (N_11396,N_11261,N_11336);
xor U11397 (N_11397,N_11291,N_11287);
xnor U11398 (N_11398,N_11365,N_11280);
or U11399 (N_11399,N_11326,N_11255);
xnor U11400 (N_11400,N_11257,N_11259);
nand U11401 (N_11401,N_11292,N_11316);
xor U11402 (N_11402,N_11317,N_11323);
xnor U11403 (N_11403,N_11266,N_11327);
and U11404 (N_11404,N_11328,N_11367);
or U11405 (N_11405,N_11351,N_11304);
nand U11406 (N_11406,N_11315,N_11362);
and U11407 (N_11407,N_11271,N_11361);
and U11408 (N_11408,N_11338,N_11337);
nor U11409 (N_11409,N_11310,N_11322);
and U11410 (N_11410,N_11331,N_11294);
nand U11411 (N_11411,N_11307,N_11339);
or U11412 (N_11412,N_11333,N_11276);
nand U11413 (N_11413,N_11357,N_11360);
nand U11414 (N_11414,N_11268,N_11285);
xor U11415 (N_11415,N_11311,N_11370);
nor U11416 (N_11416,N_11298,N_11350);
nand U11417 (N_11417,N_11279,N_11274);
nor U11418 (N_11418,N_11324,N_11369);
and U11419 (N_11419,N_11344,N_11297);
nor U11420 (N_11420,N_11263,N_11355);
or U11421 (N_11421,N_11275,N_11334);
and U11422 (N_11422,N_11264,N_11349);
and U11423 (N_11423,N_11293,N_11260);
nand U11424 (N_11424,N_11347,N_11372);
or U11425 (N_11425,N_11325,N_11269);
or U11426 (N_11426,N_11320,N_11341);
and U11427 (N_11427,N_11283,N_11371);
xnor U11428 (N_11428,N_11270,N_11282);
or U11429 (N_11429,N_11253,N_11359);
or U11430 (N_11430,N_11302,N_11308);
or U11431 (N_11431,N_11340,N_11290);
nand U11432 (N_11432,N_11356,N_11312);
nor U11433 (N_11433,N_11252,N_11303);
and U11434 (N_11434,N_11318,N_11296);
and U11435 (N_11435,N_11306,N_11288);
nor U11436 (N_11436,N_11373,N_11254);
xnor U11437 (N_11437,N_11278,N_11374);
or U11438 (N_11438,N_11293,N_11254);
nor U11439 (N_11439,N_11260,N_11336);
or U11440 (N_11440,N_11363,N_11328);
or U11441 (N_11441,N_11350,N_11287);
and U11442 (N_11442,N_11281,N_11353);
or U11443 (N_11443,N_11296,N_11290);
nand U11444 (N_11444,N_11322,N_11346);
nand U11445 (N_11445,N_11275,N_11286);
or U11446 (N_11446,N_11266,N_11299);
nor U11447 (N_11447,N_11347,N_11373);
and U11448 (N_11448,N_11309,N_11271);
or U11449 (N_11449,N_11303,N_11321);
xor U11450 (N_11450,N_11371,N_11284);
nor U11451 (N_11451,N_11309,N_11278);
nand U11452 (N_11452,N_11259,N_11363);
and U11453 (N_11453,N_11289,N_11319);
xnor U11454 (N_11454,N_11278,N_11299);
or U11455 (N_11455,N_11260,N_11323);
or U11456 (N_11456,N_11259,N_11324);
xor U11457 (N_11457,N_11273,N_11255);
nand U11458 (N_11458,N_11365,N_11291);
and U11459 (N_11459,N_11374,N_11342);
nand U11460 (N_11460,N_11296,N_11310);
xor U11461 (N_11461,N_11308,N_11310);
and U11462 (N_11462,N_11257,N_11365);
xor U11463 (N_11463,N_11300,N_11272);
or U11464 (N_11464,N_11250,N_11296);
xor U11465 (N_11465,N_11301,N_11265);
xor U11466 (N_11466,N_11361,N_11257);
or U11467 (N_11467,N_11283,N_11287);
nand U11468 (N_11468,N_11251,N_11287);
and U11469 (N_11469,N_11352,N_11315);
or U11470 (N_11470,N_11258,N_11259);
or U11471 (N_11471,N_11252,N_11261);
nand U11472 (N_11472,N_11296,N_11251);
or U11473 (N_11473,N_11310,N_11333);
nand U11474 (N_11474,N_11251,N_11326);
and U11475 (N_11475,N_11307,N_11344);
nor U11476 (N_11476,N_11281,N_11336);
or U11477 (N_11477,N_11298,N_11303);
and U11478 (N_11478,N_11294,N_11362);
xnor U11479 (N_11479,N_11347,N_11297);
or U11480 (N_11480,N_11374,N_11369);
nand U11481 (N_11481,N_11284,N_11322);
xor U11482 (N_11482,N_11313,N_11281);
and U11483 (N_11483,N_11314,N_11298);
xnor U11484 (N_11484,N_11371,N_11374);
nand U11485 (N_11485,N_11278,N_11272);
and U11486 (N_11486,N_11373,N_11261);
xnor U11487 (N_11487,N_11303,N_11295);
and U11488 (N_11488,N_11331,N_11322);
xnor U11489 (N_11489,N_11370,N_11275);
nand U11490 (N_11490,N_11356,N_11270);
and U11491 (N_11491,N_11331,N_11297);
or U11492 (N_11492,N_11292,N_11273);
xor U11493 (N_11493,N_11253,N_11314);
xnor U11494 (N_11494,N_11285,N_11368);
xnor U11495 (N_11495,N_11346,N_11332);
nor U11496 (N_11496,N_11304,N_11250);
or U11497 (N_11497,N_11301,N_11323);
xor U11498 (N_11498,N_11373,N_11328);
nand U11499 (N_11499,N_11370,N_11318);
and U11500 (N_11500,N_11459,N_11472);
xor U11501 (N_11501,N_11456,N_11403);
or U11502 (N_11502,N_11441,N_11394);
or U11503 (N_11503,N_11471,N_11436);
nor U11504 (N_11504,N_11484,N_11473);
or U11505 (N_11505,N_11375,N_11460);
xor U11506 (N_11506,N_11415,N_11464);
nand U11507 (N_11507,N_11499,N_11498);
nor U11508 (N_11508,N_11414,N_11440);
nor U11509 (N_11509,N_11425,N_11385);
or U11510 (N_11510,N_11407,N_11439);
xor U11511 (N_11511,N_11379,N_11423);
nand U11512 (N_11512,N_11452,N_11491);
and U11513 (N_11513,N_11389,N_11479);
or U11514 (N_11514,N_11381,N_11421);
nand U11515 (N_11515,N_11469,N_11477);
and U11516 (N_11516,N_11443,N_11390);
or U11517 (N_11517,N_11493,N_11466);
nor U11518 (N_11518,N_11435,N_11497);
xor U11519 (N_11519,N_11395,N_11427);
xor U11520 (N_11520,N_11400,N_11412);
xor U11521 (N_11521,N_11406,N_11428);
nor U11522 (N_11522,N_11426,N_11486);
xnor U11523 (N_11523,N_11495,N_11383);
xor U11524 (N_11524,N_11392,N_11378);
or U11525 (N_11525,N_11384,N_11430);
or U11526 (N_11526,N_11463,N_11418);
xnor U11527 (N_11527,N_11442,N_11462);
nor U11528 (N_11528,N_11481,N_11470);
or U11529 (N_11529,N_11387,N_11487);
or U11530 (N_11530,N_11434,N_11446);
xor U11531 (N_11531,N_11496,N_11417);
or U11532 (N_11532,N_11444,N_11405);
or U11533 (N_11533,N_11376,N_11492);
xor U11534 (N_11534,N_11408,N_11396);
nand U11535 (N_11535,N_11401,N_11388);
or U11536 (N_11536,N_11454,N_11437);
nand U11537 (N_11537,N_11393,N_11453);
nor U11538 (N_11538,N_11494,N_11377);
or U11539 (N_11539,N_11465,N_11476);
xnor U11540 (N_11540,N_11447,N_11419);
and U11541 (N_11541,N_11380,N_11448);
xnor U11542 (N_11542,N_11409,N_11404);
xor U11543 (N_11543,N_11483,N_11451);
nor U11544 (N_11544,N_11457,N_11485);
nor U11545 (N_11545,N_11475,N_11482);
or U11546 (N_11546,N_11391,N_11468);
xor U11547 (N_11547,N_11386,N_11413);
nor U11548 (N_11548,N_11429,N_11445);
nor U11549 (N_11549,N_11488,N_11422);
xor U11550 (N_11550,N_11467,N_11416);
xor U11551 (N_11551,N_11458,N_11461);
xor U11552 (N_11552,N_11474,N_11398);
nor U11553 (N_11553,N_11382,N_11478);
xor U11554 (N_11554,N_11489,N_11399);
xnor U11555 (N_11555,N_11420,N_11438);
nand U11556 (N_11556,N_11431,N_11402);
xor U11557 (N_11557,N_11432,N_11411);
or U11558 (N_11558,N_11490,N_11424);
or U11559 (N_11559,N_11455,N_11410);
nand U11560 (N_11560,N_11480,N_11433);
or U11561 (N_11561,N_11449,N_11397);
xnor U11562 (N_11562,N_11450,N_11398);
or U11563 (N_11563,N_11454,N_11477);
nand U11564 (N_11564,N_11499,N_11448);
and U11565 (N_11565,N_11394,N_11402);
nand U11566 (N_11566,N_11462,N_11426);
or U11567 (N_11567,N_11396,N_11415);
nor U11568 (N_11568,N_11491,N_11485);
nand U11569 (N_11569,N_11399,N_11448);
or U11570 (N_11570,N_11451,N_11498);
and U11571 (N_11571,N_11402,N_11466);
nor U11572 (N_11572,N_11453,N_11431);
nand U11573 (N_11573,N_11453,N_11456);
xor U11574 (N_11574,N_11462,N_11489);
xnor U11575 (N_11575,N_11390,N_11420);
and U11576 (N_11576,N_11435,N_11490);
nor U11577 (N_11577,N_11442,N_11467);
xnor U11578 (N_11578,N_11431,N_11495);
nand U11579 (N_11579,N_11495,N_11455);
nand U11580 (N_11580,N_11470,N_11485);
nor U11581 (N_11581,N_11395,N_11439);
or U11582 (N_11582,N_11491,N_11388);
or U11583 (N_11583,N_11441,N_11445);
xnor U11584 (N_11584,N_11499,N_11400);
xnor U11585 (N_11585,N_11490,N_11413);
nand U11586 (N_11586,N_11477,N_11438);
nand U11587 (N_11587,N_11420,N_11395);
xnor U11588 (N_11588,N_11445,N_11409);
xor U11589 (N_11589,N_11436,N_11457);
or U11590 (N_11590,N_11388,N_11493);
nand U11591 (N_11591,N_11462,N_11481);
xnor U11592 (N_11592,N_11480,N_11430);
nor U11593 (N_11593,N_11421,N_11464);
nor U11594 (N_11594,N_11440,N_11448);
nor U11595 (N_11595,N_11408,N_11445);
nand U11596 (N_11596,N_11475,N_11384);
or U11597 (N_11597,N_11380,N_11477);
xnor U11598 (N_11598,N_11428,N_11381);
xor U11599 (N_11599,N_11474,N_11392);
and U11600 (N_11600,N_11456,N_11448);
and U11601 (N_11601,N_11469,N_11409);
xor U11602 (N_11602,N_11413,N_11495);
and U11603 (N_11603,N_11391,N_11485);
nor U11604 (N_11604,N_11495,N_11407);
xor U11605 (N_11605,N_11400,N_11426);
xor U11606 (N_11606,N_11431,N_11439);
or U11607 (N_11607,N_11441,N_11456);
nand U11608 (N_11608,N_11439,N_11447);
or U11609 (N_11609,N_11488,N_11476);
nor U11610 (N_11610,N_11431,N_11472);
nand U11611 (N_11611,N_11440,N_11391);
or U11612 (N_11612,N_11481,N_11419);
nor U11613 (N_11613,N_11399,N_11452);
or U11614 (N_11614,N_11478,N_11376);
nor U11615 (N_11615,N_11390,N_11376);
and U11616 (N_11616,N_11497,N_11450);
nand U11617 (N_11617,N_11444,N_11483);
and U11618 (N_11618,N_11377,N_11397);
and U11619 (N_11619,N_11393,N_11391);
or U11620 (N_11620,N_11475,N_11442);
or U11621 (N_11621,N_11403,N_11457);
or U11622 (N_11622,N_11437,N_11431);
xor U11623 (N_11623,N_11444,N_11436);
and U11624 (N_11624,N_11484,N_11380);
xor U11625 (N_11625,N_11550,N_11598);
and U11626 (N_11626,N_11596,N_11580);
or U11627 (N_11627,N_11532,N_11599);
xnor U11628 (N_11628,N_11518,N_11562);
nand U11629 (N_11629,N_11522,N_11601);
xnor U11630 (N_11630,N_11553,N_11606);
nand U11631 (N_11631,N_11621,N_11503);
and U11632 (N_11632,N_11504,N_11527);
nand U11633 (N_11633,N_11569,N_11520);
and U11634 (N_11634,N_11531,N_11528);
or U11635 (N_11635,N_11567,N_11509);
and U11636 (N_11636,N_11540,N_11536);
nor U11637 (N_11637,N_11558,N_11548);
nand U11638 (N_11638,N_11561,N_11587);
nor U11639 (N_11639,N_11516,N_11534);
xnor U11640 (N_11640,N_11608,N_11568);
nand U11641 (N_11641,N_11581,N_11578);
nor U11642 (N_11642,N_11618,N_11533);
nand U11643 (N_11643,N_11506,N_11595);
nand U11644 (N_11644,N_11538,N_11615);
or U11645 (N_11645,N_11593,N_11526);
and U11646 (N_11646,N_11529,N_11586);
nand U11647 (N_11647,N_11565,N_11576);
and U11648 (N_11648,N_11546,N_11610);
nor U11649 (N_11649,N_11521,N_11566);
xor U11650 (N_11650,N_11537,N_11572);
nor U11651 (N_11651,N_11588,N_11541);
xnor U11652 (N_11652,N_11552,N_11614);
nor U11653 (N_11653,N_11551,N_11560);
or U11654 (N_11654,N_11623,N_11517);
xor U11655 (N_11655,N_11559,N_11555);
nand U11656 (N_11656,N_11571,N_11557);
and U11657 (N_11657,N_11619,N_11563);
nand U11658 (N_11658,N_11508,N_11514);
nand U11659 (N_11659,N_11622,N_11519);
or U11660 (N_11660,N_11554,N_11579);
and U11661 (N_11661,N_11523,N_11613);
nor U11662 (N_11662,N_11539,N_11505);
or U11663 (N_11663,N_11609,N_11510);
and U11664 (N_11664,N_11501,N_11585);
xor U11665 (N_11665,N_11591,N_11545);
nand U11666 (N_11666,N_11597,N_11544);
nand U11667 (N_11667,N_11602,N_11611);
or U11668 (N_11668,N_11574,N_11575);
or U11669 (N_11669,N_11525,N_11589);
nand U11670 (N_11670,N_11583,N_11547);
xor U11671 (N_11671,N_11524,N_11513);
or U11672 (N_11672,N_11584,N_11604);
nor U11673 (N_11673,N_11512,N_11624);
xor U11674 (N_11674,N_11535,N_11592);
xnor U11675 (N_11675,N_11502,N_11600);
nor U11676 (N_11676,N_11612,N_11507);
xnor U11677 (N_11677,N_11500,N_11542);
xnor U11678 (N_11678,N_11573,N_11617);
and U11679 (N_11679,N_11616,N_11530);
nand U11680 (N_11680,N_11577,N_11515);
or U11681 (N_11681,N_11511,N_11594);
and U11682 (N_11682,N_11570,N_11590);
xnor U11683 (N_11683,N_11556,N_11582);
nor U11684 (N_11684,N_11564,N_11607);
nand U11685 (N_11685,N_11603,N_11605);
nor U11686 (N_11686,N_11620,N_11543);
xnor U11687 (N_11687,N_11549,N_11504);
nand U11688 (N_11688,N_11514,N_11607);
xnor U11689 (N_11689,N_11507,N_11593);
and U11690 (N_11690,N_11599,N_11529);
nand U11691 (N_11691,N_11605,N_11511);
nand U11692 (N_11692,N_11525,N_11542);
and U11693 (N_11693,N_11593,N_11509);
nand U11694 (N_11694,N_11521,N_11563);
nand U11695 (N_11695,N_11549,N_11569);
or U11696 (N_11696,N_11522,N_11592);
xor U11697 (N_11697,N_11543,N_11500);
nand U11698 (N_11698,N_11501,N_11576);
xnor U11699 (N_11699,N_11502,N_11543);
nor U11700 (N_11700,N_11546,N_11543);
and U11701 (N_11701,N_11614,N_11607);
nand U11702 (N_11702,N_11535,N_11505);
xor U11703 (N_11703,N_11615,N_11571);
or U11704 (N_11704,N_11559,N_11566);
xor U11705 (N_11705,N_11516,N_11594);
and U11706 (N_11706,N_11622,N_11578);
nand U11707 (N_11707,N_11502,N_11518);
and U11708 (N_11708,N_11530,N_11509);
xor U11709 (N_11709,N_11567,N_11603);
and U11710 (N_11710,N_11528,N_11613);
nor U11711 (N_11711,N_11549,N_11565);
or U11712 (N_11712,N_11615,N_11579);
or U11713 (N_11713,N_11606,N_11605);
nor U11714 (N_11714,N_11586,N_11520);
nor U11715 (N_11715,N_11587,N_11608);
nor U11716 (N_11716,N_11517,N_11564);
and U11717 (N_11717,N_11607,N_11546);
or U11718 (N_11718,N_11507,N_11546);
nand U11719 (N_11719,N_11597,N_11524);
and U11720 (N_11720,N_11506,N_11547);
or U11721 (N_11721,N_11582,N_11599);
nand U11722 (N_11722,N_11574,N_11526);
nor U11723 (N_11723,N_11521,N_11586);
nor U11724 (N_11724,N_11515,N_11563);
nor U11725 (N_11725,N_11576,N_11548);
nand U11726 (N_11726,N_11562,N_11573);
xor U11727 (N_11727,N_11550,N_11527);
xnor U11728 (N_11728,N_11525,N_11586);
nor U11729 (N_11729,N_11593,N_11541);
or U11730 (N_11730,N_11605,N_11519);
nand U11731 (N_11731,N_11600,N_11555);
nand U11732 (N_11732,N_11569,N_11619);
or U11733 (N_11733,N_11526,N_11534);
xor U11734 (N_11734,N_11583,N_11506);
xor U11735 (N_11735,N_11537,N_11594);
and U11736 (N_11736,N_11624,N_11533);
or U11737 (N_11737,N_11579,N_11586);
or U11738 (N_11738,N_11614,N_11571);
xor U11739 (N_11739,N_11537,N_11538);
nand U11740 (N_11740,N_11578,N_11580);
nor U11741 (N_11741,N_11502,N_11612);
nor U11742 (N_11742,N_11556,N_11620);
or U11743 (N_11743,N_11509,N_11588);
xnor U11744 (N_11744,N_11564,N_11583);
xnor U11745 (N_11745,N_11586,N_11511);
nor U11746 (N_11746,N_11504,N_11599);
and U11747 (N_11747,N_11509,N_11514);
nand U11748 (N_11748,N_11526,N_11531);
nand U11749 (N_11749,N_11520,N_11523);
xor U11750 (N_11750,N_11636,N_11630);
nor U11751 (N_11751,N_11635,N_11729);
or U11752 (N_11752,N_11688,N_11678);
or U11753 (N_11753,N_11741,N_11645);
xnor U11754 (N_11754,N_11728,N_11679);
or U11755 (N_11755,N_11745,N_11639);
nand U11756 (N_11756,N_11632,N_11749);
and U11757 (N_11757,N_11656,N_11634);
or U11758 (N_11758,N_11646,N_11627);
nand U11759 (N_11759,N_11697,N_11663);
xor U11760 (N_11760,N_11653,N_11732);
or U11761 (N_11761,N_11667,N_11651);
or U11762 (N_11762,N_11735,N_11660);
xnor U11763 (N_11763,N_11746,N_11721);
nand U11764 (N_11764,N_11726,N_11637);
and U11765 (N_11765,N_11708,N_11718);
and U11766 (N_11766,N_11657,N_11683);
xor U11767 (N_11767,N_11684,N_11672);
xnor U11768 (N_11768,N_11647,N_11671);
nor U11769 (N_11769,N_11644,N_11731);
or U11770 (N_11770,N_11717,N_11669);
and U11771 (N_11771,N_11699,N_11711);
and U11772 (N_11772,N_11714,N_11687);
and U11773 (N_11773,N_11691,N_11658);
or U11774 (N_11774,N_11709,N_11725);
nor U11775 (N_11775,N_11734,N_11713);
nand U11776 (N_11776,N_11686,N_11706);
nand U11777 (N_11777,N_11747,N_11668);
nor U11778 (N_11778,N_11701,N_11674);
or U11779 (N_11779,N_11707,N_11723);
and U11780 (N_11780,N_11736,N_11705);
xor U11781 (N_11781,N_11628,N_11689);
nor U11782 (N_11782,N_11739,N_11666);
and U11783 (N_11783,N_11631,N_11648);
xor U11784 (N_11784,N_11641,N_11742);
or U11785 (N_11785,N_11694,N_11700);
or U11786 (N_11786,N_11670,N_11724);
nor U11787 (N_11787,N_11664,N_11685);
xor U11788 (N_11788,N_11716,N_11710);
nand U11789 (N_11789,N_11638,N_11719);
xnor U11790 (N_11790,N_11720,N_11676);
xnor U11791 (N_11791,N_11629,N_11733);
or U11792 (N_11792,N_11655,N_11649);
xor U11793 (N_11793,N_11695,N_11722);
and U11794 (N_11794,N_11675,N_11650);
or U11795 (N_11795,N_11703,N_11682);
nand U11796 (N_11796,N_11643,N_11673);
nor U11797 (N_11797,N_11659,N_11712);
and U11798 (N_11798,N_11665,N_11727);
nand U11799 (N_11799,N_11625,N_11744);
nor U11800 (N_11800,N_11738,N_11743);
nand U11801 (N_11801,N_11702,N_11748);
nand U11802 (N_11802,N_11661,N_11698);
or U11803 (N_11803,N_11737,N_11696);
nor U11804 (N_11804,N_11642,N_11692);
nor U11805 (N_11805,N_11680,N_11715);
xor U11806 (N_11806,N_11677,N_11633);
and U11807 (N_11807,N_11704,N_11693);
or U11808 (N_11808,N_11730,N_11740);
and U11809 (N_11809,N_11626,N_11662);
nor U11810 (N_11810,N_11690,N_11640);
xnor U11811 (N_11811,N_11652,N_11654);
nor U11812 (N_11812,N_11681,N_11742);
or U11813 (N_11813,N_11668,N_11631);
xor U11814 (N_11814,N_11734,N_11667);
nor U11815 (N_11815,N_11646,N_11700);
and U11816 (N_11816,N_11741,N_11740);
nor U11817 (N_11817,N_11706,N_11731);
and U11818 (N_11818,N_11664,N_11694);
or U11819 (N_11819,N_11724,N_11637);
nand U11820 (N_11820,N_11669,N_11644);
and U11821 (N_11821,N_11627,N_11693);
or U11822 (N_11822,N_11636,N_11663);
nand U11823 (N_11823,N_11667,N_11705);
nand U11824 (N_11824,N_11704,N_11662);
nor U11825 (N_11825,N_11735,N_11666);
nor U11826 (N_11826,N_11634,N_11746);
xnor U11827 (N_11827,N_11680,N_11710);
nand U11828 (N_11828,N_11673,N_11691);
or U11829 (N_11829,N_11713,N_11741);
nand U11830 (N_11830,N_11706,N_11662);
or U11831 (N_11831,N_11639,N_11700);
nor U11832 (N_11832,N_11677,N_11674);
nor U11833 (N_11833,N_11710,N_11749);
nand U11834 (N_11834,N_11698,N_11711);
or U11835 (N_11835,N_11745,N_11681);
nand U11836 (N_11836,N_11713,N_11685);
or U11837 (N_11837,N_11639,N_11696);
nand U11838 (N_11838,N_11723,N_11690);
nand U11839 (N_11839,N_11692,N_11747);
and U11840 (N_11840,N_11738,N_11732);
nand U11841 (N_11841,N_11748,N_11689);
and U11842 (N_11842,N_11634,N_11630);
xnor U11843 (N_11843,N_11661,N_11648);
and U11844 (N_11844,N_11661,N_11681);
and U11845 (N_11845,N_11646,N_11697);
nor U11846 (N_11846,N_11668,N_11731);
xnor U11847 (N_11847,N_11705,N_11645);
nor U11848 (N_11848,N_11687,N_11723);
and U11849 (N_11849,N_11748,N_11652);
and U11850 (N_11850,N_11671,N_11648);
nor U11851 (N_11851,N_11662,N_11728);
nor U11852 (N_11852,N_11689,N_11669);
or U11853 (N_11853,N_11651,N_11629);
nand U11854 (N_11854,N_11684,N_11702);
nand U11855 (N_11855,N_11628,N_11686);
and U11856 (N_11856,N_11639,N_11674);
nand U11857 (N_11857,N_11741,N_11725);
and U11858 (N_11858,N_11678,N_11729);
or U11859 (N_11859,N_11716,N_11742);
nor U11860 (N_11860,N_11680,N_11735);
nand U11861 (N_11861,N_11637,N_11674);
nor U11862 (N_11862,N_11749,N_11670);
xnor U11863 (N_11863,N_11746,N_11663);
nand U11864 (N_11864,N_11680,N_11698);
xor U11865 (N_11865,N_11666,N_11691);
or U11866 (N_11866,N_11639,N_11665);
nor U11867 (N_11867,N_11651,N_11707);
xor U11868 (N_11868,N_11694,N_11711);
nor U11869 (N_11869,N_11682,N_11638);
nor U11870 (N_11870,N_11742,N_11720);
or U11871 (N_11871,N_11697,N_11628);
nor U11872 (N_11872,N_11716,N_11645);
or U11873 (N_11873,N_11660,N_11741);
and U11874 (N_11874,N_11700,N_11687);
xnor U11875 (N_11875,N_11871,N_11821);
xor U11876 (N_11876,N_11798,N_11826);
nor U11877 (N_11877,N_11854,N_11841);
xor U11878 (N_11878,N_11833,N_11786);
nor U11879 (N_11879,N_11779,N_11777);
xnor U11880 (N_11880,N_11814,N_11783);
nand U11881 (N_11881,N_11867,N_11766);
xor U11882 (N_11882,N_11768,N_11767);
and U11883 (N_11883,N_11790,N_11789);
nand U11884 (N_11884,N_11813,N_11788);
and U11885 (N_11885,N_11763,N_11751);
nor U11886 (N_11886,N_11838,N_11858);
xor U11887 (N_11887,N_11754,N_11805);
nor U11888 (N_11888,N_11794,N_11866);
nand U11889 (N_11889,N_11815,N_11809);
nor U11890 (N_11890,N_11761,N_11793);
nand U11891 (N_11891,N_11784,N_11757);
and U11892 (N_11892,N_11837,N_11802);
nor U11893 (N_11893,N_11864,N_11806);
nor U11894 (N_11894,N_11834,N_11831);
and U11895 (N_11895,N_11785,N_11770);
nor U11896 (N_11896,N_11869,N_11778);
and U11897 (N_11897,N_11799,N_11810);
or U11898 (N_11898,N_11753,N_11776);
nor U11899 (N_11899,N_11843,N_11800);
xor U11900 (N_11900,N_11760,N_11860);
or U11901 (N_11901,N_11772,N_11827);
or U11902 (N_11902,N_11872,N_11762);
xor U11903 (N_11903,N_11848,N_11764);
nor U11904 (N_11904,N_11850,N_11835);
and U11905 (N_11905,N_11795,N_11853);
or U11906 (N_11906,N_11865,N_11804);
and U11907 (N_11907,N_11855,N_11874);
xor U11908 (N_11908,N_11829,N_11840);
xnor U11909 (N_11909,N_11812,N_11856);
nand U11910 (N_11910,N_11756,N_11816);
or U11911 (N_11911,N_11750,N_11873);
and U11912 (N_11912,N_11830,N_11797);
and U11913 (N_11913,N_11822,N_11765);
nand U11914 (N_11914,N_11808,N_11823);
nor U11915 (N_11915,N_11839,N_11857);
and U11916 (N_11916,N_11836,N_11819);
and U11917 (N_11917,N_11771,N_11755);
and U11918 (N_11918,N_11774,N_11868);
or U11919 (N_11919,N_11807,N_11775);
or U11920 (N_11920,N_11787,N_11792);
xnor U11921 (N_11921,N_11849,N_11842);
nor U11922 (N_11922,N_11811,N_11828);
nand U11923 (N_11923,N_11759,N_11803);
or U11924 (N_11924,N_11870,N_11758);
or U11925 (N_11925,N_11752,N_11844);
xnor U11926 (N_11926,N_11769,N_11832);
and U11927 (N_11927,N_11773,N_11851);
nor U11928 (N_11928,N_11825,N_11781);
xor U11929 (N_11929,N_11859,N_11862);
xnor U11930 (N_11930,N_11852,N_11820);
nor U11931 (N_11931,N_11863,N_11782);
nor U11932 (N_11932,N_11861,N_11817);
nand U11933 (N_11933,N_11791,N_11796);
or U11934 (N_11934,N_11818,N_11824);
or U11935 (N_11935,N_11801,N_11847);
nand U11936 (N_11936,N_11780,N_11845);
and U11937 (N_11937,N_11846,N_11767);
nor U11938 (N_11938,N_11828,N_11822);
or U11939 (N_11939,N_11799,N_11866);
nand U11940 (N_11940,N_11822,N_11836);
and U11941 (N_11941,N_11817,N_11816);
or U11942 (N_11942,N_11789,N_11785);
xnor U11943 (N_11943,N_11786,N_11764);
nand U11944 (N_11944,N_11849,N_11797);
nor U11945 (N_11945,N_11848,N_11834);
nor U11946 (N_11946,N_11791,N_11784);
and U11947 (N_11947,N_11766,N_11758);
or U11948 (N_11948,N_11812,N_11852);
and U11949 (N_11949,N_11785,N_11781);
nor U11950 (N_11950,N_11831,N_11783);
or U11951 (N_11951,N_11852,N_11825);
nand U11952 (N_11952,N_11786,N_11795);
or U11953 (N_11953,N_11854,N_11861);
nor U11954 (N_11954,N_11818,N_11807);
xnor U11955 (N_11955,N_11841,N_11853);
or U11956 (N_11956,N_11800,N_11791);
nor U11957 (N_11957,N_11781,N_11832);
or U11958 (N_11958,N_11846,N_11790);
xor U11959 (N_11959,N_11791,N_11764);
and U11960 (N_11960,N_11813,N_11823);
or U11961 (N_11961,N_11827,N_11782);
nor U11962 (N_11962,N_11793,N_11757);
nand U11963 (N_11963,N_11755,N_11866);
xnor U11964 (N_11964,N_11797,N_11811);
and U11965 (N_11965,N_11818,N_11783);
xor U11966 (N_11966,N_11762,N_11801);
nand U11967 (N_11967,N_11768,N_11828);
nand U11968 (N_11968,N_11826,N_11762);
xor U11969 (N_11969,N_11809,N_11796);
xnor U11970 (N_11970,N_11803,N_11771);
and U11971 (N_11971,N_11798,N_11774);
nand U11972 (N_11972,N_11860,N_11818);
or U11973 (N_11973,N_11855,N_11781);
or U11974 (N_11974,N_11825,N_11836);
nand U11975 (N_11975,N_11840,N_11838);
or U11976 (N_11976,N_11796,N_11841);
and U11977 (N_11977,N_11783,N_11872);
nor U11978 (N_11978,N_11762,N_11818);
nor U11979 (N_11979,N_11786,N_11867);
and U11980 (N_11980,N_11834,N_11855);
xor U11981 (N_11981,N_11819,N_11861);
and U11982 (N_11982,N_11868,N_11815);
and U11983 (N_11983,N_11813,N_11822);
xnor U11984 (N_11984,N_11798,N_11794);
or U11985 (N_11985,N_11770,N_11861);
nor U11986 (N_11986,N_11860,N_11820);
xor U11987 (N_11987,N_11812,N_11805);
nor U11988 (N_11988,N_11771,N_11853);
xnor U11989 (N_11989,N_11834,N_11782);
and U11990 (N_11990,N_11830,N_11872);
xor U11991 (N_11991,N_11775,N_11857);
or U11992 (N_11992,N_11774,N_11787);
or U11993 (N_11993,N_11785,N_11851);
nor U11994 (N_11994,N_11783,N_11851);
xor U11995 (N_11995,N_11854,N_11848);
and U11996 (N_11996,N_11780,N_11828);
and U11997 (N_11997,N_11862,N_11834);
and U11998 (N_11998,N_11800,N_11834);
nor U11999 (N_11999,N_11842,N_11871);
and U12000 (N_12000,N_11932,N_11954);
nor U12001 (N_12001,N_11925,N_11942);
nor U12002 (N_12002,N_11916,N_11980);
xor U12003 (N_12003,N_11898,N_11981);
nor U12004 (N_12004,N_11928,N_11974);
xnor U12005 (N_12005,N_11924,N_11904);
nand U12006 (N_12006,N_11902,N_11947);
or U12007 (N_12007,N_11931,N_11906);
xor U12008 (N_12008,N_11956,N_11926);
and U12009 (N_12009,N_11953,N_11948);
xnor U12010 (N_12010,N_11900,N_11959);
and U12011 (N_12011,N_11934,N_11939);
nor U12012 (N_12012,N_11937,N_11991);
and U12013 (N_12013,N_11901,N_11969);
nor U12014 (N_12014,N_11976,N_11889);
nor U12015 (N_12015,N_11892,N_11971);
nand U12016 (N_12016,N_11879,N_11883);
nand U12017 (N_12017,N_11943,N_11905);
nor U12018 (N_12018,N_11949,N_11933);
nor U12019 (N_12019,N_11982,N_11922);
nor U12020 (N_12020,N_11990,N_11945);
or U12021 (N_12021,N_11977,N_11996);
xor U12022 (N_12022,N_11936,N_11941);
and U12023 (N_12023,N_11970,N_11944);
or U12024 (N_12024,N_11997,N_11911);
nor U12025 (N_12025,N_11918,N_11927);
nand U12026 (N_12026,N_11952,N_11972);
nand U12027 (N_12027,N_11890,N_11940);
or U12028 (N_12028,N_11897,N_11903);
xor U12029 (N_12029,N_11921,N_11908);
xor U12030 (N_12030,N_11929,N_11966);
nor U12031 (N_12031,N_11995,N_11876);
and U12032 (N_12032,N_11877,N_11896);
nand U12033 (N_12033,N_11957,N_11887);
or U12034 (N_12034,N_11998,N_11888);
nor U12035 (N_12035,N_11962,N_11960);
nand U12036 (N_12036,N_11992,N_11919);
nand U12037 (N_12037,N_11978,N_11993);
nor U12038 (N_12038,N_11994,N_11913);
xnor U12039 (N_12039,N_11891,N_11907);
nand U12040 (N_12040,N_11975,N_11881);
or U12041 (N_12041,N_11984,N_11899);
and U12042 (N_12042,N_11882,N_11958);
or U12043 (N_12043,N_11964,N_11923);
xnor U12044 (N_12044,N_11986,N_11895);
nand U12045 (N_12045,N_11950,N_11987);
xnor U12046 (N_12046,N_11938,N_11917);
nor U12047 (N_12047,N_11909,N_11912);
and U12048 (N_12048,N_11884,N_11985);
and U12049 (N_12049,N_11983,N_11920);
or U12050 (N_12050,N_11989,N_11880);
and U12051 (N_12051,N_11914,N_11935);
and U12052 (N_12052,N_11946,N_11955);
or U12053 (N_12053,N_11885,N_11875);
nand U12054 (N_12054,N_11951,N_11894);
xnor U12055 (N_12055,N_11893,N_11965);
nand U12056 (N_12056,N_11988,N_11961);
or U12057 (N_12057,N_11910,N_11967);
nor U12058 (N_12058,N_11878,N_11915);
nand U12059 (N_12059,N_11886,N_11963);
xor U12060 (N_12060,N_11999,N_11930);
nor U12061 (N_12061,N_11973,N_11968);
and U12062 (N_12062,N_11979,N_11982);
xnor U12063 (N_12063,N_11942,N_11995);
nand U12064 (N_12064,N_11990,N_11966);
or U12065 (N_12065,N_11982,N_11923);
nand U12066 (N_12066,N_11910,N_11939);
or U12067 (N_12067,N_11903,N_11936);
xor U12068 (N_12068,N_11991,N_11896);
xnor U12069 (N_12069,N_11965,N_11908);
nor U12070 (N_12070,N_11977,N_11885);
nor U12071 (N_12071,N_11879,N_11960);
nor U12072 (N_12072,N_11993,N_11917);
nor U12073 (N_12073,N_11922,N_11976);
nor U12074 (N_12074,N_11938,N_11935);
or U12075 (N_12075,N_11978,N_11916);
and U12076 (N_12076,N_11932,N_11959);
or U12077 (N_12077,N_11989,N_11918);
or U12078 (N_12078,N_11958,N_11889);
nand U12079 (N_12079,N_11966,N_11989);
nand U12080 (N_12080,N_11978,N_11939);
or U12081 (N_12081,N_11959,N_11998);
nand U12082 (N_12082,N_11876,N_11880);
or U12083 (N_12083,N_11967,N_11879);
and U12084 (N_12084,N_11885,N_11876);
or U12085 (N_12085,N_11973,N_11992);
or U12086 (N_12086,N_11962,N_11983);
nor U12087 (N_12087,N_11919,N_11980);
nor U12088 (N_12088,N_11991,N_11950);
xor U12089 (N_12089,N_11929,N_11971);
nand U12090 (N_12090,N_11886,N_11877);
and U12091 (N_12091,N_11928,N_11968);
nand U12092 (N_12092,N_11925,N_11905);
or U12093 (N_12093,N_11892,N_11888);
and U12094 (N_12094,N_11920,N_11906);
xor U12095 (N_12095,N_11939,N_11901);
nor U12096 (N_12096,N_11878,N_11949);
nor U12097 (N_12097,N_11963,N_11939);
nand U12098 (N_12098,N_11945,N_11969);
nor U12099 (N_12099,N_11907,N_11951);
xnor U12100 (N_12100,N_11911,N_11954);
xnor U12101 (N_12101,N_11969,N_11924);
and U12102 (N_12102,N_11979,N_11907);
or U12103 (N_12103,N_11961,N_11915);
nand U12104 (N_12104,N_11959,N_11969);
xnor U12105 (N_12105,N_11976,N_11930);
and U12106 (N_12106,N_11923,N_11901);
nand U12107 (N_12107,N_11965,N_11939);
and U12108 (N_12108,N_11987,N_11995);
xor U12109 (N_12109,N_11991,N_11997);
nand U12110 (N_12110,N_11947,N_11944);
nor U12111 (N_12111,N_11938,N_11937);
xnor U12112 (N_12112,N_11955,N_11968);
and U12113 (N_12113,N_11947,N_11985);
nor U12114 (N_12114,N_11928,N_11960);
and U12115 (N_12115,N_11893,N_11980);
nand U12116 (N_12116,N_11997,N_11887);
and U12117 (N_12117,N_11967,N_11970);
nor U12118 (N_12118,N_11881,N_11949);
and U12119 (N_12119,N_11957,N_11962);
and U12120 (N_12120,N_11937,N_11953);
nor U12121 (N_12121,N_11985,N_11937);
and U12122 (N_12122,N_11930,N_11879);
nand U12123 (N_12123,N_11931,N_11881);
nand U12124 (N_12124,N_11979,N_11965);
xor U12125 (N_12125,N_12026,N_12100);
or U12126 (N_12126,N_12068,N_12018);
and U12127 (N_12127,N_12085,N_12077);
or U12128 (N_12128,N_12078,N_12053);
and U12129 (N_12129,N_12108,N_12020);
or U12130 (N_12130,N_12001,N_12107);
nor U12131 (N_12131,N_12052,N_12110);
nand U12132 (N_12132,N_12064,N_12013);
and U12133 (N_12133,N_12010,N_12096);
and U12134 (N_12134,N_12039,N_12051);
and U12135 (N_12135,N_12065,N_12028);
nor U12136 (N_12136,N_12092,N_12056);
nor U12137 (N_12137,N_12022,N_12043);
and U12138 (N_12138,N_12087,N_12115);
or U12139 (N_12139,N_12093,N_12038);
or U12140 (N_12140,N_12113,N_12008);
nor U12141 (N_12141,N_12016,N_12049);
or U12142 (N_12142,N_12099,N_12111);
and U12143 (N_12143,N_12014,N_12048);
nand U12144 (N_12144,N_12116,N_12103);
and U12145 (N_12145,N_12009,N_12063);
nor U12146 (N_12146,N_12044,N_12032);
xnor U12147 (N_12147,N_12124,N_12122);
xnor U12148 (N_12148,N_12035,N_12054);
nor U12149 (N_12149,N_12019,N_12101);
and U12150 (N_12150,N_12011,N_12088);
and U12151 (N_12151,N_12086,N_12042);
nor U12152 (N_12152,N_12118,N_12102);
nor U12153 (N_12153,N_12034,N_12012);
and U12154 (N_12154,N_12059,N_12120);
and U12155 (N_12155,N_12031,N_12098);
nor U12156 (N_12156,N_12074,N_12003);
or U12157 (N_12157,N_12066,N_12123);
nor U12158 (N_12158,N_12062,N_12069);
xor U12159 (N_12159,N_12109,N_12070);
or U12160 (N_12160,N_12040,N_12072);
nor U12161 (N_12161,N_12095,N_12119);
and U12162 (N_12162,N_12117,N_12084);
nor U12163 (N_12163,N_12015,N_12017);
xnor U12164 (N_12164,N_12082,N_12081);
and U12165 (N_12165,N_12036,N_12041);
nor U12166 (N_12166,N_12047,N_12079);
nor U12167 (N_12167,N_12024,N_12005);
nor U12168 (N_12168,N_12097,N_12021);
or U12169 (N_12169,N_12073,N_12106);
nand U12170 (N_12170,N_12000,N_12027);
nand U12171 (N_12171,N_12004,N_12002);
xnor U12172 (N_12172,N_12037,N_12058);
nand U12173 (N_12173,N_12030,N_12091);
and U12174 (N_12174,N_12046,N_12050);
or U12175 (N_12175,N_12083,N_12076);
nor U12176 (N_12176,N_12007,N_12075);
and U12177 (N_12177,N_12090,N_12071);
and U12178 (N_12178,N_12105,N_12029);
nand U12179 (N_12179,N_12104,N_12061);
xor U12180 (N_12180,N_12080,N_12112);
or U12181 (N_12181,N_12045,N_12025);
or U12182 (N_12182,N_12114,N_12055);
and U12183 (N_12183,N_12089,N_12067);
xor U12184 (N_12184,N_12094,N_12060);
or U12185 (N_12185,N_12033,N_12006);
nor U12186 (N_12186,N_12057,N_12023);
nor U12187 (N_12187,N_12121,N_12080);
and U12188 (N_12188,N_12031,N_12101);
nor U12189 (N_12189,N_12086,N_12049);
and U12190 (N_12190,N_12015,N_12091);
xor U12191 (N_12191,N_12078,N_12074);
xnor U12192 (N_12192,N_12065,N_12085);
and U12193 (N_12193,N_12029,N_12061);
nor U12194 (N_12194,N_12029,N_12071);
xor U12195 (N_12195,N_12004,N_12000);
and U12196 (N_12196,N_12070,N_12087);
or U12197 (N_12197,N_12000,N_12048);
nand U12198 (N_12198,N_12011,N_12092);
xnor U12199 (N_12199,N_12114,N_12030);
xor U12200 (N_12200,N_12043,N_12102);
xnor U12201 (N_12201,N_12086,N_12053);
xor U12202 (N_12202,N_12086,N_12037);
and U12203 (N_12203,N_12029,N_12056);
xor U12204 (N_12204,N_12119,N_12077);
and U12205 (N_12205,N_12048,N_12099);
and U12206 (N_12206,N_12057,N_12051);
nor U12207 (N_12207,N_12073,N_12031);
and U12208 (N_12208,N_12090,N_12037);
nor U12209 (N_12209,N_12016,N_12098);
xnor U12210 (N_12210,N_12070,N_12004);
and U12211 (N_12211,N_12070,N_12104);
nand U12212 (N_12212,N_12069,N_12113);
nand U12213 (N_12213,N_12094,N_12077);
nand U12214 (N_12214,N_12070,N_12115);
nand U12215 (N_12215,N_12078,N_12083);
xnor U12216 (N_12216,N_12040,N_12059);
and U12217 (N_12217,N_12071,N_12016);
nor U12218 (N_12218,N_12124,N_12111);
nor U12219 (N_12219,N_12115,N_12077);
and U12220 (N_12220,N_12120,N_12122);
or U12221 (N_12221,N_12056,N_12118);
xnor U12222 (N_12222,N_12018,N_12092);
or U12223 (N_12223,N_12072,N_12003);
and U12224 (N_12224,N_12110,N_12081);
or U12225 (N_12225,N_12005,N_12066);
or U12226 (N_12226,N_12027,N_12084);
nor U12227 (N_12227,N_12107,N_12096);
nand U12228 (N_12228,N_12012,N_12101);
nand U12229 (N_12229,N_12010,N_12041);
nor U12230 (N_12230,N_12015,N_12106);
nor U12231 (N_12231,N_12017,N_12072);
and U12232 (N_12232,N_12034,N_12093);
or U12233 (N_12233,N_12078,N_12105);
nand U12234 (N_12234,N_12112,N_12113);
or U12235 (N_12235,N_12039,N_12100);
and U12236 (N_12236,N_12049,N_12087);
xor U12237 (N_12237,N_12103,N_12083);
xnor U12238 (N_12238,N_12090,N_12021);
or U12239 (N_12239,N_12094,N_12089);
or U12240 (N_12240,N_12066,N_12020);
nor U12241 (N_12241,N_12114,N_12057);
or U12242 (N_12242,N_12003,N_12076);
and U12243 (N_12243,N_12030,N_12069);
and U12244 (N_12244,N_12018,N_12121);
or U12245 (N_12245,N_12038,N_12019);
nand U12246 (N_12246,N_12117,N_12088);
or U12247 (N_12247,N_12053,N_12019);
nor U12248 (N_12248,N_12046,N_12059);
xor U12249 (N_12249,N_12004,N_12071);
nand U12250 (N_12250,N_12136,N_12132);
xnor U12251 (N_12251,N_12181,N_12158);
nor U12252 (N_12252,N_12131,N_12151);
or U12253 (N_12253,N_12230,N_12229);
nor U12254 (N_12254,N_12233,N_12139);
nor U12255 (N_12255,N_12169,N_12193);
xnor U12256 (N_12256,N_12221,N_12202);
nor U12257 (N_12257,N_12200,N_12172);
nor U12258 (N_12258,N_12219,N_12125);
or U12259 (N_12259,N_12183,N_12141);
or U12260 (N_12260,N_12225,N_12189);
or U12261 (N_12261,N_12184,N_12239);
nor U12262 (N_12262,N_12155,N_12236);
and U12263 (N_12263,N_12185,N_12199);
nor U12264 (N_12264,N_12153,N_12174);
xnor U12265 (N_12265,N_12223,N_12217);
nand U12266 (N_12266,N_12138,N_12232);
or U12267 (N_12267,N_12152,N_12150);
or U12268 (N_12268,N_12245,N_12156);
or U12269 (N_12269,N_12216,N_12247);
nand U12270 (N_12270,N_12201,N_12192);
nand U12271 (N_12271,N_12171,N_12210);
or U12272 (N_12272,N_12145,N_12215);
nor U12273 (N_12273,N_12128,N_12126);
nand U12274 (N_12274,N_12157,N_12227);
and U12275 (N_12275,N_12231,N_12163);
nand U12276 (N_12276,N_12162,N_12160);
or U12277 (N_12277,N_12147,N_12148);
and U12278 (N_12278,N_12188,N_12246);
nand U12279 (N_12279,N_12127,N_12165);
xnor U12280 (N_12280,N_12242,N_12205);
xnor U12281 (N_12281,N_12191,N_12212);
or U12282 (N_12282,N_12173,N_12222);
nor U12283 (N_12283,N_12167,N_12226);
or U12284 (N_12284,N_12179,N_12135);
or U12285 (N_12285,N_12238,N_12234);
nor U12286 (N_12286,N_12220,N_12144);
and U12287 (N_12287,N_12146,N_12224);
xor U12288 (N_12288,N_12243,N_12206);
nand U12289 (N_12289,N_12197,N_12248);
xor U12290 (N_12290,N_12161,N_12213);
nor U12291 (N_12291,N_12159,N_12196);
nand U12292 (N_12292,N_12244,N_12175);
and U12293 (N_12293,N_12208,N_12235);
xor U12294 (N_12294,N_12140,N_12198);
or U12295 (N_12295,N_12207,N_12170);
or U12296 (N_12296,N_12130,N_12129);
and U12297 (N_12297,N_12190,N_12149);
xor U12298 (N_12298,N_12180,N_12168);
or U12299 (N_12299,N_12178,N_12182);
nor U12300 (N_12300,N_12187,N_12237);
xor U12301 (N_12301,N_12186,N_12228);
or U12302 (N_12302,N_12194,N_12240);
and U12303 (N_12303,N_12209,N_12177);
nand U12304 (N_12304,N_12203,N_12164);
xnor U12305 (N_12305,N_12137,N_12176);
or U12306 (N_12306,N_12241,N_12154);
and U12307 (N_12307,N_12142,N_12211);
xnor U12308 (N_12308,N_12143,N_12166);
nor U12309 (N_12309,N_12218,N_12204);
nor U12310 (N_12310,N_12195,N_12249);
and U12311 (N_12311,N_12214,N_12134);
nor U12312 (N_12312,N_12133,N_12233);
xor U12313 (N_12313,N_12199,N_12221);
or U12314 (N_12314,N_12173,N_12181);
or U12315 (N_12315,N_12180,N_12245);
and U12316 (N_12316,N_12240,N_12130);
nor U12317 (N_12317,N_12131,N_12180);
xor U12318 (N_12318,N_12127,N_12188);
nand U12319 (N_12319,N_12183,N_12166);
nor U12320 (N_12320,N_12152,N_12166);
nand U12321 (N_12321,N_12156,N_12147);
and U12322 (N_12322,N_12181,N_12127);
and U12323 (N_12323,N_12156,N_12186);
and U12324 (N_12324,N_12160,N_12191);
and U12325 (N_12325,N_12151,N_12142);
nor U12326 (N_12326,N_12179,N_12128);
xnor U12327 (N_12327,N_12173,N_12175);
nand U12328 (N_12328,N_12151,N_12146);
xnor U12329 (N_12329,N_12198,N_12163);
and U12330 (N_12330,N_12146,N_12179);
and U12331 (N_12331,N_12130,N_12150);
xor U12332 (N_12332,N_12153,N_12175);
xor U12333 (N_12333,N_12145,N_12139);
xor U12334 (N_12334,N_12167,N_12213);
or U12335 (N_12335,N_12172,N_12134);
xnor U12336 (N_12336,N_12136,N_12184);
nand U12337 (N_12337,N_12163,N_12174);
and U12338 (N_12338,N_12211,N_12187);
and U12339 (N_12339,N_12195,N_12234);
or U12340 (N_12340,N_12243,N_12234);
nor U12341 (N_12341,N_12192,N_12170);
nand U12342 (N_12342,N_12128,N_12215);
nor U12343 (N_12343,N_12209,N_12145);
xnor U12344 (N_12344,N_12143,N_12171);
nand U12345 (N_12345,N_12231,N_12190);
nor U12346 (N_12346,N_12229,N_12243);
xor U12347 (N_12347,N_12137,N_12151);
nor U12348 (N_12348,N_12220,N_12194);
xnor U12349 (N_12349,N_12202,N_12249);
nand U12350 (N_12350,N_12144,N_12244);
nand U12351 (N_12351,N_12231,N_12189);
or U12352 (N_12352,N_12228,N_12180);
or U12353 (N_12353,N_12141,N_12148);
xnor U12354 (N_12354,N_12146,N_12147);
or U12355 (N_12355,N_12240,N_12134);
nand U12356 (N_12356,N_12158,N_12204);
or U12357 (N_12357,N_12221,N_12180);
nand U12358 (N_12358,N_12223,N_12155);
xor U12359 (N_12359,N_12192,N_12156);
or U12360 (N_12360,N_12151,N_12206);
nand U12361 (N_12361,N_12222,N_12164);
nor U12362 (N_12362,N_12206,N_12135);
nand U12363 (N_12363,N_12187,N_12244);
or U12364 (N_12364,N_12221,N_12223);
nand U12365 (N_12365,N_12208,N_12142);
nand U12366 (N_12366,N_12146,N_12155);
xor U12367 (N_12367,N_12241,N_12216);
nor U12368 (N_12368,N_12215,N_12162);
or U12369 (N_12369,N_12136,N_12200);
xor U12370 (N_12370,N_12239,N_12203);
and U12371 (N_12371,N_12183,N_12227);
nand U12372 (N_12372,N_12241,N_12186);
or U12373 (N_12373,N_12217,N_12140);
nand U12374 (N_12374,N_12191,N_12143);
and U12375 (N_12375,N_12304,N_12337);
or U12376 (N_12376,N_12299,N_12352);
nor U12377 (N_12377,N_12322,N_12300);
or U12378 (N_12378,N_12265,N_12266);
and U12379 (N_12379,N_12267,N_12336);
and U12380 (N_12380,N_12294,N_12344);
or U12381 (N_12381,N_12280,N_12252);
and U12382 (N_12382,N_12319,N_12297);
xnor U12383 (N_12383,N_12274,N_12264);
xnor U12384 (N_12384,N_12276,N_12330);
nand U12385 (N_12385,N_12310,N_12347);
or U12386 (N_12386,N_12369,N_12317);
xor U12387 (N_12387,N_12298,N_12285);
and U12388 (N_12388,N_12279,N_12313);
xor U12389 (N_12389,N_12342,N_12254);
and U12390 (N_12390,N_12366,N_12282);
nor U12391 (N_12391,N_12348,N_12340);
nor U12392 (N_12392,N_12373,N_12309);
nor U12393 (N_12393,N_12316,N_12302);
nand U12394 (N_12394,N_12372,N_12341);
or U12395 (N_12395,N_12359,N_12353);
nor U12396 (N_12396,N_12354,N_12329);
nor U12397 (N_12397,N_12332,N_12368);
xor U12398 (N_12398,N_12286,N_12306);
or U12399 (N_12399,N_12360,N_12289);
xor U12400 (N_12400,N_12335,N_12260);
xor U12401 (N_12401,N_12278,N_12327);
nor U12402 (N_12402,N_12281,N_12345);
and U12403 (N_12403,N_12361,N_12270);
nor U12404 (N_12404,N_12258,N_12269);
xor U12405 (N_12405,N_12271,N_12307);
nand U12406 (N_12406,N_12293,N_12301);
and U12407 (N_12407,N_12362,N_12350);
nand U12408 (N_12408,N_12349,N_12296);
and U12409 (N_12409,N_12261,N_12331);
xnor U12410 (N_12410,N_12275,N_12268);
xor U12411 (N_12411,N_12305,N_12262);
nand U12412 (N_12412,N_12338,N_12283);
nand U12413 (N_12413,N_12277,N_12290);
xor U12414 (N_12414,N_12311,N_12291);
and U12415 (N_12415,N_12326,N_12351);
or U12416 (N_12416,N_12363,N_12323);
nor U12417 (N_12417,N_12343,N_12284);
and U12418 (N_12418,N_12355,N_12255);
nor U12419 (N_12419,N_12315,N_12288);
and U12420 (N_12420,N_12250,N_12259);
nand U12421 (N_12421,N_12320,N_12324);
nor U12422 (N_12422,N_12263,N_12321);
and U12423 (N_12423,N_12339,N_12334);
or U12424 (N_12424,N_12325,N_12333);
and U12425 (N_12425,N_12314,N_12346);
xor U12426 (N_12426,N_12371,N_12374);
xor U12427 (N_12427,N_12272,N_12287);
nand U12428 (N_12428,N_12357,N_12367);
nor U12429 (N_12429,N_12257,N_12370);
or U12430 (N_12430,N_12251,N_12292);
nand U12431 (N_12431,N_12273,N_12253);
nand U12432 (N_12432,N_12358,N_12356);
nor U12433 (N_12433,N_12295,N_12256);
xnor U12434 (N_12434,N_12312,N_12328);
nor U12435 (N_12435,N_12308,N_12364);
and U12436 (N_12436,N_12365,N_12318);
nor U12437 (N_12437,N_12303,N_12315);
and U12438 (N_12438,N_12358,N_12279);
xor U12439 (N_12439,N_12341,N_12292);
or U12440 (N_12440,N_12253,N_12325);
xor U12441 (N_12441,N_12370,N_12367);
nand U12442 (N_12442,N_12364,N_12312);
and U12443 (N_12443,N_12292,N_12327);
xnor U12444 (N_12444,N_12305,N_12288);
or U12445 (N_12445,N_12335,N_12255);
xor U12446 (N_12446,N_12361,N_12370);
nor U12447 (N_12447,N_12272,N_12321);
nand U12448 (N_12448,N_12332,N_12281);
nor U12449 (N_12449,N_12335,N_12308);
and U12450 (N_12450,N_12268,N_12277);
and U12451 (N_12451,N_12335,N_12320);
nor U12452 (N_12452,N_12271,N_12315);
or U12453 (N_12453,N_12281,N_12272);
and U12454 (N_12454,N_12319,N_12353);
xor U12455 (N_12455,N_12301,N_12296);
nor U12456 (N_12456,N_12358,N_12265);
nand U12457 (N_12457,N_12274,N_12298);
xnor U12458 (N_12458,N_12263,N_12293);
and U12459 (N_12459,N_12291,N_12350);
and U12460 (N_12460,N_12275,N_12308);
xnor U12461 (N_12461,N_12261,N_12328);
xor U12462 (N_12462,N_12295,N_12372);
xnor U12463 (N_12463,N_12357,N_12296);
or U12464 (N_12464,N_12319,N_12312);
nor U12465 (N_12465,N_12368,N_12347);
nor U12466 (N_12466,N_12250,N_12272);
nor U12467 (N_12467,N_12345,N_12356);
or U12468 (N_12468,N_12343,N_12277);
and U12469 (N_12469,N_12270,N_12351);
or U12470 (N_12470,N_12368,N_12275);
nand U12471 (N_12471,N_12262,N_12286);
nand U12472 (N_12472,N_12350,N_12329);
and U12473 (N_12473,N_12331,N_12355);
nand U12474 (N_12474,N_12256,N_12359);
nand U12475 (N_12475,N_12307,N_12360);
nand U12476 (N_12476,N_12267,N_12284);
and U12477 (N_12477,N_12356,N_12329);
nor U12478 (N_12478,N_12350,N_12317);
xnor U12479 (N_12479,N_12333,N_12364);
xnor U12480 (N_12480,N_12328,N_12342);
and U12481 (N_12481,N_12335,N_12359);
xnor U12482 (N_12482,N_12252,N_12277);
nand U12483 (N_12483,N_12290,N_12287);
xor U12484 (N_12484,N_12314,N_12358);
or U12485 (N_12485,N_12346,N_12365);
nand U12486 (N_12486,N_12318,N_12348);
or U12487 (N_12487,N_12276,N_12360);
nand U12488 (N_12488,N_12328,N_12272);
nand U12489 (N_12489,N_12333,N_12302);
xnor U12490 (N_12490,N_12317,N_12261);
or U12491 (N_12491,N_12282,N_12364);
nand U12492 (N_12492,N_12311,N_12318);
nand U12493 (N_12493,N_12328,N_12265);
xor U12494 (N_12494,N_12290,N_12352);
and U12495 (N_12495,N_12354,N_12357);
xnor U12496 (N_12496,N_12360,N_12353);
nor U12497 (N_12497,N_12280,N_12267);
or U12498 (N_12498,N_12347,N_12360);
or U12499 (N_12499,N_12312,N_12292);
or U12500 (N_12500,N_12434,N_12451);
nor U12501 (N_12501,N_12414,N_12444);
and U12502 (N_12502,N_12481,N_12454);
nor U12503 (N_12503,N_12499,N_12453);
nor U12504 (N_12504,N_12383,N_12376);
nand U12505 (N_12505,N_12385,N_12482);
or U12506 (N_12506,N_12472,N_12393);
or U12507 (N_12507,N_12448,N_12440);
nand U12508 (N_12508,N_12400,N_12394);
or U12509 (N_12509,N_12437,N_12431);
nand U12510 (N_12510,N_12496,N_12474);
nand U12511 (N_12511,N_12391,N_12486);
xnor U12512 (N_12512,N_12468,N_12413);
and U12513 (N_12513,N_12462,N_12457);
and U12514 (N_12514,N_12463,N_12450);
nor U12515 (N_12515,N_12443,N_12399);
xnor U12516 (N_12516,N_12497,N_12420);
or U12517 (N_12517,N_12470,N_12447);
or U12518 (N_12518,N_12484,N_12464);
nand U12519 (N_12519,N_12492,N_12421);
xor U12520 (N_12520,N_12422,N_12452);
or U12521 (N_12521,N_12446,N_12433);
nand U12522 (N_12522,N_12483,N_12460);
nor U12523 (N_12523,N_12398,N_12430);
and U12524 (N_12524,N_12378,N_12479);
or U12525 (N_12525,N_12487,N_12485);
nor U12526 (N_12526,N_12428,N_12379);
nor U12527 (N_12527,N_12423,N_12416);
nand U12528 (N_12528,N_12375,N_12494);
xnor U12529 (N_12529,N_12471,N_12384);
nand U12530 (N_12530,N_12445,N_12390);
nand U12531 (N_12531,N_12382,N_12466);
and U12532 (N_12532,N_12476,N_12461);
nor U12533 (N_12533,N_12396,N_12498);
nand U12534 (N_12534,N_12392,N_12402);
or U12535 (N_12535,N_12380,N_12426);
nand U12536 (N_12536,N_12418,N_12465);
nand U12537 (N_12537,N_12432,N_12439);
nand U12538 (N_12538,N_12404,N_12469);
xor U12539 (N_12539,N_12488,N_12408);
nand U12540 (N_12540,N_12417,N_12401);
nand U12541 (N_12541,N_12411,N_12456);
nor U12542 (N_12542,N_12410,N_12475);
and U12543 (N_12543,N_12403,N_12493);
xnor U12544 (N_12544,N_12395,N_12407);
nand U12545 (N_12545,N_12397,N_12389);
xnor U12546 (N_12546,N_12429,N_12377);
or U12547 (N_12547,N_12438,N_12495);
xnor U12548 (N_12548,N_12435,N_12467);
xor U12549 (N_12549,N_12386,N_12406);
and U12550 (N_12550,N_12412,N_12425);
nand U12551 (N_12551,N_12442,N_12458);
and U12552 (N_12552,N_12441,N_12405);
and U12553 (N_12553,N_12427,N_12388);
and U12554 (N_12554,N_12489,N_12477);
or U12555 (N_12555,N_12478,N_12491);
or U12556 (N_12556,N_12436,N_12473);
xor U12557 (N_12557,N_12480,N_12455);
or U12558 (N_12558,N_12419,N_12449);
or U12559 (N_12559,N_12459,N_12424);
nand U12560 (N_12560,N_12409,N_12490);
or U12561 (N_12561,N_12381,N_12387);
nand U12562 (N_12562,N_12415,N_12449);
nor U12563 (N_12563,N_12433,N_12471);
or U12564 (N_12564,N_12378,N_12416);
nor U12565 (N_12565,N_12416,N_12480);
xnor U12566 (N_12566,N_12477,N_12459);
nand U12567 (N_12567,N_12378,N_12412);
or U12568 (N_12568,N_12441,N_12385);
xor U12569 (N_12569,N_12381,N_12444);
nor U12570 (N_12570,N_12405,N_12448);
and U12571 (N_12571,N_12478,N_12476);
or U12572 (N_12572,N_12475,N_12426);
nand U12573 (N_12573,N_12443,N_12450);
or U12574 (N_12574,N_12467,N_12477);
nor U12575 (N_12575,N_12430,N_12387);
or U12576 (N_12576,N_12400,N_12417);
xor U12577 (N_12577,N_12457,N_12474);
and U12578 (N_12578,N_12448,N_12493);
xor U12579 (N_12579,N_12448,N_12390);
xnor U12580 (N_12580,N_12377,N_12477);
or U12581 (N_12581,N_12499,N_12485);
and U12582 (N_12582,N_12465,N_12388);
or U12583 (N_12583,N_12386,N_12473);
or U12584 (N_12584,N_12422,N_12480);
nand U12585 (N_12585,N_12461,N_12429);
and U12586 (N_12586,N_12488,N_12470);
nor U12587 (N_12587,N_12378,N_12462);
and U12588 (N_12588,N_12447,N_12414);
xnor U12589 (N_12589,N_12420,N_12380);
xnor U12590 (N_12590,N_12416,N_12479);
xnor U12591 (N_12591,N_12400,N_12444);
and U12592 (N_12592,N_12400,N_12469);
nand U12593 (N_12593,N_12474,N_12378);
nor U12594 (N_12594,N_12455,N_12479);
xor U12595 (N_12595,N_12406,N_12499);
nand U12596 (N_12596,N_12383,N_12445);
xnor U12597 (N_12597,N_12387,N_12463);
nand U12598 (N_12598,N_12384,N_12487);
nor U12599 (N_12599,N_12383,N_12461);
and U12600 (N_12600,N_12437,N_12482);
xor U12601 (N_12601,N_12423,N_12489);
xnor U12602 (N_12602,N_12457,N_12484);
xnor U12603 (N_12603,N_12468,N_12388);
xnor U12604 (N_12604,N_12384,N_12415);
nor U12605 (N_12605,N_12416,N_12405);
or U12606 (N_12606,N_12453,N_12376);
xor U12607 (N_12607,N_12390,N_12388);
xor U12608 (N_12608,N_12412,N_12473);
nor U12609 (N_12609,N_12418,N_12387);
or U12610 (N_12610,N_12419,N_12385);
and U12611 (N_12611,N_12435,N_12408);
and U12612 (N_12612,N_12480,N_12478);
nand U12613 (N_12613,N_12473,N_12457);
and U12614 (N_12614,N_12467,N_12485);
and U12615 (N_12615,N_12425,N_12467);
and U12616 (N_12616,N_12398,N_12451);
nor U12617 (N_12617,N_12427,N_12397);
nor U12618 (N_12618,N_12421,N_12388);
and U12619 (N_12619,N_12404,N_12390);
nand U12620 (N_12620,N_12477,N_12439);
nand U12621 (N_12621,N_12425,N_12390);
or U12622 (N_12622,N_12478,N_12432);
nor U12623 (N_12623,N_12391,N_12485);
and U12624 (N_12624,N_12430,N_12475);
or U12625 (N_12625,N_12545,N_12530);
xnor U12626 (N_12626,N_12589,N_12568);
or U12627 (N_12627,N_12553,N_12599);
xor U12628 (N_12628,N_12605,N_12604);
nand U12629 (N_12629,N_12531,N_12536);
nand U12630 (N_12630,N_12581,N_12616);
nor U12631 (N_12631,N_12597,N_12576);
and U12632 (N_12632,N_12612,N_12577);
or U12633 (N_12633,N_12611,N_12623);
nand U12634 (N_12634,N_12543,N_12600);
and U12635 (N_12635,N_12617,N_12529);
xor U12636 (N_12636,N_12548,N_12580);
or U12637 (N_12637,N_12556,N_12592);
or U12638 (N_12638,N_12512,N_12614);
xnor U12639 (N_12639,N_12560,N_12542);
or U12640 (N_12640,N_12517,N_12559);
nand U12641 (N_12641,N_12507,N_12624);
or U12642 (N_12642,N_12506,N_12569);
xor U12643 (N_12643,N_12534,N_12567);
nand U12644 (N_12644,N_12603,N_12594);
nand U12645 (N_12645,N_12610,N_12566);
and U12646 (N_12646,N_12535,N_12511);
xnor U12647 (N_12647,N_12582,N_12574);
and U12648 (N_12648,N_12565,N_12601);
nor U12649 (N_12649,N_12527,N_12561);
nand U12650 (N_12650,N_12583,N_12551);
nor U12651 (N_12651,N_12524,N_12570);
and U12652 (N_12652,N_12591,N_12547);
or U12653 (N_12653,N_12578,N_12590);
nor U12654 (N_12654,N_12584,N_12523);
nor U12655 (N_12655,N_12613,N_12595);
xor U12656 (N_12656,N_12525,N_12509);
nand U12657 (N_12657,N_12596,N_12526);
or U12658 (N_12658,N_12518,N_12502);
xnor U12659 (N_12659,N_12501,N_12621);
xnor U12660 (N_12660,N_12540,N_12552);
and U12661 (N_12661,N_12537,N_12615);
and U12662 (N_12662,N_12622,N_12516);
and U12663 (N_12663,N_12562,N_12500);
and U12664 (N_12664,N_12539,N_12522);
or U12665 (N_12665,N_12571,N_12504);
xnor U12666 (N_12666,N_12602,N_12515);
xnor U12667 (N_12667,N_12541,N_12585);
xor U12668 (N_12668,N_12532,N_12521);
xor U12669 (N_12669,N_12549,N_12519);
or U12670 (N_12670,N_12520,N_12563);
or U12671 (N_12671,N_12538,N_12586);
or U12672 (N_12672,N_12588,N_12593);
nand U12673 (N_12673,N_12544,N_12573);
and U12674 (N_12674,N_12608,N_12598);
or U12675 (N_12675,N_12510,N_12546);
or U12676 (N_12676,N_12514,N_12533);
or U12677 (N_12677,N_12607,N_12505);
and U12678 (N_12678,N_12575,N_12606);
nand U12679 (N_12679,N_12508,N_12587);
nand U12680 (N_12680,N_12564,N_12554);
or U12681 (N_12681,N_12513,N_12572);
and U12682 (N_12682,N_12555,N_12619);
nor U12683 (N_12683,N_12620,N_12528);
and U12684 (N_12684,N_12618,N_12579);
nor U12685 (N_12685,N_12558,N_12557);
and U12686 (N_12686,N_12550,N_12609);
or U12687 (N_12687,N_12503,N_12511);
or U12688 (N_12688,N_12524,N_12614);
nor U12689 (N_12689,N_12541,N_12529);
xor U12690 (N_12690,N_12513,N_12535);
xnor U12691 (N_12691,N_12530,N_12544);
xnor U12692 (N_12692,N_12507,N_12580);
nand U12693 (N_12693,N_12535,N_12558);
xnor U12694 (N_12694,N_12535,N_12574);
nor U12695 (N_12695,N_12555,N_12526);
nor U12696 (N_12696,N_12560,N_12528);
nor U12697 (N_12697,N_12535,N_12617);
xnor U12698 (N_12698,N_12540,N_12551);
nor U12699 (N_12699,N_12609,N_12501);
nor U12700 (N_12700,N_12600,N_12538);
or U12701 (N_12701,N_12596,N_12591);
and U12702 (N_12702,N_12597,N_12584);
nand U12703 (N_12703,N_12577,N_12565);
nor U12704 (N_12704,N_12530,N_12523);
nand U12705 (N_12705,N_12555,N_12512);
nor U12706 (N_12706,N_12580,N_12506);
and U12707 (N_12707,N_12574,N_12607);
xor U12708 (N_12708,N_12559,N_12500);
or U12709 (N_12709,N_12614,N_12540);
nor U12710 (N_12710,N_12623,N_12594);
and U12711 (N_12711,N_12575,N_12531);
nor U12712 (N_12712,N_12597,N_12570);
nor U12713 (N_12713,N_12504,N_12565);
and U12714 (N_12714,N_12536,N_12592);
or U12715 (N_12715,N_12562,N_12577);
xor U12716 (N_12716,N_12607,N_12530);
xnor U12717 (N_12717,N_12609,N_12614);
or U12718 (N_12718,N_12615,N_12521);
and U12719 (N_12719,N_12621,N_12554);
nor U12720 (N_12720,N_12509,N_12612);
nand U12721 (N_12721,N_12549,N_12504);
nand U12722 (N_12722,N_12524,N_12536);
nor U12723 (N_12723,N_12591,N_12590);
and U12724 (N_12724,N_12599,N_12596);
or U12725 (N_12725,N_12516,N_12514);
xor U12726 (N_12726,N_12616,N_12513);
xor U12727 (N_12727,N_12527,N_12549);
nand U12728 (N_12728,N_12592,N_12620);
or U12729 (N_12729,N_12606,N_12529);
or U12730 (N_12730,N_12590,N_12586);
nor U12731 (N_12731,N_12542,N_12599);
nand U12732 (N_12732,N_12501,N_12569);
and U12733 (N_12733,N_12612,N_12560);
nor U12734 (N_12734,N_12600,N_12554);
or U12735 (N_12735,N_12541,N_12522);
or U12736 (N_12736,N_12599,N_12514);
nand U12737 (N_12737,N_12598,N_12508);
nor U12738 (N_12738,N_12573,N_12510);
xnor U12739 (N_12739,N_12522,N_12515);
xor U12740 (N_12740,N_12591,N_12553);
xnor U12741 (N_12741,N_12563,N_12568);
nor U12742 (N_12742,N_12546,N_12611);
nand U12743 (N_12743,N_12506,N_12598);
or U12744 (N_12744,N_12512,N_12518);
and U12745 (N_12745,N_12575,N_12553);
nand U12746 (N_12746,N_12613,N_12551);
and U12747 (N_12747,N_12529,N_12539);
nor U12748 (N_12748,N_12618,N_12505);
nor U12749 (N_12749,N_12504,N_12576);
nor U12750 (N_12750,N_12625,N_12686);
and U12751 (N_12751,N_12627,N_12730);
xor U12752 (N_12752,N_12651,N_12720);
xor U12753 (N_12753,N_12644,N_12653);
xnor U12754 (N_12754,N_12682,N_12665);
nor U12755 (N_12755,N_12728,N_12749);
and U12756 (N_12756,N_12664,N_12692);
xnor U12757 (N_12757,N_12643,N_12674);
xor U12758 (N_12758,N_12701,N_12680);
nor U12759 (N_12759,N_12714,N_12628);
nor U12760 (N_12760,N_12655,N_12632);
nor U12761 (N_12761,N_12734,N_12745);
nand U12762 (N_12762,N_12725,N_12671);
or U12763 (N_12763,N_12709,N_12735);
xor U12764 (N_12764,N_12744,N_12656);
and U12765 (N_12765,N_12710,N_12652);
and U12766 (N_12766,N_12742,N_12642);
nand U12767 (N_12767,N_12741,N_12715);
and U12768 (N_12768,N_12663,N_12667);
or U12769 (N_12769,N_12717,N_12669);
nor U12770 (N_12770,N_12637,N_12641);
nand U12771 (N_12771,N_12683,N_12647);
nor U12772 (N_12772,N_12704,N_12678);
xor U12773 (N_12773,N_12706,N_12689);
xnor U12774 (N_12774,N_12646,N_12662);
xnor U12775 (N_12775,N_12740,N_12743);
or U12776 (N_12776,N_12713,N_12703);
nand U12777 (N_12777,N_12732,N_12638);
nor U12778 (N_12778,N_12648,N_12723);
xnor U12779 (N_12779,N_12731,N_12666);
nor U12780 (N_12780,N_12748,N_12718);
nand U12781 (N_12781,N_12721,N_12654);
nor U12782 (N_12782,N_12729,N_12629);
nand U12783 (N_12783,N_12691,N_12700);
and U12784 (N_12784,N_12675,N_12633);
or U12785 (N_12785,N_12702,N_12712);
xor U12786 (N_12786,N_12645,N_12636);
xor U12787 (N_12787,N_12626,N_12673);
nor U12788 (N_12788,N_12736,N_12681);
and U12789 (N_12789,N_12737,N_12658);
nor U12790 (N_12790,N_12676,N_12650);
or U12791 (N_12791,N_12733,N_12746);
and U12792 (N_12792,N_12698,N_12685);
xor U12793 (N_12793,N_12738,N_12659);
or U12794 (N_12794,N_12631,N_12679);
and U12795 (N_12795,N_12639,N_12649);
and U12796 (N_12796,N_12634,N_12640);
and U12797 (N_12797,N_12747,N_12668);
xor U12798 (N_12798,N_12697,N_12716);
nor U12799 (N_12799,N_12687,N_12707);
nand U12800 (N_12800,N_12661,N_12724);
or U12801 (N_12801,N_12699,N_12696);
or U12802 (N_12802,N_12690,N_12670);
and U12803 (N_12803,N_12677,N_12672);
nand U12804 (N_12804,N_12708,N_12711);
xor U12805 (N_12805,N_12719,N_12705);
or U12806 (N_12806,N_12657,N_12727);
and U12807 (N_12807,N_12635,N_12630);
nor U12808 (N_12808,N_12684,N_12739);
nor U12809 (N_12809,N_12722,N_12660);
and U12810 (N_12810,N_12688,N_12726);
and U12811 (N_12811,N_12693,N_12694);
or U12812 (N_12812,N_12695,N_12668);
or U12813 (N_12813,N_12668,N_12669);
and U12814 (N_12814,N_12690,N_12742);
xnor U12815 (N_12815,N_12650,N_12696);
xor U12816 (N_12816,N_12671,N_12748);
xnor U12817 (N_12817,N_12730,N_12711);
or U12818 (N_12818,N_12722,N_12652);
nor U12819 (N_12819,N_12735,N_12640);
nor U12820 (N_12820,N_12703,N_12633);
xor U12821 (N_12821,N_12671,N_12687);
xnor U12822 (N_12822,N_12720,N_12661);
or U12823 (N_12823,N_12740,N_12685);
nand U12824 (N_12824,N_12671,N_12626);
or U12825 (N_12825,N_12740,N_12625);
xor U12826 (N_12826,N_12632,N_12727);
or U12827 (N_12827,N_12670,N_12731);
xnor U12828 (N_12828,N_12745,N_12704);
xnor U12829 (N_12829,N_12717,N_12734);
and U12830 (N_12830,N_12644,N_12713);
xnor U12831 (N_12831,N_12648,N_12675);
nand U12832 (N_12832,N_12705,N_12662);
nor U12833 (N_12833,N_12660,N_12723);
and U12834 (N_12834,N_12625,N_12652);
and U12835 (N_12835,N_12736,N_12666);
nand U12836 (N_12836,N_12684,N_12729);
xor U12837 (N_12837,N_12706,N_12659);
and U12838 (N_12838,N_12687,N_12713);
and U12839 (N_12839,N_12652,N_12717);
and U12840 (N_12840,N_12665,N_12651);
nor U12841 (N_12841,N_12737,N_12672);
and U12842 (N_12842,N_12745,N_12658);
xnor U12843 (N_12843,N_12730,N_12723);
nand U12844 (N_12844,N_12716,N_12706);
or U12845 (N_12845,N_12630,N_12637);
and U12846 (N_12846,N_12626,N_12698);
nor U12847 (N_12847,N_12650,N_12681);
or U12848 (N_12848,N_12735,N_12703);
or U12849 (N_12849,N_12697,N_12701);
or U12850 (N_12850,N_12688,N_12681);
or U12851 (N_12851,N_12647,N_12737);
xor U12852 (N_12852,N_12636,N_12630);
nand U12853 (N_12853,N_12700,N_12741);
and U12854 (N_12854,N_12681,N_12675);
or U12855 (N_12855,N_12659,N_12647);
nor U12856 (N_12856,N_12686,N_12667);
nand U12857 (N_12857,N_12678,N_12642);
nor U12858 (N_12858,N_12736,N_12641);
or U12859 (N_12859,N_12677,N_12658);
and U12860 (N_12860,N_12687,N_12652);
nand U12861 (N_12861,N_12731,N_12655);
nand U12862 (N_12862,N_12630,N_12632);
nor U12863 (N_12863,N_12671,N_12630);
nand U12864 (N_12864,N_12676,N_12645);
nand U12865 (N_12865,N_12748,N_12665);
or U12866 (N_12866,N_12634,N_12688);
nand U12867 (N_12867,N_12627,N_12735);
xnor U12868 (N_12868,N_12645,N_12738);
or U12869 (N_12869,N_12741,N_12671);
xnor U12870 (N_12870,N_12688,N_12636);
or U12871 (N_12871,N_12744,N_12746);
xor U12872 (N_12872,N_12656,N_12670);
or U12873 (N_12873,N_12743,N_12648);
nor U12874 (N_12874,N_12694,N_12658);
and U12875 (N_12875,N_12871,N_12782);
and U12876 (N_12876,N_12796,N_12854);
xnor U12877 (N_12877,N_12761,N_12798);
nor U12878 (N_12878,N_12865,N_12870);
xor U12879 (N_12879,N_12751,N_12855);
or U12880 (N_12880,N_12759,N_12793);
xnor U12881 (N_12881,N_12810,N_12773);
and U12882 (N_12882,N_12815,N_12802);
nand U12883 (N_12883,N_12752,N_12840);
and U12884 (N_12884,N_12852,N_12756);
nand U12885 (N_12885,N_12801,N_12771);
or U12886 (N_12886,N_12864,N_12785);
or U12887 (N_12887,N_12857,N_12772);
or U12888 (N_12888,N_12863,N_12812);
xor U12889 (N_12889,N_12769,N_12774);
or U12890 (N_12890,N_12779,N_12862);
nor U12891 (N_12891,N_12784,N_12795);
nor U12892 (N_12892,N_12754,N_12809);
nor U12893 (N_12893,N_12816,N_12781);
nor U12894 (N_12894,N_12858,N_12755);
and U12895 (N_12895,N_12753,N_12826);
and U12896 (N_12896,N_12758,N_12853);
or U12897 (N_12897,N_12845,N_12817);
xor U12898 (N_12898,N_12834,N_12767);
or U12899 (N_12899,N_12842,N_12778);
nand U12900 (N_12900,N_12764,N_12780);
or U12901 (N_12901,N_12803,N_12804);
or U12902 (N_12902,N_12846,N_12799);
and U12903 (N_12903,N_12807,N_12860);
xor U12904 (N_12904,N_12868,N_12828);
xnor U12905 (N_12905,N_12872,N_12797);
xor U12906 (N_12906,N_12848,N_12818);
xnor U12907 (N_12907,N_12788,N_12839);
nor U12908 (N_12908,N_12841,N_12762);
nand U12909 (N_12909,N_12829,N_12859);
nor U12910 (N_12910,N_12805,N_12856);
nor U12911 (N_12911,N_12808,N_12800);
and U12912 (N_12912,N_12763,N_12844);
xor U12913 (N_12913,N_12757,N_12823);
xnor U12914 (N_12914,N_12814,N_12791);
and U12915 (N_12915,N_12819,N_12867);
nor U12916 (N_12916,N_12837,N_12849);
xor U12917 (N_12917,N_12750,N_12806);
and U12918 (N_12918,N_12873,N_12833);
or U12919 (N_12919,N_12874,N_12786);
xor U12920 (N_12920,N_12825,N_12843);
xor U12921 (N_12921,N_12811,N_12765);
nand U12922 (N_12922,N_12820,N_12813);
xnor U12923 (N_12923,N_12866,N_12775);
or U12924 (N_12924,N_12861,N_12835);
nand U12925 (N_12925,N_12787,N_12831);
nor U12926 (N_12926,N_12790,N_12776);
nor U12927 (N_12927,N_12760,N_12827);
xnor U12928 (N_12928,N_12770,N_12792);
and U12929 (N_12929,N_12822,N_12824);
nor U12930 (N_12930,N_12783,N_12766);
xor U12931 (N_12931,N_12847,N_12777);
and U12932 (N_12932,N_12821,N_12869);
nor U12933 (N_12933,N_12832,N_12836);
and U12934 (N_12934,N_12768,N_12851);
or U12935 (N_12935,N_12789,N_12830);
xnor U12936 (N_12936,N_12838,N_12794);
nand U12937 (N_12937,N_12850,N_12859);
nor U12938 (N_12938,N_12764,N_12784);
and U12939 (N_12939,N_12785,N_12856);
nor U12940 (N_12940,N_12778,N_12770);
nor U12941 (N_12941,N_12827,N_12762);
or U12942 (N_12942,N_12769,N_12829);
and U12943 (N_12943,N_12838,N_12868);
xor U12944 (N_12944,N_12831,N_12860);
or U12945 (N_12945,N_12792,N_12855);
nor U12946 (N_12946,N_12762,N_12776);
xor U12947 (N_12947,N_12772,N_12767);
xnor U12948 (N_12948,N_12810,N_12774);
or U12949 (N_12949,N_12775,N_12804);
or U12950 (N_12950,N_12861,N_12800);
and U12951 (N_12951,N_12823,N_12870);
nand U12952 (N_12952,N_12803,N_12830);
nor U12953 (N_12953,N_12779,N_12850);
xnor U12954 (N_12954,N_12824,N_12764);
and U12955 (N_12955,N_12805,N_12865);
and U12956 (N_12956,N_12823,N_12825);
nor U12957 (N_12957,N_12754,N_12805);
nor U12958 (N_12958,N_12766,N_12770);
or U12959 (N_12959,N_12827,N_12764);
nand U12960 (N_12960,N_12846,N_12756);
nand U12961 (N_12961,N_12780,N_12768);
nor U12962 (N_12962,N_12830,N_12752);
or U12963 (N_12963,N_12866,N_12779);
nor U12964 (N_12964,N_12847,N_12859);
or U12965 (N_12965,N_12838,N_12864);
xnor U12966 (N_12966,N_12837,N_12868);
nor U12967 (N_12967,N_12810,N_12869);
xor U12968 (N_12968,N_12859,N_12770);
nand U12969 (N_12969,N_12788,N_12765);
nor U12970 (N_12970,N_12790,N_12818);
nor U12971 (N_12971,N_12853,N_12830);
nand U12972 (N_12972,N_12751,N_12754);
or U12973 (N_12973,N_12766,N_12762);
nor U12974 (N_12974,N_12831,N_12760);
or U12975 (N_12975,N_12774,N_12754);
nor U12976 (N_12976,N_12834,N_12827);
nand U12977 (N_12977,N_12867,N_12802);
or U12978 (N_12978,N_12818,N_12855);
and U12979 (N_12979,N_12833,N_12870);
xor U12980 (N_12980,N_12825,N_12824);
and U12981 (N_12981,N_12860,N_12848);
or U12982 (N_12982,N_12777,N_12849);
or U12983 (N_12983,N_12797,N_12789);
or U12984 (N_12984,N_12850,N_12832);
or U12985 (N_12985,N_12812,N_12813);
nor U12986 (N_12986,N_12777,N_12843);
or U12987 (N_12987,N_12779,N_12852);
nand U12988 (N_12988,N_12842,N_12866);
xor U12989 (N_12989,N_12870,N_12755);
xnor U12990 (N_12990,N_12869,N_12809);
and U12991 (N_12991,N_12826,N_12857);
or U12992 (N_12992,N_12762,N_12781);
or U12993 (N_12993,N_12836,N_12848);
and U12994 (N_12994,N_12769,N_12816);
and U12995 (N_12995,N_12870,N_12845);
or U12996 (N_12996,N_12804,N_12809);
or U12997 (N_12997,N_12863,N_12838);
nor U12998 (N_12998,N_12832,N_12798);
nor U12999 (N_12999,N_12865,N_12758);
xor U13000 (N_13000,N_12890,N_12951);
and U13001 (N_13001,N_12918,N_12926);
xor U13002 (N_13002,N_12962,N_12914);
nand U13003 (N_13003,N_12973,N_12911);
and U13004 (N_13004,N_12898,N_12969);
nor U13005 (N_13005,N_12877,N_12909);
or U13006 (N_13006,N_12902,N_12875);
nand U13007 (N_13007,N_12976,N_12945);
nand U13008 (N_13008,N_12907,N_12982);
or U13009 (N_13009,N_12946,N_12955);
xnor U13010 (N_13010,N_12994,N_12998);
nor U13011 (N_13011,N_12983,N_12922);
nor U13012 (N_13012,N_12925,N_12903);
and U13013 (N_13013,N_12990,N_12933);
and U13014 (N_13014,N_12924,N_12993);
and U13015 (N_13015,N_12895,N_12893);
nand U13016 (N_13016,N_12901,N_12927);
or U13017 (N_13017,N_12992,N_12966);
nor U13018 (N_13018,N_12942,N_12880);
xor U13019 (N_13019,N_12931,N_12985);
or U13020 (N_13020,N_12972,N_12957);
or U13021 (N_13021,N_12935,N_12967);
xor U13022 (N_13022,N_12900,N_12944);
nor U13023 (N_13023,N_12971,N_12882);
xor U13024 (N_13024,N_12878,N_12958);
or U13025 (N_13025,N_12995,N_12965);
nor U13026 (N_13026,N_12941,N_12947);
nor U13027 (N_13027,N_12894,N_12968);
or U13028 (N_13028,N_12937,N_12889);
xor U13029 (N_13029,N_12928,N_12921);
nor U13030 (N_13030,N_12899,N_12987);
or U13031 (N_13031,N_12884,N_12879);
xor U13032 (N_13032,N_12939,N_12938);
or U13033 (N_13033,N_12930,N_12943);
xor U13034 (N_13034,N_12964,N_12940);
and U13035 (N_13035,N_12979,N_12988);
xor U13036 (N_13036,N_12991,N_12904);
nand U13037 (N_13037,N_12919,N_12963);
or U13038 (N_13038,N_12917,N_12989);
and U13039 (N_13039,N_12954,N_12913);
xor U13040 (N_13040,N_12912,N_12953);
xnor U13041 (N_13041,N_12887,N_12920);
nand U13042 (N_13042,N_12896,N_12975);
and U13043 (N_13043,N_12891,N_12950);
and U13044 (N_13044,N_12996,N_12905);
xnor U13045 (N_13045,N_12910,N_12949);
or U13046 (N_13046,N_12885,N_12908);
xnor U13047 (N_13047,N_12886,N_12888);
nor U13048 (N_13048,N_12906,N_12999);
nand U13049 (N_13049,N_12932,N_12916);
and U13050 (N_13050,N_12892,N_12978);
xor U13051 (N_13051,N_12929,N_12936);
or U13052 (N_13052,N_12881,N_12970);
and U13053 (N_13053,N_12977,N_12980);
nor U13054 (N_13054,N_12883,N_12876);
nand U13055 (N_13055,N_12934,N_12915);
or U13056 (N_13056,N_12897,N_12923);
and U13057 (N_13057,N_12959,N_12960);
nand U13058 (N_13058,N_12986,N_12997);
nand U13059 (N_13059,N_12974,N_12948);
or U13060 (N_13060,N_12956,N_12984);
xnor U13061 (N_13061,N_12952,N_12981);
or U13062 (N_13062,N_12961,N_12885);
xnor U13063 (N_13063,N_12962,N_12888);
nor U13064 (N_13064,N_12990,N_12914);
nand U13065 (N_13065,N_12981,N_12985);
nor U13066 (N_13066,N_12891,N_12928);
and U13067 (N_13067,N_12881,N_12934);
nand U13068 (N_13068,N_12942,N_12913);
xnor U13069 (N_13069,N_12894,N_12974);
or U13070 (N_13070,N_12904,N_12971);
nand U13071 (N_13071,N_12938,N_12953);
xnor U13072 (N_13072,N_12975,N_12947);
nand U13073 (N_13073,N_12935,N_12945);
xor U13074 (N_13074,N_12927,N_12961);
or U13075 (N_13075,N_12942,N_12891);
nand U13076 (N_13076,N_12938,N_12974);
nand U13077 (N_13077,N_12921,N_12927);
xor U13078 (N_13078,N_12907,N_12991);
or U13079 (N_13079,N_12884,N_12989);
or U13080 (N_13080,N_12892,N_12893);
nand U13081 (N_13081,N_12881,N_12880);
nor U13082 (N_13082,N_12987,N_12891);
xor U13083 (N_13083,N_12904,N_12875);
nor U13084 (N_13084,N_12966,N_12895);
nor U13085 (N_13085,N_12920,N_12905);
and U13086 (N_13086,N_12875,N_12990);
and U13087 (N_13087,N_12922,N_12977);
or U13088 (N_13088,N_12959,N_12896);
nand U13089 (N_13089,N_12897,N_12928);
xor U13090 (N_13090,N_12922,N_12981);
nor U13091 (N_13091,N_12903,N_12904);
nand U13092 (N_13092,N_12881,N_12964);
nor U13093 (N_13093,N_12906,N_12984);
and U13094 (N_13094,N_12929,N_12969);
xor U13095 (N_13095,N_12968,N_12958);
and U13096 (N_13096,N_12880,N_12991);
and U13097 (N_13097,N_12969,N_12930);
or U13098 (N_13098,N_12953,N_12928);
or U13099 (N_13099,N_12921,N_12924);
xor U13100 (N_13100,N_12903,N_12954);
xor U13101 (N_13101,N_12954,N_12877);
nand U13102 (N_13102,N_12897,N_12938);
or U13103 (N_13103,N_12891,N_12897);
and U13104 (N_13104,N_12883,N_12973);
or U13105 (N_13105,N_12931,N_12884);
and U13106 (N_13106,N_12971,N_12884);
nor U13107 (N_13107,N_12893,N_12975);
xnor U13108 (N_13108,N_12888,N_12988);
nor U13109 (N_13109,N_12972,N_12878);
and U13110 (N_13110,N_12905,N_12988);
or U13111 (N_13111,N_12901,N_12952);
nand U13112 (N_13112,N_12930,N_12886);
nor U13113 (N_13113,N_12955,N_12934);
and U13114 (N_13114,N_12903,N_12977);
nor U13115 (N_13115,N_12900,N_12904);
nand U13116 (N_13116,N_12930,N_12950);
and U13117 (N_13117,N_12889,N_12964);
nand U13118 (N_13118,N_12900,N_12974);
nor U13119 (N_13119,N_12913,N_12996);
and U13120 (N_13120,N_12973,N_12896);
nor U13121 (N_13121,N_12921,N_12903);
nor U13122 (N_13122,N_12965,N_12894);
and U13123 (N_13123,N_12918,N_12985);
nand U13124 (N_13124,N_12949,N_12973);
and U13125 (N_13125,N_13028,N_13116);
or U13126 (N_13126,N_13069,N_13081);
xor U13127 (N_13127,N_13009,N_13063);
xor U13128 (N_13128,N_13060,N_13035);
xnor U13129 (N_13129,N_13062,N_13108);
xnor U13130 (N_13130,N_13003,N_13054);
or U13131 (N_13131,N_13068,N_13077);
nor U13132 (N_13132,N_13061,N_13090);
nand U13133 (N_13133,N_13098,N_13095);
nor U13134 (N_13134,N_13039,N_13000);
and U13135 (N_13135,N_13008,N_13021);
nand U13136 (N_13136,N_13030,N_13002);
xnor U13137 (N_13137,N_13010,N_13111);
nand U13138 (N_13138,N_13047,N_13089);
or U13139 (N_13139,N_13087,N_13018);
nand U13140 (N_13140,N_13123,N_13092);
nand U13141 (N_13141,N_13013,N_13033);
or U13142 (N_13142,N_13056,N_13029);
nand U13143 (N_13143,N_13020,N_13122);
nor U13144 (N_13144,N_13058,N_13074);
and U13145 (N_13145,N_13079,N_13032);
and U13146 (N_13146,N_13011,N_13048);
and U13147 (N_13147,N_13042,N_13088);
nand U13148 (N_13148,N_13045,N_13104);
nor U13149 (N_13149,N_13066,N_13118);
or U13150 (N_13150,N_13076,N_13036);
xnor U13151 (N_13151,N_13043,N_13006);
nand U13152 (N_13152,N_13083,N_13073);
or U13153 (N_13153,N_13110,N_13055);
xnor U13154 (N_13154,N_13064,N_13016);
nor U13155 (N_13155,N_13014,N_13107);
nand U13156 (N_13156,N_13099,N_13115);
nand U13157 (N_13157,N_13075,N_13017);
or U13158 (N_13158,N_13001,N_13027);
nor U13159 (N_13159,N_13007,N_13019);
and U13160 (N_13160,N_13091,N_13084);
or U13161 (N_13161,N_13025,N_13094);
or U13162 (N_13162,N_13004,N_13093);
nand U13163 (N_13163,N_13080,N_13102);
xor U13164 (N_13164,N_13034,N_13112);
and U13165 (N_13165,N_13082,N_13096);
nand U13166 (N_13166,N_13109,N_13023);
nand U13167 (N_13167,N_13038,N_13057);
nand U13168 (N_13168,N_13124,N_13106);
or U13169 (N_13169,N_13051,N_13053);
nor U13170 (N_13170,N_13119,N_13072);
xnor U13171 (N_13171,N_13059,N_13067);
or U13172 (N_13172,N_13101,N_13100);
or U13173 (N_13173,N_13012,N_13050);
nor U13174 (N_13174,N_13120,N_13113);
nand U13175 (N_13175,N_13037,N_13097);
nand U13176 (N_13176,N_13078,N_13086);
and U13177 (N_13177,N_13103,N_13065);
and U13178 (N_13178,N_13117,N_13046);
or U13179 (N_13179,N_13114,N_13052);
xnor U13180 (N_13180,N_13022,N_13070);
nor U13181 (N_13181,N_13041,N_13085);
nor U13182 (N_13182,N_13105,N_13005);
nand U13183 (N_13183,N_13040,N_13044);
or U13184 (N_13184,N_13071,N_13015);
nand U13185 (N_13185,N_13049,N_13031);
nor U13186 (N_13186,N_13026,N_13024);
and U13187 (N_13187,N_13121,N_13042);
nand U13188 (N_13188,N_13027,N_13049);
and U13189 (N_13189,N_13011,N_13118);
nor U13190 (N_13190,N_13026,N_13118);
nand U13191 (N_13191,N_13069,N_13045);
nand U13192 (N_13192,N_13055,N_13015);
xor U13193 (N_13193,N_13096,N_13083);
nand U13194 (N_13194,N_13028,N_13023);
nor U13195 (N_13195,N_13115,N_13110);
or U13196 (N_13196,N_13106,N_13081);
nor U13197 (N_13197,N_13005,N_13062);
or U13198 (N_13198,N_13058,N_13008);
and U13199 (N_13199,N_13116,N_13106);
xnor U13200 (N_13200,N_13031,N_13019);
xor U13201 (N_13201,N_13104,N_13105);
xnor U13202 (N_13202,N_13114,N_13039);
or U13203 (N_13203,N_13030,N_13003);
and U13204 (N_13204,N_13010,N_13066);
or U13205 (N_13205,N_13108,N_13033);
xor U13206 (N_13206,N_13051,N_13102);
nand U13207 (N_13207,N_13112,N_13117);
or U13208 (N_13208,N_13005,N_13010);
and U13209 (N_13209,N_13029,N_13108);
nor U13210 (N_13210,N_13073,N_13070);
and U13211 (N_13211,N_13020,N_13040);
and U13212 (N_13212,N_13061,N_13046);
or U13213 (N_13213,N_13082,N_13019);
nor U13214 (N_13214,N_13011,N_13055);
or U13215 (N_13215,N_13041,N_13023);
nor U13216 (N_13216,N_13004,N_13083);
and U13217 (N_13217,N_13110,N_13071);
and U13218 (N_13218,N_13088,N_13066);
and U13219 (N_13219,N_13088,N_13046);
nand U13220 (N_13220,N_13124,N_13090);
or U13221 (N_13221,N_13067,N_13009);
nor U13222 (N_13222,N_13051,N_13030);
nand U13223 (N_13223,N_13046,N_13085);
nand U13224 (N_13224,N_13005,N_13030);
nand U13225 (N_13225,N_13057,N_13110);
nand U13226 (N_13226,N_13026,N_13039);
nand U13227 (N_13227,N_13028,N_13090);
xnor U13228 (N_13228,N_13023,N_13074);
xnor U13229 (N_13229,N_13051,N_13076);
nor U13230 (N_13230,N_13053,N_13120);
nor U13231 (N_13231,N_13017,N_13058);
or U13232 (N_13232,N_13097,N_13103);
nand U13233 (N_13233,N_13010,N_13110);
or U13234 (N_13234,N_13115,N_13020);
xnor U13235 (N_13235,N_13124,N_13052);
or U13236 (N_13236,N_13020,N_13071);
nand U13237 (N_13237,N_13060,N_13044);
xor U13238 (N_13238,N_13121,N_13103);
xor U13239 (N_13239,N_13104,N_13114);
and U13240 (N_13240,N_13005,N_13063);
and U13241 (N_13241,N_13086,N_13022);
nand U13242 (N_13242,N_13071,N_13108);
xnor U13243 (N_13243,N_13075,N_13006);
and U13244 (N_13244,N_13119,N_13014);
or U13245 (N_13245,N_13089,N_13078);
nor U13246 (N_13246,N_13062,N_13111);
nor U13247 (N_13247,N_13080,N_13001);
nand U13248 (N_13248,N_13017,N_13092);
nand U13249 (N_13249,N_13085,N_13103);
nor U13250 (N_13250,N_13198,N_13160);
nor U13251 (N_13251,N_13155,N_13159);
nor U13252 (N_13252,N_13143,N_13168);
nand U13253 (N_13253,N_13189,N_13210);
or U13254 (N_13254,N_13178,N_13208);
or U13255 (N_13255,N_13230,N_13129);
or U13256 (N_13256,N_13233,N_13206);
xnor U13257 (N_13257,N_13238,N_13172);
or U13258 (N_13258,N_13245,N_13135);
xor U13259 (N_13259,N_13185,N_13144);
nor U13260 (N_13260,N_13240,N_13153);
nor U13261 (N_13261,N_13186,N_13202);
and U13262 (N_13262,N_13215,N_13231);
or U13263 (N_13263,N_13192,N_13229);
nor U13264 (N_13264,N_13241,N_13214);
or U13265 (N_13265,N_13128,N_13145);
nor U13266 (N_13266,N_13171,N_13187);
nand U13267 (N_13267,N_13176,N_13239);
or U13268 (N_13268,N_13242,N_13223);
xnor U13269 (N_13269,N_13225,N_13209);
xnor U13270 (N_13270,N_13184,N_13150);
and U13271 (N_13271,N_13125,N_13213);
nor U13272 (N_13272,N_13181,N_13134);
and U13273 (N_13273,N_13126,N_13156);
or U13274 (N_13274,N_13132,N_13169);
nor U13275 (N_13275,N_13246,N_13152);
and U13276 (N_13276,N_13190,N_13179);
and U13277 (N_13277,N_13201,N_13147);
nand U13278 (N_13278,N_13221,N_13248);
nor U13279 (N_13279,N_13130,N_13157);
nand U13280 (N_13280,N_13235,N_13183);
or U13281 (N_13281,N_13218,N_13205);
xor U13282 (N_13282,N_13194,N_13220);
nor U13283 (N_13283,N_13149,N_13234);
and U13284 (N_13284,N_13136,N_13211);
nand U13285 (N_13285,N_13127,N_13133);
and U13286 (N_13286,N_13154,N_13222);
nand U13287 (N_13287,N_13228,N_13188);
and U13288 (N_13288,N_13217,N_13203);
xnor U13289 (N_13289,N_13139,N_13193);
nand U13290 (N_13290,N_13226,N_13164);
xnor U13291 (N_13291,N_13236,N_13174);
nor U13292 (N_13292,N_13142,N_13216);
or U13293 (N_13293,N_13244,N_13232);
and U13294 (N_13294,N_13162,N_13237);
xnor U13295 (N_13295,N_13196,N_13175);
nor U13296 (N_13296,N_13151,N_13166);
xor U13297 (N_13297,N_13195,N_13191);
nand U13298 (N_13298,N_13200,N_13141);
or U13299 (N_13299,N_13204,N_13249);
nand U13300 (N_13300,N_13167,N_13137);
or U13301 (N_13301,N_13140,N_13227);
or U13302 (N_13302,N_13197,N_13161);
xnor U13303 (N_13303,N_13138,N_13177);
nor U13304 (N_13304,N_13146,N_13131);
nand U13305 (N_13305,N_13224,N_13180);
and U13306 (N_13306,N_13207,N_13148);
and U13307 (N_13307,N_13170,N_13243);
nand U13308 (N_13308,N_13247,N_13199);
nor U13309 (N_13309,N_13219,N_13158);
nor U13310 (N_13310,N_13165,N_13212);
or U13311 (N_13311,N_13163,N_13182);
or U13312 (N_13312,N_13173,N_13241);
xnor U13313 (N_13313,N_13229,N_13181);
and U13314 (N_13314,N_13209,N_13241);
nor U13315 (N_13315,N_13137,N_13221);
and U13316 (N_13316,N_13236,N_13149);
and U13317 (N_13317,N_13228,N_13172);
or U13318 (N_13318,N_13229,N_13175);
nand U13319 (N_13319,N_13155,N_13210);
xor U13320 (N_13320,N_13221,N_13138);
and U13321 (N_13321,N_13189,N_13147);
nor U13322 (N_13322,N_13202,N_13126);
xor U13323 (N_13323,N_13157,N_13216);
xnor U13324 (N_13324,N_13227,N_13197);
and U13325 (N_13325,N_13156,N_13221);
nor U13326 (N_13326,N_13207,N_13239);
nand U13327 (N_13327,N_13225,N_13202);
xnor U13328 (N_13328,N_13185,N_13223);
nor U13329 (N_13329,N_13151,N_13132);
nand U13330 (N_13330,N_13239,N_13169);
nand U13331 (N_13331,N_13162,N_13134);
nand U13332 (N_13332,N_13212,N_13161);
nor U13333 (N_13333,N_13203,N_13214);
and U13334 (N_13334,N_13143,N_13198);
or U13335 (N_13335,N_13187,N_13166);
nor U13336 (N_13336,N_13218,N_13129);
and U13337 (N_13337,N_13204,N_13201);
or U13338 (N_13338,N_13246,N_13170);
or U13339 (N_13339,N_13133,N_13214);
nand U13340 (N_13340,N_13162,N_13222);
xor U13341 (N_13341,N_13227,N_13174);
or U13342 (N_13342,N_13186,N_13237);
and U13343 (N_13343,N_13202,N_13183);
or U13344 (N_13344,N_13230,N_13209);
xor U13345 (N_13345,N_13194,N_13128);
nor U13346 (N_13346,N_13153,N_13188);
or U13347 (N_13347,N_13208,N_13166);
or U13348 (N_13348,N_13129,N_13164);
nor U13349 (N_13349,N_13175,N_13221);
or U13350 (N_13350,N_13133,N_13168);
xnor U13351 (N_13351,N_13240,N_13195);
nand U13352 (N_13352,N_13161,N_13135);
or U13353 (N_13353,N_13220,N_13151);
and U13354 (N_13354,N_13154,N_13223);
xnor U13355 (N_13355,N_13176,N_13127);
nor U13356 (N_13356,N_13130,N_13221);
xnor U13357 (N_13357,N_13194,N_13221);
nand U13358 (N_13358,N_13218,N_13130);
and U13359 (N_13359,N_13233,N_13241);
and U13360 (N_13360,N_13228,N_13178);
or U13361 (N_13361,N_13206,N_13209);
nand U13362 (N_13362,N_13190,N_13180);
and U13363 (N_13363,N_13244,N_13233);
nand U13364 (N_13364,N_13162,N_13210);
and U13365 (N_13365,N_13204,N_13217);
xor U13366 (N_13366,N_13159,N_13143);
nand U13367 (N_13367,N_13193,N_13247);
or U13368 (N_13368,N_13212,N_13130);
nor U13369 (N_13369,N_13243,N_13247);
or U13370 (N_13370,N_13199,N_13191);
or U13371 (N_13371,N_13149,N_13202);
or U13372 (N_13372,N_13207,N_13203);
xor U13373 (N_13373,N_13156,N_13137);
and U13374 (N_13374,N_13230,N_13227);
and U13375 (N_13375,N_13339,N_13329);
and U13376 (N_13376,N_13286,N_13256);
nor U13377 (N_13377,N_13283,N_13328);
and U13378 (N_13378,N_13373,N_13290);
nor U13379 (N_13379,N_13297,N_13354);
nor U13380 (N_13380,N_13370,N_13344);
or U13381 (N_13381,N_13285,N_13306);
nand U13382 (N_13382,N_13369,N_13259);
xor U13383 (N_13383,N_13357,N_13337);
nand U13384 (N_13384,N_13257,N_13365);
or U13385 (N_13385,N_13335,N_13363);
nand U13386 (N_13386,N_13276,N_13287);
and U13387 (N_13387,N_13350,N_13308);
nand U13388 (N_13388,N_13364,N_13318);
and U13389 (N_13389,N_13343,N_13299);
or U13390 (N_13390,N_13271,N_13278);
nand U13391 (N_13391,N_13345,N_13289);
or U13392 (N_13392,N_13303,N_13347);
xor U13393 (N_13393,N_13266,N_13258);
nand U13394 (N_13394,N_13355,N_13300);
nand U13395 (N_13395,N_13307,N_13313);
and U13396 (N_13396,N_13291,N_13274);
nand U13397 (N_13397,N_13255,N_13295);
xnor U13398 (N_13398,N_13250,N_13284);
xor U13399 (N_13399,N_13314,N_13324);
nor U13400 (N_13400,N_13260,N_13315);
or U13401 (N_13401,N_13263,N_13270);
and U13402 (N_13402,N_13273,N_13342);
and U13403 (N_13403,N_13275,N_13332);
nor U13404 (N_13404,N_13262,N_13277);
xor U13405 (N_13405,N_13265,N_13305);
or U13406 (N_13406,N_13252,N_13280);
nor U13407 (N_13407,N_13288,N_13323);
nand U13408 (N_13408,N_13268,N_13272);
nand U13409 (N_13409,N_13304,N_13309);
xor U13410 (N_13410,N_13359,N_13374);
or U13411 (N_13411,N_13294,N_13341);
or U13412 (N_13412,N_13253,N_13327);
and U13413 (N_13413,N_13302,N_13367);
xor U13414 (N_13414,N_13310,N_13361);
nand U13415 (N_13415,N_13330,N_13267);
or U13416 (N_13416,N_13296,N_13311);
xor U13417 (N_13417,N_13338,N_13321);
nand U13418 (N_13418,N_13349,N_13312);
xor U13419 (N_13419,N_13322,N_13372);
and U13420 (N_13420,N_13261,N_13320);
xnor U13421 (N_13421,N_13316,N_13351);
nor U13422 (N_13422,N_13319,N_13366);
nand U13423 (N_13423,N_13356,N_13251);
nand U13424 (N_13424,N_13264,N_13281);
nand U13425 (N_13425,N_13336,N_13333);
and U13426 (N_13426,N_13279,N_13353);
and U13427 (N_13427,N_13360,N_13298);
xnor U13428 (N_13428,N_13317,N_13293);
or U13429 (N_13429,N_13292,N_13334);
nor U13430 (N_13430,N_13282,N_13362);
nor U13431 (N_13431,N_13358,N_13269);
nand U13432 (N_13432,N_13346,N_13352);
nor U13433 (N_13433,N_13371,N_13331);
or U13434 (N_13434,N_13348,N_13254);
and U13435 (N_13435,N_13368,N_13326);
nand U13436 (N_13436,N_13340,N_13301);
and U13437 (N_13437,N_13325,N_13253);
nor U13438 (N_13438,N_13345,N_13344);
or U13439 (N_13439,N_13337,N_13306);
nand U13440 (N_13440,N_13339,N_13299);
or U13441 (N_13441,N_13315,N_13341);
xnor U13442 (N_13442,N_13367,N_13328);
xnor U13443 (N_13443,N_13272,N_13322);
and U13444 (N_13444,N_13282,N_13344);
nand U13445 (N_13445,N_13315,N_13251);
or U13446 (N_13446,N_13295,N_13316);
nand U13447 (N_13447,N_13262,N_13251);
nor U13448 (N_13448,N_13329,N_13314);
xor U13449 (N_13449,N_13373,N_13372);
nand U13450 (N_13450,N_13316,N_13344);
and U13451 (N_13451,N_13326,N_13350);
xnor U13452 (N_13452,N_13316,N_13365);
nand U13453 (N_13453,N_13332,N_13305);
or U13454 (N_13454,N_13265,N_13272);
and U13455 (N_13455,N_13273,N_13373);
or U13456 (N_13456,N_13281,N_13353);
xor U13457 (N_13457,N_13328,N_13349);
nor U13458 (N_13458,N_13272,N_13273);
or U13459 (N_13459,N_13293,N_13310);
or U13460 (N_13460,N_13264,N_13288);
nand U13461 (N_13461,N_13369,N_13270);
xor U13462 (N_13462,N_13344,N_13271);
or U13463 (N_13463,N_13365,N_13301);
or U13464 (N_13464,N_13263,N_13340);
nand U13465 (N_13465,N_13350,N_13266);
xor U13466 (N_13466,N_13325,N_13298);
and U13467 (N_13467,N_13366,N_13314);
nand U13468 (N_13468,N_13300,N_13298);
or U13469 (N_13469,N_13279,N_13360);
or U13470 (N_13470,N_13328,N_13325);
and U13471 (N_13471,N_13330,N_13320);
nand U13472 (N_13472,N_13262,N_13291);
and U13473 (N_13473,N_13311,N_13325);
or U13474 (N_13474,N_13284,N_13350);
nor U13475 (N_13475,N_13275,N_13337);
and U13476 (N_13476,N_13255,N_13333);
or U13477 (N_13477,N_13335,N_13259);
or U13478 (N_13478,N_13322,N_13359);
xor U13479 (N_13479,N_13314,N_13317);
or U13480 (N_13480,N_13345,N_13368);
nand U13481 (N_13481,N_13253,N_13324);
nor U13482 (N_13482,N_13300,N_13278);
or U13483 (N_13483,N_13281,N_13261);
nor U13484 (N_13484,N_13374,N_13343);
or U13485 (N_13485,N_13273,N_13280);
xnor U13486 (N_13486,N_13340,N_13251);
xor U13487 (N_13487,N_13299,N_13341);
xor U13488 (N_13488,N_13284,N_13293);
xnor U13489 (N_13489,N_13338,N_13354);
xor U13490 (N_13490,N_13354,N_13278);
xnor U13491 (N_13491,N_13364,N_13295);
nand U13492 (N_13492,N_13355,N_13334);
and U13493 (N_13493,N_13370,N_13257);
nand U13494 (N_13494,N_13256,N_13365);
nor U13495 (N_13495,N_13286,N_13255);
or U13496 (N_13496,N_13339,N_13338);
nor U13497 (N_13497,N_13266,N_13311);
or U13498 (N_13498,N_13256,N_13346);
and U13499 (N_13499,N_13368,N_13257);
nor U13500 (N_13500,N_13399,N_13460);
nand U13501 (N_13501,N_13435,N_13420);
nand U13502 (N_13502,N_13382,N_13376);
or U13503 (N_13503,N_13419,N_13473);
nor U13504 (N_13504,N_13395,N_13384);
nand U13505 (N_13505,N_13468,N_13408);
nand U13506 (N_13506,N_13471,N_13412);
or U13507 (N_13507,N_13387,N_13409);
nor U13508 (N_13508,N_13427,N_13440);
and U13509 (N_13509,N_13451,N_13452);
xor U13510 (N_13510,N_13375,N_13443);
or U13511 (N_13511,N_13400,N_13398);
or U13512 (N_13512,N_13470,N_13441);
or U13513 (N_13513,N_13424,N_13403);
nor U13514 (N_13514,N_13458,N_13456);
nand U13515 (N_13515,N_13494,N_13411);
and U13516 (N_13516,N_13430,N_13465);
and U13517 (N_13517,N_13439,N_13428);
or U13518 (N_13518,N_13417,N_13380);
and U13519 (N_13519,N_13481,N_13394);
nand U13520 (N_13520,N_13476,N_13457);
nand U13521 (N_13521,N_13447,N_13378);
xor U13522 (N_13522,N_13423,N_13467);
xor U13523 (N_13523,N_13464,N_13461);
nor U13524 (N_13524,N_13416,N_13446);
xnor U13525 (N_13525,N_13478,N_13449);
nor U13526 (N_13526,N_13377,N_13425);
nor U13527 (N_13527,N_13491,N_13472);
or U13528 (N_13528,N_13381,N_13393);
nand U13529 (N_13529,N_13442,N_13485);
nor U13530 (N_13530,N_13407,N_13390);
nor U13531 (N_13531,N_13397,N_13421);
or U13532 (N_13532,N_13474,N_13498);
nor U13533 (N_13533,N_13492,N_13463);
nor U13534 (N_13534,N_13422,N_13448);
nand U13535 (N_13535,N_13454,N_13402);
nand U13536 (N_13536,N_13445,N_13482);
nor U13537 (N_13537,N_13405,N_13455);
nand U13538 (N_13538,N_13432,N_13396);
and U13539 (N_13539,N_13450,N_13389);
nand U13540 (N_13540,N_13386,N_13434);
xor U13541 (N_13541,N_13383,N_13486);
nand U13542 (N_13542,N_13437,N_13497);
xnor U13543 (N_13543,N_13490,N_13433);
or U13544 (N_13544,N_13436,N_13388);
and U13545 (N_13545,N_13438,N_13493);
and U13546 (N_13546,N_13410,N_13379);
xnor U13547 (N_13547,N_13431,N_13496);
nor U13548 (N_13548,N_13444,N_13499);
or U13549 (N_13549,N_13480,N_13406);
nand U13550 (N_13550,N_13426,N_13477);
xnor U13551 (N_13551,N_13466,N_13404);
or U13552 (N_13552,N_13489,N_13413);
nand U13553 (N_13553,N_13414,N_13429);
nor U13554 (N_13554,N_13392,N_13418);
and U13555 (N_13555,N_13495,N_13401);
and U13556 (N_13556,N_13479,N_13488);
or U13557 (N_13557,N_13483,N_13453);
and U13558 (N_13558,N_13415,N_13459);
nand U13559 (N_13559,N_13475,N_13391);
and U13560 (N_13560,N_13462,N_13484);
xor U13561 (N_13561,N_13469,N_13385);
xor U13562 (N_13562,N_13487,N_13489);
nand U13563 (N_13563,N_13432,N_13499);
nor U13564 (N_13564,N_13410,N_13433);
or U13565 (N_13565,N_13492,N_13447);
or U13566 (N_13566,N_13491,N_13396);
or U13567 (N_13567,N_13409,N_13453);
nand U13568 (N_13568,N_13473,N_13381);
nor U13569 (N_13569,N_13380,N_13446);
nor U13570 (N_13570,N_13428,N_13379);
nand U13571 (N_13571,N_13430,N_13443);
or U13572 (N_13572,N_13486,N_13484);
nor U13573 (N_13573,N_13434,N_13403);
or U13574 (N_13574,N_13487,N_13385);
xor U13575 (N_13575,N_13471,N_13462);
and U13576 (N_13576,N_13424,N_13426);
nand U13577 (N_13577,N_13477,N_13407);
nor U13578 (N_13578,N_13403,N_13381);
and U13579 (N_13579,N_13471,N_13409);
xor U13580 (N_13580,N_13457,N_13385);
xnor U13581 (N_13581,N_13418,N_13390);
nand U13582 (N_13582,N_13431,N_13489);
nor U13583 (N_13583,N_13427,N_13447);
nor U13584 (N_13584,N_13458,N_13386);
xor U13585 (N_13585,N_13399,N_13483);
or U13586 (N_13586,N_13473,N_13498);
or U13587 (N_13587,N_13424,N_13433);
nor U13588 (N_13588,N_13429,N_13415);
nand U13589 (N_13589,N_13438,N_13469);
nor U13590 (N_13590,N_13377,N_13452);
or U13591 (N_13591,N_13482,N_13499);
and U13592 (N_13592,N_13496,N_13449);
or U13593 (N_13593,N_13457,N_13482);
and U13594 (N_13594,N_13407,N_13487);
or U13595 (N_13595,N_13404,N_13395);
nor U13596 (N_13596,N_13474,N_13428);
and U13597 (N_13597,N_13446,N_13477);
nand U13598 (N_13598,N_13452,N_13393);
nand U13599 (N_13599,N_13421,N_13489);
and U13600 (N_13600,N_13477,N_13499);
nor U13601 (N_13601,N_13482,N_13458);
nand U13602 (N_13602,N_13491,N_13402);
or U13603 (N_13603,N_13437,N_13457);
nand U13604 (N_13604,N_13475,N_13388);
nor U13605 (N_13605,N_13430,N_13496);
and U13606 (N_13606,N_13453,N_13412);
xor U13607 (N_13607,N_13425,N_13498);
nand U13608 (N_13608,N_13481,N_13406);
and U13609 (N_13609,N_13442,N_13499);
and U13610 (N_13610,N_13498,N_13461);
nor U13611 (N_13611,N_13497,N_13480);
or U13612 (N_13612,N_13382,N_13469);
and U13613 (N_13613,N_13393,N_13453);
nand U13614 (N_13614,N_13488,N_13437);
xor U13615 (N_13615,N_13421,N_13420);
xor U13616 (N_13616,N_13474,N_13392);
or U13617 (N_13617,N_13438,N_13472);
or U13618 (N_13618,N_13380,N_13445);
and U13619 (N_13619,N_13488,N_13418);
nand U13620 (N_13620,N_13487,N_13405);
nand U13621 (N_13621,N_13427,N_13472);
and U13622 (N_13622,N_13478,N_13416);
and U13623 (N_13623,N_13461,N_13459);
nor U13624 (N_13624,N_13375,N_13432);
or U13625 (N_13625,N_13622,N_13557);
or U13626 (N_13626,N_13547,N_13507);
nand U13627 (N_13627,N_13579,N_13609);
and U13628 (N_13628,N_13518,N_13586);
xor U13629 (N_13629,N_13590,N_13504);
nor U13630 (N_13630,N_13564,N_13551);
or U13631 (N_13631,N_13555,N_13591);
or U13632 (N_13632,N_13543,N_13566);
or U13633 (N_13633,N_13620,N_13524);
xor U13634 (N_13634,N_13501,N_13554);
or U13635 (N_13635,N_13572,N_13621);
nand U13636 (N_13636,N_13599,N_13528);
or U13637 (N_13637,N_13616,N_13530);
or U13638 (N_13638,N_13596,N_13527);
nor U13639 (N_13639,N_13559,N_13526);
nor U13640 (N_13640,N_13512,N_13513);
and U13641 (N_13641,N_13511,N_13515);
or U13642 (N_13642,N_13617,N_13583);
and U13643 (N_13643,N_13537,N_13510);
nor U13644 (N_13644,N_13538,N_13624);
nand U13645 (N_13645,N_13558,N_13552);
or U13646 (N_13646,N_13540,N_13613);
xor U13647 (N_13647,N_13567,N_13506);
nor U13648 (N_13648,N_13529,N_13556);
or U13649 (N_13649,N_13517,N_13605);
and U13650 (N_13650,N_13587,N_13600);
and U13651 (N_13651,N_13536,N_13585);
nand U13652 (N_13652,N_13508,N_13604);
nor U13653 (N_13653,N_13514,N_13588);
and U13654 (N_13654,N_13595,N_13582);
nor U13655 (N_13655,N_13577,N_13568);
xnor U13656 (N_13656,N_13520,N_13581);
nor U13657 (N_13657,N_13549,N_13570);
xor U13658 (N_13658,N_13531,N_13509);
nand U13659 (N_13659,N_13603,N_13619);
nand U13660 (N_13660,N_13548,N_13541);
or U13661 (N_13661,N_13578,N_13601);
nor U13662 (N_13662,N_13542,N_13544);
nand U13663 (N_13663,N_13505,N_13575);
nand U13664 (N_13664,N_13614,N_13606);
or U13665 (N_13665,N_13618,N_13584);
and U13666 (N_13666,N_13550,N_13576);
nor U13667 (N_13667,N_13610,N_13546);
or U13668 (N_13668,N_13503,N_13592);
nand U13669 (N_13669,N_13608,N_13597);
or U13670 (N_13670,N_13561,N_13589);
or U13671 (N_13671,N_13522,N_13563);
nor U13672 (N_13672,N_13539,N_13521);
xnor U13673 (N_13673,N_13598,N_13500);
xor U13674 (N_13674,N_13532,N_13502);
nor U13675 (N_13675,N_13615,N_13569);
and U13676 (N_13676,N_13553,N_13565);
and U13677 (N_13677,N_13535,N_13602);
or U13678 (N_13678,N_13594,N_13580);
nand U13679 (N_13679,N_13593,N_13562);
xor U13680 (N_13680,N_13574,N_13611);
or U13681 (N_13681,N_13534,N_13545);
and U13682 (N_13682,N_13525,N_13607);
xnor U13683 (N_13683,N_13523,N_13623);
nor U13684 (N_13684,N_13516,N_13519);
or U13685 (N_13685,N_13571,N_13560);
or U13686 (N_13686,N_13612,N_13573);
or U13687 (N_13687,N_13533,N_13617);
nand U13688 (N_13688,N_13605,N_13622);
nor U13689 (N_13689,N_13596,N_13613);
and U13690 (N_13690,N_13510,N_13594);
xor U13691 (N_13691,N_13617,N_13607);
nand U13692 (N_13692,N_13594,N_13624);
nor U13693 (N_13693,N_13618,N_13611);
nor U13694 (N_13694,N_13558,N_13575);
and U13695 (N_13695,N_13556,N_13520);
and U13696 (N_13696,N_13508,N_13523);
nor U13697 (N_13697,N_13612,N_13567);
xnor U13698 (N_13698,N_13528,N_13561);
and U13699 (N_13699,N_13501,N_13535);
and U13700 (N_13700,N_13552,N_13588);
and U13701 (N_13701,N_13542,N_13564);
nor U13702 (N_13702,N_13562,N_13584);
nor U13703 (N_13703,N_13530,N_13535);
or U13704 (N_13704,N_13500,N_13551);
xor U13705 (N_13705,N_13599,N_13611);
or U13706 (N_13706,N_13551,N_13503);
nand U13707 (N_13707,N_13535,N_13527);
nand U13708 (N_13708,N_13516,N_13556);
or U13709 (N_13709,N_13609,N_13596);
nand U13710 (N_13710,N_13551,N_13604);
nor U13711 (N_13711,N_13581,N_13595);
and U13712 (N_13712,N_13551,N_13621);
or U13713 (N_13713,N_13538,N_13501);
or U13714 (N_13714,N_13510,N_13506);
nand U13715 (N_13715,N_13504,N_13549);
and U13716 (N_13716,N_13500,N_13563);
xnor U13717 (N_13717,N_13538,N_13517);
nor U13718 (N_13718,N_13605,N_13621);
nand U13719 (N_13719,N_13574,N_13597);
and U13720 (N_13720,N_13578,N_13528);
or U13721 (N_13721,N_13508,N_13543);
xnor U13722 (N_13722,N_13606,N_13538);
xnor U13723 (N_13723,N_13574,N_13588);
and U13724 (N_13724,N_13531,N_13560);
and U13725 (N_13725,N_13533,N_13546);
or U13726 (N_13726,N_13615,N_13619);
and U13727 (N_13727,N_13552,N_13572);
nor U13728 (N_13728,N_13618,N_13529);
xor U13729 (N_13729,N_13580,N_13579);
and U13730 (N_13730,N_13621,N_13624);
nor U13731 (N_13731,N_13539,N_13583);
or U13732 (N_13732,N_13561,N_13565);
nor U13733 (N_13733,N_13612,N_13597);
or U13734 (N_13734,N_13614,N_13564);
or U13735 (N_13735,N_13580,N_13578);
nand U13736 (N_13736,N_13504,N_13587);
nor U13737 (N_13737,N_13559,N_13527);
nor U13738 (N_13738,N_13535,N_13603);
nand U13739 (N_13739,N_13572,N_13614);
or U13740 (N_13740,N_13529,N_13597);
nor U13741 (N_13741,N_13554,N_13507);
and U13742 (N_13742,N_13612,N_13575);
nand U13743 (N_13743,N_13599,N_13527);
or U13744 (N_13744,N_13502,N_13525);
nor U13745 (N_13745,N_13509,N_13540);
and U13746 (N_13746,N_13507,N_13607);
xnor U13747 (N_13747,N_13509,N_13599);
nand U13748 (N_13748,N_13540,N_13575);
and U13749 (N_13749,N_13604,N_13610);
xor U13750 (N_13750,N_13645,N_13715);
xor U13751 (N_13751,N_13734,N_13671);
nand U13752 (N_13752,N_13695,N_13631);
and U13753 (N_13753,N_13657,N_13655);
xor U13754 (N_13754,N_13635,N_13650);
xnor U13755 (N_13755,N_13720,N_13676);
nand U13756 (N_13756,N_13706,N_13738);
nand U13757 (N_13757,N_13670,N_13730);
nand U13758 (N_13758,N_13643,N_13626);
nor U13759 (N_13759,N_13628,N_13664);
or U13760 (N_13760,N_13639,N_13694);
nor U13761 (N_13761,N_13735,N_13659);
or U13762 (N_13762,N_13651,N_13633);
or U13763 (N_13763,N_13744,N_13685);
and U13764 (N_13764,N_13711,N_13736);
or U13765 (N_13765,N_13747,N_13649);
or U13766 (N_13766,N_13731,N_13686);
xor U13767 (N_13767,N_13644,N_13681);
nor U13768 (N_13768,N_13712,N_13646);
and U13769 (N_13769,N_13724,N_13678);
nand U13770 (N_13770,N_13718,N_13669);
nor U13771 (N_13771,N_13662,N_13691);
and U13772 (N_13772,N_13742,N_13689);
nor U13773 (N_13773,N_13668,N_13699);
nand U13774 (N_13774,N_13725,N_13665);
and U13775 (N_13775,N_13654,N_13647);
and U13776 (N_13776,N_13717,N_13625);
or U13777 (N_13777,N_13704,N_13656);
nand U13778 (N_13778,N_13746,N_13713);
xor U13779 (N_13779,N_13673,N_13702);
and U13780 (N_13780,N_13707,N_13677);
nor U13781 (N_13781,N_13728,N_13696);
and U13782 (N_13782,N_13630,N_13682);
or U13783 (N_13783,N_13692,N_13721);
nor U13784 (N_13784,N_13690,N_13674);
nand U13785 (N_13785,N_13688,N_13627);
nand U13786 (N_13786,N_13716,N_13672);
and U13787 (N_13787,N_13726,N_13661);
nor U13788 (N_13788,N_13653,N_13719);
and U13789 (N_13789,N_13680,N_13642);
or U13790 (N_13790,N_13660,N_13663);
xnor U13791 (N_13791,N_13698,N_13749);
xnor U13792 (N_13792,N_13727,N_13675);
nor U13793 (N_13793,N_13658,N_13666);
and U13794 (N_13794,N_13648,N_13636);
xnor U13795 (N_13795,N_13748,N_13714);
xor U13796 (N_13796,N_13743,N_13629);
or U13797 (N_13797,N_13722,N_13637);
or U13798 (N_13798,N_13733,N_13632);
or U13799 (N_13799,N_13710,N_13687);
xor U13800 (N_13800,N_13703,N_13700);
nor U13801 (N_13801,N_13693,N_13683);
and U13802 (N_13802,N_13679,N_13741);
and U13803 (N_13803,N_13640,N_13745);
or U13804 (N_13804,N_13697,N_13708);
nor U13805 (N_13805,N_13641,N_13684);
nand U13806 (N_13806,N_13732,N_13739);
and U13807 (N_13807,N_13740,N_13723);
nor U13808 (N_13808,N_13705,N_13638);
nand U13809 (N_13809,N_13709,N_13729);
nand U13810 (N_13810,N_13634,N_13667);
and U13811 (N_13811,N_13652,N_13701);
nand U13812 (N_13812,N_13737,N_13725);
nand U13813 (N_13813,N_13741,N_13672);
xnor U13814 (N_13814,N_13682,N_13678);
nand U13815 (N_13815,N_13680,N_13687);
xor U13816 (N_13816,N_13711,N_13636);
xor U13817 (N_13817,N_13659,N_13682);
or U13818 (N_13818,N_13663,N_13634);
xor U13819 (N_13819,N_13645,N_13707);
xor U13820 (N_13820,N_13673,N_13636);
nor U13821 (N_13821,N_13671,N_13730);
and U13822 (N_13822,N_13636,N_13709);
or U13823 (N_13823,N_13658,N_13713);
and U13824 (N_13824,N_13645,N_13640);
nor U13825 (N_13825,N_13645,N_13637);
and U13826 (N_13826,N_13719,N_13723);
xor U13827 (N_13827,N_13725,N_13726);
nand U13828 (N_13828,N_13697,N_13695);
nor U13829 (N_13829,N_13626,N_13722);
xnor U13830 (N_13830,N_13709,N_13646);
nand U13831 (N_13831,N_13716,N_13632);
and U13832 (N_13832,N_13721,N_13659);
or U13833 (N_13833,N_13639,N_13686);
nand U13834 (N_13834,N_13715,N_13660);
or U13835 (N_13835,N_13722,N_13723);
and U13836 (N_13836,N_13664,N_13709);
or U13837 (N_13837,N_13635,N_13633);
and U13838 (N_13838,N_13727,N_13740);
or U13839 (N_13839,N_13641,N_13640);
xor U13840 (N_13840,N_13745,N_13734);
nor U13841 (N_13841,N_13687,N_13724);
nor U13842 (N_13842,N_13640,N_13656);
and U13843 (N_13843,N_13672,N_13736);
and U13844 (N_13844,N_13735,N_13691);
or U13845 (N_13845,N_13671,N_13653);
and U13846 (N_13846,N_13702,N_13626);
nand U13847 (N_13847,N_13647,N_13735);
xor U13848 (N_13848,N_13677,N_13719);
xor U13849 (N_13849,N_13688,N_13733);
and U13850 (N_13850,N_13668,N_13631);
or U13851 (N_13851,N_13657,N_13629);
nand U13852 (N_13852,N_13681,N_13684);
xnor U13853 (N_13853,N_13736,N_13631);
xnor U13854 (N_13854,N_13719,N_13712);
nand U13855 (N_13855,N_13641,N_13704);
or U13856 (N_13856,N_13746,N_13699);
and U13857 (N_13857,N_13705,N_13634);
and U13858 (N_13858,N_13690,N_13711);
or U13859 (N_13859,N_13737,N_13671);
and U13860 (N_13860,N_13669,N_13662);
nor U13861 (N_13861,N_13723,N_13701);
xor U13862 (N_13862,N_13745,N_13692);
xnor U13863 (N_13863,N_13716,N_13711);
and U13864 (N_13864,N_13747,N_13667);
and U13865 (N_13865,N_13725,N_13674);
and U13866 (N_13866,N_13648,N_13695);
nand U13867 (N_13867,N_13636,N_13737);
xnor U13868 (N_13868,N_13662,N_13647);
nand U13869 (N_13869,N_13745,N_13685);
nand U13870 (N_13870,N_13651,N_13681);
nand U13871 (N_13871,N_13697,N_13734);
or U13872 (N_13872,N_13641,N_13717);
nor U13873 (N_13873,N_13721,N_13634);
nor U13874 (N_13874,N_13708,N_13657);
nand U13875 (N_13875,N_13841,N_13809);
nor U13876 (N_13876,N_13874,N_13799);
nand U13877 (N_13877,N_13859,N_13860);
or U13878 (N_13878,N_13770,N_13779);
or U13879 (N_13879,N_13840,N_13758);
or U13880 (N_13880,N_13793,N_13867);
xor U13881 (N_13881,N_13836,N_13826);
or U13882 (N_13882,N_13815,N_13750);
xnor U13883 (N_13883,N_13822,N_13763);
or U13884 (N_13884,N_13846,N_13842);
nand U13885 (N_13885,N_13767,N_13791);
nand U13886 (N_13886,N_13833,N_13796);
xnor U13887 (N_13887,N_13805,N_13760);
and U13888 (N_13888,N_13832,N_13835);
and U13889 (N_13889,N_13816,N_13771);
nand U13890 (N_13890,N_13777,N_13807);
nor U13891 (N_13891,N_13800,N_13863);
nor U13892 (N_13892,N_13825,N_13795);
or U13893 (N_13893,N_13818,N_13783);
or U13894 (N_13894,N_13787,N_13873);
nor U13895 (N_13895,N_13855,N_13849);
xor U13896 (N_13896,N_13801,N_13775);
nor U13897 (N_13897,N_13798,N_13811);
or U13898 (N_13898,N_13780,N_13751);
xnor U13899 (N_13899,N_13785,N_13768);
nor U13900 (N_13900,N_13766,N_13870);
nor U13901 (N_13901,N_13872,N_13790);
nor U13902 (N_13902,N_13865,N_13792);
xor U13903 (N_13903,N_13857,N_13828);
nand U13904 (N_13904,N_13845,N_13820);
nor U13905 (N_13905,N_13789,N_13814);
xor U13906 (N_13906,N_13843,N_13856);
nor U13907 (N_13907,N_13817,N_13827);
or U13908 (N_13908,N_13852,N_13824);
and U13909 (N_13909,N_13755,N_13830);
and U13910 (N_13910,N_13823,N_13869);
or U13911 (N_13911,N_13808,N_13784);
and U13912 (N_13912,N_13848,N_13821);
nand U13913 (N_13913,N_13773,N_13864);
and U13914 (N_13914,N_13810,N_13756);
and U13915 (N_13915,N_13861,N_13871);
xor U13916 (N_13916,N_13778,N_13802);
and U13917 (N_13917,N_13839,N_13772);
nand U13918 (N_13918,N_13837,N_13804);
nand U13919 (N_13919,N_13765,N_13812);
nand U13920 (N_13920,N_13847,N_13866);
nor U13921 (N_13921,N_13850,N_13769);
nand U13922 (N_13922,N_13762,N_13776);
and U13923 (N_13923,N_13854,N_13759);
and U13924 (N_13924,N_13774,N_13853);
or U13925 (N_13925,N_13813,N_13862);
xor U13926 (N_13926,N_13797,N_13788);
xor U13927 (N_13927,N_13794,N_13803);
nor U13928 (N_13928,N_13834,N_13868);
and U13929 (N_13929,N_13851,N_13781);
xnor U13930 (N_13930,N_13752,N_13831);
nor U13931 (N_13931,N_13806,N_13844);
or U13932 (N_13932,N_13782,N_13819);
and U13933 (N_13933,N_13757,N_13786);
xor U13934 (N_13934,N_13764,N_13753);
nand U13935 (N_13935,N_13829,N_13761);
nor U13936 (N_13936,N_13858,N_13838);
and U13937 (N_13937,N_13754,N_13842);
and U13938 (N_13938,N_13852,N_13785);
nor U13939 (N_13939,N_13805,N_13768);
nand U13940 (N_13940,N_13768,N_13801);
nand U13941 (N_13941,N_13840,N_13767);
and U13942 (N_13942,N_13787,N_13869);
nor U13943 (N_13943,N_13781,N_13874);
or U13944 (N_13944,N_13827,N_13839);
and U13945 (N_13945,N_13840,N_13813);
or U13946 (N_13946,N_13758,N_13829);
or U13947 (N_13947,N_13830,N_13774);
or U13948 (N_13948,N_13756,N_13860);
xnor U13949 (N_13949,N_13798,N_13765);
xnor U13950 (N_13950,N_13828,N_13812);
and U13951 (N_13951,N_13797,N_13784);
nor U13952 (N_13952,N_13846,N_13791);
xnor U13953 (N_13953,N_13843,N_13752);
xnor U13954 (N_13954,N_13858,N_13851);
nor U13955 (N_13955,N_13837,N_13815);
xnor U13956 (N_13956,N_13864,N_13840);
nand U13957 (N_13957,N_13812,N_13822);
or U13958 (N_13958,N_13847,N_13789);
xor U13959 (N_13959,N_13809,N_13837);
or U13960 (N_13960,N_13787,N_13765);
nor U13961 (N_13961,N_13829,N_13780);
xor U13962 (N_13962,N_13787,N_13837);
xor U13963 (N_13963,N_13779,N_13846);
and U13964 (N_13964,N_13778,N_13819);
and U13965 (N_13965,N_13840,N_13873);
or U13966 (N_13966,N_13791,N_13814);
xnor U13967 (N_13967,N_13767,N_13805);
nor U13968 (N_13968,N_13871,N_13831);
or U13969 (N_13969,N_13780,N_13873);
nor U13970 (N_13970,N_13807,N_13792);
nor U13971 (N_13971,N_13768,N_13769);
and U13972 (N_13972,N_13846,N_13864);
xnor U13973 (N_13973,N_13827,N_13765);
xnor U13974 (N_13974,N_13758,N_13873);
nand U13975 (N_13975,N_13845,N_13870);
nor U13976 (N_13976,N_13773,N_13776);
nor U13977 (N_13977,N_13773,N_13808);
or U13978 (N_13978,N_13819,N_13801);
nand U13979 (N_13979,N_13781,N_13833);
or U13980 (N_13980,N_13763,N_13813);
nand U13981 (N_13981,N_13863,N_13821);
nor U13982 (N_13982,N_13772,N_13768);
xor U13983 (N_13983,N_13846,N_13758);
and U13984 (N_13984,N_13852,N_13773);
nand U13985 (N_13985,N_13871,N_13765);
nand U13986 (N_13986,N_13750,N_13814);
nand U13987 (N_13987,N_13797,N_13842);
xor U13988 (N_13988,N_13765,N_13763);
nand U13989 (N_13989,N_13843,N_13811);
nor U13990 (N_13990,N_13795,N_13766);
nor U13991 (N_13991,N_13872,N_13806);
or U13992 (N_13992,N_13790,N_13857);
xor U13993 (N_13993,N_13752,N_13836);
or U13994 (N_13994,N_13752,N_13824);
or U13995 (N_13995,N_13805,N_13842);
nor U13996 (N_13996,N_13795,N_13818);
nand U13997 (N_13997,N_13792,N_13753);
or U13998 (N_13998,N_13772,N_13833);
or U13999 (N_13999,N_13810,N_13869);
nor U14000 (N_14000,N_13950,N_13996);
nor U14001 (N_14001,N_13899,N_13880);
nor U14002 (N_14002,N_13878,N_13978);
and U14003 (N_14003,N_13957,N_13985);
xnor U14004 (N_14004,N_13891,N_13912);
xor U14005 (N_14005,N_13917,N_13926);
and U14006 (N_14006,N_13902,N_13953);
nor U14007 (N_14007,N_13879,N_13935);
xor U14008 (N_14008,N_13882,N_13955);
and U14009 (N_14009,N_13921,N_13875);
and U14010 (N_14010,N_13889,N_13940);
and U14011 (N_14011,N_13909,N_13907);
and U14012 (N_14012,N_13973,N_13934);
or U14013 (N_14013,N_13901,N_13924);
or U14014 (N_14014,N_13881,N_13987);
nor U14015 (N_14015,N_13972,N_13937);
nor U14016 (N_14016,N_13960,N_13877);
xnor U14017 (N_14017,N_13896,N_13886);
xor U14018 (N_14018,N_13995,N_13908);
and U14019 (N_14019,N_13943,N_13983);
xnor U14020 (N_14020,N_13975,N_13962);
xor U14021 (N_14021,N_13903,N_13986);
xor U14022 (N_14022,N_13948,N_13936);
and U14023 (N_14023,N_13915,N_13954);
xor U14024 (N_14024,N_13885,N_13888);
and U14025 (N_14025,N_13989,N_13916);
nand U14026 (N_14026,N_13967,N_13894);
and U14027 (N_14027,N_13991,N_13970);
nand U14028 (N_14028,N_13958,N_13922);
and U14029 (N_14029,N_13981,N_13897);
nor U14030 (N_14030,N_13910,N_13923);
xnor U14031 (N_14031,N_13927,N_13999);
or U14032 (N_14032,N_13988,N_13944);
nor U14033 (N_14033,N_13900,N_13933);
nand U14034 (N_14034,N_13956,N_13980);
xnor U14035 (N_14035,N_13945,N_13977);
nor U14036 (N_14036,N_13914,N_13959);
xnor U14037 (N_14037,N_13992,N_13952);
and U14038 (N_14038,N_13994,N_13951);
nor U14039 (N_14039,N_13974,N_13876);
and U14040 (N_14040,N_13928,N_13942);
or U14041 (N_14041,N_13968,N_13890);
or U14042 (N_14042,N_13979,N_13941);
nor U14043 (N_14043,N_13895,N_13932);
or U14044 (N_14044,N_13984,N_13982);
nand U14045 (N_14045,N_13964,N_13919);
xor U14046 (N_14046,N_13993,N_13884);
or U14047 (N_14047,N_13898,N_13976);
xnor U14048 (N_14048,N_13969,N_13905);
xnor U14049 (N_14049,N_13946,N_13947);
xnor U14050 (N_14050,N_13997,N_13971);
nand U14051 (N_14051,N_13961,N_13918);
xor U14052 (N_14052,N_13930,N_13883);
nor U14053 (N_14053,N_13939,N_13913);
nand U14054 (N_14054,N_13929,N_13925);
nand U14055 (N_14055,N_13893,N_13906);
nor U14056 (N_14056,N_13931,N_13966);
xor U14057 (N_14057,N_13911,N_13887);
nor U14058 (N_14058,N_13963,N_13949);
nand U14059 (N_14059,N_13990,N_13904);
or U14060 (N_14060,N_13938,N_13920);
nand U14061 (N_14061,N_13998,N_13892);
nand U14062 (N_14062,N_13965,N_13949);
xnor U14063 (N_14063,N_13947,N_13911);
xor U14064 (N_14064,N_13983,N_13970);
nand U14065 (N_14065,N_13972,N_13992);
xor U14066 (N_14066,N_13974,N_13949);
xnor U14067 (N_14067,N_13897,N_13982);
nand U14068 (N_14068,N_13955,N_13961);
and U14069 (N_14069,N_13884,N_13920);
or U14070 (N_14070,N_13947,N_13926);
or U14071 (N_14071,N_13934,N_13960);
nand U14072 (N_14072,N_13903,N_13922);
nand U14073 (N_14073,N_13890,N_13969);
nor U14074 (N_14074,N_13878,N_13977);
xnor U14075 (N_14075,N_13944,N_13919);
nand U14076 (N_14076,N_13935,N_13916);
and U14077 (N_14077,N_13908,N_13977);
or U14078 (N_14078,N_13887,N_13912);
nand U14079 (N_14079,N_13924,N_13918);
or U14080 (N_14080,N_13940,N_13902);
nor U14081 (N_14081,N_13967,N_13983);
or U14082 (N_14082,N_13939,N_13901);
nor U14083 (N_14083,N_13905,N_13977);
and U14084 (N_14084,N_13934,N_13925);
xor U14085 (N_14085,N_13958,N_13997);
nor U14086 (N_14086,N_13915,N_13902);
or U14087 (N_14087,N_13994,N_13982);
nand U14088 (N_14088,N_13921,N_13913);
xor U14089 (N_14089,N_13884,N_13997);
nand U14090 (N_14090,N_13932,N_13986);
and U14091 (N_14091,N_13944,N_13875);
xnor U14092 (N_14092,N_13917,N_13988);
nor U14093 (N_14093,N_13978,N_13938);
nor U14094 (N_14094,N_13911,N_13877);
xor U14095 (N_14095,N_13947,N_13918);
or U14096 (N_14096,N_13896,N_13884);
nand U14097 (N_14097,N_13876,N_13926);
and U14098 (N_14098,N_13944,N_13892);
nor U14099 (N_14099,N_13982,N_13891);
and U14100 (N_14100,N_13890,N_13996);
or U14101 (N_14101,N_13998,N_13885);
and U14102 (N_14102,N_13880,N_13979);
and U14103 (N_14103,N_13904,N_13953);
and U14104 (N_14104,N_13966,N_13942);
nand U14105 (N_14105,N_13912,N_13953);
nor U14106 (N_14106,N_13904,N_13914);
nand U14107 (N_14107,N_13949,N_13970);
nor U14108 (N_14108,N_13936,N_13908);
nand U14109 (N_14109,N_13927,N_13907);
or U14110 (N_14110,N_13892,N_13965);
nor U14111 (N_14111,N_13877,N_13910);
xor U14112 (N_14112,N_13976,N_13881);
and U14113 (N_14113,N_13961,N_13898);
nand U14114 (N_14114,N_13919,N_13949);
nand U14115 (N_14115,N_13972,N_13952);
and U14116 (N_14116,N_13908,N_13998);
xnor U14117 (N_14117,N_13946,N_13994);
and U14118 (N_14118,N_13893,N_13980);
and U14119 (N_14119,N_13963,N_13982);
and U14120 (N_14120,N_13925,N_13979);
or U14121 (N_14121,N_13958,N_13931);
nor U14122 (N_14122,N_13921,N_13939);
or U14123 (N_14123,N_13930,N_13931);
nor U14124 (N_14124,N_13994,N_13957);
xor U14125 (N_14125,N_14096,N_14061);
xor U14126 (N_14126,N_14028,N_14033);
nand U14127 (N_14127,N_14070,N_14066);
nor U14128 (N_14128,N_14042,N_14000);
nand U14129 (N_14129,N_14054,N_14073);
nor U14130 (N_14130,N_14038,N_14108);
xnor U14131 (N_14131,N_14023,N_14122);
and U14132 (N_14132,N_14052,N_14046);
nor U14133 (N_14133,N_14090,N_14034);
or U14134 (N_14134,N_14124,N_14015);
xnor U14135 (N_14135,N_14100,N_14003);
or U14136 (N_14136,N_14056,N_14104);
and U14137 (N_14137,N_14018,N_14077);
nand U14138 (N_14138,N_14089,N_14059);
nand U14139 (N_14139,N_14094,N_14017);
nand U14140 (N_14140,N_14030,N_14012);
nand U14141 (N_14141,N_14113,N_14120);
nand U14142 (N_14142,N_14092,N_14020);
nor U14143 (N_14143,N_14080,N_14075);
nor U14144 (N_14144,N_14039,N_14024);
and U14145 (N_14145,N_14064,N_14116);
or U14146 (N_14146,N_14027,N_14121);
or U14147 (N_14147,N_14032,N_14019);
nand U14148 (N_14148,N_14041,N_14119);
or U14149 (N_14149,N_14026,N_14022);
nand U14150 (N_14150,N_14044,N_14060);
xor U14151 (N_14151,N_14049,N_14053);
and U14152 (N_14152,N_14010,N_14036);
and U14153 (N_14153,N_14114,N_14040);
nor U14154 (N_14154,N_14002,N_14101);
and U14155 (N_14155,N_14093,N_14016);
nor U14156 (N_14156,N_14037,N_14123);
nand U14157 (N_14157,N_14109,N_14081);
xnor U14158 (N_14158,N_14013,N_14014);
or U14159 (N_14159,N_14103,N_14082);
or U14160 (N_14160,N_14005,N_14099);
or U14161 (N_14161,N_14078,N_14079);
nor U14162 (N_14162,N_14098,N_14047);
xor U14163 (N_14163,N_14045,N_14097);
or U14164 (N_14164,N_14007,N_14063);
and U14165 (N_14165,N_14051,N_14058);
and U14166 (N_14166,N_14117,N_14006);
nand U14167 (N_14167,N_14110,N_14069);
or U14168 (N_14168,N_14084,N_14112);
or U14169 (N_14169,N_14102,N_14050);
nor U14170 (N_14170,N_14087,N_14068);
nor U14171 (N_14171,N_14083,N_14065);
nor U14172 (N_14172,N_14004,N_14029);
xnor U14173 (N_14173,N_14025,N_14111);
xor U14174 (N_14174,N_14001,N_14008);
xnor U14175 (N_14175,N_14071,N_14043);
and U14176 (N_14176,N_14076,N_14095);
nand U14177 (N_14177,N_14085,N_14118);
nand U14178 (N_14178,N_14031,N_14115);
nand U14179 (N_14179,N_14086,N_14055);
nand U14180 (N_14180,N_14035,N_14048);
nor U14181 (N_14181,N_14088,N_14067);
xnor U14182 (N_14182,N_14105,N_14009);
and U14183 (N_14183,N_14072,N_14106);
nand U14184 (N_14184,N_14057,N_14107);
nor U14185 (N_14185,N_14062,N_14011);
and U14186 (N_14186,N_14074,N_14091);
or U14187 (N_14187,N_14021,N_14062);
or U14188 (N_14188,N_14014,N_14028);
or U14189 (N_14189,N_14041,N_14022);
xnor U14190 (N_14190,N_14013,N_14119);
and U14191 (N_14191,N_14078,N_14076);
nand U14192 (N_14192,N_14074,N_14049);
xor U14193 (N_14193,N_14121,N_14075);
nand U14194 (N_14194,N_14043,N_14036);
xnor U14195 (N_14195,N_14108,N_14070);
and U14196 (N_14196,N_14101,N_14114);
or U14197 (N_14197,N_14051,N_14105);
and U14198 (N_14198,N_14085,N_14107);
and U14199 (N_14199,N_14071,N_14114);
nor U14200 (N_14200,N_14066,N_14018);
nand U14201 (N_14201,N_14045,N_14003);
and U14202 (N_14202,N_14112,N_14077);
xor U14203 (N_14203,N_14055,N_14096);
xor U14204 (N_14204,N_14070,N_14077);
nand U14205 (N_14205,N_14113,N_14038);
and U14206 (N_14206,N_14097,N_14041);
nor U14207 (N_14207,N_14026,N_14045);
nor U14208 (N_14208,N_14033,N_14104);
and U14209 (N_14209,N_14014,N_14080);
xnor U14210 (N_14210,N_14115,N_14071);
xnor U14211 (N_14211,N_14068,N_14095);
nand U14212 (N_14212,N_14027,N_14018);
and U14213 (N_14213,N_14009,N_14061);
nand U14214 (N_14214,N_14020,N_14075);
xnor U14215 (N_14215,N_14097,N_14051);
nor U14216 (N_14216,N_14065,N_14041);
and U14217 (N_14217,N_14045,N_14094);
nand U14218 (N_14218,N_14013,N_14107);
nor U14219 (N_14219,N_14064,N_14001);
nand U14220 (N_14220,N_14116,N_14044);
nor U14221 (N_14221,N_14061,N_14065);
nor U14222 (N_14222,N_14008,N_14084);
nand U14223 (N_14223,N_14069,N_14043);
or U14224 (N_14224,N_14033,N_14032);
or U14225 (N_14225,N_14023,N_14030);
nor U14226 (N_14226,N_14046,N_14088);
and U14227 (N_14227,N_14038,N_14115);
and U14228 (N_14228,N_14059,N_14011);
xnor U14229 (N_14229,N_14076,N_14030);
and U14230 (N_14230,N_14121,N_14074);
nand U14231 (N_14231,N_14057,N_14042);
nor U14232 (N_14232,N_14123,N_14069);
nand U14233 (N_14233,N_14012,N_14035);
xnor U14234 (N_14234,N_14091,N_14068);
nor U14235 (N_14235,N_14007,N_14054);
nor U14236 (N_14236,N_14025,N_14074);
or U14237 (N_14237,N_14085,N_14019);
nand U14238 (N_14238,N_14013,N_14102);
xor U14239 (N_14239,N_14119,N_14020);
nand U14240 (N_14240,N_14085,N_14047);
and U14241 (N_14241,N_14027,N_14032);
xor U14242 (N_14242,N_14036,N_14063);
nand U14243 (N_14243,N_14003,N_14124);
nand U14244 (N_14244,N_14074,N_14048);
and U14245 (N_14245,N_14087,N_14026);
xor U14246 (N_14246,N_14036,N_14038);
nor U14247 (N_14247,N_14106,N_14080);
xor U14248 (N_14248,N_14069,N_14098);
xor U14249 (N_14249,N_14032,N_14103);
nor U14250 (N_14250,N_14133,N_14154);
xnor U14251 (N_14251,N_14147,N_14175);
xor U14252 (N_14252,N_14162,N_14235);
nand U14253 (N_14253,N_14208,N_14189);
xor U14254 (N_14254,N_14229,N_14165);
and U14255 (N_14255,N_14231,N_14245);
and U14256 (N_14256,N_14180,N_14171);
or U14257 (N_14257,N_14155,N_14159);
xnor U14258 (N_14258,N_14221,N_14146);
xnor U14259 (N_14259,N_14148,N_14134);
and U14260 (N_14260,N_14220,N_14233);
nor U14261 (N_14261,N_14181,N_14217);
xor U14262 (N_14262,N_14164,N_14161);
nor U14263 (N_14263,N_14193,N_14152);
or U14264 (N_14264,N_14135,N_14169);
xnor U14265 (N_14265,N_14210,N_14248);
or U14266 (N_14266,N_14230,N_14163);
or U14267 (N_14267,N_14138,N_14176);
xnor U14268 (N_14268,N_14128,N_14167);
or U14269 (N_14269,N_14198,N_14125);
or U14270 (N_14270,N_14194,N_14211);
nor U14271 (N_14271,N_14170,N_14127);
nor U14272 (N_14272,N_14183,N_14247);
and U14273 (N_14273,N_14212,N_14142);
xor U14274 (N_14274,N_14168,N_14219);
nor U14275 (N_14275,N_14179,N_14145);
nor U14276 (N_14276,N_14156,N_14238);
xor U14277 (N_14277,N_14144,N_14186);
or U14278 (N_14278,N_14215,N_14188);
nor U14279 (N_14279,N_14207,N_14190);
or U14280 (N_14280,N_14139,N_14246);
nand U14281 (N_14281,N_14249,N_14187);
nor U14282 (N_14282,N_14209,N_14178);
nand U14283 (N_14283,N_14243,N_14239);
nor U14284 (N_14284,N_14182,N_14140);
xor U14285 (N_14285,N_14237,N_14224);
xor U14286 (N_14286,N_14203,N_14158);
xnor U14287 (N_14287,N_14228,N_14196);
and U14288 (N_14288,N_14204,N_14172);
xor U14289 (N_14289,N_14126,N_14137);
and U14290 (N_14290,N_14205,N_14199);
nor U14291 (N_14291,N_14218,N_14136);
and U14292 (N_14292,N_14143,N_14232);
and U14293 (N_14293,N_14201,N_14160);
xnor U14294 (N_14294,N_14223,N_14149);
nand U14295 (N_14295,N_14225,N_14150);
xnor U14296 (N_14296,N_14157,N_14151);
xor U14297 (N_14297,N_14241,N_14130);
xnor U14298 (N_14298,N_14222,N_14191);
nand U14299 (N_14299,N_14197,N_14174);
or U14300 (N_14300,N_14240,N_14177);
or U14301 (N_14301,N_14227,N_14129);
nand U14302 (N_14302,N_14216,N_14200);
xnor U14303 (N_14303,N_14153,N_14173);
xor U14304 (N_14304,N_14206,N_14242);
or U14305 (N_14305,N_14141,N_14192);
xnor U14306 (N_14306,N_14131,N_14202);
or U14307 (N_14307,N_14236,N_14213);
nor U14308 (N_14308,N_14214,N_14185);
nand U14309 (N_14309,N_14166,N_14234);
xnor U14310 (N_14310,N_14226,N_14132);
nor U14311 (N_14311,N_14184,N_14244);
nor U14312 (N_14312,N_14195,N_14216);
and U14313 (N_14313,N_14135,N_14198);
or U14314 (N_14314,N_14134,N_14178);
and U14315 (N_14315,N_14131,N_14184);
nor U14316 (N_14316,N_14244,N_14147);
nor U14317 (N_14317,N_14230,N_14245);
and U14318 (N_14318,N_14128,N_14174);
or U14319 (N_14319,N_14218,N_14169);
nor U14320 (N_14320,N_14225,N_14148);
or U14321 (N_14321,N_14241,N_14185);
and U14322 (N_14322,N_14151,N_14163);
xor U14323 (N_14323,N_14243,N_14202);
nor U14324 (N_14324,N_14204,N_14219);
and U14325 (N_14325,N_14172,N_14235);
or U14326 (N_14326,N_14198,N_14206);
or U14327 (N_14327,N_14228,N_14150);
nand U14328 (N_14328,N_14151,N_14126);
or U14329 (N_14329,N_14238,N_14215);
and U14330 (N_14330,N_14137,N_14144);
and U14331 (N_14331,N_14138,N_14175);
and U14332 (N_14332,N_14146,N_14200);
or U14333 (N_14333,N_14148,N_14176);
nand U14334 (N_14334,N_14203,N_14141);
and U14335 (N_14335,N_14227,N_14177);
nand U14336 (N_14336,N_14184,N_14219);
nand U14337 (N_14337,N_14185,N_14136);
nor U14338 (N_14338,N_14169,N_14177);
xor U14339 (N_14339,N_14213,N_14148);
or U14340 (N_14340,N_14192,N_14187);
or U14341 (N_14341,N_14214,N_14206);
nor U14342 (N_14342,N_14181,N_14166);
nand U14343 (N_14343,N_14203,N_14137);
and U14344 (N_14344,N_14202,N_14167);
or U14345 (N_14345,N_14171,N_14199);
xor U14346 (N_14346,N_14214,N_14141);
or U14347 (N_14347,N_14128,N_14180);
nor U14348 (N_14348,N_14244,N_14203);
or U14349 (N_14349,N_14243,N_14181);
nor U14350 (N_14350,N_14171,N_14249);
nor U14351 (N_14351,N_14195,N_14139);
nor U14352 (N_14352,N_14152,N_14214);
nor U14353 (N_14353,N_14223,N_14221);
nand U14354 (N_14354,N_14194,N_14126);
xnor U14355 (N_14355,N_14207,N_14131);
xor U14356 (N_14356,N_14164,N_14206);
and U14357 (N_14357,N_14161,N_14175);
or U14358 (N_14358,N_14196,N_14149);
nand U14359 (N_14359,N_14166,N_14223);
and U14360 (N_14360,N_14209,N_14190);
nand U14361 (N_14361,N_14200,N_14229);
or U14362 (N_14362,N_14160,N_14156);
or U14363 (N_14363,N_14147,N_14158);
nand U14364 (N_14364,N_14195,N_14226);
nor U14365 (N_14365,N_14136,N_14132);
or U14366 (N_14366,N_14143,N_14239);
or U14367 (N_14367,N_14125,N_14234);
nand U14368 (N_14368,N_14200,N_14130);
nand U14369 (N_14369,N_14198,N_14230);
xor U14370 (N_14370,N_14174,N_14230);
and U14371 (N_14371,N_14136,N_14165);
nand U14372 (N_14372,N_14233,N_14192);
xor U14373 (N_14373,N_14182,N_14215);
and U14374 (N_14374,N_14150,N_14126);
or U14375 (N_14375,N_14278,N_14366);
xnor U14376 (N_14376,N_14303,N_14318);
xor U14377 (N_14377,N_14307,N_14285);
nand U14378 (N_14378,N_14299,N_14257);
xor U14379 (N_14379,N_14309,N_14340);
and U14380 (N_14380,N_14357,N_14300);
xor U14381 (N_14381,N_14323,N_14283);
and U14382 (N_14382,N_14273,N_14296);
nand U14383 (N_14383,N_14369,N_14253);
and U14384 (N_14384,N_14325,N_14353);
xor U14385 (N_14385,N_14356,N_14343);
nor U14386 (N_14386,N_14327,N_14295);
nor U14387 (N_14387,N_14279,N_14364);
nor U14388 (N_14388,N_14328,N_14294);
nor U14389 (N_14389,N_14312,N_14267);
nor U14390 (N_14390,N_14305,N_14250);
and U14391 (N_14391,N_14321,N_14341);
xor U14392 (N_14392,N_14320,N_14298);
xor U14393 (N_14393,N_14311,N_14284);
nor U14394 (N_14394,N_14282,N_14254);
nand U14395 (N_14395,N_14308,N_14349);
or U14396 (N_14396,N_14251,N_14301);
or U14397 (N_14397,N_14332,N_14330);
nand U14398 (N_14398,N_14261,N_14265);
nand U14399 (N_14399,N_14293,N_14339);
nand U14400 (N_14400,N_14324,N_14331);
and U14401 (N_14401,N_14276,N_14350);
nand U14402 (N_14402,N_14262,N_14362);
nor U14403 (N_14403,N_14270,N_14316);
nor U14404 (N_14404,N_14337,N_14352);
nor U14405 (N_14405,N_14292,N_14342);
and U14406 (N_14406,N_14304,N_14368);
nor U14407 (N_14407,N_14260,N_14302);
or U14408 (N_14408,N_14329,N_14358);
or U14409 (N_14409,N_14346,N_14334);
and U14410 (N_14410,N_14288,N_14286);
nor U14411 (N_14411,N_14373,N_14313);
nor U14412 (N_14412,N_14345,N_14363);
nand U14413 (N_14413,N_14354,N_14347);
xor U14414 (N_14414,N_14370,N_14322);
and U14415 (N_14415,N_14289,N_14319);
nor U14416 (N_14416,N_14372,N_14367);
and U14417 (N_14417,N_14315,N_14255);
nor U14418 (N_14418,N_14266,N_14271);
xnor U14419 (N_14419,N_14335,N_14336);
nor U14420 (N_14420,N_14264,N_14361);
and U14421 (N_14421,N_14277,N_14281);
or U14422 (N_14422,N_14287,N_14274);
nor U14423 (N_14423,N_14259,N_14338);
xnor U14424 (N_14424,N_14310,N_14371);
or U14425 (N_14425,N_14280,N_14290);
and U14426 (N_14426,N_14317,N_14351);
nor U14427 (N_14427,N_14374,N_14297);
nand U14428 (N_14428,N_14344,N_14326);
or U14429 (N_14429,N_14268,N_14359);
nor U14430 (N_14430,N_14269,N_14333);
nor U14431 (N_14431,N_14258,N_14252);
xor U14432 (N_14432,N_14256,N_14360);
xnor U14433 (N_14433,N_14306,N_14348);
nor U14434 (N_14434,N_14355,N_14275);
and U14435 (N_14435,N_14263,N_14314);
nor U14436 (N_14436,N_14291,N_14365);
nor U14437 (N_14437,N_14272,N_14309);
xnor U14438 (N_14438,N_14277,N_14327);
xnor U14439 (N_14439,N_14371,N_14327);
xor U14440 (N_14440,N_14344,N_14295);
or U14441 (N_14441,N_14312,N_14347);
xor U14442 (N_14442,N_14296,N_14314);
xor U14443 (N_14443,N_14321,N_14283);
xor U14444 (N_14444,N_14325,N_14254);
nor U14445 (N_14445,N_14318,N_14280);
nor U14446 (N_14446,N_14312,N_14357);
nand U14447 (N_14447,N_14365,N_14278);
or U14448 (N_14448,N_14366,N_14255);
xnor U14449 (N_14449,N_14372,N_14365);
nor U14450 (N_14450,N_14371,N_14276);
nand U14451 (N_14451,N_14271,N_14366);
xnor U14452 (N_14452,N_14360,N_14329);
xor U14453 (N_14453,N_14277,N_14352);
and U14454 (N_14454,N_14258,N_14286);
xnor U14455 (N_14455,N_14305,N_14331);
nor U14456 (N_14456,N_14309,N_14286);
nand U14457 (N_14457,N_14329,N_14335);
nand U14458 (N_14458,N_14284,N_14329);
nor U14459 (N_14459,N_14339,N_14367);
or U14460 (N_14460,N_14328,N_14275);
nand U14461 (N_14461,N_14329,N_14314);
or U14462 (N_14462,N_14367,N_14362);
and U14463 (N_14463,N_14312,N_14371);
nand U14464 (N_14464,N_14359,N_14295);
xor U14465 (N_14465,N_14316,N_14279);
xor U14466 (N_14466,N_14337,N_14289);
nor U14467 (N_14467,N_14271,N_14340);
nand U14468 (N_14468,N_14312,N_14296);
and U14469 (N_14469,N_14250,N_14365);
nor U14470 (N_14470,N_14296,N_14264);
and U14471 (N_14471,N_14334,N_14287);
and U14472 (N_14472,N_14308,N_14327);
and U14473 (N_14473,N_14325,N_14345);
xnor U14474 (N_14474,N_14316,N_14333);
or U14475 (N_14475,N_14258,N_14277);
xnor U14476 (N_14476,N_14262,N_14346);
xor U14477 (N_14477,N_14261,N_14345);
and U14478 (N_14478,N_14355,N_14318);
nand U14479 (N_14479,N_14348,N_14324);
nand U14480 (N_14480,N_14320,N_14307);
or U14481 (N_14481,N_14274,N_14313);
or U14482 (N_14482,N_14295,N_14316);
and U14483 (N_14483,N_14336,N_14339);
nor U14484 (N_14484,N_14348,N_14288);
and U14485 (N_14485,N_14304,N_14312);
nand U14486 (N_14486,N_14373,N_14360);
nor U14487 (N_14487,N_14286,N_14266);
xor U14488 (N_14488,N_14364,N_14304);
nand U14489 (N_14489,N_14317,N_14252);
or U14490 (N_14490,N_14353,N_14348);
xnor U14491 (N_14491,N_14260,N_14307);
nand U14492 (N_14492,N_14357,N_14353);
nor U14493 (N_14493,N_14351,N_14275);
nand U14494 (N_14494,N_14374,N_14306);
xor U14495 (N_14495,N_14367,N_14297);
nor U14496 (N_14496,N_14299,N_14365);
or U14497 (N_14497,N_14330,N_14284);
and U14498 (N_14498,N_14336,N_14331);
nand U14499 (N_14499,N_14360,N_14270);
nand U14500 (N_14500,N_14382,N_14468);
nor U14501 (N_14501,N_14440,N_14448);
xor U14502 (N_14502,N_14447,N_14484);
nor U14503 (N_14503,N_14390,N_14455);
and U14504 (N_14504,N_14460,N_14472);
nor U14505 (N_14505,N_14437,N_14419);
xor U14506 (N_14506,N_14497,N_14463);
xnor U14507 (N_14507,N_14477,N_14425);
or U14508 (N_14508,N_14422,N_14397);
nand U14509 (N_14509,N_14404,N_14485);
nand U14510 (N_14510,N_14409,N_14471);
nand U14511 (N_14511,N_14436,N_14462);
or U14512 (N_14512,N_14491,N_14439);
and U14513 (N_14513,N_14389,N_14433);
nand U14514 (N_14514,N_14407,N_14413);
nor U14515 (N_14515,N_14495,N_14399);
and U14516 (N_14516,N_14454,N_14481);
nor U14517 (N_14517,N_14416,N_14391);
nor U14518 (N_14518,N_14476,N_14446);
and U14519 (N_14519,N_14381,N_14378);
xnor U14520 (N_14520,N_14469,N_14392);
xor U14521 (N_14521,N_14421,N_14443);
nor U14522 (N_14522,N_14499,N_14474);
xor U14523 (N_14523,N_14429,N_14478);
or U14524 (N_14524,N_14492,N_14426);
nor U14525 (N_14525,N_14475,N_14435);
nand U14526 (N_14526,N_14490,N_14375);
nand U14527 (N_14527,N_14438,N_14459);
xnor U14528 (N_14528,N_14482,N_14398);
and U14529 (N_14529,N_14445,N_14417);
and U14530 (N_14530,N_14431,N_14418);
xnor U14531 (N_14531,N_14387,N_14414);
nand U14532 (N_14532,N_14386,N_14449);
nor U14533 (N_14533,N_14470,N_14383);
or U14534 (N_14534,N_14408,N_14467);
or U14535 (N_14535,N_14376,N_14496);
nand U14536 (N_14536,N_14479,N_14379);
nand U14537 (N_14537,N_14450,N_14430);
xnor U14538 (N_14538,N_14424,N_14466);
nor U14539 (N_14539,N_14406,N_14458);
nand U14540 (N_14540,N_14452,N_14488);
and U14541 (N_14541,N_14453,N_14410);
or U14542 (N_14542,N_14464,N_14394);
or U14543 (N_14543,N_14480,N_14451);
nand U14544 (N_14544,N_14380,N_14427);
or U14545 (N_14545,N_14411,N_14395);
or U14546 (N_14546,N_14400,N_14402);
and U14547 (N_14547,N_14423,N_14415);
nor U14548 (N_14548,N_14456,N_14405);
or U14549 (N_14549,N_14384,N_14494);
or U14550 (N_14550,N_14498,N_14444);
nand U14551 (N_14551,N_14396,N_14442);
or U14552 (N_14552,N_14432,N_14428);
xnor U14553 (N_14553,N_14473,N_14486);
nand U14554 (N_14554,N_14487,N_14483);
xor U14555 (N_14555,N_14403,N_14388);
xnor U14556 (N_14556,N_14401,N_14465);
and U14557 (N_14557,N_14461,N_14377);
nor U14558 (N_14558,N_14420,N_14385);
nand U14559 (N_14559,N_14493,N_14489);
nor U14560 (N_14560,N_14457,N_14412);
xnor U14561 (N_14561,N_14393,N_14434);
nor U14562 (N_14562,N_14441,N_14488);
nand U14563 (N_14563,N_14376,N_14375);
xor U14564 (N_14564,N_14450,N_14451);
nand U14565 (N_14565,N_14450,N_14498);
or U14566 (N_14566,N_14489,N_14396);
xnor U14567 (N_14567,N_14396,N_14449);
nand U14568 (N_14568,N_14402,N_14493);
nor U14569 (N_14569,N_14474,N_14475);
xor U14570 (N_14570,N_14439,N_14400);
or U14571 (N_14571,N_14377,N_14491);
xor U14572 (N_14572,N_14473,N_14419);
nor U14573 (N_14573,N_14449,N_14423);
nor U14574 (N_14574,N_14496,N_14405);
nand U14575 (N_14575,N_14446,N_14477);
nand U14576 (N_14576,N_14467,N_14496);
nand U14577 (N_14577,N_14449,N_14439);
and U14578 (N_14578,N_14499,N_14490);
or U14579 (N_14579,N_14468,N_14449);
or U14580 (N_14580,N_14400,N_14424);
or U14581 (N_14581,N_14483,N_14385);
nand U14582 (N_14582,N_14416,N_14400);
or U14583 (N_14583,N_14429,N_14418);
nand U14584 (N_14584,N_14384,N_14444);
xor U14585 (N_14585,N_14494,N_14427);
nand U14586 (N_14586,N_14439,N_14437);
nand U14587 (N_14587,N_14450,N_14434);
nand U14588 (N_14588,N_14407,N_14408);
nand U14589 (N_14589,N_14494,N_14402);
or U14590 (N_14590,N_14442,N_14375);
or U14591 (N_14591,N_14469,N_14379);
nand U14592 (N_14592,N_14444,N_14450);
xor U14593 (N_14593,N_14472,N_14453);
or U14594 (N_14594,N_14464,N_14412);
or U14595 (N_14595,N_14404,N_14426);
xor U14596 (N_14596,N_14385,N_14379);
nor U14597 (N_14597,N_14467,N_14441);
or U14598 (N_14598,N_14442,N_14422);
or U14599 (N_14599,N_14412,N_14401);
xnor U14600 (N_14600,N_14434,N_14403);
nor U14601 (N_14601,N_14384,N_14455);
and U14602 (N_14602,N_14438,N_14429);
xnor U14603 (N_14603,N_14497,N_14481);
nand U14604 (N_14604,N_14443,N_14468);
nand U14605 (N_14605,N_14492,N_14413);
nand U14606 (N_14606,N_14400,N_14442);
nor U14607 (N_14607,N_14382,N_14399);
and U14608 (N_14608,N_14494,N_14438);
xor U14609 (N_14609,N_14492,N_14396);
xor U14610 (N_14610,N_14391,N_14433);
xor U14611 (N_14611,N_14387,N_14397);
xnor U14612 (N_14612,N_14464,N_14442);
and U14613 (N_14613,N_14389,N_14466);
and U14614 (N_14614,N_14476,N_14475);
nand U14615 (N_14615,N_14394,N_14442);
and U14616 (N_14616,N_14376,N_14469);
nand U14617 (N_14617,N_14447,N_14392);
nand U14618 (N_14618,N_14421,N_14462);
or U14619 (N_14619,N_14381,N_14450);
nand U14620 (N_14620,N_14405,N_14435);
and U14621 (N_14621,N_14474,N_14409);
nand U14622 (N_14622,N_14392,N_14423);
nand U14623 (N_14623,N_14488,N_14389);
nor U14624 (N_14624,N_14469,N_14486);
or U14625 (N_14625,N_14516,N_14609);
xor U14626 (N_14626,N_14536,N_14549);
xnor U14627 (N_14627,N_14573,N_14596);
nand U14628 (N_14628,N_14502,N_14515);
nor U14629 (N_14629,N_14531,N_14575);
xnor U14630 (N_14630,N_14509,N_14558);
or U14631 (N_14631,N_14508,N_14519);
and U14632 (N_14632,N_14544,N_14597);
nand U14633 (N_14633,N_14576,N_14538);
nor U14634 (N_14634,N_14605,N_14535);
nor U14635 (N_14635,N_14512,N_14557);
or U14636 (N_14636,N_14503,N_14584);
nand U14637 (N_14637,N_14624,N_14591);
and U14638 (N_14638,N_14618,N_14540);
nand U14639 (N_14639,N_14530,N_14615);
xor U14640 (N_14640,N_14532,N_14563);
nor U14641 (N_14641,N_14553,N_14548);
xnor U14642 (N_14642,N_14552,N_14613);
xor U14643 (N_14643,N_14599,N_14518);
and U14644 (N_14644,N_14565,N_14507);
nor U14645 (N_14645,N_14537,N_14547);
nand U14646 (N_14646,N_14510,N_14529);
or U14647 (N_14647,N_14526,N_14579);
or U14648 (N_14648,N_14586,N_14587);
xor U14649 (N_14649,N_14539,N_14566);
xor U14650 (N_14650,N_14550,N_14585);
nor U14651 (N_14651,N_14501,N_14595);
nand U14652 (N_14652,N_14520,N_14589);
nor U14653 (N_14653,N_14574,N_14580);
nand U14654 (N_14654,N_14524,N_14623);
xnor U14655 (N_14655,N_14546,N_14522);
xnor U14656 (N_14656,N_14582,N_14600);
xor U14657 (N_14657,N_14578,N_14594);
nand U14658 (N_14658,N_14543,N_14621);
nand U14659 (N_14659,N_14533,N_14617);
and U14660 (N_14660,N_14504,N_14592);
and U14661 (N_14661,N_14588,N_14608);
nor U14662 (N_14662,N_14568,N_14523);
nand U14663 (N_14663,N_14572,N_14567);
or U14664 (N_14664,N_14561,N_14593);
nand U14665 (N_14665,N_14556,N_14542);
and U14666 (N_14666,N_14581,N_14577);
nand U14667 (N_14667,N_14521,N_14564);
xnor U14668 (N_14668,N_14500,N_14554);
xor U14669 (N_14669,N_14607,N_14506);
and U14670 (N_14670,N_14611,N_14569);
or U14671 (N_14671,N_14620,N_14555);
and U14672 (N_14672,N_14527,N_14562);
or U14673 (N_14673,N_14602,N_14511);
or U14674 (N_14674,N_14570,N_14606);
xor U14675 (N_14675,N_14517,N_14622);
nand U14676 (N_14676,N_14603,N_14534);
xor U14677 (N_14677,N_14559,N_14505);
nand U14678 (N_14678,N_14590,N_14583);
or U14679 (N_14679,N_14601,N_14513);
and U14680 (N_14680,N_14560,N_14598);
nand U14681 (N_14681,N_14528,N_14616);
xnor U14682 (N_14682,N_14545,N_14610);
or U14683 (N_14683,N_14541,N_14571);
or U14684 (N_14684,N_14614,N_14514);
xor U14685 (N_14685,N_14604,N_14551);
and U14686 (N_14686,N_14525,N_14619);
nor U14687 (N_14687,N_14612,N_14538);
nand U14688 (N_14688,N_14563,N_14605);
and U14689 (N_14689,N_14552,N_14556);
nand U14690 (N_14690,N_14533,N_14569);
or U14691 (N_14691,N_14519,N_14517);
and U14692 (N_14692,N_14577,N_14621);
and U14693 (N_14693,N_14586,N_14541);
and U14694 (N_14694,N_14535,N_14537);
or U14695 (N_14695,N_14597,N_14535);
nor U14696 (N_14696,N_14549,N_14554);
nand U14697 (N_14697,N_14523,N_14532);
nand U14698 (N_14698,N_14542,N_14604);
xor U14699 (N_14699,N_14520,N_14533);
nor U14700 (N_14700,N_14507,N_14501);
xnor U14701 (N_14701,N_14531,N_14550);
and U14702 (N_14702,N_14623,N_14609);
nand U14703 (N_14703,N_14555,N_14507);
and U14704 (N_14704,N_14567,N_14544);
nor U14705 (N_14705,N_14558,N_14575);
xnor U14706 (N_14706,N_14591,N_14501);
nand U14707 (N_14707,N_14545,N_14552);
or U14708 (N_14708,N_14560,N_14519);
nand U14709 (N_14709,N_14593,N_14551);
nor U14710 (N_14710,N_14606,N_14507);
nor U14711 (N_14711,N_14568,N_14574);
or U14712 (N_14712,N_14595,N_14523);
xnor U14713 (N_14713,N_14513,N_14580);
xnor U14714 (N_14714,N_14588,N_14507);
nand U14715 (N_14715,N_14598,N_14507);
and U14716 (N_14716,N_14502,N_14532);
or U14717 (N_14717,N_14564,N_14538);
xnor U14718 (N_14718,N_14599,N_14577);
nor U14719 (N_14719,N_14520,N_14515);
or U14720 (N_14720,N_14586,N_14520);
nand U14721 (N_14721,N_14563,N_14561);
or U14722 (N_14722,N_14540,N_14550);
and U14723 (N_14723,N_14531,N_14527);
and U14724 (N_14724,N_14518,N_14591);
xnor U14725 (N_14725,N_14531,N_14602);
xor U14726 (N_14726,N_14528,N_14506);
and U14727 (N_14727,N_14621,N_14541);
or U14728 (N_14728,N_14585,N_14584);
nand U14729 (N_14729,N_14575,N_14609);
or U14730 (N_14730,N_14522,N_14601);
xnor U14731 (N_14731,N_14554,N_14526);
xnor U14732 (N_14732,N_14571,N_14614);
xnor U14733 (N_14733,N_14581,N_14572);
xnor U14734 (N_14734,N_14590,N_14527);
xnor U14735 (N_14735,N_14518,N_14605);
nand U14736 (N_14736,N_14512,N_14556);
or U14737 (N_14737,N_14507,N_14537);
xor U14738 (N_14738,N_14592,N_14565);
nand U14739 (N_14739,N_14515,N_14522);
or U14740 (N_14740,N_14533,N_14535);
xnor U14741 (N_14741,N_14617,N_14525);
nor U14742 (N_14742,N_14571,N_14518);
or U14743 (N_14743,N_14535,N_14509);
xor U14744 (N_14744,N_14611,N_14516);
and U14745 (N_14745,N_14605,N_14615);
nand U14746 (N_14746,N_14621,N_14518);
and U14747 (N_14747,N_14586,N_14610);
nand U14748 (N_14748,N_14594,N_14558);
nand U14749 (N_14749,N_14514,N_14538);
and U14750 (N_14750,N_14646,N_14721);
and U14751 (N_14751,N_14720,N_14713);
and U14752 (N_14752,N_14676,N_14649);
nor U14753 (N_14753,N_14673,N_14662);
nand U14754 (N_14754,N_14664,N_14727);
xnor U14755 (N_14755,N_14719,N_14654);
and U14756 (N_14756,N_14670,N_14647);
and U14757 (N_14757,N_14740,N_14667);
or U14758 (N_14758,N_14660,N_14688);
or U14759 (N_14759,N_14640,N_14637);
nor U14760 (N_14760,N_14674,N_14703);
nand U14761 (N_14761,N_14745,N_14635);
nand U14762 (N_14762,N_14716,N_14735);
and U14763 (N_14763,N_14630,N_14632);
or U14764 (N_14764,N_14734,N_14651);
xnor U14765 (N_14765,N_14747,N_14691);
or U14766 (N_14766,N_14728,N_14636);
nand U14767 (N_14767,N_14661,N_14685);
xor U14768 (N_14768,N_14733,N_14628);
nand U14769 (N_14769,N_14665,N_14711);
or U14770 (N_14770,N_14653,N_14631);
and U14771 (N_14771,N_14710,N_14723);
and U14772 (N_14772,N_14706,N_14705);
xnor U14773 (N_14773,N_14668,N_14741);
and U14774 (N_14774,N_14749,N_14736);
xor U14775 (N_14775,N_14701,N_14678);
or U14776 (N_14776,N_14677,N_14642);
nand U14777 (N_14777,N_14700,N_14644);
nor U14778 (N_14778,N_14726,N_14690);
xor U14779 (N_14779,N_14657,N_14658);
nor U14780 (N_14780,N_14655,N_14626);
or U14781 (N_14781,N_14717,N_14748);
nor U14782 (N_14782,N_14702,N_14675);
nand U14783 (N_14783,N_14729,N_14722);
and U14784 (N_14784,N_14639,N_14712);
nor U14785 (N_14785,N_14724,N_14744);
nand U14786 (N_14786,N_14696,N_14718);
xnor U14787 (N_14787,N_14679,N_14694);
xor U14788 (N_14788,N_14669,N_14743);
or U14789 (N_14789,N_14687,N_14629);
nor U14790 (N_14790,N_14697,N_14725);
and U14791 (N_14791,N_14709,N_14693);
nor U14792 (N_14792,N_14641,N_14689);
xnor U14793 (N_14793,N_14738,N_14732);
nor U14794 (N_14794,N_14682,N_14683);
nor U14795 (N_14795,N_14731,N_14714);
nor U14796 (N_14796,N_14730,N_14680);
xor U14797 (N_14797,N_14739,N_14698);
nand U14798 (N_14798,N_14684,N_14704);
or U14799 (N_14799,N_14707,N_14746);
or U14800 (N_14800,N_14659,N_14692);
and U14801 (N_14801,N_14652,N_14663);
nor U14802 (N_14802,N_14708,N_14648);
or U14803 (N_14803,N_14645,N_14643);
nor U14804 (N_14804,N_14742,N_14686);
and U14805 (N_14805,N_14715,N_14699);
xor U14806 (N_14806,N_14625,N_14672);
nand U14807 (N_14807,N_14671,N_14737);
nor U14808 (N_14808,N_14650,N_14666);
or U14809 (N_14809,N_14656,N_14627);
nor U14810 (N_14810,N_14638,N_14633);
nand U14811 (N_14811,N_14695,N_14681);
nor U14812 (N_14812,N_14634,N_14683);
nand U14813 (N_14813,N_14700,N_14698);
or U14814 (N_14814,N_14688,N_14730);
or U14815 (N_14815,N_14655,N_14695);
xor U14816 (N_14816,N_14733,N_14706);
or U14817 (N_14817,N_14671,N_14655);
nor U14818 (N_14818,N_14739,N_14637);
xnor U14819 (N_14819,N_14699,N_14660);
or U14820 (N_14820,N_14725,N_14691);
nand U14821 (N_14821,N_14644,N_14745);
and U14822 (N_14822,N_14679,N_14710);
nor U14823 (N_14823,N_14699,N_14680);
and U14824 (N_14824,N_14666,N_14674);
or U14825 (N_14825,N_14677,N_14690);
nand U14826 (N_14826,N_14692,N_14670);
and U14827 (N_14827,N_14722,N_14674);
xnor U14828 (N_14828,N_14694,N_14699);
nand U14829 (N_14829,N_14743,N_14699);
or U14830 (N_14830,N_14746,N_14718);
or U14831 (N_14831,N_14648,N_14625);
nor U14832 (N_14832,N_14706,N_14730);
and U14833 (N_14833,N_14638,N_14746);
nor U14834 (N_14834,N_14709,N_14715);
and U14835 (N_14835,N_14640,N_14665);
or U14836 (N_14836,N_14684,N_14639);
and U14837 (N_14837,N_14710,N_14689);
xnor U14838 (N_14838,N_14649,N_14704);
xnor U14839 (N_14839,N_14716,N_14666);
and U14840 (N_14840,N_14723,N_14709);
and U14841 (N_14841,N_14712,N_14744);
nor U14842 (N_14842,N_14689,N_14672);
nand U14843 (N_14843,N_14668,N_14645);
or U14844 (N_14844,N_14719,N_14708);
and U14845 (N_14845,N_14626,N_14734);
or U14846 (N_14846,N_14730,N_14711);
xor U14847 (N_14847,N_14693,N_14630);
or U14848 (N_14848,N_14744,N_14697);
nor U14849 (N_14849,N_14727,N_14659);
or U14850 (N_14850,N_14712,N_14693);
xor U14851 (N_14851,N_14718,N_14745);
xor U14852 (N_14852,N_14667,N_14668);
or U14853 (N_14853,N_14733,N_14643);
or U14854 (N_14854,N_14681,N_14721);
or U14855 (N_14855,N_14648,N_14722);
nand U14856 (N_14856,N_14735,N_14731);
xor U14857 (N_14857,N_14711,N_14678);
xor U14858 (N_14858,N_14638,N_14738);
or U14859 (N_14859,N_14656,N_14715);
or U14860 (N_14860,N_14672,N_14734);
and U14861 (N_14861,N_14698,N_14665);
and U14862 (N_14862,N_14709,N_14637);
or U14863 (N_14863,N_14699,N_14730);
xor U14864 (N_14864,N_14654,N_14638);
or U14865 (N_14865,N_14696,N_14663);
xor U14866 (N_14866,N_14714,N_14628);
nor U14867 (N_14867,N_14677,N_14675);
nand U14868 (N_14868,N_14632,N_14703);
or U14869 (N_14869,N_14735,N_14665);
and U14870 (N_14870,N_14641,N_14733);
and U14871 (N_14871,N_14717,N_14730);
nand U14872 (N_14872,N_14687,N_14690);
and U14873 (N_14873,N_14633,N_14748);
or U14874 (N_14874,N_14726,N_14631);
nand U14875 (N_14875,N_14826,N_14813);
nor U14876 (N_14876,N_14789,N_14772);
and U14877 (N_14877,N_14816,N_14854);
or U14878 (N_14878,N_14869,N_14818);
nand U14879 (N_14879,N_14778,N_14868);
or U14880 (N_14880,N_14756,N_14837);
and U14881 (N_14881,N_14755,N_14757);
nand U14882 (N_14882,N_14862,N_14848);
and U14883 (N_14883,N_14773,N_14795);
nand U14884 (N_14884,N_14771,N_14804);
and U14885 (N_14885,N_14815,N_14836);
xor U14886 (N_14886,N_14841,N_14860);
xnor U14887 (N_14887,N_14794,N_14852);
and U14888 (N_14888,N_14865,N_14817);
or U14889 (N_14889,N_14845,N_14770);
nand U14890 (N_14890,N_14847,N_14825);
or U14891 (N_14891,N_14774,N_14751);
and U14892 (N_14892,N_14758,N_14874);
nand U14893 (N_14893,N_14827,N_14784);
and U14894 (N_14894,N_14839,N_14779);
nor U14895 (N_14895,N_14761,N_14792);
and U14896 (N_14896,N_14843,N_14796);
or U14897 (N_14897,N_14807,N_14793);
or U14898 (N_14898,N_14850,N_14803);
xnor U14899 (N_14899,N_14844,N_14859);
or U14900 (N_14900,N_14856,N_14863);
nor U14901 (N_14901,N_14753,N_14767);
or U14902 (N_14902,N_14763,N_14805);
or U14903 (N_14903,N_14840,N_14823);
and U14904 (N_14904,N_14800,N_14764);
or U14905 (N_14905,N_14821,N_14759);
or U14906 (N_14906,N_14754,N_14842);
and U14907 (N_14907,N_14783,N_14781);
and U14908 (N_14908,N_14812,N_14752);
nor U14909 (N_14909,N_14819,N_14785);
xor U14910 (N_14910,N_14824,N_14853);
and U14911 (N_14911,N_14806,N_14750);
and U14912 (N_14912,N_14765,N_14838);
and U14913 (N_14913,N_14799,N_14834);
nor U14914 (N_14914,N_14867,N_14801);
or U14915 (N_14915,N_14872,N_14762);
and U14916 (N_14916,N_14833,N_14855);
or U14917 (N_14917,N_14835,N_14766);
or U14918 (N_14918,N_14829,N_14851);
nand U14919 (N_14919,N_14846,N_14828);
and U14920 (N_14920,N_14861,N_14871);
nor U14921 (N_14921,N_14866,N_14788);
xor U14922 (N_14922,N_14870,N_14780);
xor U14923 (N_14923,N_14760,N_14808);
nor U14924 (N_14924,N_14791,N_14787);
nor U14925 (N_14925,N_14775,N_14802);
nor U14926 (N_14926,N_14831,N_14782);
or U14927 (N_14927,N_14809,N_14769);
nor U14928 (N_14928,N_14858,N_14864);
or U14929 (N_14929,N_14797,N_14790);
or U14930 (N_14930,N_14849,N_14873);
and U14931 (N_14931,N_14822,N_14830);
xnor U14932 (N_14932,N_14814,N_14776);
or U14933 (N_14933,N_14777,N_14810);
nor U14934 (N_14934,N_14857,N_14786);
or U14935 (N_14935,N_14768,N_14820);
xor U14936 (N_14936,N_14798,N_14811);
or U14937 (N_14937,N_14832,N_14783);
nand U14938 (N_14938,N_14829,N_14863);
nand U14939 (N_14939,N_14818,N_14801);
or U14940 (N_14940,N_14868,N_14848);
nand U14941 (N_14941,N_14795,N_14862);
or U14942 (N_14942,N_14819,N_14851);
nor U14943 (N_14943,N_14872,N_14796);
or U14944 (N_14944,N_14810,N_14785);
nor U14945 (N_14945,N_14771,N_14872);
nor U14946 (N_14946,N_14786,N_14768);
or U14947 (N_14947,N_14800,N_14763);
xnor U14948 (N_14948,N_14813,N_14786);
or U14949 (N_14949,N_14836,N_14785);
nor U14950 (N_14950,N_14779,N_14757);
and U14951 (N_14951,N_14769,N_14847);
nand U14952 (N_14952,N_14860,N_14805);
or U14953 (N_14953,N_14824,N_14820);
or U14954 (N_14954,N_14802,N_14830);
or U14955 (N_14955,N_14811,N_14773);
nor U14956 (N_14956,N_14818,N_14840);
xnor U14957 (N_14957,N_14846,N_14826);
nand U14958 (N_14958,N_14841,N_14791);
nand U14959 (N_14959,N_14791,N_14768);
and U14960 (N_14960,N_14758,N_14786);
nor U14961 (N_14961,N_14767,N_14795);
nor U14962 (N_14962,N_14758,N_14822);
and U14963 (N_14963,N_14783,N_14761);
xnor U14964 (N_14964,N_14860,N_14837);
and U14965 (N_14965,N_14759,N_14832);
nor U14966 (N_14966,N_14852,N_14853);
nand U14967 (N_14967,N_14825,N_14799);
xor U14968 (N_14968,N_14865,N_14819);
nor U14969 (N_14969,N_14801,N_14757);
nand U14970 (N_14970,N_14750,N_14867);
and U14971 (N_14971,N_14815,N_14781);
nor U14972 (N_14972,N_14832,N_14858);
xnor U14973 (N_14973,N_14794,N_14834);
nor U14974 (N_14974,N_14756,N_14758);
nor U14975 (N_14975,N_14861,N_14867);
nand U14976 (N_14976,N_14766,N_14753);
nor U14977 (N_14977,N_14857,N_14839);
or U14978 (N_14978,N_14826,N_14773);
or U14979 (N_14979,N_14782,N_14753);
and U14980 (N_14980,N_14840,N_14775);
and U14981 (N_14981,N_14856,N_14860);
xnor U14982 (N_14982,N_14805,N_14770);
or U14983 (N_14983,N_14797,N_14808);
and U14984 (N_14984,N_14756,N_14858);
nor U14985 (N_14985,N_14813,N_14830);
nand U14986 (N_14986,N_14790,N_14753);
nand U14987 (N_14987,N_14831,N_14774);
or U14988 (N_14988,N_14869,N_14751);
or U14989 (N_14989,N_14866,N_14828);
nor U14990 (N_14990,N_14856,N_14796);
and U14991 (N_14991,N_14781,N_14806);
and U14992 (N_14992,N_14781,N_14833);
nand U14993 (N_14993,N_14750,N_14752);
xnor U14994 (N_14994,N_14812,N_14824);
xnor U14995 (N_14995,N_14776,N_14849);
or U14996 (N_14996,N_14783,N_14790);
xnor U14997 (N_14997,N_14825,N_14774);
and U14998 (N_14998,N_14783,N_14777);
xnor U14999 (N_14999,N_14782,N_14809);
xnor UO_0 (O_0,N_14961,N_14951);
and UO_1 (O_1,N_14884,N_14907);
and UO_2 (O_2,N_14887,N_14941);
and UO_3 (O_3,N_14905,N_14964);
and UO_4 (O_4,N_14881,N_14962);
and UO_5 (O_5,N_14889,N_14918);
xnor UO_6 (O_6,N_14911,N_14926);
or UO_7 (O_7,N_14965,N_14935);
or UO_8 (O_8,N_14992,N_14921);
nand UO_9 (O_9,N_14909,N_14899);
or UO_10 (O_10,N_14966,N_14922);
nand UO_11 (O_11,N_14940,N_14981);
and UO_12 (O_12,N_14928,N_14927);
nand UO_13 (O_13,N_14897,N_14910);
or UO_14 (O_14,N_14925,N_14876);
nand UO_15 (O_15,N_14957,N_14950);
xnor UO_16 (O_16,N_14959,N_14980);
nor UO_17 (O_17,N_14877,N_14875);
xnor UO_18 (O_18,N_14947,N_14906);
nor UO_19 (O_19,N_14990,N_14985);
and UO_20 (O_20,N_14912,N_14879);
xor UO_21 (O_21,N_14969,N_14939);
nor UO_22 (O_22,N_14953,N_14920);
xor UO_23 (O_23,N_14898,N_14933);
or UO_24 (O_24,N_14930,N_14894);
xor UO_25 (O_25,N_14934,N_14937);
nand UO_26 (O_26,N_14914,N_14977);
xnor UO_27 (O_27,N_14942,N_14901);
and UO_28 (O_28,N_14916,N_14986);
xnor UO_29 (O_29,N_14956,N_14993);
xor UO_30 (O_30,N_14978,N_14974);
xor UO_31 (O_31,N_14924,N_14923);
nor UO_32 (O_32,N_14995,N_14919);
or UO_33 (O_33,N_14982,N_14900);
xnor UO_34 (O_34,N_14936,N_14896);
xnor UO_35 (O_35,N_14904,N_14952);
xnor UO_36 (O_36,N_14932,N_14878);
or UO_37 (O_37,N_14943,N_14958);
nand UO_38 (O_38,N_14979,N_14893);
and UO_39 (O_39,N_14996,N_14882);
xor UO_40 (O_40,N_14960,N_14967);
and UO_41 (O_41,N_14973,N_14915);
or UO_42 (O_42,N_14984,N_14970);
nor UO_43 (O_43,N_14948,N_14963);
or UO_44 (O_44,N_14908,N_14938);
nor UO_45 (O_45,N_14991,N_14968);
nand UO_46 (O_46,N_14903,N_14913);
nand UO_47 (O_47,N_14880,N_14917);
and UO_48 (O_48,N_14902,N_14987);
xor UO_49 (O_49,N_14994,N_14892);
nand UO_50 (O_50,N_14971,N_14954);
and UO_51 (O_51,N_14929,N_14989);
nand UO_52 (O_52,N_14955,N_14944);
nor UO_53 (O_53,N_14885,N_14988);
xor UO_54 (O_54,N_14886,N_14883);
xor UO_55 (O_55,N_14895,N_14949);
and UO_56 (O_56,N_14998,N_14997);
nor UO_57 (O_57,N_14946,N_14890);
xnor UO_58 (O_58,N_14999,N_14972);
nor UO_59 (O_59,N_14983,N_14976);
nand UO_60 (O_60,N_14975,N_14891);
nand UO_61 (O_61,N_14888,N_14945);
xnor UO_62 (O_62,N_14931,N_14984);
nand UO_63 (O_63,N_14963,N_14920);
nand UO_64 (O_64,N_14888,N_14876);
or UO_65 (O_65,N_14881,N_14928);
and UO_66 (O_66,N_14920,N_14921);
or UO_67 (O_67,N_14892,N_14979);
and UO_68 (O_68,N_14923,N_14943);
xnor UO_69 (O_69,N_14881,N_14884);
nand UO_70 (O_70,N_14899,N_14956);
or UO_71 (O_71,N_14914,N_14993);
nor UO_72 (O_72,N_14988,N_14960);
or UO_73 (O_73,N_14965,N_14962);
or UO_74 (O_74,N_14892,N_14950);
and UO_75 (O_75,N_14907,N_14995);
nand UO_76 (O_76,N_14908,N_14977);
nand UO_77 (O_77,N_14875,N_14882);
and UO_78 (O_78,N_14995,N_14938);
nor UO_79 (O_79,N_14944,N_14901);
and UO_80 (O_80,N_14951,N_14944);
or UO_81 (O_81,N_14885,N_14932);
nor UO_82 (O_82,N_14975,N_14896);
nor UO_83 (O_83,N_14938,N_14912);
nor UO_84 (O_84,N_14998,N_14924);
and UO_85 (O_85,N_14890,N_14945);
nor UO_86 (O_86,N_14934,N_14898);
or UO_87 (O_87,N_14973,N_14906);
and UO_88 (O_88,N_14969,N_14951);
nor UO_89 (O_89,N_14894,N_14968);
nand UO_90 (O_90,N_14925,N_14966);
or UO_91 (O_91,N_14878,N_14912);
nor UO_92 (O_92,N_14980,N_14969);
nand UO_93 (O_93,N_14958,N_14945);
or UO_94 (O_94,N_14973,N_14969);
and UO_95 (O_95,N_14974,N_14950);
or UO_96 (O_96,N_14914,N_14942);
nor UO_97 (O_97,N_14891,N_14993);
nor UO_98 (O_98,N_14927,N_14973);
nor UO_99 (O_99,N_14922,N_14884);
xnor UO_100 (O_100,N_14909,N_14908);
nor UO_101 (O_101,N_14935,N_14877);
or UO_102 (O_102,N_14986,N_14943);
and UO_103 (O_103,N_14986,N_14931);
nand UO_104 (O_104,N_14987,N_14970);
or UO_105 (O_105,N_14952,N_14982);
or UO_106 (O_106,N_14919,N_14877);
nor UO_107 (O_107,N_14986,N_14941);
nand UO_108 (O_108,N_14937,N_14968);
and UO_109 (O_109,N_14977,N_14956);
and UO_110 (O_110,N_14929,N_14990);
and UO_111 (O_111,N_14901,N_14986);
nor UO_112 (O_112,N_14969,N_14883);
or UO_113 (O_113,N_14879,N_14886);
nor UO_114 (O_114,N_14902,N_14942);
or UO_115 (O_115,N_14994,N_14886);
and UO_116 (O_116,N_14980,N_14987);
xor UO_117 (O_117,N_14949,N_14890);
nand UO_118 (O_118,N_14915,N_14893);
nor UO_119 (O_119,N_14936,N_14967);
nand UO_120 (O_120,N_14940,N_14943);
xnor UO_121 (O_121,N_14918,N_14901);
or UO_122 (O_122,N_14939,N_14961);
or UO_123 (O_123,N_14998,N_14973);
nand UO_124 (O_124,N_14971,N_14994);
or UO_125 (O_125,N_14958,N_14921);
xor UO_126 (O_126,N_14954,N_14948);
or UO_127 (O_127,N_14896,N_14951);
and UO_128 (O_128,N_14882,N_14951);
nand UO_129 (O_129,N_14888,N_14878);
or UO_130 (O_130,N_14955,N_14971);
nand UO_131 (O_131,N_14940,N_14925);
and UO_132 (O_132,N_14989,N_14980);
nor UO_133 (O_133,N_14966,N_14904);
xor UO_134 (O_134,N_14881,N_14956);
nand UO_135 (O_135,N_14909,N_14982);
xnor UO_136 (O_136,N_14946,N_14929);
or UO_137 (O_137,N_14883,N_14983);
xor UO_138 (O_138,N_14929,N_14963);
xor UO_139 (O_139,N_14946,N_14938);
nor UO_140 (O_140,N_14968,N_14884);
or UO_141 (O_141,N_14886,N_14964);
or UO_142 (O_142,N_14885,N_14912);
nand UO_143 (O_143,N_14923,N_14977);
or UO_144 (O_144,N_14988,N_14971);
nand UO_145 (O_145,N_14927,N_14968);
and UO_146 (O_146,N_14910,N_14997);
or UO_147 (O_147,N_14953,N_14996);
nor UO_148 (O_148,N_14881,N_14917);
xnor UO_149 (O_149,N_14960,N_14885);
nand UO_150 (O_150,N_14895,N_14990);
and UO_151 (O_151,N_14922,N_14959);
and UO_152 (O_152,N_14913,N_14968);
or UO_153 (O_153,N_14961,N_14885);
or UO_154 (O_154,N_14978,N_14890);
and UO_155 (O_155,N_14956,N_14984);
nand UO_156 (O_156,N_14924,N_14976);
nor UO_157 (O_157,N_14876,N_14933);
nor UO_158 (O_158,N_14945,N_14916);
and UO_159 (O_159,N_14887,N_14952);
and UO_160 (O_160,N_14899,N_14897);
nand UO_161 (O_161,N_14922,N_14891);
and UO_162 (O_162,N_14878,N_14970);
nor UO_163 (O_163,N_14944,N_14921);
and UO_164 (O_164,N_14897,N_14908);
nor UO_165 (O_165,N_14949,N_14919);
and UO_166 (O_166,N_14881,N_14919);
nand UO_167 (O_167,N_14910,N_14899);
nor UO_168 (O_168,N_14942,N_14935);
or UO_169 (O_169,N_14941,N_14961);
nor UO_170 (O_170,N_14962,N_14878);
nand UO_171 (O_171,N_14909,N_14931);
and UO_172 (O_172,N_14878,N_14928);
or UO_173 (O_173,N_14879,N_14913);
and UO_174 (O_174,N_14993,N_14937);
and UO_175 (O_175,N_14925,N_14898);
nor UO_176 (O_176,N_14938,N_14960);
nor UO_177 (O_177,N_14933,N_14999);
and UO_178 (O_178,N_14897,N_14998);
nand UO_179 (O_179,N_14968,N_14881);
xor UO_180 (O_180,N_14991,N_14920);
or UO_181 (O_181,N_14996,N_14965);
nand UO_182 (O_182,N_14875,N_14887);
nor UO_183 (O_183,N_14924,N_14880);
and UO_184 (O_184,N_14985,N_14890);
and UO_185 (O_185,N_14896,N_14923);
nand UO_186 (O_186,N_14920,N_14989);
and UO_187 (O_187,N_14906,N_14895);
xnor UO_188 (O_188,N_14940,N_14996);
nor UO_189 (O_189,N_14914,N_14897);
nor UO_190 (O_190,N_14900,N_14904);
nor UO_191 (O_191,N_14964,N_14919);
or UO_192 (O_192,N_14938,N_14930);
or UO_193 (O_193,N_14879,N_14946);
or UO_194 (O_194,N_14942,N_14947);
nand UO_195 (O_195,N_14968,N_14904);
and UO_196 (O_196,N_14875,N_14992);
nor UO_197 (O_197,N_14877,N_14948);
and UO_198 (O_198,N_14929,N_14914);
and UO_199 (O_199,N_14899,N_14962);
or UO_200 (O_200,N_14930,N_14959);
nor UO_201 (O_201,N_14910,N_14990);
nor UO_202 (O_202,N_14951,N_14940);
nor UO_203 (O_203,N_14972,N_14898);
and UO_204 (O_204,N_14901,N_14939);
nand UO_205 (O_205,N_14914,N_14999);
or UO_206 (O_206,N_14980,N_14902);
and UO_207 (O_207,N_14998,N_14910);
or UO_208 (O_208,N_14938,N_14881);
xor UO_209 (O_209,N_14895,N_14942);
nor UO_210 (O_210,N_14934,N_14976);
xor UO_211 (O_211,N_14998,N_14947);
xnor UO_212 (O_212,N_14880,N_14888);
xnor UO_213 (O_213,N_14910,N_14932);
and UO_214 (O_214,N_14992,N_14933);
nand UO_215 (O_215,N_14994,N_14962);
or UO_216 (O_216,N_14897,N_14993);
and UO_217 (O_217,N_14948,N_14956);
xnor UO_218 (O_218,N_14994,N_14914);
xor UO_219 (O_219,N_14904,N_14937);
nand UO_220 (O_220,N_14903,N_14952);
nor UO_221 (O_221,N_14978,N_14983);
and UO_222 (O_222,N_14959,N_14878);
xnor UO_223 (O_223,N_14951,N_14974);
xnor UO_224 (O_224,N_14909,N_14921);
xnor UO_225 (O_225,N_14961,N_14948);
nor UO_226 (O_226,N_14876,N_14975);
and UO_227 (O_227,N_14919,N_14968);
or UO_228 (O_228,N_14974,N_14967);
or UO_229 (O_229,N_14965,N_14955);
or UO_230 (O_230,N_14934,N_14971);
nand UO_231 (O_231,N_14917,N_14910);
nor UO_232 (O_232,N_14966,N_14930);
or UO_233 (O_233,N_14978,N_14884);
xnor UO_234 (O_234,N_14946,N_14987);
nor UO_235 (O_235,N_14961,N_14875);
nor UO_236 (O_236,N_14997,N_14945);
and UO_237 (O_237,N_14999,N_14973);
or UO_238 (O_238,N_14889,N_14878);
or UO_239 (O_239,N_14918,N_14958);
and UO_240 (O_240,N_14878,N_14995);
and UO_241 (O_241,N_14952,N_14917);
nand UO_242 (O_242,N_14954,N_14920);
nand UO_243 (O_243,N_14900,N_14875);
or UO_244 (O_244,N_14891,N_14941);
or UO_245 (O_245,N_14932,N_14980);
nor UO_246 (O_246,N_14946,N_14903);
and UO_247 (O_247,N_14888,N_14892);
or UO_248 (O_248,N_14895,N_14908);
nand UO_249 (O_249,N_14994,N_14993);
nor UO_250 (O_250,N_14975,N_14946);
or UO_251 (O_251,N_14881,N_14988);
and UO_252 (O_252,N_14877,N_14994);
and UO_253 (O_253,N_14892,N_14966);
nor UO_254 (O_254,N_14948,N_14929);
or UO_255 (O_255,N_14972,N_14976);
xnor UO_256 (O_256,N_14935,N_14914);
or UO_257 (O_257,N_14989,N_14982);
nor UO_258 (O_258,N_14912,N_14993);
or UO_259 (O_259,N_14889,N_14989);
nor UO_260 (O_260,N_14982,N_14902);
xnor UO_261 (O_261,N_14940,N_14887);
and UO_262 (O_262,N_14904,N_14940);
nand UO_263 (O_263,N_14881,N_14977);
and UO_264 (O_264,N_14879,N_14979);
or UO_265 (O_265,N_14997,N_14878);
xor UO_266 (O_266,N_14985,N_14883);
nor UO_267 (O_267,N_14879,N_14956);
nand UO_268 (O_268,N_14940,N_14988);
or UO_269 (O_269,N_14922,N_14941);
or UO_270 (O_270,N_14961,N_14947);
or UO_271 (O_271,N_14942,N_14887);
nand UO_272 (O_272,N_14992,N_14902);
xnor UO_273 (O_273,N_14968,N_14906);
nand UO_274 (O_274,N_14880,N_14875);
nor UO_275 (O_275,N_14923,N_14996);
and UO_276 (O_276,N_14979,N_14963);
and UO_277 (O_277,N_14947,N_14978);
nand UO_278 (O_278,N_14979,N_14877);
nand UO_279 (O_279,N_14908,N_14921);
or UO_280 (O_280,N_14965,N_14893);
xnor UO_281 (O_281,N_14882,N_14888);
nor UO_282 (O_282,N_14931,N_14903);
xnor UO_283 (O_283,N_14935,N_14943);
and UO_284 (O_284,N_14909,N_14974);
or UO_285 (O_285,N_14952,N_14971);
or UO_286 (O_286,N_14993,N_14992);
nand UO_287 (O_287,N_14992,N_14924);
and UO_288 (O_288,N_14976,N_14982);
or UO_289 (O_289,N_14927,N_14987);
or UO_290 (O_290,N_14890,N_14900);
nand UO_291 (O_291,N_14995,N_14924);
nor UO_292 (O_292,N_14946,N_14936);
or UO_293 (O_293,N_14923,N_14930);
nor UO_294 (O_294,N_14900,N_14882);
nand UO_295 (O_295,N_14987,N_14929);
or UO_296 (O_296,N_14885,N_14964);
or UO_297 (O_297,N_14882,N_14914);
nand UO_298 (O_298,N_14950,N_14982);
nand UO_299 (O_299,N_14876,N_14931);
xnor UO_300 (O_300,N_14990,N_14951);
xnor UO_301 (O_301,N_14971,N_14958);
nor UO_302 (O_302,N_14952,N_14882);
nor UO_303 (O_303,N_14880,N_14941);
or UO_304 (O_304,N_14968,N_14893);
nor UO_305 (O_305,N_14973,N_14995);
xnor UO_306 (O_306,N_14998,N_14999);
and UO_307 (O_307,N_14885,N_14927);
and UO_308 (O_308,N_14980,N_14979);
nor UO_309 (O_309,N_14936,N_14992);
xor UO_310 (O_310,N_14892,N_14881);
or UO_311 (O_311,N_14942,N_14944);
or UO_312 (O_312,N_14911,N_14882);
nor UO_313 (O_313,N_14986,N_14919);
or UO_314 (O_314,N_14948,N_14900);
nand UO_315 (O_315,N_14969,N_14916);
xor UO_316 (O_316,N_14912,N_14892);
and UO_317 (O_317,N_14910,N_14896);
and UO_318 (O_318,N_14879,N_14974);
or UO_319 (O_319,N_14897,N_14903);
and UO_320 (O_320,N_14982,N_14998);
nor UO_321 (O_321,N_14921,N_14970);
or UO_322 (O_322,N_14987,N_14925);
or UO_323 (O_323,N_14960,N_14981);
nand UO_324 (O_324,N_14947,N_14915);
and UO_325 (O_325,N_14903,N_14881);
nor UO_326 (O_326,N_14889,N_14945);
nor UO_327 (O_327,N_14940,N_14894);
nand UO_328 (O_328,N_14973,N_14981);
nor UO_329 (O_329,N_14930,N_14969);
nand UO_330 (O_330,N_14973,N_14889);
nand UO_331 (O_331,N_14960,N_14894);
nand UO_332 (O_332,N_14922,N_14978);
nand UO_333 (O_333,N_14887,N_14901);
and UO_334 (O_334,N_14956,N_14992);
nor UO_335 (O_335,N_14966,N_14895);
nor UO_336 (O_336,N_14898,N_14894);
xnor UO_337 (O_337,N_14903,N_14941);
or UO_338 (O_338,N_14985,N_14892);
and UO_339 (O_339,N_14910,N_14966);
or UO_340 (O_340,N_14919,N_14930);
and UO_341 (O_341,N_14997,N_14892);
nand UO_342 (O_342,N_14982,N_14875);
nor UO_343 (O_343,N_14899,N_14881);
nor UO_344 (O_344,N_14970,N_14998);
nor UO_345 (O_345,N_14999,N_14984);
nor UO_346 (O_346,N_14890,N_14911);
and UO_347 (O_347,N_14945,N_14923);
nand UO_348 (O_348,N_14968,N_14931);
nor UO_349 (O_349,N_14952,N_14991);
and UO_350 (O_350,N_14926,N_14995);
nand UO_351 (O_351,N_14984,N_14917);
or UO_352 (O_352,N_14989,N_14903);
or UO_353 (O_353,N_14987,N_14931);
nor UO_354 (O_354,N_14993,N_14962);
nor UO_355 (O_355,N_14950,N_14921);
or UO_356 (O_356,N_14958,N_14915);
xor UO_357 (O_357,N_14992,N_14961);
or UO_358 (O_358,N_14962,N_14887);
xnor UO_359 (O_359,N_14949,N_14979);
or UO_360 (O_360,N_14955,N_14995);
or UO_361 (O_361,N_14947,N_14982);
xor UO_362 (O_362,N_14936,N_14898);
and UO_363 (O_363,N_14990,N_14984);
nor UO_364 (O_364,N_14980,N_14930);
nand UO_365 (O_365,N_14950,N_14956);
or UO_366 (O_366,N_14995,N_14875);
and UO_367 (O_367,N_14957,N_14882);
xor UO_368 (O_368,N_14900,N_14888);
and UO_369 (O_369,N_14909,N_14993);
xor UO_370 (O_370,N_14878,N_14915);
or UO_371 (O_371,N_14984,N_14968);
nor UO_372 (O_372,N_14963,N_14919);
or UO_373 (O_373,N_14897,N_14913);
nor UO_374 (O_374,N_14913,N_14917);
nor UO_375 (O_375,N_14912,N_14959);
xnor UO_376 (O_376,N_14934,N_14936);
or UO_377 (O_377,N_14918,N_14989);
xnor UO_378 (O_378,N_14947,N_14952);
nor UO_379 (O_379,N_14978,N_14908);
and UO_380 (O_380,N_14961,N_14929);
nor UO_381 (O_381,N_14921,N_14988);
xnor UO_382 (O_382,N_14948,N_14896);
nand UO_383 (O_383,N_14922,N_14913);
or UO_384 (O_384,N_14925,N_14912);
nand UO_385 (O_385,N_14907,N_14973);
nor UO_386 (O_386,N_14929,N_14940);
or UO_387 (O_387,N_14898,N_14911);
nor UO_388 (O_388,N_14885,N_14952);
or UO_389 (O_389,N_14917,N_14971);
xor UO_390 (O_390,N_14934,N_14974);
nand UO_391 (O_391,N_14890,N_14929);
xor UO_392 (O_392,N_14977,N_14985);
nand UO_393 (O_393,N_14955,N_14890);
nor UO_394 (O_394,N_14955,N_14924);
xnor UO_395 (O_395,N_14979,N_14932);
and UO_396 (O_396,N_14969,N_14938);
nor UO_397 (O_397,N_14932,N_14933);
and UO_398 (O_398,N_14990,N_14982);
nor UO_399 (O_399,N_14972,N_14991);
and UO_400 (O_400,N_14934,N_14998);
or UO_401 (O_401,N_14931,N_14981);
or UO_402 (O_402,N_14882,N_14898);
nand UO_403 (O_403,N_14993,N_14957);
xor UO_404 (O_404,N_14885,N_14876);
or UO_405 (O_405,N_14877,N_14906);
xor UO_406 (O_406,N_14930,N_14893);
xor UO_407 (O_407,N_14920,N_14899);
xnor UO_408 (O_408,N_14886,N_14968);
nand UO_409 (O_409,N_14952,N_14906);
nor UO_410 (O_410,N_14883,N_14920);
nor UO_411 (O_411,N_14954,N_14911);
nand UO_412 (O_412,N_14901,N_14921);
nor UO_413 (O_413,N_14909,N_14936);
and UO_414 (O_414,N_14974,N_14981);
or UO_415 (O_415,N_14975,N_14996);
nor UO_416 (O_416,N_14933,N_14885);
xor UO_417 (O_417,N_14901,N_14960);
xor UO_418 (O_418,N_14963,N_14988);
nor UO_419 (O_419,N_14907,N_14963);
nand UO_420 (O_420,N_14878,N_14984);
or UO_421 (O_421,N_14980,N_14967);
and UO_422 (O_422,N_14963,N_14961);
and UO_423 (O_423,N_14917,N_14925);
nor UO_424 (O_424,N_14975,N_14971);
and UO_425 (O_425,N_14965,N_14942);
nand UO_426 (O_426,N_14912,N_14960);
or UO_427 (O_427,N_14875,N_14889);
nand UO_428 (O_428,N_14991,N_14980);
and UO_429 (O_429,N_14877,N_14882);
or UO_430 (O_430,N_14979,N_14986);
or UO_431 (O_431,N_14929,N_14939);
and UO_432 (O_432,N_14930,N_14877);
and UO_433 (O_433,N_14934,N_14880);
or UO_434 (O_434,N_14947,N_14892);
nor UO_435 (O_435,N_14933,N_14921);
nor UO_436 (O_436,N_14878,N_14894);
nand UO_437 (O_437,N_14974,N_14936);
nor UO_438 (O_438,N_14962,N_14942);
nand UO_439 (O_439,N_14914,N_14927);
nand UO_440 (O_440,N_14956,N_14922);
nor UO_441 (O_441,N_14967,N_14941);
nor UO_442 (O_442,N_14939,N_14957);
xor UO_443 (O_443,N_14911,N_14925);
and UO_444 (O_444,N_14997,N_14897);
and UO_445 (O_445,N_14982,N_14935);
and UO_446 (O_446,N_14906,N_14902);
or UO_447 (O_447,N_14968,N_14914);
and UO_448 (O_448,N_14964,N_14988);
nand UO_449 (O_449,N_14914,N_14959);
or UO_450 (O_450,N_14906,N_14909);
or UO_451 (O_451,N_14980,N_14953);
xnor UO_452 (O_452,N_14918,N_14981);
and UO_453 (O_453,N_14923,N_14892);
and UO_454 (O_454,N_14968,N_14985);
or UO_455 (O_455,N_14882,N_14936);
and UO_456 (O_456,N_14938,N_14994);
nand UO_457 (O_457,N_14945,N_14914);
nor UO_458 (O_458,N_14996,N_14945);
and UO_459 (O_459,N_14928,N_14909);
xnor UO_460 (O_460,N_14964,N_14911);
xor UO_461 (O_461,N_14902,N_14934);
or UO_462 (O_462,N_14987,N_14978);
xnor UO_463 (O_463,N_14907,N_14883);
nor UO_464 (O_464,N_14921,N_14913);
or UO_465 (O_465,N_14911,N_14880);
and UO_466 (O_466,N_14893,N_14920);
or UO_467 (O_467,N_14988,N_14980);
xnor UO_468 (O_468,N_14916,N_14962);
or UO_469 (O_469,N_14879,N_14920);
xor UO_470 (O_470,N_14925,N_14909);
and UO_471 (O_471,N_14985,N_14991);
nand UO_472 (O_472,N_14911,N_14903);
xnor UO_473 (O_473,N_14932,N_14907);
nand UO_474 (O_474,N_14892,N_14917);
nand UO_475 (O_475,N_14917,N_14908);
and UO_476 (O_476,N_14896,N_14932);
nor UO_477 (O_477,N_14912,N_14999);
nor UO_478 (O_478,N_14880,N_14930);
or UO_479 (O_479,N_14959,N_14934);
and UO_480 (O_480,N_14877,N_14881);
nand UO_481 (O_481,N_14889,N_14947);
xnor UO_482 (O_482,N_14995,N_14935);
xnor UO_483 (O_483,N_14994,N_14917);
and UO_484 (O_484,N_14877,N_14952);
xor UO_485 (O_485,N_14968,N_14938);
and UO_486 (O_486,N_14928,N_14967);
nand UO_487 (O_487,N_14941,N_14904);
nand UO_488 (O_488,N_14895,N_14877);
nor UO_489 (O_489,N_14902,N_14949);
nand UO_490 (O_490,N_14896,N_14882);
xor UO_491 (O_491,N_14942,N_14907);
nand UO_492 (O_492,N_14909,N_14948);
xnor UO_493 (O_493,N_14984,N_14924);
or UO_494 (O_494,N_14909,N_14986);
xor UO_495 (O_495,N_14976,N_14922);
and UO_496 (O_496,N_14977,N_14891);
nand UO_497 (O_497,N_14965,N_14914);
or UO_498 (O_498,N_14957,N_14897);
nor UO_499 (O_499,N_14931,N_14880);
xor UO_500 (O_500,N_14999,N_14922);
xor UO_501 (O_501,N_14941,N_14972);
or UO_502 (O_502,N_14892,N_14960);
nand UO_503 (O_503,N_14891,N_14911);
or UO_504 (O_504,N_14886,N_14924);
xnor UO_505 (O_505,N_14897,N_14950);
or UO_506 (O_506,N_14959,N_14920);
or UO_507 (O_507,N_14985,N_14936);
or UO_508 (O_508,N_14887,N_14954);
nor UO_509 (O_509,N_14882,N_14908);
nand UO_510 (O_510,N_14978,N_14881);
nand UO_511 (O_511,N_14932,N_14963);
or UO_512 (O_512,N_14890,N_14882);
nor UO_513 (O_513,N_14880,N_14986);
and UO_514 (O_514,N_14993,N_14878);
or UO_515 (O_515,N_14900,N_14976);
nor UO_516 (O_516,N_14946,N_14896);
nor UO_517 (O_517,N_14887,N_14950);
and UO_518 (O_518,N_14988,N_14876);
nand UO_519 (O_519,N_14959,N_14915);
and UO_520 (O_520,N_14895,N_14953);
or UO_521 (O_521,N_14897,N_14900);
or UO_522 (O_522,N_14915,N_14997);
nor UO_523 (O_523,N_14881,N_14933);
nor UO_524 (O_524,N_14928,N_14944);
and UO_525 (O_525,N_14957,N_14876);
nand UO_526 (O_526,N_14935,N_14913);
nor UO_527 (O_527,N_14993,N_14979);
xor UO_528 (O_528,N_14982,N_14923);
nor UO_529 (O_529,N_14993,N_14882);
nor UO_530 (O_530,N_14939,N_14995);
nor UO_531 (O_531,N_14969,N_14995);
or UO_532 (O_532,N_14984,N_14914);
xor UO_533 (O_533,N_14990,N_14893);
and UO_534 (O_534,N_14935,N_14890);
nor UO_535 (O_535,N_14896,N_14996);
and UO_536 (O_536,N_14975,N_14920);
nand UO_537 (O_537,N_14964,N_14989);
or UO_538 (O_538,N_14907,N_14916);
or UO_539 (O_539,N_14903,N_14912);
nor UO_540 (O_540,N_14957,N_14945);
nand UO_541 (O_541,N_14952,N_14949);
and UO_542 (O_542,N_14946,N_14905);
nand UO_543 (O_543,N_14977,N_14962);
or UO_544 (O_544,N_14951,N_14983);
nor UO_545 (O_545,N_14969,N_14890);
nand UO_546 (O_546,N_14892,N_14914);
or UO_547 (O_547,N_14896,N_14985);
and UO_548 (O_548,N_14961,N_14928);
or UO_549 (O_549,N_14982,N_14917);
or UO_550 (O_550,N_14890,N_14908);
or UO_551 (O_551,N_14882,N_14948);
xor UO_552 (O_552,N_14885,N_14978);
nand UO_553 (O_553,N_14961,N_14962);
or UO_554 (O_554,N_14967,N_14904);
or UO_555 (O_555,N_14907,N_14919);
nand UO_556 (O_556,N_14943,N_14931);
xor UO_557 (O_557,N_14976,N_14928);
and UO_558 (O_558,N_14936,N_14952);
nor UO_559 (O_559,N_14993,N_14876);
and UO_560 (O_560,N_14881,N_14996);
or UO_561 (O_561,N_14903,N_14963);
nor UO_562 (O_562,N_14887,N_14917);
nor UO_563 (O_563,N_14932,N_14960);
xor UO_564 (O_564,N_14913,N_14911);
and UO_565 (O_565,N_14918,N_14915);
nor UO_566 (O_566,N_14972,N_14931);
nor UO_567 (O_567,N_14981,N_14982);
nand UO_568 (O_568,N_14946,N_14995);
nand UO_569 (O_569,N_14891,N_14918);
nor UO_570 (O_570,N_14957,N_14885);
nand UO_571 (O_571,N_14988,N_14924);
xnor UO_572 (O_572,N_14904,N_14944);
nand UO_573 (O_573,N_14878,N_14875);
nor UO_574 (O_574,N_14876,N_14900);
or UO_575 (O_575,N_14978,N_14920);
xor UO_576 (O_576,N_14978,N_14909);
xor UO_577 (O_577,N_14950,N_14952);
or UO_578 (O_578,N_14896,N_14929);
nand UO_579 (O_579,N_14906,N_14975);
nand UO_580 (O_580,N_14967,N_14952);
or UO_581 (O_581,N_14981,N_14957);
and UO_582 (O_582,N_14914,N_14936);
nor UO_583 (O_583,N_14883,N_14889);
and UO_584 (O_584,N_14913,N_14885);
and UO_585 (O_585,N_14936,N_14955);
and UO_586 (O_586,N_14978,N_14977);
xnor UO_587 (O_587,N_14950,N_14955);
and UO_588 (O_588,N_14913,N_14994);
and UO_589 (O_589,N_14944,N_14936);
nor UO_590 (O_590,N_14902,N_14955);
and UO_591 (O_591,N_14991,N_14877);
nand UO_592 (O_592,N_14927,N_14904);
nor UO_593 (O_593,N_14912,N_14991);
and UO_594 (O_594,N_14906,N_14964);
nand UO_595 (O_595,N_14922,N_14889);
nor UO_596 (O_596,N_14987,N_14893);
and UO_597 (O_597,N_14906,N_14897);
nor UO_598 (O_598,N_14985,N_14998);
nand UO_599 (O_599,N_14965,N_14943);
nand UO_600 (O_600,N_14915,N_14923);
nor UO_601 (O_601,N_14901,N_14993);
nand UO_602 (O_602,N_14917,N_14996);
nor UO_603 (O_603,N_14904,N_14914);
nor UO_604 (O_604,N_14910,N_14875);
and UO_605 (O_605,N_14999,N_14930);
and UO_606 (O_606,N_14947,N_14999);
and UO_607 (O_607,N_14971,N_14914);
xnor UO_608 (O_608,N_14880,N_14884);
xor UO_609 (O_609,N_14905,N_14912);
xnor UO_610 (O_610,N_14982,N_14905);
nor UO_611 (O_611,N_14941,N_14917);
and UO_612 (O_612,N_14943,N_14891);
and UO_613 (O_613,N_14944,N_14965);
nand UO_614 (O_614,N_14997,N_14993);
nor UO_615 (O_615,N_14908,N_14995);
nor UO_616 (O_616,N_14881,N_14921);
and UO_617 (O_617,N_14908,N_14983);
nor UO_618 (O_618,N_14964,N_14946);
nor UO_619 (O_619,N_14883,N_14924);
xor UO_620 (O_620,N_14915,N_14904);
nor UO_621 (O_621,N_14978,N_14986);
and UO_622 (O_622,N_14955,N_14914);
and UO_623 (O_623,N_14949,N_14953);
or UO_624 (O_624,N_14968,N_14916);
xor UO_625 (O_625,N_14883,N_14903);
and UO_626 (O_626,N_14951,N_14981);
or UO_627 (O_627,N_14968,N_14922);
xnor UO_628 (O_628,N_14889,N_14985);
nor UO_629 (O_629,N_14884,N_14932);
nand UO_630 (O_630,N_14956,N_14934);
and UO_631 (O_631,N_14938,N_14904);
and UO_632 (O_632,N_14892,N_14913);
nand UO_633 (O_633,N_14919,N_14917);
or UO_634 (O_634,N_14960,N_14921);
nand UO_635 (O_635,N_14983,N_14980);
nand UO_636 (O_636,N_14886,N_14989);
or UO_637 (O_637,N_14922,N_14881);
and UO_638 (O_638,N_14980,N_14958);
nand UO_639 (O_639,N_14996,N_14918);
xor UO_640 (O_640,N_14903,N_14888);
and UO_641 (O_641,N_14894,N_14917);
or UO_642 (O_642,N_14960,N_14919);
and UO_643 (O_643,N_14897,N_14912);
xor UO_644 (O_644,N_14890,N_14996);
nor UO_645 (O_645,N_14876,N_14955);
and UO_646 (O_646,N_14971,N_14939);
xnor UO_647 (O_647,N_14999,N_14965);
or UO_648 (O_648,N_14883,N_14913);
xor UO_649 (O_649,N_14939,N_14886);
nor UO_650 (O_650,N_14946,N_14880);
nor UO_651 (O_651,N_14953,N_14916);
and UO_652 (O_652,N_14967,N_14939);
xor UO_653 (O_653,N_14967,N_14892);
and UO_654 (O_654,N_14972,N_14913);
nand UO_655 (O_655,N_14943,N_14938);
nand UO_656 (O_656,N_14997,N_14943);
nand UO_657 (O_657,N_14993,N_14919);
xnor UO_658 (O_658,N_14875,N_14974);
or UO_659 (O_659,N_14894,N_14992);
nor UO_660 (O_660,N_14941,N_14952);
xor UO_661 (O_661,N_14966,N_14941);
or UO_662 (O_662,N_14896,N_14903);
nor UO_663 (O_663,N_14901,N_14931);
and UO_664 (O_664,N_14992,N_14998);
xor UO_665 (O_665,N_14922,N_14932);
or UO_666 (O_666,N_14951,N_14895);
xnor UO_667 (O_667,N_14945,N_14931);
and UO_668 (O_668,N_14875,N_14901);
xor UO_669 (O_669,N_14899,N_14994);
nor UO_670 (O_670,N_14952,N_14922);
and UO_671 (O_671,N_14912,N_14992);
and UO_672 (O_672,N_14980,N_14924);
xor UO_673 (O_673,N_14957,N_14875);
nand UO_674 (O_674,N_14971,N_14981);
xor UO_675 (O_675,N_14900,N_14946);
or UO_676 (O_676,N_14899,N_14932);
nor UO_677 (O_677,N_14933,N_14949);
or UO_678 (O_678,N_14931,N_14924);
nor UO_679 (O_679,N_14913,N_14967);
nor UO_680 (O_680,N_14952,N_14905);
nor UO_681 (O_681,N_14893,N_14907);
nand UO_682 (O_682,N_14891,N_14995);
nor UO_683 (O_683,N_14979,N_14981);
and UO_684 (O_684,N_14995,N_14899);
or UO_685 (O_685,N_14912,N_14920);
or UO_686 (O_686,N_14891,N_14991);
xor UO_687 (O_687,N_14999,N_14942);
and UO_688 (O_688,N_14932,N_14939);
and UO_689 (O_689,N_14877,N_14944);
xnor UO_690 (O_690,N_14899,N_14988);
xor UO_691 (O_691,N_14975,N_14884);
nor UO_692 (O_692,N_14967,N_14959);
nor UO_693 (O_693,N_14936,N_14977);
nor UO_694 (O_694,N_14922,N_14984);
xnor UO_695 (O_695,N_14927,N_14876);
nand UO_696 (O_696,N_14910,N_14920);
or UO_697 (O_697,N_14898,N_14969);
and UO_698 (O_698,N_14884,N_14930);
or UO_699 (O_699,N_14907,N_14905);
xor UO_700 (O_700,N_14976,N_14886);
nand UO_701 (O_701,N_14884,N_14982);
nand UO_702 (O_702,N_14983,N_14879);
or UO_703 (O_703,N_14924,N_14953);
xor UO_704 (O_704,N_14951,N_14897);
or UO_705 (O_705,N_14906,N_14959);
nor UO_706 (O_706,N_14989,N_14896);
and UO_707 (O_707,N_14995,N_14951);
xnor UO_708 (O_708,N_14973,N_14879);
xor UO_709 (O_709,N_14990,N_14937);
or UO_710 (O_710,N_14972,N_14916);
or UO_711 (O_711,N_14887,N_14895);
and UO_712 (O_712,N_14921,N_14995);
or UO_713 (O_713,N_14973,N_14882);
and UO_714 (O_714,N_14922,N_14882);
nand UO_715 (O_715,N_14976,N_14921);
nor UO_716 (O_716,N_14986,N_14875);
nand UO_717 (O_717,N_14901,N_14976);
and UO_718 (O_718,N_14910,N_14938);
xnor UO_719 (O_719,N_14920,N_14880);
xor UO_720 (O_720,N_14894,N_14958);
and UO_721 (O_721,N_14984,N_14967);
and UO_722 (O_722,N_14925,N_14956);
and UO_723 (O_723,N_14989,N_14965);
or UO_724 (O_724,N_14935,N_14971);
xnor UO_725 (O_725,N_14904,N_14911);
xor UO_726 (O_726,N_14943,N_14953);
or UO_727 (O_727,N_14969,N_14993);
or UO_728 (O_728,N_14937,N_14935);
or UO_729 (O_729,N_14959,N_14885);
xor UO_730 (O_730,N_14999,N_14876);
nand UO_731 (O_731,N_14909,N_14995);
xor UO_732 (O_732,N_14876,N_14963);
nor UO_733 (O_733,N_14887,N_14906);
or UO_734 (O_734,N_14994,N_14964);
and UO_735 (O_735,N_14891,N_14877);
or UO_736 (O_736,N_14909,N_14979);
nor UO_737 (O_737,N_14912,N_14966);
xor UO_738 (O_738,N_14988,N_14991);
or UO_739 (O_739,N_14916,N_14985);
nand UO_740 (O_740,N_14988,N_14915);
nand UO_741 (O_741,N_14996,N_14926);
xor UO_742 (O_742,N_14905,N_14891);
nand UO_743 (O_743,N_14939,N_14955);
nand UO_744 (O_744,N_14910,N_14995);
or UO_745 (O_745,N_14969,N_14977);
xnor UO_746 (O_746,N_14935,N_14931);
nor UO_747 (O_747,N_14914,N_14899);
and UO_748 (O_748,N_14949,N_14966);
nor UO_749 (O_749,N_14875,N_14924);
or UO_750 (O_750,N_14924,N_14919);
and UO_751 (O_751,N_14888,N_14881);
xor UO_752 (O_752,N_14966,N_14943);
or UO_753 (O_753,N_14979,N_14882);
and UO_754 (O_754,N_14959,N_14943);
nand UO_755 (O_755,N_14971,N_14886);
or UO_756 (O_756,N_14925,N_14880);
or UO_757 (O_757,N_14962,N_14891);
nand UO_758 (O_758,N_14923,N_14960);
xnor UO_759 (O_759,N_14898,N_14964);
xor UO_760 (O_760,N_14932,N_14995);
and UO_761 (O_761,N_14903,N_14958);
or UO_762 (O_762,N_14962,N_14880);
or UO_763 (O_763,N_14991,N_14898);
nor UO_764 (O_764,N_14909,N_14885);
xnor UO_765 (O_765,N_14909,N_14965);
and UO_766 (O_766,N_14991,N_14918);
or UO_767 (O_767,N_14941,N_14988);
xor UO_768 (O_768,N_14879,N_14932);
xnor UO_769 (O_769,N_14892,N_14936);
nor UO_770 (O_770,N_14981,N_14920);
and UO_771 (O_771,N_14940,N_14928);
nand UO_772 (O_772,N_14965,N_14897);
xor UO_773 (O_773,N_14881,N_14894);
nor UO_774 (O_774,N_14899,N_14877);
nor UO_775 (O_775,N_14910,N_14878);
and UO_776 (O_776,N_14886,N_14928);
or UO_777 (O_777,N_14935,N_14920);
nand UO_778 (O_778,N_14981,N_14888);
xnor UO_779 (O_779,N_14947,N_14962);
and UO_780 (O_780,N_14915,N_14950);
nand UO_781 (O_781,N_14888,N_14926);
xnor UO_782 (O_782,N_14936,N_14913);
nor UO_783 (O_783,N_14974,N_14916);
nand UO_784 (O_784,N_14991,N_14906);
xor UO_785 (O_785,N_14877,N_14914);
or UO_786 (O_786,N_14990,N_14996);
xor UO_787 (O_787,N_14918,N_14939);
or UO_788 (O_788,N_14969,N_14936);
and UO_789 (O_789,N_14929,N_14908);
nor UO_790 (O_790,N_14886,N_14950);
nand UO_791 (O_791,N_14985,N_14980);
and UO_792 (O_792,N_14906,N_14965);
xor UO_793 (O_793,N_14895,N_14961);
or UO_794 (O_794,N_14926,N_14978);
or UO_795 (O_795,N_14899,N_14930);
nand UO_796 (O_796,N_14881,N_14898);
and UO_797 (O_797,N_14944,N_14929);
nand UO_798 (O_798,N_14916,N_14988);
nor UO_799 (O_799,N_14916,N_14891);
nand UO_800 (O_800,N_14977,N_14922);
nand UO_801 (O_801,N_14929,N_14979);
nor UO_802 (O_802,N_14893,N_14914);
nand UO_803 (O_803,N_14955,N_14906);
nor UO_804 (O_804,N_14932,N_14968);
xnor UO_805 (O_805,N_14984,N_14960);
or UO_806 (O_806,N_14884,N_14942);
and UO_807 (O_807,N_14956,N_14962);
or UO_808 (O_808,N_14949,N_14913);
nand UO_809 (O_809,N_14995,N_14956);
and UO_810 (O_810,N_14996,N_14910);
nand UO_811 (O_811,N_14992,N_14896);
and UO_812 (O_812,N_14876,N_14947);
and UO_813 (O_813,N_14987,N_14952);
and UO_814 (O_814,N_14940,N_14978);
or UO_815 (O_815,N_14924,N_14887);
nand UO_816 (O_816,N_14987,N_14959);
and UO_817 (O_817,N_14949,N_14907);
or UO_818 (O_818,N_14944,N_14940);
nand UO_819 (O_819,N_14951,N_14892);
xnor UO_820 (O_820,N_14944,N_14971);
and UO_821 (O_821,N_14907,N_14982);
and UO_822 (O_822,N_14976,N_14959);
nand UO_823 (O_823,N_14895,N_14933);
or UO_824 (O_824,N_14956,N_14987);
or UO_825 (O_825,N_14964,N_14999);
or UO_826 (O_826,N_14952,N_14932);
nor UO_827 (O_827,N_14958,N_14878);
and UO_828 (O_828,N_14917,N_14900);
nand UO_829 (O_829,N_14947,N_14923);
or UO_830 (O_830,N_14965,N_14973);
or UO_831 (O_831,N_14885,N_14963);
or UO_832 (O_832,N_14953,N_14991);
nand UO_833 (O_833,N_14998,N_14961);
nand UO_834 (O_834,N_14948,N_14950);
nand UO_835 (O_835,N_14919,N_14959);
xnor UO_836 (O_836,N_14973,N_14993);
xor UO_837 (O_837,N_14992,N_14877);
or UO_838 (O_838,N_14947,N_14920);
nor UO_839 (O_839,N_14992,N_14997);
nand UO_840 (O_840,N_14983,N_14892);
xnor UO_841 (O_841,N_14937,N_14902);
nand UO_842 (O_842,N_14894,N_14932);
or UO_843 (O_843,N_14923,N_14966);
nor UO_844 (O_844,N_14906,N_14981);
nand UO_845 (O_845,N_14907,N_14945);
nor UO_846 (O_846,N_14963,N_14985);
or UO_847 (O_847,N_14891,N_14887);
xnor UO_848 (O_848,N_14911,N_14963);
nor UO_849 (O_849,N_14975,N_14890);
nand UO_850 (O_850,N_14879,N_14916);
nor UO_851 (O_851,N_14928,N_14983);
xor UO_852 (O_852,N_14978,N_14938);
nand UO_853 (O_853,N_14921,N_14968);
or UO_854 (O_854,N_14950,N_14964);
xnor UO_855 (O_855,N_14935,N_14945);
nor UO_856 (O_856,N_14998,N_14984);
or UO_857 (O_857,N_14955,N_14985);
nand UO_858 (O_858,N_14991,N_14942);
xor UO_859 (O_859,N_14992,N_14994);
nand UO_860 (O_860,N_14927,N_14941);
nand UO_861 (O_861,N_14949,N_14899);
or UO_862 (O_862,N_14977,N_14973);
xnor UO_863 (O_863,N_14906,N_14972);
and UO_864 (O_864,N_14975,N_14918);
nand UO_865 (O_865,N_14961,N_14973);
nor UO_866 (O_866,N_14960,N_14990);
and UO_867 (O_867,N_14973,N_14997);
xor UO_868 (O_868,N_14935,N_14881);
nand UO_869 (O_869,N_14901,N_14955);
nand UO_870 (O_870,N_14953,N_14933);
xor UO_871 (O_871,N_14985,N_14920);
and UO_872 (O_872,N_14877,N_14915);
xor UO_873 (O_873,N_14985,N_14907);
and UO_874 (O_874,N_14994,N_14970);
nand UO_875 (O_875,N_14946,N_14927);
nor UO_876 (O_876,N_14957,N_14980);
or UO_877 (O_877,N_14897,N_14915);
or UO_878 (O_878,N_14884,N_14972);
xnor UO_879 (O_879,N_14884,N_14970);
xnor UO_880 (O_880,N_14969,N_14954);
or UO_881 (O_881,N_14962,N_14948);
xor UO_882 (O_882,N_14882,N_14937);
xor UO_883 (O_883,N_14901,N_14886);
and UO_884 (O_884,N_14886,N_14962);
nand UO_885 (O_885,N_14952,N_14931);
or UO_886 (O_886,N_14911,N_14907);
nand UO_887 (O_887,N_14906,N_14912);
or UO_888 (O_888,N_14875,N_14894);
and UO_889 (O_889,N_14939,N_14982);
xor UO_890 (O_890,N_14962,N_14909);
nor UO_891 (O_891,N_14968,N_14978);
nor UO_892 (O_892,N_14913,N_14933);
xor UO_893 (O_893,N_14976,N_14964);
nand UO_894 (O_894,N_14955,N_14994);
nor UO_895 (O_895,N_14900,N_14938);
xnor UO_896 (O_896,N_14993,N_14984);
or UO_897 (O_897,N_14976,N_14895);
nor UO_898 (O_898,N_14989,N_14987);
nor UO_899 (O_899,N_14951,N_14960);
and UO_900 (O_900,N_14933,N_14981);
or UO_901 (O_901,N_14889,N_14924);
and UO_902 (O_902,N_14900,N_14942);
nand UO_903 (O_903,N_14975,N_14944);
or UO_904 (O_904,N_14945,N_14893);
nand UO_905 (O_905,N_14888,N_14883);
and UO_906 (O_906,N_14952,N_14972);
xor UO_907 (O_907,N_14953,N_14898);
xor UO_908 (O_908,N_14919,N_14962);
xor UO_909 (O_909,N_14937,N_14977);
or UO_910 (O_910,N_14889,N_14998);
and UO_911 (O_911,N_14918,N_14886);
xor UO_912 (O_912,N_14966,N_14893);
or UO_913 (O_913,N_14908,N_14910);
nand UO_914 (O_914,N_14967,N_14922);
nor UO_915 (O_915,N_14927,N_14961);
or UO_916 (O_916,N_14953,N_14928);
nor UO_917 (O_917,N_14939,N_14994);
nand UO_918 (O_918,N_14986,N_14977);
nor UO_919 (O_919,N_14943,N_14975);
or UO_920 (O_920,N_14890,N_14893);
nand UO_921 (O_921,N_14924,N_14927);
xnor UO_922 (O_922,N_14965,N_14934);
and UO_923 (O_923,N_14886,N_14910);
or UO_924 (O_924,N_14876,N_14918);
xnor UO_925 (O_925,N_14973,N_14922);
nor UO_926 (O_926,N_14897,N_14945);
or UO_927 (O_927,N_14990,N_14969);
nor UO_928 (O_928,N_14897,N_14907);
nand UO_929 (O_929,N_14882,N_14953);
nand UO_930 (O_930,N_14943,N_14924);
or UO_931 (O_931,N_14955,N_14900);
or UO_932 (O_932,N_14962,N_14930);
nor UO_933 (O_933,N_14951,N_14941);
and UO_934 (O_934,N_14954,N_14987);
nor UO_935 (O_935,N_14998,N_14996);
or UO_936 (O_936,N_14907,N_14908);
xor UO_937 (O_937,N_14914,N_14956);
or UO_938 (O_938,N_14923,N_14878);
xnor UO_939 (O_939,N_14876,N_14952);
xnor UO_940 (O_940,N_14984,N_14988);
and UO_941 (O_941,N_14896,N_14927);
or UO_942 (O_942,N_14907,N_14887);
nor UO_943 (O_943,N_14996,N_14931);
or UO_944 (O_944,N_14881,N_14973);
xor UO_945 (O_945,N_14928,N_14905);
and UO_946 (O_946,N_14886,N_14927);
xnor UO_947 (O_947,N_14909,N_14940);
and UO_948 (O_948,N_14984,N_14969);
nand UO_949 (O_949,N_14934,N_14948);
nand UO_950 (O_950,N_14916,N_14996);
nor UO_951 (O_951,N_14898,N_14940);
or UO_952 (O_952,N_14935,N_14967);
nand UO_953 (O_953,N_14960,N_14903);
or UO_954 (O_954,N_14968,N_14877);
nand UO_955 (O_955,N_14877,N_14998);
and UO_956 (O_956,N_14884,N_14980);
nor UO_957 (O_957,N_14974,N_14954);
xor UO_958 (O_958,N_14980,N_14942);
and UO_959 (O_959,N_14898,N_14917);
and UO_960 (O_960,N_14928,N_14954);
nor UO_961 (O_961,N_14966,N_14884);
xnor UO_962 (O_962,N_14962,N_14931);
and UO_963 (O_963,N_14989,N_14922);
nor UO_964 (O_964,N_14930,N_14896);
nor UO_965 (O_965,N_14878,N_14941);
nor UO_966 (O_966,N_14943,N_14914);
nor UO_967 (O_967,N_14942,N_14891);
and UO_968 (O_968,N_14881,N_14906);
nor UO_969 (O_969,N_14977,N_14882);
and UO_970 (O_970,N_14957,N_14954);
or UO_971 (O_971,N_14961,N_14910);
and UO_972 (O_972,N_14975,N_14949);
xor UO_973 (O_973,N_14970,N_14939);
and UO_974 (O_974,N_14964,N_14945);
xor UO_975 (O_975,N_14972,N_14929);
nand UO_976 (O_976,N_14988,N_14932);
and UO_977 (O_977,N_14925,N_14923);
and UO_978 (O_978,N_14881,N_14880);
or UO_979 (O_979,N_14887,N_14919);
nor UO_980 (O_980,N_14934,N_14909);
xor UO_981 (O_981,N_14901,N_14946);
nand UO_982 (O_982,N_14919,N_14935);
nor UO_983 (O_983,N_14896,N_14941);
nand UO_984 (O_984,N_14952,N_14996);
nor UO_985 (O_985,N_14987,N_14949);
or UO_986 (O_986,N_14974,N_14885);
or UO_987 (O_987,N_14887,N_14889);
xor UO_988 (O_988,N_14949,N_14925);
nand UO_989 (O_989,N_14967,N_14920);
or UO_990 (O_990,N_14898,N_14883);
or UO_991 (O_991,N_14965,N_14969);
and UO_992 (O_992,N_14934,N_14929);
xnor UO_993 (O_993,N_14962,N_14929);
and UO_994 (O_994,N_14933,N_14943);
xnor UO_995 (O_995,N_14920,N_14996);
nor UO_996 (O_996,N_14981,N_14990);
nor UO_997 (O_997,N_14948,N_14996);
and UO_998 (O_998,N_14997,N_14929);
or UO_999 (O_999,N_14882,N_14933);
nor UO_1000 (O_1000,N_14989,N_14968);
or UO_1001 (O_1001,N_14958,N_14941);
or UO_1002 (O_1002,N_14989,N_14974);
nor UO_1003 (O_1003,N_14926,N_14915);
xnor UO_1004 (O_1004,N_14994,N_14949);
or UO_1005 (O_1005,N_14927,N_14930);
and UO_1006 (O_1006,N_14921,N_14954);
and UO_1007 (O_1007,N_14902,N_14915);
or UO_1008 (O_1008,N_14884,N_14892);
or UO_1009 (O_1009,N_14985,N_14942);
nand UO_1010 (O_1010,N_14980,N_14961);
or UO_1011 (O_1011,N_14917,N_14879);
nand UO_1012 (O_1012,N_14876,N_14951);
xor UO_1013 (O_1013,N_14890,N_14887);
xnor UO_1014 (O_1014,N_14935,N_14896);
nand UO_1015 (O_1015,N_14991,N_14876);
and UO_1016 (O_1016,N_14934,N_14997);
or UO_1017 (O_1017,N_14915,N_14983);
or UO_1018 (O_1018,N_14957,N_14958);
and UO_1019 (O_1019,N_14943,N_14916);
nor UO_1020 (O_1020,N_14932,N_14970);
or UO_1021 (O_1021,N_14883,N_14895);
nor UO_1022 (O_1022,N_14931,N_14929);
nand UO_1023 (O_1023,N_14940,N_14902);
nor UO_1024 (O_1024,N_14961,N_14901);
or UO_1025 (O_1025,N_14984,N_14977);
xor UO_1026 (O_1026,N_14889,N_14928);
or UO_1027 (O_1027,N_14984,N_14895);
or UO_1028 (O_1028,N_14903,N_14978);
nor UO_1029 (O_1029,N_14920,N_14924);
xnor UO_1030 (O_1030,N_14967,N_14990);
or UO_1031 (O_1031,N_14916,N_14944);
nand UO_1032 (O_1032,N_14994,N_14960);
and UO_1033 (O_1033,N_14945,N_14876);
and UO_1034 (O_1034,N_14924,N_14996);
or UO_1035 (O_1035,N_14924,N_14912);
or UO_1036 (O_1036,N_14970,N_14907);
nor UO_1037 (O_1037,N_14882,N_14984);
xor UO_1038 (O_1038,N_14953,N_14932);
or UO_1039 (O_1039,N_14969,N_14999);
nand UO_1040 (O_1040,N_14983,N_14887);
and UO_1041 (O_1041,N_14893,N_14947);
nand UO_1042 (O_1042,N_14998,N_14928);
or UO_1043 (O_1043,N_14895,N_14876);
nor UO_1044 (O_1044,N_14946,N_14944);
nor UO_1045 (O_1045,N_14988,N_14985);
nand UO_1046 (O_1046,N_14875,N_14886);
or UO_1047 (O_1047,N_14935,N_14875);
and UO_1048 (O_1048,N_14936,N_14996);
and UO_1049 (O_1049,N_14974,N_14913);
nor UO_1050 (O_1050,N_14903,N_14939);
xnor UO_1051 (O_1051,N_14997,N_14889);
or UO_1052 (O_1052,N_14947,N_14943);
and UO_1053 (O_1053,N_14901,N_14879);
and UO_1054 (O_1054,N_14964,N_14895);
or UO_1055 (O_1055,N_14883,N_14964);
and UO_1056 (O_1056,N_14982,N_14929);
nand UO_1057 (O_1057,N_14952,N_14923);
xor UO_1058 (O_1058,N_14962,N_14971);
or UO_1059 (O_1059,N_14929,N_14974);
and UO_1060 (O_1060,N_14928,N_14883);
or UO_1061 (O_1061,N_14973,N_14953);
nor UO_1062 (O_1062,N_14932,N_14911);
or UO_1063 (O_1063,N_14876,N_14917);
xnor UO_1064 (O_1064,N_14942,N_14973);
xnor UO_1065 (O_1065,N_14982,N_14919);
nor UO_1066 (O_1066,N_14968,N_14923);
or UO_1067 (O_1067,N_14920,N_14955);
or UO_1068 (O_1068,N_14948,N_14986);
and UO_1069 (O_1069,N_14998,N_14884);
nand UO_1070 (O_1070,N_14945,N_14894);
and UO_1071 (O_1071,N_14988,N_14922);
xnor UO_1072 (O_1072,N_14917,N_14943);
nor UO_1073 (O_1073,N_14941,N_14934);
xnor UO_1074 (O_1074,N_14986,N_14924);
and UO_1075 (O_1075,N_14948,N_14930);
xnor UO_1076 (O_1076,N_14918,N_14914);
xor UO_1077 (O_1077,N_14982,N_14926);
or UO_1078 (O_1078,N_14997,N_14979);
nand UO_1079 (O_1079,N_14997,N_14950);
xor UO_1080 (O_1080,N_14891,N_14903);
nand UO_1081 (O_1081,N_14904,N_14920);
nand UO_1082 (O_1082,N_14919,N_14946);
nand UO_1083 (O_1083,N_14943,N_14910);
nand UO_1084 (O_1084,N_14879,N_14955);
nand UO_1085 (O_1085,N_14915,N_14961);
nor UO_1086 (O_1086,N_14918,N_14920);
and UO_1087 (O_1087,N_14993,N_14987);
or UO_1088 (O_1088,N_14955,N_14912);
and UO_1089 (O_1089,N_14981,N_14891);
nor UO_1090 (O_1090,N_14913,N_14951);
nand UO_1091 (O_1091,N_14974,N_14994);
nor UO_1092 (O_1092,N_14894,N_14990);
and UO_1093 (O_1093,N_14902,N_14896);
or UO_1094 (O_1094,N_14940,N_14882);
nand UO_1095 (O_1095,N_14949,N_14957);
xnor UO_1096 (O_1096,N_14876,N_14980);
and UO_1097 (O_1097,N_14984,N_14923);
nand UO_1098 (O_1098,N_14958,N_14987);
xnor UO_1099 (O_1099,N_14971,N_14974);
nand UO_1100 (O_1100,N_14919,N_14893);
xor UO_1101 (O_1101,N_14981,N_14972);
nor UO_1102 (O_1102,N_14933,N_14938);
nor UO_1103 (O_1103,N_14950,N_14954);
nand UO_1104 (O_1104,N_14878,N_14939);
xor UO_1105 (O_1105,N_14958,N_14979);
nand UO_1106 (O_1106,N_14898,N_14904);
or UO_1107 (O_1107,N_14983,N_14896);
nor UO_1108 (O_1108,N_14937,N_14975);
and UO_1109 (O_1109,N_14967,N_14924);
or UO_1110 (O_1110,N_14892,N_14996);
xor UO_1111 (O_1111,N_14966,N_14982);
nand UO_1112 (O_1112,N_14937,N_14913);
xor UO_1113 (O_1113,N_14969,N_14991);
and UO_1114 (O_1114,N_14983,N_14954);
or UO_1115 (O_1115,N_14997,N_14965);
or UO_1116 (O_1116,N_14889,N_14948);
nor UO_1117 (O_1117,N_14991,N_14962);
nor UO_1118 (O_1118,N_14964,N_14878);
or UO_1119 (O_1119,N_14963,N_14934);
or UO_1120 (O_1120,N_14958,N_14999);
and UO_1121 (O_1121,N_14895,N_14994);
and UO_1122 (O_1122,N_14918,N_14982);
xnor UO_1123 (O_1123,N_14960,N_14891);
xnor UO_1124 (O_1124,N_14987,N_14951);
nor UO_1125 (O_1125,N_14952,N_14980);
nor UO_1126 (O_1126,N_14926,N_14881);
or UO_1127 (O_1127,N_14957,N_14890);
xor UO_1128 (O_1128,N_14881,N_14943);
nand UO_1129 (O_1129,N_14946,N_14952);
and UO_1130 (O_1130,N_14913,N_14880);
nand UO_1131 (O_1131,N_14898,N_14897);
nand UO_1132 (O_1132,N_14905,N_14895);
nor UO_1133 (O_1133,N_14945,N_14954);
or UO_1134 (O_1134,N_14985,N_14976);
nand UO_1135 (O_1135,N_14931,N_14975);
nand UO_1136 (O_1136,N_14946,N_14892);
or UO_1137 (O_1137,N_14897,N_14885);
or UO_1138 (O_1138,N_14944,N_14987);
nand UO_1139 (O_1139,N_14954,N_14992);
and UO_1140 (O_1140,N_14892,N_14886);
nor UO_1141 (O_1141,N_14952,N_14969);
and UO_1142 (O_1142,N_14976,N_14941);
nand UO_1143 (O_1143,N_14954,N_14962);
xor UO_1144 (O_1144,N_14983,N_14977);
xor UO_1145 (O_1145,N_14911,N_14987);
nor UO_1146 (O_1146,N_14895,N_14986);
or UO_1147 (O_1147,N_14910,N_14933);
or UO_1148 (O_1148,N_14972,N_14904);
or UO_1149 (O_1149,N_14917,N_14980);
nand UO_1150 (O_1150,N_14922,N_14995);
and UO_1151 (O_1151,N_14990,N_14997);
and UO_1152 (O_1152,N_14920,N_14915);
and UO_1153 (O_1153,N_14896,N_14980);
nor UO_1154 (O_1154,N_14908,N_14989);
or UO_1155 (O_1155,N_14896,N_14888);
xor UO_1156 (O_1156,N_14907,N_14999);
and UO_1157 (O_1157,N_14955,N_14922);
nand UO_1158 (O_1158,N_14959,N_14910);
and UO_1159 (O_1159,N_14904,N_14913);
nand UO_1160 (O_1160,N_14937,N_14950);
or UO_1161 (O_1161,N_14892,N_14980);
nor UO_1162 (O_1162,N_14912,N_14972);
nor UO_1163 (O_1163,N_14997,N_14893);
or UO_1164 (O_1164,N_14906,N_14997);
xor UO_1165 (O_1165,N_14904,N_14894);
nor UO_1166 (O_1166,N_14955,N_14897);
or UO_1167 (O_1167,N_14915,N_14984);
and UO_1168 (O_1168,N_14975,N_14898);
nand UO_1169 (O_1169,N_14902,N_14880);
nor UO_1170 (O_1170,N_14877,N_14941);
xnor UO_1171 (O_1171,N_14910,N_14926);
or UO_1172 (O_1172,N_14976,N_14992);
nor UO_1173 (O_1173,N_14916,N_14978);
nor UO_1174 (O_1174,N_14877,N_14943);
nand UO_1175 (O_1175,N_14893,N_14908);
nand UO_1176 (O_1176,N_14887,N_14923);
xor UO_1177 (O_1177,N_14893,N_14910);
or UO_1178 (O_1178,N_14894,N_14900);
or UO_1179 (O_1179,N_14879,N_14952);
xor UO_1180 (O_1180,N_14917,N_14895);
nand UO_1181 (O_1181,N_14987,N_14988);
or UO_1182 (O_1182,N_14992,N_14965);
nand UO_1183 (O_1183,N_14892,N_14889);
and UO_1184 (O_1184,N_14985,N_14879);
xnor UO_1185 (O_1185,N_14942,N_14897);
xnor UO_1186 (O_1186,N_14967,N_14997);
and UO_1187 (O_1187,N_14973,N_14954);
xor UO_1188 (O_1188,N_14971,N_14916);
nand UO_1189 (O_1189,N_14944,N_14970);
or UO_1190 (O_1190,N_14892,N_14927);
and UO_1191 (O_1191,N_14978,N_14927);
nor UO_1192 (O_1192,N_14935,N_14976);
and UO_1193 (O_1193,N_14966,N_14958);
and UO_1194 (O_1194,N_14948,N_14946);
or UO_1195 (O_1195,N_14933,N_14946);
nor UO_1196 (O_1196,N_14936,N_14948);
or UO_1197 (O_1197,N_14941,N_14987);
xnor UO_1198 (O_1198,N_14998,N_14967);
nor UO_1199 (O_1199,N_14998,N_14964);
nand UO_1200 (O_1200,N_14876,N_14992);
and UO_1201 (O_1201,N_14975,N_14980);
xnor UO_1202 (O_1202,N_14904,N_14945);
and UO_1203 (O_1203,N_14998,N_14991);
and UO_1204 (O_1204,N_14987,N_14875);
nor UO_1205 (O_1205,N_14944,N_14994);
xnor UO_1206 (O_1206,N_14938,N_14901);
or UO_1207 (O_1207,N_14922,N_14912);
or UO_1208 (O_1208,N_14926,N_14920);
and UO_1209 (O_1209,N_14892,N_14956);
and UO_1210 (O_1210,N_14957,N_14994);
nand UO_1211 (O_1211,N_14971,N_14968);
xnor UO_1212 (O_1212,N_14895,N_14979);
xnor UO_1213 (O_1213,N_14932,N_14924);
xnor UO_1214 (O_1214,N_14976,N_14975);
nand UO_1215 (O_1215,N_14882,N_14876);
or UO_1216 (O_1216,N_14897,N_14992);
nor UO_1217 (O_1217,N_14957,N_14898);
nor UO_1218 (O_1218,N_14920,N_14933);
and UO_1219 (O_1219,N_14890,N_14944);
xnor UO_1220 (O_1220,N_14937,N_14980);
nor UO_1221 (O_1221,N_14892,N_14934);
or UO_1222 (O_1222,N_14945,N_14983);
nand UO_1223 (O_1223,N_14933,N_14934);
xor UO_1224 (O_1224,N_14924,N_14917);
nor UO_1225 (O_1225,N_14998,N_14880);
and UO_1226 (O_1226,N_14892,N_14975);
nor UO_1227 (O_1227,N_14925,N_14907);
xor UO_1228 (O_1228,N_14883,N_14978);
and UO_1229 (O_1229,N_14875,N_14964);
xor UO_1230 (O_1230,N_14974,N_14920);
or UO_1231 (O_1231,N_14884,N_14973);
nand UO_1232 (O_1232,N_14895,N_14913);
xor UO_1233 (O_1233,N_14889,N_14990);
xnor UO_1234 (O_1234,N_14906,N_14941);
and UO_1235 (O_1235,N_14888,N_14957);
nor UO_1236 (O_1236,N_14963,N_14965);
and UO_1237 (O_1237,N_14906,N_14903);
nand UO_1238 (O_1238,N_14978,N_14966);
xnor UO_1239 (O_1239,N_14885,N_14881);
and UO_1240 (O_1240,N_14994,N_14909);
nor UO_1241 (O_1241,N_14997,N_14908);
nor UO_1242 (O_1242,N_14877,N_14887);
xor UO_1243 (O_1243,N_14994,N_14972);
nand UO_1244 (O_1244,N_14939,N_14876);
nand UO_1245 (O_1245,N_14981,N_14997);
nand UO_1246 (O_1246,N_14983,N_14981);
xor UO_1247 (O_1247,N_14944,N_14881);
nor UO_1248 (O_1248,N_14920,N_14922);
and UO_1249 (O_1249,N_14998,N_14990);
xor UO_1250 (O_1250,N_14943,N_14894);
and UO_1251 (O_1251,N_14984,N_14948);
nand UO_1252 (O_1252,N_14916,N_14960);
or UO_1253 (O_1253,N_14899,N_14900);
nand UO_1254 (O_1254,N_14999,N_14967);
and UO_1255 (O_1255,N_14988,N_14958);
xnor UO_1256 (O_1256,N_14973,N_14914);
nand UO_1257 (O_1257,N_14903,N_14901);
nand UO_1258 (O_1258,N_14932,N_14923);
xnor UO_1259 (O_1259,N_14883,N_14990);
nand UO_1260 (O_1260,N_14952,N_14968);
nand UO_1261 (O_1261,N_14883,N_14987);
nor UO_1262 (O_1262,N_14947,N_14908);
xor UO_1263 (O_1263,N_14925,N_14959);
nand UO_1264 (O_1264,N_14927,N_14940);
xor UO_1265 (O_1265,N_14890,N_14943);
nor UO_1266 (O_1266,N_14879,N_14937);
and UO_1267 (O_1267,N_14928,N_14901);
nand UO_1268 (O_1268,N_14973,N_14988);
nor UO_1269 (O_1269,N_14908,N_14883);
nor UO_1270 (O_1270,N_14923,N_14901);
and UO_1271 (O_1271,N_14935,N_14932);
nand UO_1272 (O_1272,N_14932,N_14981);
and UO_1273 (O_1273,N_14972,N_14922);
nor UO_1274 (O_1274,N_14895,N_14998);
and UO_1275 (O_1275,N_14878,N_14925);
or UO_1276 (O_1276,N_14933,N_14893);
nand UO_1277 (O_1277,N_14906,N_14957);
and UO_1278 (O_1278,N_14910,N_14928);
nor UO_1279 (O_1279,N_14962,N_14996);
xnor UO_1280 (O_1280,N_14991,N_14949);
and UO_1281 (O_1281,N_14983,N_14956);
or UO_1282 (O_1282,N_14932,N_14974);
xor UO_1283 (O_1283,N_14949,N_14926);
xnor UO_1284 (O_1284,N_14990,N_14995);
nor UO_1285 (O_1285,N_14941,N_14910);
nand UO_1286 (O_1286,N_14996,N_14901);
or UO_1287 (O_1287,N_14876,N_14930);
nor UO_1288 (O_1288,N_14935,N_14979);
or UO_1289 (O_1289,N_14937,N_14915);
or UO_1290 (O_1290,N_14875,N_14907);
and UO_1291 (O_1291,N_14970,N_14961);
nand UO_1292 (O_1292,N_14998,N_14976);
xor UO_1293 (O_1293,N_14923,N_14961);
nor UO_1294 (O_1294,N_14891,N_14955);
nor UO_1295 (O_1295,N_14882,N_14904);
nor UO_1296 (O_1296,N_14995,N_14986);
xor UO_1297 (O_1297,N_14894,N_14985);
xnor UO_1298 (O_1298,N_14917,N_14920);
or UO_1299 (O_1299,N_14967,N_14945);
and UO_1300 (O_1300,N_14956,N_14966);
xnor UO_1301 (O_1301,N_14890,N_14983);
nor UO_1302 (O_1302,N_14879,N_14935);
xor UO_1303 (O_1303,N_14910,N_14989);
and UO_1304 (O_1304,N_14915,N_14916);
or UO_1305 (O_1305,N_14949,N_14995);
or UO_1306 (O_1306,N_14925,N_14893);
nor UO_1307 (O_1307,N_14998,N_14978);
nand UO_1308 (O_1308,N_14979,N_14992);
or UO_1309 (O_1309,N_14943,N_14979);
nor UO_1310 (O_1310,N_14892,N_14941);
nand UO_1311 (O_1311,N_14977,N_14920);
or UO_1312 (O_1312,N_14894,N_14924);
nor UO_1313 (O_1313,N_14969,N_14997);
or UO_1314 (O_1314,N_14894,N_14944);
xor UO_1315 (O_1315,N_14895,N_14965);
xor UO_1316 (O_1316,N_14877,N_14977);
nor UO_1317 (O_1317,N_14939,N_14980);
or UO_1318 (O_1318,N_14971,N_14961);
nand UO_1319 (O_1319,N_14899,N_14923);
or UO_1320 (O_1320,N_14947,N_14953);
xor UO_1321 (O_1321,N_14958,N_14887);
and UO_1322 (O_1322,N_14948,N_14973);
and UO_1323 (O_1323,N_14914,N_14915);
xor UO_1324 (O_1324,N_14904,N_14926);
xor UO_1325 (O_1325,N_14966,N_14898);
nand UO_1326 (O_1326,N_14891,N_14967);
or UO_1327 (O_1327,N_14892,N_14928);
nor UO_1328 (O_1328,N_14957,N_14998);
nor UO_1329 (O_1329,N_14938,N_14951);
nand UO_1330 (O_1330,N_14982,N_14891);
xor UO_1331 (O_1331,N_14903,N_14914);
nor UO_1332 (O_1332,N_14909,N_14952);
or UO_1333 (O_1333,N_14937,N_14921);
nor UO_1334 (O_1334,N_14884,N_14906);
xnor UO_1335 (O_1335,N_14988,N_14961);
or UO_1336 (O_1336,N_14970,N_14940);
and UO_1337 (O_1337,N_14949,N_14958);
nand UO_1338 (O_1338,N_14886,N_14986);
xnor UO_1339 (O_1339,N_14984,N_14963);
and UO_1340 (O_1340,N_14959,N_14893);
xor UO_1341 (O_1341,N_14902,N_14967);
nor UO_1342 (O_1342,N_14927,N_14977);
xor UO_1343 (O_1343,N_14880,N_14916);
nand UO_1344 (O_1344,N_14944,N_14938);
and UO_1345 (O_1345,N_14992,N_14937);
nand UO_1346 (O_1346,N_14911,N_14965);
xnor UO_1347 (O_1347,N_14919,N_14883);
nor UO_1348 (O_1348,N_14999,N_14988);
nand UO_1349 (O_1349,N_14956,N_14926);
nor UO_1350 (O_1350,N_14956,N_14980);
nor UO_1351 (O_1351,N_14932,N_14957);
xor UO_1352 (O_1352,N_14919,N_14981);
xnor UO_1353 (O_1353,N_14913,N_14890);
xor UO_1354 (O_1354,N_14981,N_14947);
nand UO_1355 (O_1355,N_14879,N_14928);
or UO_1356 (O_1356,N_14952,N_14943);
nor UO_1357 (O_1357,N_14883,N_14973);
xnor UO_1358 (O_1358,N_14976,N_14947);
xor UO_1359 (O_1359,N_14956,N_14927);
nand UO_1360 (O_1360,N_14936,N_14981);
or UO_1361 (O_1361,N_14962,N_14875);
or UO_1362 (O_1362,N_14978,N_14954);
or UO_1363 (O_1363,N_14915,N_14925);
nand UO_1364 (O_1364,N_14921,N_14923);
nor UO_1365 (O_1365,N_14999,N_14886);
nor UO_1366 (O_1366,N_14961,N_14959);
and UO_1367 (O_1367,N_14877,N_14937);
xnor UO_1368 (O_1368,N_14947,N_14880);
and UO_1369 (O_1369,N_14878,N_14955);
nor UO_1370 (O_1370,N_14985,N_14970);
nand UO_1371 (O_1371,N_14940,N_14961);
xor UO_1372 (O_1372,N_14930,N_14983);
nand UO_1373 (O_1373,N_14958,N_14890);
or UO_1374 (O_1374,N_14956,N_14944);
xnor UO_1375 (O_1375,N_14880,N_14951);
or UO_1376 (O_1376,N_14899,N_14904);
xor UO_1377 (O_1377,N_14963,N_14993);
nand UO_1378 (O_1378,N_14948,N_14947);
xnor UO_1379 (O_1379,N_14924,N_14913);
and UO_1380 (O_1380,N_14894,N_14921);
nand UO_1381 (O_1381,N_14922,N_14926);
and UO_1382 (O_1382,N_14901,N_14878);
xor UO_1383 (O_1383,N_14963,N_14908);
and UO_1384 (O_1384,N_14935,N_14921);
xor UO_1385 (O_1385,N_14912,N_14923);
or UO_1386 (O_1386,N_14920,N_14951);
xnor UO_1387 (O_1387,N_14880,N_14988);
and UO_1388 (O_1388,N_14904,N_14917);
or UO_1389 (O_1389,N_14901,N_14956);
or UO_1390 (O_1390,N_14990,N_14993);
nor UO_1391 (O_1391,N_14967,N_14911);
or UO_1392 (O_1392,N_14963,N_14976);
xnor UO_1393 (O_1393,N_14947,N_14990);
and UO_1394 (O_1394,N_14875,N_14956);
and UO_1395 (O_1395,N_14959,N_14960);
and UO_1396 (O_1396,N_14939,N_14934);
and UO_1397 (O_1397,N_14879,N_14887);
nor UO_1398 (O_1398,N_14947,N_14955);
nand UO_1399 (O_1399,N_14916,N_14983);
nand UO_1400 (O_1400,N_14927,N_14935);
nor UO_1401 (O_1401,N_14973,N_14890);
nand UO_1402 (O_1402,N_14962,N_14924);
xor UO_1403 (O_1403,N_14999,N_14901);
or UO_1404 (O_1404,N_14888,N_14985);
xnor UO_1405 (O_1405,N_14977,N_14972);
and UO_1406 (O_1406,N_14959,N_14968);
or UO_1407 (O_1407,N_14921,N_14896);
nor UO_1408 (O_1408,N_14970,N_14965);
nor UO_1409 (O_1409,N_14941,N_14932);
xnor UO_1410 (O_1410,N_14928,N_14941);
nand UO_1411 (O_1411,N_14955,N_14933);
nand UO_1412 (O_1412,N_14885,N_14926);
nor UO_1413 (O_1413,N_14950,N_14958);
nand UO_1414 (O_1414,N_14933,N_14905);
nand UO_1415 (O_1415,N_14941,N_14956);
and UO_1416 (O_1416,N_14876,N_14881);
nor UO_1417 (O_1417,N_14959,N_14972);
xnor UO_1418 (O_1418,N_14932,N_14969);
or UO_1419 (O_1419,N_14936,N_14940);
or UO_1420 (O_1420,N_14935,N_14956);
or UO_1421 (O_1421,N_14917,N_14975);
and UO_1422 (O_1422,N_14912,N_14929);
nor UO_1423 (O_1423,N_14940,N_14958);
or UO_1424 (O_1424,N_14899,N_14944);
nand UO_1425 (O_1425,N_14998,N_14977);
nand UO_1426 (O_1426,N_14886,N_14916);
nor UO_1427 (O_1427,N_14981,N_14896);
and UO_1428 (O_1428,N_14905,N_14999);
or UO_1429 (O_1429,N_14996,N_14904);
and UO_1430 (O_1430,N_14904,N_14963);
xor UO_1431 (O_1431,N_14881,N_14960);
nand UO_1432 (O_1432,N_14976,N_14955);
xnor UO_1433 (O_1433,N_14991,N_14983);
nor UO_1434 (O_1434,N_14996,N_14879);
nor UO_1435 (O_1435,N_14881,N_14883);
xnor UO_1436 (O_1436,N_14937,N_14930);
xnor UO_1437 (O_1437,N_14936,N_14875);
or UO_1438 (O_1438,N_14882,N_14955);
xor UO_1439 (O_1439,N_14908,N_14974);
nand UO_1440 (O_1440,N_14920,N_14993);
nor UO_1441 (O_1441,N_14918,N_14934);
nor UO_1442 (O_1442,N_14922,N_14982);
and UO_1443 (O_1443,N_14912,N_14934);
and UO_1444 (O_1444,N_14890,N_14936);
xnor UO_1445 (O_1445,N_14948,N_14977);
and UO_1446 (O_1446,N_14938,N_14909);
or UO_1447 (O_1447,N_14887,N_14900);
or UO_1448 (O_1448,N_14943,N_14963);
xor UO_1449 (O_1449,N_14898,N_14923);
or UO_1450 (O_1450,N_14909,N_14879);
and UO_1451 (O_1451,N_14915,N_14882);
nor UO_1452 (O_1452,N_14918,N_14992);
xnor UO_1453 (O_1453,N_14967,N_14934);
xnor UO_1454 (O_1454,N_14996,N_14932);
nand UO_1455 (O_1455,N_14877,N_14945);
and UO_1456 (O_1456,N_14884,N_14939);
xor UO_1457 (O_1457,N_14956,N_14986);
nand UO_1458 (O_1458,N_14995,N_14967);
and UO_1459 (O_1459,N_14895,N_14940);
and UO_1460 (O_1460,N_14978,N_14979);
nand UO_1461 (O_1461,N_14876,N_14938);
nand UO_1462 (O_1462,N_14950,N_14966);
xnor UO_1463 (O_1463,N_14961,N_14969);
xor UO_1464 (O_1464,N_14942,N_14992);
nor UO_1465 (O_1465,N_14954,N_14931);
or UO_1466 (O_1466,N_14893,N_14892);
xor UO_1467 (O_1467,N_14884,N_14936);
nor UO_1468 (O_1468,N_14946,N_14888);
xor UO_1469 (O_1469,N_14997,N_14962);
nand UO_1470 (O_1470,N_14978,N_14907);
or UO_1471 (O_1471,N_14967,N_14926);
or UO_1472 (O_1472,N_14881,N_14925);
xnor UO_1473 (O_1473,N_14989,N_14928);
nand UO_1474 (O_1474,N_14915,N_14876);
nor UO_1475 (O_1475,N_14977,N_14955);
nor UO_1476 (O_1476,N_14981,N_14938);
xor UO_1477 (O_1477,N_14923,N_14946);
xor UO_1478 (O_1478,N_14959,N_14981);
nand UO_1479 (O_1479,N_14887,N_14980);
nor UO_1480 (O_1480,N_14908,N_14987);
and UO_1481 (O_1481,N_14914,N_14964);
nand UO_1482 (O_1482,N_14945,N_14933);
and UO_1483 (O_1483,N_14919,N_14905);
nand UO_1484 (O_1484,N_14952,N_14937);
nor UO_1485 (O_1485,N_14897,N_14880);
xnor UO_1486 (O_1486,N_14900,N_14968);
nor UO_1487 (O_1487,N_14908,N_14915);
nand UO_1488 (O_1488,N_14894,N_14987);
and UO_1489 (O_1489,N_14917,N_14911);
xor UO_1490 (O_1490,N_14885,N_14955);
or UO_1491 (O_1491,N_14962,N_14879);
nand UO_1492 (O_1492,N_14919,N_14977);
or UO_1493 (O_1493,N_14989,N_14883);
nor UO_1494 (O_1494,N_14995,N_14900);
and UO_1495 (O_1495,N_14907,N_14891);
nor UO_1496 (O_1496,N_14902,N_14988);
nand UO_1497 (O_1497,N_14933,N_14912);
xor UO_1498 (O_1498,N_14984,N_14947);
nor UO_1499 (O_1499,N_14902,N_14933);
nand UO_1500 (O_1500,N_14996,N_14957);
and UO_1501 (O_1501,N_14930,N_14956);
and UO_1502 (O_1502,N_14922,N_14946);
nand UO_1503 (O_1503,N_14916,N_14925);
nor UO_1504 (O_1504,N_14923,N_14954);
nor UO_1505 (O_1505,N_14997,N_14957);
nand UO_1506 (O_1506,N_14921,N_14959);
or UO_1507 (O_1507,N_14917,N_14922);
nand UO_1508 (O_1508,N_14959,N_14918);
xor UO_1509 (O_1509,N_14986,N_14938);
nor UO_1510 (O_1510,N_14898,N_14987);
or UO_1511 (O_1511,N_14893,N_14989);
or UO_1512 (O_1512,N_14940,N_14892);
nand UO_1513 (O_1513,N_14877,N_14921);
xnor UO_1514 (O_1514,N_14990,N_14926);
xor UO_1515 (O_1515,N_14990,N_14921);
nand UO_1516 (O_1516,N_14886,N_14920);
xor UO_1517 (O_1517,N_14919,N_14894);
or UO_1518 (O_1518,N_14918,N_14953);
or UO_1519 (O_1519,N_14922,N_14876);
nor UO_1520 (O_1520,N_14887,N_14943);
and UO_1521 (O_1521,N_14924,N_14911);
and UO_1522 (O_1522,N_14888,N_14970);
and UO_1523 (O_1523,N_14906,N_14999);
xnor UO_1524 (O_1524,N_14878,N_14954);
xor UO_1525 (O_1525,N_14991,N_14880);
or UO_1526 (O_1526,N_14881,N_14970);
or UO_1527 (O_1527,N_14892,N_14958);
nand UO_1528 (O_1528,N_14965,N_14950);
xor UO_1529 (O_1529,N_14899,N_14985);
nor UO_1530 (O_1530,N_14941,N_14900);
or UO_1531 (O_1531,N_14907,N_14914);
nor UO_1532 (O_1532,N_14982,N_14987);
nor UO_1533 (O_1533,N_14995,N_14957);
or UO_1534 (O_1534,N_14885,N_14986);
nand UO_1535 (O_1535,N_14957,N_14975);
nand UO_1536 (O_1536,N_14914,N_14937);
nor UO_1537 (O_1537,N_14964,N_14888);
nor UO_1538 (O_1538,N_14954,N_14937);
nand UO_1539 (O_1539,N_14991,N_14974);
xor UO_1540 (O_1540,N_14951,N_14883);
or UO_1541 (O_1541,N_14914,N_14900);
nor UO_1542 (O_1542,N_14997,N_14896);
nor UO_1543 (O_1543,N_14898,N_14949);
or UO_1544 (O_1544,N_14912,N_14884);
nand UO_1545 (O_1545,N_14980,N_14900);
nor UO_1546 (O_1546,N_14915,N_14943);
nor UO_1547 (O_1547,N_14975,N_14923);
or UO_1548 (O_1548,N_14879,N_14940);
nand UO_1549 (O_1549,N_14987,N_14999);
nand UO_1550 (O_1550,N_14902,N_14886);
nand UO_1551 (O_1551,N_14950,N_14909);
nand UO_1552 (O_1552,N_14907,N_14921);
or UO_1553 (O_1553,N_14959,N_14897);
and UO_1554 (O_1554,N_14931,N_14991);
nand UO_1555 (O_1555,N_14996,N_14919);
or UO_1556 (O_1556,N_14928,N_14926);
nor UO_1557 (O_1557,N_14952,N_14970);
nand UO_1558 (O_1558,N_14981,N_14995);
nand UO_1559 (O_1559,N_14924,N_14916);
xnor UO_1560 (O_1560,N_14908,N_14906);
or UO_1561 (O_1561,N_14974,N_14904);
nor UO_1562 (O_1562,N_14998,N_14960);
nor UO_1563 (O_1563,N_14893,N_14970);
or UO_1564 (O_1564,N_14911,N_14897);
xor UO_1565 (O_1565,N_14978,N_14967);
xnor UO_1566 (O_1566,N_14956,N_14893);
and UO_1567 (O_1567,N_14948,N_14965);
and UO_1568 (O_1568,N_14967,N_14954);
nand UO_1569 (O_1569,N_14990,N_14901);
xnor UO_1570 (O_1570,N_14978,N_14904);
or UO_1571 (O_1571,N_14913,N_14906);
nor UO_1572 (O_1572,N_14963,N_14969);
nand UO_1573 (O_1573,N_14891,N_14898);
nand UO_1574 (O_1574,N_14877,N_14959);
nor UO_1575 (O_1575,N_14918,N_14956);
nand UO_1576 (O_1576,N_14889,N_14905);
or UO_1577 (O_1577,N_14967,N_14894);
xor UO_1578 (O_1578,N_14984,N_14983);
and UO_1579 (O_1579,N_14932,N_14936);
or UO_1580 (O_1580,N_14906,N_14876);
and UO_1581 (O_1581,N_14996,N_14951);
and UO_1582 (O_1582,N_14932,N_14978);
nor UO_1583 (O_1583,N_14940,N_14907);
and UO_1584 (O_1584,N_14909,N_14945);
or UO_1585 (O_1585,N_14948,N_14974);
or UO_1586 (O_1586,N_14964,N_14929);
and UO_1587 (O_1587,N_14999,N_14923);
and UO_1588 (O_1588,N_14966,N_14900);
nand UO_1589 (O_1589,N_14951,N_14993);
or UO_1590 (O_1590,N_14969,N_14904);
or UO_1591 (O_1591,N_14910,N_14934);
nand UO_1592 (O_1592,N_14955,N_14990);
xnor UO_1593 (O_1593,N_14957,N_14920);
nand UO_1594 (O_1594,N_14978,N_14911);
and UO_1595 (O_1595,N_14971,N_14933);
or UO_1596 (O_1596,N_14946,N_14990);
and UO_1597 (O_1597,N_14952,N_14939);
and UO_1598 (O_1598,N_14967,N_14983);
and UO_1599 (O_1599,N_14947,N_14989);
and UO_1600 (O_1600,N_14988,N_14944);
xnor UO_1601 (O_1601,N_14909,N_14992);
nor UO_1602 (O_1602,N_14995,N_14975);
nand UO_1603 (O_1603,N_14889,N_14882);
and UO_1604 (O_1604,N_14999,N_14900);
xor UO_1605 (O_1605,N_14945,N_14949);
and UO_1606 (O_1606,N_14876,N_14996);
xor UO_1607 (O_1607,N_14886,N_14919);
and UO_1608 (O_1608,N_14943,N_14896);
xnor UO_1609 (O_1609,N_14886,N_14996);
or UO_1610 (O_1610,N_14973,N_14985);
nand UO_1611 (O_1611,N_14929,N_14919);
or UO_1612 (O_1612,N_14983,N_14962);
and UO_1613 (O_1613,N_14899,N_14960);
xnor UO_1614 (O_1614,N_14919,N_14947);
and UO_1615 (O_1615,N_14962,N_14922);
xnor UO_1616 (O_1616,N_14989,N_14943);
or UO_1617 (O_1617,N_14990,N_14924);
nor UO_1618 (O_1618,N_14883,N_14896);
and UO_1619 (O_1619,N_14950,N_14920);
and UO_1620 (O_1620,N_14878,N_14887);
nor UO_1621 (O_1621,N_14883,N_14877);
nand UO_1622 (O_1622,N_14957,N_14893);
nand UO_1623 (O_1623,N_14879,N_14938);
nor UO_1624 (O_1624,N_14986,N_14950);
xnor UO_1625 (O_1625,N_14939,N_14926);
or UO_1626 (O_1626,N_14988,N_14945);
xnor UO_1627 (O_1627,N_14950,N_14998);
nor UO_1628 (O_1628,N_14924,N_14882);
nor UO_1629 (O_1629,N_14924,N_14884);
xnor UO_1630 (O_1630,N_14981,N_14966);
or UO_1631 (O_1631,N_14943,N_14960);
xnor UO_1632 (O_1632,N_14904,N_14881);
or UO_1633 (O_1633,N_14892,N_14962);
nor UO_1634 (O_1634,N_14999,N_14929);
nand UO_1635 (O_1635,N_14969,N_14877);
and UO_1636 (O_1636,N_14901,N_14937);
and UO_1637 (O_1637,N_14946,N_14878);
and UO_1638 (O_1638,N_14918,N_14893);
xor UO_1639 (O_1639,N_14876,N_14970);
and UO_1640 (O_1640,N_14981,N_14952);
or UO_1641 (O_1641,N_14934,N_14928);
nand UO_1642 (O_1642,N_14954,N_14935);
or UO_1643 (O_1643,N_14952,N_14900);
nand UO_1644 (O_1644,N_14903,N_14900);
or UO_1645 (O_1645,N_14949,N_14940);
and UO_1646 (O_1646,N_14999,N_14976);
nand UO_1647 (O_1647,N_14952,N_14878);
nor UO_1648 (O_1648,N_14921,N_14977);
and UO_1649 (O_1649,N_14931,N_14989);
or UO_1650 (O_1650,N_14916,N_14931);
nor UO_1651 (O_1651,N_14899,N_14921);
xor UO_1652 (O_1652,N_14916,N_14911);
or UO_1653 (O_1653,N_14944,N_14907);
and UO_1654 (O_1654,N_14905,N_14886);
nand UO_1655 (O_1655,N_14979,N_14939);
xor UO_1656 (O_1656,N_14929,N_14915);
nand UO_1657 (O_1657,N_14955,N_14952);
xnor UO_1658 (O_1658,N_14891,N_14925);
nand UO_1659 (O_1659,N_14900,N_14949);
and UO_1660 (O_1660,N_14900,N_14974);
nand UO_1661 (O_1661,N_14911,N_14956);
xnor UO_1662 (O_1662,N_14878,N_14900);
xnor UO_1663 (O_1663,N_14932,N_14946);
and UO_1664 (O_1664,N_14995,N_14974);
nand UO_1665 (O_1665,N_14878,N_14940);
and UO_1666 (O_1666,N_14893,N_14964);
nor UO_1667 (O_1667,N_14903,N_14884);
xor UO_1668 (O_1668,N_14969,N_14897);
or UO_1669 (O_1669,N_14926,N_14951);
nand UO_1670 (O_1670,N_14985,N_14951);
or UO_1671 (O_1671,N_14987,N_14940);
or UO_1672 (O_1672,N_14910,N_14976);
and UO_1673 (O_1673,N_14968,N_14911);
xor UO_1674 (O_1674,N_14915,N_14932);
and UO_1675 (O_1675,N_14938,N_14987);
and UO_1676 (O_1676,N_14885,N_14892);
nand UO_1677 (O_1677,N_14935,N_14902);
nand UO_1678 (O_1678,N_14957,N_14889);
nor UO_1679 (O_1679,N_14948,N_14982);
nor UO_1680 (O_1680,N_14963,N_14966);
xor UO_1681 (O_1681,N_14964,N_14980);
nand UO_1682 (O_1682,N_14955,N_14909);
xor UO_1683 (O_1683,N_14916,N_14902);
xor UO_1684 (O_1684,N_14940,N_14939);
nand UO_1685 (O_1685,N_14957,N_14917);
nand UO_1686 (O_1686,N_14931,N_14922);
xnor UO_1687 (O_1687,N_14929,N_14954);
xor UO_1688 (O_1688,N_14885,N_14956);
nand UO_1689 (O_1689,N_14896,N_14964);
or UO_1690 (O_1690,N_14884,N_14944);
or UO_1691 (O_1691,N_14968,N_14924);
nand UO_1692 (O_1692,N_14888,N_14891);
xnor UO_1693 (O_1693,N_14986,N_14968);
or UO_1694 (O_1694,N_14967,N_14948);
nor UO_1695 (O_1695,N_14917,N_14988);
nor UO_1696 (O_1696,N_14899,N_14953);
xnor UO_1697 (O_1697,N_14886,N_14990);
nor UO_1698 (O_1698,N_14918,N_14967);
or UO_1699 (O_1699,N_14992,N_14945);
nor UO_1700 (O_1700,N_14921,N_14966);
and UO_1701 (O_1701,N_14955,N_14932);
xnor UO_1702 (O_1702,N_14890,N_14950);
or UO_1703 (O_1703,N_14924,N_14892);
and UO_1704 (O_1704,N_14931,N_14884);
nand UO_1705 (O_1705,N_14902,N_14957);
and UO_1706 (O_1706,N_14880,N_14960);
xor UO_1707 (O_1707,N_14968,N_14930);
xnor UO_1708 (O_1708,N_14946,N_14891);
and UO_1709 (O_1709,N_14884,N_14893);
nand UO_1710 (O_1710,N_14933,N_14950);
nand UO_1711 (O_1711,N_14954,N_14972);
and UO_1712 (O_1712,N_14987,N_14922);
or UO_1713 (O_1713,N_14934,N_14947);
xor UO_1714 (O_1714,N_14950,N_14883);
and UO_1715 (O_1715,N_14995,N_14906);
nor UO_1716 (O_1716,N_14893,N_14977);
nor UO_1717 (O_1717,N_14994,N_14995);
or UO_1718 (O_1718,N_14968,N_14957);
nor UO_1719 (O_1719,N_14950,N_14992);
nor UO_1720 (O_1720,N_14967,N_14881);
nand UO_1721 (O_1721,N_14994,N_14991);
or UO_1722 (O_1722,N_14991,N_14990);
nand UO_1723 (O_1723,N_14965,N_14985);
nand UO_1724 (O_1724,N_14960,N_14876);
and UO_1725 (O_1725,N_14885,N_14886);
xnor UO_1726 (O_1726,N_14957,N_14931);
xor UO_1727 (O_1727,N_14951,N_14959);
or UO_1728 (O_1728,N_14930,N_14886);
and UO_1729 (O_1729,N_14877,N_14897);
or UO_1730 (O_1730,N_14974,N_14972);
xnor UO_1731 (O_1731,N_14948,N_14976);
nand UO_1732 (O_1732,N_14975,N_14914);
and UO_1733 (O_1733,N_14930,N_14918);
and UO_1734 (O_1734,N_14903,N_14909);
and UO_1735 (O_1735,N_14918,N_14971);
nand UO_1736 (O_1736,N_14975,N_14942);
or UO_1737 (O_1737,N_14946,N_14965);
and UO_1738 (O_1738,N_14881,N_14905);
xnor UO_1739 (O_1739,N_14995,N_14954);
and UO_1740 (O_1740,N_14970,N_14967);
or UO_1741 (O_1741,N_14986,N_14928);
or UO_1742 (O_1742,N_14932,N_14909);
nand UO_1743 (O_1743,N_14894,N_14952);
xor UO_1744 (O_1744,N_14919,N_14958);
or UO_1745 (O_1745,N_14998,N_14883);
xor UO_1746 (O_1746,N_14875,N_14937);
nor UO_1747 (O_1747,N_14904,N_14981);
and UO_1748 (O_1748,N_14929,N_14967);
xnor UO_1749 (O_1749,N_14891,N_14875);
nor UO_1750 (O_1750,N_14881,N_14948);
nor UO_1751 (O_1751,N_14883,N_14977);
xnor UO_1752 (O_1752,N_14960,N_14989);
or UO_1753 (O_1753,N_14997,N_14963);
or UO_1754 (O_1754,N_14925,N_14981);
nand UO_1755 (O_1755,N_14996,N_14877);
xnor UO_1756 (O_1756,N_14886,N_14946);
nor UO_1757 (O_1757,N_14936,N_14997);
nor UO_1758 (O_1758,N_14970,N_14957);
nor UO_1759 (O_1759,N_14886,N_14954);
nor UO_1760 (O_1760,N_14896,N_14899);
nor UO_1761 (O_1761,N_14983,N_14931);
nand UO_1762 (O_1762,N_14989,N_14921);
xnor UO_1763 (O_1763,N_14987,N_14947);
xor UO_1764 (O_1764,N_14937,N_14942);
and UO_1765 (O_1765,N_14982,N_14888);
nor UO_1766 (O_1766,N_14963,N_14972);
xor UO_1767 (O_1767,N_14936,N_14894);
nor UO_1768 (O_1768,N_14891,N_14894);
nand UO_1769 (O_1769,N_14928,N_14887);
nand UO_1770 (O_1770,N_14971,N_14976);
or UO_1771 (O_1771,N_14961,N_14936);
nor UO_1772 (O_1772,N_14882,N_14894);
or UO_1773 (O_1773,N_14999,N_14919);
or UO_1774 (O_1774,N_14913,N_14995);
or UO_1775 (O_1775,N_14983,N_14906);
or UO_1776 (O_1776,N_14985,N_14900);
nor UO_1777 (O_1777,N_14914,N_14905);
nor UO_1778 (O_1778,N_14909,N_14897);
and UO_1779 (O_1779,N_14884,N_14993);
and UO_1780 (O_1780,N_14923,N_14942);
or UO_1781 (O_1781,N_14983,N_14921);
and UO_1782 (O_1782,N_14912,N_14880);
and UO_1783 (O_1783,N_14891,N_14883);
or UO_1784 (O_1784,N_14921,N_14967);
or UO_1785 (O_1785,N_14881,N_14979);
or UO_1786 (O_1786,N_14885,N_14938);
or UO_1787 (O_1787,N_14959,N_14903);
xnor UO_1788 (O_1788,N_14882,N_14961);
and UO_1789 (O_1789,N_14976,N_14914);
or UO_1790 (O_1790,N_14958,N_14990);
nand UO_1791 (O_1791,N_14939,N_14887);
or UO_1792 (O_1792,N_14935,N_14970);
and UO_1793 (O_1793,N_14907,N_14950);
and UO_1794 (O_1794,N_14955,N_14954);
or UO_1795 (O_1795,N_14976,N_14906);
and UO_1796 (O_1796,N_14961,N_14900);
nor UO_1797 (O_1797,N_14892,N_14922);
and UO_1798 (O_1798,N_14938,N_14892);
nand UO_1799 (O_1799,N_14958,N_14922);
and UO_1800 (O_1800,N_14985,N_14978);
and UO_1801 (O_1801,N_14970,N_14917);
nand UO_1802 (O_1802,N_14965,N_14993);
nand UO_1803 (O_1803,N_14910,N_14877);
or UO_1804 (O_1804,N_14879,N_14998);
or UO_1805 (O_1805,N_14911,N_14877);
or UO_1806 (O_1806,N_14907,N_14895);
and UO_1807 (O_1807,N_14919,N_14899);
or UO_1808 (O_1808,N_14952,N_14986);
xnor UO_1809 (O_1809,N_14945,N_14978);
or UO_1810 (O_1810,N_14889,N_14893);
and UO_1811 (O_1811,N_14936,N_14942);
nor UO_1812 (O_1812,N_14927,N_14991);
nor UO_1813 (O_1813,N_14985,N_14904);
nor UO_1814 (O_1814,N_14935,N_14950);
xor UO_1815 (O_1815,N_14937,N_14943);
nand UO_1816 (O_1816,N_14937,N_14970);
or UO_1817 (O_1817,N_14999,N_14985);
or UO_1818 (O_1818,N_14876,N_14944);
nand UO_1819 (O_1819,N_14959,N_14958);
and UO_1820 (O_1820,N_14959,N_14984);
or UO_1821 (O_1821,N_14881,N_14981);
or UO_1822 (O_1822,N_14890,N_14892);
or UO_1823 (O_1823,N_14970,N_14966);
or UO_1824 (O_1824,N_14975,N_14895);
xor UO_1825 (O_1825,N_14988,N_14974);
or UO_1826 (O_1826,N_14968,N_14961);
or UO_1827 (O_1827,N_14880,N_14961);
or UO_1828 (O_1828,N_14952,N_14919);
and UO_1829 (O_1829,N_14908,N_14991);
xor UO_1830 (O_1830,N_14960,N_14978);
nor UO_1831 (O_1831,N_14990,N_14944);
and UO_1832 (O_1832,N_14910,N_14919);
nand UO_1833 (O_1833,N_14923,N_14993);
nand UO_1834 (O_1834,N_14890,N_14965);
or UO_1835 (O_1835,N_14950,N_14900);
nand UO_1836 (O_1836,N_14998,N_14954);
xnor UO_1837 (O_1837,N_14922,N_14919);
and UO_1838 (O_1838,N_14888,N_14994);
and UO_1839 (O_1839,N_14881,N_14879);
and UO_1840 (O_1840,N_14968,N_14958);
nor UO_1841 (O_1841,N_14902,N_14948);
and UO_1842 (O_1842,N_14887,N_14896);
and UO_1843 (O_1843,N_14969,N_14970);
nor UO_1844 (O_1844,N_14879,N_14934);
or UO_1845 (O_1845,N_14953,N_14945);
xnor UO_1846 (O_1846,N_14961,N_14905);
and UO_1847 (O_1847,N_14902,N_14918);
xnor UO_1848 (O_1848,N_14939,N_14936);
nand UO_1849 (O_1849,N_14952,N_14992);
xnor UO_1850 (O_1850,N_14900,N_14991);
and UO_1851 (O_1851,N_14883,N_14882);
nor UO_1852 (O_1852,N_14982,N_14956);
or UO_1853 (O_1853,N_14985,N_14934);
and UO_1854 (O_1854,N_14927,N_14980);
xnor UO_1855 (O_1855,N_14944,N_14932);
or UO_1856 (O_1856,N_14968,N_14944);
nor UO_1857 (O_1857,N_14915,N_14930);
or UO_1858 (O_1858,N_14961,N_14902);
and UO_1859 (O_1859,N_14897,N_14881);
and UO_1860 (O_1860,N_14961,N_14911);
nand UO_1861 (O_1861,N_14900,N_14930);
nor UO_1862 (O_1862,N_14916,N_14890);
nor UO_1863 (O_1863,N_14951,N_14875);
xor UO_1864 (O_1864,N_14934,N_14962);
and UO_1865 (O_1865,N_14938,N_14931);
nand UO_1866 (O_1866,N_14999,N_14982);
or UO_1867 (O_1867,N_14988,N_14975);
or UO_1868 (O_1868,N_14905,N_14930);
nor UO_1869 (O_1869,N_14933,N_14907);
nor UO_1870 (O_1870,N_14884,N_14937);
or UO_1871 (O_1871,N_14964,N_14951);
xnor UO_1872 (O_1872,N_14907,N_14980);
nand UO_1873 (O_1873,N_14896,N_14928);
or UO_1874 (O_1874,N_14935,N_14946);
or UO_1875 (O_1875,N_14894,N_14955);
xor UO_1876 (O_1876,N_14974,N_14955);
and UO_1877 (O_1877,N_14928,N_14891);
and UO_1878 (O_1878,N_14917,N_14927);
nand UO_1879 (O_1879,N_14898,N_14982);
nor UO_1880 (O_1880,N_14994,N_14883);
and UO_1881 (O_1881,N_14984,N_14918);
nor UO_1882 (O_1882,N_14943,N_14901);
or UO_1883 (O_1883,N_14884,N_14985);
xor UO_1884 (O_1884,N_14925,N_14986);
or UO_1885 (O_1885,N_14993,N_14903);
nor UO_1886 (O_1886,N_14918,N_14943);
or UO_1887 (O_1887,N_14926,N_14880);
nor UO_1888 (O_1888,N_14948,N_14918);
nand UO_1889 (O_1889,N_14963,N_14888);
and UO_1890 (O_1890,N_14894,N_14957);
and UO_1891 (O_1891,N_14958,N_14910);
and UO_1892 (O_1892,N_14907,N_14959);
or UO_1893 (O_1893,N_14966,N_14953);
nand UO_1894 (O_1894,N_14961,N_14916);
nand UO_1895 (O_1895,N_14976,N_14915);
nor UO_1896 (O_1896,N_14898,N_14999);
and UO_1897 (O_1897,N_14968,N_14905);
nand UO_1898 (O_1898,N_14998,N_14956);
nand UO_1899 (O_1899,N_14984,N_14892);
and UO_1900 (O_1900,N_14912,N_14994);
or UO_1901 (O_1901,N_14877,N_14966);
nor UO_1902 (O_1902,N_14943,N_14996);
nor UO_1903 (O_1903,N_14982,N_14885);
or UO_1904 (O_1904,N_14888,N_14949);
xnor UO_1905 (O_1905,N_14949,N_14968);
nor UO_1906 (O_1906,N_14981,N_14883);
xnor UO_1907 (O_1907,N_14985,N_14995);
and UO_1908 (O_1908,N_14916,N_14930);
nor UO_1909 (O_1909,N_14957,N_14927);
nor UO_1910 (O_1910,N_14941,N_14995);
xor UO_1911 (O_1911,N_14927,N_14903);
or UO_1912 (O_1912,N_14888,N_14980);
and UO_1913 (O_1913,N_14948,N_14955);
or UO_1914 (O_1914,N_14939,N_14954);
nand UO_1915 (O_1915,N_14942,N_14932);
xor UO_1916 (O_1916,N_14950,N_14995);
xor UO_1917 (O_1917,N_14925,N_14875);
nand UO_1918 (O_1918,N_14924,N_14935);
xnor UO_1919 (O_1919,N_14879,N_14911);
nand UO_1920 (O_1920,N_14966,N_14902);
nor UO_1921 (O_1921,N_14965,N_14983);
or UO_1922 (O_1922,N_14947,N_14878);
and UO_1923 (O_1923,N_14957,N_14936);
xnor UO_1924 (O_1924,N_14969,N_14906);
nor UO_1925 (O_1925,N_14975,N_14939);
nor UO_1926 (O_1926,N_14971,N_14965);
xnor UO_1927 (O_1927,N_14925,N_14928);
and UO_1928 (O_1928,N_14889,N_14968);
nor UO_1929 (O_1929,N_14992,N_14955);
and UO_1930 (O_1930,N_14885,N_14907);
nand UO_1931 (O_1931,N_14876,N_14894);
nor UO_1932 (O_1932,N_14927,N_14944);
nand UO_1933 (O_1933,N_14972,N_14908);
and UO_1934 (O_1934,N_14900,N_14954);
xnor UO_1935 (O_1935,N_14920,N_14900);
nor UO_1936 (O_1936,N_14970,N_14890);
xnor UO_1937 (O_1937,N_14946,N_14993);
and UO_1938 (O_1938,N_14885,N_14882);
nor UO_1939 (O_1939,N_14995,N_14894);
nor UO_1940 (O_1940,N_14941,N_14937);
and UO_1941 (O_1941,N_14977,N_14987);
nand UO_1942 (O_1942,N_14988,N_14923);
and UO_1943 (O_1943,N_14911,N_14901);
or UO_1944 (O_1944,N_14919,N_14991);
nand UO_1945 (O_1945,N_14959,N_14926);
nand UO_1946 (O_1946,N_14883,N_14884);
nor UO_1947 (O_1947,N_14931,N_14887);
and UO_1948 (O_1948,N_14893,N_14909);
nor UO_1949 (O_1949,N_14910,N_14979);
xnor UO_1950 (O_1950,N_14983,N_14994);
and UO_1951 (O_1951,N_14979,N_14923);
and UO_1952 (O_1952,N_14980,N_14928);
nor UO_1953 (O_1953,N_14900,N_14962);
nor UO_1954 (O_1954,N_14997,N_14996);
nand UO_1955 (O_1955,N_14999,N_14962);
or UO_1956 (O_1956,N_14976,N_14987);
nor UO_1957 (O_1957,N_14969,N_14964);
or UO_1958 (O_1958,N_14986,N_14951);
and UO_1959 (O_1959,N_14931,N_14940);
nor UO_1960 (O_1960,N_14902,N_14879);
or UO_1961 (O_1961,N_14889,N_14879);
nor UO_1962 (O_1962,N_14894,N_14920);
xor UO_1963 (O_1963,N_14984,N_14940);
xnor UO_1964 (O_1964,N_14956,N_14906);
or UO_1965 (O_1965,N_14954,N_14889);
nor UO_1966 (O_1966,N_14911,N_14908);
nor UO_1967 (O_1967,N_14940,N_14983);
or UO_1968 (O_1968,N_14973,N_14945);
nand UO_1969 (O_1969,N_14922,N_14906);
xnor UO_1970 (O_1970,N_14969,N_14920);
nor UO_1971 (O_1971,N_14979,N_14974);
xor UO_1972 (O_1972,N_14898,N_14910);
xnor UO_1973 (O_1973,N_14953,N_14954);
and UO_1974 (O_1974,N_14976,N_14942);
nor UO_1975 (O_1975,N_14910,N_14987);
nor UO_1976 (O_1976,N_14919,N_14943);
or UO_1977 (O_1977,N_14990,N_14878);
or UO_1978 (O_1978,N_14982,N_14890);
or UO_1979 (O_1979,N_14939,N_14964);
nor UO_1980 (O_1980,N_14998,N_14952);
nand UO_1981 (O_1981,N_14938,N_14922);
nor UO_1982 (O_1982,N_14988,N_14925);
and UO_1983 (O_1983,N_14932,N_14994);
nor UO_1984 (O_1984,N_14990,N_14887);
xnor UO_1985 (O_1985,N_14896,N_14944);
nand UO_1986 (O_1986,N_14966,N_14876);
and UO_1987 (O_1987,N_14977,N_14904);
or UO_1988 (O_1988,N_14937,N_14997);
and UO_1989 (O_1989,N_14968,N_14951);
or UO_1990 (O_1990,N_14927,N_14910);
nor UO_1991 (O_1991,N_14934,N_14906);
or UO_1992 (O_1992,N_14969,N_14948);
xor UO_1993 (O_1993,N_14901,N_14893);
or UO_1994 (O_1994,N_14975,N_14974);
xor UO_1995 (O_1995,N_14967,N_14957);
xnor UO_1996 (O_1996,N_14889,N_14956);
xor UO_1997 (O_1997,N_14928,N_14884);
or UO_1998 (O_1998,N_14903,N_14935);
xor UO_1999 (O_1999,N_14993,N_14932);
endmodule