module basic_750_5000_1000_50_levels_2xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
and U0 (N_0,In_473,In_327);
nand U1 (N_1,In_262,In_730);
or U2 (N_2,In_412,In_352);
and U3 (N_3,In_388,In_711);
or U4 (N_4,In_384,In_715);
nand U5 (N_5,In_84,In_54);
xor U6 (N_6,In_496,In_680);
nand U7 (N_7,In_230,In_266);
nor U8 (N_8,In_56,In_294);
or U9 (N_9,In_96,In_251);
nor U10 (N_10,In_426,In_374);
nor U11 (N_11,In_112,In_149);
or U12 (N_12,In_695,In_623);
and U13 (N_13,In_539,In_127);
and U14 (N_14,In_3,In_208);
nor U15 (N_15,In_318,In_47);
nand U16 (N_16,In_238,In_583);
and U17 (N_17,In_261,In_9);
nand U18 (N_18,In_717,In_351);
or U19 (N_19,In_236,In_228);
nor U20 (N_20,In_507,In_105);
and U21 (N_21,In_706,In_661);
or U22 (N_22,In_551,In_687);
nand U23 (N_23,In_283,In_281);
and U24 (N_24,In_296,In_285);
nor U25 (N_25,In_381,In_182);
nand U26 (N_26,In_137,In_532);
or U27 (N_27,In_650,In_557);
nor U28 (N_28,In_475,In_91);
nor U29 (N_29,In_253,In_494);
and U30 (N_30,In_274,In_598);
or U31 (N_31,In_187,In_93);
and U32 (N_32,In_134,In_663);
or U33 (N_33,In_447,In_631);
and U34 (N_34,In_737,In_684);
or U35 (N_35,In_662,In_647);
or U36 (N_36,In_470,In_39);
and U37 (N_37,In_75,In_309);
nor U38 (N_38,In_368,In_406);
nor U39 (N_39,In_728,In_697);
nand U40 (N_40,In_659,In_584);
or U41 (N_41,In_122,In_675);
or U42 (N_42,In_104,In_257);
nand U43 (N_43,In_245,In_652);
or U44 (N_44,In_171,In_682);
nand U45 (N_45,In_702,In_548);
nand U46 (N_46,In_59,In_355);
nor U47 (N_47,In_681,In_674);
and U48 (N_48,In_32,In_546);
nor U49 (N_49,In_567,In_461);
nor U50 (N_50,In_547,In_160);
or U51 (N_51,In_608,In_118);
nor U52 (N_52,In_341,In_704);
nor U53 (N_53,In_272,In_747);
and U54 (N_54,In_424,In_739);
nand U55 (N_55,In_568,In_367);
xor U56 (N_56,In_648,In_657);
nor U57 (N_57,In_1,In_30);
or U58 (N_58,In_499,In_535);
nand U59 (N_59,In_521,In_353);
or U60 (N_60,In_577,In_326);
or U61 (N_61,In_52,In_218);
or U62 (N_62,In_8,In_375);
nor U63 (N_63,In_17,In_502);
nand U64 (N_64,In_354,In_265);
nand U65 (N_65,In_254,In_308);
nor U66 (N_66,In_313,In_175);
and U67 (N_67,In_744,In_268);
xor U68 (N_68,In_78,In_94);
or U69 (N_69,In_206,In_544);
nor U70 (N_70,In_537,In_64);
or U71 (N_71,In_13,In_370);
nor U72 (N_72,In_333,In_701);
nor U73 (N_73,In_242,In_414);
nand U74 (N_74,In_128,In_685);
or U75 (N_75,In_348,In_106);
and U76 (N_76,In_627,In_514);
nor U77 (N_77,In_22,In_220);
nor U78 (N_78,In_305,In_436);
nor U79 (N_79,In_234,In_519);
nor U80 (N_80,In_88,In_154);
nand U81 (N_81,In_655,In_58);
and U82 (N_82,In_481,In_85);
nand U83 (N_83,In_362,In_497);
or U84 (N_84,In_376,In_530);
xnor U85 (N_85,In_562,In_307);
or U86 (N_86,In_738,In_511);
and U87 (N_87,In_269,In_212);
nand U88 (N_88,In_329,In_536);
nand U89 (N_89,In_637,In_332);
or U90 (N_90,In_203,In_732);
or U91 (N_91,In_231,In_724);
and U92 (N_92,In_446,In_714);
nor U93 (N_93,In_45,In_19);
and U94 (N_94,In_700,In_144);
nor U95 (N_95,In_81,In_259);
or U96 (N_96,In_735,In_334);
nor U97 (N_97,In_719,In_188);
nand U98 (N_98,In_31,In_115);
nor U99 (N_99,In_382,In_450);
nor U100 (N_100,In_435,In_18);
nand U101 (N_101,In_428,In_438);
nor U102 (N_102,In_72,In_491);
nor U103 (N_103,In_696,In_713);
and U104 (N_104,In_71,In_552);
or U105 (N_105,In_99,In_44);
nand U106 (N_106,In_397,In_310);
nand U107 (N_107,In_559,In_503);
or U108 (N_108,In_545,In_12);
or U109 (N_109,In_596,In_26);
or U110 (N_110,In_664,In_169);
nand U111 (N_111,In_191,In_315);
nor U112 (N_112,In_364,In_574);
nor U113 (N_113,In_512,N_71);
nor U114 (N_114,In_540,In_404);
nor U115 (N_115,In_459,In_145);
and U116 (N_116,In_600,In_287);
xnor U117 (N_117,In_566,In_138);
or U118 (N_118,In_229,In_194);
or U119 (N_119,N_81,In_217);
nand U120 (N_120,In_418,In_179);
nor U121 (N_121,In_90,In_727);
and U122 (N_122,In_27,In_526);
nand U123 (N_123,In_692,N_91);
or U124 (N_124,In_184,In_410);
nor U125 (N_125,N_1,In_298);
nor U126 (N_126,In_79,In_746);
and U127 (N_127,In_485,In_299);
or U128 (N_128,In_226,In_133);
xor U129 (N_129,In_304,In_195);
nand U130 (N_130,In_603,In_135);
nand U131 (N_131,In_158,In_394);
or U132 (N_132,N_50,In_156);
nor U133 (N_133,In_89,In_634);
nand U134 (N_134,In_189,In_660);
or U135 (N_135,In_162,In_103);
or U136 (N_136,In_716,N_77);
nand U137 (N_137,N_79,N_8);
and U138 (N_138,In_143,In_139);
nand U139 (N_139,In_508,In_462);
nor U140 (N_140,In_455,In_369);
nor U141 (N_141,In_98,In_466);
nand U142 (N_142,In_431,N_57);
nand U143 (N_143,In_300,In_258);
nand U144 (N_144,N_90,N_69);
nand U145 (N_145,In_672,In_155);
nor U146 (N_146,In_34,In_87);
and U147 (N_147,In_55,In_642);
nand U148 (N_148,In_407,In_534);
nor U149 (N_149,In_482,In_250);
and U150 (N_150,In_358,In_211);
nand U151 (N_151,N_21,In_319);
nor U152 (N_152,In_159,N_59);
nor U153 (N_153,N_20,In_51);
or U154 (N_154,In_243,In_301);
and U155 (N_155,In_60,In_606);
or U156 (N_156,In_282,In_177);
nor U157 (N_157,In_399,In_342);
nor U158 (N_158,In_213,In_669);
nand U159 (N_159,N_34,In_325);
or U160 (N_160,In_43,In_323);
or U161 (N_161,N_99,N_66);
nand U162 (N_162,N_70,In_553);
or U163 (N_163,In_260,N_58);
or U164 (N_164,N_14,In_723);
nand U165 (N_165,In_201,In_641);
or U166 (N_166,In_338,In_693);
and U167 (N_167,In_560,In_237);
xnor U168 (N_168,In_136,In_40);
nor U169 (N_169,In_186,In_667);
and U170 (N_170,In_378,In_252);
and U171 (N_171,In_20,In_405);
or U172 (N_172,In_620,In_501);
nand U173 (N_173,In_564,In_518);
nor U174 (N_174,In_288,In_267);
or U175 (N_175,In_6,N_41);
nand U176 (N_176,N_35,In_76);
and U177 (N_177,In_232,In_277);
nor U178 (N_178,In_176,N_75);
xor U179 (N_179,N_23,In_63);
and U180 (N_180,In_463,In_644);
nor U181 (N_181,N_80,In_690);
nand U182 (N_182,In_82,In_581);
nor U183 (N_183,In_411,In_636);
nor U184 (N_184,In_357,In_689);
nor U185 (N_185,In_726,N_19);
and U186 (N_186,N_11,In_400);
xor U187 (N_187,In_359,In_164);
xor U188 (N_188,In_50,In_556);
or U189 (N_189,N_46,In_522);
nor U190 (N_190,In_295,In_233);
xor U191 (N_191,In_586,In_247);
or U192 (N_192,In_500,In_453);
nor U193 (N_193,In_597,In_484);
nor U194 (N_194,N_85,In_542);
nor U195 (N_195,In_671,In_677);
nand U196 (N_196,In_588,In_227);
xnor U197 (N_197,In_256,In_83);
and U198 (N_198,In_360,In_246);
and U199 (N_199,N_13,In_477);
or U200 (N_200,N_167,In_422);
and U201 (N_201,In_490,In_209);
nor U202 (N_202,In_74,In_616);
and U203 (N_203,In_569,In_0);
or U204 (N_204,In_28,In_293);
nand U205 (N_205,In_224,N_181);
nand U206 (N_206,In_244,In_488);
nand U207 (N_207,In_621,In_14);
nor U208 (N_208,N_125,In_480);
nor U209 (N_209,In_114,N_160);
and U210 (N_210,In_688,In_38);
and U211 (N_211,In_330,In_452);
and U212 (N_212,In_423,In_415);
or U213 (N_213,In_699,In_36);
or U214 (N_214,In_457,In_205);
xor U215 (N_215,In_167,In_125);
and U216 (N_216,In_361,In_53);
and U217 (N_217,N_130,In_192);
or U218 (N_218,N_171,In_70);
nand U219 (N_219,In_168,In_345);
or U220 (N_220,In_95,N_139);
nand U221 (N_221,In_151,In_392);
nor U222 (N_222,N_26,In_391);
and U223 (N_223,N_131,N_56);
or U224 (N_224,In_193,In_386);
xnor U225 (N_225,N_37,N_127);
nand U226 (N_226,In_132,In_339);
xor U227 (N_227,In_401,N_141);
nand U228 (N_228,N_152,In_336);
or U229 (N_229,In_486,In_207);
nor U230 (N_230,In_430,In_441);
and U231 (N_231,In_694,N_117);
or U232 (N_232,In_601,N_119);
nand U233 (N_233,In_23,In_183);
or U234 (N_234,In_73,In_248);
nor U235 (N_235,In_742,In_42);
or U236 (N_236,In_311,In_582);
and U237 (N_237,In_347,In_276);
nor U238 (N_238,N_96,In_487);
and U239 (N_239,N_116,N_126);
nor U240 (N_240,N_101,In_204);
and U241 (N_241,In_395,In_185);
nand U242 (N_242,N_38,N_49);
and U243 (N_243,N_142,N_42);
nor U244 (N_244,In_492,In_541);
or U245 (N_245,In_77,In_617);
nand U246 (N_246,In_673,N_166);
or U247 (N_247,In_614,In_421);
nand U248 (N_248,In_445,In_222);
nor U249 (N_249,In_736,N_65);
nand U250 (N_250,N_45,In_398);
and U251 (N_251,In_721,In_147);
nor U252 (N_252,In_196,N_169);
or U253 (N_253,N_29,In_474);
nor U254 (N_254,N_172,In_123);
or U255 (N_255,In_613,In_712);
nand U256 (N_256,In_314,In_214);
and U257 (N_257,In_61,In_380);
and U258 (N_258,In_478,In_202);
or U259 (N_259,N_118,In_385);
nand U260 (N_260,In_312,In_420);
and U261 (N_261,In_725,In_350);
and U262 (N_262,N_121,In_278);
and U263 (N_263,In_297,In_303);
nand U264 (N_264,In_456,N_173);
or U265 (N_265,N_165,In_622);
and U266 (N_266,N_148,In_29);
and U267 (N_267,In_174,In_146);
and U268 (N_268,In_324,In_656);
or U269 (N_269,N_18,In_589);
nor U270 (N_270,In_396,In_126);
nor U271 (N_271,N_193,In_483);
nor U272 (N_272,In_2,In_571);
nand U273 (N_273,In_594,In_591);
or U274 (N_274,In_538,N_196);
nand U275 (N_275,N_25,In_528);
or U276 (N_276,In_383,In_554);
nand U277 (N_277,In_745,N_140);
and U278 (N_278,In_340,N_187);
and U279 (N_279,In_280,In_679);
and U280 (N_280,In_219,N_109);
nor U281 (N_281,In_172,In_654);
nor U282 (N_282,In_109,In_121);
or U283 (N_283,In_469,In_249);
xnor U284 (N_284,N_10,In_170);
nor U285 (N_285,N_157,In_624);
or U286 (N_286,In_604,N_155);
or U287 (N_287,In_565,In_615);
nor U288 (N_288,N_191,In_264);
or U289 (N_289,In_629,In_416);
and U290 (N_290,In_199,In_638);
xnor U291 (N_291,In_523,In_216);
nor U292 (N_292,N_12,In_402);
or U293 (N_293,In_417,In_97);
nand U294 (N_294,N_82,In_49);
and U295 (N_295,In_197,In_190);
or U296 (N_296,In_157,In_449);
or U297 (N_297,In_433,In_549);
nor U298 (N_298,In_729,In_460);
nand U299 (N_299,In_467,N_176);
nand U300 (N_300,N_195,N_224);
or U301 (N_301,In_676,In_708);
nor U302 (N_302,In_68,In_377);
nand U303 (N_303,N_282,N_55);
and U304 (N_304,N_164,N_104);
nand U305 (N_305,In_612,N_73);
nor U306 (N_306,In_639,N_103);
and U307 (N_307,N_245,In_645);
or U308 (N_308,In_320,In_221);
nor U309 (N_309,N_184,N_183);
nor U310 (N_310,N_235,N_286);
nor U311 (N_311,N_260,In_148);
or U312 (N_312,In_741,N_27);
and U313 (N_313,N_72,In_322);
and U314 (N_314,In_150,N_237);
nand U315 (N_315,N_163,In_198);
nor U316 (N_316,In_665,N_253);
or U317 (N_317,In_640,In_271);
nor U318 (N_318,N_92,N_52);
nand U319 (N_319,In_578,In_344);
nor U320 (N_320,In_107,In_678);
nor U321 (N_321,In_670,N_15);
or U322 (N_322,In_510,N_146);
nor U323 (N_323,N_133,In_579);
and U324 (N_324,In_493,N_158);
nand U325 (N_325,In_722,N_230);
nor U326 (N_326,N_98,N_194);
or U327 (N_327,N_87,In_709);
nor U328 (N_328,N_257,In_210);
and U329 (N_329,In_572,In_442);
nor U330 (N_330,In_16,N_264);
or U331 (N_331,N_262,In_111);
or U332 (N_332,In_46,In_163);
nor U333 (N_333,In_513,N_234);
and U334 (N_334,In_524,In_102);
nand U335 (N_335,In_720,N_68);
nor U336 (N_336,N_277,N_203);
nor U337 (N_337,N_272,N_170);
nand U338 (N_338,N_24,N_251);
and U339 (N_339,N_281,N_47);
or U340 (N_340,In_550,In_215);
nand U341 (N_341,N_283,In_279);
or U342 (N_342,In_718,N_226);
nor U343 (N_343,N_132,In_129);
or U344 (N_344,N_280,N_239);
and U345 (N_345,N_84,In_451);
nand U346 (N_346,In_240,N_124);
or U347 (N_347,In_292,N_243);
nor U348 (N_348,N_174,In_335);
or U349 (N_349,In_328,N_95);
or U350 (N_350,In_625,In_471);
nor U351 (N_351,N_108,N_178);
xor U352 (N_352,In_563,In_707);
or U353 (N_353,In_611,In_101);
nor U354 (N_354,In_703,N_274);
nand U355 (N_355,In_113,In_57);
nand U356 (N_356,N_32,N_151);
nor U357 (N_357,N_210,N_89);
nor U358 (N_358,In_80,N_211);
nor U359 (N_359,N_93,N_259);
and U360 (N_360,In_15,In_387);
nand U361 (N_361,In_4,N_159);
and U362 (N_362,N_292,N_223);
xnor U363 (N_363,In_605,N_36);
nor U364 (N_364,In_626,In_587);
nand U365 (N_365,In_454,N_175);
nor U366 (N_366,In_69,In_585);
or U367 (N_367,In_11,N_112);
or U368 (N_368,N_199,In_200);
or U369 (N_369,In_289,In_165);
nor U370 (N_370,In_363,N_273);
nand U371 (N_371,In_686,N_252);
or U372 (N_372,In_425,In_413);
and U373 (N_373,In_643,N_214);
and U374 (N_374,N_30,In_740);
or U375 (N_375,In_291,In_25);
and U376 (N_376,N_122,In_349);
or U377 (N_377,N_28,N_44);
nor U378 (N_378,N_238,N_61);
or U379 (N_379,In_468,In_517);
nand U380 (N_380,N_299,In_284);
nand U381 (N_381,N_220,N_231);
nor U382 (N_382,N_217,N_6);
and U383 (N_383,N_107,N_275);
nor U384 (N_384,N_51,N_48);
nor U385 (N_385,In_543,In_630);
or U386 (N_386,N_247,In_365);
or U387 (N_387,N_17,N_31);
nor U388 (N_388,In_108,N_9);
and U389 (N_389,In_633,In_607);
and U390 (N_390,In_161,In_62);
nor U391 (N_391,N_145,In_748);
or U392 (N_392,N_111,In_427);
nand U393 (N_393,In_575,In_346);
nand U394 (N_394,In_152,N_254);
nand U395 (N_395,In_316,N_106);
or U396 (N_396,In_389,In_476);
nand U397 (N_397,N_295,N_94);
nor U398 (N_398,N_120,N_78);
nand U399 (N_399,N_154,N_213);
and U400 (N_400,In_628,N_105);
or U401 (N_401,N_215,N_137);
nand U402 (N_402,N_385,In_263);
and U403 (N_403,N_209,In_618);
nor U404 (N_404,In_683,In_731);
and U405 (N_405,In_653,N_391);
nor U406 (N_406,N_261,In_131);
nor U407 (N_407,In_649,In_472);
nor U408 (N_408,In_239,In_124);
nand U409 (N_409,In_698,N_135);
or U410 (N_410,N_325,N_369);
and U411 (N_411,In_33,N_216);
nand U412 (N_412,N_180,N_394);
and U413 (N_413,N_343,N_22);
nor U414 (N_414,In_448,N_134);
and U415 (N_415,N_289,N_156);
or U416 (N_416,N_360,N_138);
and U417 (N_417,In_140,N_39);
or U418 (N_418,N_316,N_123);
nand U419 (N_419,In_65,In_173);
or U420 (N_420,N_387,In_7);
nand U421 (N_421,In_529,N_374);
or U422 (N_422,In_658,N_97);
nand U423 (N_423,N_315,N_4);
and U424 (N_424,In_635,N_86);
nand U425 (N_425,In_506,N_361);
and U426 (N_426,In_743,N_182);
nand U427 (N_427,N_60,In_302);
or U428 (N_428,In_592,N_185);
nand U429 (N_429,In_86,N_329);
nand U430 (N_430,N_392,N_268);
nor U431 (N_431,In_24,In_439);
and U432 (N_432,In_178,In_181);
nor U433 (N_433,In_595,N_205);
nor U434 (N_434,N_354,N_53);
or U435 (N_435,N_302,N_186);
nor U436 (N_436,N_357,N_389);
and U437 (N_437,N_296,N_340);
and U438 (N_438,N_320,N_143);
and U439 (N_439,In_440,In_130);
xnor U440 (N_440,In_666,N_168);
nand U441 (N_441,In_520,In_10);
and U442 (N_442,N_240,N_284);
nand U443 (N_443,N_294,N_149);
and U444 (N_444,N_388,N_372);
nor U445 (N_445,In_580,N_352);
nand U446 (N_446,N_246,N_3);
nor U447 (N_447,N_212,N_276);
xor U448 (N_448,In_734,N_248);
nand U449 (N_449,In_505,N_335);
or U450 (N_450,N_128,In_691);
nand U451 (N_451,N_144,N_342);
nand U452 (N_452,In_444,N_229);
or U453 (N_453,In_180,In_5);
nand U454 (N_454,N_0,N_386);
and U455 (N_455,In_41,N_74);
xnor U456 (N_456,N_378,N_221);
nand U457 (N_457,N_312,N_227);
or U458 (N_458,N_395,N_313);
nand U459 (N_459,N_338,N_16);
nand U460 (N_460,In_570,In_437);
nand U461 (N_461,N_114,N_397);
nor U462 (N_462,N_62,N_298);
or U463 (N_463,N_54,N_332);
and U464 (N_464,N_305,In_142);
nor U465 (N_465,N_236,N_207);
and U466 (N_466,In_504,N_337);
and U467 (N_467,In_393,In_531);
or U468 (N_468,N_301,In_479);
nor U469 (N_469,N_265,N_300);
nand U470 (N_470,N_365,In_465);
or U471 (N_471,N_189,N_304);
or U472 (N_472,N_390,In_458);
or U473 (N_473,N_303,In_525);
and U474 (N_474,In_646,In_379);
nand U475 (N_475,In_366,N_375);
nor U476 (N_476,In_403,N_258);
nand U477 (N_477,N_308,N_76);
and U478 (N_478,In_495,N_310);
nor U479 (N_479,In_619,In_373);
xnor U480 (N_480,In_733,N_250);
and U481 (N_481,N_370,N_198);
and U482 (N_482,In_390,In_489);
and U483 (N_483,N_83,N_355);
or U484 (N_484,In_337,In_225);
and U485 (N_485,N_88,N_366);
nor U486 (N_486,In_255,N_347);
and U487 (N_487,In_576,N_317);
nand U488 (N_488,N_242,N_314);
nand U489 (N_489,N_244,In_593);
nand U490 (N_490,N_271,In_434);
nor U491 (N_491,N_269,N_222);
or U492 (N_492,N_373,N_381);
nor U493 (N_493,In_408,N_345);
and U494 (N_494,In_141,N_399);
or U495 (N_495,N_331,N_318);
nand U496 (N_496,In_555,N_256);
or U497 (N_497,N_364,N_344);
and U498 (N_498,N_197,In_515);
and U499 (N_499,N_241,In_432);
or U500 (N_500,In_498,In_749);
nand U501 (N_501,In_100,In_117);
xor U502 (N_502,N_287,N_288);
and U503 (N_503,N_377,N_263);
nand U504 (N_504,N_356,N_454);
and U505 (N_505,N_327,N_228);
and U506 (N_506,N_418,N_279);
nand U507 (N_507,N_492,N_450);
nor U508 (N_508,N_225,N_417);
nand U509 (N_509,In_321,N_147);
nand U510 (N_510,N_497,N_465);
or U511 (N_511,In_67,In_286);
xor U512 (N_512,N_192,N_434);
xor U513 (N_513,N_136,N_477);
xor U514 (N_514,N_188,In_120);
or U515 (N_515,In_275,N_179);
or U516 (N_516,N_306,N_333);
and U517 (N_517,N_416,N_443);
nor U518 (N_518,N_384,N_328);
nand U519 (N_519,N_398,In_119);
xor U520 (N_520,N_309,In_527);
and U521 (N_521,N_404,N_446);
or U522 (N_522,N_452,N_115);
and U523 (N_523,N_150,N_379);
and U524 (N_524,N_311,N_7);
nor U525 (N_525,In_343,In_116);
nor U526 (N_526,N_421,N_480);
and U527 (N_527,N_432,N_349);
and U528 (N_528,N_419,N_113);
nor U529 (N_529,In_610,In_372);
or U530 (N_530,In_561,N_449);
and U531 (N_531,N_440,In_331);
nor U532 (N_532,N_322,N_346);
nand U533 (N_533,N_376,In_273);
and U534 (N_534,N_359,N_267);
nor U535 (N_535,N_491,N_350);
and U536 (N_536,N_218,In_573);
or U537 (N_537,N_401,In_153);
or U538 (N_538,N_479,N_202);
and U539 (N_539,N_490,N_436);
nor U540 (N_540,In_509,N_368);
nand U541 (N_541,N_430,N_472);
nand U542 (N_542,N_43,N_473);
nand U543 (N_543,N_439,N_307);
and U544 (N_544,N_424,N_423);
or U545 (N_545,N_362,N_400);
and U546 (N_546,N_441,In_705);
and U547 (N_547,In_429,In_241);
nand U548 (N_548,In_602,N_433);
nor U549 (N_549,N_468,In_609);
nor U550 (N_550,N_407,N_5);
or U551 (N_551,N_40,N_448);
nand U552 (N_552,N_499,N_422);
nand U553 (N_553,N_285,N_319);
nor U554 (N_554,N_481,N_153);
or U555 (N_555,N_429,N_478);
nand U556 (N_556,In_37,In_66);
nor U557 (N_557,N_129,N_371);
or U558 (N_558,N_467,In_419);
and U559 (N_559,In_590,N_474);
and U560 (N_560,N_482,N_380);
nand U561 (N_561,N_498,N_334);
nor U562 (N_562,N_270,N_382);
or U563 (N_563,N_496,N_326);
nor U564 (N_564,N_455,N_201);
or U565 (N_565,In_651,N_470);
nand U566 (N_566,N_396,In_223);
and U567 (N_567,N_321,N_412);
nand U568 (N_568,N_451,In_35);
or U569 (N_569,In_533,In_409);
or U570 (N_570,N_367,N_464);
or U571 (N_571,N_484,N_393);
and U572 (N_572,N_495,N_291);
nor U573 (N_573,In_516,In_21);
or U574 (N_574,N_459,In_166);
nand U575 (N_575,N_339,N_100);
and U576 (N_576,N_431,N_204);
and U577 (N_577,N_488,N_348);
nand U578 (N_578,N_405,N_290);
nor U579 (N_579,N_445,N_249);
or U580 (N_580,N_447,N_457);
or U581 (N_581,N_402,In_599);
and U582 (N_582,N_33,N_410);
or U583 (N_583,In_235,N_493);
or U584 (N_584,N_428,In_668);
nand U585 (N_585,N_278,N_444);
nor U586 (N_586,N_266,N_475);
nand U587 (N_587,N_190,N_442);
and U588 (N_588,N_200,N_426);
nor U589 (N_589,N_161,N_453);
and U590 (N_590,In_443,N_2);
nand U591 (N_591,N_219,N_358);
nor U592 (N_592,In_48,N_323);
nor U593 (N_593,N_487,N_64);
nor U594 (N_594,N_456,N_476);
nand U595 (N_595,N_363,N_489);
and U596 (N_596,In_317,N_463);
and U597 (N_597,N_353,N_206);
or U598 (N_598,N_483,N_336);
xnor U599 (N_599,N_461,N_324);
nand U600 (N_600,N_415,N_566);
or U601 (N_601,N_510,N_297);
or U602 (N_602,In_110,N_528);
or U603 (N_603,N_514,N_588);
nand U604 (N_604,In_710,N_571);
and U605 (N_605,N_513,In_371);
nand U606 (N_606,In_464,N_177);
nand U607 (N_607,N_589,N_537);
nand U608 (N_608,N_504,N_466);
nor U609 (N_609,N_383,N_538);
nand U610 (N_610,N_560,N_554);
nor U611 (N_611,N_293,N_505);
or U612 (N_612,N_420,N_437);
and U613 (N_613,N_435,N_547);
or U614 (N_614,In_92,N_579);
and U615 (N_615,N_507,N_585);
or U616 (N_616,N_425,N_595);
and U617 (N_617,N_330,N_561);
and U618 (N_618,In_306,N_162);
nor U619 (N_619,N_406,N_580);
and U620 (N_620,N_592,N_517);
and U621 (N_621,N_550,N_520);
or U622 (N_622,N_559,N_408);
and U623 (N_623,N_500,N_403);
nand U624 (N_624,N_574,In_558);
nand U625 (N_625,N_351,N_506);
or U626 (N_626,N_427,N_67);
or U627 (N_627,N_509,N_591);
and U628 (N_628,N_522,N_341);
xnor U629 (N_629,N_462,N_576);
or U630 (N_630,In_356,N_460);
nand U631 (N_631,N_411,N_555);
nand U632 (N_632,N_519,N_558);
or U633 (N_633,N_545,N_556);
and U634 (N_634,N_543,N_414);
and U635 (N_635,N_469,N_586);
nor U636 (N_636,N_438,N_553);
and U637 (N_637,N_255,N_532);
nand U638 (N_638,N_529,N_409);
or U639 (N_639,N_518,N_569);
nand U640 (N_640,N_570,N_549);
and U641 (N_641,N_531,N_572);
nor U642 (N_642,N_593,N_534);
or U643 (N_643,N_542,N_521);
nand U644 (N_644,N_516,N_508);
nor U645 (N_645,N_584,N_587);
nand U646 (N_646,N_485,N_552);
xnor U647 (N_647,N_515,N_502);
nor U648 (N_648,In_290,N_546);
and U649 (N_649,N_599,N_512);
nand U650 (N_650,N_102,N_578);
or U651 (N_651,N_581,N_471);
nand U652 (N_652,N_535,N_232);
nand U653 (N_653,N_63,N_524);
nand U654 (N_654,N_596,N_594);
and U655 (N_655,N_503,N_577);
and U656 (N_656,N_564,N_526);
nor U657 (N_657,N_567,N_557);
and U658 (N_658,N_208,N_233);
nor U659 (N_659,N_590,N_568);
or U660 (N_660,N_540,N_413);
or U661 (N_661,N_551,N_110);
nand U662 (N_662,N_458,N_536);
nor U663 (N_663,N_582,N_583);
and U664 (N_664,N_527,N_563);
nand U665 (N_665,N_575,In_632);
or U666 (N_666,N_548,N_501);
and U667 (N_667,N_598,N_525);
or U668 (N_668,N_539,In_270);
or U669 (N_669,N_486,N_541);
nor U670 (N_670,N_597,N_573);
or U671 (N_671,N_533,N_544);
or U672 (N_672,N_494,N_511);
and U673 (N_673,N_565,N_530);
or U674 (N_674,N_562,N_523);
and U675 (N_675,N_555,N_560);
nor U676 (N_676,N_544,N_425);
nor U677 (N_677,N_592,N_518);
nand U678 (N_678,N_409,N_542);
nand U679 (N_679,N_564,N_588);
nor U680 (N_680,N_466,N_500);
nand U681 (N_681,N_462,N_548);
nand U682 (N_682,N_517,In_92);
or U683 (N_683,N_545,N_513);
and U684 (N_684,N_587,N_552);
and U685 (N_685,N_589,N_543);
and U686 (N_686,N_462,N_460);
xor U687 (N_687,N_506,N_550);
or U688 (N_688,N_589,N_533);
or U689 (N_689,N_110,N_553);
and U690 (N_690,N_526,N_403);
nand U691 (N_691,In_356,N_597);
and U692 (N_692,N_595,N_582);
or U693 (N_693,N_547,In_270);
or U694 (N_694,N_587,In_306);
and U695 (N_695,N_577,N_506);
nor U696 (N_696,N_563,N_553);
and U697 (N_697,N_67,N_535);
nor U698 (N_698,N_293,N_528);
and U699 (N_699,N_593,N_539);
nor U700 (N_700,N_600,N_684);
nor U701 (N_701,N_643,N_664);
nor U702 (N_702,N_605,N_602);
nor U703 (N_703,N_680,N_645);
nand U704 (N_704,N_633,N_668);
and U705 (N_705,N_607,N_649);
and U706 (N_706,N_630,N_626);
nand U707 (N_707,N_636,N_603);
or U708 (N_708,N_621,N_646);
nand U709 (N_709,N_609,N_669);
nand U710 (N_710,N_687,N_658);
xnor U711 (N_711,N_642,N_653);
and U712 (N_712,N_625,N_688);
and U713 (N_713,N_637,N_611);
and U714 (N_714,N_631,N_627);
nand U715 (N_715,N_675,N_650);
nand U716 (N_716,N_629,N_686);
or U717 (N_717,N_651,N_635);
nand U718 (N_718,N_695,N_612);
nor U719 (N_719,N_659,N_652);
and U720 (N_720,N_656,N_689);
nor U721 (N_721,N_615,N_674);
nand U722 (N_722,N_685,N_690);
and U723 (N_723,N_681,N_644);
and U724 (N_724,N_673,N_610);
and U725 (N_725,N_655,N_618);
or U726 (N_726,N_624,N_677);
or U727 (N_727,N_614,N_657);
or U728 (N_728,N_683,N_623);
nand U729 (N_729,N_619,N_692);
nand U730 (N_730,N_666,N_661);
nand U731 (N_731,N_678,N_620);
nor U732 (N_732,N_699,N_604);
or U733 (N_733,N_662,N_616);
and U734 (N_734,N_667,N_693);
and U735 (N_735,N_608,N_660);
nor U736 (N_736,N_632,N_676);
nand U737 (N_737,N_671,N_606);
nand U738 (N_738,N_639,N_663);
and U739 (N_739,N_697,N_696);
nor U740 (N_740,N_641,N_654);
nand U741 (N_741,N_691,N_665);
xor U742 (N_742,N_634,N_679);
nand U743 (N_743,N_647,N_638);
and U744 (N_744,N_682,N_648);
or U745 (N_745,N_622,N_601);
nand U746 (N_746,N_613,N_640);
nand U747 (N_747,N_617,N_698);
or U748 (N_748,N_672,N_694);
nand U749 (N_749,N_628,N_670);
nand U750 (N_750,N_606,N_693);
and U751 (N_751,N_669,N_619);
nor U752 (N_752,N_663,N_621);
nor U753 (N_753,N_656,N_676);
nor U754 (N_754,N_613,N_673);
nor U755 (N_755,N_669,N_689);
and U756 (N_756,N_682,N_621);
nand U757 (N_757,N_634,N_642);
or U758 (N_758,N_618,N_634);
or U759 (N_759,N_619,N_633);
or U760 (N_760,N_688,N_646);
and U761 (N_761,N_657,N_620);
nand U762 (N_762,N_699,N_679);
xnor U763 (N_763,N_622,N_684);
or U764 (N_764,N_653,N_629);
nand U765 (N_765,N_676,N_607);
nor U766 (N_766,N_625,N_607);
and U767 (N_767,N_696,N_627);
or U768 (N_768,N_697,N_621);
and U769 (N_769,N_657,N_608);
nand U770 (N_770,N_637,N_651);
or U771 (N_771,N_657,N_656);
or U772 (N_772,N_653,N_665);
nand U773 (N_773,N_602,N_622);
nor U774 (N_774,N_619,N_650);
nor U775 (N_775,N_631,N_639);
or U776 (N_776,N_603,N_660);
and U777 (N_777,N_652,N_624);
nor U778 (N_778,N_612,N_606);
nor U779 (N_779,N_604,N_680);
or U780 (N_780,N_624,N_632);
nor U781 (N_781,N_689,N_617);
nand U782 (N_782,N_646,N_685);
or U783 (N_783,N_650,N_646);
nand U784 (N_784,N_647,N_639);
nand U785 (N_785,N_600,N_680);
or U786 (N_786,N_671,N_634);
or U787 (N_787,N_658,N_685);
nor U788 (N_788,N_622,N_664);
xor U789 (N_789,N_690,N_616);
nand U790 (N_790,N_664,N_616);
and U791 (N_791,N_672,N_654);
or U792 (N_792,N_650,N_651);
or U793 (N_793,N_676,N_622);
or U794 (N_794,N_642,N_602);
or U795 (N_795,N_688,N_662);
or U796 (N_796,N_641,N_689);
nor U797 (N_797,N_600,N_646);
nor U798 (N_798,N_680,N_696);
nor U799 (N_799,N_635,N_681);
nor U800 (N_800,N_717,N_738);
nor U801 (N_801,N_794,N_749);
or U802 (N_802,N_701,N_784);
and U803 (N_803,N_767,N_783);
or U804 (N_804,N_785,N_751);
nand U805 (N_805,N_728,N_753);
and U806 (N_806,N_731,N_702);
and U807 (N_807,N_711,N_745);
nor U808 (N_808,N_713,N_718);
nand U809 (N_809,N_725,N_780);
or U810 (N_810,N_732,N_758);
nor U811 (N_811,N_776,N_733);
or U812 (N_812,N_747,N_781);
nand U813 (N_813,N_740,N_787);
xnor U814 (N_814,N_797,N_766);
and U815 (N_815,N_791,N_704);
nand U816 (N_816,N_750,N_789);
xnor U817 (N_817,N_708,N_700);
nand U818 (N_818,N_778,N_719);
nor U819 (N_819,N_737,N_754);
or U820 (N_820,N_710,N_774);
nor U821 (N_821,N_771,N_741);
or U822 (N_822,N_786,N_743);
nor U823 (N_823,N_796,N_721);
or U824 (N_824,N_792,N_775);
and U825 (N_825,N_770,N_757);
nor U826 (N_826,N_788,N_798);
nor U827 (N_827,N_735,N_795);
and U828 (N_828,N_729,N_764);
nor U829 (N_829,N_761,N_782);
or U830 (N_830,N_793,N_712);
nand U831 (N_831,N_716,N_705);
and U832 (N_832,N_755,N_707);
or U833 (N_833,N_714,N_760);
nor U834 (N_834,N_706,N_742);
nor U835 (N_835,N_736,N_790);
and U836 (N_836,N_703,N_772);
and U837 (N_837,N_720,N_773);
or U838 (N_838,N_765,N_779);
and U839 (N_839,N_734,N_722);
nor U840 (N_840,N_799,N_759);
xnor U841 (N_841,N_726,N_768);
and U842 (N_842,N_777,N_739);
or U843 (N_843,N_730,N_769);
or U844 (N_844,N_723,N_715);
nand U845 (N_845,N_763,N_752);
nor U846 (N_846,N_746,N_709);
and U847 (N_847,N_762,N_724);
or U848 (N_848,N_748,N_727);
nand U849 (N_849,N_744,N_756);
xnor U850 (N_850,N_762,N_737);
nor U851 (N_851,N_796,N_748);
nor U852 (N_852,N_710,N_726);
and U853 (N_853,N_716,N_711);
nand U854 (N_854,N_795,N_737);
or U855 (N_855,N_702,N_784);
nor U856 (N_856,N_778,N_755);
nor U857 (N_857,N_779,N_707);
nor U858 (N_858,N_781,N_767);
and U859 (N_859,N_793,N_766);
nand U860 (N_860,N_766,N_707);
or U861 (N_861,N_789,N_727);
and U862 (N_862,N_746,N_787);
nand U863 (N_863,N_733,N_782);
and U864 (N_864,N_762,N_728);
nand U865 (N_865,N_783,N_743);
and U866 (N_866,N_784,N_730);
nor U867 (N_867,N_787,N_725);
nand U868 (N_868,N_759,N_760);
nor U869 (N_869,N_741,N_738);
or U870 (N_870,N_770,N_706);
or U871 (N_871,N_737,N_790);
and U872 (N_872,N_795,N_791);
nand U873 (N_873,N_723,N_710);
and U874 (N_874,N_741,N_798);
nand U875 (N_875,N_774,N_739);
and U876 (N_876,N_740,N_728);
and U877 (N_877,N_716,N_781);
or U878 (N_878,N_721,N_755);
or U879 (N_879,N_734,N_771);
or U880 (N_880,N_706,N_757);
nand U881 (N_881,N_740,N_796);
or U882 (N_882,N_712,N_705);
nand U883 (N_883,N_791,N_708);
xnor U884 (N_884,N_734,N_743);
xor U885 (N_885,N_749,N_751);
and U886 (N_886,N_722,N_711);
nor U887 (N_887,N_772,N_769);
or U888 (N_888,N_744,N_701);
and U889 (N_889,N_740,N_749);
nor U890 (N_890,N_720,N_747);
and U891 (N_891,N_767,N_730);
or U892 (N_892,N_785,N_736);
nor U893 (N_893,N_788,N_776);
nor U894 (N_894,N_700,N_753);
nand U895 (N_895,N_776,N_714);
or U896 (N_896,N_726,N_715);
and U897 (N_897,N_763,N_795);
nor U898 (N_898,N_702,N_778);
nand U899 (N_899,N_780,N_756);
and U900 (N_900,N_880,N_817);
and U901 (N_901,N_870,N_856);
nand U902 (N_902,N_846,N_815);
or U903 (N_903,N_875,N_858);
or U904 (N_904,N_816,N_804);
and U905 (N_905,N_831,N_887);
and U906 (N_906,N_863,N_840);
nor U907 (N_907,N_847,N_800);
nor U908 (N_908,N_869,N_805);
or U909 (N_909,N_835,N_890);
or U910 (N_910,N_892,N_855);
and U911 (N_911,N_864,N_891);
xor U912 (N_912,N_829,N_857);
xnor U913 (N_913,N_823,N_814);
or U914 (N_914,N_834,N_867);
nor U915 (N_915,N_841,N_873);
or U916 (N_916,N_894,N_828);
and U917 (N_917,N_885,N_813);
nand U918 (N_918,N_899,N_861);
nor U919 (N_919,N_803,N_812);
or U920 (N_920,N_844,N_839);
nor U921 (N_921,N_801,N_884);
nand U922 (N_922,N_898,N_811);
nor U923 (N_923,N_827,N_862);
nand U924 (N_924,N_874,N_802);
or U925 (N_925,N_836,N_833);
or U926 (N_926,N_809,N_886);
and U927 (N_927,N_830,N_878);
xnor U928 (N_928,N_848,N_888);
nor U929 (N_929,N_806,N_842);
nand U930 (N_930,N_881,N_879);
and U931 (N_931,N_849,N_821);
nand U932 (N_932,N_859,N_818);
nand U933 (N_933,N_819,N_824);
nand U934 (N_934,N_889,N_810);
nor U935 (N_935,N_860,N_838);
nand U936 (N_936,N_871,N_882);
nand U937 (N_937,N_876,N_825);
or U938 (N_938,N_851,N_808);
or U939 (N_939,N_837,N_895);
nor U940 (N_940,N_893,N_845);
nor U941 (N_941,N_897,N_854);
nand U942 (N_942,N_868,N_832);
and U943 (N_943,N_826,N_820);
and U944 (N_944,N_883,N_866);
and U945 (N_945,N_843,N_865);
or U946 (N_946,N_877,N_807);
nand U947 (N_947,N_852,N_896);
nand U948 (N_948,N_850,N_822);
nor U949 (N_949,N_853,N_872);
nor U950 (N_950,N_849,N_869);
nand U951 (N_951,N_878,N_832);
nand U952 (N_952,N_811,N_845);
nand U953 (N_953,N_804,N_822);
nand U954 (N_954,N_807,N_851);
and U955 (N_955,N_892,N_848);
or U956 (N_956,N_811,N_831);
or U957 (N_957,N_846,N_887);
or U958 (N_958,N_862,N_810);
nand U959 (N_959,N_810,N_882);
nor U960 (N_960,N_898,N_872);
nand U961 (N_961,N_830,N_834);
and U962 (N_962,N_886,N_856);
xor U963 (N_963,N_820,N_877);
and U964 (N_964,N_828,N_811);
and U965 (N_965,N_860,N_862);
or U966 (N_966,N_848,N_879);
nor U967 (N_967,N_867,N_813);
nor U968 (N_968,N_843,N_834);
nor U969 (N_969,N_814,N_879);
nand U970 (N_970,N_847,N_821);
or U971 (N_971,N_888,N_865);
or U972 (N_972,N_860,N_808);
nand U973 (N_973,N_889,N_805);
nor U974 (N_974,N_818,N_863);
or U975 (N_975,N_835,N_858);
or U976 (N_976,N_871,N_874);
or U977 (N_977,N_808,N_889);
xor U978 (N_978,N_836,N_829);
nor U979 (N_979,N_810,N_815);
nor U980 (N_980,N_880,N_892);
and U981 (N_981,N_890,N_894);
nor U982 (N_982,N_896,N_858);
nor U983 (N_983,N_896,N_890);
or U984 (N_984,N_855,N_899);
nor U985 (N_985,N_822,N_861);
or U986 (N_986,N_842,N_844);
or U987 (N_987,N_862,N_896);
or U988 (N_988,N_848,N_891);
nand U989 (N_989,N_838,N_867);
nand U990 (N_990,N_810,N_887);
xor U991 (N_991,N_836,N_817);
nand U992 (N_992,N_867,N_839);
or U993 (N_993,N_887,N_886);
nor U994 (N_994,N_882,N_853);
nor U995 (N_995,N_885,N_867);
nand U996 (N_996,N_860,N_834);
or U997 (N_997,N_811,N_863);
nand U998 (N_998,N_815,N_889);
nor U999 (N_999,N_801,N_855);
nand U1000 (N_1000,N_904,N_971);
nor U1001 (N_1001,N_911,N_956);
xnor U1002 (N_1002,N_905,N_984);
and U1003 (N_1003,N_998,N_977);
or U1004 (N_1004,N_951,N_985);
and U1005 (N_1005,N_903,N_982);
and U1006 (N_1006,N_953,N_991);
or U1007 (N_1007,N_983,N_946);
or U1008 (N_1008,N_947,N_974);
or U1009 (N_1009,N_918,N_959);
nand U1010 (N_1010,N_919,N_950);
nor U1011 (N_1011,N_928,N_997);
nand U1012 (N_1012,N_975,N_938);
nand U1013 (N_1013,N_987,N_962);
and U1014 (N_1014,N_966,N_912);
and U1015 (N_1015,N_941,N_995);
nand U1016 (N_1016,N_964,N_976);
nand U1017 (N_1017,N_907,N_996);
xor U1018 (N_1018,N_934,N_948);
and U1019 (N_1019,N_972,N_980);
or U1020 (N_1020,N_942,N_937);
or U1021 (N_1021,N_901,N_986);
nand U1022 (N_1022,N_917,N_940);
and U1023 (N_1023,N_958,N_920);
and U1024 (N_1024,N_936,N_978);
xor U1025 (N_1025,N_955,N_990);
and U1026 (N_1026,N_925,N_922);
nand U1027 (N_1027,N_988,N_967);
nor U1028 (N_1028,N_932,N_923);
nand U1029 (N_1029,N_909,N_944);
nor U1030 (N_1030,N_930,N_949);
nand U1031 (N_1031,N_915,N_954);
xnor U1032 (N_1032,N_969,N_926);
nor U1033 (N_1033,N_989,N_900);
nand U1034 (N_1034,N_957,N_963);
and U1035 (N_1035,N_968,N_994);
nand U1036 (N_1036,N_970,N_965);
nor U1037 (N_1037,N_906,N_992);
nor U1038 (N_1038,N_945,N_916);
and U1039 (N_1039,N_931,N_914);
or U1040 (N_1040,N_973,N_943);
and U1041 (N_1041,N_921,N_952);
or U1042 (N_1042,N_902,N_927);
or U1043 (N_1043,N_979,N_908);
and U1044 (N_1044,N_933,N_960);
nor U1045 (N_1045,N_999,N_913);
nor U1046 (N_1046,N_910,N_929);
nor U1047 (N_1047,N_993,N_961);
or U1048 (N_1048,N_981,N_935);
or U1049 (N_1049,N_924,N_939);
nor U1050 (N_1050,N_960,N_996);
nor U1051 (N_1051,N_953,N_918);
and U1052 (N_1052,N_938,N_921);
and U1053 (N_1053,N_981,N_972);
or U1054 (N_1054,N_967,N_921);
nor U1055 (N_1055,N_967,N_971);
nand U1056 (N_1056,N_938,N_982);
or U1057 (N_1057,N_919,N_989);
nand U1058 (N_1058,N_937,N_944);
or U1059 (N_1059,N_940,N_906);
nor U1060 (N_1060,N_967,N_944);
nor U1061 (N_1061,N_953,N_933);
or U1062 (N_1062,N_915,N_930);
or U1063 (N_1063,N_926,N_955);
nand U1064 (N_1064,N_924,N_966);
nor U1065 (N_1065,N_958,N_918);
or U1066 (N_1066,N_936,N_984);
and U1067 (N_1067,N_950,N_959);
nand U1068 (N_1068,N_929,N_966);
or U1069 (N_1069,N_917,N_994);
nand U1070 (N_1070,N_926,N_902);
or U1071 (N_1071,N_933,N_952);
nor U1072 (N_1072,N_905,N_901);
nand U1073 (N_1073,N_997,N_945);
and U1074 (N_1074,N_939,N_943);
nand U1075 (N_1075,N_980,N_963);
and U1076 (N_1076,N_967,N_915);
and U1077 (N_1077,N_935,N_988);
nor U1078 (N_1078,N_968,N_961);
or U1079 (N_1079,N_910,N_934);
or U1080 (N_1080,N_903,N_957);
xnor U1081 (N_1081,N_906,N_997);
nor U1082 (N_1082,N_908,N_996);
nand U1083 (N_1083,N_982,N_953);
nor U1084 (N_1084,N_944,N_981);
nor U1085 (N_1085,N_982,N_951);
nand U1086 (N_1086,N_967,N_924);
nor U1087 (N_1087,N_915,N_968);
nor U1088 (N_1088,N_951,N_911);
or U1089 (N_1089,N_920,N_986);
nand U1090 (N_1090,N_966,N_982);
xor U1091 (N_1091,N_967,N_934);
nand U1092 (N_1092,N_904,N_998);
nand U1093 (N_1093,N_911,N_996);
or U1094 (N_1094,N_924,N_983);
nand U1095 (N_1095,N_986,N_991);
or U1096 (N_1096,N_966,N_942);
or U1097 (N_1097,N_933,N_944);
xor U1098 (N_1098,N_901,N_994);
and U1099 (N_1099,N_932,N_918);
nand U1100 (N_1100,N_1020,N_1023);
or U1101 (N_1101,N_1084,N_1041);
nor U1102 (N_1102,N_1057,N_1096);
or U1103 (N_1103,N_1016,N_1055);
or U1104 (N_1104,N_1074,N_1073);
nand U1105 (N_1105,N_1099,N_1043);
or U1106 (N_1106,N_1097,N_1076);
nor U1107 (N_1107,N_1086,N_1051);
and U1108 (N_1108,N_1068,N_1054);
and U1109 (N_1109,N_1026,N_1080);
nand U1110 (N_1110,N_1036,N_1038);
xnor U1111 (N_1111,N_1030,N_1040);
nand U1112 (N_1112,N_1077,N_1079);
nor U1113 (N_1113,N_1039,N_1063);
nor U1114 (N_1114,N_1029,N_1082);
nand U1115 (N_1115,N_1003,N_1048);
and U1116 (N_1116,N_1059,N_1083);
nor U1117 (N_1117,N_1058,N_1049);
nor U1118 (N_1118,N_1044,N_1098);
or U1119 (N_1119,N_1065,N_1067);
or U1120 (N_1120,N_1093,N_1006);
or U1121 (N_1121,N_1085,N_1027);
or U1122 (N_1122,N_1010,N_1031);
and U1123 (N_1123,N_1094,N_1066);
or U1124 (N_1124,N_1009,N_1034);
and U1125 (N_1125,N_1037,N_1081);
nor U1126 (N_1126,N_1091,N_1005);
and U1127 (N_1127,N_1033,N_1008);
nand U1128 (N_1128,N_1011,N_1002);
nand U1129 (N_1129,N_1013,N_1000);
nand U1130 (N_1130,N_1001,N_1050);
or U1131 (N_1131,N_1025,N_1035);
nor U1132 (N_1132,N_1052,N_1014);
nor U1133 (N_1133,N_1028,N_1012);
or U1134 (N_1134,N_1070,N_1022);
and U1135 (N_1135,N_1007,N_1092);
and U1136 (N_1136,N_1072,N_1018);
and U1137 (N_1137,N_1075,N_1042);
nand U1138 (N_1138,N_1004,N_1032);
and U1139 (N_1139,N_1019,N_1062);
nand U1140 (N_1140,N_1015,N_1069);
or U1141 (N_1141,N_1053,N_1095);
nand U1142 (N_1142,N_1060,N_1047);
nand U1143 (N_1143,N_1090,N_1088);
and U1144 (N_1144,N_1021,N_1061);
or U1145 (N_1145,N_1017,N_1064);
and U1146 (N_1146,N_1087,N_1078);
and U1147 (N_1147,N_1071,N_1046);
nand U1148 (N_1148,N_1056,N_1045);
or U1149 (N_1149,N_1089,N_1024);
and U1150 (N_1150,N_1028,N_1033);
nand U1151 (N_1151,N_1092,N_1021);
and U1152 (N_1152,N_1000,N_1096);
nor U1153 (N_1153,N_1088,N_1065);
or U1154 (N_1154,N_1075,N_1065);
and U1155 (N_1155,N_1065,N_1042);
or U1156 (N_1156,N_1006,N_1025);
nand U1157 (N_1157,N_1061,N_1083);
nor U1158 (N_1158,N_1044,N_1011);
and U1159 (N_1159,N_1008,N_1010);
or U1160 (N_1160,N_1096,N_1066);
and U1161 (N_1161,N_1034,N_1017);
or U1162 (N_1162,N_1002,N_1012);
nand U1163 (N_1163,N_1025,N_1092);
or U1164 (N_1164,N_1038,N_1032);
nor U1165 (N_1165,N_1001,N_1067);
or U1166 (N_1166,N_1097,N_1053);
nor U1167 (N_1167,N_1045,N_1014);
nor U1168 (N_1168,N_1025,N_1001);
and U1169 (N_1169,N_1060,N_1075);
and U1170 (N_1170,N_1023,N_1064);
nor U1171 (N_1171,N_1062,N_1084);
nand U1172 (N_1172,N_1095,N_1081);
and U1173 (N_1173,N_1018,N_1083);
nand U1174 (N_1174,N_1034,N_1069);
nand U1175 (N_1175,N_1005,N_1011);
nand U1176 (N_1176,N_1016,N_1096);
nor U1177 (N_1177,N_1079,N_1084);
nand U1178 (N_1178,N_1078,N_1025);
and U1179 (N_1179,N_1050,N_1092);
and U1180 (N_1180,N_1034,N_1060);
or U1181 (N_1181,N_1021,N_1086);
and U1182 (N_1182,N_1038,N_1053);
or U1183 (N_1183,N_1029,N_1024);
nand U1184 (N_1184,N_1027,N_1039);
and U1185 (N_1185,N_1073,N_1012);
nand U1186 (N_1186,N_1067,N_1005);
nand U1187 (N_1187,N_1072,N_1041);
nor U1188 (N_1188,N_1039,N_1037);
and U1189 (N_1189,N_1094,N_1020);
nand U1190 (N_1190,N_1049,N_1004);
nand U1191 (N_1191,N_1002,N_1033);
nand U1192 (N_1192,N_1097,N_1090);
nor U1193 (N_1193,N_1008,N_1044);
or U1194 (N_1194,N_1036,N_1078);
or U1195 (N_1195,N_1012,N_1091);
nand U1196 (N_1196,N_1040,N_1054);
nand U1197 (N_1197,N_1069,N_1033);
or U1198 (N_1198,N_1092,N_1068);
nor U1199 (N_1199,N_1072,N_1057);
nand U1200 (N_1200,N_1154,N_1121);
or U1201 (N_1201,N_1131,N_1134);
nor U1202 (N_1202,N_1187,N_1105);
xor U1203 (N_1203,N_1186,N_1137);
or U1204 (N_1204,N_1133,N_1144);
nand U1205 (N_1205,N_1123,N_1164);
and U1206 (N_1206,N_1115,N_1104);
xor U1207 (N_1207,N_1153,N_1119);
nand U1208 (N_1208,N_1168,N_1191);
nor U1209 (N_1209,N_1155,N_1157);
nand U1210 (N_1210,N_1100,N_1116);
nand U1211 (N_1211,N_1101,N_1114);
nor U1212 (N_1212,N_1128,N_1174);
nor U1213 (N_1213,N_1142,N_1199);
nand U1214 (N_1214,N_1169,N_1183);
or U1215 (N_1215,N_1149,N_1161);
nand U1216 (N_1216,N_1130,N_1127);
nor U1217 (N_1217,N_1112,N_1192);
nand U1218 (N_1218,N_1176,N_1136);
nor U1219 (N_1219,N_1189,N_1143);
or U1220 (N_1220,N_1170,N_1138);
or U1221 (N_1221,N_1167,N_1177);
nand U1222 (N_1222,N_1194,N_1120);
or U1223 (N_1223,N_1106,N_1113);
nor U1224 (N_1224,N_1159,N_1160);
nor U1225 (N_1225,N_1141,N_1162);
and U1226 (N_1226,N_1173,N_1126);
and U1227 (N_1227,N_1178,N_1111);
or U1228 (N_1228,N_1193,N_1195);
nor U1229 (N_1229,N_1125,N_1184);
and U1230 (N_1230,N_1109,N_1196);
xnor U1231 (N_1231,N_1145,N_1107);
and U1232 (N_1232,N_1158,N_1182);
or U1233 (N_1233,N_1163,N_1139);
nor U1234 (N_1234,N_1147,N_1140);
or U1235 (N_1235,N_1124,N_1165);
and U1236 (N_1236,N_1197,N_1148);
or U1237 (N_1237,N_1118,N_1172);
or U1238 (N_1238,N_1108,N_1175);
nor U1239 (N_1239,N_1166,N_1103);
and U1240 (N_1240,N_1122,N_1117);
nor U1241 (N_1241,N_1198,N_1171);
or U1242 (N_1242,N_1151,N_1146);
nor U1243 (N_1243,N_1180,N_1135);
and U1244 (N_1244,N_1181,N_1156);
nand U1245 (N_1245,N_1179,N_1185);
or U1246 (N_1246,N_1132,N_1150);
nor U1247 (N_1247,N_1152,N_1190);
nor U1248 (N_1248,N_1102,N_1129);
nor U1249 (N_1249,N_1110,N_1188);
nand U1250 (N_1250,N_1135,N_1197);
and U1251 (N_1251,N_1199,N_1158);
nand U1252 (N_1252,N_1100,N_1155);
or U1253 (N_1253,N_1179,N_1124);
and U1254 (N_1254,N_1163,N_1119);
and U1255 (N_1255,N_1142,N_1151);
nand U1256 (N_1256,N_1103,N_1132);
or U1257 (N_1257,N_1139,N_1198);
or U1258 (N_1258,N_1190,N_1199);
nand U1259 (N_1259,N_1163,N_1186);
nor U1260 (N_1260,N_1178,N_1198);
or U1261 (N_1261,N_1145,N_1195);
and U1262 (N_1262,N_1195,N_1125);
nand U1263 (N_1263,N_1133,N_1177);
xor U1264 (N_1264,N_1111,N_1184);
nand U1265 (N_1265,N_1141,N_1128);
nand U1266 (N_1266,N_1103,N_1154);
and U1267 (N_1267,N_1130,N_1112);
nor U1268 (N_1268,N_1136,N_1137);
nor U1269 (N_1269,N_1178,N_1174);
or U1270 (N_1270,N_1141,N_1198);
and U1271 (N_1271,N_1171,N_1191);
nand U1272 (N_1272,N_1134,N_1132);
nand U1273 (N_1273,N_1142,N_1116);
nor U1274 (N_1274,N_1151,N_1175);
nor U1275 (N_1275,N_1135,N_1111);
and U1276 (N_1276,N_1106,N_1112);
nor U1277 (N_1277,N_1114,N_1122);
and U1278 (N_1278,N_1161,N_1111);
nand U1279 (N_1279,N_1138,N_1149);
and U1280 (N_1280,N_1155,N_1163);
nand U1281 (N_1281,N_1162,N_1197);
nor U1282 (N_1282,N_1114,N_1139);
and U1283 (N_1283,N_1159,N_1161);
nor U1284 (N_1284,N_1158,N_1167);
or U1285 (N_1285,N_1137,N_1131);
or U1286 (N_1286,N_1143,N_1173);
and U1287 (N_1287,N_1199,N_1162);
nor U1288 (N_1288,N_1163,N_1150);
and U1289 (N_1289,N_1165,N_1184);
or U1290 (N_1290,N_1153,N_1167);
and U1291 (N_1291,N_1112,N_1121);
nand U1292 (N_1292,N_1180,N_1188);
or U1293 (N_1293,N_1186,N_1129);
nand U1294 (N_1294,N_1132,N_1149);
nor U1295 (N_1295,N_1168,N_1120);
and U1296 (N_1296,N_1169,N_1189);
nor U1297 (N_1297,N_1183,N_1196);
nor U1298 (N_1298,N_1157,N_1179);
nand U1299 (N_1299,N_1131,N_1113);
or U1300 (N_1300,N_1212,N_1293);
nor U1301 (N_1301,N_1280,N_1285);
and U1302 (N_1302,N_1282,N_1242);
nor U1303 (N_1303,N_1259,N_1240);
nand U1304 (N_1304,N_1279,N_1232);
or U1305 (N_1305,N_1203,N_1222);
or U1306 (N_1306,N_1251,N_1233);
and U1307 (N_1307,N_1260,N_1208);
or U1308 (N_1308,N_1207,N_1268);
nand U1309 (N_1309,N_1278,N_1249);
or U1310 (N_1310,N_1254,N_1218);
or U1311 (N_1311,N_1291,N_1277);
or U1312 (N_1312,N_1294,N_1246);
nor U1313 (N_1313,N_1248,N_1299);
and U1314 (N_1314,N_1243,N_1200);
or U1315 (N_1315,N_1226,N_1221);
nor U1316 (N_1316,N_1234,N_1284);
or U1317 (N_1317,N_1247,N_1269);
nand U1318 (N_1318,N_1295,N_1271);
nand U1319 (N_1319,N_1244,N_1252);
nand U1320 (N_1320,N_1227,N_1217);
nand U1321 (N_1321,N_1250,N_1224);
nand U1322 (N_1322,N_1290,N_1264);
nand U1323 (N_1323,N_1253,N_1241);
nor U1324 (N_1324,N_1286,N_1215);
nand U1325 (N_1325,N_1229,N_1230);
nand U1326 (N_1326,N_1298,N_1255);
or U1327 (N_1327,N_1273,N_1283);
or U1328 (N_1328,N_1267,N_1238);
and U1329 (N_1329,N_1214,N_1275);
or U1330 (N_1330,N_1201,N_1239);
nor U1331 (N_1331,N_1206,N_1292);
nand U1332 (N_1332,N_1272,N_1261);
nand U1333 (N_1333,N_1205,N_1263);
nand U1334 (N_1334,N_1274,N_1209);
nor U1335 (N_1335,N_1256,N_1296);
or U1336 (N_1336,N_1216,N_1262);
nand U1337 (N_1337,N_1236,N_1287);
or U1338 (N_1338,N_1231,N_1220);
nand U1339 (N_1339,N_1258,N_1210);
or U1340 (N_1340,N_1281,N_1219);
and U1341 (N_1341,N_1213,N_1276);
nand U1342 (N_1342,N_1289,N_1211);
and U1343 (N_1343,N_1257,N_1223);
and U1344 (N_1344,N_1225,N_1245);
nor U1345 (N_1345,N_1202,N_1266);
and U1346 (N_1346,N_1204,N_1228);
and U1347 (N_1347,N_1265,N_1297);
nand U1348 (N_1348,N_1288,N_1270);
or U1349 (N_1349,N_1237,N_1235);
nor U1350 (N_1350,N_1271,N_1218);
nor U1351 (N_1351,N_1267,N_1201);
and U1352 (N_1352,N_1256,N_1248);
or U1353 (N_1353,N_1200,N_1211);
and U1354 (N_1354,N_1281,N_1201);
nor U1355 (N_1355,N_1288,N_1297);
and U1356 (N_1356,N_1221,N_1246);
or U1357 (N_1357,N_1253,N_1270);
or U1358 (N_1358,N_1207,N_1215);
nor U1359 (N_1359,N_1286,N_1238);
and U1360 (N_1360,N_1206,N_1201);
and U1361 (N_1361,N_1221,N_1200);
or U1362 (N_1362,N_1223,N_1242);
or U1363 (N_1363,N_1291,N_1299);
or U1364 (N_1364,N_1227,N_1234);
or U1365 (N_1365,N_1295,N_1268);
and U1366 (N_1366,N_1234,N_1277);
nor U1367 (N_1367,N_1215,N_1256);
or U1368 (N_1368,N_1248,N_1271);
nor U1369 (N_1369,N_1202,N_1201);
nand U1370 (N_1370,N_1288,N_1223);
or U1371 (N_1371,N_1265,N_1226);
xor U1372 (N_1372,N_1251,N_1249);
nor U1373 (N_1373,N_1273,N_1284);
or U1374 (N_1374,N_1214,N_1286);
nand U1375 (N_1375,N_1266,N_1217);
nor U1376 (N_1376,N_1289,N_1255);
or U1377 (N_1377,N_1251,N_1298);
xnor U1378 (N_1378,N_1252,N_1283);
nand U1379 (N_1379,N_1252,N_1200);
or U1380 (N_1380,N_1200,N_1245);
or U1381 (N_1381,N_1264,N_1286);
xor U1382 (N_1382,N_1210,N_1234);
or U1383 (N_1383,N_1228,N_1262);
nor U1384 (N_1384,N_1240,N_1288);
and U1385 (N_1385,N_1241,N_1209);
and U1386 (N_1386,N_1287,N_1226);
and U1387 (N_1387,N_1274,N_1256);
nand U1388 (N_1388,N_1249,N_1288);
and U1389 (N_1389,N_1267,N_1271);
and U1390 (N_1390,N_1203,N_1256);
and U1391 (N_1391,N_1248,N_1201);
and U1392 (N_1392,N_1206,N_1277);
and U1393 (N_1393,N_1263,N_1212);
nor U1394 (N_1394,N_1250,N_1202);
or U1395 (N_1395,N_1294,N_1223);
xor U1396 (N_1396,N_1287,N_1246);
nand U1397 (N_1397,N_1274,N_1223);
and U1398 (N_1398,N_1223,N_1218);
and U1399 (N_1399,N_1279,N_1298);
nor U1400 (N_1400,N_1355,N_1317);
nand U1401 (N_1401,N_1377,N_1375);
and U1402 (N_1402,N_1387,N_1337);
nor U1403 (N_1403,N_1346,N_1368);
nor U1404 (N_1404,N_1394,N_1338);
nand U1405 (N_1405,N_1342,N_1303);
nor U1406 (N_1406,N_1331,N_1334);
nand U1407 (N_1407,N_1341,N_1376);
xnor U1408 (N_1408,N_1339,N_1391);
or U1409 (N_1409,N_1371,N_1388);
nand U1410 (N_1410,N_1301,N_1305);
nand U1411 (N_1411,N_1300,N_1392);
or U1412 (N_1412,N_1309,N_1313);
or U1413 (N_1413,N_1359,N_1365);
or U1414 (N_1414,N_1328,N_1353);
or U1415 (N_1415,N_1350,N_1327);
nor U1416 (N_1416,N_1310,N_1347);
and U1417 (N_1417,N_1393,N_1367);
nand U1418 (N_1418,N_1399,N_1369);
nor U1419 (N_1419,N_1326,N_1374);
or U1420 (N_1420,N_1370,N_1381);
nand U1421 (N_1421,N_1372,N_1319);
nor U1422 (N_1422,N_1366,N_1318);
nor U1423 (N_1423,N_1361,N_1325);
and U1424 (N_1424,N_1311,N_1329);
or U1425 (N_1425,N_1356,N_1373);
nor U1426 (N_1426,N_1322,N_1323);
nor U1427 (N_1427,N_1336,N_1343);
and U1428 (N_1428,N_1321,N_1320);
nor U1429 (N_1429,N_1364,N_1315);
or U1430 (N_1430,N_1324,N_1348);
or U1431 (N_1431,N_1335,N_1316);
nand U1432 (N_1432,N_1386,N_1380);
nor U1433 (N_1433,N_1302,N_1333);
nor U1434 (N_1434,N_1349,N_1352);
nor U1435 (N_1435,N_1344,N_1330);
nand U1436 (N_1436,N_1345,N_1390);
and U1437 (N_1437,N_1360,N_1385);
nand U1438 (N_1438,N_1307,N_1358);
and U1439 (N_1439,N_1308,N_1382);
or U1440 (N_1440,N_1378,N_1354);
nor U1441 (N_1441,N_1351,N_1383);
and U1442 (N_1442,N_1363,N_1396);
or U1443 (N_1443,N_1357,N_1398);
and U1444 (N_1444,N_1384,N_1397);
or U1445 (N_1445,N_1362,N_1332);
and U1446 (N_1446,N_1306,N_1395);
nand U1447 (N_1447,N_1312,N_1314);
nor U1448 (N_1448,N_1340,N_1389);
and U1449 (N_1449,N_1304,N_1379);
nand U1450 (N_1450,N_1367,N_1322);
or U1451 (N_1451,N_1358,N_1342);
nor U1452 (N_1452,N_1329,N_1368);
nor U1453 (N_1453,N_1317,N_1351);
and U1454 (N_1454,N_1353,N_1332);
nand U1455 (N_1455,N_1352,N_1338);
nor U1456 (N_1456,N_1391,N_1356);
or U1457 (N_1457,N_1389,N_1396);
nor U1458 (N_1458,N_1358,N_1393);
or U1459 (N_1459,N_1348,N_1382);
or U1460 (N_1460,N_1351,N_1382);
nor U1461 (N_1461,N_1318,N_1395);
nand U1462 (N_1462,N_1340,N_1353);
nor U1463 (N_1463,N_1315,N_1365);
nand U1464 (N_1464,N_1355,N_1349);
or U1465 (N_1465,N_1372,N_1345);
and U1466 (N_1466,N_1367,N_1377);
nand U1467 (N_1467,N_1317,N_1336);
or U1468 (N_1468,N_1305,N_1376);
or U1469 (N_1469,N_1366,N_1300);
or U1470 (N_1470,N_1374,N_1305);
and U1471 (N_1471,N_1383,N_1307);
or U1472 (N_1472,N_1304,N_1369);
nor U1473 (N_1473,N_1329,N_1312);
nand U1474 (N_1474,N_1376,N_1355);
nand U1475 (N_1475,N_1322,N_1391);
or U1476 (N_1476,N_1339,N_1300);
nor U1477 (N_1477,N_1382,N_1342);
nor U1478 (N_1478,N_1328,N_1380);
or U1479 (N_1479,N_1339,N_1322);
or U1480 (N_1480,N_1378,N_1389);
or U1481 (N_1481,N_1320,N_1330);
and U1482 (N_1482,N_1357,N_1367);
nand U1483 (N_1483,N_1389,N_1316);
nand U1484 (N_1484,N_1346,N_1394);
and U1485 (N_1485,N_1315,N_1321);
nand U1486 (N_1486,N_1349,N_1358);
and U1487 (N_1487,N_1354,N_1329);
and U1488 (N_1488,N_1300,N_1337);
or U1489 (N_1489,N_1323,N_1377);
or U1490 (N_1490,N_1355,N_1370);
and U1491 (N_1491,N_1327,N_1399);
and U1492 (N_1492,N_1387,N_1362);
or U1493 (N_1493,N_1374,N_1310);
nand U1494 (N_1494,N_1325,N_1356);
and U1495 (N_1495,N_1328,N_1330);
and U1496 (N_1496,N_1378,N_1396);
and U1497 (N_1497,N_1333,N_1395);
nor U1498 (N_1498,N_1338,N_1354);
nor U1499 (N_1499,N_1395,N_1315);
nand U1500 (N_1500,N_1482,N_1472);
nor U1501 (N_1501,N_1494,N_1468);
and U1502 (N_1502,N_1401,N_1480);
xor U1503 (N_1503,N_1434,N_1411);
or U1504 (N_1504,N_1441,N_1404);
or U1505 (N_1505,N_1474,N_1431);
nor U1506 (N_1506,N_1495,N_1471);
nor U1507 (N_1507,N_1440,N_1406);
xor U1508 (N_1508,N_1455,N_1432);
and U1509 (N_1509,N_1442,N_1417);
or U1510 (N_1510,N_1438,N_1463);
nor U1511 (N_1511,N_1429,N_1402);
nand U1512 (N_1512,N_1462,N_1436);
nand U1513 (N_1513,N_1477,N_1497);
nor U1514 (N_1514,N_1457,N_1461);
and U1515 (N_1515,N_1448,N_1420);
or U1516 (N_1516,N_1487,N_1493);
nand U1517 (N_1517,N_1486,N_1426);
or U1518 (N_1518,N_1435,N_1430);
and U1519 (N_1519,N_1449,N_1422);
or U1520 (N_1520,N_1444,N_1483);
or U1521 (N_1521,N_1445,N_1479);
nand U1522 (N_1522,N_1405,N_1467);
xnor U1523 (N_1523,N_1425,N_1439);
or U1524 (N_1524,N_1443,N_1466);
nand U1525 (N_1525,N_1476,N_1481);
and U1526 (N_1526,N_1418,N_1460);
or U1527 (N_1527,N_1424,N_1407);
and U1528 (N_1528,N_1419,N_1412);
or U1529 (N_1529,N_1496,N_1427);
nand U1530 (N_1530,N_1403,N_1452);
nand U1531 (N_1531,N_1453,N_1414);
or U1532 (N_1532,N_1416,N_1465);
and U1533 (N_1533,N_1456,N_1491);
and U1534 (N_1534,N_1433,N_1447);
nand U1535 (N_1535,N_1413,N_1421);
and U1536 (N_1536,N_1409,N_1464);
nor U1537 (N_1537,N_1446,N_1469);
or U1538 (N_1538,N_1485,N_1415);
and U1539 (N_1539,N_1489,N_1490);
nand U1540 (N_1540,N_1459,N_1400);
nand U1541 (N_1541,N_1408,N_1484);
nor U1542 (N_1542,N_1428,N_1499);
nand U1543 (N_1543,N_1450,N_1492);
and U1544 (N_1544,N_1451,N_1423);
nor U1545 (N_1545,N_1470,N_1454);
or U1546 (N_1546,N_1475,N_1458);
and U1547 (N_1547,N_1498,N_1488);
nor U1548 (N_1548,N_1410,N_1478);
or U1549 (N_1549,N_1473,N_1437);
and U1550 (N_1550,N_1420,N_1407);
and U1551 (N_1551,N_1420,N_1475);
nor U1552 (N_1552,N_1480,N_1451);
xor U1553 (N_1553,N_1460,N_1482);
or U1554 (N_1554,N_1415,N_1438);
or U1555 (N_1555,N_1451,N_1405);
nor U1556 (N_1556,N_1469,N_1473);
or U1557 (N_1557,N_1499,N_1449);
or U1558 (N_1558,N_1487,N_1412);
nor U1559 (N_1559,N_1475,N_1451);
nor U1560 (N_1560,N_1422,N_1484);
or U1561 (N_1561,N_1458,N_1484);
or U1562 (N_1562,N_1441,N_1435);
and U1563 (N_1563,N_1427,N_1456);
or U1564 (N_1564,N_1419,N_1455);
or U1565 (N_1565,N_1415,N_1434);
or U1566 (N_1566,N_1492,N_1493);
and U1567 (N_1567,N_1408,N_1473);
or U1568 (N_1568,N_1491,N_1457);
or U1569 (N_1569,N_1470,N_1472);
and U1570 (N_1570,N_1468,N_1474);
or U1571 (N_1571,N_1416,N_1432);
and U1572 (N_1572,N_1486,N_1460);
and U1573 (N_1573,N_1476,N_1427);
and U1574 (N_1574,N_1482,N_1405);
and U1575 (N_1575,N_1425,N_1404);
nor U1576 (N_1576,N_1467,N_1416);
nor U1577 (N_1577,N_1409,N_1405);
nand U1578 (N_1578,N_1464,N_1442);
xnor U1579 (N_1579,N_1430,N_1498);
nand U1580 (N_1580,N_1439,N_1483);
and U1581 (N_1581,N_1496,N_1466);
and U1582 (N_1582,N_1417,N_1473);
nor U1583 (N_1583,N_1485,N_1447);
xor U1584 (N_1584,N_1471,N_1424);
nor U1585 (N_1585,N_1437,N_1408);
nor U1586 (N_1586,N_1409,N_1407);
nand U1587 (N_1587,N_1489,N_1403);
nor U1588 (N_1588,N_1405,N_1459);
nor U1589 (N_1589,N_1486,N_1474);
or U1590 (N_1590,N_1434,N_1462);
xnor U1591 (N_1591,N_1456,N_1443);
and U1592 (N_1592,N_1460,N_1409);
nor U1593 (N_1593,N_1432,N_1427);
and U1594 (N_1594,N_1401,N_1402);
nand U1595 (N_1595,N_1431,N_1455);
and U1596 (N_1596,N_1490,N_1477);
nand U1597 (N_1597,N_1400,N_1426);
nand U1598 (N_1598,N_1416,N_1477);
xnor U1599 (N_1599,N_1487,N_1419);
and U1600 (N_1600,N_1502,N_1543);
nor U1601 (N_1601,N_1528,N_1516);
and U1602 (N_1602,N_1569,N_1529);
and U1603 (N_1603,N_1599,N_1521);
or U1604 (N_1604,N_1554,N_1522);
and U1605 (N_1605,N_1519,N_1570);
or U1606 (N_1606,N_1545,N_1583);
nand U1607 (N_1607,N_1547,N_1571);
nand U1608 (N_1608,N_1594,N_1596);
nand U1609 (N_1609,N_1588,N_1534);
nor U1610 (N_1610,N_1518,N_1532);
or U1611 (N_1611,N_1580,N_1506);
or U1612 (N_1612,N_1536,N_1514);
xnor U1613 (N_1613,N_1513,N_1559);
nand U1614 (N_1614,N_1579,N_1577);
nand U1615 (N_1615,N_1589,N_1560);
or U1616 (N_1616,N_1531,N_1568);
nor U1617 (N_1617,N_1558,N_1540);
nor U1618 (N_1618,N_1526,N_1578);
or U1619 (N_1619,N_1548,N_1517);
nand U1620 (N_1620,N_1525,N_1591);
and U1621 (N_1621,N_1562,N_1592);
xnor U1622 (N_1622,N_1505,N_1574);
nand U1623 (N_1623,N_1509,N_1550);
or U1624 (N_1624,N_1527,N_1551);
and U1625 (N_1625,N_1507,N_1561);
nand U1626 (N_1626,N_1564,N_1524);
nor U1627 (N_1627,N_1553,N_1535);
and U1628 (N_1628,N_1501,N_1555);
nand U1629 (N_1629,N_1576,N_1567);
and U1630 (N_1630,N_1539,N_1552);
nor U1631 (N_1631,N_1523,N_1504);
nand U1632 (N_1632,N_1508,N_1541);
nor U1633 (N_1633,N_1597,N_1520);
and U1634 (N_1634,N_1530,N_1581);
and U1635 (N_1635,N_1538,N_1546);
nor U1636 (N_1636,N_1586,N_1512);
nor U1637 (N_1637,N_1503,N_1587);
nor U1638 (N_1638,N_1582,N_1595);
or U1639 (N_1639,N_1533,N_1537);
nor U1640 (N_1640,N_1511,N_1549);
nand U1641 (N_1641,N_1585,N_1572);
nand U1642 (N_1642,N_1542,N_1590);
xor U1643 (N_1643,N_1557,N_1544);
or U1644 (N_1644,N_1575,N_1598);
and U1645 (N_1645,N_1563,N_1593);
and U1646 (N_1646,N_1515,N_1500);
nand U1647 (N_1647,N_1566,N_1565);
nor U1648 (N_1648,N_1584,N_1510);
and U1649 (N_1649,N_1573,N_1556);
nor U1650 (N_1650,N_1565,N_1584);
nand U1651 (N_1651,N_1586,N_1559);
nand U1652 (N_1652,N_1591,N_1558);
nand U1653 (N_1653,N_1504,N_1517);
or U1654 (N_1654,N_1503,N_1562);
nor U1655 (N_1655,N_1577,N_1515);
and U1656 (N_1656,N_1581,N_1550);
nor U1657 (N_1657,N_1503,N_1518);
and U1658 (N_1658,N_1504,N_1505);
nand U1659 (N_1659,N_1501,N_1551);
and U1660 (N_1660,N_1513,N_1574);
nand U1661 (N_1661,N_1574,N_1563);
and U1662 (N_1662,N_1530,N_1525);
nor U1663 (N_1663,N_1551,N_1553);
or U1664 (N_1664,N_1524,N_1540);
nand U1665 (N_1665,N_1546,N_1537);
nand U1666 (N_1666,N_1570,N_1542);
and U1667 (N_1667,N_1557,N_1506);
and U1668 (N_1668,N_1591,N_1585);
nor U1669 (N_1669,N_1519,N_1558);
nor U1670 (N_1670,N_1561,N_1504);
nor U1671 (N_1671,N_1505,N_1564);
xnor U1672 (N_1672,N_1503,N_1597);
nor U1673 (N_1673,N_1544,N_1529);
nand U1674 (N_1674,N_1572,N_1547);
nand U1675 (N_1675,N_1579,N_1555);
or U1676 (N_1676,N_1547,N_1552);
nand U1677 (N_1677,N_1563,N_1514);
nand U1678 (N_1678,N_1578,N_1513);
nor U1679 (N_1679,N_1532,N_1510);
and U1680 (N_1680,N_1548,N_1510);
nor U1681 (N_1681,N_1577,N_1524);
nand U1682 (N_1682,N_1536,N_1537);
nor U1683 (N_1683,N_1581,N_1516);
or U1684 (N_1684,N_1580,N_1543);
nor U1685 (N_1685,N_1555,N_1544);
and U1686 (N_1686,N_1562,N_1591);
and U1687 (N_1687,N_1519,N_1530);
or U1688 (N_1688,N_1513,N_1525);
and U1689 (N_1689,N_1544,N_1570);
nand U1690 (N_1690,N_1568,N_1583);
or U1691 (N_1691,N_1563,N_1579);
and U1692 (N_1692,N_1521,N_1551);
xnor U1693 (N_1693,N_1591,N_1530);
and U1694 (N_1694,N_1550,N_1517);
and U1695 (N_1695,N_1514,N_1517);
and U1696 (N_1696,N_1594,N_1583);
or U1697 (N_1697,N_1572,N_1593);
nor U1698 (N_1698,N_1552,N_1523);
and U1699 (N_1699,N_1552,N_1553);
nor U1700 (N_1700,N_1670,N_1635);
and U1701 (N_1701,N_1624,N_1656);
or U1702 (N_1702,N_1658,N_1645);
nor U1703 (N_1703,N_1662,N_1697);
nor U1704 (N_1704,N_1649,N_1600);
or U1705 (N_1705,N_1668,N_1696);
nor U1706 (N_1706,N_1628,N_1679);
and U1707 (N_1707,N_1673,N_1678);
nand U1708 (N_1708,N_1604,N_1691);
nand U1709 (N_1709,N_1699,N_1630);
and U1710 (N_1710,N_1616,N_1688);
or U1711 (N_1711,N_1605,N_1622);
nand U1712 (N_1712,N_1685,N_1666);
nor U1713 (N_1713,N_1633,N_1611);
and U1714 (N_1714,N_1634,N_1651);
nor U1715 (N_1715,N_1613,N_1626);
nor U1716 (N_1716,N_1674,N_1621);
or U1717 (N_1717,N_1639,N_1650);
xor U1718 (N_1718,N_1643,N_1655);
and U1719 (N_1719,N_1682,N_1676);
and U1720 (N_1720,N_1672,N_1661);
and U1721 (N_1721,N_1647,N_1606);
or U1722 (N_1722,N_1680,N_1664);
nand U1723 (N_1723,N_1687,N_1677);
or U1724 (N_1724,N_1637,N_1614);
nor U1725 (N_1725,N_1690,N_1623);
nor U1726 (N_1726,N_1636,N_1601);
nor U1727 (N_1727,N_1653,N_1654);
nor U1728 (N_1728,N_1612,N_1684);
nand U1729 (N_1729,N_1602,N_1669);
nand U1730 (N_1730,N_1686,N_1660);
nor U1731 (N_1731,N_1694,N_1652);
nand U1732 (N_1732,N_1619,N_1657);
nand U1733 (N_1733,N_1617,N_1648);
and U1734 (N_1734,N_1667,N_1608);
or U1735 (N_1735,N_1629,N_1610);
and U1736 (N_1736,N_1627,N_1620);
nor U1737 (N_1737,N_1659,N_1640);
and U1738 (N_1738,N_1644,N_1692);
and U1739 (N_1739,N_1609,N_1625);
or U1740 (N_1740,N_1698,N_1693);
nor U1741 (N_1741,N_1675,N_1665);
nand U1742 (N_1742,N_1695,N_1631);
and U1743 (N_1743,N_1671,N_1683);
or U1744 (N_1744,N_1618,N_1607);
nand U1745 (N_1745,N_1689,N_1642);
nand U1746 (N_1746,N_1603,N_1646);
nor U1747 (N_1747,N_1663,N_1641);
and U1748 (N_1748,N_1681,N_1638);
nand U1749 (N_1749,N_1615,N_1632);
nor U1750 (N_1750,N_1635,N_1623);
and U1751 (N_1751,N_1628,N_1654);
or U1752 (N_1752,N_1655,N_1672);
or U1753 (N_1753,N_1678,N_1633);
xnor U1754 (N_1754,N_1659,N_1671);
or U1755 (N_1755,N_1675,N_1608);
nor U1756 (N_1756,N_1692,N_1600);
nand U1757 (N_1757,N_1691,N_1617);
and U1758 (N_1758,N_1698,N_1682);
or U1759 (N_1759,N_1618,N_1659);
or U1760 (N_1760,N_1689,N_1630);
and U1761 (N_1761,N_1631,N_1648);
and U1762 (N_1762,N_1699,N_1683);
nor U1763 (N_1763,N_1613,N_1650);
or U1764 (N_1764,N_1603,N_1681);
and U1765 (N_1765,N_1684,N_1600);
nand U1766 (N_1766,N_1609,N_1643);
and U1767 (N_1767,N_1668,N_1618);
nand U1768 (N_1768,N_1639,N_1679);
and U1769 (N_1769,N_1631,N_1673);
nand U1770 (N_1770,N_1694,N_1650);
nand U1771 (N_1771,N_1614,N_1681);
nor U1772 (N_1772,N_1691,N_1697);
or U1773 (N_1773,N_1610,N_1648);
and U1774 (N_1774,N_1620,N_1619);
and U1775 (N_1775,N_1687,N_1661);
nand U1776 (N_1776,N_1693,N_1619);
and U1777 (N_1777,N_1671,N_1678);
and U1778 (N_1778,N_1614,N_1632);
and U1779 (N_1779,N_1638,N_1648);
nand U1780 (N_1780,N_1632,N_1683);
or U1781 (N_1781,N_1602,N_1682);
or U1782 (N_1782,N_1663,N_1646);
and U1783 (N_1783,N_1659,N_1644);
nor U1784 (N_1784,N_1684,N_1634);
and U1785 (N_1785,N_1635,N_1647);
nor U1786 (N_1786,N_1683,N_1652);
xor U1787 (N_1787,N_1687,N_1667);
and U1788 (N_1788,N_1678,N_1666);
and U1789 (N_1789,N_1611,N_1650);
and U1790 (N_1790,N_1677,N_1683);
nand U1791 (N_1791,N_1666,N_1611);
and U1792 (N_1792,N_1640,N_1645);
and U1793 (N_1793,N_1698,N_1662);
nor U1794 (N_1794,N_1628,N_1641);
xnor U1795 (N_1795,N_1621,N_1684);
or U1796 (N_1796,N_1641,N_1600);
nand U1797 (N_1797,N_1671,N_1636);
or U1798 (N_1798,N_1689,N_1670);
and U1799 (N_1799,N_1606,N_1632);
and U1800 (N_1800,N_1793,N_1711);
or U1801 (N_1801,N_1700,N_1740);
nor U1802 (N_1802,N_1703,N_1778);
and U1803 (N_1803,N_1741,N_1795);
and U1804 (N_1804,N_1717,N_1723);
nor U1805 (N_1805,N_1713,N_1704);
nand U1806 (N_1806,N_1785,N_1769);
nor U1807 (N_1807,N_1774,N_1777);
and U1808 (N_1808,N_1734,N_1766);
or U1809 (N_1809,N_1714,N_1798);
or U1810 (N_1810,N_1738,N_1782);
nand U1811 (N_1811,N_1780,N_1792);
nand U1812 (N_1812,N_1767,N_1771);
or U1813 (N_1813,N_1787,N_1721);
nand U1814 (N_1814,N_1705,N_1729);
or U1815 (N_1815,N_1761,N_1726);
nor U1816 (N_1816,N_1733,N_1745);
xnor U1817 (N_1817,N_1731,N_1790);
xor U1818 (N_1818,N_1765,N_1747);
and U1819 (N_1819,N_1779,N_1770);
or U1820 (N_1820,N_1756,N_1781);
and U1821 (N_1821,N_1737,N_1708);
and U1822 (N_1822,N_1716,N_1796);
nand U1823 (N_1823,N_1776,N_1742);
or U1824 (N_1824,N_1755,N_1743);
nand U1825 (N_1825,N_1728,N_1702);
xnor U1826 (N_1826,N_1754,N_1759);
nand U1827 (N_1827,N_1715,N_1752);
nand U1828 (N_1828,N_1749,N_1753);
and U1829 (N_1829,N_1763,N_1724);
or U1830 (N_1830,N_1748,N_1768);
or U1831 (N_1831,N_1797,N_1751);
nand U1832 (N_1832,N_1701,N_1718);
nand U1833 (N_1833,N_1773,N_1722);
nand U1834 (N_1834,N_1709,N_1746);
nor U1835 (N_1835,N_1791,N_1775);
and U1836 (N_1836,N_1744,N_1784);
or U1837 (N_1837,N_1730,N_1758);
and U1838 (N_1838,N_1783,N_1712);
or U1839 (N_1839,N_1739,N_1772);
nand U1840 (N_1840,N_1736,N_1750);
nand U1841 (N_1841,N_1710,N_1719);
nand U1842 (N_1842,N_1757,N_1732);
or U1843 (N_1843,N_1727,N_1707);
nand U1844 (N_1844,N_1706,N_1789);
xor U1845 (N_1845,N_1720,N_1725);
xnor U1846 (N_1846,N_1794,N_1764);
and U1847 (N_1847,N_1735,N_1786);
nor U1848 (N_1848,N_1762,N_1760);
nand U1849 (N_1849,N_1788,N_1799);
or U1850 (N_1850,N_1735,N_1737);
and U1851 (N_1851,N_1779,N_1797);
and U1852 (N_1852,N_1724,N_1771);
nor U1853 (N_1853,N_1727,N_1792);
nand U1854 (N_1854,N_1775,N_1782);
or U1855 (N_1855,N_1703,N_1768);
nor U1856 (N_1856,N_1710,N_1727);
and U1857 (N_1857,N_1727,N_1741);
nand U1858 (N_1858,N_1718,N_1790);
nor U1859 (N_1859,N_1717,N_1731);
nand U1860 (N_1860,N_1799,N_1733);
or U1861 (N_1861,N_1750,N_1730);
nand U1862 (N_1862,N_1729,N_1768);
nand U1863 (N_1863,N_1751,N_1726);
or U1864 (N_1864,N_1755,N_1749);
nor U1865 (N_1865,N_1733,N_1706);
nor U1866 (N_1866,N_1706,N_1737);
or U1867 (N_1867,N_1736,N_1760);
nor U1868 (N_1868,N_1787,N_1715);
or U1869 (N_1869,N_1720,N_1727);
xor U1870 (N_1870,N_1786,N_1725);
nand U1871 (N_1871,N_1746,N_1740);
nand U1872 (N_1872,N_1722,N_1739);
nand U1873 (N_1873,N_1795,N_1705);
nor U1874 (N_1874,N_1797,N_1777);
nand U1875 (N_1875,N_1740,N_1779);
nand U1876 (N_1876,N_1733,N_1759);
or U1877 (N_1877,N_1755,N_1787);
nand U1878 (N_1878,N_1777,N_1713);
or U1879 (N_1879,N_1744,N_1724);
nor U1880 (N_1880,N_1768,N_1707);
and U1881 (N_1881,N_1727,N_1721);
nand U1882 (N_1882,N_1749,N_1744);
nor U1883 (N_1883,N_1771,N_1738);
and U1884 (N_1884,N_1767,N_1788);
and U1885 (N_1885,N_1780,N_1727);
or U1886 (N_1886,N_1748,N_1771);
nand U1887 (N_1887,N_1720,N_1783);
and U1888 (N_1888,N_1724,N_1750);
or U1889 (N_1889,N_1771,N_1732);
and U1890 (N_1890,N_1722,N_1784);
and U1891 (N_1891,N_1708,N_1792);
and U1892 (N_1892,N_1748,N_1700);
xor U1893 (N_1893,N_1754,N_1765);
nand U1894 (N_1894,N_1728,N_1745);
nand U1895 (N_1895,N_1778,N_1784);
nor U1896 (N_1896,N_1777,N_1793);
nand U1897 (N_1897,N_1702,N_1766);
or U1898 (N_1898,N_1737,N_1751);
or U1899 (N_1899,N_1729,N_1762);
nand U1900 (N_1900,N_1827,N_1802);
nor U1901 (N_1901,N_1883,N_1847);
nand U1902 (N_1902,N_1892,N_1875);
or U1903 (N_1903,N_1870,N_1867);
nor U1904 (N_1904,N_1877,N_1894);
nand U1905 (N_1905,N_1860,N_1889);
or U1906 (N_1906,N_1817,N_1861);
nand U1907 (N_1907,N_1873,N_1813);
and U1908 (N_1908,N_1890,N_1898);
nand U1909 (N_1909,N_1800,N_1834);
and U1910 (N_1910,N_1872,N_1812);
and U1911 (N_1911,N_1830,N_1823);
or U1912 (N_1912,N_1869,N_1864);
nand U1913 (N_1913,N_1849,N_1824);
or U1914 (N_1914,N_1835,N_1833);
and U1915 (N_1915,N_1853,N_1806);
and U1916 (N_1916,N_1874,N_1855);
or U1917 (N_1917,N_1803,N_1895);
and U1918 (N_1918,N_1816,N_1819);
and U1919 (N_1919,N_1840,N_1815);
xnor U1920 (N_1920,N_1888,N_1859);
and U1921 (N_1921,N_1825,N_1871);
nand U1922 (N_1922,N_1887,N_1810);
nor U1923 (N_1923,N_1846,N_1868);
nand U1924 (N_1924,N_1856,N_1891);
and U1925 (N_1925,N_1826,N_1881);
or U1926 (N_1926,N_1879,N_1828);
nand U1927 (N_1927,N_1897,N_1808);
nand U1928 (N_1928,N_1899,N_1880);
nand U1929 (N_1929,N_1832,N_1852);
and U1930 (N_1930,N_1851,N_1893);
and U1931 (N_1931,N_1884,N_1822);
nor U1932 (N_1932,N_1804,N_1820);
nand U1933 (N_1933,N_1876,N_1896);
nor U1934 (N_1934,N_1845,N_1862);
nor U1935 (N_1935,N_1829,N_1885);
or U1936 (N_1936,N_1866,N_1837);
nand U1937 (N_1937,N_1882,N_1854);
xor U1938 (N_1938,N_1807,N_1858);
and U1939 (N_1939,N_1848,N_1811);
and U1940 (N_1940,N_1839,N_1821);
or U1941 (N_1941,N_1801,N_1842);
nand U1942 (N_1942,N_1843,N_1805);
nor U1943 (N_1943,N_1886,N_1831);
or U1944 (N_1944,N_1844,N_1850);
or U1945 (N_1945,N_1838,N_1809);
or U1946 (N_1946,N_1818,N_1863);
nand U1947 (N_1947,N_1841,N_1878);
nand U1948 (N_1948,N_1814,N_1836);
nand U1949 (N_1949,N_1865,N_1857);
and U1950 (N_1950,N_1898,N_1846);
and U1951 (N_1951,N_1823,N_1895);
or U1952 (N_1952,N_1829,N_1834);
or U1953 (N_1953,N_1812,N_1817);
or U1954 (N_1954,N_1883,N_1867);
or U1955 (N_1955,N_1860,N_1869);
or U1956 (N_1956,N_1874,N_1862);
nor U1957 (N_1957,N_1874,N_1898);
or U1958 (N_1958,N_1849,N_1865);
and U1959 (N_1959,N_1830,N_1899);
or U1960 (N_1960,N_1883,N_1827);
and U1961 (N_1961,N_1841,N_1863);
nor U1962 (N_1962,N_1815,N_1873);
and U1963 (N_1963,N_1806,N_1885);
and U1964 (N_1964,N_1817,N_1867);
nor U1965 (N_1965,N_1848,N_1851);
or U1966 (N_1966,N_1840,N_1882);
nand U1967 (N_1967,N_1857,N_1889);
or U1968 (N_1968,N_1804,N_1826);
xnor U1969 (N_1969,N_1808,N_1864);
nand U1970 (N_1970,N_1879,N_1812);
nor U1971 (N_1971,N_1845,N_1840);
nor U1972 (N_1972,N_1800,N_1824);
nor U1973 (N_1973,N_1806,N_1867);
nand U1974 (N_1974,N_1896,N_1855);
nand U1975 (N_1975,N_1805,N_1898);
or U1976 (N_1976,N_1806,N_1892);
nand U1977 (N_1977,N_1855,N_1862);
nand U1978 (N_1978,N_1826,N_1801);
nand U1979 (N_1979,N_1893,N_1831);
nand U1980 (N_1980,N_1856,N_1893);
nor U1981 (N_1981,N_1861,N_1880);
or U1982 (N_1982,N_1851,N_1876);
xnor U1983 (N_1983,N_1861,N_1829);
nor U1984 (N_1984,N_1833,N_1889);
and U1985 (N_1985,N_1866,N_1851);
or U1986 (N_1986,N_1876,N_1899);
nand U1987 (N_1987,N_1802,N_1808);
nor U1988 (N_1988,N_1866,N_1867);
nand U1989 (N_1989,N_1881,N_1847);
or U1990 (N_1990,N_1822,N_1836);
xor U1991 (N_1991,N_1843,N_1816);
nor U1992 (N_1992,N_1889,N_1884);
nor U1993 (N_1993,N_1817,N_1801);
or U1994 (N_1994,N_1879,N_1839);
or U1995 (N_1995,N_1839,N_1880);
or U1996 (N_1996,N_1823,N_1854);
nor U1997 (N_1997,N_1823,N_1892);
nand U1998 (N_1998,N_1899,N_1828);
nand U1999 (N_1999,N_1811,N_1869);
and U2000 (N_2000,N_1964,N_1966);
or U2001 (N_2001,N_1961,N_1942);
nor U2002 (N_2002,N_1923,N_1949);
xor U2003 (N_2003,N_1935,N_1977);
and U2004 (N_2004,N_1978,N_1919);
and U2005 (N_2005,N_1960,N_1957);
and U2006 (N_2006,N_1903,N_1946);
nor U2007 (N_2007,N_1995,N_1900);
nor U2008 (N_2008,N_1973,N_1908);
and U2009 (N_2009,N_1906,N_1941);
nor U2010 (N_2010,N_1974,N_1927);
xnor U2011 (N_2011,N_1948,N_1969);
nand U2012 (N_2012,N_1939,N_1918);
nor U2013 (N_2013,N_1956,N_1920);
or U2014 (N_2014,N_1965,N_1982);
or U2015 (N_2015,N_1975,N_1952);
nand U2016 (N_2016,N_1953,N_1909);
or U2017 (N_2017,N_1917,N_1922);
nor U2018 (N_2018,N_1929,N_1991);
nand U2019 (N_2019,N_1943,N_1968);
and U2020 (N_2020,N_1913,N_1998);
or U2021 (N_2021,N_1985,N_1902);
and U2022 (N_2022,N_1955,N_1981);
or U2023 (N_2023,N_1996,N_1915);
or U2024 (N_2024,N_1933,N_1931);
nand U2025 (N_2025,N_1962,N_1934);
nor U2026 (N_2026,N_1990,N_1901);
or U2027 (N_2027,N_1951,N_1992);
nor U2028 (N_2028,N_1936,N_1986);
and U2029 (N_2029,N_1938,N_1954);
xnor U2030 (N_2030,N_1967,N_1916);
or U2031 (N_2031,N_1993,N_1950);
nand U2032 (N_2032,N_1930,N_1921);
and U2033 (N_2033,N_1987,N_1972);
or U2034 (N_2034,N_1914,N_1937);
or U2035 (N_2035,N_1911,N_1976);
or U2036 (N_2036,N_1907,N_1988);
nor U2037 (N_2037,N_1926,N_1945);
and U2038 (N_2038,N_1925,N_1910);
and U2039 (N_2039,N_1983,N_1947);
and U2040 (N_2040,N_1963,N_1997);
nor U2041 (N_2041,N_1959,N_1958);
or U2042 (N_2042,N_1971,N_1994);
xor U2043 (N_2043,N_1904,N_1944);
and U2044 (N_2044,N_1980,N_1932);
nor U2045 (N_2045,N_1940,N_1970);
or U2046 (N_2046,N_1905,N_1984);
and U2047 (N_2047,N_1924,N_1989);
nand U2048 (N_2048,N_1999,N_1928);
and U2049 (N_2049,N_1912,N_1979);
and U2050 (N_2050,N_1924,N_1966);
and U2051 (N_2051,N_1926,N_1960);
or U2052 (N_2052,N_1976,N_1956);
nand U2053 (N_2053,N_1999,N_1910);
and U2054 (N_2054,N_1955,N_1940);
nor U2055 (N_2055,N_1971,N_1914);
or U2056 (N_2056,N_1967,N_1952);
nor U2057 (N_2057,N_1994,N_1987);
nand U2058 (N_2058,N_1941,N_1933);
nand U2059 (N_2059,N_1900,N_1912);
nand U2060 (N_2060,N_1904,N_1957);
and U2061 (N_2061,N_1923,N_1987);
and U2062 (N_2062,N_1922,N_1986);
nand U2063 (N_2063,N_1934,N_1941);
nor U2064 (N_2064,N_1946,N_1984);
and U2065 (N_2065,N_1989,N_1914);
nor U2066 (N_2066,N_1976,N_1928);
and U2067 (N_2067,N_1961,N_1945);
and U2068 (N_2068,N_1943,N_1969);
nor U2069 (N_2069,N_1926,N_1901);
nor U2070 (N_2070,N_1902,N_1919);
or U2071 (N_2071,N_1919,N_1913);
xnor U2072 (N_2072,N_1991,N_1987);
nand U2073 (N_2073,N_1979,N_1934);
nand U2074 (N_2074,N_1956,N_1984);
nor U2075 (N_2075,N_1978,N_1935);
or U2076 (N_2076,N_1916,N_1973);
or U2077 (N_2077,N_1924,N_1967);
nand U2078 (N_2078,N_1930,N_1980);
nand U2079 (N_2079,N_1909,N_1938);
nand U2080 (N_2080,N_1908,N_1937);
nand U2081 (N_2081,N_1954,N_1987);
nor U2082 (N_2082,N_1976,N_1926);
and U2083 (N_2083,N_1961,N_1916);
nand U2084 (N_2084,N_1931,N_1994);
nand U2085 (N_2085,N_1914,N_1955);
nor U2086 (N_2086,N_1943,N_1929);
nand U2087 (N_2087,N_1901,N_1946);
or U2088 (N_2088,N_1934,N_1983);
and U2089 (N_2089,N_1960,N_1903);
nor U2090 (N_2090,N_1950,N_1977);
nand U2091 (N_2091,N_1960,N_1974);
nor U2092 (N_2092,N_1901,N_1996);
and U2093 (N_2093,N_1999,N_1908);
nor U2094 (N_2094,N_1968,N_1973);
nor U2095 (N_2095,N_1971,N_1909);
or U2096 (N_2096,N_1936,N_1999);
nand U2097 (N_2097,N_1938,N_1983);
nand U2098 (N_2098,N_1978,N_1977);
and U2099 (N_2099,N_1955,N_1979);
nand U2100 (N_2100,N_2007,N_2002);
nand U2101 (N_2101,N_2053,N_2014);
and U2102 (N_2102,N_2030,N_2071);
nand U2103 (N_2103,N_2084,N_2097);
and U2104 (N_2104,N_2001,N_2093);
nand U2105 (N_2105,N_2036,N_2009);
and U2106 (N_2106,N_2033,N_2058);
nor U2107 (N_2107,N_2072,N_2065);
or U2108 (N_2108,N_2016,N_2087);
or U2109 (N_2109,N_2057,N_2079);
nor U2110 (N_2110,N_2035,N_2043);
or U2111 (N_2111,N_2067,N_2026);
or U2112 (N_2112,N_2069,N_2040);
nor U2113 (N_2113,N_2089,N_2078);
nor U2114 (N_2114,N_2077,N_2017);
nor U2115 (N_2115,N_2098,N_2099);
and U2116 (N_2116,N_2041,N_2024);
or U2117 (N_2117,N_2063,N_2042);
nor U2118 (N_2118,N_2010,N_2082);
and U2119 (N_2119,N_2039,N_2095);
nand U2120 (N_2120,N_2023,N_2013);
xor U2121 (N_2121,N_2019,N_2025);
or U2122 (N_2122,N_2032,N_2006);
and U2123 (N_2123,N_2031,N_2045);
nand U2124 (N_2124,N_2059,N_2088);
nand U2125 (N_2125,N_2076,N_2021);
nor U2126 (N_2126,N_2028,N_2056);
and U2127 (N_2127,N_2061,N_2055);
and U2128 (N_2128,N_2046,N_2049);
and U2129 (N_2129,N_2064,N_2060);
nand U2130 (N_2130,N_2073,N_2005);
nand U2131 (N_2131,N_2047,N_2081);
or U2132 (N_2132,N_2000,N_2054);
and U2133 (N_2133,N_2034,N_2074);
or U2134 (N_2134,N_2075,N_2094);
or U2135 (N_2135,N_2027,N_2004);
nor U2136 (N_2136,N_2050,N_2052);
and U2137 (N_2137,N_2048,N_2080);
nor U2138 (N_2138,N_2085,N_2070);
nand U2139 (N_2139,N_2068,N_2011);
nor U2140 (N_2140,N_2044,N_2022);
and U2141 (N_2141,N_2018,N_2086);
nand U2142 (N_2142,N_2015,N_2037);
nor U2143 (N_2143,N_2029,N_2051);
and U2144 (N_2144,N_2090,N_2038);
or U2145 (N_2145,N_2066,N_2020);
and U2146 (N_2146,N_2062,N_2096);
nor U2147 (N_2147,N_2092,N_2091);
nand U2148 (N_2148,N_2003,N_2008);
nor U2149 (N_2149,N_2012,N_2083);
or U2150 (N_2150,N_2028,N_2050);
nor U2151 (N_2151,N_2040,N_2032);
nor U2152 (N_2152,N_2049,N_2041);
nor U2153 (N_2153,N_2025,N_2018);
nand U2154 (N_2154,N_2091,N_2096);
or U2155 (N_2155,N_2070,N_2034);
or U2156 (N_2156,N_2048,N_2068);
or U2157 (N_2157,N_2027,N_2073);
nand U2158 (N_2158,N_2064,N_2000);
nor U2159 (N_2159,N_2064,N_2011);
and U2160 (N_2160,N_2020,N_2047);
nand U2161 (N_2161,N_2023,N_2008);
or U2162 (N_2162,N_2004,N_2053);
and U2163 (N_2163,N_2044,N_2031);
and U2164 (N_2164,N_2030,N_2033);
and U2165 (N_2165,N_2017,N_2069);
nand U2166 (N_2166,N_2032,N_2029);
nand U2167 (N_2167,N_2087,N_2098);
nor U2168 (N_2168,N_2038,N_2039);
or U2169 (N_2169,N_2009,N_2053);
nor U2170 (N_2170,N_2037,N_2097);
nor U2171 (N_2171,N_2050,N_2009);
nand U2172 (N_2172,N_2076,N_2027);
nor U2173 (N_2173,N_2040,N_2001);
nand U2174 (N_2174,N_2071,N_2044);
nand U2175 (N_2175,N_2038,N_2013);
nor U2176 (N_2176,N_2060,N_2078);
nor U2177 (N_2177,N_2019,N_2041);
nand U2178 (N_2178,N_2001,N_2021);
nor U2179 (N_2179,N_2051,N_2052);
nand U2180 (N_2180,N_2097,N_2073);
and U2181 (N_2181,N_2025,N_2077);
nand U2182 (N_2182,N_2072,N_2030);
nor U2183 (N_2183,N_2066,N_2069);
nand U2184 (N_2184,N_2016,N_2041);
nor U2185 (N_2185,N_2051,N_2043);
and U2186 (N_2186,N_2060,N_2015);
nor U2187 (N_2187,N_2063,N_2035);
or U2188 (N_2188,N_2003,N_2084);
and U2189 (N_2189,N_2020,N_2082);
or U2190 (N_2190,N_2086,N_2021);
and U2191 (N_2191,N_2062,N_2098);
nand U2192 (N_2192,N_2039,N_2013);
xor U2193 (N_2193,N_2068,N_2090);
and U2194 (N_2194,N_2087,N_2064);
or U2195 (N_2195,N_2083,N_2096);
or U2196 (N_2196,N_2070,N_2095);
or U2197 (N_2197,N_2033,N_2059);
and U2198 (N_2198,N_2006,N_2041);
nand U2199 (N_2199,N_2089,N_2098);
and U2200 (N_2200,N_2125,N_2192);
and U2201 (N_2201,N_2137,N_2126);
and U2202 (N_2202,N_2199,N_2139);
or U2203 (N_2203,N_2152,N_2108);
or U2204 (N_2204,N_2191,N_2165);
nor U2205 (N_2205,N_2194,N_2174);
nand U2206 (N_2206,N_2109,N_2101);
and U2207 (N_2207,N_2121,N_2130);
nor U2208 (N_2208,N_2124,N_2113);
or U2209 (N_2209,N_2164,N_2160);
nor U2210 (N_2210,N_2102,N_2143);
and U2211 (N_2211,N_2180,N_2112);
nor U2212 (N_2212,N_2140,N_2154);
or U2213 (N_2213,N_2127,N_2120);
xnor U2214 (N_2214,N_2155,N_2153);
or U2215 (N_2215,N_2158,N_2182);
or U2216 (N_2216,N_2106,N_2115);
and U2217 (N_2217,N_2144,N_2185);
or U2218 (N_2218,N_2161,N_2162);
or U2219 (N_2219,N_2147,N_2178);
and U2220 (N_2220,N_2173,N_2184);
and U2221 (N_2221,N_2189,N_2183);
or U2222 (N_2222,N_2169,N_2156);
nor U2223 (N_2223,N_2104,N_2151);
and U2224 (N_2224,N_2105,N_2188);
or U2225 (N_2225,N_2132,N_2146);
or U2226 (N_2226,N_2171,N_2122);
or U2227 (N_2227,N_2141,N_2129);
and U2228 (N_2228,N_2119,N_2145);
nor U2229 (N_2229,N_2172,N_2100);
nor U2230 (N_2230,N_2138,N_2163);
nor U2231 (N_2231,N_2167,N_2196);
nand U2232 (N_2232,N_2136,N_2116);
or U2233 (N_2233,N_2131,N_2193);
and U2234 (N_2234,N_2181,N_2114);
and U2235 (N_2235,N_2134,N_2133);
and U2236 (N_2236,N_2177,N_2179);
nor U2237 (N_2237,N_2128,N_2148);
and U2238 (N_2238,N_2157,N_2168);
and U2239 (N_2239,N_2118,N_2175);
or U2240 (N_2240,N_2159,N_2149);
nand U2241 (N_2241,N_2150,N_2187);
and U2242 (N_2242,N_2195,N_2111);
and U2243 (N_2243,N_2197,N_2103);
and U2244 (N_2244,N_2142,N_2198);
and U2245 (N_2245,N_2117,N_2190);
nor U2246 (N_2246,N_2110,N_2123);
nor U2247 (N_2247,N_2166,N_2107);
nor U2248 (N_2248,N_2176,N_2135);
nand U2249 (N_2249,N_2186,N_2170);
nand U2250 (N_2250,N_2107,N_2120);
nor U2251 (N_2251,N_2153,N_2192);
or U2252 (N_2252,N_2110,N_2139);
or U2253 (N_2253,N_2118,N_2148);
nor U2254 (N_2254,N_2115,N_2159);
and U2255 (N_2255,N_2179,N_2182);
xor U2256 (N_2256,N_2108,N_2172);
and U2257 (N_2257,N_2108,N_2146);
nor U2258 (N_2258,N_2181,N_2178);
nor U2259 (N_2259,N_2196,N_2171);
and U2260 (N_2260,N_2114,N_2151);
or U2261 (N_2261,N_2107,N_2171);
nor U2262 (N_2262,N_2119,N_2197);
nor U2263 (N_2263,N_2138,N_2136);
and U2264 (N_2264,N_2112,N_2106);
and U2265 (N_2265,N_2161,N_2143);
or U2266 (N_2266,N_2153,N_2145);
nand U2267 (N_2267,N_2121,N_2140);
nor U2268 (N_2268,N_2150,N_2133);
nand U2269 (N_2269,N_2122,N_2108);
nor U2270 (N_2270,N_2187,N_2165);
nor U2271 (N_2271,N_2183,N_2117);
and U2272 (N_2272,N_2192,N_2135);
or U2273 (N_2273,N_2113,N_2167);
nand U2274 (N_2274,N_2119,N_2113);
or U2275 (N_2275,N_2184,N_2158);
nand U2276 (N_2276,N_2120,N_2182);
or U2277 (N_2277,N_2154,N_2190);
nor U2278 (N_2278,N_2158,N_2117);
and U2279 (N_2279,N_2184,N_2167);
nor U2280 (N_2280,N_2194,N_2114);
nor U2281 (N_2281,N_2165,N_2164);
nor U2282 (N_2282,N_2196,N_2129);
nand U2283 (N_2283,N_2174,N_2186);
or U2284 (N_2284,N_2110,N_2128);
and U2285 (N_2285,N_2109,N_2164);
and U2286 (N_2286,N_2190,N_2116);
nor U2287 (N_2287,N_2102,N_2181);
and U2288 (N_2288,N_2105,N_2107);
nor U2289 (N_2289,N_2139,N_2137);
and U2290 (N_2290,N_2196,N_2108);
nor U2291 (N_2291,N_2176,N_2145);
and U2292 (N_2292,N_2138,N_2123);
and U2293 (N_2293,N_2140,N_2174);
or U2294 (N_2294,N_2181,N_2106);
nor U2295 (N_2295,N_2116,N_2198);
nor U2296 (N_2296,N_2155,N_2176);
and U2297 (N_2297,N_2157,N_2183);
nand U2298 (N_2298,N_2147,N_2137);
or U2299 (N_2299,N_2114,N_2199);
nand U2300 (N_2300,N_2245,N_2221);
nand U2301 (N_2301,N_2237,N_2270);
and U2302 (N_2302,N_2242,N_2203);
or U2303 (N_2303,N_2206,N_2251);
nor U2304 (N_2304,N_2285,N_2264);
nor U2305 (N_2305,N_2277,N_2220);
and U2306 (N_2306,N_2209,N_2298);
or U2307 (N_2307,N_2260,N_2223);
nor U2308 (N_2308,N_2282,N_2243);
nand U2309 (N_2309,N_2238,N_2248);
or U2310 (N_2310,N_2240,N_2293);
nand U2311 (N_2311,N_2274,N_2296);
nand U2312 (N_2312,N_2287,N_2257);
nor U2313 (N_2313,N_2273,N_2253);
nor U2314 (N_2314,N_2278,N_2275);
nand U2315 (N_2315,N_2241,N_2249);
nand U2316 (N_2316,N_2201,N_2266);
nand U2317 (N_2317,N_2267,N_2268);
and U2318 (N_2318,N_2219,N_2232);
nor U2319 (N_2319,N_2239,N_2231);
and U2320 (N_2320,N_2297,N_2292);
and U2321 (N_2321,N_2204,N_2288);
or U2322 (N_2322,N_2236,N_2263);
nor U2323 (N_2323,N_2217,N_2254);
nand U2324 (N_2324,N_2281,N_2207);
nand U2325 (N_2325,N_2289,N_2269);
nand U2326 (N_2326,N_2208,N_2228);
or U2327 (N_2327,N_2225,N_2256);
nor U2328 (N_2328,N_2234,N_2212);
and U2329 (N_2329,N_2290,N_2216);
nor U2330 (N_2330,N_2218,N_2222);
nor U2331 (N_2331,N_2230,N_2200);
nand U2332 (N_2332,N_2227,N_2244);
nand U2333 (N_2333,N_2246,N_2280);
nand U2334 (N_2334,N_2262,N_2283);
or U2335 (N_2335,N_2276,N_2291);
and U2336 (N_2336,N_2226,N_2265);
and U2337 (N_2337,N_2272,N_2271);
nor U2338 (N_2338,N_2255,N_2252);
nor U2339 (N_2339,N_2211,N_2233);
or U2340 (N_2340,N_2210,N_2202);
nand U2341 (N_2341,N_2299,N_2259);
and U2342 (N_2342,N_2284,N_2205);
and U2343 (N_2343,N_2215,N_2224);
nand U2344 (N_2344,N_2261,N_2235);
or U2345 (N_2345,N_2294,N_2214);
nor U2346 (N_2346,N_2250,N_2247);
nand U2347 (N_2347,N_2258,N_2213);
and U2348 (N_2348,N_2295,N_2279);
nand U2349 (N_2349,N_2229,N_2286);
and U2350 (N_2350,N_2282,N_2228);
or U2351 (N_2351,N_2202,N_2209);
xor U2352 (N_2352,N_2207,N_2267);
nor U2353 (N_2353,N_2233,N_2266);
xor U2354 (N_2354,N_2266,N_2240);
nand U2355 (N_2355,N_2257,N_2244);
and U2356 (N_2356,N_2272,N_2225);
and U2357 (N_2357,N_2220,N_2248);
nand U2358 (N_2358,N_2288,N_2290);
xnor U2359 (N_2359,N_2224,N_2201);
and U2360 (N_2360,N_2251,N_2222);
nand U2361 (N_2361,N_2224,N_2209);
nor U2362 (N_2362,N_2273,N_2248);
and U2363 (N_2363,N_2272,N_2224);
or U2364 (N_2364,N_2288,N_2265);
or U2365 (N_2365,N_2286,N_2262);
nand U2366 (N_2366,N_2295,N_2206);
nand U2367 (N_2367,N_2281,N_2227);
nand U2368 (N_2368,N_2264,N_2255);
or U2369 (N_2369,N_2217,N_2249);
or U2370 (N_2370,N_2283,N_2257);
nand U2371 (N_2371,N_2211,N_2292);
nand U2372 (N_2372,N_2291,N_2251);
nand U2373 (N_2373,N_2233,N_2210);
and U2374 (N_2374,N_2220,N_2299);
nor U2375 (N_2375,N_2269,N_2238);
or U2376 (N_2376,N_2218,N_2278);
nor U2377 (N_2377,N_2284,N_2279);
or U2378 (N_2378,N_2239,N_2228);
or U2379 (N_2379,N_2210,N_2212);
nand U2380 (N_2380,N_2205,N_2206);
xnor U2381 (N_2381,N_2234,N_2227);
nand U2382 (N_2382,N_2276,N_2299);
or U2383 (N_2383,N_2267,N_2209);
and U2384 (N_2384,N_2209,N_2295);
nand U2385 (N_2385,N_2261,N_2297);
and U2386 (N_2386,N_2293,N_2222);
and U2387 (N_2387,N_2269,N_2288);
or U2388 (N_2388,N_2254,N_2233);
nand U2389 (N_2389,N_2233,N_2228);
or U2390 (N_2390,N_2265,N_2273);
and U2391 (N_2391,N_2298,N_2269);
nor U2392 (N_2392,N_2232,N_2231);
nand U2393 (N_2393,N_2226,N_2250);
nand U2394 (N_2394,N_2247,N_2218);
nand U2395 (N_2395,N_2242,N_2249);
and U2396 (N_2396,N_2233,N_2271);
nand U2397 (N_2397,N_2283,N_2244);
nand U2398 (N_2398,N_2212,N_2203);
nor U2399 (N_2399,N_2208,N_2285);
or U2400 (N_2400,N_2381,N_2328);
nand U2401 (N_2401,N_2340,N_2362);
or U2402 (N_2402,N_2393,N_2317);
and U2403 (N_2403,N_2367,N_2390);
nand U2404 (N_2404,N_2392,N_2313);
or U2405 (N_2405,N_2350,N_2380);
and U2406 (N_2406,N_2332,N_2306);
and U2407 (N_2407,N_2398,N_2347);
or U2408 (N_2408,N_2324,N_2386);
or U2409 (N_2409,N_2315,N_2397);
xnor U2410 (N_2410,N_2389,N_2365);
or U2411 (N_2411,N_2366,N_2325);
xnor U2412 (N_2412,N_2327,N_2383);
nor U2413 (N_2413,N_2318,N_2391);
nand U2414 (N_2414,N_2333,N_2351);
nor U2415 (N_2415,N_2355,N_2312);
and U2416 (N_2416,N_2387,N_2395);
nor U2417 (N_2417,N_2336,N_2323);
nand U2418 (N_2418,N_2337,N_2378);
or U2419 (N_2419,N_2374,N_2379);
nor U2420 (N_2420,N_2341,N_2385);
or U2421 (N_2421,N_2349,N_2343);
xor U2422 (N_2422,N_2358,N_2310);
or U2423 (N_2423,N_2373,N_2384);
nand U2424 (N_2424,N_2322,N_2370);
or U2425 (N_2425,N_2348,N_2346);
nand U2426 (N_2426,N_2388,N_2334);
nor U2427 (N_2427,N_2308,N_2368);
nor U2428 (N_2428,N_2357,N_2371);
nor U2429 (N_2429,N_2302,N_2353);
or U2430 (N_2430,N_2309,N_2376);
and U2431 (N_2431,N_2305,N_2335);
and U2432 (N_2432,N_2356,N_2377);
or U2433 (N_2433,N_2320,N_2352);
nor U2434 (N_2434,N_2359,N_2360);
xor U2435 (N_2435,N_2339,N_2345);
nand U2436 (N_2436,N_2375,N_2319);
or U2437 (N_2437,N_2304,N_2314);
nor U2438 (N_2438,N_2331,N_2321);
xor U2439 (N_2439,N_2303,N_2369);
and U2440 (N_2440,N_2394,N_2329);
or U2441 (N_2441,N_2342,N_2300);
nand U2442 (N_2442,N_2344,N_2354);
or U2443 (N_2443,N_2361,N_2316);
nor U2444 (N_2444,N_2396,N_2382);
and U2445 (N_2445,N_2364,N_2399);
nor U2446 (N_2446,N_2326,N_2372);
nor U2447 (N_2447,N_2307,N_2338);
nand U2448 (N_2448,N_2330,N_2363);
nand U2449 (N_2449,N_2311,N_2301);
and U2450 (N_2450,N_2367,N_2363);
and U2451 (N_2451,N_2370,N_2324);
or U2452 (N_2452,N_2398,N_2362);
nor U2453 (N_2453,N_2395,N_2329);
nor U2454 (N_2454,N_2398,N_2381);
nand U2455 (N_2455,N_2397,N_2326);
nor U2456 (N_2456,N_2318,N_2394);
or U2457 (N_2457,N_2317,N_2341);
nor U2458 (N_2458,N_2331,N_2346);
and U2459 (N_2459,N_2372,N_2386);
nor U2460 (N_2460,N_2382,N_2344);
nor U2461 (N_2461,N_2309,N_2344);
nor U2462 (N_2462,N_2343,N_2397);
and U2463 (N_2463,N_2376,N_2360);
or U2464 (N_2464,N_2311,N_2381);
nand U2465 (N_2465,N_2388,N_2357);
and U2466 (N_2466,N_2369,N_2364);
nor U2467 (N_2467,N_2324,N_2368);
nand U2468 (N_2468,N_2334,N_2367);
and U2469 (N_2469,N_2324,N_2361);
nor U2470 (N_2470,N_2316,N_2367);
nor U2471 (N_2471,N_2341,N_2351);
or U2472 (N_2472,N_2306,N_2345);
nor U2473 (N_2473,N_2376,N_2322);
xor U2474 (N_2474,N_2359,N_2334);
and U2475 (N_2475,N_2309,N_2393);
or U2476 (N_2476,N_2312,N_2323);
nand U2477 (N_2477,N_2392,N_2399);
or U2478 (N_2478,N_2338,N_2358);
nor U2479 (N_2479,N_2368,N_2354);
xnor U2480 (N_2480,N_2337,N_2311);
nand U2481 (N_2481,N_2385,N_2353);
and U2482 (N_2482,N_2311,N_2365);
and U2483 (N_2483,N_2387,N_2376);
nand U2484 (N_2484,N_2338,N_2327);
nor U2485 (N_2485,N_2345,N_2346);
nand U2486 (N_2486,N_2308,N_2346);
or U2487 (N_2487,N_2302,N_2313);
or U2488 (N_2488,N_2333,N_2330);
nor U2489 (N_2489,N_2356,N_2315);
nand U2490 (N_2490,N_2354,N_2316);
nand U2491 (N_2491,N_2347,N_2357);
nor U2492 (N_2492,N_2376,N_2375);
or U2493 (N_2493,N_2337,N_2397);
nand U2494 (N_2494,N_2398,N_2373);
or U2495 (N_2495,N_2325,N_2377);
nand U2496 (N_2496,N_2391,N_2336);
and U2497 (N_2497,N_2348,N_2307);
nand U2498 (N_2498,N_2384,N_2363);
nor U2499 (N_2499,N_2378,N_2328);
nor U2500 (N_2500,N_2489,N_2432);
or U2501 (N_2501,N_2447,N_2407);
nor U2502 (N_2502,N_2416,N_2435);
and U2503 (N_2503,N_2470,N_2494);
nand U2504 (N_2504,N_2482,N_2459);
nand U2505 (N_2505,N_2428,N_2463);
and U2506 (N_2506,N_2423,N_2434);
or U2507 (N_2507,N_2491,N_2478);
or U2508 (N_2508,N_2448,N_2485);
nand U2509 (N_2509,N_2471,N_2467);
and U2510 (N_2510,N_2405,N_2497);
and U2511 (N_2511,N_2412,N_2465);
nand U2512 (N_2512,N_2411,N_2477);
or U2513 (N_2513,N_2444,N_2469);
and U2514 (N_2514,N_2484,N_2410);
xnor U2515 (N_2515,N_2453,N_2413);
nand U2516 (N_2516,N_2474,N_2409);
nor U2517 (N_2517,N_2454,N_2495);
and U2518 (N_2518,N_2402,N_2490);
and U2519 (N_2519,N_2424,N_2488);
or U2520 (N_2520,N_2401,N_2446);
nor U2521 (N_2521,N_2440,N_2403);
and U2522 (N_2522,N_2487,N_2451);
and U2523 (N_2523,N_2493,N_2457);
nand U2524 (N_2524,N_2473,N_2481);
or U2525 (N_2525,N_2452,N_2430);
or U2526 (N_2526,N_2449,N_2472);
and U2527 (N_2527,N_2422,N_2439);
nand U2528 (N_2528,N_2421,N_2420);
and U2529 (N_2529,N_2492,N_2414);
or U2530 (N_2530,N_2468,N_2475);
and U2531 (N_2531,N_2419,N_2427);
and U2532 (N_2532,N_2455,N_2404);
or U2533 (N_2533,N_2431,N_2479);
and U2534 (N_2534,N_2466,N_2462);
and U2535 (N_2535,N_2458,N_2417);
nand U2536 (N_2536,N_2499,N_2418);
and U2537 (N_2537,N_2456,N_2441);
nor U2538 (N_2538,N_2425,N_2464);
and U2539 (N_2539,N_2408,N_2429);
and U2540 (N_2540,N_2450,N_2442);
nand U2541 (N_2541,N_2406,N_2486);
nand U2542 (N_2542,N_2415,N_2480);
nor U2543 (N_2543,N_2443,N_2483);
xor U2544 (N_2544,N_2445,N_2436);
nand U2545 (N_2545,N_2460,N_2496);
and U2546 (N_2546,N_2461,N_2476);
nand U2547 (N_2547,N_2437,N_2400);
and U2548 (N_2548,N_2438,N_2498);
nand U2549 (N_2549,N_2433,N_2426);
and U2550 (N_2550,N_2459,N_2414);
or U2551 (N_2551,N_2456,N_2442);
nor U2552 (N_2552,N_2426,N_2450);
nor U2553 (N_2553,N_2494,N_2437);
nand U2554 (N_2554,N_2420,N_2407);
and U2555 (N_2555,N_2438,N_2430);
or U2556 (N_2556,N_2458,N_2403);
nor U2557 (N_2557,N_2437,N_2455);
and U2558 (N_2558,N_2429,N_2466);
nor U2559 (N_2559,N_2423,N_2471);
nand U2560 (N_2560,N_2476,N_2418);
nand U2561 (N_2561,N_2478,N_2490);
and U2562 (N_2562,N_2494,N_2462);
nand U2563 (N_2563,N_2425,N_2449);
and U2564 (N_2564,N_2443,N_2449);
nand U2565 (N_2565,N_2462,N_2413);
and U2566 (N_2566,N_2402,N_2462);
or U2567 (N_2567,N_2424,N_2432);
nor U2568 (N_2568,N_2428,N_2422);
or U2569 (N_2569,N_2405,N_2468);
nor U2570 (N_2570,N_2419,N_2420);
nor U2571 (N_2571,N_2404,N_2437);
or U2572 (N_2572,N_2497,N_2498);
nor U2573 (N_2573,N_2446,N_2489);
or U2574 (N_2574,N_2444,N_2448);
or U2575 (N_2575,N_2481,N_2485);
nor U2576 (N_2576,N_2420,N_2424);
nor U2577 (N_2577,N_2402,N_2415);
or U2578 (N_2578,N_2473,N_2434);
nand U2579 (N_2579,N_2445,N_2473);
and U2580 (N_2580,N_2427,N_2463);
nand U2581 (N_2581,N_2422,N_2406);
or U2582 (N_2582,N_2413,N_2479);
and U2583 (N_2583,N_2423,N_2405);
and U2584 (N_2584,N_2443,N_2405);
or U2585 (N_2585,N_2447,N_2483);
xor U2586 (N_2586,N_2482,N_2403);
and U2587 (N_2587,N_2413,N_2429);
nor U2588 (N_2588,N_2457,N_2434);
xor U2589 (N_2589,N_2457,N_2467);
nor U2590 (N_2590,N_2402,N_2450);
or U2591 (N_2591,N_2462,N_2493);
nor U2592 (N_2592,N_2489,N_2466);
and U2593 (N_2593,N_2481,N_2409);
or U2594 (N_2594,N_2442,N_2493);
nand U2595 (N_2595,N_2403,N_2489);
nand U2596 (N_2596,N_2435,N_2447);
and U2597 (N_2597,N_2414,N_2448);
and U2598 (N_2598,N_2431,N_2400);
and U2599 (N_2599,N_2479,N_2426);
and U2600 (N_2600,N_2579,N_2516);
nor U2601 (N_2601,N_2548,N_2510);
nand U2602 (N_2602,N_2526,N_2559);
nor U2603 (N_2603,N_2549,N_2582);
and U2604 (N_2604,N_2551,N_2508);
or U2605 (N_2605,N_2545,N_2547);
nor U2606 (N_2606,N_2598,N_2558);
and U2607 (N_2607,N_2538,N_2562);
nand U2608 (N_2608,N_2534,N_2500);
and U2609 (N_2609,N_2520,N_2536);
and U2610 (N_2610,N_2581,N_2573);
or U2611 (N_2611,N_2546,N_2568);
nand U2612 (N_2612,N_2530,N_2543);
nor U2613 (N_2613,N_2523,N_2586);
and U2614 (N_2614,N_2594,N_2511);
nor U2615 (N_2615,N_2599,N_2552);
or U2616 (N_2616,N_2576,N_2541);
or U2617 (N_2617,N_2565,N_2567);
nand U2618 (N_2618,N_2506,N_2553);
and U2619 (N_2619,N_2577,N_2585);
nand U2620 (N_2620,N_2560,N_2563);
nand U2621 (N_2621,N_2596,N_2580);
or U2622 (N_2622,N_2517,N_2504);
nand U2623 (N_2623,N_2509,N_2505);
or U2624 (N_2624,N_2525,N_2539);
nor U2625 (N_2625,N_2540,N_2529);
nor U2626 (N_2626,N_2589,N_2521);
nand U2627 (N_2627,N_2518,N_2519);
or U2628 (N_2628,N_2590,N_2593);
nand U2629 (N_2629,N_2595,N_2527);
nor U2630 (N_2630,N_2575,N_2592);
and U2631 (N_2631,N_2569,N_2515);
nand U2632 (N_2632,N_2564,N_2555);
and U2633 (N_2633,N_2556,N_2584);
and U2634 (N_2634,N_2561,N_2597);
nor U2635 (N_2635,N_2507,N_2542);
and U2636 (N_2636,N_2501,N_2566);
nand U2637 (N_2637,N_2570,N_2535);
nor U2638 (N_2638,N_2532,N_2578);
nor U2639 (N_2639,N_2557,N_2503);
nor U2640 (N_2640,N_2524,N_2588);
nor U2641 (N_2641,N_2583,N_2544);
nand U2642 (N_2642,N_2533,N_2574);
nand U2643 (N_2643,N_2522,N_2531);
nor U2644 (N_2644,N_2513,N_2512);
and U2645 (N_2645,N_2572,N_2571);
nand U2646 (N_2646,N_2591,N_2537);
nor U2647 (N_2647,N_2528,N_2514);
nand U2648 (N_2648,N_2587,N_2554);
or U2649 (N_2649,N_2502,N_2550);
and U2650 (N_2650,N_2521,N_2566);
or U2651 (N_2651,N_2582,N_2554);
nand U2652 (N_2652,N_2553,N_2564);
nor U2653 (N_2653,N_2585,N_2541);
nand U2654 (N_2654,N_2508,N_2528);
and U2655 (N_2655,N_2565,N_2532);
nand U2656 (N_2656,N_2581,N_2594);
or U2657 (N_2657,N_2518,N_2517);
or U2658 (N_2658,N_2533,N_2522);
nor U2659 (N_2659,N_2538,N_2593);
or U2660 (N_2660,N_2553,N_2598);
nor U2661 (N_2661,N_2507,N_2547);
or U2662 (N_2662,N_2519,N_2501);
or U2663 (N_2663,N_2558,N_2530);
nand U2664 (N_2664,N_2573,N_2549);
or U2665 (N_2665,N_2581,N_2561);
nand U2666 (N_2666,N_2528,N_2583);
and U2667 (N_2667,N_2560,N_2549);
and U2668 (N_2668,N_2596,N_2539);
and U2669 (N_2669,N_2575,N_2524);
nand U2670 (N_2670,N_2534,N_2559);
or U2671 (N_2671,N_2523,N_2508);
or U2672 (N_2672,N_2562,N_2570);
nor U2673 (N_2673,N_2571,N_2516);
nor U2674 (N_2674,N_2553,N_2500);
nor U2675 (N_2675,N_2542,N_2517);
nand U2676 (N_2676,N_2501,N_2598);
nand U2677 (N_2677,N_2575,N_2580);
xor U2678 (N_2678,N_2500,N_2516);
and U2679 (N_2679,N_2590,N_2549);
nand U2680 (N_2680,N_2550,N_2525);
nor U2681 (N_2681,N_2554,N_2569);
and U2682 (N_2682,N_2533,N_2541);
or U2683 (N_2683,N_2521,N_2586);
or U2684 (N_2684,N_2576,N_2552);
and U2685 (N_2685,N_2504,N_2544);
and U2686 (N_2686,N_2583,N_2587);
and U2687 (N_2687,N_2531,N_2516);
nand U2688 (N_2688,N_2593,N_2534);
and U2689 (N_2689,N_2564,N_2595);
and U2690 (N_2690,N_2561,N_2571);
and U2691 (N_2691,N_2575,N_2531);
or U2692 (N_2692,N_2570,N_2548);
or U2693 (N_2693,N_2577,N_2560);
nand U2694 (N_2694,N_2518,N_2503);
nor U2695 (N_2695,N_2572,N_2579);
nor U2696 (N_2696,N_2501,N_2595);
and U2697 (N_2697,N_2508,N_2566);
and U2698 (N_2698,N_2528,N_2504);
nand U2699 (N_2699,N_2585,N_2522);
or U2700 (N_2700,N_2650,N_2610);
or U2701 (N_2701,N_2632,N_2600);
or U2702 (N_2702,N_2624,N_2684);
nand U2703 (N_2703,N_2601,N_2682);
nand U2704 (N_2704,N_2667,N_2635);
nand U2705 (N_2705,N_2604,N_2665);
or U2706 (N_2706,N_2683,N_2607);
nor U2707 (N_2707,N_2660,N_2686);
or U2708 (N_2708,N_2664,N_2655);
and U2709 (N_2709,N_2688,N_2637);
xor U2710 (N_2710,N_2623,N_2649);
or U2711 (N_2711,N_2681,N_2657);
and U2712 (N_2712,N_2695,N_2697);
and U2713 (N_2713,N_2631,N_2689);
and U2714 (N_2714,N_2673,N_2612);
and U2715 (N_2715,N_2619,N_2617);
nor U2716 (N_2716,N_2616,N_2621);
nor U2717 (N_2717,N_2634,N_2652);
or U2718 (N_2718,N_2608,N_2620);
nand U2719 (N_2719,N_2696,N_2609);
nor U2720 (N_2720,N_2671,N_2685);
nor U2721 (N_2721,N_2691,N_2602);
or U2722 (N_2722,N_2653,N_2666);
and U2723 (N_2723,N_2692,N_2639);
nor U2724 (N_2724,N_2618,N_2614);
or U2725 (N_2725,N_2676,N_2641);
xnor U2726 (N_2726,N_2626,N_2611);
or U2727 (N_2727,N_2645,N_2669);
nor U2728 (N_2728,N_2663,N_2662);
nand U2729 (N_2729,N_2656,N_2613);
or U2730 (N_2730,N_2627,N_2605);
nand U2731 (N_2731,N_2625,N_2658);
nor U2732 (N_2732,N_2675,N_2698);
nor U2733 (N_2733,N_2678,N_2651);
nor U2734 (N_2734,N_2668,N_2638);
and U2735 (N_2735,N_2687,N_2647);
nand U2736 (N_2736,N_2661,N_2615);
or U2737 (N_2737,N_2674,N_2690);
and U2738 (N_2738,N_2636,N_2606);
nand U2739 (N_2739,N_2622,N_2699);
nand U2740 (N_2740,N_2640,N_2654);
nand U2741 (N_2741,N_2644,N_2677);
nor U2742 (N_2742,N_2633,N_2648);
or U2743 (N_2743,N_2643,N_2630);
and U2744 (N_2744,N_2680,N_2603);
nand U2745 (N_2745,N_2646,N_2672);
and U2746 (N_2746,N_2642,N_2693);
and U2747 (N_2747,N_2629,N_2670);
nor U2748 (N_2748,N_2694,N_2679);
or U2749 (N_2749,N_2659,N_2628);
nor U2750 (N_2750,N_2672,N_2648);
or U2751 (N_2751,N_2620,N_2631);
or U2752 (N_2752,N_2635,N_2689);
and U2753 (N_2753,N_2610,N_2683);
and U2754 (N_2754,N_2642,N_2602);
or U2755 (N_2755,N_2633,N_2675);
or U2756 (N_2756,N_2624,N_2618);
and U2757 (N_2757,N_2632,N_2618);
nor U2758 (N_2758,N_2657,N_2617);
and U2759 (N_2759,N_2687,N_2677);
and U2760 (N_2760,N_2631,N_2678);
nand U2761 (N_2761,N_2625,N_2672);
nand U2762 (N_2762,N_2632,N_2670);
nor U2763 (N_2763,N_2608,N_2643);
nand U2764 (N_2764,N_2686,N_2648);
nor U2765 (N_2765,N_2614,N_2615);
and U2766 (N_2766,N_2608,N_2653);
and U2767 (N_2767,N_2690,N_2695);
nand U2768 (N_2768,N_2609,N_2677);
and U2769 (N_2769,N_2681,N_2612);
and U2770 (N_2770,N_2658,N_2600);
nand U2771 (N_2771,N_2652,N_2673);
nand U2772 (N_2772,N_2604,N_2633);
nand U2773 (N_2773,N_2697,N_2647);
or U2774 (N_2774,N_2623,N_2643);
nand U2775 (N_2775,N_2636,N_2691);
and U2776 (N_2776,N_2617,N_2651);
or U2777 (N_2777,N_2694,N_2620);
nand U2778 (N_2778,N_2607,N_2622);
nand U2779 (N_2779,N_2621,N_2630);
nand U2780 (N_2780,N_2644,N_2637);
nand U2781 (N_2781,N_2687,N_2627);
nand U2782 (N_2782,N_2654,N_2682);
nand U2783 (N_2783,N_2603,N_2691);
nand U2784 (N_2784,N_2626,N_2652);
and U2785 (N_2785,N_2611,N_2629);
nand U2786 (N_2786,N_2609,N_2681);
nand U2787 (N_2787,N_2667,N_2611);
and U2788 (N_2788,N_2656,N_2660);
or U2789 (N_2789,N_2661,N_2650);
nand U2790 (N_2790,N_2660,N_2687);
or U2791 (N_2791,N_2682,N_2642);
or U2792 (N_2792,N_2638,N_2676);
nand U2793 (N_2793,N_2664,N_2638);
or U2794 (N_2794,N_2653,N_2603);
and U2795 (N_2795,N_2689,N_2665);
nor U2796 (N_2796,N_2664,N_2673);
or U2797 (N_2797,N_2682,N_2602);
and U2798 (N_2798,N_2655,N_2663);
or U2799 (N_2799,N_2606,N_2625);
or U2800 (N_2800,N_2781,N_2776);
and U2801 (N_2801,N_2730,N_2753);
nor U2802 (N_2802,N_2784,N_2747);
and U2803 (N_2803,N_2794,N_2721);
nand U2804 (N_2804,N_2704,N_2739);
or U2805 (N_2805,N_2765,N_2760);
nand U2806 (N_2806,N_2718,N_2745);
and U2807 (N_2807,N_2738,N_2716);
xnor U2808 (N_2808,N_2751,N_2795);
and U2809 (N_2809,N_2700,N_2740);
nor U2810 (N_2810,N_2702,N_2759);
and U2811 (N_2811,N_2722,N_2723);
nor U2812 (N_2812,N_2785,N_2779);
nand U2813 (N_2813,N_2772,N_2758);
or U2814 (N_2814,N_2742,N_2797);
and U2815 (N_2815,N_2725,N_2729);
nor U2816 (N_2816,N_2790,N_2769);
nand U2817 (N_2817,N_2706,N_2782);
nand U2818 (N_2818,N_2787,N_2791);
and U2819 (N_2819,N_2752,N_2703);
nand U2820 (N_2820,N_2728,N_2712);
nand U2821 (N_2821,N_2735,N_2707);
nor U2822 (N_2822,N_2720,N_2708);
nor U2823 (N_2823,N_2799,N_2770);
or U2824 (N_2824,N_2748,N_2749);
and U2825 (N_2825,N_2762,N_2793);
or U2826 (N_2826,N_2701,N_2789);
and U2827 (N_2827,N_2757,N_2746);
nor U2828 (N_2828,N_2744,N_2750);
and U2829 (N_2829,N_2768,N_2713);
nand U2830 (N_2830,N_2777,N_2775);
nand U2831 (N_2831,N_2788,N_2798);
and U2832 (N_2832,N_2705,N_2796);
xor U2833 (N_2833,N_2755,N_2754);
and U2834 (N_2834,N_2764,N_2724);
or U2835 (N_2835,N_2732,N_2743);
and U2836 (N_2836,N_2773,N_2778);
nand U2837 (N_2837,N_2715,N_2786);
and U2838 (N_2838,N_2726,N_2763);
and U2839 (N_2839,N_2719,N_2741);
nor U2840 (N_2840,N_2737,N_2792);
nor U2841 (N_2841,N_2774,N_2767);
nor U2842 (N_2842,N_2771,N_2717);
nor U2843 (N_2843,N_2727,N_2734);
nand U2844 (N_2844,N_2756,N_2733);
nand U2845 (N_2845,N_2761,N_2783);
nand U2846 (N_2846,N_2710,N_2731);
nor U2847 (N_2847,N_2736,N_2711);
nor U2848 (N_2848,N_2714,N_2780);
and U2849 (N_2849,N_2766,N_2709);
or U2850 (N_2850,N_2785,N_2700);
or U2851 (N_2851,N_2744,N_2756);
or U2852 (N_2852,N_2712,N_2718);
or U2853 (N_2853,N_2765,N_2732);
nand U2854 (N_2854,N_2741,N_2793);
nand U2855 (N_2855,N_2739,N_2738);
nor U2856 (N_2856,N_2723,N_2798);
or U2857 (N_2857,N_2791,N_2799);
nor U2858 (N_2858,N_2779,N_2763);
nand U2859 (N_2859,N_2771,N_2733);
nand U2860 (N_2860,N_2777,N_2798);
or U2861 (N_2861,N_2713,N_2712);
nor U2862 (N_2862,N_2779,N_2781);
nand U2863 (N_2863,N_2738,N_2755);
or U2864 (N_2864,N_2709,N_2759);
or U2865 (N_2865,N_2787,N_2751);
xor U2866 (N_2866,N_2769,N_2725);
or U2867 (N_2867,N_2776,N_2712);
or U2868 (N_2868,N_2730,N_2783);
or U2869 (N_2869,N_2746,N_2720);
or U2870 (N_2870,N_2746,N_2778);
nand U2871 (N_2871,N_2730,N_2760);
and U2872 (N_2872,N_2708,N_2779);
or U2873 (N_2873,N_2776,N_2788);
and U2874 (N_2874,N_2789,N_2707);
or U2875 (N_2875,N_2730,N_2715);
nor U2876 (N_2876,N_2725,N_2782);
nor U2877 (N_2877,N_2733,N_2760);
nand U2878 (N_2878,N_2718,N_2765);
and U2879 (N_2879,N_2710,N_2705);
nand U2880 (N_2880,N_2711,N_2752);
and U2881 (N_2881,N_2746,N_2716);
xnor U2882 (N_2882,N_2754,N_2717);
or U2883 (N_2883,N_2747,N_2769);
and U2884 (N_2884,N_2792,N_2794);
nor U2885 (N_2885,N_2714,N_2705);
or U2886 (N_2886,N_2793,N_2740);
or U2887 (N_2887,N_2744,N_2776);
nand U2888 (N_2888,N_2782,N_2761);
and U2889 (N_2889,N_2715,N_2773);
nand U2890 (N_2890,N_2774,N_2784);
nand U2891 (N_2891,N_2701,N_2787);
nor U2892 (N_2892,N_2723,N_2771);
nand U2893 (N_2893,N_2789,N_2775);
nor U2894 (N_2894,N_2729,N_2794);
or U2895 (N_2895,N_2775,N_2788);
nand U2896 (N_2896,N_2763,N_2783);
nor U2897 (N_2897,N_2715,N_2737);
xor U2898 (N_2898,N_2765,N_2738);
nor U2899 (N_2899,N_2701,N_2752);
and U2900 (N_2900,N_2859,N_2888);
or U2901 (N_2901,N_2869,N_2872);
and U2902 (N_2902,N_2808,N_2829);
nor U2903 (N_2903,N_2825,N_2819);
nor U2904 (N_2904,N_2827,N_2890);
nor U2905 (N_2905,N_2842,N_2867);
and U2906 (N_2906,N_2856,N_2866);
nand U2907 (N_2907,N_2857,N_2870);
and U2908 (N_2908,N_2868,N_2881);
nand U2909 (N_2909,N_2811,N_2886);
nand U2910 (N_2910,N_2839,N_2863);
nand U2911 (N_2911,N_2826,N_2802);
nand U2912 (N_2912,N_2899,N_2845);
or U2913 (N_2913,N_2891,N_2816);
and U2914 (N_2914,N_2847,N_2836);
nand U2915 (N_2915,N_2882,N_2851);
and U2916 (N_2916,N_2805,N_2848);
nand U2917 (N_2917,N_2879,N_2835);
xor U2918 (N_2918,N_2806,N_2804);
nor U2919 (N_2919,N_2817,N_2850);
nor U2920 (N_2920,N_2831,N_2852);
or U2921 (N_2921,N_2821,N_2801);
nand U2922 (N_2922,N_2858,N_2897);
nor U2923 (N_2923,N_2815,N_2889);
nor U2924 (N_2924,N_2840,N_2885);
and U2925 (N_2925,N_2873,N_2834);
or U2926 (N_2926,N_2832,N_2828);
nand U2927 (N_2927,N_2853,N_2824);
or U2928 (N_2928,N_2895,N_2864);
or U2929 (N_2929,N_2841,N_2818);
nor U2930 (N_2930,N_2896,N_2855);
and U2931 (N_2931,N_2862,N_2875);
or U2932 (N_2932,N_2878,N_2844);
or U2933 (N_2933,N_2830,N_2813);
nand U2934 (N_2934,N_2894,N_2838);
or U2935 (N_2935,N_2860,N_2800);
nor U2936 (N_2936,N_2849,N_2874);
xor U2937 (N_2937,N_2837,N_2861);
or U2938 (N_2938,N_2898,N_2820);
nor U2939 (N_2939,N_2871,N_2883);
or U2940 (N_2940,N_2876,N_2865);
or U2941 (N_2941,N_2803,N_2822);
or U2942 (N_2942,N_2810,N_2812);
nand U2943 (N_2943,N_2807,N_2884);
or U2944 (N_2944,N_2823,N_2880);
nor U2945 (N_2945,N_2814,N_2809);
nor U2946 (N_2946,N_2843,N_2887);
or U2947 (N_2947,N_2833,N_2877);
nand U2948 (N_2948,N_2892,N_2893);
and U2949 (N_2949,N_2854,N_2846);
nor U2950 (N_2950,N_2835,N_2820);
nand U2951 (N_2951,N_2855,N_2885);
nand U2952 (N_2952,N_2844,N_2813);
xnor U2953 (N_2953,N_2828,N_2892);
nor U2954 (N_2954,N_2886,N_2802);
nand U2955 (N_2955,N_2854,N_2899);
nor U2956 (N_2956,N_2851,N_2830);
nand U2957 (N_2957,N_2892,N_2817);
or U2958 (N_2958,N_2898,N_2801);
and U2959 (N_2959,N_2804,N_2865);
nand U2960 (N_2960,N_2836,N_2818);
or U2961 (N_2961,N_2813,N_2895);
and U2962 (N_2962,N_2834,N_2801);
nor U2963 (N_2963,N_2856,N_2807);
nor U2964 (N_2964,N_2814,N_2807);
nand U2965 (N_2965,N_2879,N_2860);
nor U2966 (N_2966,N_2884,N_2849);
xnor U2967 (N_2967,N_2814,N_2826);
nand U2968 (N_2968,N_2812,N_2878);
and U2969 (N_2969,N_2892,N_2867);
nand U2970 (N_2970,N_2853,N_2802);
or U2971 (N_2971,N_2886,N_2819);
or U2972 (N_2972,N_2807,N_2836);
nor U2973 (N_2973,N_2869,N_2803);
nor U2974 (N_2974,N_2859,N_2803);
xor U2975 (N_2975,N_2893,N_2888);
nand U2976 (N_2976,N_2854,N_2872);
nor U2977 (N_2977,N_2866,N_2884);
nand U2978 (N_2978,N_2830,N_2872);
xor U2979 (N_2979,N_2842,N_2852);
and U2980 (N_2980,N_2856,N_2877);
or U2981 (N_2981,N_2834,N_2857);
nand U2982 (N_2982,N_2830,N_2806);
nand U2983 (N_2983,N_2876,N_2846);
nand U2984 (N_2984,N_2881,N_2857);
and U2985 (N_2985,N_2878,N_2891);
nand U2986 (N_2986,N_2822,N_2807);
xnor U2987 (N_2987,N_2869,N_2810);
and U2988 (N_2988,N_2878,N_2862);
and U2989 (N_2989,N_2860,N_2867);
nand U2990 (N_2990,N_2863,N_2879);
and U2991 (N_2991,N_2875,N_2872);
and U2992 (N_2992,N_2847,N_2844);
nor U2993 (N_2993,N_2890,N_2826);
or U2994 (N_2994,N_2880,N_2834);
or U2995 (N_2995,N_2867,N_2854);
and U2996 (N_2996,N_2842,N_2800);
and U2997 (N_2997,N_2823,N_2831);
or U2998 (N_2998,N_2811,N_2825);
and U2999 (N_2999,N_2866,N_2800);
nor U3000 (N_3000,N_2906,N_2907);
or U3001 (N_3001,N_2961,N_2989);
nor U3002 (N_3002,N_2995,N_2946);
nor U3003 (N_3003,N_2918,N_2978);
nand U3004 (N_3004,N_2936,N_2986);
and U3005 (N_3005,N_2937,N_2925);
or U3006 (N_3006,N_2968,N_2956);
and U3007 (N_3007,N_2940,N_2941);
nor U3008 (N_3008,N_2972,N_2900);
nand U3009 (N_3009,N_2947,N_2950);
nor U3010 (N_3010,N_2911,N_2929);
nor U3011 (N_3011,N_2930,N_2966);
and U3012 (N_3012,N_2970,N_2903);
nor U3013 (N_3013,N_2938,N_2928);
or U3014 (N_3014,N_2908,N_2943);
and U3015 (N_3015,N_2902,N_2931);
and U3016 (N_3016,N_2951,N_2987);
or U3017 (N_3017,N_2960,N_2959);
and U3018 (N_3018,N_2957,N_2990);
nor U3019 (N_3019,N_2975,N_2965);
nor U3020 (N_3020,N_2953,N_2915);
nor U3021 (N_3021,N_2998,N_2922);
nor U3022 (N_3022,N_2955,N_2916);
nand U3023 (N_3023,N_2949,N_2919);
and U3024 (N_3024,N_2923,N_2969);
nor U3025 (N_3025,N_2948,N_2981);
or U3026 (N_3026,N_2927,N_2997);
nor U3027 (N_3027,N_2985,N_2991);
or U3028 (N_3028,N_2952,N_2934);
or U3029 (N_3029,N_2958,N_2994);
and U3030 (N_3030,N_2914,N_2942);
nand U3031 (N_3031,N_2973,N_2904);
xor U3032 (N_3032,N_2912,N_2976);
nand U3033 (N_3033,N_2963,N_2993);
xor U3034 (N_3034,N_2984,N_2982);
nor U3035 (N_3035,N_2996,N_2910);
nand U3036 (N_3036,N_2974,N_2962);
and U3037 (N_3037,N_2920,N_2980);
nor U3038 (N_3038,N_2905,N_2979);
nand U3039 (N_3039,N_2935,N_2945);
and U3040 (N_3040,N_2932,N_2901);
and U3041 (N_3041,N_2924,N_2999);
and U3042 (N_3042,N_2964,N_2926);
and U3043 (N_3043,N_2917,N_2954);
and U3044 (N_3044,N_2921,N_2944);
nand U3045 (N_3045,N_2913,N_2971);
and U3046 (N_3046,N_2983,N_2909);
nor U3047 (N_3047,N_2967,N_2977);
or U3048 (N_3048,N_2939,N_2933);
nand U3049 (N_3049,N_2992,N_2988);
and U3050 (N_3050,N_2973,N_2965);
or U3051 (N_3051,N_2917,N_2913);
or U3052 (N_3052,N_2943,N_2961);
or U3053 (N_3053,N_2940,N_2963);
or U3054 (N_3054,N_2926,N_2942);
and U3055 (N_3055,N_2917,N_2973);
and U3056 (N_3056,N_2952,N_2979);
or U3057 (N_3057,N_2993,N_2905);
nand U3058 (N_3058,N_2946,N_2991);
and U3059 (N_3059,N_2915,N_2911);
or U3060 (N_3060,N_2949,N_2954);
and U3061 (N_3061,N_2986,N_2924);
or U3062 (N_3062,N_2942,N_2917);
nand U3063 (N_3063,N_2937,N_2948);
nand U3064 (N_3064,N_2977,N_2910);
nand U3065 (N_3065,N_2907,N_2989);
nand U3066 (N_3066,N_2925,N_2927);
nand U3067 (N_3067,N_2999,N_2931);
xor U3068 (N_3068,N_2975,N_2995);
nand U3069 (N_3069,N_2985,N_2957);
and U3070 (N_3070,N_2950,N_2960);
nand U3071 (N_3071,N_2900,N_2930);
nor U3072 (N_3072,N_2941,N_2956);
and U3073 (N_3073,N_2949,N_2930);
nor U3074 (N_3074,N_2956,N_2985);
nand U3075 (N_3075,N_2987,N_2969);
or U3076 (N_3076,N_2912,N_2924);
nand U3077 (N_3077,N_2903,N_2906);
or U3078 (N_3078,N_2967,N_2973);
nand U3079 (N_3079,N_2970,N_2995);
nand U3080 (N_3080,N_2954,N_2981);
and U3081 (N_3081,N_2914,N_2925);
nor U3082 (N_3082,N_2939,N_2976);
nand U3083 (N_3083,N_2959,N_2951);
and U3084 (N_3084,N_2938,N_2924);
and U3085 (N_3085,N_2943,N_2916);
nor U3086 (N_3086,N_2948,N_2980);
and U3087 (N_3087,N_2988,N_2932);
and U3088 (N_3088,N_2909,N_2962);
and U3089 (N_3089,N_2947,N_2936);
nand U3090 (N_3090,N_2977,N_2965);
nand U3091 (N_3091,N_2977,N_2958);
and U3092 (N_3092,N_2967,N_2991);
nor U3093 (N_3093,N_2937,N_2907);
xnor U3094 (N_3094,N_2946,N_2992);
or U3095 (N_3095,N_2930,N_2982);
nand U3096 (N_3096,N_2989,N_2954);
and U3097 (N_3097,N_2950,N_2962);
nor U3098 (N_3098,N_2913,N_2938);
nand U3099 (N_3099,N_2964,N_2912);
or U3100 (N_3100,N_3093,N_3044);
nor U3101 (N_3101,N_3096,N_3089);
and U3102 (N_3102,N_3055,N_3019);
nor U3103 (N_3103,N_3039,N_3078);
nand U3104 (N_3104,N_3016,N_3068);
or U3105 (N_3105,N_3061,N_3099);
nand U3106 (N_3106,N_3015,N_3037);
xor U3107 (N_3107,N_3080,N_3018);
and U3108 (N_3108,N_3077,N_3069);
or U3109 (N_3109,N_3053,N_3084);
and U3110 (N_3110,N_3074,N_3057);
and U3111 (N_3111,N_3064,N_3028);
nor U3112 (N_3112,N_3088,N_3027);
nand U3113 (N_3113,N_3030,N_3000);
or U3114 (N_3114,N_3052,N_3009);
or U3115 (N_3115,N_3058,N_3004);
and U3116 (N_3116,N_3091,N_3050);
nor U3117 (N_3117,N_3014,N_3083);
nor U3118 (N_3118,N_3040,N_3070);
and U3119 (N_3119,N_3081,N_3076);
nand U3120 (N_3120,N_3048,N_3001);
nor U3121 (N_3121,N_3042,N_3003);
nor U3122 (N_3122,N_3063,N_3094);
or U3123 (N_3123,N_3007,N_3033);
or U3124 (N_3124,N_3060,N_3002);
and U3125 (N_3125,N_3022,N_3087);
or U3126 (N_3126,N_3034,N_3082);
xor U3127 (N_3127,N_3097,N_3046);
or U3128 (N_3128,N_3059,N_3073);
or U3129 (N_3129,N_3056,N_3035);
nand U3130 (N_3130,N_3049,N_3013);
nor U3131 (N_3131,N_3086,N_3006);
nand U3132 (N_3132,N_3010,N_3023);
and U3133 (N_3133,N_3026,N_3036);
or U3134 (N_3134,N_3067,N_3072);
or U3135 (N_3135,N_3085,N_3017);
and U3136 (N_3136,N_3062,N_3054);
nor U3137 (N_3137,N_3098,N_3071);
nand U3138 (N_3138,N_3038,N_3045);
and U3139 (N_3139,N_3025,N_3079);
and U3140 (N_3140,N_3075,N_3065);
nor U3141 (N_3141,N_3051,N_3047);
or U3142 (N_3142,N_3066,N_3029);
nand U3143 (N_3143,N_3092,N_3024);
nand U3144 (N_3144,N_3032,N_3031);
nor U3145 (N_3145,N_3012,N_3005);
or U3146 (N_3146,N_3090,N_3095);
nand U3147 (N_3147,N_3008,N_3011);
and U3148 (N_3148,N_3020,N_3041);
or U3149 (N_3149,N_3021,N_3043);
nor U3150 (N_3150,N_3080,N_3088);
xnor U3151 (N_3151,N_3028,N_3095);
nor U3152 (N_3152,N_3067,N_3005);
nor U3153 (N_3153,N_3069,N_3098);
or U3154 (N_3154,N_3014,N_3088);
nand U3155 (N_3155,N_3085,N_3043);
and U3156 (N_3156,N_3093,N_3025);
and U3157 (N_3157,N_3040,N_3029);
or U3158 (N_3158,N_3069,N_3078);
nor U3159 (N_3159,N_3011,N_3057);
or U3160 (N_3160,N_3082,N_3087);
or U3161 (N_3161,N_3066,N_3088);
and U3162 (N_3162,N_3071,N_3024);
nand U3163 (N_3163,N_3083,N_3055);
nand U3164 (N_3164,N_3030,N_3029);
and U3165 (N_3165,N_3081,N_3096);
and U3166 (N_3166,N_3053,N_3063);
nand U3167 (N_3167,N_3058,N_3073);
and U3168 (N_3168,N_3038,N_3087);
nor U3169 (N_3169,N_3011,N_3065);
nor U3170 (N_3170,N_3039,N_3066);
and U3171 (N_3171,N_3000,N_3036);
nor U3172 (N_3172,N_3066,N_3061);
or U3173 (N_3173,N_3084,N_3072);
and U3174 (N_3174,N_3039,N_3058);
and U3175 (N_3175,N_3088,N_3054);
xor U3176 (N_3176,N_3012,N_3042);
nor U3177 (N_3177,N_3025,N_3009);
nand U3178 (N_3178,N_3078,N_3050);
and U3179 (N_3179,N_3076,N_3016);
xnor U3180 (N_3180,N_3046,N_3013);
nand U3181 (N_3181,N_3009,N_3033);
nor U3182 (N_3182,N_3094,N_3004);
or U3183 (N_3183,N_3085,N_3057);
or U3184 (N_3184,N_3039,N_3064);
or U3185 (N_3185,N_3059,N_3068);
nand U3186 (N_3186,N_3051,N_3046);
and U3187 (N_3187,N_3088,N_3030);
or U3188 (N_3188,N_3002,N_3094);
nor U3189 (N_3189,N_3011,N_3084);
nand U3190 (N_3190,N_3065,N_3026);
and U3191 (N_3191,N_3097,N_3091);
and U3192 (N_3192,N_3027,N_3064);
nor U3193 (N_3193,N_3056,N_3009);
or U3194 (N_3194,N_3015,N_3096);
nand U3195 (N_3195,N_3005,N_3026);
nor U3196 (N_3196,N_3051,N_3049);
and U3197 (N_3197,N_3092,N_3022);
nand U3198 (N_3198,N_3081,N_3070);
nand U3199 (N_3199,N_3054,N_3066);
nand U3200 (N_3200,N_3138,N_3104);
or U3201 (N_3201,N_3133,N_3171);
nand U3202 (N_3202,N_3111,N_3153);
or U3203 (N_3203,N_3178,N_3145);
or U3204 (N_3204,N_3136,N_3164);
or U3205 (N_3205,N_3193,N_3137);
nor U3206 (N_3206,N_3198,N_3119);
nor U3207 (N_3207,N_3156,N_3143);
nand U3208 (N_3208,N_3194,N_3184);
nand U3209 (N_3209,N_3157,N_3146);
nand U3210 (N_3210,N_3185,N_3165);
nand U3211 (N_3211,N_3160,N_3162);
or U3212 (N_3212,N_3181,N_3106);
nor U3213 (N_3213,N_3199,N_3112);
and U3214 (N_3214,N_3100,N_3115);
or U3215 (N_3215,N_3192,N_3182);
or U3216 (N_3216,N_3109,N_3187);
xor U3217 (N_3217,N_3150,N_3188);
and U3218 (N_3218,N_3173,N_3159);
nand U3219 (N_3219,N_3113,N_3129);
or U3220 (N_3220,N_3121,N_3183);
and U3221 (N_3221,N_3147,N_3167);
and U3222 (N_3222,N_3132,N_3124);
or U3223 (N_3223,N_3120,N_3176);
and U3224 (N_3224,N_3148,N_3102);
nor U3225 (N_3225,N_3174,N_3128);
and U3226 (N_3226,N_3114,N_3131);
or U3227 (N_3227,N_3170,N_3149);
nand U3228 (N_3228,N_3186,N_3158);
or U3229 (N_3229,N_3126,N_3155);
or U3230 (N_3230,N_3175,N_3168);
and U3231 (N_3231,N_3135,N_3172);
or U3232 (N_3232,N_3134,N_3130);
or U3233 (N_3233,N_3141,N_3118);
and U3234 (N_3234,N_3161,N_3169);
and U3235 (N_3235,N_3179,N_3108);
nand U3236 (N_3236,N_3196,N_3177);
xnor U3237 (N_3237,N_3140,N_3125);
nor U3238 (N_3238,N_3152,N_3122);
nand U3239 (N_3239,N_3117,N_3189);
xnor U3240 (N_3240,N_3144,N_3197);
or U3241 (N_3241,N_3116,N_3190);
nor U3242 (N_3242,N_3123,N_3166);
nand U3243 (N_3243,N_3154,N_3105);
nor U3244 (N_3244,N_3142,N_3195);
or U3245 (N_3245,N_3139,N_3191);
nor U3246 (N_3246,N_3151,N_3180);
nand U3247 (N_3247,N_3163,N_3103);
nand U3248 (N_3248,N_3107,N_3110);
nand U3249 (N_3249,N_3127,N_3101);
or U3250 (N_3250,N_3133,N_3112);
or U3251 (N_3251,N_3143,N_3155);
or U3252 (N_3252,N_3179,N_3123);
nor U3253 (N_3253,N_3129,N_3135);
nand U3254 (N_3254,N_3137,N_3126);
nand U3255 (N_3255,N_3142,N_3175);
nand U3256 (N_3256,N_3154,N_3199);
nor U3257 (N_3257,N_3162,N_3157);
nor U3258 (N_3258,N_3128,N_3184);
nand U3259 (N_3259,N_3101,N_3166);
and U3260 (N_3260,N_3133,N_3136);
or U3261 (N_3261,N_3139,N_3138);
nand U3262 (N_3262,N_3166,N_3127);
or U3263 (N_3263,N_3106,N_3171);
and U3264 (N_3264,N_3106,N_3199);
nand U3265 (N_3265,N_3193,N_3183);
nor U3266 (N_3266,N_3132,N_3102);
and U3267 (N_3267,N_3114,N_3126);
nor U3268 (N_3268,N_3118,N_3134);
nand U3269 (N_3269,N_3147,N_3120);
nor U3270 (N_3270,N_3197,N_3173);
or U3271 (N_3271,N_3133,N_3124);
nand U3272 (N_3272,N_3156,N_3118);
or U3273 (N_3273,N_3137,N_3100);
nor U3274 (N_3274,N_3123,N_3195);
or U3275 (N_3275,N_3167,N_3108);
or U3276 (N_3276,N_3129,N_3187);
and U3277 (N_3277,N_3174,N_3175);
or U3278 (N_3278,N_3185,N_3121);
and U3279 (N_3279,N_3197,N_3112);
nand U3280 (N_3280,N_3113,N_3140);
and U3281 (N_3281,N_3166,N_3109);
or U3282 (N_3282,N_3170,N_3107);
xor U3283 (N_3283,N_3135,N_3158);
or U3284 (N_3284,N_3181,N_3129);
or U3285 (N_3285,N_3185,N_3173);
nor U3286 (N_3286,N_3146,N_3126);
nor U3287 (N_3287,N_3102,N_3159);
or U3288 (N_3288,N_3105,N_3125);
nand U3289 (N_3289,N_3141,N_3110);
or U3290 (N_3290,N_3128,N_3126);
nor U3291 (N_3291,N_3179,N_3142);
and U3292 (N_3292,N_3144,N_3137);
nor U3293 (N_3293,N_3188,N_3152);
nand U3294 (N_3294,N_3111,N_3132);
and U3295 (N_3295,N_3154,N_3126);
nand U3296 (N_3296,N_3117,N_3121);
or U3297 (N_3297,N_3170,N_3106);
nor U3298 (N_3298,N_3187,N_3140);
nor U3299 (N_3299,N_3185,N_3149);
nand U3300 (N_3300,N_3266,N_3209);
nor U3301 (N_3301,N_3274,N_3220);
and U3302 (N_3302,N_3207,N_3256);
nor U3303 (N_3303,N_3296,N_3286);
nor U3304 (N_3304,N_3257,N_3270);
and U3305 (N_3305,N_3239,N_3252);
or U3306 (N_3306,N_3201,N_3290);
or U3307 (N_3307,N_3234,N_3268);
and U3308 (N_3308,N_3240,N_3203);
nor U3309 (N_3309,N_3253,N_3284);
and U3310 (N_3310,N_3247,N_3244);
or U3311 (N_3311,N_3227,N_3219);
and U3312 (N_3312,N_3226,N_3200);
xnor U3313 (N_3313,N_3213,N_3288);
nand U3314 (N_3314,N_3229,N_3235);
nand U3315 (N_3315,N_3275,N_3269);
nor U3316 (N_3316,N_3242,N_3254);
nor U3317 (N_3317,N_3230,N_3285);
and U3318 (N_3318,N_3211,N_3264);
and U3319 (N_3319,N_3204,N_3221);
or U3320 (N_3320,N_3214,N_3251);
nand U3321 (N_3321,N_3293,N_3261);
nand U3322 (N_3322,N_3263,N_3238);
nor U3323 (N_3323,N_3262,N_3278);
and U3324 (N_3324,N_3218,N_3250);
nor U3325 (N_3325,N_3231,N_3280);
nand U3326 (N_3326,N_3271,N_3297);
or U3327 (N_3327,N_3210,N_3259);
and U3328 (N_3328,N_3249,N_3291);
or U3329 (N_3329,N_3292,N_3289);
nand U3330 (N_3330,N_3237,N_3279);
nor U3331 (N_3331,N_3287,N_3298);
and U3332 (N_3332,N_3265,N_3258);
nand U3333 (N_3333,N_3243,N_3248);
and U3334 (N_3334,N_3255,N_3276);
or U3335 (N_3335,N_3224,N_3245);
xnor U3336 (N_3336,N_3222,N_3212);
or U3337 (N_3337,N_3217,N_3208);
or U3338 (N_3338,N_3241,N_3294);
or U3339 (N_3339,N_3246,N_3205);
nor U3340 (N_3340,N_3216,N_3295);
nand U3341 (N_3341,N_3283,N_3273);
nand U3342 (N_3342,N_3232,N_3202);
or U3343 (N_3343,N_3260,N_3299);
nand U3344 (N_3344,N_3282,N_3277);
and U3345 (N_3345,N_3228,N_3267);
nor U3346 (N_3346,N_3233,N_3225);
nor U3347 (N_3347,N_3206,N_3223);
nor U3348 (N_3348,N_3236,N_3272);
nand U3349 (N_3349,N_3215,N_3281);
and U3350 (N_3350,N_3284,N_3277);
nor U3351 (N_3351,N_3282,N_3268);
or U3352 (N_3352,N_3268,N_3261);
and U3353 (N_3353,N_3292,N_3259);
or U3354 (N_3354,N_3283,N_3240);
or U3355 (N_3355,N_3294,N_3260);
nand U3356 (N_3356,N_3213,N_3216);
and U3357 (N_3357,N_3280,N_3258);
and U3358 (N_3358,N_3215,N_3210);
nor U3359 (N_3359,N_3296,N_3292);
and U3360 (N_3360,N_3280,N_3278);
and U3361 (N_3361,N_3239,N_3277);
nor U3362 (N_3362,N_3299,N_3288);
or U3363 (N_3363,N_3237,N_3218);
nor U3364 (N_3364,N_3299,N_3251);
nand U3365 (N_3365,N_3267,N_3278);
or U3366 (N_3366,N_3290,N_3247);
nand U3367 (N_3367,N_3296,N_3298);
nand U3368 (N_3368,N_3295,N_3292);
xnor U3369 (N_3369,N_3241,N_3245);
and U3370 (N_3370,N_3202,N_3214);
nor U3371 (N_3371,N_3211,N_3246);
nand U3372 (N_3372,N_3248,N_3272);
or U3373 (N_3373,N_3292,N_3266);
nor U3374 (N_3374,N_3236,N_3208);
nand U3375 (N_3375,N_3225,N_3206);
nand U3376 (N_3376,N_3287,N_3278);
nor U3377 (N_3377,N_3217,N_3222);
xnor U3378 (N_3378,N_3210,N_3240);
nand U3379 (N_3379,N_3262,N_3246);
and U3380 (N_3380,N_3204,N_3220);
nand U3381 (N_3381,N_3221,N_3251);
or U3382 (N_3382,N_3233,N_3295);
and U3383 (N_3383,N_3222,N_3210);
nand U3384 (N_3384,N_3256,N_3258);
and U3385 (N_3385,N_3265,N_3236);
or U3386 (N_3386,N_3253,N_3283);
nand U3387 (N_3387,N_3299,N_3274);
or U3388 (N_3388,N_3203,N_3272);
or U3389 (N_3389,N_3225,N_3220);
nor U3390 (N_3390,N_3246,N_3242);
or U3391 (N_3391,N_3247,N_3228);
nand U3392 (N_3392,N_3267,N_3235);
nor U3393 (N_3393,N_3200,N_3259);
nand U3394 (N_3394,N_3276,N_3208);
and U3395 (N_3395,N_3273,N_3236);
nor U3396 (N_3396,N_3202,N_3250);
or U3397 (N_3397,N_3232,N_3278);
nor U3398 (N_3398,N_3286,N_3248);
and U3399 (N_3399,N_3221,N_3281);
nor U3400 (N_3400,N_3320,N_3381);
and U3401 (N_3401,N_3359,N_3383);
or U3402 (N_3402,N_3350,N_3343);
and U3403 (N_3403,N_3384,N_3395);
nor U3404 (N_3404,N_3339,N_3329);
or U3405 (N_3405,N_3304,N_3382);
and U3406 (N_3406,N_3313,N_3327);
nand U3407 (N_3407,N_3371,N_3365);
nand U3408 (N_3408,N_3314,N_3335);
nand U3409 (N_3409,N_3363,N_3390);
or U3410 (N_3410,N_3328,N_3333);
and U3411 (N_3411,N_3379,N_3348);
and U3412 (N_3412,N_3388,N_3345);
or U3413 (N_3413,N_3394,N_3337);
or U3414 (N_3414,N_3300,N_3370);
and U3415 (N_3415,N_3369,N_3342);
or U3416 (N_3416,N_3357,N_3316);
nor U3417 (N_3417,N_3354,N_3308);
nor U3418 (N_3418,N_3336,N_3380);
or U3419 (N_3419,N_3302,N_3374);
and U3420 (N_3420,N_3311,N_3331);
nand U3421 (N_3421,N_3301,N_3346);
nor U3422 (N_3422,N_3325,N_3397);
nor U3423 (N_3423,N_3378,N_3355);
nor U3424 (N_3424,N_3385,N_3368);
and U3425 (N_3425,N_3367,N_3372);
nor U3426 (N_3426,N_3373,N_3347);
and U3427 (N_3427,N_3340,N_3366);
and U3428 (N_3428,N_3332,N_3360);
nand U3429 (N_3429,N_3389,N_3376);
or U3430 (N_3430,N_3353,N_3392);
and U3431 (N_3431,N_3303,N_3334);
nor U3432 (N_3432,N_3393,N_3375);
nand U3433 (N_3433,N_3306,N_3344);
nand U3434 (N_3434,N_3312,N_3351);
and U3435 (N_3435,N_3358,N_3361);
or U3436 (N_3436,N_3307,N_3323);
and U3437 (N_3437,N_3362,N_3387);
nand U3438 (N_3438,N_3396,N_3364);
nor U3439 (N_3439,N_3356,N_3386);
nor U3440 (N_3440,N_3398,N_3352);
nor U3441 (N_3441,N_3341,N_3319);
nor U3442 (N_3442,N_3330,N_3326);
and U3443 (N_3443,N_3324,N_3318);
and U3444 (N_3444,N_3321,N_3399);
nand U3445 (N_3445,N_3309,N_3322);
xor U3446 (N_3446,N_3349,N_3391);
or U3447 (N_3447,N_3377,N_3315);
nand U3448 (N_3448,N_3310,N_3317);
or U3449 (N_3449,N_3338,N_3305);
nand U3450 (N_3450,N_3372,N_3301);
or U3451 (N_3451,N_3366,N_3352);
nor U3452 (N_3452,N_3364,N_3308);
nor U3453 (N_3453,N_3308,N_3317);
and U3454 (N_3454,N_3398,N_3364);
or U3455 (N_3455,N_3348,N_3334);
and U3456 (N_3456,N_3312,N_3336);
and U3457 (N_3457,N_3322,N_3396);
nor U3458 (N_3458,N_3375,N_3335);
or U3459 (N_3459,N_3391,N_3367);
nand U3460 (N_3460,N_3395,N_3380);
nand U3461 (N_3461,N_3363,N_3376);
nor U3462 (N_3462,N_3308,N_3383);
or U3463 (N_3463,N_3347,N_3313);
or U3464 (N_3464,N_3330,N_3357);
nor U3465 (N_3465,N_3372,N_3321);
and U3466 (N_3466,N_3313,N_3363);
nand U3467 (N_3467,N_3359,N_3314);
and U3468 (N_3468,N_3346,N_3347);
or U3469 (N_3469,N_3333,N_3352);
nor U3470 (N_3470,N_3341,N_3390);
and U3471 (N_3471,N_3338,N_3339);
or U3472 (N_3472,N_3315,N_3348);
and U3473 (N_3473,N_3380,N_3333);
nand U3474 (N_3474,N_3307,N_3316);
nor U3475 (N_3475,N_3338,N_3341);
or U3476 (N_3476,N_3379,N_3383);
or U3477 (N_3477,N_3367,N_3360);
and U3478 (N_3478,N_3341,N_3343);
nor U3479 (N_3479,N_3314,N_3343);
or U3480 (N_3480,N_3371,N_3398);
and U3481 (N_3481,N_3360,N_3321);
nor U3482 (N_3482,N_3389,N_3306);
or U3483 (N_3483,N_3376,N_3384);
and U3484 (N_3484,N_3315,N_3392);
nor U3485 (N_3485,N_3307,N_3312);
or U3486 (N_3486,N_3361,N_3335);
nand U3487 (N_3487,N_3309,N_3314);
nor U3488 (N_3488,N_3332,N_3364);
nand U3489 (N_3489,N_3347,N_3395);
or U3490 (N_3490,N_3344,N_3395);
nand U3491 (N_3491,N_3300,N_3337);
nand U3492 (N_3492,N_3326,N_3301);
nand U3493 (N_3493,N_3305,N_3383);
nand U3494 (N_3494,N_3378,N_3309);
or U3495 (N_3495,N_3382,N_3360);
nor U3496 (N_3496,N_3369,N_3304);
or U3497 (N_3497,N_3357,N_3313);
nand U3498 (N_3498,N_3379,N_3338);
and U3499 (N_3499,N_3348,N_3325);
and U3500 (N_3500,N_3446,N_3445);
nand U3501 (N_3501,N_3470,N_3415);
nand U3502 (N_3502,N_3427,N_3426);
nor U3503 (N_3503,N_3480,N_3410);
and U3504 (N_3504,N_3412,N_3498);
or U3505 (N_3505,N_3494,N_3423);
nor U3506 (N_3506,N_3497,N_3452);
or U3507 (N_3507,N_3419,N_3424);
or U3508 (N_3508,N_3425,N_3443);
and U3509 (N_3509,N_3431,N_3486);
xor U3510 (N_3510,N_3441,N_3409);
xnor U3511 (N_3511,N_3400,N_3459);
nor U3512 (N_3512,N_3422,N_3428);
and U3513 (N_3513,N_3457,N_3477);
or U3514 (N_3514,N_3456,N_3491);
nand U3515 (N_3515,N_3478,N_3436);
nor U3516 (N_3516,N_3416,N_3453);
nor U3517 (N_3517,N_3458,N_3449);
nor U3518 (N_3518,N_3430,N_3421);
or U3519 (N_3519,N_3466,N_3489);
or U3520 (N_3520,N_3434,N_3493);
nor U3521 (N_3521,N_3495,N_3476);
nand U3522 (N_3522,N_3487,N_3469);
nand U3523 (N_3523,N_3488,N_3467);
nor U3524 (N_3524,N_3461,N_3448);
nand U3525 (N_3525,N_3439,N_3414);
nand U3526 (N_3526,N_3462,N_3442);
and U3527 (N_3527,N_3429,N_3435);
or U3528 (N_3528,N_3483,N_3482);
or U3529 (N_3529,N_3432,N_3451);
nor U3530 (N_3530,N_3411,N_3472);
nor U3531 (N_3531,N_3479,N_3481);
and U3532 (N_3532,N_3499,N_3454);
nor U3533 (N_3533,N_3455,N_3468);
nand U3534 (N_3534,N_3401,N_3471);
nand U3535 (N_3535,N_3420,N_3417);
or U3536 (N_3536,N_3496,N_3402);
nor U3537 (N_3537,N_3463,N_3464);
and U3538 (N_3538,N_3460,N_3485);
nand U3539 (N_3539,N_3447,N_3484);
or U3540 (N_3540,N_3440,N_3465);
or U3541 (N_3541,N_3444,N_3404);
and U3542 (N_3542,N_3418,N_3437);
and U3543 (N_3543,N_3413,N_3433);
nand U3544 (N_3544,N_3403,N_3406);
nand U3545 (N_3545,N_3405,N_3490);
nand U3546 (N_3546,N_3450,N_3408);
or U3547 (N_3547,N_3473,N_3492);
and U3548 (N_3548,N_3474,N_3407);
and U3549 (N_3549,N_3438,N_3475);
and U3550 (N_3550,N_3494,N_3465);
or U3551 (N_3551,N_3430,N_3419);
nand U3552 (N_3552,N_3453,N_3496);
or U3553 (N_3553,N_3469,N_3429);
nand U3554 (N_3554,N_3472,N_3463);
nand U3555 (N_3555,N_3449,N_3407);
nand U3556 (N_3556,N_3445,N_3415);
or U3557 (N_3557,N_3465,N_3431);
or U3558 (N_3558,N_3463,N_3413);
nand U3559 (N_3559,N_3458,N_3444);
nand U3560 (N_3560,N_3483,N_3441);
nor U3561 (N_3561,N_3442,N_3446);
nor U3562 (N_3562,N_3457,N_3486);
or U3563 (N_3563,N_3467,N_3497);
nand U3564 (N_3564,N_3428,N_3438);
or U3565 (N_3565,N_3481,N_3416);
nor U3566 (N_3566,N_3452,N_3400);
nand U3567 (N_3567,N_3454,N_3439);
nand U3568 (N_3568,N_3481,N_3442);
or U3569 (N_3569,N_3431,N_3489);
or U3570 (N_3570,N_3402,N_3456);
nand U3571 (N_3571,N_3480,N_3443);
nand U3572 (N_3572,N_3412,N_3474);
or U3573 (N_3573,N_3441,N_3482);
or U3574 (N_3574,N_3424,N_3441);
nor U3575 (N_3575,N_3455,N_3467);
nand U3576 (N_3576,N_3463,N_3474);
nor U3577 (N_3577,N_3474,N_3403);
nand U3578 (N_3578,N_3462,N_3452);
nand U3579 (N_3579,N_3426,N_3445);
nand U3580 (N_3580,N_3478,N_3426);
nand U3581 (N_3581,N_3423,N_3408);
and U3582 (N_3582,N_3444,N_3485);
nand U3583 (N_3583,N_3402,N_3436);
or U3584 (N_3584,N_3467,N_3474);
nand U3585 (N_3585,N_3423,N_3434);
or U3586 (N_3586,N_3438,N_3424);
and U3587 (N_3587,N_3487,N_3453);
nand U3588 (N_3588,N_3431,N_3495);
and U3589 (N_3589,N_3459,N_3458);
xor U3590 (N_3590,N_3435,N_3472);
and U3591 (N_3591,N_3401,N_3466);
nor U3592 (N_3592,N_3442,N_3456);
nor U3593 (N_3593,N_3459,N_3454);
nor U3594 (N_3594,N_3454,N_3461);
nor U3595 (N_3595,N_3483,N_3492);
nand U3596 (N_3596,N_3494,N_3403);
or U3597 (N_3597,N_3482,N_3464);
nand U3598 (N_3598,N_3411,N_3438);
nand U3599 (N_3599,N_3415,N_3482);
or U3600 (N_3600,N_3580,N_3530);
nor U3601 (N_3601,N_3559,N_3593);
and U3602 (N_3602,N_3592,N_3578);
or U3603 (N_3603,N_3587,N_3534);
nand U3604 (N_3604,N_3591,N_3549);
or U3605 (N_3605,N_3537,N_3569);
or U3606 (N_3606,N_3566,N_3515);
or U3607 (N_3607,N_3507,N_3539);
or U3608 (N_3608,N_3511,N_3532);
or U3609 (N_3609,N_3518,N_3519);
nand U3610 (N_3610,N_3528,N_3586);
nor U3611 (N_3611,N_3563,N_3513);
nor U3612 (N_3612,N_3582,N_3536);
and U3613 (N_3613,N_3547,N_3523);
nor U3614 (N_3614,N_3508,N_3502);
and U3615 (N_3615,N_3505,N_3581);
nor U3616 (N_3616,N_3520,N_3521);
nand U3617 (N_3617,N_3542,N_3571);
and U3618 (N_3618,N_3583,N_3576);
nor U3619 (N_3619,N_3510,N_3585);
nand U3620 (N_3620,N_3522,N_3565);
nand U3621 (N_3621,N_3567,N_3554);
nand U3622 (N_3622,N_3541,N_3500);
nor U3623 (N_3623,N_3527,N_3538);
nor U3624 (N_3624,N_3535,N_3589);
nand U3625 (N_3625,N_3560,N_3551);
and U3626 (N_3626,N_3543,N_3552);
and U3627 (N_3627,N_3562,N_3597);
nor U3628 (N_3628,N_3540,N_3504);
and U3629 (N_3629,N_3564,N_3577);
and U3630 (N_3630,N_3524,N_3509);
nand U3631 (N_3631,N_3590,N_3529);
nand U3632 (N_3632,N_3545,N_3544);
nand U3633 (N_3633,N_3594,N_3558);
and U3634 (N_3634,N_3598,N_3546);
nor U3635 (N_3635,N_3555,N_3596);
nand U3636 (N_3636,N_3575,N_3516);
and U3637 (N_3637,N_3599,N_3573);
nand U3638 (N_3638,N_3550,N_3514);
nor U3639 (N_3639,N_3517,N_3553);
and U3640 (N_3640,N_3512,N_3572);
nand U3641 (N_3641,N_3584,N_3568);
nand U3642 (N_3642,N_3579,N_3557);
or U3643 (N_3643,N_3595,N_3574);
nand U3644 (N_3644,N_3561,N_3526);
or U3645 (N_3645,N_3531,N_3588);
nand U3646 (N_3646,N_3506,N_3570);
and U3647 (N_3647,N_3556,N_3548);
and U3648 (N_3648,N_3533,N_3525);
or U3649 (N_3649,N_3503,N_3501);
nor U3650 (N_3650,N_3568,N_3530);
or U3651 (N_3651,N_3567,N_3558);
nor U3652 (N_3652,N_3508,N_3589);
and U3653 (N_3653,N_3586,N_3598);
xnor U3654 (N_3654,N_3513,N_3522);
nor U3655 (N_3655,N_3501,N_3533);
and U3656 (N_3656,N_3550,N_3528);
and U3657 (N_3657,N_3595,N_3539);
nand U3658 (N_3658,N_3511,N_3520);
nor U3659 (N_3659,N_3594,N_3515);
or U3660 (N_3660,N_3508,N_3552);
nor U3661 (N_3661,N_3501,N_3532);
nand U3662 (N_3662,N_3548,N_3570);
or U3663 (N_3663,N_3570,N_3510);
and U3664 (N_3664,N_3525,N_3572);
and U3665 (N_3665,N_3519,N_3508);
nand U3666 (N_3666,N_3555,N_3559);
nor U3667 (N_3667,N_3582,N_3521);
and U3668 (N_3668,N_3533,N_3564);
nor U3669 (N_3669,N_3522,N_3558);
nor U3670 (N_3670,N_3579,N_3526);
nand U3671 (N_3671,N_3539,N_3592);
or U3672 (N_3672,N_3540,N_3564);
nand U3673 (N_3673,N_3544,N_3540);
and U3674 (N_3674,N_3546,N_3555);
or U3675 (N_3675,N_3523,N_3585);
or U3676 (N_3676,N_3582,N_3509);
nor U3677 (N_3677,N_3562,N_3522);
and U3678 (N_3678,N_3583,N_3544);
or U3679 (N_3679,N_3557,N_3558);
and U3680 (N_3680,N_3506,N_3564);
nor U3681 (N_3681,N_3509,N_3598);
xnor U3682 (N_3682,N_3566,N_3529);
nor U3683 (N_3683,N_3539,N_3577);
nand U3684 (N_3684,N_3538,N_3553);
nand U3685 (N_3685,N_3504,N_3503);
or U3686 (N_3686,N_3565,N_3552);
nand U3687 (N_3687,N_3544,N_3585);
nor U3688 (N_3688,N_3533,N_3592);
and U3689 (N_3689,N_3580,N_3511);
nor U3690 (N_3690,N_3584,N_3509);
and U3691 (N_3691,N_3574,N_3509);
and U3692 (N_3692,N_3536,N_3577);
or U3693 (N_3693,N_3578,N_3504);
nor U3694 (N_3694,N_3553,N_3564);
and U3695 (N_3695,N_3511,N_3500);
nand U3696 (N_3696,N_3596,N_3549);
xnor U3697 (N_3697,N_3557,N_3519);
and U3698 (N_3698,N_3593,N_3528);
nor U3699 (N_3699,N_3529,N_3508);
nor U3700 (N_3700,N_3697,N_3679);
and U3701 (N_3701,N_3664,N_3628);
nor U3702 (N_3702,N_3638,N_3658);
nor U3703 (N_3703,N_3619,N_3692);
nand U3704 (N_3704,N_3680,N_3696);
nand U3705 (N_3705,N_3605,N_3698);
and U3706 (N_3706,N_3623,N_3603);
or U3707 (N_3707,N_3662,N_3661);
nand U3708 (N_3708,N_3685,N_3610);
nor U3709 (N_3709,N_3651,N_3601);
or U3710 (N_3710,N_3667,N_3650);
and U3711 (N_3711,N_3663,N_3612);
or U3712 (N_3712,N_3686,N_3644);
nor U3713 (N_3713,N_3694,N_3688);
nand U3714 (N_3714,N_3627,N_3608);
nor U3715 (N_3715,N_3616,N_3634);
or U3716 (N_3716,N_3671,N_3657);
nand U3717 (N_3717,N_3668,N_3656);
or U3718 (N_3718,N_3655,N_3672);
or U3719 (N_3719,N_3624,N_3665);
nor U3720 (N_3720,N_3646,N_3626);
nor U3721 (N_3721,N_3669,N_3617);
and U3722 (N_3722,N_3611,N_3607);
nand U3723 (N_3723,N_3648,N_3691);
or U3724 (N_3724,N_3604,N_3654);
nand U3725 (N_3725,N_3684,N_3677);
nor U3726 (N_3726,N_3600,N_3659);
nor U3727 (N_3727,N_3699,N_3670);
nand U3728 (N_3728,N_3687,N_3674);
nand U3729 (N_3729,N_3632,N_3666);
or U3730 (N_3730,N_3606,N_3682);
nor U3731 (N_3731,N_3639,N_3652);
and U3732 (N_3732,N_3614,N_3645);
or U3733 (N_3733,N_3622,N_3629);
nor U3734 (N_3734,N_3678,N_3637);
or U3735 (N_3735,N_3635,N_3636);
and U3736 (N_3736,N_3633,N_3631);
nor U3737 (N_3737,N_3683,N_3690);
or U3738 (N_3738,N_3630,N_3673);
and U3739 (N_3739,N_3609,N_3693);
or U3740 (N_3740,N_3675,N_3681);
or U3741 (N_3741,N_3641,N_3625);
and U3742 (N_3742,N_3647,N_3649);
or U3743 (N_3743,N_3695,N_3620);
nand U3744 (N_3744,N_3653,N_3618);
nor U3745 (N_3745,N_3640,N_3660);
nand U3746 (N_3746,N_3676,N_3642);
xnor U3747 (N_3747,N_3615,N_3621);
nand U3748 (N_3748,N_3689,N_3613);
and U3749 (N_3749,N_3643,N_3602);
or U3750 (N_3750,N_3609,N_3671);
and U3751 (N_3751,N_3671,N_3648);
nand U3752 (N_3752,N_3637,N_3688);
nor U3753 (N_3753,N_3627,N_3667);
nand U3754 (N_3754,N_3617,N_3645);
or U3755 (N_3755,N_3662,N_3693);
and U3756 (N_3756,N_3657,N_3692);
nor U3757 (N_3757,N_3621,N_3696);
nor U3758 (N_3758,N_3664,N_3668);
xor U3759 (N_3759,N_3643,N_3606);
nand U3760 (N_3760,N_3631,N_3612);
and U3761 (N_3761,N_3656,N_3676);
nor U3762 (N_3762,N_3616,N_3690);
nor U3763 (N_3763,N_3660,N_3639);
nor U3764 (N_3764,N_3696,N_3629);
and U3765 (N_3765,N_3622,N_3627);
or U3766 (N_3766,N_3637,N_3650);
nand U3767 (N_3767,N_3625,N_3685);
and U3768 (N_3768,N_3651,N_3665);
or U3769 (N_3769,N_3657,N_3662);
nor U3770 (N_3770,N_3637,N_3695);
nand U3771 (N_3771,N_3669,N_3611);
or U3772 (N_3772,N_3678,N_3652);
nor U3773 (N_3773,N_3699,N_3664);
or U3774 (N_3774,N_3653,N_3682);
or U3775 (N_3775,N_3682,N_3646);
or U3776 (N_3776,N_3603,N_3628);
nand U3777 (N_3777,N_3614,N_3662);
nand U3778 (N_3778,N_3639,N_3614);
and U3779 (N_3779,N_3600,N_3650);
and U3780 (N_3780,N_3663,N_3627);
and U3781 (N_3781,N_3686,N_3609);
nand U3782 (N_3782,N_3600,N_3610);
nand U3783 (N_3783,N_3649,N_3691);
nor U3784 (N_3784,N_3686,N_3643);
nand U3785 (N_3785,N_3681,N_3635);
or U3786 (N_3786,N_3688,N_3628);
nand U3787 (N_3787,N_3615,N_3622);
nor U3788 (N_3788,N_3696,N_3642);
nor U3789 (N_3789,N_3641,N_3685);
nor U3790 (N_3790,N_3618,N_3686);
xnor U3791 (N_3791,N_3646,N_3663);
or U3792 (N_3792,N_3604,N_3668);
and U3793 (N_3793,N_3629,N_3665);
xor U3794 (N_3794,N_3652,N_3671);
and U3795 (N_3795,N_3626,N_3670);
and U3796 (N_3796,N_3617,N_3607);
and U3797 (N_3797,N_3601,N_3613);
or U3798 (N_3798,N_3604,N_3657);
and U3799 (N_3799,N_3641,N_3679);
nor U3800 (N_3800,N_3775,N_3728);
nand U3801 (N_3801,N_3744,N_3750);
or U3802 (N_3802,N_3732,N_3769);
nand U3803 (N_3803,N_3793,N_3794);
nand U3804 (N_3804,N_3770,N_3799);
and U3805 (N_3805,N_3760,N_3797);
and U3806 (N_3806,N_3704,N_3772);
nor U3807 (N_3807,N_3778,N_3748);
or U3808 (N_3808,N_3713,N_3781);
and U3809 (N_3809,N_3700,N_3783);
nand U3810 (N_3810,N_3721,N_3717);
nor U3811 (N_3811,N_3738,N_3718);
and U3812 (N_3812,N_3712,N_3773);
nor U3813 (N_3813,N_3739,N_3791);
nor U3814 (N_3814,N_3707,N_3749);
nand U3815 (N_3815,N_3779,N_3761);
nand U3816 (N_3816,N_3703,N_3714);
or U3817 (N_3817,N_3771,N_3796);
nor U3818 (N_3818,N_3701,N_3731);
nand U3819 (N_3819,N_3795,N_3710);
and U3820 (N_3820,N_3752,N_3751);
nor U3821 (N_3821,N_3706,N_3719);
and U3822 (N_3822,N_3757,N_3780);
xnor U3823 (N_3823,N_3792,N_3722);
and U3824 (N_3824,N_3755,N_3708);
nor U3825 (N_3825,N_3776,N_3798);
nand U3826 (N_3826,N_3753,N_3730);
or U3827 (N_3827,N_3711,N_3787);
and U3828 (N_3828,N_3766,N_3754);
nand U3829 (N_3829,N_3782,N_3765);
nor U3830 (N_3830,N_3725,N_3777);
and U3831 (N_3831,N_3767,N_3734);
and U3832 (N_3832,N_3786,N_3743);
nor U3833 (N_3833,N_3762,N_3763);
nor U3834 (N_3834,N_3742,N_3733);
nor U3835 (N_3835,N_3745,N_3764);
and U3836 (N_3836,N_3747,N_3735);
nand U3837 (N_3837,N_3774,N_3759);
nand U3838 (N_3838,N_3720,N_3724);
and U3839 (N_3839,N_3768,N_3737);
or U3840 (N_3840,N_3740,N_3716);
nand U3841 (N_3841,N_3789,N_3723);
and U3842 (N_3842,N_3741,N_3736);
or U3843 (N_3843,N_3729,N_3788);
nand U3844 (N_3844,N_3746,N_3702);
or U3845 (N_3845,N_3727,N_3784);
or U3846 (N_3846,N_3756,N_3726);
or U3847 (N_3847,N_3785,N_3709);
or U3848 (N_3848,N_3705,N_3758);
nand U3849 (N_3849,N_3715,N_3790);
and U3850 (N_3850,N_3751,N_3735);
and U3851 (N_3851,N_3709,N_3746);
nor U3852 (N_3852,N_3740,N_3783);
nand U3853 (N_3853,N_3759,N_3748);
or U3854 (N_3854,N_3752,N_3724);
nand U3855 (N_3855,N_3716,N_3729);
and U3856 (N_3856,N_3755,N_3781);
nor U3857 (N_3857,N_3776,N_3712);
or U3858 (N_3858,N_3701,N_3703);
xnor U3859 (N_3859,N_3761,N_3775);
or U3860 (N_3860,N_3790,N_3716);
or U3861 (N_3861,N_3709,N_3702);
or U3862 (N_3862,N_3737,N_3790);
or U3863 (N_3863,N_3786,N_3740);
and U3864 (N_3864,N_3721,N_3748);
or U3865 (N_3865,N_3716,N_3760);
and U3866 (N_3866,N_3762,N_3775);
and U3867 (N_3867,N_3753,N_3727);
and U3868 (N_3868,N_3789,N_3781);
nand U3869 (N_3869,N_3755,N_3717);
or U3870 (N_3870,N_3760,N_3775);
or U3871 (N_3871,N_3716,N_3746);
or U3872 (N_3872,N_3738,N_3796);
nand U3873 (N_3873,N_3739,N_3757);
nor U3874 (N_3874,N_3742,N_3771);
nand U3875 (N_3875,N_3737,N_3777);
nand U3876 (N_3876,N_3701,N_3754);
or U3877 (N_3877,N_3702,N_3719);
or U3878 (N_3878,N_3760,N_3787);
nor U3879 (N_3879,N_3741,N_3743);
nor U3880 (N_3880,N_3751,N_3785);
or U3881 (N_3881,N_3726,N_3775);
nor U3882 (N_3882,N_3702,N_3700);
nand U3883 (N_3883,N_3717,N_3738);
nor U3884 (N_3884,N_3783,N_3725);
or U3885 (N_3885,N_3712,N_3746);
nor U3886 (N_3886,N_3773,N_3771);
and U3887 (N_3887,N_3704,N_3748);
or U3888 (N_3888,N_3735,N_3743);
and U3889 (N_3889,N_3715,N_3703);
and U3890 (N_3890,N_3756,N_3788);
and U3891 (N_3891,N_3759,N_3788);
nor U3892 (N_3892,N_3708,N_3741);
nand U3893 (N_3893,N_3749,N_3757);
nand U3894 (N_3894,N_3785,N_3756);
or U3895 (N_3895,N_3739,N_3783);
and U3896 (N_3896,N_3714,N_3753);
and U3897 (N_3897,N_3780,N_3754);
nor U3898 (N_3898,N_3744,N_3752);
nand U3899 (N_3899,N_3757,N_3711);
nand U3900 (N_3900,N_3851,N_3823);
nand U3901 (N_3901,N_3817,N_3891);
or U3902 (N_3902,N_3830,N_3858);
nor U3903 (N_3903,N_3874,N_3863);
nand U3904 (N_3904,N_3829,N_3846);
or U3905 (N_3905,N_3890,N_3880);
nand U3906 (N_3906,N_3803,N_3862);
and U3907 (N_3907,N_3839,N_3827);
and U3908 (N_3908,N_3853,N_3888);
and U3909 (N_3909,N_3868,N_3814);
nor U3910 (N_3910,N_3864,N_3835);
nor U3911 (N_3911,N_3898,N_3822);
nor U3912 (N_3912,N_3894,N_3807);
and U3913 (N_3913,N_3802,N_3804);
nand U3914 (N_3914,N_3887,N_3895);
or U3915 (N_3915,N_3806,N_3856);
or U3916 (N_3916,N_3881,N_3833);
nor U3917 (N_3917,N_3838,N_3870);
and U3918 (N_3918,N_3818,N_3840);
or U3919 (N_3919,N_3886,N_3843);
or U3920 (N_3920,N_3885,N_3801);
or U3921 (N_3921,N_3805,N_3869);
nor U3922 (N_3922,N_3867,N_3893);
and U3923 (N_3923,N_3811,N_3810);
and U3924 (N_3924,N_3837,N_3899);
nor U3925 (N_3925,N_3859,N_3879);
nor U3926 (N_3926,N_3866,N_3865);
or U3927 (N_3927,N_3821,N_3809);
and U3928 (N_3928,N_3820,N_3896);
nand U3929 (N_3929,N_3842,N_3808);
nor U3930 (N_3930,N_3860,N_3884);
nor U3931 (N_3931,N_3834,N_3883);
and U3932 (N_3932,N_3882,N_3850);
nor U3933 (N_3933,N_3889,N_3848);
or U3934 (N_3934,N_3812,N_3819);
nor U3935 (N_3935,N_3826,N_3845);
nor U3936 (N_3936,N_3849,N_3831);
or U3937 (N_3937,N_3825,N_3857);
or U3938 (N_3938,N_3875,N_3878);
or U3939 (N_3939,N_3828,N_3844);
nand U3940 (N_3940,N_3861,N_3892);
or U3941 (N_3941,N_3813,N_3872);
or U3942 (N_3942,N_3871,N_3877);
or U3943 (N_3943,N_3876,N_3873);
or U3944 (N_3944,N_3854,N_3852);
nand U3945 (N_3945,N_3841,N_3824);
nand U3946 (N_3946,N_3816,N_3897);
nor U3947 (N_3947,N_3847,N_3800);
and U3948 (N_3948,N_3815,N_3836);
nand U3949 (N_3949,N_3855,N_3832);
and U3950 (N_3950,N_3890,N_3813);
and U3951 (N_3951,N_3814,N_3845);
or U3952 (N_3952,N_3830,N_3827);
nor U3953 (N_3953,N_3824,N_3802);
nor U3954 (N_3954,N_3807,N_3822);
xnor U3955 (N_3955,N_3883,N_3802);
nand U3956 (N_3956,N_3895,N_3885);
or U3957 (N_3957,N_3801,N_3841);
nand U3958 (N_3958,N_3801,N_3837);
nor U3959 (N_3959,N_3807,N_3808);
or U3960 (N_3960,N_3892,N_3839);
nand U3961 (N_3961,N_3818,N_3859);
xor U3962 (N_3962,N_3814,N_3818);
nor U3963 (N_3963,N_3846,N_3881);
nor U3964 (N_3964,N_3825,N_3886);
nand U3965 (N_3965,N_3861,N_3877);
nand U3966 (N_3966,N_3841,N_3821);
and U3967 (N_3967,N_3821,N_3836);
nand U3968 (N_3968,N_3832,N_3815);
nor U3969 (N_3969,N_3874,N_3814);
and U3970 (N_3970,N_3898,N_3812);
and U3971 (N_3971,N_3849,N_3860);
nand U3972 (N_3972,N_3837,N_3890);
and U3973 (N_3973,N_3836,N_3881);
nor U3974 (N_3974,N_3846,N_3831);
nand U3975 (N_3975,N_3831,N_3806);
nand U3976 (N_3976,N_3849,N_3846);
or U3977 (N_3977,N_3860,N_3807);
and U3978 (N_3978,N_3839,N_3882);
nand U3979 (N_3979,N_3844,N_3803);
nand U3980 (N_3980,N_3889,N_3859);
nand U3981 (N_3981,N_3895,N_3804);
or U3982 (N_3982,N_3855,N_3862);
or U3983 (N_3983,N_3866,N_3804);
nor U3984 (N_3984,N_3833,N_3822);
or U3985 (N_3985,N_3847,N_3879);
or U3986 (N_3986,N_3897,N_3826);
nor U3987 (N_3987,N_3860,N_3879);
nor U3988 (N_3988,N_3812,N_3860);
or U3989 (N_3989,N_3875,N_3845);
nor U3990 (N_3990,N_3892,N_3865);
nand U3991 (N_3991,N_3828,N_3887);
nor U3992 (N_3992,N_3879,N_3856);
or U3993 (N_3993,N_3804,N_3853);
and U3994 (N_3994,N_3819,N_3856);
or U3995 (N_3995,N_3851,N_3839);
nand U3996 (N_3996,N_3878,N_3823);
and U3997 (N_3997,N_3866,N_3883);
nor U3998 (N_3998,N_3861,N_3899);
nand U3999 (N_3999,N_3842,N_3817);
or U4000 (N_4000,N_3959,N_3936);
and U4001 (N_4001,N_3915,N_3914);
and U4002 (N_4002,N_3962,N_3932);
or U4003 (N_4003,N_3949,N_3908);
or U4004 (N_4004,N_3933,N_3987);
xor U4005 (N_4005,N_3989,N_3931);
nor U4006 (N_4006,N_3907,N_3990);
or U4007 (N_4007,N_3921,N_3997);
nor U4008 (N_4008,N_3970,N_3951);
nand U4009 (N_4009,N_3946,N_3977);
nor U4010 (N_4010,N_3945,N_3918);
or U4011 (N_4011,N_3961,N_3909);
or U4012 (N_4012,N_3967,N_3944);
and U4013 (N_4013,N_3937,N_3963);
xnor U4014 (N_4014,N_3928,N_3976);
and U4015 (N_4015,N_3979,N_3982);
nor U4016 (N_4016,N_3953,N_3998);
nand U4017 (N_4017,N_3988,N_3983);
or U4018 (N_4018,N_3994,N_3923);
nand U4019 (N_4019,N_3948,N_3972);
nand U4020 (N_4020,N_3916,N_3995);
or U4021 (N_4021,N_3968,N_3929);
nand U4022 (N_4022,N_3917,N_3971);
and U4023 (N_4023,N_3939,N_3956);
nor U4024 (N_4024,N_3950,N_3985);
nor U4025 (N_4025,N_3902,N_3930);
and U4026 (N_4026,N_3980,N_3952);
xor U4027 (N_4027,N_3981,N_3974);
and U4028 (N_4028,N_3958,N_3960);
or U4029 (N_4029,N_3911,N_3991);
nand U4030 (N_4030,N_3966,N_3969);
or U4031 (N_4031,N_3913,N_3954);
and U4032 (N_4032,N_3938,N_3965);
or U4033 (N_4033,N_3935,N_3942);
nor U4034 (N_4034,N_3925,N_3978);
nor U4035 (N_4035,N_3943,N_3940);
nand U4036 (N_4036,N_3919,N_3900);
or U4037 (N_4037,N_3986,N_3912);
nor U4038 (N_4038,N_3964,N_3905);
xnor U4039 (N_4039,N_3955,N_3999);
and U4040 (N_4040,N_3957,N_3993);
or U4041 (N_4041,N_3904,N_3926);
xor U4042 (N_4042,N_3973,N_3920);
nor U4043 (N_4043,N_3922,N_3927);
and U4044 (N_4044,N_3947,N_3975);
nor U4045 (N_4045,N_3941,N_3901);
nor U4046 (N_4046,N_3924,N_3906);
and U4047 (N_4047,N_3903,N_3996);
and U4048 (N_4048,N_3992,N_3934);
and U4049 (N_4049,N_3984,N_3910);
nor U4050 (N_4050,N_3901,N_3962);
and U4051 (N_4051,N_3946,N_3918);
or U4052 (N_4052,N_3980,N_3987);
nor U4053 (N_4053,N_3935,N_3953);
and U4054 (N_4054,N_3989,N_3968);
and U4055 (N_4055,N_3977,N_3931);
and U4056 (N_4056,N_3956,N_3988);
or U4057 (N_4057,N_3954,N_3972);
or U4058 (N_4058,N_3969,N_3972);
and U4059 (N_4059,N_3957,N_3935);
nand U4060 (N_4060,N_3931,N_3961);
or U4061 (N_4061,N_3981,N_3906);
and U4062 (N_4062,N_3934,N_3914);
nor U4063 (N_4063,N_3922,N_3921);
or U4064 (N_4064,N_3979,N_3912);
or U4065 (N_4065,N_3926,N_3912);
and U4066 (N_4066,N_3919,N_3968);
and U4067 (N_4067,N_3950,N_3983);
and U4068 (N_4068,N_3947,N_3955);
nand U4069 (N_4069,N_3975,N_3990);
nand U4070 (N_4070,N_3976,N_3953);
and U4071 (N_4071,N_3988,N_3969);
and U4072 (N_4072,N_3996,N_3973);
and U4073 (N_4073,N_3945,N_3906);
or U4074 (N_4074,N_3935,N_3903);
nand U4075 (N_4075,N_3991,N_3929);
xnor U4076 (N_4076,N_3955,N_3941);
and U4077 (N_4077,N_3930,N_3919);
nand U4078 (N_4078,N_3907,N_3936);
and U4079 (N_4079,N_3952,N_3927);
or U4080 (N_4080,N_3941,N_3940);
nor U4081 (N_4081,N_3930,N_3964);
nor U4082 (N_4082,N_3974,N_3920);
or U4083 (N_4083,N_3969,N_3932);
xor U4084 (N_4084,N_3977,N_3970);
nor U4085 (N_4085,N_3990,N_3965);
and U4086 (N_4086,N_3960,N_3993);
and U4087 (N_4087,N_3963,N_3968);
or U4088 (N_4088,N_3973,N_3988);
and U4089 (N_4089,N_3919,N_3978);
nand U4090 (N_4090,N_3959,N_3981);
and U4091 (N_4091,N_3943,N_3951);
and U4092 (N_4092,N_3970,N_3953);
or U4093 (N_4093,N_3998,N_3978);
and U4094 (N_4094,N_3929,N_3939);
nand U4095 (N_4095,N_3996,N_3994);
or U4096 (N_4096,N_3955,N_3932);
nand U4097 (N_4097,N_3916,N_3934);
or U4098 (N_4098,N_3953,N_3979);
or U4099 (N_4099,N_3988,N_3972);
or U4100 (N_4100,N_4043,N_4081);
nor U4101 (N_4101,N_4056,N_4087);
or U4102 (N_4102,N_4055,N_4060);
and U4103 (N_4103,N_4012,N_4062);
and U4104 (N_4104,N_4007,N_4044);
nand U4105 (N_4105,N_4000,N_4021);
or U4106 (N_4106,N_4077,N_4039);
nand U4107 (N_4107,N_4067,N_4093);
nand U4108 (N_4108,N_4031,N_4019);
and U4109 (N_4109,N_4038,N_4002);
nor U4110 (N_4110,N_4070,N_4063);
nor U4111 (N_4111,N_4091,N_4008);
and U4112 (N_4112,N_4088,N_4090);
or U4113 (N_4113,N_4041,N_4075);
and U4114 (N_4114,N_4053,N_4082);
xnor U4115 (N_4115,N_4004,N_4071);
and U4116 (N_4116,N_4006,N_4058);
and U4117 (N_4117,N_4035,N_4092);
nor U4118 (N_4118,N_4042,N_4020);
nor U4119 (N_4119,N_4078,N_4037);
nand U4120 (N_4120,N_4069,N_4011);
or U4121 (N_4121,N_4034,N_4098);
nor U4122 (N_4122,N_4032,N_4083);
and U4123 (N_4123,N_4080,N_4089);
or U4124 (N_4124,N_4076,N_4029);
or U4125 (N_4125,N_4049,N_4096);
nor U4126 (N_4126,N_4025,N_4016);
nor U4127 (N_4127,N_4033,N_4066);
and U4128 (N_4128,N_4001,N_4024);
xor U4129 (N_4129,N_4027,N_4086);
or U4130 (N_4130,N_4072,N_4095);
nand U4131 (N_4131,N_4040,N_4005);
or U4132 (N_4132,N_4017,N_4085);
xnor U4133 (N_4133,N_4048,N_4057);
and U4134 (N_4134,N_4074,N_4052);
xor U4135 (N_4135,N_4015,N_4022);
and U4136 (N_4136,N_4073,N_4028);
and U4137 (N_4137,N_4051,N_4061);
nor U4138 (N_4138,N_4030,N_4065);
nand U4139 (N_4139,N_4013,N_4059);
or U4140 (N_4140,N_4054,N_4068);
xor U4141 (N_4141,N_4099,N_4010);
or U4142 (N_4142,N_4014,N_4023);
and U4143 (N_4143,N_4026,N_4047);
nor U4144 (N_4144,N_4050,N_4097);
and U4145 (N_4145,N_4003,N_4045);
or U4146 (N_4146,N_4036,N_4009);
nor U4147 (N_4147,N_4084,N_4094);
or U4148 (N_4148,N_4064,N_4018);
nand U4149 (N_4149,N_4079,N_4046);
xor U4150 (N_4150,N_4048,N_4040);
and U4151 (N_4151,N_4095,N_4038);
nor U4152 (N_4152,N_4098,N_4057);
nand U4153 (N_4153,N_4096,N_4025);
nand U4154 (N_4154,N_4071,N_4085);
and U4155 (N_4155,N_4080,N_4045);
and U4156 (N_4156,N_4076,N_4008);
or U4157 (N_4157,N_4084,N_4005);
or U4158 (N_4158,N_4009,N_4058);
and U4159 (N_4159,N_4039,N_4014);
or U4160 (N_4160,N_4064,N_4095);
or U4161 (N_4161,N_4023,N_4042);
or U4162 (N_4162,N_4000,N_4018);
nor U4163 (N_4163,N_4013,N_4071);
or U4164 (N_4164,N_4026,N_4081);
nand U4165 (N_4165,N_4085,N_4050);
nand U4166 (N_4166,N_4049,N_4047);
nand U4167 (N_4167,N_4070,N_4000);
nand U4168 (N_4168,N_4086,N_4065);
and U4169 (N_4169,N_4026,N_4038);
nand U4170 (N_4170,N_4065,N_4035);
nor U4171 (N_4171,N_4059,N_4046);
or U4172 (N_4172,N_4070,N_4054);
and U4173 (N_4173,N_4033,N_4070);
and U4174 (N_4174,N_4045,N_4004);
or U4175 (N_4175,N_4082,N_4039);
nand U4176 (N_4176,N_4013,N_4023);
and U4177 (N_4177,N_4063,N_4031);
nand U4178 (N_4178,N_4006,N_4096);
nor U4179 (N_4179,N_4047,N_4034);
and U4180 (N_4180,N_4073,N_4044);
nor U4181 (N_4181,N_4045,N_4085);
or U4182 (N_4182,N_4020,N_4083);
or U4183 (N_4183,N_4003,N_4079);
and U4184 (N_4184,N_4069,N_4010);
and U4185 (N_4185,N_4029,N_4023);
nor U4186 (N_4186,N_4083,N_4070);
nand U4187 (N_4187,N_4048,N_4077);
nor U4188 (N_4188,N_4052,N_4091);
or U4189 (N_4189,N_4087,N_4086);
nand U4190 (N_4190,N_4099,N_4008);
nor U4191 (N_4191,N_4018,N_4080);
and U4192 (N_4192,N_4028,N_4015);
or U4193 (N_4193,N_4086,N_4069);
and U4194 (N_4194,N_4064,N_4092);
and U4195 (N_4195,N_4044,N_4059);
nand U4196 (N_4196,N_4074,N_4045);
or U4197 (N_4197,N_4095,N_4017);
and U4198 (N_4198,N_4062,N_4049);
nor U4199 (N_4199,N_4068,N_4060);
nand U4200 (N_4200,N_4135,N_4183);
and U4201 (N_4201,N_4174,N_4182);
or U4202 (N_4202,N_4197,N_4125);
or U4203 (N_4203,N_4185,N_4104);
and U4204 (N_4204,N_4143,N_4168);
nand U4205 (N_4205,N_4198,N_4184);
or U4206 (N_4206,N_4131,N_4130);
nand U4207 (N_4207,N_4188,N_4172);
or U4208 (N_4208,N_4190,N_4186);
and U4209 (N_4209,N_4140,N_4121);
nor U4210 (N_4210,N_4189,N_4133);
nor U4211 (N_4211,N_4180,N_4160);
and U4212 (N_4212,N_4128,N_4167);
nand U4213 (N_4213,N_4196,N_4175);
and U4214 (N_4214,N_4100,N_4195);
xnor U4215 (N_4215,N_4142,N_4187);
nand U4216 (N_4216,N_4129,N_4113);
nand U4217 (N_4217,N_4155,N_4132);
or U4218 (N_4218,N_4134,N_4116);
and U4219 (N_4219,N_4136,N_4153);
and U4220 (N_4220,N_4192,N_4106);
or U4221 (N_4221,N_4165,N_4146);
and U4222 (N_4222,N_4157,N_4191);
and U4223 (N_4223,N_4179,N_4193);
nor U4224 (N_4224,N_4139,N_4117);
nand U4225 (N_4225,N_4166,N_4199);
and U4226 (N_4226,N_4101,N_4111);
nor U4227 (N_4227,N_4127,N_4105);
xor U4228 (N_4228,N_4162,N_4178);
and U4229 (N_4229,N_4158,N_4163);
and U4230 (N_4230,N_4177,N_4123);
and U4231 (N_4231,N_4181,N_4119);
and U4232 (N_4232,N_4102,N_4108);
or U4233 (N_4233,N_4103,N_4194);
nand U4234 (N_4234,N_4114,N_4161);
nand U4235 (N_4235,N_4152,N_4122);
or U4236 (N_4236,N_4159,N_4124);
or U4237 (N_4237,N_4109,N_4147);
nand U4238 (N_4238,N_4126,N_4173);
and U4239 (N_4239,N_4171,N_4138);
or U4240 (N_4240,N_4170,N_4151);
or U4241 (N_4241,N_4120,N_4107);
nand U4242 (N_4242,N_4141,N_4144);
or U4243 (N_4243,N_4110,N_4115);
nand U4244 (N_4244,N_4156,N_4112);
nor U4245 (N_4245,N_4148,N_4176);
or U4246 (N_4246,N_4150,N_4137);
nand U4247 (N_4247,N_4118,N_4169);
nand U4248 (N_4248,N_4145,N_4149);
or U4249 (N_4249,N_4164,N_4154);
and U4250 (N_4250,N_4191,N_4169);
and U4251 (N_4251,N_4178,N_4119);
nor U4252 (N_4252,N_4130,N_4148);
or U4253 (N_4253,N_4189,N_4107);
and U4254 (N_4254,N_4192,N_4131);
or U4255 (N_4255,N_4187,N_4126);
and U4256 (N_4256,N_4126,N_4123);
nand U4257 (N_4257,N_4187,N_4198);
nand U4258 (N_4258,N_4166,N_4171);
nor U4259 (N_4259,N_4106,N_4190);
nand U4260 (N_4260,N_4142,N_4158);
nor U4261 (N_4261,N_4183,N_4103);
nand U4262 (N_4262,N_4184,N_4143);
nor U4263 (N_4263,N_4150,N_4103);
and U4264 (N_4264,N_4138,N_4157);
nor U4265 (N_4265,N_4108,N_4195);
or U4266 (N_4266,N_4126,N_4110);
and U4267 (N_4267,N_4162,N_4128);
nor U4268 (N_4268,N_4156,N_4182);
and U4269 (N_4269,N_4165,N_4160);
nand U4270 (N_4270,N_4104,N_4101);
nand U4271 (N_4271,N_4111,N_4143);
nand U4272 (N_4272,N_4167,N_4159);
and U4273 (N_4273,N_4109,N_4170);
or U4274 (N_4274,N_4146,N_4115);
or U4275 (N_4275,N_4119,N_4198);
or U4276 (N_4276,N_4122,N_4140);
xnor U4277 (N_4277,N_4148,N_4163);
and U4278 (N_4278,N_4195,N_4170);
nand U4279 (N_4279,N_4197,N_4195);
and U4280 (N_4280,N_4178,N_4128);
nand U4281 (N_4281,N_4106,N_4168);
or U4282 (N_4282,N_4122,N_4182);
nand U4283 (N_4283,N_4112,N_4122);
nand U4284 (N_4284,N_4138,N_4174);
or U4285 (N_4285,N_4122,N_4169);
nand U4286 (N_4286,N_4126,N_4128);
nor U4287 (N_4287,N_4122,N_4165);
and U4288 (N_4288,N_4172,N_4136);
and U4289 (N_4289,N_4170,N_4185);
and U4290 (N_4290,N_4139,N_4127);
nor U4291 (N_4291,N_4107,N_4182);
or U4292 (N_4292,N_4106,N_4133);
and U4293 (N_4293,N_4143,N_4120);
nor U4294 (N_4294,N_4113,N_4100);
or U4295 (N_4295,N_4122,N_4119);
nand U4296 (N_4296,N_4198,N_4131);
or U4297 (N_4297,N_4102,N_4139);
and U4298 (N_4298,N_4118,N_4189);
nand U4299 (N_4299,N_4195,N_4112);
or U4300 (N_4300,N_4279,N_4203);
nor U4301 (N_4301,N_4291,N_4285);
and U4302 (N_4302,N_4264,N_4266);
xor U4303 (N_4303,N_4241,N_4276);
or U4304 (N_4304,N_4207,N_4222);
nand U4305 (N_4305,N_4284,N_4280);
nor U4306 (N_4306,N_4243,N_4258);
and U4307 (N_4307,N_4263,N_4296);
nand U4308 (N_4308,N_4287,N_4227);
and U4309 (N_4309,N_4240,N_4267);
and U4310 (N_4310,N_4239,N_4261);
and U4311 (N_4311,N_4225,N_4244);
nand U4312 (N_4312,N_4255,N_4271);
nor U4313 (N_4313,N_4208,N_4228);
nand U4314 (N_4314,N_4262,N_4235);
or U4315 (N_4315,N_4217,N_4253);
xor U4316 (N_4316,N_4234,N_4297);
nor U4317 (N_4317,N_4272,N_4277);
nor U4318 (N_4318,N_4251,N_4299);
or U4319 (N_4319,N_4212,N_4286);
and U4320 (N_4320,N_4221,N_4250);
nand U4321 (N_4321,N_4273,N_4238);
or U4322 (N_4322,N_4206,N_4282);
nor U4323 (N_4323,N_4205,N_4211);
and U4324 (N_4324,N_4278,N_4213);
nand U4325 (N_4325,N_4254,N_4233);
nand U4326 (N_4326,N_4204,N_4293);
xnor U4327 (N_4327,N_4281,N_4220);
nor U4328 (N_4328,N_4265,N_4236);
nor U4329 (N_4329,N_4200,N_4256);
nor U4330 (N_4330,N_4298,N_4230);
and U4331 (N_4331,N_4210,N_4215);
nand U4332 (N_4332,N_4229,N_4214);
and U4333 (N_4333,N_4275,N_4226);
and U4334 (N_4334,N_4223,N_4219);
nand U4335 (N_4335,N_4290,N_4202);
nand U4336 (N_4336,N_4295,N_4231);
or U4337 (N_4337,N_4283,N_4209);
or U4338 (N_4338,N_4237,N_4292);
xor U4339 (N_4339,N_4245,N_4216);
nand U4340 (N_4340,N_4288,N_4232);
or U4341 (N_4341,N_4257,N_4248);
nor U4342 (N_4342,N_4224,N_4246);
or U4343 (N_4343,N_4201,N_4249);
or U4344 (N_4344,N_4268,N_4269);
or U4345 (N_4345,N_4247,N_4252);
nand U4346 (N_4346,N_4259,N_4289);
and U4347 (N_4347,N_4242,N_4274);
or U4348 (N_4348,N_4218,N_4260);
nor U4349 (N_4349,N_4294,N_4270);
or U4350 (N_4350,N_4270,N_4203);
and U4351 (N_4351,N_4278,N_4252);
xor U4352 (N_4352,N_4247,N_4283);
and U4353 (N_4353,N_4236,N_4205);
nor U4354 (N_4354,N_4238,N_4284);
nor U4355 (N_4355,N_4276,N_4250);
nand U4356 (N_4356,N_4283,N_4255);
or U4357 (N_4357,N_4285,N_4258);
or U4358 (N_4358,N_4216,N_4275);
or U4359 (N_4359,N_4265,N_4254);
and U4360 (N_4360,N_4202,N_4283);
nor U4361 (N_4361,N_4257,N_4252);
nand U4362 (N_4362,N_4285,N_4208);
or U4363 (N_4363,N_4221,N_4202);
nor U4364 (N_4364,N_4247,N_4265);
and U4365 (N_4365,N_4223,N_4251);
and U4366 (N_4366,N_4247,N_4235);
or U4367 (N_4367,N_4265,N_4223);
xnor U4368 (N_4368,N_4275,N_4237);
or U4369 (N_4369,N_4245,N_4200);
and U4370 (N_4370,N_4243,N_4290);
or U4371 (N_4371,N_4258,N_4219);
or U4372 (N_4372,N_4271,N_4208);
or U4373 (N_4373,N_4275,N_4262);
nand U4374 (N_4374,N_4209,N_4259);
nor U4375 (N_4375,N_4215,N_4250);
and U4376 (N_4376,N_4226,N_4228);
nand U4377 (N_4377,N_4288,N_4257);
or U4378 (N_4378,N_4203,N_4233);
nor U4379 (N_4379,N_4293,N_4236);
xnor U4380 (N_4380,N_4271,N_4235);
nor U4381 (N_4381,N_4244,N_4284);
and U4382 (N_4382,N_4260,N_4298);
or U4383 (N_4383,N_4210,N_4289);
xnor U4384 (N_4384,N_4203,N_4255);
nor U4385 (N_4385,N_4211,N_4224);
or U4386 (N_4386,N_4211,N_4287);
xnor U4387 (N_4387,N_4291,N_4225);
xnor U4388 (N_4388,N_4260,N_4263);
nor U4389 (N_4389,N_4204,N_4225);
and U4390 (N_4390,N_4267,N_4218);
and U4391 (N_4391,N_4247,N_4289);
nor U4392 (N_4392,N_4220,N_4230);
nor U4393 (N_4393,N_4242,N_4243);
and U4394 (N_4394,N_4211,N_4264);
or U4395 (N_4395,N_4258,N_4274);
nor U4396 (N_4396,N_4257,N_4256);
nor U4397 (N_4397,N_4209,N_4268);
and U4398 (N_4398,N_4256,N_4208);
xnor U4399 (N_4399,N_4297,N_4204);
nand U4400 (N_4400,N_4391,N_4369);
and U4401 (N_4401,N_4322,N_4388);
nor U4402 (N_4402,N_4397,N_4337);
nand U4403 (N_4403,N_4310,N_4350);
and U4404 (N_4404,N_4329,N_4316);
nor U4405 (N_4405,N_4303,N_4398);
or U4406 (N_4406,N_4300,N_4336);
nand U4407 (N_4407,N_4338,N_4343);
nand U4408 (N_4408,N_4395,N_4304);
nand U4409 (N_4409,N_4357,N_4371);
nand U4410 (N_4410,N_4354,N_4335);
and U4411 (N_4411,N_4373,N_4379);
and U4412 (N_4412,N_4325,N_4380);
and U4413 (N_4413,N_4306,N_4334);
and U4414 (N_4414,N_4314,N_4364);
and U4415 (N_4415,N_4309,N_4392);
xnor U4416 (N_4416,N_4356,N_4313);
and U4417 (N_4417,N_4341,N_4361);
or U4418 (N_4418,N_4358,N_4345);
or U4419 (N_4419,N_4349,N_4312);
and U4420 (N_4420,N_4365,N_4321);
nor U4421 (N_4421,N_4377,N_4319);
and U4422 (N_4422,N_4372,N_4347);
nand U4423 (N_4423,N_4307,N_4352);
and U4424 (N_4424,N_4340,N_4390);
nand U4425 (N_4425,N_4318,N_4393);
or U4426 (N_4426,N_4368,N_4315);
nor U4427 (N_4427,N_4359,N_4374);
or U4428 (N_4428,N_4311,N_4389);
and U4429 (N_4429,N_4387,N_4330);
and U4430 (N_4430,N_4383,N_4396);
nand U4431 (N_4431,N_4376,N_4360);
or U4432 (N_4432,N_4399,N_4332);
or U4433 (N_4433,N_4339,N_4326);
or U4434 (N_4434,N_4301,N_4344);
nand U4435 (N_4435,N_4348,N_4385);
nor U4436 (N_4436,N_4302,N_4317);
nor U4437 (N_4437,N_4320,N_4308);
nand U4438 (N_4438,N_4346,N_4381);
or U4439 (N_4439,N_4386,N_4362);
nor U4440 (N_4440,N_4355,N_4384);
nor U4441 (N_4441,N_4323,N_4324);
nand U4442 (N_4442,N_4363,N_4305);
nor U4443 (N_4443,N_4351,N_4333);
or U4444 (N_4444,N_4353,N_4375);
and U4445 (N_4445,N_4327,N_4382);
nand U4446 (N_4446,N_4342,N_4394);
nand U4447 (N_4447,N_4328,N_4331);
nand U4448 (N_4448,N_4366,N_4370);
nor U4449 (N_4449,N_4367,N_4378);
nand U4450 (N_4450,N_4393,N_4353);
nor U4451 (N_4451,N_4317,N_4359);
nand U4452 (N_4452,N_4321,N_4346);
and U4453 (N_4453,N_4312,N_4329);
or U4454 (N_4454,N_4327,N_4362);
and U4455 (N_4455,N_4358,N_4361);
and U4456 (N_4456,N_4333,N_4352);
or U4457 (N_4457,N_4396,N_4308);
nor U4458 (N_4458,N_4307,N_4396);
and U4459 (N_4459,N_4321,N_4392);
nand U4460 (N_4460,N_4354,N_4370);
nor U4461 (N_4461,N_4363,N_4322);
nand U4462 (N_4462,N_4397,N_4323);
nor U4463 (N_4463,N_4348,N_4365);
and U4464 (N_4464,N_4317,N_4385);
or U4465 (N_4465,N_4396,N_4325);
nand U4466 (N_4466,N_4305,N_4354);
nor U4467 (N_4467,N_4388,N_4319);
or U4468 (N_4468,N_4340,N_4333);
nor U4469 (N_4469,N_4302,N_4307);
or U4470 (N_4470,N_4388,N_4339);
or U4471 (N_4471,N_4380,N_4305);
nor U4472 (N_4472,N_4354,N_4394);
or U4473 (N_4473,N_4330,N_4331);
and U4474 (N_4474,N_4399,N_4300);
nor U4475 (N_4475,N_4366,N_4330);
nor U4476 (N_4476,N_4384,N_4372);
nor U4477 (N_4477,N_4323,N_4361);
or U4478 (N_4478,N_4388,N_4329);
or U4479 (N_4479,N_4384,N_4382);
or U4480 (N_4480,N_4373,N_4348);
and U4481 (N_4481,N_4352,N_4335);
and U4482 (N_4482,N_4312,N_4371);
and U4483 (N_4483,N_4341,N_4332);
and U4484 (N_4484,N_4352,N_4327);
nor U4485 (N_4485,N_4368,N_4387);
nand U4486 (N_4486,N_4362,N_4329);
nand U4487 (N_4487,N_4334,N_4339);
nor U4488 (N_4488,N_4300,N_4317);
or U4489 (N_4489,N_4310,N_4319);
nor U4490 (N_4490,N_4317,N_4378);
nor U4491 (N_4491,N_4309,N_4380);
or U4492 (N_4492,N_4323,N_4339);
nand U4493 (N_4493,N_4329,N_4347);
or U4494 (N_4494,N_4343,N_4360);
nor U4495 (N_4495,N_4392,N_4343);
nor U4496 (N_4496,N_4312,N_4305);
or U4497 (N_4497,N_4301,N_4319);
xnor U4498 (N_4498,N_4328,N_4361);
nand U4499 (N_4499,N_4352,N_4377);
or U4500 (N_4500,N_4471,N_4438);
nand U4501 (N_4501,N_4470,N_4402);
nor U4502 (N_4502,N_4497,N_4465);
or U4503 (N_4503,N_4466,N_4439);
and U4504 (N_4504,N_4425,N_4432);
or U4505 (N_4505,N_4445,N_4426);
or U4506 (N_4506,N_4490,N_4441);
nor U4507 (N_4507,N_4417,N_4488);
and U4508 (N_4508,N_4420,N_4481);
nand U4509 (N_4509,N_4403,N_4416);
nor U4510 (N_4510,N_4472,N_4469);
or U4511 (N_4511,N_4468,N_4491);
nand U4512 (N_4512,N_4463,N_4429);
and U4513 (N_4513,N_4419,N_4460);
or U4514 (N_4514,N_4428,N_4440);
nand U4515 (N_4515,N_4480,N_4482);
nor U4516 (N_4516,N_4452,N_4450);
or U4517 (N_4517,N_4489,N_4431);
or U4518 (N_4518,N_4492,N_4442);
or U4519 (N_4519,N_4476,N_4479);
or U4520 (N_4520,N_4404,N_4436);
nand U4521 (N_4521,N_4462,N_4493);
and U4522 (N_4522,N_4412,N_4443);
or U4523 (N_4523,N_4449,N_4422);
or U4524 (N_4524,N_4483,N_4401);
nand U4525 (N_4525,N_4499,N_4487);
or U4526 (N_4526,N_4459,N_4477);
and U4527 (N_4527,N_4451,N_4434);
nor U4528 (N_4528,N_4427,N_4409);
and U4529 (N_4529,N_4411,N_4444);
nor U4530 (N_4530,N_4474,N_4400);
or U4531 (N_4531,N_4475,N_4458);
nor U4532 (N_4532,N_4486,N_4455);
and U4533 (N_4533,N_4430,N_4495);
nand U4534 (N_4534,N_4435,N_4405);
nand U4535 (N_4535,N_4485,N_4484);
xnor U4536 (N_4536,N_4457,N_4446);
nand U4537 (N_4537,N_4496,N_4467);
nand U4538 (N_4538,N_4454,N_4494);
nand U4539 (N_4539,N_4473,N_4478);
xor U4540 (N_4540,N_4456,N_4423);
nor U4541 (N_4541,N_4437,N_4447);
or U4542 (N_4542,N_4453,N_4406);
nor U4543 (N_4543,N_4421,N_4408);
and U4544 (N_4544,N_4418,N_4464);
nand U4545 (N_4545,N_4461,N_4413);
and U4546 (N_4546,N_4415,N_4407);
or U4547 (N_4547,N_4414,N_4448);
nand U4548 (N_4548,N_4433,N_4410);
nor U4549 (N_4549,N_4498,N_4424);
nor U4550 (N_4550,N_4442,N_4441);
and U4551 (N_4551,N_4421,N_4440);
and U4552 (N_4552,N_4433,N_4425);
nor U4553 (N_4553,N_4459,N_4469);
or U4554 (N_4554,N_4489,N_4400);
nand U4555 (N_4555,N_4452,N_4457);
nand U4556 (N_4556,N_4440,N_4490);
nor U4557 (N_4557,N_4425,N_4479);
or U4558 (N_4558,N_4405,N_4454);
and U4559 (N_4559,N_4463,N_4405);
nor U4560 (N_4560,N_4459,N_4497);
nor U4561 (N_4561,N_4421,N_4468);
or U4562 (N_4562,N_4463,N_4487);
or U4563 (N_4563,N_4494,N_4418);
and U4564 (N_4564,N_4436,N_4426);
nor U4565 (N_4565,N_4415,N_4421);
or U4566 (N_4566,N_4480,N_4416);
nand U4567 (N_4567,N_4494,N_4440);
and U4568 (N_4568,N_4460,N_4482);
nor U4569 (N_4569,N_4477,N_4423);
nand U4570 (N_4570,N_4401,N_4482);
and U4571 (N_4571,N_4426,N_4486);
or U4572 (N_4572,N_4463,N_4418);
nand U4573 (N_4573,N_4424,N_4443);
nand U4574 (N_4574,N_4472,N_4414);
and U4575 (N_4575,N_4456,N_4475);
or U4576 (N_4576,N_4496,N_4437);
nand U4577 (N_4577,N_4443,N_4441);
nand U4578 (N_4578,N_4427,N_4403);
nand U4579 (N_4579,N_4423,N_4470);
nor U4580 (N_4580,N_4437,N_4416);
and U4581 (N_4581,N_4437,N_4450);
nor U4582 (N_4582,N_4468,N_4436);
nand U4583 (N_4583,N_4496,N_4492);
nand U4584 (N_4584,N_4431,N_4420);
nand U4585 (N_4585,N_4462,N_4403);
and U4586 (N_4586,N_4484,N_4481);
nor U4587 (N_4587,N_4443,N_4493);
nor U4588 (N_4588,N_4458,N_4401);
nor U4589 (N_4589,N_4456,N_4496);
and U4590 (N_4590,N_4411,N_4476);
nor U4591 (N_4591,N_4433,N_4475);
nand U4592 (N_4592,N_4435,N_4475);
nor U4593 (N_4593,N_4442,N_4486);
nand U4594 (N_4594,N_4475,N_4419);
or U4595 (N_4595,N_4418,N_4402);
nor U4596 (N_4596,N_4426,N_4442);
nor U4597 (N_4597,N_4435,N_4497);
and U4598 (N_4598,N_4461,N_4454);
nand U4599 (N_4599,N_4418,N_4437);
and U4600 (N_4600,N_4558,N_4553);
xnor U4601 (N_4601,N_4550,N_4561);
and U4602 (N_4602,N_4521,N_4584);
xnor U4603 (N_4603,N_4568,N_4589);
nand U4604 (N_4604,N_4531,N_4504);
or U4605 (N_4605,N_4534,N_4503);
and U4606 (N_4606,N_4572,N_4585);
nand U4607 (N_4607,N_4583,N_4586);
and U4608 (N_4608,N_4559,N_4508);
nor U4609 (N_4609,N_4519,N_4501);
or U4610 (N_4610,N_4563,N_4565);
or U4611 (N_4611,N_4515,N_4543);
and U4612 (N_4612,N_4540,N_4510);
or U4613 (N_4613,N_4556,N_4577);
and U4614 (N_4614,N_4535,N_4537);
nor U4615 (N_4615,N_4576,N_4598);
nand U4616 (N_4616,N_4520,N_4555);
or U4617 (N_4617,N_4545,N_4505);
nor U4618 (N_4618,N_4595,N_4599);
or U4619 (N_4619,N_4530,N_4554);
nor U4620 (N_4620,N_4526,N_4588);
xnor U4621 (N_4621,N_4529,N_4513);
and U4622 (N_4622,N_4516,N_4523);
and U4623 (N_4623,N_4567,N_4549);
nor U4624 (N_4624,N_4581,N_4594);
nor U4625 (N_4625,N_4564,N_4551);
xnor U4626 (N_4626,N_4542,N_4566);
or U4627 (N_4627,N_4514,N_4578);
nor U4628 (N_4628,N_4596,N_4591);
and U4629 (N_4629,N_4570,N_4597);
nor U4630 (N_4630,N_4552,N_4541);
nand U4631 (N_4631,N_4507,N_4582);
or U4632 (N_4632,N_4517,N_4506);
nor U4633 (N_4633,N_4546,N_4532);
nand U4634 (N_4634,N_4569,N_4580);
or U4635 (N_4635,N_4502,N_4511);
or U4636 (N_4636,N_4574,N_4538);
nor U4637 (N_4637,N_4524,N_4575);
or U4638 (N_4638,N_4557,N_4500);
xor U4639 (N_4639,N_4547,N_4527);
or U4640 (N_4640,N_4539,N_4590);
and U4641 (N_4641,N_4522,N_4560);
and U4642 (N_4642,N_4536,N_4593);
and U4643 (N_4643,N_4571,N_4509);
nand U4644 (N_4644,N_4544,N_4512);
or U4645 (N_4645,N_4579,N_4562);
nor U4646 (N_4646,N_4587,N_4525);
nor U4647 (N_4647,N_4533,N_4592);
nor U4648 (N_4648,N_4528,N_4548);
and U4649 (N_4649,N_4573,N_4518);
xnor U4650 (N_4650,N_4538,N_4519);
nor U4651 (N_4651,N_4597,N_4501);
and U4652 (N_4652,N_4558,N_4547);
and U4653 (N_4653,N_4560,N_4506);
nand U4654 (N_4654,N_4555,N_4585);
or U4655 (N_4655,N_4591,N_4541);
nor U4656 (N_4656,N_4576,N_4587);
nor U4657 (N_4657,N_4571,N_4584);
nor U4658 (N_4658,N_4580,N_4507);
and U4659 (N_4659,N_4513,N_4586);
or U4660 (N_4660,N_4522,N_4588);
nor U4661 (N_4661,N_4516,N_4565);
nor U4662 (N_4662,N_4502,N_4593);
nor U4663 (N_4663,N_4536,N_4517);
nand U4664 (N_4664,N_4598,N_4591);
xnor U4665 (N_4665,N_4586,N_4576);
and U4666 (N_4666,N_4545,N_4503);
or U4667 (N_4667,N_4507,N_4590);
nand U4668 (N_4668,N_4584,N_4553);
or U4669 (N_4669,N_4556,N_4574);
or U4670 (N_4670,N_4556,N_4582);
nand U4671 (N_4671,N_4573,N_4533);
nor U4672 (N_4672,N_4505,N_4510);
nand U4673 (N_4673,N_4522,N_4546);
nand U4674 (N_4674,N_4536,N_4589);
nand U4675 (N_4675,N_4502,N_4571);
or U4676 (N_4676,N_4503,N_4509);
and U4677 (N_4677,N_4591,N_4543);
or U4678 (N_4678,N_4539,N_4508);
or U4679 (N_4679,N_4508,N_4596);
or U4680 (N_4680,N_4569,N_4581);
or U4681 (N_4681,N_4575,N_4572);
nand U4682 (N_4682,N_4591,N_4594);
nor U4683 (N_4683,N_4587,N_4552);
or U4684 (N_4684,N_4553,N_4554);
nor U4685 (N_4685,N_4548,N_4524);
nor U4686 (N_4686,N_4559,N_4561);
xor U4687 (N_4687,N_4527,N_4594);
and U4688 (N_4688,N_4506,N_4570);
nand U4689 (N_4689,N_4540,N_4548);
nand U4690 (N_4690,N_4553,N_4588);
nand U4691 (N_4691,N_4519,N_4566);
nand U4692 (N_4692,N_4504,N_4551);
nor U4693 (N_4693,N_4580,N_4531);
nor U4694 (N_4694,N_4592,N_4525);
and U4695 (N_4695,N_4589,N_4502);
and U4696 (N_4696,N_4516,N_4533);
or U4697 (N_4697,N_4549,N_4584);
and U4698 (N_4698,N_4560,N_4586);
nand U4699 (N_4699,N_4547,N_4514);
and U4700 (N_4700,N_4688,N_4608);
or U4701 (N_4701,N_4694,N_4671);
nor U4702 (N_4702,N_4636,N_4692);
nor U4703 (N_4703,N_4675,N_4605);
nor U4704 (N_4704,N_4622,N_4614);
nand U4705 (N_4705,N_4691,N_4640);
and U4706 (N_4706,N_4615,N_4647);
nand U4707 (N_4707,N_4612,N_4646);
nor U4708 (N_4708,N_4634,N_4649);
or U4709 (N_4709,N_4655,N_4613);
nand U4710 (N_4710,N_4616,N_4681);
nor U4711 (N_4711,N_4641,N_4629);
and U4712 (N_4712,N_4673,N_4624);
and U4713 (N_4713,N_4623,N_4603);
or U4714 (N_4714,N_4672,N_4696);
nand U4715 (N_4715,N_4630,N_4682);
or U4716 (N_4716,N_4621,N_4697);
nand U4717 (N_4717,N_4650,N_4663);
nor U4718 (N_4718,N_4674,N_4678);
or U4719 (N_4719,N_4658,N_4618);
xor U4720 (N_4720,N_4652,N_4627);
nand U4721 (N_4721,N_4637,N_4687);
nand U4722 (N_4722,N_4644,N_4679);
nand U4723 (N_4723,N_4668,N_4643);
and U4724 (N_4724,N_4632,N_4662);
nor U4725 (N_4725,N_4653,N_4659);
nor U4726 (N_4726,N_4695,N_4628);
or U4727 (N_4727,N_4656,N_4683);
or U4728 (N_4728,N_4689,N_4690);
nand U4729 (N_4729,N_4617,N_4638);
and U4730 (N_4730,N_4664,N_4699);
or U4731 (N_4731,N_4669,N_4600);
and U4732 (N_4732,N_4633,N_4670);
xor U4733 (N_4733,N_4642,N_4625);
nor U4734 (N_4734,N_4604,N_4665);
or U4735 (N_4735,N_4680,N_4610);
and U4736 (N_4736,N_4645,N_4684);
nor U4737 (N_4737,N_4609,N_4635);
or U4738 (N_4738,N_4619,N_4611);
nor U4739 (N_4739,N_4620,N_4606);
and U4740 (N_4740,N_4698,N_4654);
and U4741 (N_4741,N_4685,N_4666);
and U4742 (N_4742,N_4607,N_4631);
or U4743 (N_4743,N_4661,N_4639);
nand U4744 (N_4744,N_4626,N_4657);
nand U4745 (N_4745,N_4677,N_4667);
xnor U4746 (N_4746,N_4686,N_4602);
and U4747 (N_4747,N_4601,N_4660);
nand U4748 (N_4748,N_4693,N_4651);
nand U4749 (N_4749,N_4676,N_4648);
nor U4750 (N_4750,N_4600,N_4678);
nand U4751 (N_4751,N_4639,N_4660);
or U4752 (N_4752,N_4600,N_4666);
or U4753 (N_4753,N_4613,N_4629);
nor U4754 (N_4754,N_4682,N_4609);
nand U4755 (N_4755,N_4675,N_4678);
nand U4756 (N_4756,N_4614,N_4644);
nand U4757 (N_4757,N_4658,N_4647);
nand U4758 (N_4758,N_4654,N_4610);
nand U4759 (N_4759,N_4695,N_4665);
and U4760 (N_4760,N_4654,N_4618);
nand U4761 (N_4761,N_4661,N_4618);
and U4762 (N_4762,N_4624,N_4613);
or U4763 (N_4763,N_4653,N_4605);
nand U4764 (N_4764,N_4665,N_4620);
nor U4765 (N_4765,N_4607,N_4671);
or U4766 (N_4766,N_4639,N_4695);
nand U4767 (N_4767,N_4600,N_4667);
or U4768 (N_4768,N_4664,N_4640);
or U4769 (N_4769,N_4604,N_4657);
or U4770 (N_4770,N_4627,N_4636);
nor U4771 (N_4771,N_4640,N_4686);
nand U4772 (N_4772,N_4649,N_4640);
nand U4773 (N_4773,N_4605,N_4609);
nor U4774 (N_4774,N_4635,N_4676);
and U4775 (N_4775,N_4646,N_4652);
nor U4776 (N_4776,N_4639,N_4680);
nand U4777 (N_4777,N_4630,N_4695);
nand U4778 (N_4778,N_4667,N_4619);
and U4779 (N_4779,N_4620,N_4636);
nor U4780 (N_4780,N_4623,N_4649);
or U4781 (N_4781,N_4606,N_4621);
nor U4782 (N_4782,N_4662,N_4698);
or U4783 (N_4783,N_4602,N_4661);
nor U4784 (N_4784,N_4667,N_4632);
and U4785 (N_4785,N_4666,N_4678);
nand U4786 (N_4786,N_4604,N_4685);
and U4787 (N_4787,N_4605,N_4634);
nor U4788 (N_4788,N_4651,N_4672);
and U4789 (N_4789,N_4637,N_4608);
and U4790 (N_4790,N_4656,N_4607);
and U4791 (N_4791,N_4637,N_4628);
or U4792 (N_4792,N_4630,N_4693);
and U4793 (N_4793,N_4606,N_4672);
and U4794 (N_4794,N_4659,N_4630);
nand U4795 (N_4795,N_4697,N_4640);
or U4796 (N_4796,N_4658,N_4641);
nor U4797 (N_4797,N_4646,N_4665);
nor U4798 (N_4798,N_4609,N_4658);
nand U4799 (N_4799,N_4647,N_4673);
or U4800 (N_4800,N_4717,N_4751);
or U4801 (N_4801,N_4779,N_4796);
or U4802 (N_4802,N_4724,N_4787);
nand U4803 (N_4803,N_4754,N_4708);
and U4804 (N_4804,N_4721,N_4767);
nor U4805 (N_4805,N_4748,N_4734);
or U4806 (N_4806,N_4784,N_4781);
nor U4807 (N_4807,N_4740,N_4762);
nor U4808 (N_4808,N_4770,N_4798);
or U4809 (N_4809,N_4722,N_4750);
and U4810 (N_4810,N_4714,N_4725);
nor U4811 (N_4811,N_4764,N_4704);
nand U4812 (N_4812,N_4755,N_4732);
xnor U4813 (N_4813,N_4774,N_4705);
nor U4814 (N_4814,N_4752,N_4726);
and U4815 (N_4815,N_4793,N_4733);
nand U4816 (N_4816,N_4744,N_4749);
or U4817 (N_4817,N_4735,N_4706);
nor U4818 (N_4818,N_4763,N_4707);
nand U4819 (N_4819,N_4772,N_4747);
nand U4820 (N_4820,N_4701,N_4777);
nand U4821 (N_4821,N_4765,N_4775);
or U4822 (N_4822,N_4757,N_4745);
and U4823 (N_4823,N_4761,N_4753);
nor U4824 (N_4824,N_4795,N_4728);
and U4825 (N_4825,N_4758,N_4737);
nand U4826 (N_4826,N_4746,N_4743);
and U4827 (N_4827,N_4742,N_4771);
nor U4828 (N_4828,N_4785,N_4778);
and U4829 (N_4829,N_4712,N_4716);
or U4830 (N_4830,N_4790,N_4702);
or U4831 (N_4831,N_4703,N_4782);
or U4832 (N_4832,N_4792,N_4719);
xor U4833 (N_4833,N_4715,N_4760);
nor U4834 (N_4834,N_4768,N_4731);
nand U4835 (N_4835,N_4710,N_4700);
nor U4836 (N_4836,N_4730,N_4723);
or U4837 (N_4837,N_4729,N_4736);
nand U4838 (N_4838,N_4739,N_4759);
and U4839 (N_4839,N_4797,N_4791);
or U4840 (N_4840,N_4766,N_4738);
xnor U4841 (N_4841,N_4788,N_4794);
xor U4842 (N_4842,N_4783,N_4769);
and U4843 (N_4843,N_4727,N_4718);
or U4844 (N_4844,N_4720,N_4786);
nor U4845 (N_4845,N_4773,N_4756);
nor U4846 (N_4846,N_4741,N_4711);
or U4847 (N_4847,N_4713,N_4780);
or U4848 (N_4848,N_4799,N_4776);
or U4849 (N_4849,N_4709,N_4789);
or U4850 (N_4850,N_4720,N_4714);
or U4851 (N_4851,N_4704,N_4761);
nor U4852 (N_4852,N_4732,N_4707);
or U4853 (N_4853,N_4703,N_4728);
nand U4854 (N_4854,N_4799,N_4761);
or U4855 (N_4855,N_4706,N_4769);
nand U4856 (N_4856,N_4766,N_4798);
or U4857 (N_4857,N_4757,N_4732);
and U4858 (N_4858,N_4703,N_4766);
or U4859 (N_4859,N_4732,N_4713);
nand U4860 (N_4860,N_4740,N_4731);
and U4861 (N_4861,N_4764,N_4777);
xnor U4862 (N_4862,N_4720,N_4776);
or U4863 (N_4863,N_4700,N_4727);
nor U4864 (N_4864,N_4726,N_4715);
or U4865 (N_4865,N_4798,N_4748);
or U4866 (N_4866,N_4789,N_4705);
nand U4867 (N_4867,N_4760,N_4707);
or U4868 (N_4868,N_4706,N_4763);
or U4869 (N_4869,N_4765,N_4777);
nand U4870 (N_4870,N_4779,N_4773);
nor U4871 (N_4871,N_4731,N_4757);
or U4872 (N_4872,N_4795,N_4774);
or U4873 (N_4873,N_4799,N_4716);
nor U4874 (N_4874,N_4722,N_4771);
nor U4875 (N_4875,N_4799,N_4709);
or U4876 (N_4876,N_4792,N_4795);
nor U4877 (N_4877,N_4753,N_4732);
nand U4878 (N_4878,N_4740,N_4759);
nor U4879 (N_4879,N_4707,N_4781);
nor U4880 (N_4880,N_4785,N_4788);
nor U4881 (N_4881,N_4714,N_4749);
nand U4882 (N_4882,N_4783,N_4799);
and U4883 (N_4883,N_4763,N_4764);
nor U4884 (N_4884,N_4738,N_4764);
nor U4885 (N_4885,N_4711,N_4713);
nand U4886 (N_4886,N_4752,N_4750);
and U4887 (N_4887,N_4755,N_4763);
and U4888 (N_4888,N_4775,N_4782);
and U4889 (N_4889,N_4745,N_4772);
nand U4890 (N_4890,N_4798,N_4740);
and U4891 (N_4891,N_4799,N_4770);
and U4892 (N_4892,N_4742,N_4728);
and U4893 (N_4893,N_4777,N_4797);
xor U4894 (N_4894,N_4777,N_4729);
nand U4895 (N_4895,N_4738,N_4781);
or U4896 (N_4896,N_4706,N_4788);
and U4897 (N_4897,N_4781,N_4745);
or U4898 (N_4898,N_4769,N_4724);
nand U4899 (N_4899,N_4785,N_4728);
nand U4900 (N_4900,N_4833,N_4856);
and U4901 (N_4901,N_4841,N_4842);
nor U4902 (N_4902,N_4837,N_4851);
and U4903 (N_4903,N_4810,N_4883);
and U4904 (N_4904,N_4882,N_4878);
or U4905 (N_4905,N_4846,N_4891);
or U4906 (N_4906,N_4864,N_4853);
nand U4907 (N_4907,N_4821,N_4879);
nand U4908 (N_4908,N_4824,N_4835);
nand U4909 (N_4909,N_4805,N_4844);
nand U4910 (N_4910,N_4814,N_4852);
or U4911 (N_4911,N_4880,N_4802);
and U4912 (N_4912,N_4872,N_4830);
or U4913 (N_4913,N_4800,N_4858);
or U4914 (N_4914,N_4867,N_4850);
and U4915 (N_4915,N_4893,N_4827);
nand U4916 (N_4916,N_4801,N_4874);
or U4917 (N_4917,N_4855,N_4897);
nor U4918 (N_4918,N_4848,N_4825);
nand U4919 (N_4919,N_4899,N_4840);
or U4920 (N_4920,N_4888,N_4822);
nand U4921 (N_4921,N_4873,N_4826);
nand U4922 (N_4922,N_4804,N_4843);
or U4923 (N_4923,N_4865,N_4859);
nor U4924 (N_4924,N_4871,N_4870);
or U4925 (N_4925,N_4807,N_4890);
nand U4926 (N_4926,N_4887,N_4886);
nand U4927 (N_4927,N_4839,N_4862);
nand U4928 (N_4928,N_4817,N_4892);
and U4929 (N_4929,N_4863,N_4895);
nor U4930 (N_4930,N_4828,N_4815);
nand U4931 (N_4931,N_4884,N_4838);
or U4932 (N_4932,N_4806,N_4829);
and U4933 (N_4933,N_4877,N_4894);
and U4934 (N_4934,N_4803,N_4866);
nor U4935 (N_4935,N_4818,N_4869);
nor U4936 (N_4936,N_4868,N_4831);
or U4937 (N_4937,N_4898,N_4896);
or U4938 (N_4938,N_4836,N_4813);
nor U4939 (N_4939,N_4808,N_4816);
or U4940 (N_4940,N_4857,N_4811);
nand U4941 (N_4941,N_4812,N_4876);
or U4942 (N_4942,N_4889,N_4885);
and U4943 (N_4943,N_4819,N_4860);
nand U4944 (N_4944,N_4823,N_4849);
or U4945 (N_4945,N_4861,N_4875);
and U4946 (N_4946,N_4845,N_4834);
or U4947 (N_4947,N_4854,N_4881);
or U4948 (N_4948,N_4809,N_4847);
or U4949 (N_4949,N_4832,N_4820);
nand U4950 (N_4950,N_4830,N_4899);
nor U4951 (N_4951,N_4845,N_4838);
or U4952 (N_4952,N_4853,N_4861);
nand U4953 (N_4953,N_4847,N_4807);
nor U4954 (N_4954,N_4847,N_4827);
nand U4955 (N_4955,N_4893,N_4871);
and U4956 (N_4956,N_4850,N_4880);
nand U4957 (N_4957,N_4832,N_4880);
nor U4958 (N_4958,N_4887,N_4831);
or U4959 (N_4959,N_4863,N_4869);
or U4960 (N_4960,N_4858,N_4812);
nor U4961 (N_4961,N_4830,N_4833);
nand U4962 (N_4962,N_4873,N_4886);
nor U4963 (N_4963,N_4892,N_4894);
and U4964 (N_4964,N_4833,N_4859);
and U4965 (N_4965,N_4828,N_4827);
or U4966 (N_4966,N_4860,N_4811);
nand U4967 (N_4967,N_4828,N_4871);
nand U4968 (N_4968,N_4876,N_4840);
or U4969 (N_4969,N_4858,N_4804);
or U4970 (N_4970,N_4858,N_4861);
and U4971 (N_4971,N_4897,N_4869);
nand U4972 (N_4972,N_4811,N_4835);
nand U4973 (N_4973,N_4805,N_4853);
nor U4974 (N_4974,N_4809,N_4854);
nand U4975 (N_4975,N_4857,N_4886);
nand U4976 (N_4976,N_4830,N_4879);
nor U4977 (N_4977,N_4802,N_4814);
or U4978 (N_4978,N_4865,N_4802);
nor U4979 (N_4979,N_4895,N_4807);
and U4980 (N_4980,N_4852,N_4808);
nor U4981 (N_4981,N_4834,N_4830);
nand U4982 (N_4982,N_4845,N_4872);
and U4983 (N_4983,N_4883,N_4817);
nor U4984 (N_4984,N_4877,N_4814);
or U4985 (N_4985,N_4878,N_4811);
nor U4986 (N_4986,N_4889,N_4871);
nor U4987 (N_4987,N_4803,N_4873);
and U4988 (N_4988,N_4801,N_4806);
nand U4989 (N_4989,N_4889,N_4803);
and U4990 (N_4990,N_4825,N_4896);
and U4991 (N_4991,N_4899,N_4880);
nand U4992 (N_4992,N_4821,N_4814);
or U4993 (N_4993,N_4868,N_4842);
or U4994 (N_4994,N_4896,N_4877);
nand U4995 (N_4995,N_4857,N_4819);
or U4996 (N_4996,N_4870,N_4880);
xor U4997 (N_4997,N_4839,N_4824);
nand U4998 (N_4998,N_4855,N_4867);
or U4999 (N_4999,N_4822,N_4831);
nand UO_0 (O_0,N_4948,N_4922);
nand UO_1 (O_1,N_4928,N_4979);
and UO_2 (O_2,N_4972,N_4907);
or UO_3 (O_3,N_4967,N_4943);
and UO_4 (O_4,N_4906,N_4952);
or UO_5 (O_5,N_4926,N_4921);
nor UO_6 (O_6,N_4959,N_4991);
and UO_7 (O_7,N_4932,N_4912);
or UO_8 (O_8,N_4960,N_4949);
nand UO_9 (O_9,N_4974,N_4951);
or UO_10 (O_10,N_4930,N_4913);
or UO_11 (O_11,N_4941,N_4973);
nand UO_12 (O_12,N_4953,N_4929);
xor UO_13 (O_13,N_4900,N_4927);
xor UO_14 (O_14,N_4999,N_4924);
or UO_15 (O_15,N_4918,N_4919);
xor UO_16 (O_16,N_4954,N_4980);
and UO_17 (O_17,N_4997,N_4984);
or UO_18 (O_18,N_4988,N_4917);
or UO_19 (O_19,N_4940,N_4990);
nor UO_20 (O_20,N_4944,N_4933);
or UO_21 (O_21,N_4904,N_4942);
nor UO_22 (O_22,N_4986,N_4958);
or UO_23 (O_23,N_4946,N_4910);
and UO_24 (O_24,N_4903,N_4985);
nand UO_25 (O_25,N_4905,N_4908);
nor UO_26 (O_26,N_4971,N_4966);
nand UO_27 (O_27,N_4982,N_4992);
nor UO_28 (O_28,N_4976,N_4996);
nand UO_29 (O_29,N_4938,N_4931);
nor UO_30 (O_30,N_4975,N_4947);
and UO_31 (O_31,N_4920,N_4995);
nand UO_32 (O_32,N_4935,N_4977);
nand UO_33 (O_33,N_4945,N_4969);
nor UO_34 (O_34,N_4978,N_4909);
and UO_35 (O_35,N_4939,N_4925);
or UO_36 (O_36,N_4911,N_4989);
nor UO_37 (O_37,N_4970,N_4957);
nor UO_38 (O_38,N_4998,N_4923);
nor UO_39 (O_39,N_4902,N_4901);
xnor UO_40 (O_40,N_4983,N_4987);
or UO_41 (O_41,N_4962,N_4968);
or UO_42 (O_42,N_4964,N_4950);
nor UO_43 (O_43,N_4937,N_4961);
nand UO_44 (O_44,N_4915,N_4963);
nor UO_45 (O_45,N_4934,N_4993);
nand UO_46 (O_46,N_4916,N_4981);
or UO_47 (O_47,N_4994,N_4956);
or UO_48 (O_48,N_4936,N_4955);
nor UO_49 (O_49,N_4914,N_4965);
nor UO_50 (O_50,N_4905,N_4931);
and UO_51 (O_51,N_4911,N_4967);
or UO_52 (O_52,N_4952,N_4932);
or UO_53 (O_53,N_4917,N_4921);
nor UO_54 (O_54,N_4920,N_4935);
nor UO_55 (O_55,N_4991,N_4901);
nand UO_56 (O_56,N_4920,N_4983);
and UO_57 (O_57,N_4981,N_4982);
xor UO_58 (O_58,N_4940,N_4937);
nand UO_59 (O_59,N_4973,N_4926);
or UO_60 (O_60,N_4944,N_4962);
nor UO_61 (O_61,N_4942,N_4917);
nand UO_62 (O_62,N_4915,N_4996);
nor UO_63 (O_63,N_4953,N_4984);
nor UO_64 (O_64,N_4907,N_4986);
xnor UO_65 (O_65,N_4979,N_4946);
and UO_66 (O_66,N_4972,N_4984);
nor UO_67 (O_67,N_4906,N_4964);
or UO_68 (O_68,N_4973,N_4922);
and UO_69 (O_69,N_4958,N_4963);
nand UO_70 (O_70,N_4960,N_4911);
and UO_71 (O_71,N_4907,N_4966);
nand UO_72 (O_72,N_4937,N_4921);
nor UO_73 (O_73,N_4901,N_4912);
nand UO_74 (O_74,N_4924,N_4907);
nor UO_75 (O_75,N_4904,N_4949);
or UO_76 (O_76,N_4934,N_4982);
or UO_77 (O_77,N_4979,N_4986);
nand UO_78 (O_78,N_4905,N_4918);
and UO_79 (O_79,N_4964,N_4959);
nand UO_80 (O_80,N_4973,N_4901);
and UO_81 (O_81,N_4963,N_4986);
nand UO_82 (O_82,N_4903,N_4933);
nand UO_83 (O_83,N_4960,N_4928);
nand UO_84 (O_84,N_4938,N_4966);
or UO_85 (O_85,N_4920,N_4919);
and UO_86 (O_86,N_4985,N_4937);
nand UO_87 (O_87,N_4962,N_4955);
nor UO_88 (O_88,N_4931,N_4980);
nor UO_89 (O_89,N_4999,N_4972);
nand UO_90 (O_90,N_4927,N_4962);
nand UO_91 (O_91,N_4904,N_4935);
and UO_92 (O_92,N_4908,N_4997);
xor UO_93 (O_93,N_4915,N_4923);
and UO_94 (O_94,N_4900,N_4968);
nand UO_95 (O_95,N_4989,N_4909);
nor UO_96 (O_96,N_4988,N_4928);
and UO_97 (O_97,N_4909,N_4963);
or UO_98 (O_98,N_4961,N_4972);
nor UO_99 (O_99,N_4993,N_4994);
or UO_100 (O_100,N_4909,N_4986);
nand UO_101 (O_101,N_4994,N_4923);
or UO_102 (O_102,N_4902,N_4996);
nor UO_103 (O_103,N_4988,N_4960);
xor UO_104 (O_104,N_4968,N_4944);
and UO_105 (O_105,N_4980,N_4977);
or UO_106 (O_106,N_4978,N_4958);
nand UO_107 (O_107,N_4935,N_4973);
or UO_108 (O_108,N_4939,N_4952);
nand UO_109 (O_109,N_4977,N_4999);
and UO_110 (O_110,N_4975,N_4920);
nand UO_111 (O_111,N_4961,N_4903);
nand UO_112 (O_112,N_4942,N_4976);
or UO_113 (O_113,N_4953,N_4961);
or UO_114 (O_114,N_4911,N_4939);
nand UO_115 (O_115,N_4968,N_4987);
nor UO_116 (O_116,N_4909,N_4999);
xor UO_117 (O_117,N_4921,N_4959);
or UO_118 (O_118,N_4958,N_4980);
nand UO_119 (O_119,N_4943,N_4945);
nand UO_120 (O_120,N_4972,N_4955);
or UO_121 (O_121,N_4904,N_4901);
nor UO_122 (O_122,N_4941,N_4919);
or UO_123 (O_123,N_4916,N_4900);
and UO_124 (O_124,N_4960,N_4909);
or UO_125 (O_125,N_4903,N_4964);
nand UO_126 (O_126,N_4900,N_4974);
nand UO_127 (O_127,N_4984,N_4985);
and UO_128 (O_128,N_4922,N_4938);
nand UO_129 (O_129,N_4971,N_4947);
or UO_130 (O_130,N_4902,N_4958);
nand UO_131 (O_131,N_4976,N_4904);
nor UO_132 (O_132,N_4982,N_4994);
and UO_133 (O_133,N_4974,N_4991);
nor UO_134 (O_134,N_4918,N_4910);
nor UO_135 (O_135,N_4969,N_4904);
nor UO_136 (O_136,N_4932,N_4974);
nand UO_137 (O_137,N_4904,N_4943);
nor UO_138 (O_138,N_4961,N_4984);
and UO_139 (O_139,N_4923,N_4946);
nor UO_140 (O_140,N_4980,N_4975);
and UO_141 (O_141,N_4999,N_4941);
or UO_142 (O_142,N_4943,N_4902);
or UO_143 (O_143,N_4993,N_4958);
and UO_144 (O_144,N_4922,N_4911);
nor UO_145 (O_145,N_4976,N_4975);
xor UO_146 (O_146,N_4922,N_4993);
nand UO_147 (O_147,N_4958,N_4985);
nand UO_148 (O_148,N_4962,N_4926);
nand UO_149 (O_149,N_4975,N_4951);
or UO_150 (O_150,N_4916,N_4936);
nand UO_151 (O_151,N_4963,N_4987);
or UO_152 (O_152,N_4987,N_4992);
or UO_153 (O_153,N_4972,N_4928);
nand UO_154 (O_154,N_4903,N_4945);
nand UO_155 (O_155,N_4917,N_4939);
xnor UO_156 (O_156,N_4912,N_4900);
and UO_157 (O_157,N_4956,N_4999);
nor UO_158 (O_158,N_4952,N_4962);
or UO_159 (O_159,N_4927,N_4983);
or UO_160 (O_160,N_4924,N_4979);
nand UO_161 (O_161,N_4909,N_4979);
or UO_162 (O_162,N_4915,N_4911);
or UO_163 (O_163,N_4903,N_4976);
nor UO_164 (O_164,N_4964,N_4973);
and UO_165 (O_165,N_4966,N_4956);
or UO_166 (O_166,N_4960,N_4975);
or UO_167 (O_167,N_4967,N_4984);
nand UO_168 (O_168,N_4942,N_4907);
nand UO_169 (O_169,N_4976,N_4957);
xor UO_170 (O_170,N_4972,N_4952);
nand UO_171 (O_171,N_4906,N_4961);
xor UO_172 (O_172,N_4916,N_4914);
and UO_173 (O_173,N_4986,N_4906);
and UO_174 (O_174,N_4991,N_4912);
or UO_175 (O_175,N_4904,N_4987);
nand UO_176 (O_176,N_4922,N_4999);
nor UO_177 (O_177,N_4922,N_4950);
or UO_178 (O_178,N_4985,N_4961);
and UO_179 (O_179,N_4963,N_4941);
nor UO_180 (O_180,N_4965,N_4998);
nor UO_181 (O_181,N_4920,N_4922);
nor UO_182 (O_182,N_4929,N_4957);
and UO_183 (O_183,N_4921,N_4972);
or UO_184 (O_184,N_4943,N_4927);
and UO_185 (O_185,N_4994,N_4954);
xnor UO_186 (O_186,N_4908,N_4921);
and UO_187 (O_187,N_4908,N_4907);
nor UO_188 (O_188,N_4970,N_4968);
nand UO_189 (O_189,N_4919,N_4987);
and UO_190 (O_190,N_4902,N_4949);
xor UO_191 (O_191,N_4995,N_4901);
or UO_192 (O_192,N_4958,N_4983);
nand UO_193 (O_193,N_4935,N_4962);
nand UO_194 (O_194,N_4987,N_4947);
and UO_195 (O_195,N_4991,N_4953);
nor UO_196 (O_196,N_4985,N_4983);
and UO_197 (O_197,N_4910,N_4938);
nor UO_198 (O_198,N_4912,N_4911);
nand UO_199 (O_199,N_4985,N_4975);
nor UO_200 (O_200,N_4998,N_4902);
nor UO_201 (O_201,N_4912,N_4960);
nand UO_202 (O_202,N_4939,N_4919);
or UO_203 (O_203,N_4963,N_4983);
nand UO_204 (O_204,N_4923,N_4922);
nor UO_205 (O_205,N_4965,N_4948);
and UO_206 (O_206,N_4909,N_4982);
and UO_207 (O_207,N_4924,N_4908);
nand UO_208 (O_208,N_4958,N_4956);
nand UO_209 (O_209,N_4925,N_4910);
and UO_210 (O_210,N_4986,N_4950);
and UO_211 (O_211,N_4987,N_4962);
xor UO_212 (O_212,N_4952,N_4949);
nor UO_213 (O_213,N_4919,N_4950);
and UO_214 (O_214,N_4933,N_4917);
or UO_215 (O_215,N_4977,N_4962);
or UO_216 (O_216,N_4949,N_4989);
and UO_217 (O_217,N_4912,N_4981);
or UO_218 (O_218,N_4987,N_4981);
nor UO_219 (O_219,N_4964,N_4914);
nor UO_220 (O_220,N_4922,N_4967);
and UO_221 (O_221,N_4916,N_4913);
nor UO_222 (O_222,N_4904,N_4910);
nor UO_223 (O_223,N_4986,N_4994);
or UO_224 (O_224,N_4998,N_4977);
nand UO_225 (O_225,N_4996,N_4927);
and UO_226 (O_226,N_4928,N_4938);
and UO_227 (O_227,N_4916,N_4922);
or UO_228 (O_228,N_4967,N_4903);
or UO_229 (O_229,N_4924,N_4917);
or UO_230 (O_230,N_4959,N_4950);
nor UO_231 (O_231,N_4934,N_4974);
nand UO_232 (O_232,N_4935,N_4921);
or UO_233 (O_233,N_4984,N_4992);
nand UO_234 (O_234,N_4974,N_4975);
nor UO_235 (O_235,N_4929,N_4937);
nor UO_236 (O_236,N_4984,N_4921);
nor UO_237 (O_237,N_4900,N_4998);
nand UO_238 (O_238,N_4933,N_4925);
and UO_239 (O_239,N_4904,N_4914);
nand UO_240 (O_240,N_4972,N_4903);
nor UO_241 (O_241,N_4921,N_4933);
or UO_242 (O_242,N_4914,N_4929);
nand UO_243 (O_243,N_4906,N_4955);
nor UO_244 (O_244,N_4945,N_4905);
and UO_245 (O_245,N_4918,N_4986);
nand UO_246 (O_246,N_4946,N_4936);
xor UO_247 (O_247,N_4916,N_4908);
or UO_248 (O_248,N_4997,N_4976);
and UO_249 (O_249,N_4952,N_4976);
nand UO_250 (O_250,N_4967,N_4924);
xnor UO_251 (O_251,N_4993,N_4975);
and UO_252 (O_252,N_4937,N_4953);
or UO_253 (O_253,N_4952,N_4969);
nand UO_254 (O_254,N_4916,N_4938);
and UO_255 (O_255,N_4930,N_4949);
nand UO_256 (O_256,N_4922,N_4915);
or UO_257 (O_257,N_4982,N_4943);
xor UO_258 (O_258,N_4969,N_4920);
nand UO_259 (O_259,N_4978,N_4902);
and UO_260 (O_260,N_4936,N_4930);
and UO_261 (O_261,N_4915,N_4913);
or UO_262 (O_262,N_4954,N_4928);
nand UO_263 (O_263,N_4915,N_4916);
nor UO_264 (O_264,N_4916,N_4973);
or UO_265 (O_265,N_4903,N_4932);
nor UO_266 (O_266,N_4987,N_4933);
nor UO_267 (O_267,N_4956,N_4930);
and UO_268 (O_268,N_4969,N_4993);
nand UO_269 (O_269,N_4970,N_4918);
or UO_270 (O_270,N_4923,N_4958);
nand UO_271 (O_271,N_4987,N_4964);
xnor UO_272 (O_272,N_4917,N_4975);
nand UO_273 (O_273,N_4953,N_4915);
and UO_274 (O_274,N_4928,N_4937);
or UO_275 (O_275,N_4979,N_4978);
or UO_276 (O_276,N_4947,N_4904);
nor UO_277 (O_277,N_4970,N_4926);
nor UO_278 (O_278,N_4977,N_4947);
and UO_279 (O_279,N_4947,N_4914);
or UO_280 (O_280,N_4907,N_4961);
nand UO_281 (O_281,N_4974,N_4942);
nand UO_282 (O_282,N_4911,N_4959);
and UO_283 (O_283,N_4924,N_4912);
nor UO_284 (O_284,N_4975,N_4946);
nand UO_285 (O_285,N_4985,N_4970);
or UO_286 (O_286,N_4917,N_4934);
or UO_287 (O_287,N_4990,N_4950);
and UO_288 (O_288,N_4924,N_4998);
and UO_289 (O_289,N_4943,N_4957);
nor UO_290 (O_290,N_4956,N_4976);
nor UO_291 (O_291,N_4929,N_4911);
nand UO_292 (O_292,N_4926,N_4984);
or UO_293 (O_293,N_4910,N_4978);
and UO_294 (O_294,N_4914,N_4910);
nor UO_295 (O_295,N_4934,N_4954);
or UO_296 (O_296,N_4929,N_4919);
nand UO_297 (O_297,N_4917,N_4948);
and UO_298 (O_298,N_4950,N_4968);
nand UO_299 (O_299,N_4927,N_4967);
and UO_300 (O_300,N_4921,N_4999);
nor UO_301 (O_301,N_4960,N_4997);
nor UO_302 (O_302,N_4928,N_4909);
nor UO_303 (O_303,N_4967,N_4934);
and UO_304 (O_304,N_4938,N_4994);
nand UO_305 (O_305,N_4981,N_4904);
nor UO_306 (O_306,N_4984,N_4932);
or UO_307 (O_307,N_4911,N_4934);
or UO_308 (O_308,N_4910,N_4972);
nor UO_309 (O_309,N_4982,N_4900);
or UO_310 (O_310,N_4960,N_4921);
nand UO_311 (O_311,N_4967,N_4925);
nand UO_312 (O_312,N_4952,N_4942);
or UO_313 (O_313,N_4952,N_4984);
nor UO_314 (O_314,N_4942,N_4994);
nand UO_315 (O_315,N_4915,N_4959);
or UO_316 (O_316,N_4911,N_4979);
xnor UO_317 (O_317,N_4993,N_4952);
or UO_318 (O_318,N_4987,N_4939);
and UO_319 (O_319,N_4921,N_4962);
nand UO_320 (O_320,N_4945,N_4938);
nor UO_321 (O_321,N_4991,N_4975);
and UO_322 (O_322,N_4980,N_4953);
nand UO_323 (O_323,N_4976,N_4984);
and UO_324 (O_324,N_4969,N_4984);
and UO_325 (O_325,N_4928,N_4922);
or UO_326 (O_326,N_4935,N_4947);
or UO_327 (O_327,N_4948,N_4920);
nand UO_328 (O_328,N_4934,N_4994);
and UO_329 (O_329,N_4993,N_4974);
nor UO_330 (O_330,N_4905,N_4928);
nor UO_331 (O_331,N_4952,N_4973);
and UO_332 (O_332,N_4961,N_4962);
nor UO_333 (O_333,N_4933,N_4956);
nand UO_334 (O_334,N_4903,N_4994);
nor UO_335 (O_335,N_4908,N_4981);
or UO_336 (O_336,N_4902,N_4935);
nand UO_337 (O_337,N_4926,N_4969);
nor UO_338 (O_338,N_4942,N_4968);
and UO_339 (O_339,N_4968,N_4936);
nand UO_340 (O_340,N_4952,N_4902);
or UO_341 (O_341,N_4966,N_4924);
or UO_342 (O_342,N_4942,N_4909);
or UO_343 (O_343,N_4960,N_4966);
nand UO_344 (O_344,N_4987,N_4988);
and UO_345 (O_345,N_4906,N_4933);
or UO_346 (O_346,N_4993,N_4989);
or UO_347 (O_347,N_4989,N_4995);
nand UO_348 (O_348,N_4964,N_4980);
nor UO_349 (O_349,N_4944,N_4919);
nand UO_350 (O_350,N_4910,N_4986);
or UO_351 (O_351,N_4970,N_4910);
or UO_352 (O_352,N_4928,N_4949);
or UO_353 (O_353,N_4922,N_4968);
and UO_354 (O_354,N_4917,N_4967);
nand UO_355 (O_355,N_4983,N_4907);
and UO_356 (O_356,N_4998,N_4937);
and UO_357 (O_357,N_4909,N_4952);
and UO_358 (O_358,N_4927,N_4914);
and UO_359 (O_359,N_4990,N_4903);
xnor UO_360 (O_360,N_4953,N_4954);
nor UO_361 (O_361,N_4930,N_4940);
and UO_362 (O_362,N_4989,N_4903);
or UO_363 (O_363,N_4970,N_4931);
and UO_364 (O_364,N_4979,N_4900);
nor UO_365 (O_365,N_4901,N_4972);
and UO_366 (O_366,N_4939,N_4905);
nor UO_367 (O_367,N_4990,N_4913);
nor UO_368 (O_368,N_4995,N_4974);
or UO_369 (O_369,N_4983,N_4960);
xor UO_370 (O_370,N_4981,N_4936);
or UO_371 (O_371,N_4955,N_4961);
nand UO_372 (O_372,N_4972,N_4956);
and UO_373 (O_373,N_4974,N_4926);
nand UO_374 (O_374,N_4977,N_4931);
or UO_375 (O_375,N_4904,N_4998);
or UO_376 (O_376,N_4980,N_4900);
and UO_377 (O_377,N_4950,N_4963);
and UO_378 (O_378,N_4991,N_4931);
or UO_379 (O_379,N_4905,N_4927);
and UO_380 (O_380,N_4903,N_4914);
and UO_381 (O_381,N_4900,N_4947);
and UO_382 (O_382,N_4966,N_4977);
or UO_383 (O_383,N_4991,N_4923);
nor UO_384 (O_384,N_4973,N_4986);
and UO_385 (O_385,N_4937,N_4992);
nand UO_386 (O_386,N_4960,N_4990);
and UO_387 (O_387,N_4938,N_4997);
nor UO_388 (O_388,N_4980,N_4948);
and UO_389 (O_389,N_4956,N_4959);
or UO_390 (O_390,N_4946,N_4913);
and UO_391 (O_391,N_4917,N_4981);
xnor UO_392 (O_392,N_4928,N_4991);
nor UO_393 (O_393,N_4962,N_4996);
nand UO_394 (O_394,N_4931,N_4997);
and UO_395 (O_395,N_4998,N_4985);
nor UO_396 (O_396,N_4986,N_4937);
nand UO_397 (O_397,N_4934,N_4922);
nor UO_398 (O_398,N_4985,N_4913);
nor UO_399 (O_399,N_4951,N_4925);
nor UO_400 (O_400,N_4963,N_4912);
or UO_401 (O_401,N_4906,N_4947);
and UO_402 (O_402,N_4909,N_4931);
nand UO_403 (O_403,N_4931,N_4941);
or UO_404 (O_404,N_4964,N_4979);
nor UO_405 (O_405,N_4912,N_4998);
nor UO_406 (O_406,N_4953,N_4998);
or UO_407 (O_407,N_4922,N_4986);
nand UO_408 (O_408,N_4952,N_4988);
nand UO_409 (O_409,N_4947,N_4911);
nor UO_410 (O_410,N_4987,N_4984);
nand UO_411 (O_411,N_4921,N_4987);
xnor UO_412 (O_412,N_4926,N_4916);
nor UO_413 (O_413,N_4963,N_4927);
or UO_414 (O_414,N_4911,N_4971);
and UO_415 (O_415,N_4918,N_4992);
nor UO_416 (O_416,N_4992,N_4922);
xnor UO_417 (O_417,N_4938,N_4943);
nand UO_418 (O_418,N_4989,N_4921);
xor UO_419 (O_419,N_4967,N_4994);
and UO_420 (O_420,N_4925,N_4913);
and UO_421 (O_421,N_4950,N_4999);
and UO_422 (O_422,N_4979,N_4980);
nor UO_423 (O_423,N_4998,N_4922);
nor UO_424 (O_424,N_4973,N_4997);
or UO_425 (O_425,N_4953,N_4993);
nor UO_426 (O_426,N_4915,N_4975);
nor UO_427 (O_427,N_4932,N_4966);
and UO_428 (O_428,N_4947,N_4910);
nor UO_429 (O_429,N_4976,N_4922);
nand UO_430 (O_430,N_4924,N_4965);
and UO_431 (O_431,N_4968,N_4930);
nand UO_432 (O_432,N_4956,N_4916);
or UO_433 (O_433,N_4986,N_4926);
nand UO_434 (O_434,N_4900,N_4961);
and UO_435 (O_435,N_4942,N_4963);
and UO_436 (O_436,N_4981,N_4929);
or UO_437 (O_437,N_4916,N_4923);
nor UO_438 (O_438,N_4962,N_4971);
and UO_439 (O_439,N_4925,N_4907);
or UO_440 (O_440,N_4981,N_4945);
nand UO_441 (O_441,N_4951,N_4940);
nor UO_442 (O_442,N_4918,N_4944);
and UO_443 (O_443,N_4965,N_4922);
nor UO_444 (O_444,N_4985,N_4935);
or UO_445 (O_445,N_4965,N_4994);
nand UO_446 (O_446,N_4940,N_4931);
xor UO_447 (O_447,N_4987,N_4927);
nand UO_448 (O_448,N_4973,N_4971);
nand UO_449 (O_449,N_4984,N_4902);
nand UO_450 (O_450,N_4920,N_4991);
nor UO_451 (O_451,N_4965,N_4974);
or UO_452 (O_452,N_4939,N_4910);
nor UO_453 (O_453,N_4994,N_4963);
and UO_454 (O_454,N_4941,N_4993);
nand UO_455 (O_455,N_4904,N_4971);
nand UO_456 (O_456,N_4906,N_4918);
nand UO_457 (O_457,N_4946,N_4956);
nor UO_458 (O_458,N_4927,N_4940);
nor UO_459 (O_459,N_4993,N_4933);
and UO_460 (O_460,N_4999,N_4969);
and UO_461 (O_461,N_4950,N_4945);
and UO_462 (O_462,N_4933,N_4911);
and UO_463 (O_463,N_4901,N_4970);
and UO_464 (O_464,N_4945,N_4944);
or UO_465 (O_465,N_4955,N_4903);
and UO_466 (O_466,N_4987,N_4951);
or UO_467 (O_467,N_4908,N_4923);
nand UO_468 (O_468,N_4962,N_4937);
nand UO_469 (O_469,N_4982,N_4988);
nand UO_470 (O_470,N_4951,N_4914);
nand UO_471 (O_471,N_4970,N_4945);
xor UO_472 (O_472,N_4991,N_4995);
or UO_473 (O_473,N_4944,N_4973);
and UO_474 (O_474,N_4953,N_4982);
or UO_475 (O_475,N_4983,N_4967);
or UO_476 (O_476,N_4932,N_4991);
and UO_477 (O_477,N_4926,N_4903);
nor UO_478 (O_478,N_4977,N_4948);
and UO_479 (O_479,N_4962,N_4904);
or UO_480 (O_480,N_4999,N_4931);
nand UO_481 (O_481,N_4929,N_4907);
nor UO_482 (O_482,N_4909,N_4919);
and UO_483 (O_483,N_4923,N_4971);
nor UO_484 (O_484,N_4936,N_4953);
or UO_485 (O_485,N_4993,N_4992);
or UO_486 (O_486,N_4921,N_4993);
or UO_487 (O_487,N_4924,N_4925);
and UO_488 (O_488,N_4959,N_4960);
and UO_489 (O_489,N_4934,N_4972);
or UO_490 (O_490,N_4993,N_4926);
nand UO_491 (O_491,N_4908,N_4940);
or UO_492 (O_492,N_4907,N_4946);
nor UO_493 (O_493,N_4925,N_4929);
nand UO_494 (O_494,N_4902,N_4991);
nor UO_495 (O_495,N_4938,N_4900);
and UO_496 (O_496,N_4975,N_4958);
and UO_497 (O_497,N_4972,N_4947);
and UO_498 (O_498,N_4959,N_4930);
or UO_499 (O_499,N_4919,N_4999);
and UO_500 (O_500,N_4986,N_4908);
nor UO_501 (O_501,N_4997,N_4943);
and UO_502 (O_502,N_4967,N_4986);
or UO_503 (O_503,N_4919,N_4938);
and UO_504 (O_504,N_4909,N_4964);
nor UO_505 (O_505,N_4942,N_4973);
nand UO_506 (O_506,N_4939,N_4962);
or UO_507 (O_507,N_4956,N_4982);
or UO_508 (O_508,N_4949,N_4905);
nor UO_509 (O_509,N_4955,N_4921);
nand UO_510 (O_510,N_4975,N_4969);
or UO_511 (O_511,N_4978,N_4932);
nor UO_512 (O_512,N_4978,N_4984);
nand UO_513 (O_513,N_4994,N_4961);
nand UO_514 (O_514,N_4973,N_4960);
and UO_515 (O_515,N_4960,N_4971);
nor UO_516 (O_516,N_4907,N_4965);
nand UO_517 (O_517,N_4900,N_4911);
nand UO_518 (O_518,N_4953,N_4971);
xnor UO_519 (O_519,N_4999,N_4985);
and UO_520 (O_520,N_4981,N_4975);
and UO_521 (O_521,N_4996,N_4924);
nor UO_522 (O_522,N_4916,N_4949);
or UO_523 (O_523,N_4973,N_4949);
or UO_524 (O_524,N_4922,N_4980);
and UO_525 (O_525,N_4974,N_4901);
nor UO_526 (O_526,N_4996,N_4988);
and UO_527 (O_527,N_4957,N_4960);
nand UO_528 (O_528,N_4935,N_4932);
nand UO_529 (O_529,N_4932,N_4982);
nand UO_530 (O_530,N_4929,N_4949);
and UO_531 (O_531,N_4929,N_4916);
nand UO_532 (O_532,N_4969,N_4910);
nand UO_533 (O_533,N_4963,N_4935);
nor UO_534 (O_534,N_4991,N_4944);
nand UO_535 (O_535,N_4928,N_4935);
nand UO_536 (O_536,N_4911,N_4949);
or UO_537 (O_537,N_4980,N_4924);
nor UO_538 (O_538,N_4984,N_4938);
nand UO_539 (O_539,N_4979,N_4955);
or UO_540 (O_540,N_4999,N_4982);
or UO_541 (O_541,N_4918,N_4911);
nand UO_542 (O_542,N_4942,N_4984);
or UO_543 (O_543,N_4958,N_4912);
nand UO_544 (O_544,N_4913,N_4976);
or UO_545 (O_545,N_4971,N_4985);
and UO_546 (O_546,N_4941,N_4955);
xnor UO_547 (O_547,N_4916,N_4907);
nand UO_548 (O_548,N_4955,N_4970);
nand UO_549 (O_549,N_4970,N_4921);
or UO_550 (O_550,N_4958,N_4931);
nand UO_551 (O_551,N_4951,N_4956);
nand UO_552 (O_552,N_4916,N_4980);
and UO_553 (O_553,N_4947,N_4951);
nor UO_554 (O_554,N_4912,N_4957);
or UO_555 (O_555,N_4937,N_4954);
and UO_556 (O_556,N_4970,N_4940);
nand UO_557 (O_557,N_4995,N_4922);
nor UO_558 (O_558,N_4935,N_4905);
or UO_559 (O_559,N_4918,N_4960);
nand UO_560 (O_560,N_4943,N_4998);
nor UO_561 (O_561,N_4999,N_4945);
and UO_562 (O_562,N_4957,N_4987);
or UO_563 (O_563,N_4970,N_4972);
or UO_564 (O_564,N_4906,N_4982);
nor UO_565 (O_565,N_4943,N_4978);
nor UO_566 (O_566,N_4921,N_4915);
or UO_567 (O_567,N_4958,N_4935);
and UO_568 (O_568,N_4932,N_4997);
and UO_569 (O_569,N_4931,N_4946);
or UO_570 (O_570,N_4932,N_4945);
nand UO_571 (O_571,N_4960,N_4910);
nor UO_572 (O_572,N_4988,N_4916);
or UO_573 (O_573,N_4900,N_4965);
nor UO_574 (O_574,N_4913,N_4932);
nand UO_575 (O_575,N_4919,N_4995);
nor UO_576 (O_576,N_4949,N_4956);
nor UO_577 (O_577,N_4929,N_4951);
or UO_578 (O_578,N_4981,N_4991);
nor UO_579 (O_579,N_4942,N_4972);
nor UO_580 (O_580,N_4916,N_4933);
nand UO_581 (O_581,N_4934,N_4912);
xor UO_582 (O_582,N_4951,N_4954);
and UO_583 (O_583,N_4972,N_4988);
and UO_584 (O_584,N_4929,N_4903);
or UO_585 (O_585,N_4958,N_4927);
and UO_586 (O_586,N_4969,N_4965);
and UO_587 (O_587,N_4942,N_4938);
nor UO_588 (O_588,N_4995,N_4929);
and UO_589 (O_589,N_4908,N_4944);
and UO_590 (O_590,N_4916,N_4977);
nand UO_591 (O_591,N_4902,N_4909);
nor UO_592 (O_592,N_4923,N_4979);
and UO_593 (O_593,N_4916,N_4918);
and UO_594 (O_594,N_4981,N_4978);
or UO_595 (O_595,N_4956,N_4919);
nor UO_596 (O_596,N_4962,N_4922);
nand UO_597 (O_597,N_4974,N_4977);
and UO_598 (O_598,N_4992,N_4957);
nor UO_599 (O_599,N_4925,N_4931);
nand UO_600 (O_600,N_4938,N_4960);
nor UO_601 (O_601,N_4975,N_4961);
and UO_602 (O_602,N_4902,N_4974);
and UO_603 (O_603,N_4978,N_4983);
and UO_604 (O_604,N_4942,N_4993);
and UO_605 (O_605,N_4980,N_4971);
or UO_606 (O_606,N_4956,N_4997);
and UO_607 (O_607,N_4901,N_4992);
and UO_608 (O_608,N_4946,N_4916);
and UO_609 (O_609,N_4934,N_4921);
nand UO_610 (O_610,N_4997,N_4952);
nand UO_611 (O_611,N_4906,N_4917);
or UO_612 (O_612,N_4995,N_4985);
nand UO_613 (O_613,N_4970,N_4911);
nand UO_614 (O_614,N_4940,N_4914);
or UO_615 (O_615,N_4993,N_4961);
xor UO_616 (O_616,N_4912,N_4975);
nand UO_617 (O_617,N_4960,N_4958);
and UO_618 (O_618,N_4975,N_4955);
nor UO_619 (O_619,N_4925,N_4916);
nor UO_620 (O_620,N_4913,N_4960);
nand UO_621 (O_621,N_4990,N_4991);
and UO_622 (O_622,N_4986,N_4940);
or UO_623 (O_623,N_4904,N_4920);
nor UO_624 (O_624,N_4959,N_4999);
nor UO_625 (O_625,N_4921,N_4912);
and UO_626 (O_626,N_4923,N_4910);
and UO_627 (O_627,N_4959,N_4914);
or UO_628 (O_628,N_4924,N_4926);
nand UO_629 (O_629,N_4946,N_4912);
or UO_630 (O_630,N_4921,N_4979);
nor UO_631 (O_631,N_4919,N_4992);
and UO_632 (O_632,N_4969,N_4980);
or UO_633 (O_633,N_4981,N_4906);
and UO_634 (O_634,N_4964,N_4943);
xnor UO_635 (O_635,N_4918,N_4968);
nor UO_636 (O_636,N_4910,N_4921);
and UO_637 (O_637,N_4904,N_4908);
nor UO_638 (O_638,N_4910,N_4911);
nor UO_639 (O_639,N_4937,N_4909);
nor UO_640 (O_640,N_4950,N_4989);
nor UO_641 (O_641,N_4922,N_4933);
and UO_642 (O_642,N_4948,N_4934);
or UO_643 (O_643,N_4937,N_4989);
nor UO_644 (O_644,N_4905,N_4914);
nor UO_645 (O_645,N_4912,N_4940);
nor UO_646 (O_646,N_4947,N_4993);
or UO_647 (O_647,N_4985,N_4943);
nand UO_648 (O_648,N_4948,N_4983);
or UO_649 (O_649,N_4958,N_4968);
nand UO_650 (O_650,N_4964,N_4928);
and UO_651 (O_651,N_4963,N_4919);
nand UO_652 (O_652,N_4908,N_4938);
nor UO_653 (O_653,N_4914,N_4971);
nand UO_654 (O_654,N_4981,N_4938);
nor UO_655 (O_655,N_4971,N_4982);
nor UO_656 (O_656,N_4992,N_4906);
and UO_657 (O_657,N_4977,N_4954);
and UO_658 (O_658,N_4946,N_4971);
xnor UO_659 (O_659,N_4901,N_4945);
and UO_660 (O_660,N_4901,N_4989);
and UO_661 (O_661,N_4931,N_4955);
or UO_662 (O_662,N_4981,N_4986);
or UO_663 (O_663,N_4975,N_4992);
and UO_664 (O_664,N_4909,N_4923);
or UO_665 (O_665,N_4953,N_4950);
and UO_666 (O_666,N_4929,N_4986);
or UO_667 (O_667,N_4946,N_4977);
and UO_668 (O_668,N_4996,N_4921);
nand UO_669 (O_669,N_4997,N_4970);
and UO_670 (O_670,N_4972,N_4940);
and UO_671 (O_671,N_4911,N_4994);
or UO_672 (O_672,N_4952,N_4935);
and UO_673 (O_673,N_4910,N_4958);
and UO_674 (O_674,N_4959,N_4954);
nor UO_675 (O_675,N_4993,N_4955);
and UO_676 (O_676,N_4932,N_4969);
xnor UO_677 (O_677,N_4982,N_4965);
and UO_678 (O_678,N_4910,N_4957);
or UO_679 (O_679,N_4914,N_4995);
and UO_680 (O_680,N_4976,N_4934);
and UO_681 (O_681,N_4953,N_4903);
and UO_682 (O_682,N_4913,N_4968);
nor UO_683 (O_683,N_4914,N_4989);
xor UO_684 (O_684,N_4993,N_4948);
and UO_685 (O_685,N_4942,N_4921);
nor UO_686 (O_686,N_4944,N_4998);
nand UO_687 (O_687,N_4917,N_4904);
and UO_688 (O_688,N_4939,N_4947);
or UO_689 (O_689,N_4981,N_4947);
nor UO_690 (O_690,N_4949,N_4922);
or UO_691 (O_691,N_4956,N_4917);
and UO_692 (O_692,N_4964,N_4937);
nor UO_693 (O_693,N_4910,N_4987);
or UO_694 (O_694,N_4991,N_4952);
or UO_695 (O_695,N_4931,N_4973);
nor UO_696 (O_696,N_4991,N_4972);
nor UO_697 (O_697,N_4986,N_4965);
nand UO_698 (O_698,N_4956,N_4931);
or UO_699 (O_699,N_4913,N_4987);
nand UO_700 (O_700,N_4988,N_4976);
or UO_701 (O_701,N_4954,N_4909);
or UO_702 (O_702,N_4987,N_4903);
or UO_703 (O_703,N_4990,N_4939);
nor UO_704 (O_704,N_4973,N_4919);
or UO_705 (O_705,N_4972,N_4922);
or UO_706 (O_706,N_4905,N_4915);
nor UO_707 (O_707,N_4998,N_4959);
nor UO_708 (O_708,N_4950,N_4935);
and UO_709 (O_709,N_4992,N_4952);
nand UO_710 (O_710,N_4982,N_4912);
nor UO_711 (O_711,N_4943,N_4933);
or UO_712 (O_712,N_4980,N_4918);
nor UO_713 (O_713,N_4964,N_4932);
nand UO_714 (O_714,N_4949,N_4924);
and UO_715 (O_715,N_4961,N_4944);
nor UO_716 (O_716,N_4992,N_4976);
nand UO_717 (O_717,N_4935,N_4984);
nand UO_718 (O_718,N_4960,N_4962);
nor UO_719 (O_719,N_4912,N_4939);
nor UO_720 (O_720,N_4972,N_4958);
and UO_721 (O_721,N_4953,N_4958);
nand UO_722 (O_722,N_4939,N_4955);
and UO_723 (O_723,N_4937,N_4917);
or UO_724 (O_724,N_4992,N_4947);
and UO_725 (O_725,N_4947,N_4908);
xor UO_726 (O_726,N_4951,N_4990);
and UO_727 (O_727,N_4906,N_4977);
nor UO_728 (O_728,N_4909,N_4969);
and UO_729 (O_729,N_4929,N_4964);
or UO_730 (O_730,N_4990,N_4959);
nand UO_731 (O_731,N_4940,N_4919);
nor UO_732 (O_732,N_4954,N_4945);
nand UO_733 (O_733,N_4953,N_4992);
nand UO_734 (O_734,N_4970,N_4969);
nand UO_735 (O_735,N_4999,N_4915);
nor UO_736 (O_736,N_4958,N_4936);
nor UO_737 (O_737,N_4972,N_4949);
nor UO_738 (O_738,N_4903,N_4905);
and UO_739 (O_739,N_4972,N_4948);
nor UO_740 (O_740,N_4955,N_4958);
nor UO_741 (O_741,N_4933,N_4991);
nand UO_742 (O_742,N_4991,N_4993);
or UO_743 (O_743,N_4972,N_4929);
nor UO_744 (O_744,N_4966,N_4980);
or UO_745 (O_745,N_4995,N_4945);
nand UO_746 (O_746,N_4901,N_4990);
and UO_747 (O_747,N_4925,N_4964);
and UO_748 (O_748,N_4934,N_4963);
nand UO_749 (O_749,N_4998,N_4911);
nand UO_750 (O_750,N_4923,N_4920);
nor UO_751 (O_751,N_4985,N_4956);
and UO_752 (O_752,N_4979,N_4970);
or UO_753 (O_753,N_4935,N_4989);
nand UO_754 (O_754,N_4960,N_4901);
nor UO_755 (O_755,N_4920,N_4916);
or UO_756 (O_756,N_4963,N_4964);
xor UO_757 (O_757,N_4931,N_4987);
or UO_758 (O_758,N_4915,N_4987);
nor UO_759 (O_759,N_4989,N_4987);
xnor UO_760 (O_760,N_4935,N_4906);
nand UO_761 (O_761,N_4946,N_4978);
and UO_762 (O_762,N_4952,N_4947);
or UO_763 (O_763,N_4992,N_4936);
nor UO_764 (O_764,N_4980,N_4928);
and UO_765 (O_765,N_4906,N_4941);
nand UO_766 (O_766,N_4927,N_4902);
and UO_767 (O_767,N_4938,N_4925);
and UO_768 (O_768,N_4928,N_4925);
or UO_769 (O_769,N_4966,N_4963);
nand UO_770 (O_770,N_4948,N_4969);
nor UO_771 (O_771,N_4973,N_4987);
nand UO_772 (O_772,N_4998,N_4995);
nor UO_773 (O_773,N_4972,N_4909);
or UO_774 (O_774,N_4921,N_4954);
xnor UO_775 (O_775,N_4916,N_4945);
and UO_776 (O_776,N_4958,N_4966);
and UO_777 (O_777,N_4909,N_4932);
and UO_778 (O_778,N_4948,N_4911);
or UO_779 (O_779,N_4933,N_4957);
or UO_780 (O_780,N_4966,N_4912);
nand UO_781 (O_781,N_4913,N_4955);
and UO_782 (O_782,N_4907,N_4963);
and UO_783 (O_783,N_4980,N_4961);
and UO_784 (O_784,N_4919,N_4952);
or UO_785 (O_785,N_4967,N_4902);
nor UO_786 (O_786,N_4987,N_4986);
nor UO_787 (O_787,N_4916,N_4963);
nor UO_788 (O_788,N_4937,N_4906);
or UO_789 (O_789,N_4939,N_4982);
nor UO_790 (O_790,N_4928,N_4962);
and UO_791 (O_791,N_4918,N_4927);
and UO_792 (O_792,N_4956,N_4969);
nor UO_793 (O_793,N_4988,N_4981);
nor UO_794 (O_794,N_4976,N_4954);
nor UO_795 (O_795,N_4945,N_4949);
nor UO_796 (O_796,N_4971,N_4931);
nand UO_797 (O_797,N_4909,N_4955);
or UO_798 (O_798,N_4958,N_4911);
nand UO_799 (O_799,N_4909,N_4900);
and UO_800 (O_800,N_4991,N_4930);
and UO_801 (O_801,N_4998,N_4967);
nand UO_802 (O_802,N_4918,N_4948);
nor UO_803 (O_803,N_4954,N_4906);
or UO_804 (O_804,N_4994,N_4996);
nor UO_805 (O_805,N_4985,N_4955);
or UO_806 (O_806,N_4905,N_4916);
nor UO_807 (O_807,N_4967,N_4936);
and UO_808 (O_808,N_4956,N_4968);
and UO_809 (O_809,N_4913,N_4959);
or UO_810 (O_810,N_4934,N_4956);
nor UO_811 (O_811,N_4915,N_4904);
or UO_812 (O_812,N_4985,N_4957);
xnor UO_813 (O_813,N_4965,N_4931);
or UO_814 (O_814,N_4954,N_4985);
and UO_815 (O_815,N_4956,N_4983);
nand UO_816 (O_816,N_4986,N_4901);
nand UO_817 (O_817,N_4913,N_4943);
nor UO_818 (O_818,N_4956,N_4909);
nor UO_819 (O_819,N_4926,N_4946);
or UO_820 (O_820,N_4990,N_4976);
or UO_821 (O_821,N_4928,N_4916);
and UO_822 (O_822,N_4917,N_4927);
or UO_823 (O_823,N_4953,N_4999);
nand UO_824 (O_824,N_4934,N_4918);
nor UO_825 (O_825,N_4943,N_4972);
nor UO_826 (O_826,N_4953,N_4942);
nor UO_827 (O_827,N_4951,N_4958);
nor UO_828 (O_828,N_4954,N_4955);
or UO_829 (O_829,N_4950,N_4997);
nor UO_830 (O_830,N_4980,N_4987);
xor UO_831 (O_831,N_4937,N_4923);
or UO_832 (O_832,N_4993,N_4978);
and UO_833 (O_833,N_4951,N_4999);
and UO_834 (O_834,N_4981,N_4973);
and UO_835 (O_835,N_4971,N_4939);
or UO_836 (O_836,N_4980,N_4965);
nor UO_837 (O_837,N_4940,N_4955);
and UO_838 (O_838,N_4913,N_4996);
nor UO_839 (O_839,N_4922,N_4903);
or UO_840 (O_840,N_4964,N_4927);
nor UO_841 (O_841,N_4982,N_4902);
and UO_842 (O_842,N_4985,N_4977);
nand UO_843 (O_843,N_4950,N_4927);
and UO_844 (O_844,N_4967,N_4950);
or UO_845 (O_845,N_4944,N_4982);
nor UO_846 (O_846,N_4910,N_4997);
nor UO_847 (O_847,N_4975,N_4966);
nand UO_848 (O_848,N_4914,N_4912);
and UO_849 (O_849,N_4959,N_4952);
or UO_850 (O_850,N_4919,N_4990);
nor UO_851 (O_851,N_4966,N_4919);
xor UO_852 (O_852,N_4900,N_4922);
nand UO_853 (O_853,N_4954,N_4981);
and UO_854 (O_854,N_4911,N_4950);
and UO_855 (O_855,N_4976,N_4915);
or UO_856 (O_856,N_4942,N_4991);
xnor UO_857 (O_857,N_4920,N_4921);
nand UO_858 (O_858,N_4935,N_4903);
nand UO_859 (O_859,N_4963,N_4928);
nand UO_860 (O_860,N_4900,N_4972);
nor UO_861 (O_861,N_4987,N_4936);
nand UO_862 (O_862,N_4963,N_4985);
xnor UO_863 (O_863,N_4973,N_4976);
and UO_864 (O_864,N_4992,N_4912);
and UO_865 (O_865,N_4989,N_4977);
and UO_866 (O_866,N_4942,N_4913);
nor UO_867 (O_867,N_4939,N_4916);
nor UO_868 (O_868,N_4962,N_4963);
or UO_869 (O_869,N_4910,N_4950);
nand UO_870 (O_870,N_4974,N_4920);
nand UO_871 (O_871,N_4966,N_4939);
or UO_872 (O_872,N_4943,N_4973);
and UO_873 (O_873,N_4998,N_4960);
nand UO_874 (O_874,N_4995,N_4924);
nand UO_875 (O_875,N_4986,N_4914);
nand UO_876 (O_876,N_4900,N_4970);
and UO_877 (O_877,N_4993,N_4935);
nor UO_878 (O_878,N_4936,N_4979);
nand UO_879 (O_879,N_4940,N_4969);
and UO_880 (O_880,N_4920,N_4953);
or UO_881 (O_881,N_4940,N_4963);
or UO_882 (O_882,N_4906,N_4983);
and UO_883 (O_883,N_4936,N_4980);
nor UO_884 (O_884,N_4922,N_4937);
nor UO_885 (O_885,N_4988,N_4921);
and UO_886 (O_886,N_4956,N_4965);
nand UO_887 (O_887,N_4983,N_4913);
nor UO_888 (O_888,N_4923,N_4936);
or UO_889 (O_889,N_4918,N_4963);
nand UO_890 (O_890,N_4963,N_4993);
and UO_891 (O_891,N_4911,N_4902);
nand UO_892 (O_892,N_4921,N_4977);
nand UO_893 (O_893,N_4970,N_4930);
and UO_894 (O_894,N_4906,N_4938);
nor UO_895 (O_895,N_4974,N_4961);
nor UO_896 (O_896,N_4997,N_4983);
nor UO_897 (O_897,N_4967,N_4912);
nor UO_898 (O_898,N_4977,N_4938);
nand UO_899 (O_899,N_4985,N_4987);
or UO_900 (O_900,N_4926,N_4936);
nand UO_901 (O_901,N_4987,N_4923);
nand UO_902 (O_902,N_4970,N_4960);
and UO_903 (O_903,N_4948,N_4921);
nand UO_904 (O_904,N_4958,N_4907);
and UO_905 (O_905,N_4991,N_4913);
nand UO_906 (O_906,N_4924,N_4946);
and UO_907 (O_907,N_4953,N_4996);
and UO_908 (O_908,N_4960,N_4977);
xor UO_909 (O_909,N_4948,N_4963);
or UO_910 (O_910,N_4923,N_4988);
nand UO_911 (O_911,N_4983,N_4999);
nand UO_912 (O_912,N_4957,N_4911);
or UO_913 (O_913,N_4991,N_4963);
nor UO_914 (O_914,N_4958,N_4970);
nand UO_915 (O_915,N_4991,N_4903);
or UO_916 (O_916,N_4984,N_4941);
nand UO_917 (O_917,N_4993,N_4996);
nand UO_918 (O_918,N_4943,N_4965);
nor UO_919 (O_919,N_4996,N_4941);
nand UO_920 (O_920,N_4920,N_4932);
or UO_921 (O_921,N_4991,N_4982);
nand UO_922 (O_922,N_4976,N_4916);
and UO_923 (O_923,N_4906,N_4930);
and UO_924 (O_924,N_4967,N_4931);
nor UO_925 (O_925,N_4930,N_4946);
nand UO_926 (O_926,N_4930,N_4947);
nand UO_927 (O_927,N_4912,N_4954);
nand UO_928 (O_928,N_4994,N_4929);
and UO_929 (O_929,N_4950,N_4991);
nor UO_930 (O_930,N_4912,N_4916);
and UO_931 (O_931,N_4919,N_4928);
and UO_932 (O_932,N_4941,N_4982);
nor UO_933 (O_933,N_4931,N_4981);
or UO_934 (O_934,N_4978,N_4962);
and UO_935 (O_935,N_4992,N_4905);
nand UO_936 (O_936,N_4946,N_4966);
xor UO_937 (O_937,N_4923,N_4976);
nor UO_938 (O_938,N_4940,N_4923);
nor UO_939 (O_939,N_4959,N_4983);
or UO_940 (O_940,N_4925,N_4923);
nor UO_941 (O_941,N_4994,N_4913);
or UO_942 (O_942,N_4979,N_4957);
and UO_943 (O_943,N_4934,N_4989);
and UO_944 (O_944,N_4975,N_4987);
and UO_945 (O_945,N_4923,N_4900);
and UO_946 (O_946,N_4910,N_4944);
and UO_947 (O_947,N_4916,N_4986);
nor UO_948 (O_948,N_4922,N_4943);
nand UO_949 (O_949,N_4969,N_4954);
nor UO_950 (O_950,N_4972,N_4927);
and UO_951 (O_951,N_4965,N_4906);
xnor UO_952 (O_952,N_4993,N_4966);
and UO_953 (O_953,N_4999,N_4908);
nand UO_954 (O_954,N_4991,N_4945);
or UO_955 (O_955,N_4963,N_4939);
and UO_956 (O_956,N_4911,N_4964);
or UO_957 (O_957,N_4948,N_4938);
or UO_958 (O_958,N_4934,N_4919);
nor UO_959 (O_959,N_4990,N_4981);
and UO_960 (O_960,N_4951,N_4961);
nand UO_961 (O_961,N_4937,N_4957);
nor UO_962 (O_962,N_4976,N_4948);
nor UO_963 (O_963,N_4988,N_4914);
and UO_964 (O_964,N_4962,N_4956);
or UO_965 (O_965,N_4952,N_4930);
nor UO_966 (O_966,N_4954,N_4910);
nor UO_967 (O_967,N_4927,N_4973);
and UO_968 (O_968,N_4965,N_4972);
or UO_969 (O_969,N_4965,N_4911);
nand UO_970 (O_970,N_4923,N_4985);
and UO_971 (O_971,N_4945,N_4917);
or UO_972 (O_972,N_4905,N_4988);
or UO_973 (O_973,N_4908,N_4954);
and UO_974 (O_974,N_4953,N_4987);
nand UO_975 (O_975,N_4977,N_4925);
nor UO_976 (O_976,N_4957,N_4946);
and UO_977 (O_977,N_4979,N_4983);
nand UO_978 (O_978,N_4994,N_4900);
nor UO_979 (O_979,N_4933,N_4977);
nor UO_980 (O_980,N_4963,N_4938);
or UO_981 (O_981,N_4930,N_4961);
nor UO_982 (O_982,N_4956,N_4980);
or UO_983 (O_983,N_4993,N_4971);
nand UO_984 (O_984,N_4920,N_4911);
and UO_985 (O_985,N_4964,N_4997);
nand UO_986 (O_986,N_4956,N_4975);
and UO_987 (O_987,N_4908,N_4962);
nor UO_988 (O_988,N_4945,N_4926);
and UO_989 (O_989,N_4927,N_4941);
and UO_990 (O_990,N_4924,N_4940);
nand UO_991 (O_991,N_4934,N_4925);
and UO_992 (O_992,N_4961,N_4977);
xor UO_993 (O_993,N_4957,N_4917);
and UO_994 (O_994,N_4918,N_4923);
nor UO_995 (O_995,N_4959,N_4969);
nand UO_996 (O_996,N_4995,N_4961);
nor UO_997 (O_997,N_4969,N_4911);
nor UO_998 (O_998,N_4901,N_4915);
and UO_999 (O_999,N_4916,N_4934);
endmodule