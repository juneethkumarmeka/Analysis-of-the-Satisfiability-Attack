module basic_750_5000_1000_50_levels_10xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
or U0 (N_0,In_32,In_573);
nand U1 (N_1,In_211,In_296);
or U2 (N_2,In_234,In_617);
xor U3 (N_3,In_142,In_448);
or U4 (N_4,In_375,In_29);
nor U5 (N_5,In_107,In_416);
nor U6 (N_6,In_614,In_1);
xor U7 (N_7,In_84,In_559);
and U8 (N_8,In_315,In_701);
or U9 (N_9,In_620,In_724);
or U10 (N_10,In_399,In_449);
or U11 (N_11,In_447,In_453);
xor U12 (N_12,In_450,In_38);
and U13 (N_13,In_293,In_540);
nor U14 (N_14,In_340,In_597);
nor U15 (N_15,In_305,In_100);
nor U16 (N_16,In_477,In_121);
nand U17 (N_17,In_420,In_373);
nand U18 (N_18,In_455,In_680);
nor U19 (N_19,In_630,In_226);
xor U20 (N_20,In_446,In_529);
xnor U21 (N_21,In_213,In_516);
nand U22 (N_22,In_564,In_596);
xor U23 (N_23,In_370,In_642);
or U24 (N_24,In_191,In_321);
and U25 (N_25,In_451,In_598);
or U26 (N_26,In_671,In_35);
xnor U27 (N_27,In_616,In_587);
or U28 (N_28,In_716,In_282);
nand U29 (N_29,In_688,In_271);
or U30 (N_30,In_437,In_498);
and U31 (N_31,In_524,In_388);
nand U32 (N_32,In_552,In_394);
nor U33 (N_33,In_436,In_183);
nor U34 (N_34,In_155,In_23);
and U35 (N_35,In_555,In_6);
nor U36 (N_36,In_212,In_503);
nor U37 (N_37,In_472,In_55);
xor U38 (N_38,In_415,In_104);
xor U39 (N_39,In_297,In_138);
nor U40 (N_40,In_53,In_641);
or U41 (N_41,In_274,In_194);
xor U42 (N_42,In_623,In_433);
or U43 (N_43,In_726,In_576);
or U44 (N_44,In_290,In_160);
nand U45 (N_45,In_329,In_300);
and U46 (N_46,In_563,In_273);
nand U47 (N_47,In_568,In_124);
and U48 (N_48,In_203,In_607);
nand U49 (N_49,In_389,In_270);
and U50 (N_50,In_77,In_34);
and U51 (N_51,In_75,In_214);
or U52 (N_52,In_640,In_654);
nor U53 (N_53,In_462,In_380);
or U54 (N_54,In_600,In_391);
nand U55 (N_55,In_217,In_426);
or U56 (N_56,In_429,In_515);
or U57 (N_57,In_200,In_737);
or U58 (N_58,In_506,In_99);
nor U59 (N_59,In_149,In_268);
xnor U60 (N_60,In_281,In_513);
xnor U61 (N_61,In_255,In_180);
xor U62 (N_62,In_624,In_478);
or U63 (N_63,In_626,In_357);
nor U64 (N_64,In_311,In_510);
nor U65 (N_65,In_280,In_66);
nor U66 (N_66,In_250,In_251);
or U67 (N_67,In_424,In_589);
and U68 (N_68,In_692,In_725);
xor U69 (N_69,In_245,In_502);
nor U70 (N_70,In_523,In_122);
or U71 (N_71,In_7,In_405);
nand U72 (N_72,In_26,In_358);
or U73 (N_73,In_661,In_728);
xnor U74 (N_74,In_537,In_699);
nor U75 (N_75,In_491,In_461);
and U76 (N_76,In_583,In_153);
and U77 (N_77,In_417,In_238);
xor U78 (N_78,In_743,In_209);
xor U79 (N_79,In_590,In_474);
xor U80 (N_80,In_714,In_495);
or U81 (N_81,In_60,In_628);
or U82 (N_82,In_56,In_143);
nand U83 (N_83,In_223,In_276);
nand U84 (N_84,In_658,In_93);
nor U85 (N_85,In_560,In_289);
nor U86 (N_86,In_79,In_619);
and U87 (N_87,In_158,In_704);
nor U88 (N_88,In_186,In_298);
and U89 (N_89,In_507,In_468);
nand U90 (N_90,In_229,In_254);
xnor U91 (N_91,In_685,In_599);
nand U92 (N_92,In_98,In_567);
and U93 (N_93,In_206,In_356);
nand U94 (N_94,In_132,In_427);
nand U95 (N_95,In_224,In_662);
xnor U96 (N_96,In_593,In_65);
or U97 (N_97,In_412,In_479);
and U98 (N_98,In_738,In_54);
and U99 (N_99,In_5,In_177);
and U100 (N_100,In_525,In_185);
xnor U101 (N_101,N_68,In_249);
nand U102 (N_102,N_82,In_706);
and U103 (N_103,In_456,In_246);
or U104 (N_104,In_74,In_258);
or U105 (N_105,In_664,N_79);
nor U106 (N_106,In_371,In_639);
nand U107 (N_107,In_444,In_42);
xnor U108 (N_108,In_611,In_409);
and U109 (N_109,In_253,In_591);
and U110 (N_110,N_44,N_20);
nand U111 (N_111,In_168,In_228);
and U112 (N_112,In_361,In_39);
or U113 (N_113,In_328,N_12);
or U114 (N_114,In_196,In_635);
and U115 (N_115,In_128,In_719);
and U116 (N_116,In_647,In_88);
or U117 (N_117,In_667,In_485);
xor U118 (N_118,In_398,In_721);
xnor U119 (N_119,In_291,In_579);
and U120 (N_120,In_154,In_663);
and U121 (N_121,In_202,In_260);
or U122 (N_122,In_126,N_99);
or U123 (N_123,In_172,In_182);
xor U124 (N_124,In_13,In_313);
or U125 (N_125,In_693,N_97);
nand U126 (N_126,In_201,In_316);
and U127 (N_127,In_277,In_494);
nand U128 (N_128,In_720,In_683);
nand U129 (N_129,In_331,In_569);
nor U130 (N_130,N_58,In_670);
or U131 (N_131,In_25,In_225);
or U132 (N_132,In_638,In_592);
or U133 (N_133,In_376,In_164);
or U134 (N_134,In_14,In_92);
or U135 (N_135,In_86,In_476);
or U136 (N_136,In_272,In_404);
or U137 (N_137,In_410,In_395);
xor U138 (N_138,In_78,In_440);
nand U139 (N_139,In_146,In_156);
and U140 (N_140,In_733,N_3);
xnor U141 (N_141,In_570,In_689);
and U142 (N_142,In_551,In_163);
xor U143 (N_143,In_500,In_364);
nand U144 (N_144,In_324,In_95);
nand U145 (N_145,In_428,In_602);
or U146 (N_146,N_50,In_644);
or U147 (N_147,In_730,In_267);
or U148 (N_148,In_369,In_480);
nand U149 (N_149,In_216,N_92);
and U150 (N_150,In_11,In_118);
xor U151 (N_151,In_709,In_505);
xor U152 (N_152,In_94,In_530);
or U153 (N_153,N_29,In_204);
nor U154 (N_154,N_46,N_81);
or U155 (N_155,In_252,In_345);
or U156 (N_156,In_115,In_207);
and U157 (N_157,In_130,N_47);
nor U158 (N_158,In_443,In_80);
or U159 (N_159,In_501,In_463);
nor U160 (N_160,In_423,In_534);
and U161 (N_161,In_59,In_702);
nor U162 (N_162,In_269,In_30);
and U163 (N_163,In_621,In_393);
or U164 (N_164,N_89,N_6);
nor U165 (N_165,In_17,In_601);
nor U166 (N_166,In_317,In_347);
or U167 (N_167,In_656,In_711);
xor U168 (N_168,In_546,In_565);
or U169 (N_169,In_707,In_432);
or U170 (N_170,In_337,In_262);
or U171 (N_171,In_136,In_105);
nor U172 (N_172,In_8,N_0);
xor U173 (N_173,In_16,In_648);
nor U174 (N_174,In_220,In_96);
and U175 (N_175,In_715,In_208);
nor U176 (N_176,In_244,In_594);
nor U177 (N_177,In_586,In_181);
and U178 (N_178,In_27,In_323);
xor U179 (N_179,In_117,In_673);
nor U180 (N_180,In_401,In_520);
nand U181 (N_181,In_40,In_400);
nand U182 (N_182,In_350,In_613);
or U183 (N_183,In_547,In_562);
and U184 (N_184,In_379,In_744);
xor U185 (N_185,In_90,In_64);
nand U186 (N_186,In_218,In_452);
nand U187 (N_187,In_386,In_486);
nand U188 (N_188,In_230,In_346);
xnor U189 (N_189,In_622,N_38);
nor U190 (N_190,In_418,In_381);
and U191 (N_191,In_575,In_694);
and U192 (N_192,In_91,N_37);
nand U193 (N_193,In_745,In_722);
or U194 (N_194,In_10,In_483);
xnor U195 (N_195,In_102,In_384);
xnor U196 (N_196,In_286,N_67);
nor U197 (N_197,N_9,In_669);
nand U198 (N_198,N_14,In_574);
nor U199 (N_199,In_278,In_336);
and U200 (N_200,N_167,In_314);
xor U201 (N_201,In_141,N_106);
nand U202 (N_202,In_604,N_93);
nand U203 (N_203,In_167,In_655);
or U204 (N_204,In_522,In_385);
nor U205 (N_205,In_548,In_33);
nor U206 (N_206,In_261,N_192);
or U207 (N_207,N_62,N_72);
xor U208 (N_208,In_499,N_117);
or U209 (N_209,In_301,N_133);
and U210 (N_210,In_668,In_12);
nand U211 (N_211,In_749,In_741);
xnor U212 (N_212,N_18,In_174);
nor U213 (N_213,In_509,In_43);
nand U214 (N_214,In_512,In_488);
nor U215 (N_215,N_184,In_518);
and U216 (N_216,In_698,In_553);
and U217 (N_217,In_279,In_431);
and U218 (N_218,In_199,N_135);
nor U219 (N_219,In_577,In_731);
or U220 (N_220,In_101,In_554);
xor U221 (N_221,N_178,In_588);
xnor U222 (N_222,In_333,In_434);
xor U223 (N_223,N_124,N_130);
xnor U224 (N_224,In_189,N_179);
and U225 (N_225,In_435,N_143);
xnor U226 (N_226,In_539,In_465);
xnor U227 (N_227,In_705,In_578);
nor U228 (N_228,In_471,In_377);
nand U229 (N_229,N_128,In_89);
and U230 (N_230,In_442,N_150);
nor U231 (N_231,In_292,In_28);
nand U232 (N_232,In_351,In_46);
nor U233 (N_233,N_27,In_58);
and U234 (N_234,In_490,In_325);
and U235 (N_235,N_19,N_51);
nor U236 (N_236,In_354,N_153);
and U237 (N_237,N_34,In_542);
nand U238 (N_238,In_372,N_17);
and U239 (N_239,In_265,In_649);
or U240 (N_240,N_22,In_425);
xor U241 (N_241,In_114,In_533);
nor U242 (N_242,In_20,In_161);
and U243 (N_243,In_627,In_341);
and U244 (N_244,In_367,In_157);
and U245 (N_245,N_108,In_116);
nand U246 (N_246,N_88,In_227);
or U247 (N_247,N_87,In_71);
and U248 (N_248,In_646,N_103);
nand U249 (N_249,In_308,N_199);
or U250 (N_250,N_142,N_4);
nand U251 (N_251,In_166,In_343);
and U252 (N_252,In_454,In_113);
and U253 (N_253,N_90,In_475);
and U254 (N_254,In_295,In_69);
and U255 (N_255,In_580,In_309);
xor U256 (N_256,In_411,In_441);
nand U257 (N_257,N_10,In_684);
and U258 (N_258,In_460,N_115);
nor U259 (N_259,In_481,In_205);
nor U260 (N_260,N_36,In_188);
and U261 (N_261,N_105,N_49);
nor U262 (N_262,In_469,In_275);
nand U263 (N_263,In_430,N_95);
and U264 (N_264,N_112,In_110);
and U265 (N_265,N_66,N_123);
and U266 (N_266,In_243,N_11);
nor U267 (N_267,In_193,N_74);
xor U268 (N_268,In_363,In_61);
and U269 (N_269,N_174,N_45);
nor U270 (N_270,In_727,In_544);
or U271 (N_271,In_657,In_215);
or U272 (N_272,In_184,N_100);
xnor U273 (N_273,In_549,In_402);
xnor U274 (N_274,N_65,In_210);
nand U275 (N_275,N_98,N_116);
xnor U276 (N_276,In_397,In_713);
and U277 (N_277,In_742,In_304);
nand U278 (N_278,N_15,N_160);
or U279 (N_279,N_77,In_68);
and U280 (N_280,In_18,N_94);
xnor U281 (N_281,In_595,In_535);
and U282 (N_282,In_691,N_104);
nor U283 (N_283,In_144,In_165);
xor U284 (N_284,In_242,In_125);
nor U285 (N_285,N_159,In_2);
xor U286 (N_286,In_482,In_335);
and U287 (N_287,In_746,In_152);
nand U288 (N_288,In_414,In_72);
nor U289 (N_289,In_241,In_162);
or U290 (N_290,In_748,In_15);
nor U291 (N_291,In_710,In_190);
xor U292 (N_292,In_349,In_679);
and U293 (N_293,In_637,In_556);
or U294 (N_294,N_109,N_132);
or U295 (N_295,In_545,In_51);
or U296 (N_296,In_632,In_284);
or U297 (N_297,N_31,In_4);
and U298 (N_298,In_303,In_392);
nor U299 (N_299,In_195,In_703);
and U300 (N_300,In_532,In_247);
nor U301 (N_301,In_326,In_729);
and U302 (N_302,N_164,N_261);
and U303 (N_303,N_83,In_52);
nor U304 (N_304,In_21,N_260);
and U305 (N_305,In_359,In_526);
nor U306 (N_306,N_282,N_190);
and U307 (N_307,In_631,In_57);
and U308 (N_308,In_135,N_180);
and U309 (N_309,N_129,N_194);
nor U310 (N_310,N_70,N_292);
or U311 (N_311,N_208,N_231);
nor U312 (N_312,In_82,In_368);
nand U313 (N_313,N_225,In_633);
xnor U314 (N_314,N_23,N_176);
or U315 (N_315,In_173,In_259);
xor U316 (N_316,N_134,N_157);
or U317 (N_317,N_131,In_151);
nor U318 (N_318,In_634,N_212);
or U319 (N_319,In_263,In_736);
or U320 (N_320,In_717,N_188);
nor U321 (N_321,In_603,In_231);
nor U322 (N_322,N_290,N_195);
and U323 (N_323,In_123,N_113);
or U324 (N_324,In_687,In_362);
xor U325 (N_325,In_383,N_149);
nor U326 (N_326,In_127,N_273);
xnor U327 (N_327,N_266,N_56);
and U328 (N_328,In_170,N_262);
nor U329 (N_329,In_572,N_234);
nor U330 (N_330,N_274,In_718);
and U331 (N_331,In_541,N_86);
xnor U332 (N_332,In_723,In_473);
xor U333 (N_333,In_45,N_288);
xnor U334 (N_334,In_585,In_531);
and U335 (N_335,In_708,N_64);
xor U336 (N_336,N_147,N_218);
xnor U337 (N_337,In_466,N_213);
nor U338 (N_338,N_215,N_28);
and U339 (N_339,N_120,In_73);
nor U340 (N_340,N_110,N_127);
and U341 (N_341,In_651,In_690);
xnor U342 (N_342,In_256,In_83);
nand U343 (N_343,N_59,In_665);
nor U344 (N_344,N_268,N_161);
and U345 (N_345,N_263,N_244);
and U346 (N_346,N_42,In_299);
nor U347 (N_347,In_408,N_295);
and U348 (N_348,N_210,In_62);
nor U349 (N_349,In_171,In_47);
and U350 (N_350,In_322,In_467);
and U351 (N_351,In_396,N_205);
and U352 (N_352,In_103,N_5);
nand U353 (N_353,In_332,N_101);
nor U354 (N_354,In_439,N_223);
and U355 (N_355,N_39,In_111);
or U356 (N_356,In_137,In_240);
nor U357 (N_357,N_73,In_606);
xnor U358 (N_358,N_2,In_248);
or U359 (N_359,N_84,In_85);
xnor U360 (N_360,In_528,In_464);
nand U361 (N_361,N_236,N_33);
and U362 (N_362,In_41,N_237);
nor U363 (N_363,In_22,In_739);
nor U364 (N_364,N_294,In_239);
xor U365 (N_365,In_283,In_527);
xnor U366 (N_366,In_348,N_25);
nand U367 (N_367,N_272,N_126);
or U368 (N_368,In_63,N_214);
xor U369 (N_369,N_201,In_320);
or U370 (N_370,In_686,In_87);
nor U371 (N_371,N_216,N_26);
nor U372 (N_372,In_339,In_285);
nand U373 (N_373,In_31,N_281);
nor U374 (N_374,N_144,In_366);
or U375 (N_375,N_137,N_258);
nand U376 (N_376,N_251,N_253);
nand U377 (N_377,N_43,N_148);
nand U378 (N_378,N_257,N_165);
xor U379 (N_379,N_48,N_299);
nor U380 (N_380,In_197,N_152);
nor U381 (N_381,N_246,In_561);
or U382 (N_382,In_97,N_7);
nand U383 (N_383,N_222,N_166);
nor U384 (N_384,In_330,N_232);
nand U385 (N_385,N_287,In_558);
nor U386 (N_386,In_489,N_21);
nand U387 (N_387,N_259,N_209);
or U388 (N_388,N_114,N_193);
nor U389 (N_389,In_674,N_55);
nor U390 (N_390,N_228,N_170);
and U391 (N_391,N_69,In_378);
xor U392 (N_392,In_131,N_156);
nor U393 (N_393,N_173,In_382);
nor U394 (N_394,N_271,N_284);
nor U395 (N_395,N_252,N_63);
and U396 (N_396,In_612,N_235);
nor U397 (N_397,N_270,In_735);
and U398 (N_398,N_277,In_584);
or U399 (N_399,In_198,N_233);
and U400 (N_400,In_360,N_304);
or U401 (N_401,N_399,In_338);
and U402 (N_402,In_732,N_352);
nor U403 (N_403,N_217,N_76);
nor U404 (N_404,N_322,In_636);
or U405 (N_405,N_35,N_334);
xnor U406 (N_406,N_249,In_438);
xnor U407 (N_407,In_327,N_311);
or U408 (N_408,In_618,In_140);
nand U409 (N_409,In_571,In_49);
and U410 (N_410,In_387,In_581);
nor U411 (N_411,N_187,In_678);
or U412 (N_412,In_0,In_615);
nand U413 (N_413,N_380,In_287);
xor U414 (N_414,In_3,N_151);
xor U415 (N_415,N_360,N_346);
nand U416 (N_416,In_219,N_227);
xor U417 (N_417,N_363,N_296);
nor U418 (N_418,N_40,In_288);
xor U419 (N_419,In_133,N_255);
nand U420 (N_420,In_233,In_294);
or U421 (N_421,N_344,In_352);
or U422 (N_422,In_696,In_179);
nand U423 (N_423,N_310,In_48);
or U424 (N_424,N_265,N_285);
nor U425 (N_425,N_308,In_445);
and U426 (N_426,In_36,In_487);
xnor U427 (N_427,In_237,N_327);
xnor U428 (N_428,N_107,In_610);
nor U429 (N_429,In_413,N_338);
nor U430 (N_430,In_257,In_457);
nand U431 (N_431,N_183,N_138);
nor U432 (N_432,In_521,N_96);
and U433 (N_433,N_136,In_176);
xor U434 (N_434,N_367,N_305);
nor U435 (N_435,N_242,In_307);
nand U436 (N_436,In_355,N_102);
nand U437 (N_437,In_169,N_203);
nor U438 (N_438,In_134,N_378);
and U439 (N_439,N_269,N_189);
nand U440 (N_440,In_106,N_350);
xor U441 (N_441,N_139,N_140);
nor U442 (N_442,In_266,N_181);
xnor U443 (N_443,In_676,N_254);
nand U444 (N_444,In_519,N_278);
nor U445 (N_445,N_13,N_300);
nor U446 (N_446,In_582,In_740);
and U447 (N_447,N_241,N_85);
or U448 (N_448,In_236,In_652);
or U449 (N_449,N_320,In_514);
nor U450 (N_450,N_240,In_310);
nand U451 (N_451,N_366,In_643);
and U452 (N_452,In_543,In_508);
or U453 (N_453,N_307,N_52);
nand U454 (N_454,N_185,N_118);
or U455 (N_455,N_158,N_1);
or U456 (N_456,In_511,In_318);
nor U457 (N_457,In_119,In_609);
nand U458 (N_458,N_335,N_293);
nand U459 (N_459,N_75,N_230);
or U460 (N_460,N_396,N_369);
xor U461 (N_461,In_470,N_286);
nor U462 (N_462,N_313,N_397);
xnor U463 (N_463,N_393,N_154);
nand U464 (N_464,In_422,N_356);
nand U465 (N_465,N_388,N_30);
nand U466 (N_466,N_341,In_459);
or U467 (N_467,N_202,N_331);
nor U468 (N_468,N_111,In_538);
or U469 (N_469,N_191,N_204);
xnor U470 (N_470,N_394,N_351);
nand U471 (N_471,In_566,N_381);
or U472 (N_472,N_383,N_119);
or U473 (N_473,N_386,N_8);
nand U474 (N_474,N_211,N_326);
or U475 (N_475,N_220,N_60);
nand U476 (N_476,N_41,N_186);
nand U477 (N_477,N_389,In_147);
nor U478 (N_478,In_497,N_298);
nand U479 (N_479,In_625,N_343);
nand U480 (N_480,N_221,N_276);
nand U481 (N_481,N_169,N_219);
nor U482 (N_482,N_54,N_16);
nand U483 (N_483,N_332,N_238);
or U484 (N_484,N_328,In_145);
nand U485 (N_485,In_353,In_306);
xor U486 (N_486,N_339,N_355);
nand U487 (N_487,In_19,N_372);
and U488 (N_488,N_376,N_91);
nand U489 (N_489,In_44,N_374);
nand U490 (N_490,N_330,In_557);
or U491 (N_491,In_493,In_653);
xor U492 (N_492,N_71,N_171);
or U493 (N_493,N_61,N_302);
xnor U494 (N_494,N_243,In_517);
or U495 (N_495,N_390,N_168);
or U496 (N_496,In_605,In_24);
or U497 (N_497,N_155,N_317);
and U498 (N_498,N_175,N_125);
nand U499 (N_499,In_550,N_358);
and U500 (N_500,In_302,N_483);
xnor U501 (N_501,In_712,N_489);
nand U502 (N_502,In_697,N_426);
xnor U503 (N_503,In_37,N_370);
nor U504 (N_504,N_479,N_319);
xnor U505 (N_505,N_375,N_451);
nor U506 (N_506,N_438,N_446);
nor U507 (N_507,N_465,N_340);
or U508 (N_508,N_444,N_475);
and U509 (N_509,N_467,N_373);
or U510 (N_510,N_368,N_122);
or U511 (N_511,N_391,N_309);
and U512 (N_512,In_109,N_401);
nand U513 (N_513,N_406,N_454);
nand U514 (N_514,N_78,N_385);
and U515 (N_515,N_414,N_459);
xor U516 (N_516,N_80,In_608);
nor U517 (N_517,N_405,N_472);
or U518 (N_518,N_403,N_456);
and U519 (N_519,In_187,N_353);
nor U520 (N_520,N_432,N_229);
nand U521 (N_521,N_404,In_365);
or U522 (N_522,In_650,In_458);
and U523 (N_523,N_411,N_354);
or U524 (N_524,N_24,N_362);
or U525 (N_525,N_484,In_484);
xnor U526 (N_526,N_172,N_342);
nor U527 (N_527,N_297,N_325);
nor U528 (N_528,In_67,N_424);
or U529 (N_529,N_435,In_232);
and U530 (N_530,In_139,N_392);
or U531 (N_531,In_682,N_466);
nor U532 (N_532,N_141,N_57);
or U533 (N_533,N_224,N_336);
nor U534 (N_534,N_196,N_162);
and U535 (N_535,N_314,N_497);
nor U536 (N_536,N_425,N_267);
nand U537 (N_537,N_464,N_427);
nand U538 (N_538,In_178,N_419);
xor U539 (N_539,In_148,N_488);
xnor U540 (N_540,N_371,N_442);
or U541 (N_541,N_410,N_447);
nand U542 (N_542,In_319,N_333);
or U543 (N_543,N_395,N_279);
and U544 (N_544,N_478,In_129);
nand U545 (N_545,N_471,N_458);
and U546 (N_546,N_486,N_377);
or U547 (N_547,N_347,N_163);
or U548 (N_548,N_441,In_50);
or U549 (N_549,N_32,N_283);
and U550 (N_550,N_206,In_700);
xor U551 (N_551,N_198,N_291);
or U552 (N_552,In_407,N_239);
or U553 (N_553,In_421,N_473);
and U554 (N_554,N_145,N_357);
xor U555 (N_555,N_382,N_321);
or U556 (N_556,N_485,N_431);
xor U557 (N_557,N_430,N_387);
nor U558 (N_558,N_492,In_747);
or U559 (N_559,N_345,N_197);
nor U560 (N_560,N_450,In_120);
nor U561 (N_561,N_318,N_247);
and U562 (N_562,N_449,N_359);
nor U563 (N_563,N_476,N_289);
or U564 (N_564,In_76,In_666);
nor U565 (N_565,N_312,N_248);
nand U566 (N_566,N_280,In_734);
and U567 (N_567,N_453,In_81);
or U568 (N_568,N_412,N_423);
or U569 (N_569,N_461,N_182);
or U570 (N_570,N_480,N_491);
xor U571 (N_571,N_365,N_301);
nor U572 (N_572,N_457,N_413);
or U573 (N_573,In_681,N_256);
xnor U574 (N_574,N_462,N_121);
xnor U575 (N_575,N_460,N_384);
or U576 (N_576,N_337,N_400);
xnor U577 (N_577,N_324,N_398);
and U578 (N_578,N_452,N_146);
and U579 (N_579,In_150,In_159);
nand U580 (N_580,N_379,N_494);
nor U581 (N_581,N_306,N_329);
and U582 (N_582,In_108,In_221);
xnor U583 (N_583,N_436,N_482);
and U584 (N_584,N_364,N_316);
nor U585 (N_585,In_695,N_349);
nor U586 (N_586,In_419,N_417);
nor U587 (N_587,N_470,N_409);
and U588 (N_588,In_9,N_468);
nand U589 (N_589,In_629,In_175);
and U590 (N_590,N_250,N_315);
xnor U591 (N_591,N_498,N_407);
xor U592 (N_592,N_434,N_402);
and U593 (N_593,N_429,N_474);
and U594 (N_594,In_406,N_200);
nor U595 (N_595,N_490,N_487);
nand U596 (N_596,In_312,In_536);
nor U597 (N_597,N_439,N_455);
nand U598 (N_598,N_440,N_408);
or U599 (N_599,In_492,N_348);
xnor U600 (N_600,In_672,N_590);
or U601 (N_601,N_495,In_235);
or U602 (N_602,N_420,In_222);
nor U603 (N_603,N_507,N_526);
nor U604 (N_604,N_568,In_112);
xnor U605 (N_605,N_577,N_561);
nand U606 (N_606,N_443,N_589);
nor U607 (N_607,N_591,N_445);
nor U608 (N_608,N_560,N_481);
xnor U609 (N_609,N_564,N_525);
or U610 (N_610,N_583,N_599);
and U611 (N_611,N_531,N_415);
or U612 (N_612,N_566,N_275);
nor U613 (N_613,N_552,N_584);
nor U614 (N_614,In_645,N_585);
or U615 (N_615,N_565,N_586);
nand U616 (N_616,N_587,N_575);
nand U617 (N_617,N_177,N_523);
nor U618 (N_618,In_675,N_540);
or U619 (N_619,N_594,N_422);
nor U620 (N_620,N_516,N_571);
nor U621 (N_621,N_574,N_539);
or U622 (N_622,N_563,N_535);
or U623 (N_623,N_578,In_70);
and U624 (N_624,N_581,N_264);
and U625 (N_625,N_500,In_334);
and U626 (N_626,N_514,N_506);
or U627 (N_627,N_572,In_504);
nand U628 (N_628,N_521,N_520);
nor U629 (N_629,N_538,N_524);
and U630 (N_630,N_579,N_555);
and U631 (N_631,N_511,N_496);
xor U632 (N_632,N_548,N_510);
or U633 (N_633,N_421,N_509);
nor U634 (N_634,N_553,N_598);
or U635 (N_635,N_501,In_390);
nor U636 (N_636,N_595,In_660);
nor U637 (N_637,N_418,N_515);
or U638 (N_638,N_549,N_536);
nand U639 (N_639,N_559,In_374);
and U640 (N_640,N_508,N_570);
xor U641 (N_641,N_463,N_547);
and U642 (N_642,N_469,N_529);
nor U643 (N_643,N_567,N_544);
nand U644 (N_644,N_597,N_517);
nor U645 (N_645,N_593,N_588);
nor U646 (N_646,N_573,In_264);
and U647 (N_647,N_513,N_533);
nor U648 (N_648,N_502,N_416);
or U649 (N_649,N_527,N_582);
nand U650 (N_650,In_659,N_537);
nor U651 (N_651,N_504,N_528);
xnor U652 (N_652,N_580,N_512);
and U653 (N_653,N_592,N_477);
and U654 (N_654,N_303,N_543);
nand U655 (N_655,N_546,N_207);
xor U656 (N_656,N_551,N_499);
nand U657 (N_657,N_556,N_542);
nand U658 (N_658,N_596,In_344);
nand U659 (N_659,N_437,N_562);
and U660 (N_660,N_519,N_361);
nand U661 (N_661,N_576,N_522);
and U662 (N_662,N_428,In_403);
nor U663 (N_663,N_503,N_53);
nand U664 (N_664,N_569,In_342);
or U665 (N_665,In_192,N_554);
or U666 (N_666,N_530,N_532);
or U667 (N_667,N_493,N_534);
and U668 (N_668,N_518,N_505);
or U669 (N_669,N_550,N_226);
or U670 (N_670,N_433,In_677);
or U671 (N_671,N_541,N_245);
nand U672 (N_672,In_496,N_448);
nand U673 (N_673,N_557,N_545);
nor U674 (N_674,N_558,N_323);
nand U675 (N_675,N_551,N_567);
nor U676 (N_676,N_275,N_564);
or U677 (N_677,N_544,N_512);
or U678 (N_678,N_517,N_587);
nor U679 (N_679,In_192,N_570);
nand U680 (N_680,N_571,N_585);
or U681 (N_681,N_546,N_516);
nand U682 (N_682,N_428,N_576);
and U683 (N_683,N_538,N_421);
xor U684 (N_684,In_390,In_344);
and U685 (N_685,In_645,N_595);
nand U686 (N_686,N_448,In_645);
or U687 (N_687,N_560,N_558);
nor U688 (N_688,In_496,N_499);
xnor U689 (N_689,N_557,N_514);
nor U690 (N_690,N_594,N_569);
nand U691 (N_691,N_496,N_519);
or U692 (N_692,N_587,N_418);
or U693 (N_693,N_559,N_537);
and U694 (N_694,N_526,N_463);
or U695 (N_695,N_592,N_597);
and U696 (N_696,N_590,In_677);
or U697 (N_697,N_593,In_672);
nand U698 (N_698,N_443,N_564);
nand U699 (N_699,N_323,In_403);
xnor U700 (N_700,N_650,N_619);
xnor U701 (N_701,N_630,N_657);
and U702 (N_702,N_661,N_673);
and U703 (N_703,N_683,N_635);
or U704 (N_704,N_666,N_620);
or U705 (N_705,N_684,N_680);
xor U706 (N_706,N_631,N_600);
nor U707 (N_707,N_627,N_669);
or U708 (N_708,N_693,N_668);
and U709 (N_709,N_679,N_678);
nor U710 (N_710,N_639,N_665);
xnor U711 (N_711,N_629,N_646);
nor U712 (N_712,N_653,N_672);
nand U713 (N_713,N_645,N_676);
nor U714 (N_714,N_626,N_663);
and U715 (N_715,N_652,N_697);
and U716 (N_716,N_604,N_698);
nor U717 (N_717,N_617,N_675);
nor U718 (N_718,N_642,N_677);
or U719 (N_719,N_649,N_692);
or U720 (N_720,N_662,N_611);
xnor U721 (N_721,N_644,N_608);
and U722 (N_722,N_637,N_605);
nand U723 (N_723,N_625,N_659);
or U724 (N_724,N_658,N_660);
xnor U725 (N_725,N_602,N_643);
nor U726 (N_726,N_615,N_695);
xnor U727 (N_727,N_628,N_689);
or U728 (N_728,N_682,N_694);
nor U729 (N_729,N_654,N_641);
xnor U730 (N_730,N_656,N_651);
and U731 (N_731,N_696,N_674);
xor U732 (N_732,N_622,N_690);
or U733 (N_733,N_647,N_618);
xnor U734 (N_734,N_670,N_607);
xor U735 (N_735,N_614,N_638);
nor U736 (N_736,N_613,N_621);
or U737 (N_737,N_616,N_606);
or U738 (N_738,N_671,N_664);
nor U739 (N_739,N_603,N_609);
nand U740 (N_740,N_624,N_699);
and U741 (N_741,N_633,N_667);
xnor U742 (N_742,N_612,N_648);
xnor U743 (N_743,N_632,N_623);
and U744 (N_744,N_685,N_655);
nand U745 (N_745,N_610,N_681);
nand U746 (N_746,N_634,N_636);
or U747 (N_747,N_640,N_686);
and U748 (N_748,N_687,N_691);
nor U749 (N_749,N_688,N_601);
or U750 (N_750,N_615,N_694);
nand U751 (N_751,N_678,N_681);
and U752 (N_752,N_674,N_641);
nor U753 (N_753,N_638,N_640);
xnor U754 (N_754,N_685,N_698);
nand U755 (N_755,N_666,N_681);
and U756 (N_756,N_685,N_636);
and U757 (N_757,N_654,N_630);
or U758 (N_758,N_656,N_626);
or U759 (N_759,N_698,N_680);
and U760 (N_760,N_668,N_658);
xor U761 (N_761,N_643,N_661);
nor U762 (N_762,N_644,N_668);
nand U763 (N_763,N_635,N_673);
nand U764 (N_764,N_664,N_629);
nor U765 (N_765,N_667,N_647);
or U766 (N_766,N_642,N_627);
and U767 (N_767,N_642,N_625);
nor U768 (N_768,N_685,N_669);
and U769 (N_769,N_688,N_624);
or U770 (N_770,N_660,N_670);
nand U771 (N_771,N_676,N_652);
and U772 (N_772,N_620,N_668);
nand U773 (N_773,N_621,N_667);
or U774 (N_774,N_689,N_617);
xor U775 (N_775,N_667,N_626);
and U776 (N_776,N_675,N_613);
nor U777 (N_777,N_670,N_688);
nand U778 (N_778,N_617,N_613);
nor U779 (N_779,N_623,N_670);
nand U780 (N_780,N_648,N_697);
nand U781 (N_781,N_676,N_635);
xor U782 (N_782,N_664,N_633);
nand U783 (N_783,N_632,N_690);
nor U784 (N_784,N_633,N_684);
nand U785 (N_785,N_654,N_688);
nand U786 (N_786,N_610,N_643);
xor U787 (N_787,N_674,N_680);
nor U788 (N_788,N_604,N_601);
nor U789 (N_789,N_613,N_673);
xor U790 (N_790,N_616,N_695);
or U791 (N_791,N_659,N_686);
or U792 (N_792,N_652,N_686);
and U793 (N_793,N_650,N_697);
nor U794 (N_794,N_605,N_612);
or U795 (N_795,N_699,N_610);
or U796 (N_796,N_671,N_627);
nor U797 (N_797,N_636,N_669);
nor U798 (N_798,N_666,N_646);
or U799 (N_799,N_697,N_678);
nand U800 (N_800,N_752,N_780);
nand U801 (N_801,N_756,N_707);
nand U802 (N_802,N_773,N_733);
nor U803 (N_803,N_720,N_718);
xor U804 (N_804,N_732,N_777);
or U805 (N_805,N_751,N_791);
or U806 (N_806,N_762,N_783);
nand U807 (N_807,N_750,N_723);
or U808 (N_808,N_743,N_747);
nand U809 (N_809,N_709,N_794);
nand U810 (N_810,N_706,N_782);
xnor U811 (N_811,N_785,N_736);
nand U812 (N_812,N_708,N_767);
or U813 (N_813,N_705,N_768);
nand U814 (N_814,N_769,N_795);
nand U815 (N_815,N_760,N_711);
or U816 (N_816,N_734,N_753);
nor U817 (N_817,N_724,N_740);
nand U818 (N_818,N_717,N_754);
nand U819 (N_819,N_744,N_738);
nor U820 (N_820,N_755,N_786);
nand U821 (N_821,N_742,N_796);
nor U822 (N_822,N_731,N_775);
xnor U823 (N_823,N_797,N_715);
xor U824 (N_824,N_778,N_725);
nor U825 (N_825,N_758,N_764);
nand U826 (N_826,N_766,N_771);
and U827 (N_827,N_722,N_713);
and U828 (N_828,N_799,N_721);
or U829 (N_829,N_714,N_745);
nand U830 (N_830,N_757,N_726);
or U831 (N_831,N_716,N_792);
or U832 (N_832,N_727,N_703);
nand U833 (N_833,N_761,N_788);
or U834 (N_834,N_748,N_710);
nor U835 (N_835,N_793,N_700);
and U836 (N_836,N_776,N_701);
or U837 (N_837,N_739,N_729);
and U838 (N_838,N_774,N_789);
nor U839 (N_839,N_702,N_781);
and U840 (N_840,N_737,N_787);
xor U841 (N_841,N_728,N_730);
nand U842 (N_842,N_712,N_704);
nor U843 (N_843,N_759,N_719);
nor U844 (N_844,N_746,N_735);
xor U845 (N_845,N_772,N_763);
nand U846 (N_846,N_749,N_784);
nor U847 (N_847,N_779,N_770);
nand U848 (N_848,N_765,N_790);
and U849 (N_849,N_741,N_798);
and U850 (N_850,N_798,N_704);
xnor U851 (N_851,N_773,N_743);
nor U852 (N_852,N_715,N_789);
and U853 (N_853,N_761,N_784);
xnor U854 (N_854,N_753,N_754);
or U855 (N_855,N_777,N_746);
and U856 (N_856,N_751,N_757);
or U857 (N_857,N_795,N_782);
or U858 (N_858,N_751,N_755);
nand U859 (N_859,N_793,N_777);
xnor U860 (N_860,N_736,N_787);
nand U861 (N_861,N_748,N_798);
nand U862 (N_862,N_775,N_766);
nand U863 (N_863,N_754,N_736);
nand U864 (N_864,N_703,N_719);
or U865 (N_865,N_758,N_744);
nand U866 (N_866,N_780,N_742);
or U867 (N_867,N_729,N_766);
or U868 (N_868,N_701,N_715);
and U869 (N_869,N_703,N_705);
xnor U870 (N_870,N_780,N_745);
nor U871 (N_871,N_786,N_711);
nor U872 (N_872,N_742,N_708);
xnor U873 (N_873,N_729,N_718);
nor U874 (N_874,N_732,N_771);
or U875 (N_875,N_778,N_739);
nand U876 (N_876,N_780,N_732);
and U877 (N_877,N_780,N_776);
and U878 (N_878,N_740,N_714);
nand U879 (N_879,N_718,N_711);
xor U880 (N_880,N_702,N_765);
nor U881 (N_881,N_723,N_744);
nand U882 (N_882,N_792,N_771);
or U883 (N_883,N_796,N_760);
nor U884 (N_884,N_798,N_797);
xor U885 (N_885,N_710,N_723);
nand U886 (N_886,N_734,N_754);
nor U887 (N_887,N_702,N_703);
nand U888 (N_888,N_777,N_709);
xor U889 (N_889,N_764,N_737);
or U890 (N_890,N_785,N_753);
nand U891 (N_891,N_780,N_715);
and U892 (N_892,N_753,N_752);
and U893 (N_893,N_750,N_756);
xor U894 (N_894,N_769,N_789);
nor U895 (N_895,N_767,N_751);
nor U896 (N_896,N_762,N_718);
nor U897 (N_897,N_786,N_796);
xnor U898 (N_898,N_781,N_740);
and U899 (N_899,N_767,N_762);
nor U900 (N_900,N_867,N_856);
nand U901 (N_901,N_878,N_851);
xor U902 (N_902,N_869,N_807);
or U903 (N_903,N_829,N_859);
or U904 (N_904,N_804,N_892);
nand U905 (N_905,N_899,N_811);
nand U906 (N_906,N_832,N_837);
nand U907 (N_907,N_815,N_805);
nor U908 (N_908,N_884,N_814);
nor U909 (N_909,N_886,N_868);
and U910 (N_910,N_849,N_887);
or U911 (N_911,N_896,N_853);
or U912 (N_912,N_857,N_828);
or U913 (N_913,N_803,N_844);
and U914 (N_914,N_898,N_835);
nor U915 (N_915,N_840,N_838);
and U916 (N_916,N_865,N_860);
nor U917 (N_917,N_891,N_879);
xnor U918 (N_918,N_895,N_827);
nor U919 (N_919,N_877,N_881);
and U920 (N_920,N_862,N_897);
nand U921 (N_921,N_818,N_858);
nand U922 (N_922,N_872,N_809);
or U923 (N_923,N_873,N_801);
or U924 (N_924,N_819,N_883);
and U925 (N_925,N_833,N_816);
or U926 (N_926,N_880,N_817);
or U927 (N_927,N_852,N_864);
nor U928 (N_928,N_810,N_836);
and U929 (N_929,N_893,N_846);
xor U930 (N_930,N_863,N_890);
xor U931 (N_931,N_850,N_802);
and U932 (N_932,N_813,N_888);
xnor U933 (N_933,N_825,N_841);
or U934 (N_934,N_821,N_894);
and U935 (N_935,N_847,N_842);
or U936 (N_936,N_823,N_808);
xnor U937 (N_937,N_812,N_855);
nor U938 (N_938,N_885,N_871);
or U939 (N_939,N_875,N_854);
and U940 (N_940,N_889,N_843);
and U941 (N_941,N_861,N_882);
xor U942 (N_942,N_848,N_806);
xor U943 (N_943,N_824,N_826);
or U944 (N_944,N_876,N_845);
or U945 (N_945,N_870,N_874);
or U946 (N_946,N_834,N_820);
nor U947 (N_947,N_800,N_866);
nor U948 (N_948,N_831,N_839);
and U949 (N_949,N_822,N_830);
nor U950 (N_950,N_834,N_831);
xnor U951 (N_951,N_802,N_855);
xnor U952 (N_952,N_865,N_864);
nand U953 (N_953,N_831,N_893);
nor U954 (N_954,N_830,N_810);
nand U955 (N_955,N_863,N_888);
nor U956 (N_956,N_867,N_801);
and U957 (N_957,N_895,N_821);
nor U958 (N_958,N_897,N_842);
nand U959 (N_959,N_800,N_811);
xnor U960 (N_960,N_812,N_810);
or U961 (N_961,N_884,N_818);
nor U962 (N_962,N_841,N_890);
or U963 (N_963,N_853,N_854);
or U964 (N_964,N_818,N_841);
or U965 (N_965,N_839,N_881);
nor U966 (N_966,N_811,N_847);
nand U967 (N_967,N_827,N_804);
nor U968 (N_968,N_882,N_818);
or U969 (N_969,N_895,N_843);
and U970 (N_970,N_865,N_875);
nor U971 (N_971,N_867,N_837);
nor U972 (N_972,N_888,N_850);
nor U973 (N_973,N_817,N_804);
nor U974 (N_974,N_832,N_891);
xnor U975 (N_975,N_885,N_898);
xnor U976 (N_976,N_806,N_841);
nor U977 (N_977,N_815,N_804);
nor U978 (N_978,N_888,N_865);
and U979 (N_979,N_879,N_810);
nor U980 (N_980,N_813,N_802);
or U981 (N_981,N_808,N_829);
xnor U982 (N_982,N_868,N_837);
nor U983 (N_983,N_845,N_891);
nor U984 (N_984,N_825,N_858);
or U985 (N_985,N_833,N_881);
nor U986 (N_986,N_814,N_862);
and U987 (N_987,N_856,N_817);
and U988 (N_988,N_897,N_894);
xor U989 (N_989,N_811,N_891);
and U990 (N_990,N_885,N_891);
nor U991 (N_991,N_817,N_811);
nor U992 (N_992,N_896,N_891);
and U993 (N_993,N_865,N_898);
and U994 (N_994,N_803,N_845);
nor U995 (N_995,N_816,N_817);
and U996 (N_996,N_890,N_818);
and U997 (N_997,N_869,N_841);
nor U998 (N_998,N_812,N_868);
nor U999 (N_999,N_859,N_822);
and U1000 (N_1000,N_950,N_913);
xnor U1001 (N_1001,N_965,N_989);
nand U1002 (N_1002,N_906,N_933);
or U1003 (N_1003,N_901,N_991);
nand U1004 (N_1004,N_932,N_981);
or U1005 (N_1005,N_928,N_945);
nor U1006 (N_1006,N_948,N_993);
or U1007 (N_1007,N_909,N_942);
xnor U1008 (N_1008,N_935,N_929);
and U1009 (N_1009,N_967,N_927);
nor U1010 (N_1010,N_995,N_934);
nor U1011 (N_1011,N_976,N_940);
or U1012 (N_1012,N_911,N_925);
and U1013 (N_1013,N_919,N_956);
and U1014 (N_1014,N_960,N_990);
and U1015 (N_1015,N_915,N_983);
xnor U1016 (N_1016,N_997,N_984);
and U1017 (N_1017,N_931,N_979);
and U1018 (N_1018,N_996,N_947);
nor U1019 (N_1019,N_994,N_971);
nand U1020 (N_1020,N_985,N_982);
nand U1021 (N_1021,N_914,N_930);
xnor U1022 (N_1022,N_961,N_907);
nor U1023 (N_1023,N_951,N_905);
and U1024 (N_1024,N_910,N_938);
nor U1025 (N_1025,N_972,N_980);
nor U1026 (N_1026,N_949,N_975);
xor U1027 (N_1027,N_968,N_966);
nor U1028 (N_1028,N_921,N_963);
or U1029 (N_1029,N_987,N_957);
xnor U1030 (N_1030,N_977,N_992);
and U1031 (N_1031,N_999,N_953);
nand U1032 (N_1032,N_923,N_926);
or U1033 (N_1033,N_922,N_969);
nand U1034 (N_1034,N_924,N_970);
nor U1035 (N_1035,N_939,N_900);
nor U1036 (N_1036,N_912,N_998);
and U1037 (N_1037,N_903,N_958);
xor U1038 (N_1038,N_941,N_988);
nor U1039 (N_1039,N_973,N_943);
nor U1040 (N_1040,N_902,N_916);
and U1041 (N_1041,N_959,N_978);
or U1042 (N_1042,N_962,N_944);
or U1043 (N_1043,N_946,N_937);
nand U1044 (N_1044,N_974,N_904);
and U1045 (N_1045,N_920,N_908);
nand U1046 (N_1046,N_955,N_918);
nand U1047 (N_1047,N_954,N_917);
or U1048 (N_1048,N_986,N_952);
nor U1049 (N_1049,N_936,N_964);
or U1050 (N_1050,N_922,N_970);
nand U1051 (N_1051,N_911,N_930);
and U1052 (N_1052,N_936,N_915);
nand U1053 (N_1053,N_901,N_988);
nor U1054 (N_1054,N_961,N_970);
nand U1055 (N_1055,N_977,N_944);
or U1056 (N_1056,N_980,N_902);
nor U1057 (N_1057,N_904,N_954);
or U1058 (N_1058,N_917,N_909);
or U1059 (N_1059,N_988,N_989);
or U1060 (N_1060,N_920,N_939);
nand U1061 (N_1061,N_975,N_953);
and U1062 (N_1062,N_900,N_985);
nor U1063 (N_1063,N_987,N_914);
and U1064 (N_1064,N_967,N_963);
nand U1065 (N_1065,N_918,N_913);
nor U1066 (N_1066,N_928,N_921);
and U1067 (N_1067,N_984,N_921);
xor U1068 (N_1068,N_972,N_971);
nor U1069 (N_1069,N_957,N_931);
nor U1070 (N_1070,N_963,N_908);
nor U1071 (N_1071,N_943,N_908);
or U1072 (N_1072,N_995,N_943);
nor U1073 (N_1073,N_926,N_972);
nor U1074 (N_1074,N_999,N_932);
nand U1075 (N_1075,N_923,N_974);
or U1076 (N_1076,N_992,N_915);
nor U1077 (N_1077,N_979,N_976);
and U1078 (N_1078,N_908,N_909);
or U1079 (N_1079,N_908,N_983);
xor U1080 (N_1080,N_969,N_982);
and U1081 (N_1081,N_942,N_930);
or U1082 (N_1082,N_975,N_917);
xor U1083 (N_1083,N_984,N_991);
nand U1084 (N_1084,N_943,N_957);
xor U1085 (N_1085,N_935,N_915);
and U1086 (N_1086,N_942,N_902);
and U1087 (N_1087,N_998,N_927);
nand U1088 (N_1088,N_952,N_964);
nand U1089 (N_1089,N_911,N_939);
nor U1090 (N_1090,N_955,N_965);
and U1091 (N_1091,N_910,N_930);
xnor U1092 (N_1092,N_982,N_994);
nand U1093 (N_1093,N_963,N_988);
nor U1094 (N_1094,N_929,N_988);
and U1095 (N_1095,N_956,N_915);
xor U1096 (N_1096,N_990,N_981);
or U1097 (N_1097,N_920,N_914);
nor U1098 (N_1098,N_908,N_995);
and U1099 (N_1099,N_954,N_965);
and U1100 (N_1100,N_1075,N_1085);
nand U1101 (N_1101,N_1091,N_1052);
and U1102 (N_1102,N_1079,N_1068);
or U1103 (N_1103,N_1096,N_1039);
nor U1104 (N_1104,N_1058,N_1057);
or U1105 (N_1105,N_1086,N_1060);
xor U1106 (N_1106,N_1070,N_1094);
xor U1107 (N_1107,N_1082,N_1099);
xnor U1108 (N_1108,N_1072,N_1069);
or U1109 (N_1109,N_1066,N_1008);
nand U1110 (N_1110,N_1071,N_1064);
and U1111 (N_1111,N_1097,N_1017);
xor U1112 (N_1112,N_1024,N_1005);
nand U1113 (N_1113,N_1003,N_1048);
and U1114 (N_1114,N_1073,N_1049);
and U1115 (N_1115,N_1027,N_1046);
and U1116 (N_1116,N_1083,N_1009);
nor U1117 (N_1117,N_1090,N_1016);
xor U1118 (N_1118,N_1015,N_1004);
nor U1119 (N_1119,N_1010,N_1001);
and U1120 (N_1120,N_1012,N_1040);
and U1121 (N_1121,N_1032,N_1019);
or U1122 (N_1122,N_1030,N_1020);
xor U1123 (N_1123,N_1007,N_1088);
and U1124 (N_1124,N_1098,N_1081);
xor U1125 (N_1125,N_1006,N_1018);
xor U1126 (N_1126,N_1033,N_1053);
or U1127 (N_1127,N_1089,N_1054);
xor U1128 (N_1128,N_1038,N_1036);
or U1129 (N_1129,N_1034,N_1095);
xnor U1130 (N_1130,N_1045,N_1011);
nor U1131 (N_1131,N_1029,N_1031);
nor U1132 (N_1132,N_1067,N_1014);
and U1133 (N_1133,N_1002,N_1021);
nand U1134 (N_1134,N_1065,N_1077);
xor U1135 (N_1135,N_1092,N_1080);
nor U1136 (N_1136,N_1074,N_1047);
nand U1137 (N_1137,N_1055,N_1056);
nand U1138 (N_1138,N_1093,N_1059);
xor U1139 (N_1139,N_1025,N_1044);
nand U1140 (N_1140,N_1043,N_1084);
xor U1141 (N_1141,N_1026,N_1013);
nor U1142 (N_1142,N_1035,N_1078);
xnor U1143 (N_1143,N_1087,N_1062);
nand U1144 (N_1144,N_1023,N_1076);
and U1145 (N_1145,N_1063,N_1061);
nor U1146 (N_1146,N_1041,N_1000);
and U1147 (N_1147,N_1042,N_1050);
or U1148 (N_1148,N_1051,N_1022);
or U1149 (N_1149,N_1037,N_1028);
nor U1150 (N_1150,N_1051,N_1089);
xor U1151 (N_1151,N_1057,N_1070);
nand U1152 (N_1152,N_1027,N_1079);
and U1153 (N_1153,N_1022,N_1041);
and U1154 (N_1154,N_1024,N_1059);
nor U1155 (N_1155,N_1096,N_1098);
nand U1156 (N_1156,N_1071,N_1023);
or U1157 (N_1157,N_1062,N_1022);
xnor U1158 (N_1158,N_1034,N_1059);
xor U1159 (N_1159,N_1092,N_1020);
nor U1160 (N_1160,N_1008,N_1006);
nor U1161 (N_1161,N_1004,N_1076);
and U1162 (N_1162,N_1099,N_1024);
nor U1163 (N_1163,N_1007,N_1065);
nand U1164 (N_1164,N_1047,N_1072);
and U1165 (N_1165,N_1072,N_1079);
nor U1166 (N_1166,N_1087,N_1080);
or U1167 (N_1167,N_1003,N_1088);
and U1168 (N_1168,N_1068,N_1074);
and U1169 (N_1169,N_1079,N_1046);
nor U1170 (N_1170,N_1051,N_1056);
or U1171 (N_1171,N_1083,N_1054);
xnor U1172 (N_1172,N_1017,N_1088);
xnor U1173 (N_1173,N_1065,N_1021);
and U1174 (N_1174,N_1005,N_1017);
nor U1175 (N_1175,N_1082,N_1048);
or U1176 (N_1176,N_1076,N_1044);
nor U1177 (N_1177,N_1046,N_1088);
nand U1178 (N_1178,N_1052,N_1092);
and U1179 (N_1179,N_1005,N_1011);
and U1180 (N_1180,N_1034,N_1079);
or U1181 (N_1181,N_1035,N_1089);
and U1182 (N_1182,N_1052,N_1012);
nor U1183 (N_1183,N_1015,N_1013);
and U1184 (N_1184,N_1056,N_1073);
and U1185 (N_1185,N_1026,N_1011);
xor U1186 (N_1186,N_1096,N_1045);
xnor U1187 (N_1187,N_1045,N_1010);
xor U1188 (N_1188,N_1021,N_1052);
and U1189 (N_1189,N_1064,N_1070);
nor U1190 (N_1190,N_1038,N_1081);
nand U1191 (N_1191,N_1028,N_1014);
nor U1192 (N_1192,N_1044,N_1016);
nor U1193 (N_1193,N_1033,N_1040);
or U1194 (N_1194,N_1062,N_1026);
nand U1195 (N_1195,N_1020,N_1014);
or U1196 (N_1196,N_1036,N_1061);
or U1197 (N_1197,N_1097,N_1058);
nand U1198 (N_1198,N_1054,N_1008);
and U1199 (N_1199,N_1088,N_1098);
or U1200 (N_1200,N_1133,N_1192);
or U1201 (N_1201,N_1167,N_1189);
and U1202 (N_1202,N_1197,N_1187);
nor U1203 (N_1203,N_1177,N_1171);
nand U1204 (N_1204,N_1118,N_1176);
nor U1205 (N_1205,N_1141,N_1159);
or U1206 (N_1206,N_1140,N_1185);
nor U1207 (N_1207,N_1155,N_1135);
and U1208 (N_1208,N_1165,N_1158);
or U1209 (N_1209,N_1138,N_1109);
and U1210 (N_1210,N_1117,N_1134);
or U1211 (N_1211,N_1143,N_1175);
or U1212 (N_1212,N_1128,N_1150);
nor U1213 (N_1213,N_1132,N_1183);
nor U1214 (N_1214,N_1179,N_1121);
nand U1215 (N_1215,N_1152,N_1160);
and U1216 (N_1216,N_1195,N_1145);
nor U1217 (N_1217,N_1180,N_1119);
nor U1218 (N_1218,N_1182,N_1108);
nand U1219 (N_1219,N_1125,N_1169);
nand U1220 (N_1220,N_1123,N_1115);
and U1221 (N_1221,N_1153,N_1111);
xnor U1222 (N_1222,N_1144,N_1101);
or U1223 (N_1223,N_1164,N_1194);
nor U1224 (N_1224,N_1139,N_1100);
xnor U1225 (N_1225,N_1199,N_1148);
and U1226 (N_1226,N_1120,N_1154);
nor U1227 (N_1227,N_1191,N_1196);
or U1228 (N_1228,N_1114,N_1126);
nand U1229 (N_1229,N_1146,N_1124);
nor U1230 (N_1230,N_1113,N_1110);
or U1231 (N_1231,N_1162,N_1137);
nand U1232 (N_1232,N_1156,N_1188);
nand U1233 (N_1233,N_1178,N_1147);
and U1234 (N_1234,N_1190,N_1127);
or U1235 (N_1235,N_1136,N_1181);
nor U1236 (N_1236,N_1173,N_1172);
nand U1237 (N_1237,N_1157,N_1161);
nor U1238 (N_1238,N_1112,N_1170);
nor U1239 (N_1239,N_1174,N_1105);
nand U1240 (N_1240,N_1103,N_1104);
and U1241 (N_1241,N_1163,N_1184);
nor U1242 (N_1242,N_1131,N_1106);
nand U1243 (N_1243,N_1122,N_1186);
nand U1244 (N_1244,N_1149,N_1107);
xor U1245 (N_1245,N_1151,N_1166);
xnor U1246 (N_1246,N_1142,N_1193);
nor U1247 (N_1247,N_1130,N_1102);
nor U1248 (N_1248,N_1198,N_1168);
nor U1249 (N_1249,N_1116,N_1129);
and U1250 (N_1250,N_1111,N_1131);
nor U1251 (N_1251,N_1169,N_1187);
nor U1252 (N_1252,N_1138,N_1116);
and U1253 (N_1253,N_1198,N_1112);
and U1254 (N_1254,N_1108,N_1160);
nor U1255 (N_1255,N_1118,N_1160);
and U1256 (N_1256,N_1130,N_1183);
nand U1257 (N_1257,N_1177,N_1170);
or U1258 (N_1258,N_1182,N_1155);
and U1259 (N_1259,N_1102,N_1148);
nor U1260 (N_1260,N_1171,N_1142);
nand U1261 (N_1261,N_1171,N_1133);
nand U1262 (N_1262,N_1152,N_1173);
nand U1263 (N_1263,N_1121,N_1113);
or U1264 (N_1264,N_1192,N_1136);
or U1265 (N_1265,N_1123,N_1179);
xor U1266 (N_1266,N_1186,N_1180);
and U1267 (N_1267,N_1114,N_1133);
or U1268 (N_1268,N_1179,N_1195);
and U1269 (N_1269,N_1125,N_1170);
nand U1270 (N_1270,N_1167,N_1125);
and U1271 (N_1271,N_1135,N_1173);
and U1272 (N_1272,N_1168,N_1121);
nor U1273 (N_1273,N_1168,N_1167);
and U1274 (N_1274,N_1132,N_1112);
and U1275 (N_1275,N_1111,N_1121);
nand U1276 (N_1276,N_1114,N_1178);
xor U1277 (N_1277,N_1133,N_1116);
xnor U1278 (N_1278,N_1152,N_1193);
or U1279 (N_1279,N_1190,N_1165);
and U1280 (N_1280,N_1134,N_1162);
nand U1281 (N_1281,N_1106,N_1165);
nand U1282 (N_1282,N_1184,N_1183);
nor U1283 (N_1283,N_1172,N_1163);
or U1284 (N_1284,N_1135,N_1156);
or U1285 (N_1285,N_1184,N_1107);
nor U1286 (N_1286,N_1188,N_1187);
and U1287 (N_1287,N_1156,N_1163);
and U1288 (N_1288,N_1136,N_1120);
or U1289 (N_1289,N_1103,N_1121);
xor U1290 (N_1290,N_1135,N_1171);
xor U1291 (N_1291,N_1176,N_1149);
and U1292 (N_1292,N_1131,N_1108);
and U1293 (N_1293,N_1175,N_1191);
or U1294 (N_1294,N_1142,N_1105);
xor U1295 (N_1295,N_1155,N_1192);
nor U1296 (N_1296,N_1118,N_1131);
xor U1297 (N_1297,N_1146,N_1106);
nor U1298 (N_1298,N_1153,N_1124);
xor U1299 (N_1299,N_1163,N_1145);
xor U1300 (N_1300,N_1245,N_1289);
and U1301 (N_1301,N_1241,N_1299);
xnor U1302 (N_1302,N_1253,N_1249);
nor U1303 (N_1303,N_1217,N_1247);
nand U1304 (N_1304,N_1292,N_1270);
xor U1305 (N_1305,N_1295,N_1294);
or U1306 (N_1306,N_1236,N_1282);
nand U1307 (N_1307,N_1229,N_1237);
and U1308 (N_1308,N_1269,N_1223);
xor U1309 (N_1309,N_1286,N_1268);
nor U1310 (N_1310,N_1202,N_1218);
nand U1311 (N_1311,N_1257,N_1291);
xor U1312 (N_1312,N_1204,N_1279);
or U1313 (N_1313,N_1285,N_1220);
xor U1314 (N_1314,N_1200,N_1243);
and U1315 (N_1315,N_1227,N_1224);
or U1316 (N_1316,N_1272,N_1281);
nor U1317 (N_1317,N_1238,N_1297);
or U1318 (N_1318,N_1276,N_1298);
nor U1319 (N_1319,N_1209,N_1266);
or U1320 (N_1320,N_1273,N_1251);
nor U1321 (N_1321,N_1221,N_1275);
nand U1322 (N_1322,N_1230,N_1232);
nand U1323 (N_1323,N_1240,N_1284);
or U1324 (N_1324,N_1214,N_1296);
nor U1325 (N_1325,N_1203,N_1225);
xor U1326 (N_1326,N_1256,N_1248);
or U1327 (N_1327,N_1239,N_1264);
or U1328 (N_1328,N_1280,N_1246);
and U1329 (N_1329,N_1231,N_1288);
nor U1330 (N_1330,N_1205,N_1207);
and U1331 (N_1331,N_1219,N_1254);
nor U1332 (N_1332,N_1262,N_1290);
nand U1333 (N_1333,N_1252,N_1265);
nand U1334 (N_1334,N_1287,N_1208);
and U1335 (N_1335,N_1278,N_1216);
nand U1336 (N_1336,N_1250,N_1201);
and U1337 (N_1337,N_1244,N_1234);
or U1338 (N_1338,N_1258,N_1260);
and U1339 (N_1339,N_1255,N_1215);
nor U1340 (N_1340,N_1267,N_1274);
nor U1341 (N_1341,N_1263,N_1226);
and U1342 (N_1342,N_1211,N_1210);
nand U1343 (N_1343,N_1259,N_1283);
or U1344 (N_1344,N_1235,N_1206);
or U1345 (N_1345,N_1293,N_1222);
nor U1346 (N_1346,N_1277,N_1242);
and U1347 (N_1347,N_1261,N_1271);
or U1348 (N_1348,N_1212,N_1233);
xor U1349 (N_1349,N_1228,N_1213);
nand U1350 (N_1350,N_1228,N_1230);
xnor U1351 (N_1351,N_1283,N_1249);
and U1352 (N_1352,N_1224,N_1276);
and U1353 (N_1353,N_1259,N_1251);
nor U1354 (N_1354,N_1236,N_1220);
and U1355 (N_1355,N_1228,N_1218);
nor U1356 (N_1356,N_1253,N_1297);
nor U1357 (N_1357,N_1293,N_1245);
nand U1358 (N_1358,N_1291,N_1285);
nand U1359 (N_1359,N_1206,N_1222);
nand U1360 (N_1360,N_1239,N_1218);
or U1361 (N_1361,N_1287,N_1213);
or U1362 (N_1362,N_1287,N_1288);
nor U1363 (N_1363,N_1226,N_1284);
and U1364 (N_1364,N_1231,N_1233);
xnor U1365 (N_1365,N_1284,N_1225);
nor U1366 (N_1366,N_1265,N_1271);
and U1367 (N_1367,N_1271,N_1287);
nand U1368 (N_1368,N_1265,N_1227);
nand U1369 (N_1369,N_1235,N_1285);
xnor U1370 (N_1370,N_1248,N_1250);
nand U1371 (N_1371,N_1223,N_1292);
and U1372 (N_1372,N_1228,N_1288);
xnor U1373 (N_1373,N_1203,N_1288);
or U1374 (N_1374,N_1274,N_1294);
or U1375 (N_1375,N_1260,N_1291);
nand U1376 (N_1376,N_1278,N_1203);
nand U1377 (N_1377,N_1239,N_1210);
nand U1378 (N_1378,N_1267,N_1299);
nor U1379 (N_1379,N_1274,N_1277);
nor U1380 (N_1380,N_1274,N_1211);
nor U1381 (N_1381,N_1206,N_1255);
nand U1382 (N_1382,N_1216,N_1281);
nand U1383 (N_1383,N_1247,N_1258);
and U1384 (N_1384,N_1286,N_1238);
nor U1385 (N_1385,N_1200,N_1221);
or U1386 (N_1386,N_1206,N_1299);
nor U1387 (N_1387,N_1294,N_1226);
or U1388 (N_1388,N_1262,N_1250);
nor U1389 (N_1389,N_1224,N_1265);
or U1390 (N_1390,N_1218,N_1274);
nand U1391 (N_1391,N_1234,N_1218);
and U1392 (N_1392,N_1245,N_1299);
nor U1393 (N_1393,N_1295,N_1256);
xnor U1394 (N_1394,N_1239,N_1225);
xor U1395 (N_1395,N_1222,N_1239);
xor U1396 (N_1396,N_1254,N_1244);
xor U1397 (N_1397,N_1281,N_1201);
xor U1398 (N_1398,N_1220,N_1258);
and U1399 (N_1399,N_1276,N_1282);
nand U1400 (N_1400,N_1344,N_1361);
xnor U1401 (N_1401,N_1324,N_1365);
or U1402 (N_1402,N_1360,N_1338);
and U1403 (N_1403,N_1398,N_1349);
xnor U1404 (N_1404,N_1363,N_1376);
xnor U1405 (N_1405,N_1326,N_1356);
xor U1406 (N_1406,N_1304,N_1350);
xnor U1407 (N_1407,N_1325,N_1354);
xor U1408 (N_1408,N_1319,N_1332);
nor U1409 (N_1409,N_1369,N_1303);
or U1410 (N_1410,N_1381,N_1373);
and U1411 (N_1411,N_1339,N_1394);
and U1412 (N_1412,N_1371,N_1358);
xor U1413 (N_1413,N_1382,N_1367);
xor U1414 (N_1414,N_1374,N_1393);
nor U1415 (N_1415,N_1334,N_1375);
xnor U1416 (N_1416,N_1352,N_1387);
and U1417 (N_1417,N_1336,N_1312);
or U1418 (N_1418,N_1359,N_1335);
xor U1419 (N_1419,N_1309,N_1306);
and U1420 (N_1420,N_1337,N_1355);
xor U1421 (N_1421,N_1330,N_1321);
and U1422 (N_1422,N_1311,N_1397);
nor U1423 (N_1423,N_1341,N_1351);
nor U1424 (N_1424,N_1362,N_1378);
xnor U1425 (N_1425,N_1300,N_1315);
or U1426 (N_1426,N_1328,N_1379);
xnor U1427 (N_1427,N_1310,N_1392);
and U1428 (N_1428,N_1316,N_1372);
or U1429 (N_1429,N_1389,N_1391);
and U1430 (N_1430,N_1345,N_1384);
nand U1431 (N_1431,N_1364,N_1323);
nand U1432 (N_1432,N_1386,N_1340);
nor U1433 (N_1433,N_1353,N_1308);
or U1434 (N_1434,N_1327,N_1318);
nor U1435 (N_1435,N_1343,N_1390);
nand U1436 (N_1436,N_1347,N_1380);
nor U1437 (N_1437,N_1333,N_1301);
xnor U1438 (N_1438,N_1346,N_1317);
or U1439 (N_1439,N_1314,N_1366);
xor U1440 (N_1440,N_1329,N_1322);
xor U1441 (N_1441,N_1395,N_1399);
and U1442 (N_1442,N_1302,N_1357);
xnor U1443 (N_1443,N_1305,N_1385);
nand U1444 (N_1444,N_1370,N_1383);
nand U1445 (N_1445,N_1396,N_1307);
nor U1446 (N_1446,N_1368,N_1342);
or U1447 (N_1447,N_1313,N_1320);
xnor U1448 (N_1448,N_1388,N_1348);
nand U1449 (N_1449,N_1331,N_1377);
and U1450 (N_1450,N_1369,N_1334);
and U1451 (N_1451,N_1365,N_1361);
nand U1452 (N_1452,N_1372,N_1373);
or U1453 (N_1453,N_1305,N_1375);
nor U1454 (N_1454,N_1399,N_1341);
nor U1455 (N_1455,N_1351,N_1313);
nor U1456 (N_1456,N_1327,N_1332);
nor U1457 (N_1457,N_1324,N_1363);
xor U1458 (N_1458,N_1328,N_1362);
nand U1459 (N_1459,N_1334,N_1350);
and U1460 (N_1460,N_1386,N_1314);
or U1461 (N_1461,N_1389,N_1383);
xnor U1462 (N_1462,N_1353,N_1397);
and U1463 (N_1463,N_1392,N_1340);
nor U1464 (N_1464,N_1331,N_1371);
nor U1465 (N_1465,N_1350,N_1337);
nor U1466 (N_1466,N_1332,N_1378);
and U1467 (N_1467,N_1383,N_1323);
nor U1468 (N_1468,N_1358,N_1350);
or U1469 (N_1469,N_1315,N_1349);
or U1470 (N_1470,N_1328,N_1360);
nand U1471 (N_1471,N_1349,N_1399);
or U1472 (N_1472,N_1303,N_1317);
or U1473 (N_1473,N_1325,N_1369);
nand U1474 (N_1474,N_1323,N_1351);
and U1475 (N_1475,N_1341,N_1376);
and U1476 (N_1476,N_1394,N_1398);
xnor U1477 (N_1477,N_1338,N_1335);
nor U1478 (N_1478,N_1345,N_1367);
xnor U1479 (N_1479,N_1329,N_1378);
nor U1480 (N_1480,N_1326,N_1375);
nor U1481 (N_1481,N_1396,N_1385);
and U1482 (N_1482,N_1385,N_1334);
nand U1483 (N_1483,N_1384,N_1301);
nand U1484 (N_1484,N_1310,N_1365);
or U1485 (N_1485,N_1329,N_1363);
nor U1486 (N_1486,N_1397,N_1361);
nand U1487 (N_1487,N_1384,N_1387);
and U1488 (N_1488,N_1354,N_1308);
nor U1489 (N_1489,N_1370,N_1384);
and U1490 (N_1490,N_1310,N_1315);
nand U1491 (N_1491,N_1349,N_1393);
nand U1492 (N_1492,N_1305,N_1384);
or U1493 (N_1493,N_1315,N_1338);
nand U1494 (N_1494,N_1355,N_1368);
nand U1495 (N_1495,N_1329,N_1387);
xnor U1496 (N_1496,N_1310,N_1303);
nand U1497 (N_1497,N_1392,N_1364);
xor U1498 (N_1498,N_1377,N_1323);
and U1499 (N_1499,N_1364,N_1336);
nand U1500 (N_1500,N_1408,N_1453);
nor U1501 (N_1501,N_1406,N_1468);
nand U1502 (N_1502,N_1439,N_1437);
nor U1503 (N_1503,N_1411,N_1438);
and U1504 (N_1504,N_1479,N_1455);
nand U1505 (N_1505,N_1445,N_1498);
nand U1506 (N_1506,N_1414,N_1451);
nor U1507 (N_1507,N_1422,N_1407);
and U1508 (N_1508,N_1450,N_1475);
and U1509 (N_1509,N_1456,N_1476);
or U1510 (N_1510,N_1416,N_1490);
nand U1511 (N_1511,N_1458,N_1442);
and U1512 (N_1512,N_1412,N_1457);
and U1513 (N_1513,N_1461,N_1469);
nand U1514 (N_1514,N_1425,N_1499);
or U1515 (N_1515,N_1403,N_1477);
xnor U1516 (N_1516,N_1415,N_1418);
nand U1517 (N_1517,N_1428,N_1410);
xor U1518 (N_1518,N_1473,N_1478);
and U1519 (N_1519,N_1452,N_1459);
and U1520 (N_1520,N_1474,N_1436);
xor U1521 (N_1521,N_1417,N_1482);
xor U1522 (N_1522,N_1423,N_1470);
nor U1523 (N_1523,N_1462,N_1449);
or U1524 (N_1524,N_1448,N_1487);
nor U1525 (N_1525,N_1467,N_1464);
nor U1526 (N_1526,N_1444,N_1430);
and U1527 (N_1527,N_1491,N_1494);
nand U1528 (N_1528,N_1486,N_1447);
nand U1529 (N_1529,N_1402,N_1484);
and U1530 (N_1530,N_1463,N_1480);
or U1531 (N_1531,N_1481,N_1426);
nand U1532 (N_1532,N_1400,N_1413);
and U1533 (N_1533,N_1472,N_1440);
or U1534 (N_1534,N_1431,N_1419);
and U1535 (N_1535,N_1424,N_1483);
nor U1536 (N_1536,N_1401,N_1488);
and U1537 (N_1537,N_1432,N_1421);
nor U1538 (N_1538,N_1405,N_1460);
xor U1539 (N_1539,N_1434,N_1446);
or U1540 (N_1540,N_1485,N_1429);
xor U1541 (N_1541,N_1497,N_1409);
xnor U1542 (N_1542,N_1441,N_1435);
xor U1543 (N_1543,N_1492,N_1493);
nor U1544 (N_1544,N_1454,N_1465);
nor U1545 (N_1545,N_1496,N_1433);
or U1546 (N_1546,N_1495,N_1427);
nor U1547 (N_1547,N_1471,N_1404);
nor U1548 (N_1548,N_1420,N_1466);
nor U1549 (N_1549,N_1443,N_1489);
nor U1550 (N_1550,N_1453,N_1466);
xor U1551 (N_1551,N_1451,N_1479);
nand U1552 (N_1552,N_1483,N_1409);
xnor U1553 (N_1553,N_1475,N_1490);
and U1554 (N_1554,N_1443,N_1451);
and U1555 (N_1555,N_1425,N_1481);
nor U1556 (N_1556,N_1437,N_1426);
or U1557 (N_1557,N_1492,N_1434);
nor U1558 (N_1558,N_1472,N_1420);
or U1559 (N_1559,N_1439,N_1476);
and U1560 (N_1560,N_1403,N_1485);
and U1561 (N_1561,N_1478,N_1431);
nand U1562 (N_1562,N_1497,N_1421);
nor U1563 (N_1563,N_1437,N_1486);
and U1564 (N_1564,N_1446,N_1452);
or U1565 (N_1565,N_1460,N_1484);
or U1566 (N_1566,N_1443,N_1484);
and U1567 (N_1567,N_1409,N_1417);
nand U1568 (N_1568,N_1485,N_1480);
nand U1569 (N_1569,N_1428,N_1433);
nand U1570 (N_1570,N_1418,N_1452);
or U1571 (N_1571,N_1426,N_1458);
and U1572 (N_1572,N_1458,N_1400);
or U1573 (N_1573,N_1440,N_1441);
nor U1574 (N_1574,N_1486,N_1494);
or U1575 (N_1575,N_1425,N_1408);
nand U1576 (N_1576,N_1499,N_1486);
or U1577 (N_1577,N_1428,N_1472);
nand U1578 (N_1578,N_1415,N_1409);
nand U1579 (N_1579,N_1451,N_1458);
nand U1580 (N_1580,N_1432,N_1496);
or U1581 (N_1581,N_1451,N_1424);
nor U1582 (N_1582,N_1490,N_1436);
xor U1583 (N_1583,N_1442,N_1425);
nor U1584 (N_1584,N_1406,N_1435);
xnor U1585 (N_1585,N_1425,N_1414);
or U1586 (N_1586,N_1476,N_1442);
or U1587 (N_1587,N_1467,N_1443);
nor U1588 (N_1588,N_1489,N_1421);
or U1589 (N_1589,N_1458,N_1453);
nand U1590 (N_1590,N_1445,N_1460);
nand U1591 (N_1591,N_1496,N_1424);
xnor U1592 (N_1592,N_1441,N_1464);
or U1593 (N_1593,N_1498,N_1474);
xnor U1594 (N_1594,N_1429,N_1471);
or U1595 (N_1595,N_1411,N_1418);
xor U1596 (N_1596,N_1416,N_1436);
nand U1597 (N_1597,N_1413,N_1458);
nor U1598 (N_1598,N_1443,N_1403);
and U1599 (N_1599,N_1406,N_1478);
xor U1600 (N_1600,N_1517,N_1594);
or U1601 (N_1601,N_1570,N_1585);
nor U1602 (N_1602,N_1520,N_1550);
and U1603 (N_1603,N_1590,N_1574);
nand U1604 (N_1604,N_1547,N_1527);
and U1605 (N_1605,N_1571,N_1515);
nand U1606 (N_1606,N_1524,N_1521);
and U1607 (N_1607,N_1561,N_1579);
xor U1608 (N_1608,N_1516,N_1511);
and U1609 (N_1609,N_1539,N_1531);
nand U1610 (N_1610,N_1540,N_1564);
nor U1611 (N_1611,N_1541,N_1592);
and U1612 (N_1612,N_1587,N_1510);
nand U1613 (N_1613,N_1591,N_1513);
nor U1614 (N_1614,N_1536,N_1584);
nand U1615 (N_1615,N_1502,N_1582);
xor U1616 (N_1616,N_1577,N_1503);
xor U1617 (N_1617,N_1528,N_1545);
or U1618 (N_1618,N_1558,N_1573);
nand U1619 (N_1619,N_1538,N_1522);
or U1620 (N_1620,N_1578,N_1544);
xor U1621 (N_1621,N_1559,N_1518);
and U1622 (N_1622,N_1580,N_1549);
or U1623 (N_1623,N_1525,N_1598);
nand U1624 (N_1624,N_1551,N_1501);
nor U1625 (N_1625,N_1529,N_1568);
nand U1626 (N_1626,N_1504,N_1555);
nand U1627 (N_1627,N_1546,N_1523);
or U1628 (N_1628,N_1556,N_1567);
nor U1629 (N_1629,N_1553,N_1596);
xnor U1630 (N_1630,N_1560,N_1557);
and U1631 (N_1631,N_1569,N_1588);
or U1632 (N_1632,N_1563,N_1509);
and U1633 (N_1633,N_1581,N_1506);
nand U1634 (N_1634,N_1599,N_1519);
and U1635 (N_1635,N_1500,N_1508);
and U1636 (N_1636,N_1537,N_1552);
and U1637 (N_1637,N_1507,N_1514);
nor U1638 (N_1638,N_1534,N_1583);
and U1639 (N_1639,N_1543,N_1532);
and U1640 (N_1640,N_1589,N_1562);
or U1641 (N_1641,N_1548,N_1512);
xnor U1642 (N_1642,N_1575,N_1576);
nor U1643 (N_1643,N_1526,N_1542);
xor U1644 (N_1644,N_1530,N_1566);
or U1645 (N_1645,N_1595,N_1533);
nand U1646 (N_1646,N_1565,N_1597);
or U1647 (N_1647,N_1554,N_1572);
or U1648 (N_1648,N_1593,N_1535);
and U1649 (N_1649,N_1505,N_1586);
nand U1650 (N_1650,N_1576,N_1513);
nor U1651 (N_1651,N_1503,N_1540);
xor U1652 (N_1652,N_1585,N_1515);
nand U1653 (N_1653,N_1534,N_1572);
xnor U1654 (N_1654,N_1522,N_1513);
xnor U1655 (N_1655,N_1504,N_1523);
and U1656 (N_1656,N_1575,N_1506);
nand U1657 (N_1657,N_1531,N_1527);
nand U1658 (N_1658,N_1534,N_1589);
or U1659 (N_1659,N_1528,N_1522);
or U1660 (N_1660,N_1599,N_1588);
and U1661 (N_1661,N_1522,N_1556);
or U1662 (N_1662,N_1548,N_1556);
xor U1663 (N_1663,N_1589,N_1542);
nor U1664 (N_1664,N_1543,N_1531);
xor U1665 (N_1665,N_1553,N_1519);
and U1666 (N_1666,N_1571,N_1544);
or U1667 (N_1667,N_1564,N_1524);
nor U1668 (N_1668,N_1588,N_1581);
nand U1669 (N_1669,N_1517,N_1528);
xor U1670 (N_1670,N_1543,N_1508);
and U1671 (N_1671,N_1545,N_1590);
and U1672 (N_1672,N_1546,N_1545);
xnor U1673 (N_1673,N_1586,N_1591);
or U1674 (N_1674,N_1555,N_1514);
or U1675 (N_1675,N_1577,N_1580);
and U1676 (N_1676,N_1532,N_1578);
or U1677 (N_1677,N_1525,N_1510);
nand U1678 (N_1678,N_1598,N_1508);
and U1679 (N_1679,N_1513,N_1530);
and U1680 (N_1680,N_1550,N_1563);
or U1681 (N_1681,N_1575,N_1557);
nor U1682 (N_1682,N_1535,N_1573);
or U1683 (N_1683,N_1547,N_1562);
nor U1684 (N_1684,N_1576,N_1584);
xnor U1685 (N_1685,N_1558,N_1583);
or U1686 (N_1686,N_1508,N_1557);
nand U1687 (N_1687,N_1518,N_1542);
nor U1688 (N_1688,N_1594,N_1529);
nand U1689 (N_1689,N_1594,N_1521);
nor U1690 (N_1690,N_1512,N_1577);
nand U1691 (N_1691,N_1538,N_1524);
and U1692 (N_1692,N_1542,N_1596);
or U1693 (N_1693,N_1504,N_1508);
nand U1694 (N_1694,N_1538,N_1515);
nand U1695 (N_1695,N_1527,N_1580);
nand U1696 (N_1696,N_1513,N_1534);
xor U1697 (N_1697,N_1566,N_1539);
nand U1698 (N_1698,N_1533,N_1596);
or U1699 (N_1699,N_1512,N_1591);
nor U1700 (N_1700,N_1673,N_1672);
nor U1701 (N_1701,N_1658,N_1628);
xnor U1702 (N_1702,N_1692,N_1675);
nor U1703 (N_1703,N_1683,N_1629);
nand U1704 (N_1704,N_1642,N_1698);
nand U1705 (N_1705,N_1609,N_1652);
xor U1706 (N_1706,N_1678,N_1646);
nand U1707 (N_1707,N_1688,N_1643);
xnor U1708 (N_1708,N_1659,N_1621);
or U1709 (N_1709,N_1685,N_1641);
and U1710 (N_1710,N_1699,N_1644);
or U1711 (N_1711,N_1633,N_1661);
nor U1712 (N_1712,N_1687,N_1679);
nor U1713 (N_1713,N_1622,N_1639);
nor U1714 (N_1714,N_1649,N_1668);
and U1715 (N_1715,N_1696,N_1601);
xnor U1716 (N_1716,N_1657,N_1610);
nor U1717 (N_1717,N_1623,N_1604);
xor U1718 (N_1718,N_1682,N_1614);
and U1719 (N_1719,N_1686,N_1697);
or U1720 (N_1720,N_1611,N_1636);
or U1721 (N_1721,N_1600,N_1620);
and U1722 (N_1722,N_1606,N_1653);
xor U1723 (N_1723,N_1645,N_1626);
nand U1724 (N_1724,N_1613,N_1663);
xor U1725 (N_1725,N_1608,N_1640);
nand U1726 (N_1726,N_1632,N_1617);
nor U1727 (N_1727,N_1695,N_1676);
nand U1728 (N_1728,N_1605,N_1615);
nand U1729 (N_1729,N_1619,N_1665);
nor U1730 (N_1730,N_1669,N_1660);
nand U1731 (N_1731,N_1662,N_1651);
nor U1732 (N_1732,N_1624,N_1603);
and U1733 (N_1733,N_1631,N_1681);
nor U1734 (N_1734,N_1691,N_1671);
nor U1735 (N_1735,N_1648,N_1627);
nand U1736 (N_1736,N_1670,N_1625);
nor U1737 (N_1737,N_1667,N_1635);
nand U1738 (N_1738,N_1618,N_1656);
nand U1739 (N_1739,N_1630,N_1664);
or U1740 (N_1740,N_1607,N_1690);
nand U1741 (N_1741,N_1680,N_1650);
and U1742 (N_1742,N_1693,N_1689);
and U1743 (N_1743,N_1654,N_1634);
xnor U1744 (N_1744,N_1638,N_1616);
and U1745 (N_1745,N_1694,N_1612);
nand U1746 (N_1746,N_1684,N_1647);
nor U1747 (N_1747,N_1637,N_1655);
xnor U1748 (N_1748,N_1677,N_1666);
or U1749 (N_1749,N_1602,N_1674);
or U1750 (N_1750,N_1696,N_1633);
or U1751 (N_1751,N_1613,N_1608);
xnor U1752 (N_1752,N_1648,N_1692);
xnor U1753 (N_1753,N_1645,N_1630);
nand U1754 (N_1754,N_1688,N_1661);
nor U1755 (N_1755,N_1697,N_1630);
xnor U1756 (N_1756,N_1646,N_1635);
or U1757 (N_1757,N_1679,N_1671);
nor U1758 (N_1758,N_1656,N_1624);
and U1759 (N_1759,N_1674,N_1699);
nand U1760 (N_1760,N_1698,N_1656);
nor U1761 (N_1761,N_1642,N_1607);
xor U1762 (N_1762,N_1668,N_1644);
xor U1763 (N_1763,N_1628,N_1647);
nand U1764 (N_1764,N_1609,N_1680);
nand U1765 (N_1765,N_1624,N_1684);
or U1766 (N_1766,N_1637,N_1669);
nand U1767 (N_1767,N_1646,N_1621);
and U1768 (N_1768,N_1693,N_1690);
or U1769 (N_1769,N_1627,N_1605);
or U1770 (N_1770,N_1680,N_1639);
xor U1771 (N_1771,N_1605,N_1626);
and U1772 (N_1772,N_1605,N_1648);
nor U1773 (N_1773,N_1601,N_1688);
or U1774 (N_1774,N_1644,N_1610);
and U1775 (N_1775,N_1626,N_1672);
nand U1776 (N_1776,N_1628,N_1673);
or U1777 (N_1777,N_1660,N_1602);
xnor U1778 (N_1778,N_1657,N_1614);
and U1779 (N_1779,N_1608,N_1685);
and U1780 (N_1780,N_1689,N_1616);
nand U1781 (N_1781,N_1668,N_1621);
nor U1782 (N_1782,N_1660,N_1655);
nor U1783 (N_1783,N_1641,N_1647);
or U1784 (N_1784,N_1684,N_1639);
and U1785 (N_1785,N_1670,N_1679);
or U1786 (N_1786,N_1637,N_1685);
xnor U1787 (N_1787,N_1684,N_1692);
or U1788 (N_1788,N_1697,N_1682);
nand U1789 (N_1789,N_1629,N_1661);
and U1790 (N_1790,N_1612,N_1655);
nor U1791 (N_1791,N_1651,N_1668);
and U1792 (N_1792,N_1637,N_1647);
or U1793 (N_1793,N_1607,N_1666);
and U1794 (N_1794,N_1662,N_1653);
xor U1795 (N_1795,N_1692,N_1625);
or U1796 (N_1796,N_1621,N_1652);
nor U1797 (N_1797,N_1673,N_1694);
xnor U1798 (N_1798,N_1695,N_1603);
xor U1799 (N_1799,N_1694,N_1635);
xor U1800 (N_1800,N_1785,N_1754);
and U1801 (N_1801,N_1708,N_1751);
xor U1802 (N_1802,N_1781,N_1777);
and U1803 (N_1803,N_1755,N_1728);
nor U1804 (N_1804,N_1734,N_1723);
or U1805 (N_1805,N_1768,N_1707);
or U1806 (N_1806,N_1786,N_1745);
or U1807 (N_1807,N_1749,N_1722);
and U1808 (N_1808,N_1703,N_1729);
nor U1809 (N_1809,N_1775,N_1796);
xnor U1810 (N_1810,N_1750,N_1763);
nor U1811 (N_1811,N_1760,N_1773);
nand U1812 (N_1812,N_1787,N_1742);
nand U1813 (N_1813,N_1782,N_1744);
xor U1814 (N_1814,N_1727,N_1736);
and U1815 (N_1815,N_1718,N_1770);
or U1816 (N_1816,N_1790,N_1712);
nor U1817 (N_1817,N_1779,N_1731);
and U1818 (N_1818,N_1743,N_1778);
nor U1819 (N_1819,N_1733,N_1776);
or U1820 (N_1820,N_1724,N_1761);
xor U1821 (N_1821,N_1720,N_1753);
or U1822 (N_1822,N_1794,N_1737);
nand U1823 (N_1823,N_1746,N_1799);
xor U1824 (N_1824,N_1735,N_1711);
nor U1825 (N_1825,N_1769,N_1772);
nand U1826 (N_1826,N_1713,N_1756);
xor U1827 (N_1827,N_1792,N_1766);
and U1828 (N_1828,N_1738,N_1797);
nor U1829 (N_1829,N_1771,N_1780);
xor U1830 (N_1830,N_1706,N_1767);
or U1831 (N_1831,N_1757,N_1759);
and U1832 (N_1832,N_1702,N_1739);
xor U1833 (N_1833,N_1747,N_1764);
or U1834 (N_1834,N_1715,N_1719);
nor U1835 (N_1835,N_1795,N_1714);
xnor U1836 (N_1836,N_1752,N_1717);
nor U1837 (N_1837,N_1788,N_1710);
and U1838 (N_1838,N_1758,N_1765);
nand U1839 (N_1839,N_1701,N_1725);
xnor U1840 (N_1840,N_1730,N_1732);
xnor U1841 (N_1841,N_1748,N_1721);
or U1842 (N_1842,N_1700,N_1741);
or U1843 (N_1843,N_1784,N_1704);
and U1844 (N_1844,N_1716,N_1774);
xnor U1845 (N_1845,N_1791,N_1726);
nor U1846 (N_1846,N_1705,N_1762);
or U1847 (N_1847,N_1793,N_1789);
and U1848 (N_1848,N_1709,N_1783);
nand U1849 (N_1849,N_1740,N_1798);
and U1850 (N_1850,N_1701,N_1732);
or U1851 (N_1851,N_1734,N_1702);
or U1852 (N_1852,N_1700,N_1780);
nor U1853 (N_1853,N_1757,N_1798);
and U1854 (N_1854,N_1752,N_1781);
or U1855 (N_1855,N_1773,N_1720);
nand U1856 (N_1856,N_1738,N_1730);
or U1857 (N_1857,N_1738,N_1778);
and U1858 (N_1858,N_1752,N_1765);
and U1859 (N_1859,N_1779,N_1758);
and U1860 (N_1860,N_1791,N_1700);
or U1861 (N_1861,N_1734,N_1795);
nor U1862 (N_1862,N_1739,N_1789);
nor U1863 (N_1863,N_1796,N_1728);
xor U1864 (N_1864,N_1784,N_1713);
and U1865 (N_1865,N_1748,N_1723);
nand U1866 (N_1866,N_1744,N_1747);
xnor U1867 (N_1867,N_1701,N_1730);
nand U1868 (N_1868,N_1750,N_1739);
or U1869 (N_1869,N_1773,N_1766);
nand U1870 (N_1870,N_1769,N_1783);
and U1871 (N_1871,N_1712,N_1711);
nor U1872 (N_1872,N_1788,N_1708);
nor U1873 (N_1873,N_1704,N_1731);
nand U1874 (N_1874,N_1765,N_1732);
or U1875 (N_1875,N_1767,N_1719);
nor U1876 (N_1876,N_1753,N_1700);
and U1877 (N_1877,N_1776,N_1764);
xor U1878 (N_1878,N_1713,N_1745);
or U1879 (N_1879,N_1746,N_1704);
nor U1880 (N_1880,N_1770,N_1783);
nand U1881 (N_1881,N_1717,N_1710);
nand U1882 (N_1882,N_1704,N_1711);
nand U1883 (N_1883,N_1761,N_1770);
nand U1884 (N_1884,N_1757,N_1756);
xor U1885 (N_1885,N_1799,N_1792);
xor U1886 (N_1886,N_1761,N_1703);
and U1887 (N_1887,N_1716,N_1712);
nand U1888 (N_1888,N_1724,N_1783);
nor U1889 (N_1889,N_1760,N_1714);
or U1890 (N_1890,N_1762,N_1776);
or U1891 (N_1891,N_1787,N_1769);
and U1892 (N_1892,N_1760,N_1784);
or U1893 (N_1893,N_1709,N_1770);
or U1894 (N_1894,N_1746,N_1715);
nor U1895 (N_1895,N_1747,N_1709);
or U1896 (N_1896,N_1743,N_1751);
nand U1897 (N_1897,N_1754,N_1746);
or U1898 (N_1898,N_1744,N_1759);
or U1899 (N_1899,N_1757,N_1782);
nor U1900 (N_1900,N_1894,N_1841);
nand U1901 (N_1901,N_1803,N_1896);
and U1902 (N_1902,N_1812,N_1873);
or U1903 (N_1903,N_1857,N_1827);
nand U1904 (N_1904,N_1872,N_1847);
and U1905 (N_1905,N_1815,N_1811);
and U1906 (N_1906,N_1869,N_1855);
and U1907 (N_1907,N_1883,N_1868);
nand U1908 (N_1908,N_1890,N_1810);
or U1909 (N_1909,N_1878,N_1843);
or U1910 (N_1910,N_1853,N_1880);
or U1911 (N_1911,N_1826,N_1840);
nand U1912 (N_1912,N_1886,N_1842);
nand U1913 (N_1913,N_1859,N_1837);
or U1914 (N_1914,N_1808,N_1899);
and U1915 (N_1915,N_1825,N_1865);
xor U1916 (N_1916,N_1889,N_1833);
nor U1917 (N_1917,N_1881,N_1858);
nor U1918 (N_1918,N_1820,N_1882);
and U1919 (N_1919,N_1836,N_1852);
and U1920 (N_1920,N_1834,N_1864);
xnor U1921 (N_1921,N_1844,N_1823);
nand U1922 (N_1922,N_1818,N_1832);
nor U1923 (N_1923,N_1814,N_1822);
nand U1924 (N_1924,N_1849,N_1888);
xnor U1925 (N_1925,N_1856,N_1851);
nand U1926 (N_1926,N_1835,N_1830);
nor U1927 (N_1927,N_1877,N_1875);
xnor U1928 (N_1928,N_1806,N_1893);
nor U1929 (N_1929,N_1804,N_1850);
nand U1930 (N_1930,N_1871,N_1831);
and U1931 (N_1931,N_1829,N_1828);
nor U1932 (N_1932,N_1854,N_1874);
nor U1933 (N_1933,N_1805,N_1895);
or U1934 (N_1934,N_1891,N_1885);
nor U1935 (N_1935,N_1845,N_1839);
nand U1936 (N_1936,N_1898,N_1801);
nand U1937 (N_1937,N_1867,N_1816);
or U1938 (N_1938,N_1807,N_1862);
and U1939 (N_1939,N_1809,N_1838);
xnor U1940 (N_1940,N_1846,N_1824);
or U1941 (N_1941,N_1866,N_1870);
nand U1942 (N_1942,N_1861,N_1887);
and U1943 (N_1943,N_1819,N_1802);
xnor U1944 (N_1944,N_1817,N_1879);
and U1945 (N_1945,N_1821,N_1884);
nand U1946 (N_1946,N_1892,N_1813);
nor U1947 (N_1947,N_1860,N_1848);
or U1948 (N_1948,N_1800,N_1863);
xor U1949 (N_1949,N_1876,N_1897);
or U1950 (N_1950,N_1811,N_1878);
xor U1951 (N_1951,N_1824,N_1845);
or U1952 (N_1952,N_1885,N_1807);
xor U1953 (N_1953,N_1832,N_1824);
xnor U1954 (N_1954,N_1897,N_1857);
xnor U1955 (N_1955,N_1863,N_1877);
and U1956 (N_1956,N_1846,N_1825);
or U1957 (N_1957,N_1801,N_1840);
or U1958 (N_1958,N_1820,N_1839);
nor U1959 (N_1959,N_1802,N_1864);
or U1960 (N_1960,N_1899,N_1834);
nor U1961 (N_1961,N_1868,N_1880);
or U1962 (N_1962,N_1875,N_1848);
nand U1963 (N_1963,N_1846,N_1810);
and U1964 (N_1964,N_1808,N_1866);
nor U1965 (N_1965,N_1815,N_1827);
nand U1966 (N_1966,N_1818,N_1805);
nand U1967 (N_1967,N_1881,N_1848);
xor U1968 (N_1968,N_1814,N_1831);
and U1969 (N_1969,N_1823,N_1847);
nand U1970 (N_1970,N_1896,N_1843);
xor U1971 (N_1971,N_1851,N_1881);
nor U1972 (N_1972,N_1878,N_1849);
nor U1973 (N_1973,N_1870,N_1898);
xnor U1974 (N_1974,N_1860,N_1868);
or U1975 (N_1975,N_1859,N_1891);
or U1976 (N_1976,N_1892,N_1881);
or U1977 (N_1977,N_1880,N_1809);
xnor U1978 (N_1978,N_1889,N_1896);
xor U1979 (N_1979,N_1814,N_1875);
nand U1980 (N_1980,N_1820,N_1869);
nor U1981 (N_1981,N_1869,N_1814);
and U1982 (N_1982,N_1888,N_1883);
nor U1983 (N_1983,N_1897,N_1878);
nor U1984 (N_1984,N_1897,N_1838);
and U1985 (N_1985,N_1803,N_1870);
nor U1986 (N_1986,N_1884,N_1812);
xnor U1987 (N_1987,N_1873,N_1823);
nor U1988 (N_1988,N_1870,N_1871);
nor U1989 (N_1989,N_1871,N_1867);
xnor U1990 (N_1990,N_1834,N_1813);
and U1991 (N_1991,N_1863,N_1859);
nand U1992 (N_1992,N_1877,N_1864);
xnor U1993 (N_1993,N_1810,N_1813);
xnor U1994 (N_1994,N_1827,N_1873);
and U1995 (N_1995,N_1818,N_1845);
nor U1996 (N_1996,N_1878,N_1832);
nor U1997 (N_1997,N_1815,N_1890);
nor U1998 (N_1998,N_1822,N_1810);
and U1999 (N_1999,N_1879,N_1841);
nor U2000 (N_2000,N_1987,N_1925);
and U2001 (N_2001,N_1907,N_1918);
nor U2002 (N_2002,N_1955,N_1981);
or U2003 (N_2003,N_1938,N_1930);
and U2004 (N_2004,N_1959,N_1951);
nor U2005 (N_2005,N_1921,N_1904);
xor U2006 (N_2006,N_1971,N_1931);
nor U2007 (N_2007,N_1913,N_1915);
nand U2008 (N_2008,N_1986,N_1927);
nand U2009 (N_2009,N_1917,N_1970);
and U2010 (N_2010,N_1978,N_1929);
xor U2011 (N_2011,N_1982,N_1924);
and U2012 (N_2012,N_1946,N_1936);
nor U2013 (N_2013,N_1960,N_1932);
nand U2014 (N_2014,N_1995,N_1952);
and U2015 (N_2015,N_1956,N_1916);
xnor U2016 (N_2016,N_1984,N_1906);
and U2017 (N_2017,N_1997,N_1993);
nor U2018 (N_2018,N_1994,N_1928);
nor U2019 (N_2019,N_1998,N_1919);
or U2020 (N_2020,N_1908,N_1976);
nand U2021 (N_2021,N_1912,N_1991);
and U2022 (N_2022,N_1974,N_1941);
nand U2023 (N_2023,N_1923,N_1968);
nand U2024 (N_2024,N_1980,N_1937);
nor U2025 (N_2025,N_1958,N_1969);
or U2026 (N_2026,N_1944,N_1999);
xnor U2027 (N_2027,N_1954,N_1996);
and U2028 (N_2028,N_1900,N_1911);
nand U2029 (N_2029,N_1967,N_1975);
nor U2030 (N_2030,N_1945,N_1920);
xor U2031 (N_2031,N_1962,N_1942);
or U2032 (N_2032,N_1914,N_1973);
nand U2033 (N_2033,N_1979,N_1933);
or U2034 (N_2034,N_1902,N_1901);
nor U2035 (N_2035,N_1972,N_1926);
nor U2036 (N_2036,N_1950,N_1963);
nand U2037 (N_2037,N_1988,N_1990);
xor U2038 (N_2038,N_1948,N_1909);
and U2039 (N_2039,N_1966,N_1903);
nand U2040 (N_2040,N_1949,N_1992);
and U2041 (N_2041,N_1939,N_1943);
xor U2042 (N_2042,N_1905,N_1940);
nand U2043 (N_2043,N_1953,N_1964);
and U2044 (N_2044,N_1934,N_1961);
nand U2045 (N_2045,N_1922,N_1977);
nor U2046 (N_2046,N_1989,N_1910);
and U2047 (N_2047,N_1985,N_1935);
xor U2048 (N_2048,N_1983,N_1957);
and U2049 (N_2049,N_1947,N_1965);
and U2050 (N_2050,N_1901,N_1948);
nand U2051 (N_2051,N_1981,N_1997);
nor U2052 (N_2052,N_1989,N_1943);
or U2053 (N_2053,N_1906,N_1958);
xor U2054 (N_2054,N_1972,N_1961);
and U2055 (N_2055,N_1972,N_1907);
xor U2056 (N_2056,N_1942,N_1911);
nor U2057 (N_2057,N_1901,N_1936);
or U2058 (N_2058,N_1925,N_1931);
or U2059 (N_2059,N_1955,N_1994);
xor U2060 (N_2060,N_1980,N_1939);
nand U2061 (N_2061,N_1998,N_1957);
and U2062 (N_2062,N_1990,N_1913);
nor U2063 (N_2063,N_1979,N_1947);
xnor U2064 (N_2064,N_1923,N_1976);
and U2065 (N_2065,N_1981,N_1965);
xor U2066 (N_2066,N_1989,N_1976);
nor U2067 (N_2067,N_1924,N_1978);
nor U2068 (N_2068,N_1955,N_1963);
and U2069 (N_2069,N_1974,N_1971);
or U2070 (N_2070,N_1913,N_1984);
xor U2071 (N_2071,N_1950,N_1901);
and U2072 (N_2072,N_1915,N_1978);
nor U2073 (N_2073,N_1923,N_1972);
nor U2074 (N_2074,N_1957,N_1927);
nand U2075 (N_2075,N_1977,N_1989);
xor U2076 (N_2076,N_1984,N_1994);
xnor U2077 (N_2077,N_1944,N_1966);
xnor U2078 (N_2078,N_1968,N_1973);
nand U2079 (N_2079,N_1975,N_1920);
nor U2080 (N_2080,N_1980,N_1986);
or U2081 (N_2081,N_1945,N_1925);
and U2082 (N_2082,N_1980,N_1965);
or U2083 (N_2083,N_1927,N_1980);
or U2084 (N_2084,N_1902,N_1900);
xnor U2085 (N_2085,N_1998,N_1989);
and U2086 (N_2086,N_1955,N_1933);
and U2087 (N_2087,N_1920,N_1953);
and U2088 (N_2088,N_1994,N_1930);
and U2089 (N_2089,N_1991,N_1917);
or U2090 (N_2090,N_1953,N_1930);
nand U2091 (N_2091,N_1984,N_1948);
and U2092 (N_2092,N_1921,N_1910);
and U2093 (N_2093,N_1922,N_1926);
xnor U2094 (N_2094,N_1919,N_1943);
or U2095 (N_2095,N_1949,N_1912);
and U2096 (N_2096,N_1967,N_1920);
or U2097 (N_2097,N_1961,N_1943);
xnor U2098 (N_2098,N_1999,N_1900);
nor U2099 (N_2099,N_1918,N_1930);
xor U2100 (N_2100,N_2064,N_2009);
and U2101 (N_2101,N_2050,N_2062);
nor U2102 (N_2102,N_2065,N_2038);
nor U2103 (N_2103,N_2024,N_2082);
nand U2104 (N_2104,N_2011,N_2025);
and U2105 (N_2105,N_2077,N_2063);
and U2106 (N_2106,N_2083,N_2034);
or U2107 (N_2107,N_2066,N_2031);
xnor U2108 (N_2108,N_2061,N_2092);
and U2109 (N_2109,N_2069,N_2051);
nor U2110 (N_2110,N_2096,N_2014);
nor U2111 (N_2111,N_2093,N_2040);
nor U2112 (N_2112,N_2087,N_2013);
nor U2113 (N_2113,N_2052,N_2047);
and U2114 (N_2114,N_2070,N_2088);
nor U2115 (N_2115,N_2059,N_2078);
nand U2116 (N_2116,N_2023,N_2022);
or U2117 (N_2117,N_2039,N_2081);
nor U2118 (N_2118,N_2004,N_2091);
and U2119 (N_2119,N_2074,N_2029);
or U2120 (N_2120,N_2058,N_2057);
and U2121 (N_2121,N_2072,N_2002);
nand U2122 (N_2122,N_2003,N_2045);
nand U2123 (N_2123,N_2055,N_2033);
xnor U2124 (N_2124,N_2007,N_2071);
nor U2125 (N_2125,N_2042,N_2080);
xnor U2126 (N_2126,N_2067,N_2075);
nor U2127 (N_2127,N_2017,N_2056);
nand U2128 (N_2128,N_2068,N_2030);
or U2129 (N_2129,N_2041,N_2086);
xor U2130 (N_2130,N_2001,N_2018);
or U2131 (N_2131,N_2053,N_2073);
nand U2132 (N_2132,N_2019,N_2049);
or U2133 (N_2133,N_2016,N_2060);
and U2134 (N_2134,N_2028,N_2095);
xnor U2135 (N_2135,N_2043,N_2027);
nor U2136 (N_2136,N_2097,N_2085);
nand U2137 (N_2137,N_2000,N_2008);
nand U2138 (N_2138,N_2054,N_2046);
xnor U2139 (N_2139,N_2037,N_2021);
xnor U2140 (N_2140,N_2098,N_2048);
or U2141 (N_2141,N_2005,N_2076);
or U2142 (N_2142,N_2084,N_2012);
nor U2143 (N_2143,N_2089,N_2015);
or U2144 (N_2144,N_2026,N_2010);
or U2145 (N_2145,N_2035,N_2090);
nor U2146 (N_2146,N_2044,N_2032);
or U2147 (N_2147,N_2094,N_2079);
xnor U2148 (N_2148,N_2036,N_2006);
and U2149 (N_2149,N_2099,N_2020);
or U2150 (N_2150,N_2014,N_2045);
and U2151 (N_2151,N_2059,N_2077);
nor U2152 (N_2152,N_2085,N_2060);
nand U2153 (N_2153,N_2078,N_2012);
nor U2154 (N_2154,N_2039,N_2031);
and U2155 (N_2155,N_2043,N_2080);
nor U2156 (N_2156,N_2064,N_2067);
nand U2157 (N_2157,N_2038,N_2011);
nor U2158 (N_2158,N_2081,N_2066);
and U2159 (N_2159,N_2068,N_2011);
xnor U2160 (N_2160,N_2002,N_2061);
nand U2161 (N_2161,N_2054,N_2014);
and U2162 (N_2162,N_2036,N_2070);
xnor U2163 (N_2163,N_2088,N_2094);
nand U2164 (N_2164,N_2021,N_2066);
xnor U2165 (N_2165,N_2010,N_2008);
or U2166 (N_2166,N_2040,N_2028);
and U2167 (N_2167,N_2007,N_2040);
or U2168 (N_2168,N_2030,N_2002);
nand U2169 (N_2169,N_2045,N_2036);
and U2170 (N_2170,N_2016,N_2058);
or U2171 (N_2171,N_2045,N_2008);
nor U2172 (N_2172,N_2063,N_2086);
nand U2173 (N_2173,N_2094,N_2037);
or U2174 (N_2174,N_2053,N_2032);
and U2175 (N_2175,N_2002,N_2020);
xnor U2176 (N_2176,N_2029,N_2021);
or U2177 (N_2177,N_2013,N_2050);
or U2178 (N_2178,N_2023,N_2003);
and U2179 (N_2179,N_2038,N_2019);
and U2180 (N_2180,N_2072,N_2017);
nand U2181 (N_2181,N_2006,N_2078);
and U2182 (N_2182,N_2057,N_2082);
xor U2183 (N_2183,N_2085,N_2058);
nand U2184 (N_2184,N_2039,N_2093);
or U2185 (N_2185,N_2008,N_2075);
and U2186 (N_2186,N_2019,N_2092);
and U2187 (N_2187,N_2032,N_2045);
nor U2188 (N_2188,N_2008,N_2063);
xnor U2189 (N_2189,N_2006,N_2066);
or U2190 (N_2190,N_2096,N_2077);
nor U2191 (N_2191,N_2027,N_2058);
xor U2192 (N_2192,N_2009,N_2093);
xor U2193 (N_2193,N_2069,N_2098);
or U2194 (N_2194,N_2039,N_2094);
nand U2195 (N_2195,N_2011,N_2047);
or U2196 (N_2196,N_2060,N_2077);
or U2197 (N_2197,N_2014,N_2018);
and U2198 (N_2198,N_2004,N_2015);
and U2199 (N_2199,N_2092,N_2040);
nand U2200 (N_2200,N_2178,N_2179);
and U2201 (N_2201,N_2102,N_2115);
nand U2202 (N_2202,N_2167,N_2106);
xor U2203 (N_2203,N_2196,N_2198);
or U2204 (N_2204,N_2112,N_2156);
and U2205 (N_2205,N_2188,N_2187);
and U2206 (N_2206,N_2150,N_2158);
and U2207 (N_2207,N_2169,N_2133);
and U2208 (N_2208,N_2146,N_2171);
or U2209 (N_2209,N_2141,N_2173);
xor U2210 (N_2210,N_2137,N_2103);
and U2211 (N_2211,N_2101,N_2139);
xnor U2212 (N_2212,N_2125,N_2168);
nor U2213 (N_2213,N_2116,N_2136);
nand U2214 (N_2214,N_2134,N_2113);
or U2215 (N_2215,N_2160,N_2162);
or U2216 (N_2216,N_2174,N_2132);
xnor U2217 (N_2217,N_2184,N_2155);
nand U2218 (N_2218,N_2194,N_2157);
or U2219 (N_2219,N_2107,N_2143);
nor U2220 (N_2220,N_2170,N_2185);
nor U2221 (N_2221,N_2127,N_2109);
and U2222 (N_2222,N_2131,N_2135);
nor U2223 (N_2223,N_2190,N_2195);
xor U2224 (N_2224,N_2140,N_2197);
nand U2225 (N_2225,N_2186,N_2108);
or U2226 (N_2226,N_2183,N_2161);
and U2227 (N_2227,N_2189,N_2118);
nor U2228 (N_2228,N_2182,N_2121);
xor U2229 (N_2229,N_2119,N_2172);
xor U2230 (N_2230,N_2147,N_2154);
and U2231 (N_2231,N_2130,N_2151);
nand U2232 (N_2232,N_2110,N_2148);
or U2233 (N_2233,N_2153,N_2100);
nand U2234 (N_2234,N_2180,N_2181);
or U2235 (N_2235,N_2191,N_2163);
or U2236 (N_2236,N_2111,N_2105);
xnor U2237 (N_2237,N_2117,N_2104);
nor U2238 (N_2238,N_2164,N_2177);
or U2239 (N_2239,N_2152,N_2165);
nand U2240 (N_2240,N_2114,N_2192);
xnor U2241 (N_2241,N_2166,N_2142);
and U2242 (N_2242,N_2122,N_2138);
xnor U2243 (N_2243,N_2193,N_2123);
xor U2244 (N_2244,N_2126,N_2175);
nor U2245 (N_2245,N_2149,N_2124);
xnor U2246 (N_2246,N_2129,N_2159);
nand U2247 (N_2247,N_2145,N_2144);
nor U2248 (N_2248,N_2120,N_2199);
nand U2249 (N_2249,N_2176,N_2128);
nand U2250 (N_2250,N_2102,N_2101);
and U2251 (N_2251,N_2114,N_2179);
or U2252 (N_2252,N_2135,N_2117);
xor U2253 (N_2253,N_2146,N_2176);
xor U2254 (N_2254,N_2123,N_2172);
and U2255 (N_2255,N_2158,N_2120);
nand U2256 (N_2256,N_2192,N_2147);
xnor U2257 (N_2257,N_2113,N_2135);
xor U2258 (N_2258,N_2120,N_2150);
or U2259 (N_2259,N_2111,N_2152);
or U2260 (N_2260,N_2125,N_2104);
or U2261 (N_2261,N_2151,N_2119);
and U2262 (N_2262,N_2157,N_2154);
nand U2263 (N_2263,N_2175,N_2189);
or U2264 (N_2264,N_2103,N_2178);
nor U2265 (N_2265,N_2158,N_2179);
or U2266 (N_2266,N_2174,N_2112);
or U2267 (N_2267,N_2122,N_2136);
nor U2268 (N_2268,N_2195,N_2135);
or U2269 (N_2269,N_2103,N_2171);
and U2270 (N_2270,N_2151,N_2162);
and U2271 (N_2271,N_2157,N_2161);
xnor U2272 (N_2272,N_2109,N_2182);
xnor U2273 (N_2273,N_2191,N_2102);
nor U2274 (N_2274,N_2189,N_2143);
or U2275 (N_2275,N_2161,N_2160);
nor U2276 (N_2276,N_2122,N_2130);
and U2277 (N_2277,N_2115,N_2160);
nand U2278 (N_2278,N_2178,N_2104);
nor U2279 (N_2279,N_2128,N_2142);
nand U2280 (N_2280,N_2157,N_2153);
nor U2281 (N_2281,N_2186,N_2119);
xor U2282 (N_2282,N_2177,N_2187);
nor U2283 (N_2283,N_2155,N_2175);
or U2284 (N_2284,N_2156,N_2107);
or U2285 (N_2285,N_2179,N_2159);
nand U2286 (N_2286,N_2116,N_2161);
xnor U2287 (N_2287,N_2184,N_2106);
or U2288 (N_2288,N_2189,N_2185);
and U2289 (N_2289,N_2193,N_2196);
xnor U2290 (N_2290,N_2177,N_2123);
nor U2291 (N_2291,N_2113,N_2136);
xor U2292 (N_2292,N_2151,N_2107);
xnor U2293 (N_2293,N_2116,N_2159);
nand U2294 (N_2294,N_2164,N_2171);
and U2295 (N_2295,N_2168,N_2175);
and U2296 (N_2296,N_2145,N_2134);
xor U2297 (N_2297,N_2126,N_2149);
xor U2298 (N_2298,N_2154,N_2123);
xor U2299 (N_2299,N_2169,N_2187);
nand U2300 (N_2300,N_2239,N_2229);
nand U2301 (N_2301,N_2203,N_2227);
or U2302 (N_2302,N_2270,N_2210);
nand U2303 (N_2303,N_2258,N_2278);
or U2304 (N_2304,N_2286,N_2209);
xor U2305 (N_2305,N_2213,N_2262);
and U2306 (N_2306,N_2240,N_2241);
or U2307 (N_2307,N_2224,N_2218);
nand U2308 (N_2308,N_2291,N_2214);
or U2309 (N_2309,N_2280,N_2211);
nand U2310 (N_2310,N_2261,N_2207);
nand U2311 (N_2311,N_2294,N_2265);
or U2312 (N_2312,N_2237,N_2269);
nor U2313 (N_2313,N_2230,N_2245);
and U2314 (N_2314,N_2281,N_2297);
xnor U2315 (N_2315,N_2216,N_2250);
nor U2316 (N_2316,N_2290,N_2244);
xnor U2317 (N_2317,N_2263,N_2220);
and U2318 (N_2318,N_2212,N_2264);
or U2319 (N_2319,N_2200,N_2228);
nand U2320 (N_2320,N_2298,N_2202);
nor U2321 (N_2321,N_2282,N_2201);
and U2322 (N_2322,N_2232,N_2231);
nor U2323 (N_2323,N_2287,N_2266);
xor U2324 (N_2324,N_2277,N_2288);
xor U2325 (N_2325,N_2293,N_2275);
and U2326 (N_2326,N_2226,N_2222);
or U2327 (N_2327,N_2254,N_2252);
nor U2328 (N_2328,N_2238,N_2233);
nor U2329 (N_2329,N_2219,N_2296);
xnor U2330 (N_2330,N_2247,N_2208);
nand U2331 (N_2331,N_2268,N_2279);
nand U2332 (N_2332,N_2221,N_2295);
and U2333 (N_2333,N_2251,N_2248);
and U2334 (N_2334,N_2215,N_2223);
and U2335 (N_2335,N_2246,N_2284);
or U2336 (N_2336,N_2256,N_2236);
or U2337 (N_2337,N_2283,N_2235);
xor U2338 (N_2338,N_2259,N_2205);
nor U2339 (N_2339,N_2225,N_2255);
nand U2340 (N_2340,N_2243,N_2267);
nor U2341 (N_2341,N_2206,N_2271);
and U2342 (N_2342,N_2272,N_2204);
and U2343 (N_2343,N_2260,N_2217);
nand U2344 (N_2344,N_2249,N_2242);
xor U2345 (N_2345,N_2289,N_2292);
nand U2346 (N_2346,N_2276,N_2274);
or U2347 (N_2347,N_2257,N_2253);
or U2348 (N_2348,N_2273,N_2299);
and U2349 (N_2349,N_2285,N_2234);
xnor U2350 (N_2350,N_2254,N_2231);
or U2351 (N_2351,N_2246,N_2288);
and U2352 (N_2352,N_2291,N_2260);
nor U2353 (N_2353,N_2256,N_2207);
and U2354 (N_2354,N_2287,N_2204);
nor U2355 (N_2355,N_2269,N_2238);
xnor U2356 (N_2356,N_2239,N_2231);
nand U2357 (N_2357,N_2237,N_2294);
nand U2358 (N_2358,N_2298,N_2243);
or U2359 (N_2359,N_2213,N_2238);
nand U2360 (N_2360,N_2222,N_2255);
nand U2361 (N_2361,N_2213,N_2283);
nand U2362 (N_2362,N_2269,N_2231);
nand U2363 (N_2363,N_2286,N_2234);
nor U2364 (N_2364,N_2205,N_2298);
nand U2365 (N_2365,N_2272,N_2275);
xnor U2366 (N_2366,N_2206,N_2248);
nor U2367 (N_2367,N_2262,N_2232);
nand U2368 (N_2368,N_2256,N_2204);
nand U2369 (N_2369,N_2227,N_2260);
xnor U2370 (N_2370,N_2253,N_2228);
xnor U2371 (N_2371,N_2262,N_2212);
or U2372 (N_2372,N_2289,N_2284);
and U2373 (N_2373,N_2207,N_2279);
and U2374 (N_2374,N_2261,N_2234);
xnor U2375 (N_2375,N_2210,N_2229);
and U2376 (N_2376,N_2248,N_2290);
nor U2377 (N_2377,N_2250,N_2215);
nor U2378 (N_2378,N_2296,N_2211);
or U2379 (N_2379,N_2233,N_2263);
nor U2380 (N_2380,N_2271,N_2297);
nor U2381 (N_2381,N_2292,N_2265);
xnor U2382 (N_2382,N_2273,N_2296);
or U2383 (N_2383,N_2260,N_2234);
nand U2384 (N_2384,N_2268,N_2241);
and U2385 (N_2385,N_2237,N_2256);
xnor U2386 (N_2386,N_2208,N_2241);
nand U2387 (N_2387,N_2216,N_2253);
and U2388 (N_2388,N_2227,N_2202);
nor U2389 (N_2389,N_2226,N_2248);
xnor U2390 (N_2390,N_2212,N_2284);
nand U2391 (N_2391,N_2273,N_2234);
nand U2392 (N_2392,N_2291,N_2233);
and U2393 (N_2393,N_2230,N_2228);
or U2394 (N_2394,N_2225,N_2260);
xor U2395 (N_2395,N_2225,N_2233);
and U2396 (N_2396,N_2273,N_2229);
nand U2397 (N_2397,N_2280,N_2224);
nand U2398 (N_2398,N_2239,N_2205);
nor U2399 (N_2399,N_2239,N_2271);
or U2400 (N_2400,N_2379,N_2354);
nand U2401 (N_2401,N_2361,N_2306);
nand U2402 (N_2402,N_2357,N_2355);
and U2403 (N_2403,N_2352,N_2326);
nor U2404 (N_2404,N_2387,N_2347);
nor U2405 (N_2405,N_2329,N_2315);
or U2406 (N_2406,N_2317,N_2338);
nand U2407 (N_2407,N_2399,N_2324);
or U2408 (N_2408,N_2381,N_2301);
nor U2409 (N_2409,N_2363,N_2328);
nand U2410 (N_2410,N_2382,N_2373);
xor U2411 (N_2411,N_2318,N_2321);
nor U2412 (N_2412,N_2376,N_2353);
nor U2413 (N_2413,N_2325,N_2383);
or U2414 (N_2414,N_2307,N_2358);
xor U2415 (N_2415,N_2345,N_2367);
and U2416 (N_2416,N_2330,N_2341);
nor U2417 (N_2417,N_2384,N_2333);
nor U2418 (N_2418,N_2300,N_2336);
xor U2419 (N_2419,N_2389,N_2375);
or U2420 (N_2420,N_2346,N_2393);
nor U2421 (N_2421,N_2377,N_2343);
nand U2422 (N_2422,N_2335,N_2312);
or U2423 (N_2423,N_2316,N_2348);
nor U2424 (N_2424,N_2395,N_2327);
nand U2425 (N_2425,N_2304,N_2380);
or U2426 (N_2426,N_2308,N_2388);
nor U2427 (N_2427,N_2344,N_2391);
and U2428 (N_2428,N_2392,N_2372);
and U2429 (N_2429,N_2356,N_2390);
nor U2430 (N_2430,N_2337,N_2351);
or U2431 (N_2431,N_2310,N_2374);
nor U2432 (N_2432,N_2350,N_2334);
and U2433 (N_2433,N_2360,N_2386);
and U2434 (N_2434,N_2369,N_2362);
and U2435 (N_2435,N_2359,N_2311);
or U2436 (N_2436,N_2323,N_2340);
nand U2437 (N_2437,N_2309,N_2370);
nor U2438 (N_2438,N_2303,N_2368);
nand U2439 (N_2439,N_2365,N_2339);
xor U2440 (N_2440,N_2342,N_2302);
and U2441 (N_2441,N_2332,N_2398);
or U2442 (N_2442,N_2305,N_2349);
and U2443 (N_2443,N_2378,N_2371);
xnor U2444 (N_2444,N_2385,N_2320);
xor U2445 (N_2445,N_2331,N_2366);
or U2446 (N_2446,N_2322,N_2313);
and U2447 (N_2447,N_2394,N_2364);
xor U2448 (N_2448,N_2319,N_2396);
or U2449 (N_2449,N_2397,N_2314);
nor U2450 (N_2450,N_2379,N_2322);
xnor U2451 (N_2451,N_2335,N_2385);
xor U2452 (N_2452,N_2377,N_2333);
or U2453 (N_2453,N_2355,N_2368);
nand U2454 (N_2454,N_2344,N_2334);
and U2455 (N_2455,N_2313,N_2367);
or U2456 (N_2456,N_2389,N_2360);
xor U2457 (N_2457,N_2355,N_2323);
and U2458 (N_2458,N_2389,N_2337);
nand U2459 (N_2459,N_2324,N_2398);
xnor U2460 (N_2460,N_2344,N_2312);
and U2461 (N_2461,N_2331,N_2321);
or U2462 (N_2462,N_2315,N_2395);
and U2463 (N_2463,N_2317,N_2383);
or U2464 (N_2464,N_2377,N_2331);
and U2465 (N_2465,N_2380,N_2359);
nor U2466 (N_2466,N_2367,N_2361);
nand U2467 (N_2467,N_2381,N_2396);
nand U2468 (N_2468,N_2379,N_2302);
nand U2469 (N_2469,N_2356,N_2351);
nand U2470 (N_2470,N_2355,N_2393);
nand U2471 (N_2471,N_2313,N_2324);
and U2472 (N_2472,N_2330,N_2325);
xor U2473 (N_2473,N_2355,N_2375);
or U2474 (N_2474,N_2337,N_2309);
xnor U2475 (N_2475,N_2369,N_2340);
nand U2476 (N_2476,N_2327,N_2306);
nor U2477 (N_2477,N_2356,N_2363);
nor U2478 (N_2478,N_2381,N_2320);
nand U2479 (N_2479,N_2366,N_2336);
nand U2480 (N_2480,N_2376,N_2394);
nor U2481 (N_2481,N_2352,N_2335);
xor U2482 (N_2482,N_2318,N_2322);
or U2483 (N_2483,N_2366,N_2370);
or U2484 (N_2484,N_2303,N_2387);
nand U2485 (N_2485,N_2314,N_2396);
xnor U2486 (N_2486,N_2315,N_2369);
nor U2487 (N_2487,N_2399,N_2336);
nand U2488 (N_2488,N_2374,N_2361);
nand U2489 (N_2489,N_2365,N_2314);
or U2490 (N_2490,N_2395,N_2340);
nand U2491 (N_2491,N_2388,N_2311);
and U2492 (N_2492,N_2353,N_2393);
xor U2493 (N_2493,N_2339,N_2374);
and U2494 (N_2494,N_2354,N_2368);
nand U2495 (N_2495,N_2353,N_2355);
and U2496 (N_2496,N_2332,N_2318);
nor U2497 (N_2497,N_2335,N_2394);
xor U2498 (N_2498,N_2369,N_2322);
nand U2499 (N_2499,N_2368,N_2328);
or U2500 (N_2500,N_2442,N_2497);
xor U2501 (N_2501,N_2485,N_2447);
xnor U2502 (N_2502,N_2448,N_2486);
nand U2503 (N_2503,N_2478,N_2483);
xnor U2504 (N_2504,N_2434,N_2401);
or U2505 (N_2505,N_2498,N_2410);
nand U2506 (N_2506,N_2496,N_2494);
and U2507 (N_2507,N_2490,N_2450);
nand U2508 (N_2508,N_2418,N_2441);
and U2509 (N_2509,N_2461,N_2423);
nand U2510 (N_2510,N_2403,N_2404);
xor U2511 (N_2511,N_2428,N_2471);
nand U2512 (N_2512,N_2430,N_2433);
and U2513 (N_2513,N_2451,N_2472);
xnor U2514 (N_2514,N_2446,N_2405);
xnor U2515 (N_2515,N_2409,N_2402);
nor U2516 (N_2516,N_2437,N_2466);
xor U2517 (N_2517,N_2462,N_2422);
nor U2518 (N_2518,N_2468,N_2495);
or U2519 (N_2519,N_2477,N_2426);
nor U2520 (N_2520,N_2476,N_2419);
or U2521 (N_2521,N_2411,N_2470);
nor U2522 (N_2522,N_2439,N_2481);
nand U2523 (N_2523,N_2489,N_2436);
xnor U2524 (N_2524,N_2453,N_2488);
xnor U2525 (N_2525,N_2444,N_2449);
and U2526 (N_2526,N_2473,N_2458);
and U2527 (N_2527,N_2456,N_2491);
or U2528 (N_2528,N_2414,N_2424);
or U2529 (N_2529,N_2420,N_2499);
xnor U2530 (N_2530,N_2400,N_2435);
and U2531 (N_2531,N_2432,N_2454);
or U2532 (N_2532,N_2429,N_2455);
xor U2533 (N_2533,N_2438,N_2459);
and U2534 (N_2534,N_2480,N_2475);
nand U2535 (N_2535,N_2415,N_2487);
and U2536 (N_2536,N_2427,N_2452);
xnor U2537 (N_2537,N_2406,N_2445);
nand U2538 (N_2538,N_2407,N_2460);
and U2539 (N_2539,N_2440,N_2464);
nand U2540 (N_2540,N_2431,N_2425);
and U2541 (N_2541,N_2443,N_2412);
nor U2542 (N_2542,N_2408,N_2463);
nand U2543 (N_2543,N_2467,N_2457);
nand U2544 (N_2544,N_2413,N_2492);
nor U2545 (N_2545,N_2482,N_2416);
or U2546 (N_2546,N_2484,N_2469);
and U2547 (N_2547,N_2465,N_2479);
xor U2548 (N_2548,N_2417,N_2421);
nor U2549 (N_2549,N_2474,N_2493);
nand U2550 (N_2550,N_2445,N_2425);
and U2551 (N_2551,N_2403,N_2461);
nand U2552 (N_2552,N_2467,N_2419);
and U2553 (N_2553,N_2497,N_2472);
nor U2554 (N_2554,N_2443,N_2461);
or U2555 (N_2555,N_2423,N_2442);
or U2556 (N_2556,N_2490,N_2436);
and U2557 (N_2557,N_2412,N_2418);
xor U2558 (N_2558,N_2436,N_2446);
nor U2559 (N_2559,N_2489,N_2461);
xor U2560 (N_2560,N_2400,N_2483);
and U2561 (N_2561,N_2442,N_2419);
xnor U2562 (N_2562,N_2483,N_2440);
xnor U2563 (N_2563,N_2490,N_2403);
nor U2564 (N_2564,N_2437,N_2485);
nor U2565 (N_2565,N_2492,N_2434);
nor U2566 (N_2566,N_2486,N_2445);
or U2567 (N_2567,N_2410,N_2420);
nand U2568 (N_2568,N_2441,N_2482);
and U2569 (N_2569,N_2410,N_2496);
xnor U2570 (N_2570,N_2473,N_2419);
nor U2571 (N_2571,N_2456,N_2437);
xor U2572 (N_2572,N_2489,N_2427);
nand U2573 (N_2573,N_2430,N_2467);
nand U2574 (N_2574,N_2436,N_2481);
xor U2575 (N_2575,N_2469,N_2438);
nand U2576 (N_2576,N_2437,N_2400);
nand U2577 (N_2577,N_2454,N_2484);
nand U2578 (N_2578,N_2407,N_2404);
and U2579 (N_2579,N_2455,N_2432);
nand U2580 (N_2580,N_2467,N_2426);
xnor U2581 (N_2581,N_2454,N_2475);
nand U2582 (N_2582,N_2445,N_2485);
nor U2583 (N_2583,N_2427,N_2421);
and U2584 (N_2584,N_2457,N_2405);
or U2585 (N_2585,N_2416,N_2461);
nand U2586 (N_2586,N_2473,N_2415);
xnor U2587 (N_2587,N_2405,N_2420);
and U2588 (N_2588,N_2449,N_2456);
nand U2589 (N_2589,N_2474,N_2497);
and U2590 (N_2590,N_2402,N_2471);
or U2591 (N_2591,N_2481,N_2443);
nor U2592 (N_2592,N_2424,N_2429);
xnor U2593 (N_2593,N_2480,N_2419);
nand U2594 (N_2594,N_2476,N_2439);
nand U2595 (N_2595,N_2474,N_2478);
and U2596 (N_2596,N_2493,N_2472);
or U2597 (N_2597,N_2468,N_2432);
or U2598 (N_2598,N_2494,N_2403);
nor U2599 (N_2599,N_2417,N_2434);
nor U2600 (N_2600,N_2591,N_2577);
xor U2601 (N_2601,N_2540,N_2574);
nand U2602 (N_2602,N_2500,N_2513);
and U2603 (N_2603,N_2536,N_2533);
nand U2604 (N_2604,N_2537,N_2521);
nand U2605 (N_2605,N_2572,N_2588);
xnor U2606 (N_2606,N_2516,N_2555);
and U2607 (N_2607,N_2598,N_2584);
or U2608 (N_2608,N_2597,N_2561);
and U2609 (N_2609,N_2520,N_2594);
or U2610 (N_2610,N_2586,N_2557);
xor U2611 (N_2611,N_2539,N_2587);
or U2612 (N_2612,N_2592,N_2535);
or U2613 (N_2613,N_2599,N_2563);
nand U2614 (N_2614,N_2504,N_2501);
nand U2615 (N_2615,N_2548,N_2567);
nand U2616 (N_2616,N_2559,N_2525);
xor U2617 (N_2617,N_2511,N_2579);
or U2618 (N_2618,N_2560,N_2576);
nand U2619 (N_2619,N_2510,N_2509);
nor U2620 (N_2620,N_2580,N_2523);
and U2621 (N_2621,N_2570,N_2512);
and U2622 (N_2622,N_2519,N_2590);
or U2623 (N_2623,N_2527,N_2552);
xnor U2624 (N_2624,N_2514,N_2564);
nor U2625 (N_2625,N_2551,N_2569);
nor U2626 (N_2626,N_2554,N_2573);
nor U2627 (N_2627,N_2506,N_2524);
nor U2628 (N_2628,N_2502,N_2532);
nor U2629 (N_2629,N_2589,N_2581);
nor U2630 (N_2630,N_2582,N_2522);
or U2631 (N_2631,N_2541,N_2566);
or U2632 (N_2632,N_2547,N_2507);
and U2633 (N_2633,N_2517,N_2528);
or U2634 (N_2634,N_2593,N_2545);
nand U2635 (N_2635,N_2550,N_2553);
or U2636 (N_2636,N_2565,N_2558);
xor U2637 (N_2637,N_2534,N_2531);
xor U2638 (N_2638,N_2562,N_2503);
xnor U2639 (N_2639,N_2578,N_2583);
nand U2640 (N_2640,N_2596,N_2505);
xor U2641 (N_2641,N_2556,N_2530);
xor U2642 (N_2642,N_2518,N_2585);
nand U2643 (N_2643,N_2568,N_2549);
nand U2644 (N_2644,N_2526,N_2571);
nor U2645 (N_2645,N_2546,N_2543);
nor U2646 (N_2646,N_2542,N_2575);
nand U2647 (N_2647,N_2515,N_2544);
nand U2648 (N_2648,N_2508,N_2529);
and U2649 (N_2649,N_2538,N_2595);
nor U2650 (N_2650,N_2540,N_2514);
xor U2651 (N_2651,N_2586,N_2539);
xor U2652 (N_2652,N_2504,N_2561);
and U2653 (N_2653,N_2515,N_2564);
xnor U2654 (N_2654,N_2541,N_2568);
and U2655 (N_2655,N_2540,N_2527);
xnor U2656 (N_2656,N_2543,N_2548);
nand U2657 (N_2657,N_2594,N_2593);
nand U2658 (N_2658,N_2555,N_2500);
and U2659 (N_2659,N_2588,N_2565);
nand U2660 (N_2660,N_2576,N_2523);
xor U2661 (N_2661,N_2554,N_2558);
xnor U2662 (N_2662,N_2545,N_2505);
nor U2663 (N_2663,N_2548,N_2532);
xor U2664 (N_2664,N_2503,N_2513);
nand U2665 (N_2665,N_2525,N_2530);
and U2666 (N_2666,N_2573,N_2592);
nor U2667 (N_2667,N_2535,N_2547);
xor U2668 (N_2668,N_2583,N_2505);
nor U2669 (N_2669,N_2500,N_2588);
nor U2670 (N_2670,N_2596,N_2562);
or U2671 (N_2671,N_2578,N_2509);
or U2672 (N_2672,N_2541,N_2559);
or U2673 (N_2673,N_2552,N_2504);
nand U2674 (N_2674,N_2526,N_2569);
xor U2675 (N_2675,N_2598,N_2504);
nor U2676 (N_2676,N_2517,N_2500);
or U2677 (N_2677,N_2547,N_2512);
and U2678 (N_2678,N_2541,N_2550);
and U2679 (N_2679,N_2560,N_2553);
nor U2680 (N_2680,N_2512,N_2553);
nand U2681 (N_2681,N_2562,N_2513);
nand U2682 (N_2682,N_2586,N_2566);
or U2683 (N_2683,N_2539,N_2559);
or U2684 (N_2684,N_2557,N_2589);
xor U2685 (N_2685,N_2534,N_2552);
and U2686 (N_2686,N_2532,N_2550);
nand U2687 (N_2687,N_2531,N_2599);
nor U2688 (N_2688,N_2582,N_2535);
and U2689 (N_2689,N_2510,N_2535);
xnor U2690 (N_2690,N_2525,N_2546);
nor U2691 (N_2691,N_2541,N_2599);
or U2692 (N_2692,N_2519,N_2522);
nand U2693 (N_2693,N_2584,N_2517);
and U2694 (N_2694,N_2557,N_2534);
and U2695 (N_2695,N_2575,N_2586);
xnor U2696 (N_2696,N_2501,N_2561);
or U2697 (N_2697,N_2569,N_2560);
nand U2698 (N_2698,N_2523,N_2557);
or U2699 (N_2699,N_2599,N_2522);
or U2700 (N_2700,N_2690,N_2642);
nor U2701 (N_2701,N_2617,N_2626);
nand U2702 (N_2702,N_2687,N_2644);
and U2703 (N_2703,N_2654,N_2600);
and U2704 (N_2704,N_2618,N_2691);
nand U2705 (N_2705,N_2609,N_2652);
nand U2706 (N_2706,N_2605,N_2657);
nor U2707 (N_2707,N_2624,N_2673);
and U2708 (N_2708,N_2662,N_2663);
nand U2709 (N_2709,N_2631,N_2655);
or U2710 (N_2710,N_2683,N_2668);
xor U2711 (N_2711,N_2613,N_2692);
nand U2712 (N_2712,N_2675,N_2679);
nand U2713 (N_2713,N_2620,N_2603);
or U2714 (N_2714,N_2627,N_2659);
nand U2715 (N_2715,N_2608,N_2614);
or U2716 (N_2716,N_2688,N_2639);
and U2717 (N_2717,N_2686,N_2638);
nor U2718 (N_2718,N_2623,N_2622);
and U2719 (N_2719,N_2672,N_2602);
or U2720 (N_2720,N_2615,N_2640);
nor U2721 (N_2721,N_2666,N_2619);
or U2722 (N_2722,N_2610,N_2669);
nand U2723 (N_2723,N_2607,N_2693);
or U2724 (N_2724,N_2635,N_2604);
nor U2725 (N_2725,N_2697,N_2696);
xnor U2726 (N_2726,N_2625,N_2653);
and U2727 (N_2727,N_2648,N_2606);
xnor U2728 (N_2728,N_2689,N_2634);
xor U2729 (N_2729,N_2612,N_2630);
xor U2730 (N_2730,N_2660,N_2636);
or U2731 (N_2731,N_2694,N_2671);
nand U2732 (N_2732,N_2680,N_2682);
and U2733 (N_2733,N_2658,N_2678);
nand U2734 (N_2734,N_2685,N_2611);
and U2735 (N_2735,N_2628,N_2645);
and U2736 (N_2736,N_2656,N_2665);
or U2737 (N_2737,N_2633,N_2698);
and U2738 (N_2738,N_2684,N_2661);
and U2739 (N_2739,N_2681,N_2651);
nand U2740 (N_2740,N_2664,N_2650);
nand U2741 (N_2741,N_2676,N_2699);
nand U2742 (N_2742,N_2695,N_2621);
xor U2743 (N_2743,N_2616,N_2641);
nand U2744 (N_2744,N_2677,N_2649);
and U2745 (N_2745,N_2674,N_2643);
nand U2746 (N_2746,N_2667,N_2629);
nor U2747 (N_2747,N_2647,N_2601);
nor U2748 (N_2748,N_2632,N_2637);
and U2749 (N_2749,N_2670,N_2646);
nand U2750 (N_2750,N_2637,N_2688);
and U2751 (N_2751,N_2668,N_2682);
or U2752 (N_2752,N_2683,N_2697);
or U2753 (N_2753,N_2644,N_2621);
nor U2754 (N_2754,N_2667,N_2621);
xor U2755 (N_2755,N_2638,N_2609);
xnor U2756 (N_2756,N_2672,N_2677);
nand U2757 (N_2757,N_2619,N_2617);
nor U2758 (N_2758,N_2682,N_2692);
nand U2759 (N_2759,N_2625,N_2663);
nor U2760 (N_2760,N_2636,N_2678);
nor U2761 (N_2761,N_2663,N_2651);
or U2762 (N_2762,N_2639,N_2647);
and U2763 (N_2763,N_2698,N_2673);
nand U2764 (N_2764,N_2667,N_2633);
or U2765 (N_2765,N_2693,N_2656);
or U2766 (N_2766,N_2628,N_2658);
nor U2767 (N_2767,N_2680,N_2628);
nor U2768 (N_2768,N_2640,N_2648);
and U2769 (N_2769,N_2654,N_2674);
and U2770 (N_2770,N_2654,N_2664);
xor U2771 (N_2771,N_2603,N_2640);
xnor U2772 (N_2772,N_2634,N_2622);
nand U2773 (N_2773,N_2635,N_2687);
and U2774 (N_2774,N_2617,N_2677);
xor U2775 (N_2775,N_2650,N_2619);
xor U2776 (N_2776,N_2676,N_2621);
xor U2777 (N_2777,N_2690,N_2639);
nor U2778 (N_2778,N_2616,N_2653);
nand U2779 (N_2779,N_2674,N_2653);
and U2780 (N_2780,N_2695,N_2693);
or U2781 (N_2781,N_2607,N_2615);
and U2782 (N_2782,N_2645,N_2627);
nor U2783 (N_2783,N_2691,N_2668);
nand U2784 (N_2784,N_2683,N_2619);
and U2785 (N_2785,N_2652,N_2699);
nand U2786 (N_2786,N_2608,N_2684);
nor U2787 (N_2787,N_2660,N_2664);
nor U2788 (N_2788,N_2686,N_2658);
xor U2789 (N_2789,N_2626,N_2606);
nor U2790 (N_2790,N_2696,N_2626);
or U2791 (N_2791,N_2601,N_2657);
or U2792 (N_2792,N_2626,N_2622);
or U2793 (N_2793,N_2657,N_2637);
xnor U2794 (N_2794,N_2646,N_2693);
and U2795 (N_2795,N_2610,N_2661);
and U2796 (N_2796,N_2616,N_2672);
nor U2797 (N_2797,N_2608,N_2644);
nand U2798 (N_2798,N_2603,N_2660);
nor U2799 (N_2799,N_2688,N_2684);
xnor U2800 (N_2800,N_2724,N_2793);
nand U2801 (N_2801,N_2788,N_2733);
nand U2802 (N_2802,N_2741,N_2719);
nand U2803 (N_2803,N_2753,N_2762);
or U2804 (N_2804,N_2728,N_2730);
or U2805 (N_2805,N_2744,N_2766);
nor U2806 (N_2806,N_2713,N_2736);
and U2807 (N_2807,N_2721,N_2740);
nand U2808 (N_2808,N_2745,N_2764);
nand U2809 (N_2809,N_2769,N_2742);
or U2810 (N_2810,N_2726,N_2770);
xnor U2811 (N_2811,N_2774,N_2795);
or U2812 (N_2812,N_2761,N_2789);
xnor U2813 (N_2813,N_2747,N_2752);
xnor U2814 (N_2814,N_2706,N_2751);
or U2815 (N_2815,N_2755,N_2715);
and U2816 (N_2816,N_2743,N_2796);
and U2817 (N_2817,N_2708,N_2702);
xor U2818 (N_2818,N_2705,N_2704);
and U2819 (N_2819,N_2799,N_2739);
and U2820 (N_2820,N_2716,N_2738);
and U2821 (N_2821,N_2717,N_2765);
and U2822 (N_2822,N_2758,N_2776);
nor U2823 (N_2823,N_2750,N_2777);
xor U2824 (N_2824,N_2783,N_2798);
nand U2825 (N_2825,N_2757,N_2781);
or U2826 (N_2826,N_2768,N_2773);
or U2827 (N_2827,N_2729,N_2703);
xnor U2828 (N_2828,N_2707,N_2787);
nor U2829 (N_2829,N_2797,N_2732);
xor U2830 (N_2830,N_2771,N_2714);
xor U2831 (N_2831,N_2756,N_2701);
xor U2832 (N_2832,N_2709,N_2737);
nand U2833 (N_2833,N_2794,N_2720);
nor U2834 (N_2834,N_2767,N_2711);
xor U2835 (N_2835,N_2725,N_2727);
and U2836 (N_2836,N_2722,N_2700);
nand U2837 (N_2837,N_2790,N_2760);
nor U2838 (N_2838,N_2748,N_2731);
and U2839 (N_2839,N_2763,N_2772);
nor U2840 (N_2840,N_2723,N_2746);
and U2841 (N_2841,N_2779,N_2712);
or U2842 (N_2842,N_2735,N_2782);
nand U2843 (N_2843,N_2778,N_2749);
or U2844 (N_2844,N_2792,N_2775);
nor U2845 (N_2845,N_2784,N_2718);
xnor U2846 (N_2846,N_2759,N_2780);
or U2847 (N_2847,N_2791,N_2734);
nand U2848 (N_2848,N_2785,N_2710);
and U2849 (N_2849,N_2754,N_2786);
nor U2850 (N_2850,N_2775,N_2772);
nor U2851 (N_2851,N_2771,N_2783);
xnor U2852 (N_2852,N_2795,N_2758);
or U2853 (N_2853,N_2715,N_2796);
and U2854 (N_2854,N_2785,N_2731);
xnor U2855 (N_2855,N_2744,N_2789);
xnor U2856 (N_2856,N_2793,N_2774);
nor U2857 (N_2857,N_2724,N_2706);
nand U2858 (N_2858,N_2768,N_2729);
xor U2859 (N_2859,N_2740,N_2739);
xnor U2860 (N_2860,N_2798,N_2758);
or U2861 (N_2861,N_2713,N_2703);
or U2862 (N_2862,N_2798,N_2750);
and U2863 (N_2863,N_2739,N_2708);
nand U2864 (N_2864,N_2774,N_2755);
nand U2865 (N_2865,N_2702,N_2738);
and U2866 (N_2866,N_2780,N_2733);
nor U2867 (N_2867,N_2757,N_2744);
or U2868 (N_2868,N_2708,N_2758);
nand U2869 (N_2869,N_2725,N_2707);
or U2870 (N_2870,N_2704,N_2709);
and U2871 (N_2871,N_2735,N_2785);
nor U2872 (N_2872,N_2718,N_2755);
nand U2873 (N_2873,N_2727,N_2757);
xnor U2874 (N_2874,N_2747,N_2734);
or U2875 (N_2875,N_2765,N_2721);
and U2876 (N_2876,N_2769,N_2739);
nand U2877 (N_2877,N_2777,N_2773);
or U2878 (N_2878,N_2715,N_2788);
xor U2879 (N_2879,N_2783,N_2724);
nand U2880 (N_2880,N_2749,N_2770);
nor U2881 (N_2881,N_2736,N_2768);
and U2882 (N_2882,N_2726,N_2702);
nor U2883 (N_2883,N_2773,N_2730);
and U2884 (N_2884,N_2772,N_2702);
nand U2885 (N_2885,N_2718,N_2771);
nor U2886 (N_2886,N_2765,N_2781);
nand U2887 (N_2887,N_2738,N_2701);
or U2888 (N_2888,N_2746,N_2721);
or U2889 (N_2889,N_2727,N_2783);
or U2890 (N_2890,N_2705,N_2753);
and U2891 (N_2891,N_2717,N_2758);
nand U2892 (N_2892,N_2748,N_2777);
xor U2893 (N_2893,N_2757,N_2749);
or U2894 (N_2894,N_2724,N_2770);
nand U2895 (N_2895,N_2730,N_2726);
or U2896 (N_2896,N_2718,N_2781);
or U2897 (N_2897,N_2742,N_2799);
nor U2898 (N_2898,N_2793,N_2797);
and U2899 (N_2899,N_2790,N_2763);
xnor U2900 (N_2900,N_2874,N_2898);
xor U2901 (N_2901,N_2861,N_2825);
xnor U2902 (N_2902,N_2802,N_2884);
and U2903 (N_2903,N_2896,N_2869);
xnor U2904 (N_2904,N_2834,N_2819);
nor U2905 (N_2905,N_2879,N_2870);
nand U2906 (N_2906,N_2816,N_2892);
nor U2907 (N_2907,N_2863,N_2860);
xnor U2908 (N_2908,N_2831,N_2810);
nor U2909 (N_2909,N_2803,N_2865);
and U2910 (N_2910,N_2844,N_2826);
nand U2911 (N_2911,N_2823,N_2885);
xnor U2912 (N_2912,N_2817,N_2837);
nand U2913 (N_2913,N_2897,N_2830);
xnor U2914 (N_2914,N_2887,N_2846);
nand U2915 (N_2915,N_2838,N_2873);
or U2916 (N_2916,N_2822,N_2852);
or U2917 (N_2917,N_2849,N_2848);
or U2918 (N_2918,N_2818,N_2836);
or U2919 (N_2919,N_2877,N_2842);
and U2920 (N_2920,N_2883,N_2805);
nor U2921 (N_2921,N_2856,N_2827);
xor U2922 (N_2922,N_2881,N_2821);
and U2923 (N_2923,N_2807,N_2886);
or U2924 (N_2924,N_2895,N_2813);
and U2925 (N_2925,N_2840,N_2845);
nor U2926 (N_2926,N_2857,N_2882);
or U2927 (N_2927,N_2811,N_2862);
nor U2928 (N_2928,N_2875,N_2893);
or U2929 (N_2929,N_2858,N_2829);
nor U2930 (N_2930,N_2894,N_2828);
xor U2931 (N_2931,N_2809,N_2878);
and U2932 (N_2932,N_2800,N_2815);
nand U2933 (N_2933,N_2853,N_2839);
nor U2934 (N_2934,N_2872,N_2880);
or U2935 (N_2935,N_2843,N_2899);
or U2936 (N_2936,N_2851,N_2871);
xnor U2937 (N_2937,N_2876,N_2806);
nand U2938 (N_2938,N_2841,N_2890);
xnor U2939 (N_2939,N_2864,N_2854);
nand U2940 (N_2940,N_2867,N_2847);
nand U2941 (N_2941,N_2859,N_2888);
nand U2942 (N_2942,N_2804,N_2808);
nor U2943 (N_2943,N_2889,N_2868);
nand U2944 (N_2944,N_2835,N_2812);
nand U2945 (N_2945,N_2824,N_2832);
nor U2946 (N_2946,N_2855,N_2866);
xnor U2947 (N_2947,N_2814,N_2833);
xor U2948 (N_2948,N_2891,N_2801);
xor U2949 (N_2949,N_2850,N_2820);
and U2950 (N_2950,N_2813,N_2897);
and U2951 (N_2951,N_2819,N_2825);
nand U2952 (N_2952,N_2874,N_2804);
nor U2953 (N_2953,N_2839,N_2812);
or U2954 (N_2954,N_2814,N_2864);
xor U2955 (N_2955,N_2837,N_2844);
and U2956 (N_2956,N_2847,N_2826);
xnor U2957 (N_2957,N_2840,N_2892);
or U2958 (N_2958,N_2844,N_2818);
or U2959 (N_2959,N_2843,N_2814);
xnor U2960 (N_2960,N_2830,N_2856);
or U2961 (N_2961,N_2835,N_2832);
xor U2962 (N_2962,N_2873,N_2894);
nor U2963 (N_2963,N_2865,N_2869);
or U2964 (N_2964,N_2877,N_2821);
and U2965 (N_2965,N_2893,N_2829);
and U2966 (N_2966,N_2833,N_2809);
nand U2967 (N_2967,N_2823,N_2889);
nand U2968 (N_2968,N_2817,N_2866);
nor U2969 (N_2969,N_2881,N_2891);
nand U2970 (N_2970,N_2806,N_2880);
or U2971 (N_2971,N_2845,N_2897);
nand U2972 (N_2972,N_2868,N_2888);
xor U2973 (N_2973,N_2800,N_2865);
or U2974 (N_2974,N_2892,N_2804);
xor U2975 (N_2975,N_2838,N_2856);
or U2976 (N_2976,N_2856,N_2886);
nor U2977 (N_2977,N_2878,N_2885);
nor U2978 (N_2978,N_2853,N_2850);
nand U2979 (N_2979,N_2840,N_2881);
and U2980 (N_2980,N_2804,N_2851);
nand U2981 (N_2981,N_2870,N_2809);
and U2982 (N_2982,N_2898,N_2846);
xor U2983 (N_2983,N_2874,N_2899);
nor U2984 (N_2984,N_2855,N_2856);
nor U2985 (N_2985,N_2881,N_2856);
or U2986 (N_2986,N_2827,N_2812);
nand U2987 (N_2987,N_2883,N_2846);
xnor U2988 (N_2988,N_2855,N_2822);
or U2989 (N_2989,N_2841,N_2884);
nand U2990 (N_2990,N_2893,N_2850);
or U2991 (N_2991,N_2894,N_2846);
nand U2992 (N_2992,N_2838,N_2894);
or U2993 (N_2993,N_2841,N_2843);
nand U2994 (N_2994,N_2805,N_2848);
and U2995 (N_2995,N_2845,N_2863);
and U2996 (N_2996,N_2866,N_2865);
nor U2997 (N_2997,N_2865,N_2824);
xor U2998 (N_2998,N_2826,N_2845);
and U2999 (N_2999,N_2899,N_2875);
nand U3000 (N_3000,N_2987,N_2930);
nand U3001 (N_3001,N_2956,N_2968);
or U3002 (N_3002,N_2967,N_2963);
xnor U3003 (N_3003,N_2938,N_2998);
and U3004 (N_3004,N_2985,N_2961);
and U3005 (N_3005,N_2900,N_2953);
or U3006 (N_3006,N_2941,N_2936);
and U3007 (N_3007,N_2969,N_2984);
nand U3008 (N_3008,N_2957,N_2971);
nand U3009 (N_3009,N_2997,N_2929);
and U3010 (N_3010,N_2964,N_2990);
nand U3011 (N_3011,N_2973,N_2918);
xor U3012 (N_3012,N_2912,N_2996);
or U3013 (N_3013,N_2906,N_2960);
nor U3014 (N_3014,N_2911,N_2928);
nand U3015 (N_3015,N_2945,N_2901);
nor U3016 (N_3016,N_2940,N_2903);
xor U3017 (N_3017,N_2991,N_2917);
nand U3018 (N_3018,N_2981,N_2946);
nand U3019 (N_3019,N_2979,N_2944);
or U3020 (N_3020,N_2986,N_2924);
xnor U3021 (N_3021,N_2908,N_2980);
or U3022 (N_3022,N_2992,N_2916);
xor U3023 (N_3023,N_2943,N_2937);
xor U3024 (N_3024,N_2915,N_2927);
xnor U3025 (N_3025,N_2999,N_2910);
xnor U3026 (N_3026,N_2965,N_2934);
and U3027 (N_3027,N_2959,N_2921);
or U3028 (N_3028,N_2962,N_2922);
or U3029 (N_3029,N_2907,N_2978);
xor U3030 (N_3030,N_2951,N_2977);
nand U3031 (N_3031,N_2925,N_2972);
or U3032 (N_3032,N_2988,N_2948);
nand U3033 (N_3033,N_2909,N_2942);
or U3034 (N_3034,N_2958,N_2982);
or U3035 (N_3035,N_2970,N_2905);
xnor U3036 (N_3036,N_2975,N_2920);
xor U3037 (N_3037,N_2923,N_2935);
xor U3038 (N_3038,N_2950,N_2932);
and U3039 (N_3039,N_2931,N_2983);
and U3040 (N_3040,N_2995,N_2949);
nor U3041 (N_3041,N_2966,N_2994);
nor U3042 (N_3042,N_2989,N_2954);
and U3043 (N_3043,N_2914,N_2993);
or U3044 (N_3044,N_2976,N_2974);
nor U3045 (N_3045,N_2952,N_2919);
and U3046 (N_3046,N_2913,N_2902);
xor U3047 (N_3047,N_2947,N_2939);
or U3048 (N_3048,N_2904,N_2933);
xnor U3049 (N_3049,N_2955,N_2926);
nand U3050 (N_3050,N_2918,N_2982);
and U3051 (N_3051,N_2999,N_2948);
nand U3052 (N_3052,N_2924,N_2963);
nand U3053 (N_3053,N_2987,N_2958);
nand U3054 (N_3054,N_2985,N_2962);
or U3055 (N_3055,N_2912,N_2976);
or U3056 (N_3056,N_2921,N_2914);
nor U3057 (N_3057,N_2976,N_2938);
nor U3058 (N_3058,N_2965,N_2984);
and U3059 (N_3059,N_2944,N_2958);
nand U3060 (N_3060,N_2997,N_2982);
nor U3061 (N_3061,N_2950,N_2965);
and U3062 (N_3062,N_2911,N_2912);
nand U3063 (N_3063,N_2975,N_2924);
or U3064 (N_3064,N_2932,N_2923);
xor U3065 (N_3065,N_2952,N_2950);
nand U3066 (N_3066,N_2902,N_2936);
nor U3067 (N_3067,N_2986,N_2958);
nand U3068 (N_3068,N_2989,N_2928);
xnor U3069 (N_3069,N_2952,N_2968);
or U3070 (N_3070,N_2964,N_2988);
xor U3071 (N_3071,N_2923,N_2992);
or U3072 (N_3072,N_2936,N_2954);
xnor U3073 (N_3073,N_2941,N_2984);
xnor U3074 (N_3074,N_2932,N_2920);
nor U3075 (N_3075,N_2908,N_2973);
or U3076 (N_3076,N_2989,N_2999);
nand U3077 (N_3077,N_2947,N_2924);
xor U3078 (N_3078,N_2999,N_2951);
nor U3079 (N_3079,N_2950,N_2911);
or U3080 (N_3080,N_2981,N_2968);
and U3081 (N_3081,N_2988,N_2943);
or U3082 (N_3082,N_2902,N_2995);
and U3083 (N_3083,N_2989,N_2988);
nand U3084 (N_3084,N_2976,N_2994);
xor U3085 (N_3085,N_2978,N_2922);
or U3086 (N_3086,N_2971,N_2960);
and U3087 (N_3087,N_2938,N_2909);
xnor U3088 (N_3088,N_2953,N_2932);
xor U3089 (N_3089,N_2986,N_2969);
xor U3090 (N_3090,N_2924,N_2973);
xnor U3091 (N_3091,N_2949,N_2975);
xnor U3092 (N_3092,N_2975,N_2910);
and U3093 (N_3093,N_2999,N_2976);
and U3094 (N_3094,N_2937,N_2976);
or U3095 (N_3095,N_2911,N_2961);
xor U3096 (N_3096,N_2961,N_2952);
xnor U3097 (N_3097,N_2972,N_2986);
xor U3098 (N_3098,N_2977,N_2927);
or U3099 (N_3099,N_2965,N_2982);
or U3100 (N_3100,N_3076,N_3017);
nor U3101 (N_3101,N_3066,N_3003);
nand U3102 (N_3102,N_3010,N_3071);
or U3103 (N_3103,N_3070,N_3068);
or U3104 (N_3104,N_3075,N_3019);
nor U3105 (N_3105,N_3047,N_3034);
or U3106 (N_3106,N_3038,N_3004);
or U3107 (N_3107,N_3063,N_3018);
and U3108 (N_3108,N_3037,N_3043);
xor U3109 (N_3109,N_3036,N_3007);
or U3110 (N_3110,N_3058,N_3069);
xor U3111 (N_3111,N_3077,N_3082);
nand U3112 (N_3112,N_3040,N_3064);
xor U3113 (N_3113,N_3095,N_3094);
xor U3114 (N_3114,N_3041,N_3097);
xor U3115 (N_3115,N_3005,N_3009);
xor U3116 (N_3116,N_3090,N_3000);
and U3117 (N_3117,N_3025,N_3021);
xor U3118 (N_3118,N_3093,N_3065);
and U3119 (N_3119,N_3096,N_3083);
or U3120 (N_3120,N_3061,N_3074);
nor U3121 (N_3121,N_3054,N_3046);
nand U3122 (N_3122,N_3024,N_3023);
or U3123 (N_3123,N_3032,N_3039);
or U3124 (N_3124,N_3013,N_3031);
nor U3125 (N_3125,N_3044,N_3050);
and U3126 (N_3126,N_3042,N_3086);
or U3127 (N_3127,N_3098,N_3091);
or U3128 (N_3128,N_3027,N_3099);
nand U3129 (N_3129,N_3002,N_3067);
nand U3130 (N_3130,N_3006,N_3045);
and U3131 (N_3131,N_3030,N_3011);
and U3132 (N_3132,N_3051,N_3016);
nand U3133 (N_3133,N_3029,N_3056);
xnor U3134 (N_3134,N_3012,N_3080);
nor U3135 (N_3135,N_3035,N_3092);
nand U3136 (N_3136,N_3022,N_3028);
xnor U3137 (N_3137,N_3085,N_3088);
and U3138 (N_3138,N_3060,N_3057);
xnor U3139 (N_3139,N_3062,N_3081);
xnor U3140 (N_3140,N_3089,N_3020);
and U3141 (N_3141,N_3015,N_3049);
xnor U3142 (N_3142,N_3008,N_3052);
nor U3143 (N_3143,N_3084,N_3059);
nand U3144 (N_3144,N_3079,N_3026);
and U3145 (N_3145,N_3048,N_3072);
and U3146 (N_3146,N_3073,N_3033);
nor U3147 (N_3147,N_3055,N_3001);
nand U3148 (N_3148,N_3078,N_3053);
and U3149 (N_3149,N_3014,N_3087);
xor U3150 (N_3150,N_3049,N_3097);
nand U3151 (N_3151,N_3047,N_3090);
xor U3152 (N_3152,N_3076,N_3023);
nor U3153 (N_3153,N_3019,N_3095);
xnor U3154 (N_3154,N_3038,N_3079);
nand U3155 (N_3155,N_3005,N_3002);
and U3156 (N_3156,N_3047,N_3051);
or U3157 (N_3157,N_3068,N_3007);
nand U3158 (N_3158,N_3068,N_3095);
xnor U3159 (N_3159,N_3071,N_3036);
xnor U3160 (N_3160,N_3055,N_3062);
or U3161 (N_3161,N_3084,N_3055);
nor U3162 (N_3162,N_3019,N_3064);
nand U3163 (N_3163,N_3097,N_3020);
and U3164 (N_3164,N_3069,N_3074);
nand U3165 (N_3165,N_3054,N_3008);
nand U3166 (N_3166,N_3014,N_3063);
or U3167 (N_3167,N_3058,N_3032);
xor U3168 (N_3168,N_3045,N_3008);
xor U3169 (N_3169,N_3032,N_3052);
xor U3170 (N_3170,N_3096,N_3017);
and U3171 (N_3171,N_3062,N_3076);
and U3172 (N_3172,N_3021,N_3064);
nor U3173 (N_3173,N_3014,N_3005);
or U3174 (N_3174,N_3094,N_3027);
nand U3175 (N_3175,N_3078,N_3038);
xor U3176 (N_3176,N_3002,N_3012);
xnor U3177 (N_3177,N_3006,N_3069);
nor U3178 (N_3178,N_3084,N_3002);
and U3179 (N_3179,N_3037,N_3092);
nand U3180 (N_3180,N_3061,N_3028);
and U3181 (N_3181,N_3083,N_3019);
xor U3182 (N_3182,N_3094,N_3092);
nand U3183 (N_3183,N_3034,N_3031);
and U3184 (N_3184,N_3079,N_3016);
or U3185 (N_3185,N_3048,N_3089);
nand U3186 (N_3186,N_3013,N_3075);
xor U3187 (N_3187,N_3085,N_3001);
xor U3188 (N_3188,N_3070,N_3078);
nor U3189 (N_3189,N_3001,N_3024);
nand U3190 (N_3190,N_3063,N_3006);
and U3191 (N_3191,N_3008,N_3048);
and U3192 (N_3192,N_3066,N_3090);
and U3193 (N_3193,N_3007,N_3003);
nand U3194 (N_3194,N_3030,N_3050);
nor U3195 (N_3195,N_3054,N_3041);
nand U3196 (N_3196,N_3021,N_3059);
nor U3197 (N_3197,N_3070,N_3081);
xor U3198 (N_3198,N_3075,N_3089);
or U3199 (N_3199,N_3066,N_3085);
nand U3200 (N_3200,N_3125,N_3184);
nand U3201 (N_3201,N_3161,N_3189);
and U3202 (N_3202,N_3170,N_3152);
or U3203 (N_3203,N_3148,N_3142);
nor U3204 (N_3204,N_3160,N_3182);
xor U3205 (N_3205,N_3144,N_3130);
nor U3206 (N_3206,N_3107,N_3164);
and U3207 (N_3207,N_3122,N_3169);
nor U3208 (N_3208,N_3187,N_3186);
nand U3209 (N_3209,N_3135,N_3132);
xor U3210 (N_3210,N_3139,N_3115);
xnor U3211 (N_3211,N_3171,N_3176);
or U3212 (N_3212,N_3194,N_3150);
xor U3213 (N_3213,N_3157,N_3198);
or U3214 (N_3214,N_3102,N_3149);
xnor U3215 (N_3215,N_3101,N_3117);
or U3216 (N_3216,N_3128,N_3188);
nor U3217 (N_3217,N_3116,N_3195);
nand U3218 (N_3218,N_3145,N_3147);
and U3219 (N_3219,N_3168,N_3167);
and U3220 (N_3220,N_3162,N_3105);
and U3221 (N_3221,N_3190,N_3154);
or U3222 (N_3222,N_3114,N_3192);
and U3223 (N_3223,N_3134,N_3112);
xor U3224 (N_3224,N_3146,N_3177);
or U3225 (N_3225,N_3118,N_3183);
and U3226 (N_3226,N_3156,N_3126);
and U3227 (N_3227,N_3165,N_3119);
nor U3228 (N_3228,N_3138,N_3159);
xnor U3229 (N_3229,N_3104,N_3131);
and U3230 (N_3230,N_3185,N_3191);
and U3231 (N_3231,N_3129,N_3140);
xnor U3232 (N_3232,N_3166,N_3109);
nor U3233 (N_3233,N_3133,N_3172);
xnor U3234 (N_3234,N_3197,N_3141);
xnor U3235 (N_3235,N_3111,N_3120);
xnor U3236 (N_3236,N_3143,N_3199);
or U3237 (N_3237,N_3137,N_3174);
and U3238 (N_3238,N_3173,N_3155);
and U3239 (N_3239,N_3100,N_3178);
or U3240 (N_3240,N_3103,N_3136);
nor U3241 (N_3241,N_3106,N_3175);
or U3242 (N_3242,N_3124,N_3127);
nand U3243 (N_3243,N_3196,N_3123);
xor U3244 (N_3244,N_3151,N_3193);
nand U3245 (N_3245,N_3153,N_3108);
nor U3246 (N_3246,N_3181,N_3110);
nor U3247 (N_3247,N_3180,N_3121);
nand U3248 (N_3248,N_3179,N_3163);
or U3249 (N_3249,N_3113,N_3158);
xor U3250 (N_3250,N_3188,N_3197);
xnor U3251 (N_3251,N_3169,N_3120);
and U3252 (N_3252,N_3118,N_3180);
and U3253 (N_3253,N_3191,N_3189);
or U3254 (N_3254,N_3103,N_3107);
or U3255 (N_3255,N_3131,N_3122);
nand U3256 (N_3256,N_3158,N_3195);
nand U3257 (N_3257,N_3197,N_3103);
or U3258 (N_3258,N_3153,N_3109);
or U3259 (N_3259,N_3151,N_3185);
xnor U3260 (N_3260,N_3188,N_3137);
or U3261 (N_3261,N_3139,N_3103);
xor U3262 (N_3262,N_3153,N_3148);
or U3263 (N_3263,N_3199,N_3181);
xor U3264 (N_3264,N_3107,N_3124);
or U3265 (N_3265,N_3183,N_3113);
xor U3266 (N_3266,N_3135,N_3182);
nand U3267 (N_3267,N_3125,N_3131);
or U3268 (N_3268,N_3122,N_3111);
or U3269 (N_3269,N_3182,N_3161);
xor U3270 (N_3270,N_3175,N_3196);
or U3271 (N_3271,N_3189,N_3159);
or U3272 (N_3272,N_3139,N_3163);
nor U3273 (N_3273,N_3126,N_3150);
or U3274 (N_3274,N_3148,N_3140);
xnor U3275 (N_3275,N_3145,N_3100);
nor U3276 (N_3276,N_3141,N_3163);
or U3277 (N_3277,N_3117,N_3109);
or U3278 (N_3278,N_3135,N_3129);
nand U3279 (N_3279,N_3111,N_3121);
and U3280 (N_3280,N_3135,N_3139);
and U3281 (N_3281,N_3147,N_3159);
or U3282 (N_3282,N_3118,N_3163);
and U3283 (N_3283,N_3151,N_3167);
nand U3284 (N_3284,N_3105,N_3148);
nor U3285 (N_3285,N_3102,N_3169);
and U3286 (N_3286,N_3191,N_3119);
nand U3287 (N_3287,N_3175,N_3179);
or U3288 (N_3288,N_3154,N_3168);
nand U3289 (N_3289,N_3116,N_3149);
or U3290 (N_3290,N_3130,N_3102);
xor U3291 (N_3291,N_3115,N_3155);
nor U3292 (N_3292,N_3145,N_3105);
xor U3293 (N_3293,N_3113,N_3114);
nand U3294 (N_3294,N_3164,N_3181);
or U3295 (N_3295,N_3163,N_3145);
and U3296 (N_3296,N_3186,N_3148);
xnor U3297 (N_3297,N_3142,N_3128);
xor U3298 (N_3298,N_3113,N_3130);
xor U3299 (N_3299,N_3124,N_3159);
xnor U3300 (N_3300,N_3239,N_3248);
or U3301 (N_3301,N_3231,N_3234);
nand U3302 (N_3302,N_3237,N_3219);
xor U3303 (N_3303,N_3226,N_3252);
nor U3304 (N_3304,N_3260,N_3285);
nor U3305 (N_3305,N_3222,N_3200);
xnor U3306 (N_3306,N_3203,N_3242);
nor U3307 (N_3307,N_3251,N_3295);
xnor U3308 (N_3308,N_3270,N_3213);
or U3309 (N_3309,N_3292,N_3299);
nand U3310 (N_3310,N_3223,N_3291);
and U3311 (N_3311,N_3293,N_3281);
or U3312 (N_3312,N_3256,N_3258);
xor U3313 (N_3313,N_3298,N_3230);
or U3314 (N_3314,N_3272,N_3246);
or U3315 (N_3315,N_3263,N_3288);
nand U3316 (N_3316,N_3275,N_3279);
nand U3317 (N_3317,N_3243,N_3216);
nor U3318 (N_3318,N_3294,N_3262);
xor U3319 (N_3319,N_3276,N_3241);
nand U3320 (N_3320,N_3296,N_3290);
or U3321 (N_3321,N_3254,N_3210);
nor U3322 (N_3322,N_3225,N_3249);
nor U3323 (N_3323,N_3267,N_3218);
nand U3324 (N_3324,N_3232,N_3229);
nor U3325 (N_3325,N_3240,N_3221);
and U3326 (N_3326,N_3269,N_3250);
nand U3327 (N_3327,N_3233,N_3202);
xnor U3328 (N_3328,N_3205,N_3289);
or U3329 (N_3329,N_3215,N_3208);
nand U3330 (N_3330,N_3255,N_3257);
nor U3331 (N_3331,N_3261,N_3212);
or U3332 (N_3332,N_3206,N_3274);
nand U3333 (N_3333,N_3204,N_3238);
nor U3334 (N_3334,N_3282,N_3297);
nand U3335 (N_3335,N_3277,N_3278);
nor U3336 (N_3336,N_3228,N_3214);
nor U3337 (N_3337,N_3280,N_3284);
xor U3338 (N_3338,N_3253,N_3271);
and U3339 (N_3339,N_3265,N_3211);
and U3340 (N_3340,N_3244,N_3236);
xnor U3341 (N_3341,N_3209,N_3273);
xor U3342 (N_3342,N_3245,N_3220);
xor U3343 (N_3343,N_3268,N_3235);
nand U3344 (N_3344,N_3283,N_3224);
xor U3345 (N_3345,N_3287,N_3201);
nor U3346 (N_3346,N_3247,N_3259);
xor U3347 (N_3347,N_3286,N_3266);
or U3348 (N_3348,N_3227,N_3217);
or U3349 (N_3349,N_3264,N_3207);
or U3350 (N_3350,N_3241,N_3219);
nand U3351 (N_3351,N_3250,N_3219);
or U3352 (N_3352,N_3200,N_3219);
nand U3353 (N_3353,N_3286,N_3227);
xnor U3354 (N_3354,N_3265,N_3231);
xnor U3355 (N_3355,N_3241,N_3296);
xor U3356 (N_3356,N_3283,N_3252);
nand U3357 (N_3357,N_3230,N_3280);
or U3358 (N_3358,N_3270,N_3207);
nor U3359 (N_3359,N_3284,N_3210);
nand U3360 (N_3360,N_3214,N_3290);
nand U3361 (N_3361,N_3200,N_3273);
or U3362 (N_3362,N_3289,N_3285);
or U3363 (N_3363,N_3258,N_3253);
nand U3364 (N_3364,N_3250,N_3294);
nand U3365 (N_3365,N_3284,N_3216);
or U3366 (N_3366,N_3209,N_3277);
nand U3367 (N_3367,N_3219,N_3295);
xnor U3368 (N_3368,N_3248,N_3270);
and U3369 (N_3369,N_3239,N_3219);
and U3370 (N_3370,N_3273,N_3247);
nand U3371 (N_3371,N_3275,N_3236);
nor U3372 (N_3372,N_3242,N_3202);
nand U3373 (N_3373,N_3205,N_3255);
or U3374 (N_3374,N_3296,N_3295);
or U3375 (N_3375,N_3240,N_3288);
xor U3376 (N_3376,N_3201,N_3241);
nand U3377 (N_3377,N_3255,N_3286);
and U3378 (N_3378,N_3238,N_3292);
xor U3379 (N_3379,N_3299,N_3211);
nand U3380 (N_3380,N_3294,N_3242);
or U3381 (N_3381,N_3200,N_3275);
nand U3382 (N_3382,N_3266,N_3297);
nor U3383 (N_3383,N_3287,N_3284);
or U3384 (N_3384,N_3224,N_3230);
and U3385 (N_3385,N_3273,N_3252);
or U3386 (N_3386,N_3241,N_3220);
nand U3387 (N_3387,N_3256,N_3273);
xnor U3388 (N_3388,N_3293,N_3278);
and U3389 (N_3389,N_3258,N_3278);
or U3390 (N_3390,N_3271,N_3257);
and U3391 (N_3391,N_3271,N_3284);
nor U3392 (N_3392,N_3269,N_3224);
or U3393 (N_3393,N_3243,N_3208);
nor U3394 (N_3394,N_3212,N_3294);
nor U3395 (N_3395,N_3260,N_3211);
nand U3396 (N_3396,N_3201,N_3223);
nand U3397 (N_3397,N_3262,N_3277);
xor U3398 (N_3398,N_3280,N_3246);
or U3399 (N_3399,N_3289,N_3235);
and U3400 (N_3400,N_3385,N_3388);
xnor U3401 (N_3401,N_3358,N_3334);
nand U3402 (N_3402,N_3389,N_3386);
or U3403 (N_3403,N_3398,N_3333);
nor U3404 (N_3404,N_3352,N_3374);
nor U3405 (N_3405,N_3345,N_3335);
nand U3406 (N_3406,N_3338,N_3399);
xor U3407 (N_3407,N_3365,N_3331);
or U3408 (N_3408,N_3311,N_3381);
and U3409 (N_3409,N_3305,N_3394);
xor U3410 (N_3410,N_3319,N_3326);
nand U3411 (N_3411,N_3350,N_3306);
xnor U3412 (N_3412,N_3375,N_3327);
nor U3413 (N_3413,N_3322,N_3384);
nor U3414 (N_3414,N_3393,N_3336);
nand U3415 (N_3415,N_3392,N_3321);
nand U3416 (N_3416,N_3387,N_3301);
nor U3417 (N_3417,N_3360,N_3348);
nand U3418 (N_3418,N_3342,N_3320);
nand U3419 (N_3419,N_3373,N_3390);
nor U3420 (N_3420,N_3341,N_3304);
nand U3421 (N_3421,N_3377,N_3300);
xnor U3422 (N_3422,N_3353,N_3396);
and U3423 (N_3423,N_3339,N_3329);
or U3424 (N_3424,N_3378,N_3303);
nand U3425 (N_3425,N_3328,N_3309);
and U3426 (N_3426,N_3356,N_3343);
nor U3427 (N_3427,N_3351,N_3325);
nor U3428 (N_3428,N_3330,N_3364);
xnor U3429 (N_3429,N_3317,N_3370);
nor U3430 (N_3430,N_3395,N_3382);
or U3431 (N_3431,N_3313,N_3316);
or U3432 (N_3432,N_3368,N_3362);
xor U3433 (N_3433,N_3372,N_3366);
and U3434 (N_3434,N_3332,N_3347);
nor U3435 (N_3435,N_3361,N_3310);
and U3436 (N_3436,N_3312,N_3355);
nand U3437 (N_3437,N_3359,N_3323);
or U3438 (N_3438,N_3363,N_3369);
nor U3439 (N_3439,N_3367,N_3391);
and U3440 (N_3440,N_3376,N_3380);
or U3441 (N_3441,N_3340,N_3318);
nor U3442 (N_3442,N_3307,N_3383);
xnor U3443 (N_3443,N_3337,N_3314);
nand U3444 (N_3444,N_3354,N_3379);
xor U3445 (N_3445,N_3357,N_3324);
nand U3446 (N_3446,N_3397,N_3346);
and U3447 (N_3447,N_3344,N_3302);
nand U3448 (N_3448,N_3371,N_3315);
nor U3449 (N_3449,N_3349,N_3308);
xor U3450 (N_3450,N_3345,N_3374);
xor U3451 (N_3451,N_3374,N_3386);
or U3452 (N_3452,N_3361,N_3354);
xnor U3453 (N_3453,N_3382,N_3363);
nand U3454 (N_3454,N_3323,N_3390);
or U3455 (N_3455,N_3340,N_3333);
and U3456 (N_3456,N_3349,N_3372);
xor U3457 (N_3457,N_3346,N_3369);
and U3458 (N_3458,N_3375,N_3386);
xnor U3459 (N_3459,N_3382,N_3347);
xnor U3460 (N_3460,N_3320,N_3388);
nor U3461 (N_3461,N_3305,N_3351);
nand U3462 (N_3462,N_3323,N_3366);
nand U3463 (N_3463,N_3354,N_3373);
and U3464 (N_3464,N_3375,N_3380);
or U3465 (N_3465,N_3312,N_3352);
or U3466 (N_3466,N_3316,N_3323);
or U3467 (N_3467,N_3322,N_3326);
or U3468 (N_3468,N_3370,N_3325);
or U3469 (N_3469,N_3314,N_3396);
or U3470 (N_3470,N_3379,N_3375);
nand U3471 (N_3471,N_3327,N_3395);
and U3472 (N_3472,N_3314,N_3307);
nand U3473 (N_3473,N_3366,N_3338);
nand U3474 (N_3474,N_3308,N_3373);
and U3475 (N_3475,N_3342,N_3393);
xnor U3476 (N_3476,N_3364,N_3344);
xnor U3477 (N_3477,N_3306,N_3363);
nand U3478 (N_3478,N_3380,N_3301);
and U3479 (N_3479,N_3367,N_3329);
and U3480 (N_3480,N_3333,N_3392);
nand U3481 (N_3481,N_3345,N_3382);
or U3482 (N_3482,N_3385,N_3360);
xor U3483 (N_3483,N_3333,N_3384);
nor U3484 (N_3484,N_3362,N_3392);
xnor U3485 (N_3485,N_3384,N_3393);
nand U3486 (N_3486,N_3325,N_3377);
nor U3487 (N_3487,N_3394,N_3390);
or U3488 (N_3488,N_3331,N_3375);
xor U3489 (N_3489,N_3344,N_3337);
and U3490 (N_3490,N_3342,N_3318);
nand U3491 (N_3491,N_3312,N_3328);
and U3492 (N_3492,N_3386,N_3381);
nor U3493 (N_3493,N_3399,N_3363);
and U3494 (N_3494,N_3393,N_3396);
xnor U3495 (N_3495,N_3309,N_3319);
or U3496 (N_3496,N_3354,N_3369);
xor U3497 (N_3497,N_3357,N_3306);
and U3498 (N_3498,N_3321,N_3316);
nand U3499 (N_3499,N_3392,N_3332);
nor U3500 (N_3500,N_3460,N_3409);
or U3501 (N_3501,N_3459,N_3412);
or U3502 (N_3502,N_3447,N_3470);
xor U3503 (N_3503,N_3457,N_3466);
nor U3504 (N_3504,N_3429,N_3446);
and U3505 (N_3505,N_3404,N_3431);
or U3506 (N_3506,N_3481,N_3467);
xor U3507 (N_3507,N_3433,N_3454);
and U3508 (N_3508,N_3406,N_3495);
xor U3509 (N_3509,N_3441,N_3477);
nand U3510 (N_3510,N_3487,N_3438);
nor U3511 (N_3511,N_3469,N_3453);
xor U3512 (N_3512,N_3475,N_3462);
nor U3513 (N_3513,N_3449,N_3483);
xor U3514 (N_3514,N_3430,N_3484);
and U3515 (N_3515,N_3499,N_3417);
nand U3516 (N_3516,N_3480,N_3408);
xor U3517 (N_3517,N_3405,N_3497);
or U3518 (N_3518,N_3472,N_3420);
nor U3519 (N_3519,N_3456,N_3452);
and U3520 (N_3520,N_3491,N_3415);
nand U3521 (N_3521,N_3434,N_3473);
xor U3522 (N_3522,N_3437,N_3465);
nand U3523 (N_3523,N_3440,N_3458);
xor U3524 (N_3524,N_3471,N_3479);
or U3525 (N_3525,N_3427,N_3402);
and U3526 (N_3526,N_3476,N_3451);
nor U3527 (N_3527,N_3489,N_3486);
and U3528 (N_3528,N_3442,N_3403);
xor U3529 (N_3529,N_3474,N_3401);
and U3530 (N_3530,N_3439,N_3468);
and U3531 (N_3531,N_3422,N_3461);
nor U3532 (N_3532,N_3419,N_3496);
xor U3533 (N_3533,N_3410,N_3463);
and U3534 (N_3534,N_3418,N_3478);
nor U3535 (N_3535,N_3492,N_3455);
or U3536 (N_3536,N_3423,N_3413);
nand U3537 (N_3537,N_3407,N_3421);
or U3538 (N_3538,N_3443,N_3416);
nor U3539 (N_3539,N_3424,N_3411);
nor U3540 (N_3540,N_3485,N_3400);
nand U3541 (N_3541,N_3490,N_3436);
nand U3542 (N_3542,N_3432,N_3448);
or U3543 (N_3543,N_3494,N_3444);
xnor U3544 (N_3544,N_3425,N_3450);
xnor U3545 (N_3545,N_3464,N_3435);
xor U3546 (N_3546,N_3445,N_3493);
xnor U3547 (N_3547,N_3414,N_3426);
and U3548 (N_3548,N_3498,N_3488);
or U3549 (N_3549,N_3428,N_3482);
or U3550 (N_3550,N_3401,N_3482);
nand U3551 (N_3551,N_3425,N_3404);
xnor U3552 (N_3552,N_3432,N_3480);
and U3553 (N_3553,N_3458,N_3417);
or U3554 (N_3554,N_3473,N_3437);
or U3555 (N_3555,N_3443,N_3456);
xor U3556 (N_3556,N_3428,N_3460);
xnor U3557 (N_3557,N_3471,N_3447);
nor U3558 (N_3558,N_3466,N_3416);
and U3559 (N_3559,N_3418,N_3414);
nor U3560 (N_3560,N_3432,N_3411);
nor U3561 (N_3561,N_3488,N_3470);
or U3562 (N_3562,N_3424,N_3486);
or U3563 (N_3563,N_3417,N_3416);
xor U3564 (N_3564,N_3419,N_3426);
xnor U3565 (N_3565,N_3408,N_3430);
xnor U3566 (N_3566,N_3467,N_3498);
and U3567 (N_3567,N_3433,N_3403);
xnor U3568 (N_3568,N_3426,N_3425);
xnor U3569 (N_3569,N_3473,N_3423);
nand U3570 (N_3570,N_3405,N_3464);
or U3571 (N_3571,N_3441,N_3491);
nand U3572 (N_3572,N_3449,N_3496);
nor U3573 (N_3573,N_3415,N_3482);
and U3574 (N_3574,N_3463,N_3455);
nor U3575 (N_3575,N_3467,N_3440);
and U3576 (N_3576,N_3415,N_3424);
or U3577 (N_3577,N_3453,N_3433);
or U3578 (N_3578,N_3435,N_3457);
or U3579 (N_3579,N_3428,N_3401);
xnor U3580 (N_3580,N_3451,N_3430);
nand U3581 (N_3581,N_3497,N_3459);
nor U3582 (N_3582,N_3443,N_3457);
nor U3583 (N_3583,N_3452,N_3462);
nor U3584 (N_3584,N_3462,N_3490);
xnor U3585 (N_3585,N_3492,N_3447);
nor U3586 (N_3586,N_3463,N_3464);
nand U3587 (N_3587,N_3479,N_3468);
or U3588 (N_3588,N_3445,N_3427);
or U3589 (N_3589,N_3481,N_3495);
and U3590 (N_3590,N_3452,N_3482);
or U3591 (N_3591,N_3451,N_3470);
and U3592 (N_3592,N_3483,N_3460);
and U3593 (N_3593,N_3450,N_3415);
or U3594 (N_3594,N_3446,N_3480);
xor U3595 (N_3595,N_3484,N_3485);
and U3596 (N_3596,N_3450,N_3408);
and U3597 (N_3597,N_3487,N_3448);
xor U3598 (N_3598,N_3486,N_3464);
xor U3599 (N_3599,N_3414,N_3489);
or U3600 (N_3600,N_3570,N_3546);
xor U3601 (N_3601,N_3502,N_3573);
and U3602 (N_3602,N_3555,N_3562);
xnor U3603 (N_3603,N_3557,N_3592);
nand U3604 (N_3604,N_3520,N_3582);
and U3605 (N_3605,N_3561,N_3579);
or U3606 (N_3606,N_3585,N_3524);
and U3607 (N_3607,N_3556,N_3537);
nand U3608 (N_3608,N_3558,N_3541);
and U3609 (N_3609,N_3594,N_3506);
and U3610 (N_3610,N_3547,N_3580);
xor U3611 (N_3611,N_3574,N_3563);
xnor U3612 (N_3612,N_3587,N_3503);
nor U3613 (N_3613,N_3581,N_3545);
and U3614 (N_3614,N_3518,N_3598);
nand U3615 (N_3615,N_3593,N_3571);
nand U3616 (N_3616,N_3522,N_3559);
nor U3617 (N_3617,N_3554,N_3508);
nand U3618 (N_3618,N_3523,N_3517);
xnor U3619 (N_3619,N_3532,N_3536);
xnor U3620 (N_3620,N_3516,N_3577);
or U3621 (N_3621,N_3501,N_3514);
or U3622 (N_3622,N_3560,N_3567);
and U3623 (N_3623,N_3507,N_3564);
or U3624 (N_3624,N_3565,N_3540);
and U3625 (N_3625,N_3529,N_3599);
nor U3626 (N_3626,N_3586,N_3500);
and U3627 (N_3627,N_3569,N_3504);
nand U3628 (N_3628,N_3597,N_3591);
xnor U3629 (N_3629,N_3530,N_3596);
nand U3630 (N_3630,N_3544,N_3505);
or U3631 (N_3631,N_3512,N_3589);
and U3632 (N_3632,N_3509,N_3566);
or U3633 (N_3633,N_3552,N_3576);
nor U3634 (N_3634,N_3553,N_3551);
nor U3635 (N_3635,N_3568,N_3542);
nor U3636 (N_3636,N_3548,N_3526);
nor U3637 (N_3637,N_3525,N_3535);
or U3638 (N_3638,N_3550,N_3527);
xnor U3639 (N_3639,N_3521,N_3584);
nor U3640 (N_3640,N_3588,N_3513);
nor U3641 (N_3641,N_3519,N_3511);
nor U3642 (N_3642,N_3590,N_3549);
nor U3643 (N_3643,N_3534,N_3538);
xor U3644 (N_3644,N_3539,N_3510);
and U3645 (N_3645,N_3583,N_3572);
nor U3646 (N_3646,N_3575,N_3528);
xnor U3647 (N_3647,N_3543,N_3578);
xnor U3648 (N_3648,N_3531,N_3515);
xor U3649 (N_3649,N_3595,N_3533);
nor U3650 (N_3650,N_3599,N_3558);
nor U3651 (N_3651,N_3575,N_3508);
or U3652 (N_3652,N_3580,N_3566);
nor U3653 (N_3653,N_3540,N_3502);
nor U3654 (N_3654,N_3504,N_3586);
nand U3655 (N_3655,N_3550,N_3588);
nand U3656 (N_3656,N_3584,N_3546);
and U3657 (N_3657,N_3512,N_3525);
nand U3658 (N_3658,N_3564,N_3514);
nor U3659 (N_3659,N_3599,N_3560);
nand U3660 (N_3660,N_3527,N_3546);
nand U3661 (N_3661,N_3504,N_3568);
and U3662 (N_3662,N_3594,N_3547);
or U3663 (N_3663,N_3563,N_3515);
xnor U3664 (N_3664,N_3577,N_3556);
xor U3665 (N_3665,N_3543,N_3566);
or U3666 (N_3666,N_3597,N_3584);
and U3667 (N_3667,N_3552,N_3572);
or U3668 (N_3668,N_3551,N_3580);
or U3669 (N_3669,N_3529,N_3551);
and U3670 (N_3670,N_3517,N_3559);
or U3671 (N_3671,N_3577,N_3558);
nor U3672 (N_3672,N_3556,N_3524);
nor U3673 (N_3673,N_3543,N_3575);
xnor U3674 (N_3674,N_3599,N_3593);
and U3675 (N_3675,N_3537,N_3573);
nand U3676 (N_3676,N_3545,N_3537);
nor U3677 (N_3677,N_3570,N_3530);
nand U3678 (N_3678,N_3520,N_3559);
and U3679 (N_3679,N_3569,N_3508);
xor U3680 (N_3680,N_3541,N_3578);
xnor U3681 (N_3681,N_3574,N_3581);
or U3682 (N_3682,N_3531,N_3570);
nand U3683 (N_3683,N_3537,N_3514);
and U3684 (N_3684,N_3560,N_3571);
and U3685 (N_3685,N_3518,N_3592);
and U3686 (N_3686,N_3503,N_3550);
nor U3687 (N_3687,N_3581,N_3521);
or U3688 (N_3688,N_3572,N_3595);
and U3689 (N_3689,N_3575,N_3566);
or U3690 (N_3690,N_3585,N_3583);
and U3691 (N_3691,N_3533,N_3568);
xor U3692 (N_3692,N_3537,N_3560);
xor U3693 (N_3693,N_3574,N_3569);
xor U3694 (N_3694,N_3558,N_3556);
nor U3695 (N_3695,N_3573,N_3554);
xnor U3696 (N_3696,N_3522,N_3550);
and U3697 (N_3697,N_3524,N_3555);
nand U3698 (N_3698,N_3551,N_3550);
and U3699 (N_3699,N_3576,N_3515);
xnor U3700 (N_3700,N_3634,N_3605);
or U3701 (N_3701,N_3620,N_3696);
xnor U3702 (N_3702,N_3642,N_3655);
nor U3703 (N_3703,N_3691,N_3659);
and U3704 (N_3704,N_3680,N_3638);
and U3705 (N_3705,N_3650,N_3619);
nand U3706 (N_3706,N_3686,N_3673);
or U3707 (N_3707,N_3643,N_3630);
or U3708 (N_3708,N_3617,N_3623);
nor U3709 (N_3709,N_3684,N_3667);
nor U3710 (N_3710,N_3645,N_3669);
xor U3711 (N_3711,N_3687,N_3690);
xnor U3712 (N_3712,N_3639,N_3657);
and U3713 (N_3713,N_3651,N_3612);
nand U3714 (N_3714,N_3616,N_3604);
nand U3715 (N_3715,N_3636,N_3683);
nand U3716 (N_3716,N_3609,N_3661);
xnor U3717 (N_3717,N_3675,N_3664);
and U3718 (N_3718,N_3640,N_3637);
nor U3719 (N_3719,N_3633,N_3693);
nor U3720 (N_3720,N_3628,N_3694);
and U3721 (N_3721,N_3629,N_3649);
or U3722 (N_3722,N_3666,N_3646);
and U3723 (N_3723,N_3656,N_3648);
nand U3724 (N_3724,N_3615,N_3603);
nor U3725 (N_3725,N_3662,N_3607);
nand U3726 (N_3726,N_3695,N_3610);
nand U3727 (N_3727,N_3613,N_3608);
xor U3728 (N_3728,N_3600,N_3674);
nand U3729 (N_3729,N_3676,N_3631);
and U3730 (N_3730,N_3626,N_3625);
xnor U3731 (N_3731,N_3681,N_3624);
or U3732 (N_3732,N_3632,N_3652);
xnor U3733 (N_3733,N_3601,N_3622);
and U3734 (N_3734,N_3665,N_3621);
or U3735 (N_3735,N_3602,N_3682);
nor U3736 (N_3736,N_3671,N_3611);
and U3737 (N_3737,N_3654,N_3698);
xor U3738 (N_3738,N_3697,N_3658);
xnor U3739 (N_3739,N_3668,N_3688);
nor U3740 (N_3740,N_3653,N_3614);
nor U3741 (N_3741,N_3641,N_3660);
xor U3742 (N_3742,N_3699,N_3692);
or U3743 (N_3743,N_3618,N_3663);
nor U3744 (N_3744,N_3606,N_3635);
nand U3745 (N_3745,N_3677,N_3670);
or U3746 (N_3746,N_3644,N_3678);
or U3747 (N_3747,N_3627,N_3672);
nand U3748 (N_3748,N_3647,N_3679);
xnor U3749 (N_3749,N_3685,N_3689);
or U3750 (N_3750,N_3631,N_3697);
or U3751 (N_3751,N_3620,N_3694);
xnor U3752 (N_3752,N_3641,N_3645);
nand U3753 (N_3753,N_3617,N_3657);
and U3754 (N_3754,N_3669,N_3623);
xor U3755 (N_3755,N_3615,N_3692);
nand U3756 (N_3756,N_3621,N_3670);
or U3757 (N_3757,N_3641,N_3642);
and U3758 (N_3758,N_3670,N_3615);
nor U3759 (N_3759,N_3690,N_3658);
xnor U3760 (N_3760,N_3671,N_3665);
or U3761 (N_3761,N_3618,N_3682);
and U3762 (N_3762,N_3678,N_3658);
and U3763 (N_3763,N_3602,N_3621);
nand U3764 (N_3764,N_3643,N_3698);
nand U3765 (N_3765,N_3617,N_3675);
xnor U3766 (N_3766,N_3627,N_3696);
nor U3767 (N_3767,N_3651,N_3699);
and U3768 (N_3768,N_3637,N_3664);
and U3769 (N_3769,N_3638,N_3637);
or U3770 (N_3770,N_3617,N_3669);
nand U3771 (N_3771,N_3608,N_3666);
nand U3772 (N_3772,N_3694,N_3677);
xnor U3773 (N_3773,N_3672,N_3684);
and U3774 (N_3774,N_3617,N_3699);
xor U3775 (N_3775,N_3676,N_3658);
xor U3776 (N_3776,N_3617,N_3687);
or U3777 (N_3777,N_3675,N_3643);
or U3778 (N_3778,N_3631,N_3648);
nand U3779 (N_3779,N_3681,N_3604);
nand U3780 (N_3780,N_3604,N_3641);
xnor U3781 (N_3781,N_3619,N_3661);
nor U3782 (N_3782,N_3600,N_3650);
and U3783 (N_3783,N_3660,N_3611);
and U3784 (N_3784,N_3697,N_3681);
or U3785 (N_3785,N_3661,N_3649);
or U3786 (N_3786,N_3685,N_3677);
nor U3787 (N_3787,N_3693,N_3654);
nor U3788 (N_3788,N_3639,N_3653);
xnor U3789 (N_3789,N_3630,N_3679);
xnor U3790 (N_3790,N_3635,N_3634);
and U3791 (N_3791,N_3685,N_3698);
nand U3792 (N_3792,N_3643,N_3689);
or U3793 (N_3793,N_3677,N_3644);
or U3794 (N_3794,N_3621,N_3674);
or U3795 (N_3795,N_3681,N_3647);
nand U3796 (N_3796,N_3670,N_3694);
and U3797 (N_3797,N_3634,N_3637);
xor U3798 (N_3798,N_3631,N_3655);
nor U3799 (N_3799,N_3694,N_3629);
and U3800 (N_3800,N_3786,N_3704);
or U3801 (N_3801,N_3796,N_3740);
nor U3802 (N_3802,N_3788,N_3729);
xnor U3803 (N_3803,N_3714,N_3752);
nand U3804 (N_3804,N_3747,N_3793);
xnor U3805 (N_3805,N_3741,N_3719);
nor U3806 (N_3806,N_3773,N_3718);
and U3807 (N_3807,N_3790,N_3727);
and U3808 (N_3808,N_3724,N_3759);
nor U3809 (N_3809,N_3709,N_3787);
nor U3810 (N_3810,N_3776,N_3792);
nor U3811 (N_3811,N_3750,N_3725);
nand U3812 (N_3812,N_3763,N_3721);
nand U3813 (N_3813,N_3748,N_3780);
xor U3814 (N_3814,N_3798,N_3743);
nor U3815 (N_3815,N_3702,N_3771);
xor U3816 (N_3816,N_3795,N_3738);
xor U3817 (N_3817,N_3784,N_3713);
xor U3818 (N_3818,N_3770,N_3799);
or U3819 (N_3819,N_3716,N_3711);
or U3820 (N_3820,N_3757,N_3735);
and U3821 (N_3821,N_3737,N_3730);
xnor U3822 (N_3822,N_3785,N_3736);
xor U3823 (N_3823,N_3746,N_3708);
and U3824 (N_3824,N_3783,N_3710);
nor U3825 (N_3825,N_3717,N_3779);
nand U3826 (N_3826,N_3728,N_3703);
and U3827 (N_3827,N_3722,N_3731);
nand U3828 (N_3828,N_3745,N_3766);
or U3829 (N_3829,N_3700,N_3715);
or U3830 (N_3830,N_3705,N_3797);
and U3831 (N_3831,N_3712,N_3756);
nand U3832 (N_3832,N_3791,N_3767);
nor U3833 (N_3833,N_3755,N_3701);
nand U3834 (N_3834,N_3781,N_3762);
or U3835 (N_3835,N_3765,N_3753);
xor U3836 (N_3836,N_3751,N_3760);
and U3837 (N_3837,N_3723,N_3772);
nand U3838 (N_3838,N_3744,N_3794);
and U3839 (N_3839,N_3707,N_3742);
nor U3840 (N_3840,N_3774,N_3754);
nor U3841 (N_3841,N_3758,N_3782);
nor U3842 (N_3842,N_3764,N_3739);
and U3843 (N_3843,N_3733,N_3720);
and U3844 (N_3844,N_3789,N_3749);
or U3845 (N_3845,N_3778,N_3775);
nor U3846 (N_3846,N_3726,N_3768);
xor U3847 (N_3847,N_3777,N_3761);
nor U3848 (N_3848,N_3769,N_3732);
nand U3849 (N_3849,N_3706,N_3734);
nand U3850 (N_3850,N_3718,N_3743);
nand U3851 (N_3851,N_3727,N_3750);
nand U3852 (N_3852,N_3704,N_3793);
xor U3853 (N_3853,N_3727,N_3761);
nand U3854 (N_3854,N_3753,N_3792);
or U3855 (N_3855,N_3719,N_3754);
or U3856 (N_3856,N_3798,N_3706);
or U3857 (N_3857,N_3728,N_3758);
nor U3858 (N_3858,N_3728,N_3787);
nand U3859 (N_3859,N_3728,N_3707);
xnor U3860 (N_3860,N_3787,N_3790);
nor U3861 (N_3861,N_3773,N_3706);
and U3862 (N_3862,N_3765,N_3701);
nor U3863 (N_3863,N_3789,N_3704);
nor U3864 (N_3864,N_3732,N_3775);
nor U3865 (N_3865,N_3730,N_3759);
xor U3866 (N_3866,N_3765,N_3782);
nor U3867 (N_3867,N_3729,N_3787);
or U3868 (N_3868,N_3746,N_3793);
nor U3869 (N_3869,N_3713,N_3703);
and U3870 (N_3870,N_3781,N_3703);
nor U3871 (N_3871,N_3739,N_3726);
nor U3872 (N_3872,N_3704,N_3748);
and U3873 (N_3873,N_3756,N_3736);
nand U3874 (N_3874,N_3791,N_3766);
and U3875 (N_3875,N_3790,N_3706);
xor U3876 (N_3876,N_3775,N_3710);
and U3877 (N_3877,N_3757,N_3727);
xnor U3878 (N_3878,N_3739,N_3746);
or U3879 (N_3879,N_3736,N_3794);
xnor U3880 (N_3880,N_3737,N_3755);
and U3881 (N_3881,N_3765,N_3703);
or U3882 (N_3882,N_3768,N_3784);
and U3883 (N_3883,N_3755,N_3727);
nand U3884 (N_3884,N_3762,N_3772);
or U3885 (N_3885,N_3762,N_3740);
nor U3886 (N_3886,N_3784,N_3723);
nor U3887 (N_3887,N_3724,N_3775);
nand U3888 (N_3888,N_3753,N_3799);
nor U3889 (N_3889,N_3784,N_3738);
or U3890 (N_3890,N_3790,N_3750);
and U3891 (N_3891,N_3733,N_3740);
and U3892 (N_3892,N_3715,N_3751);
nand U3893 (N_3893,N_3741,N_3750);
and U3894 (N_3894,N_3706,N_3718);
nand U3895 (N_3895,N_3789,N_3706);
nand U3896 (N_3896,N_3730,N_3727);
nand U3897 (N_3897,N_3759,N_3750);
nor U3898 (N_3898,N_3737,N_3766);
or U3899 (N_3899,N_3713,N_3774);
nor U3900 (N_3900,N_3839,N_3854);
nand U3901 (N_3901,N_3898,N_3894);
nor U3902 (N_3902,N_3881,N_3802);
xor U3903 (N_3903,N_3870,N_3863);
nand U3904 (N_3904,N_3880,N_3812);
or U3905 (N_3905,N_3851,N_3869);
xor U3906 (N_3906,N_3836,N_3805);
nand U3907 (N_3907,N_3885,N_3819);
nand U3908 (N_3908,N_3865,N_3879);
and U3909 (N_3909,N_3821,N_3848);
xor U3910 (N_3910,N_3832,N_3893);
nor U3911 (N_3911,N_3842,N_3849);
nor U3912 (N_3912,N_3822,N_3878);
xor U3913 (N_3913,N_3871,N_3857);
nand U3914 (N_3914,N_3897,N_3824);
nor U3915 (N_3915,N_3872,N_3862);
xor U3916 (N_3916,N_3803,N_3856);
or U3917 (N_3917,N_3852,N_3874);
xnor U3918 (N_3918,N_3831,N_3886);
xnor U3919 (N_3919,N_3808,N_3841);
nor U3920 (N_3920,N_3835,N_3801);
or U3921 (N_3921,N_3888,N_3844);
xor U3922 (N_3922,N_3864,N_3800);
nand U3923 (N_3923,N_3833,N_3899);
nand U3924 (N_3924,N_3896,N_3818);
nand U3925 (N_3925,N_3887,N_3884);
nand U3926 (N_3926,N_3876,N_3814);
xor U3927 (N_3927,N_3866,N_3809);
xnor U3928 (N_3928,N_3807,N_3817);
nor U3929 (N_3929,N_3859,N_3875);
xor U3930 (N_3930,N_3837,N_3873);
xnor U3931 (N_3931,N_3811,N_3861);
xnor U3932 (N_3932,N_3813,N_3820);
nand U3933 (N_3933,N_3891,N_3892);
nand U3934 (N_3934,N_3882,N_3829);
and U3935 (N_3935,N_3868,N_3830);
nand U3936 (N_3936,N_3853,N_3858);
xnor U3937 (N_3937,N_3804,N_3816);
nor U3938 (N_3938,N_3850,N_3877);
xor U3939 (N_3939,N_3838,N_3867);
and U3940 (N_3940,N_3825,N_3855);
xor U3941 (N_3941,N_3890,N_3823);
and U3942 (N_3942,N_3815,N_3889);
xnor U3943 (N_3943,N_3895,N_3834);
or U3944 (N_3944,N_3828,N_3845);
or U3945 (N_3945,N_3827,N_3883);
or U3946 (N_3946,N_3846,N_3860);
nor U3947 (N_3947,N_3847,N_3810);
or U3948 (N_3948,N_3843,N_3826);
nor U3949 (N_3949,N_3840,N_3806);
nand U3950 (N_3950,N_3895,N_3827);
or U3951 (N_3951,N_3889,N_3858);
nor U3952 (N_3952,N_3884,N_3896);
and U3953 (N_3953,N_3829,N_3812);
nor U3954 (N_3954,N_3889,N_3899);
and U3955 (N_3955,N_3873,N_3883);
and U3956 (N_3956,N_3866,N_3814);
and U3957 (N_3957,N_3817,N_3857);
nand U3958 (N_3958,N_3866,N_3884);
xnor U3959 (N_3959,N_3841,N_3833);
and U3960 (N_3960,N_3810,N_3866);
nand U3961 (N_3961,N_3892,N_3889);
and U3962 (N_3962,N_3853,N_3886);
nor U3963 (N_3963,N_3853,N_3891);
nor U3964 (N_3964,N_3854,N_3860);
and U3965 (N_3965,N_3837,N_3881);
nor U3966 (N_3966,N_3854,N_3816);
and U3967 (N_3967,N_3845,N_3847);
and U3968 (N_3968,N_3807,N_3833);
nand U3969 (N_3969,N_3882,N_3811);
and U3970 (N_3970,N_3874,N_3829);
or U3971 (N_3971,N_3888,N_3813);
and U3972 (N_3972,N_3849,N_3819);
nor U3973 (N_3973,N_3836,N_3828);
xnor U3974 (N_3974,N_3812,N_3883);
nand U3975 (N_3975,N_3838,N_3808);
nand U3976 (N_3976,N_3811,N_3892);
and U3977 (N_3977,N_3871,N_3883);
nand U3978 (N_3978,N_3892,N_3809);
xnor U3979 (N_3979,N_3853,N_3816);
nor U3980 (N_3980,N_3872,N_3899);
nand U3981 (N_3981,N_3827,N_3896);
nand U3982 (N_3982,N_3826,N_3838);
nor U3983 (N_3983,N_3821,N_3875);
and U3984 (N_3984,N_3843,N_3807);
nor U3985 (N_3985,N_3864,N_3845);
nor U3986 (N_3986,N_3825,N_3873);
nand U3987 (N_3987,N_3877,N_3823);
and U3988 (N_3988,N_3890,N_3893);
or U3989 (N_3989,N_3895,N_3867);
nor U3990 (N_3990,N_3860,N_3896);
nor U3991 (N_3991,N_3826,N_3845);
or U3992 (N_3992,N_3896,N_3808);
or U3993 (N_3993,N_3896,N_3887);
and U3994 (N_3994,N_3875,N_3804);
and U3995 (N_3995,N_3863,N_3864);
nor U3996 (N_3996,N_3864,N_3891);
and U3997 (N_3997,N_3813,N_3869);
xor U3998 (N_3998,N_3870,N_3810);
xor U3999 (N_3999,N_3882,N_3836);
and U4000 (N_4000,N_3914,N_3975);
and U4001 (N_4001,N_3962,N_3900);
nand U4002 (N_4002,N_3907,N_3923);
nor U4003 (N_4003,N_3974,N_3927);
nor U4004 (N_4004,N_3904,N_3970);
nand U4005 (N_4005,N_3976,N_3950);
and U4006 (N_4006,N_3930,N_3973);
or U4007 (N_4007,N_3958,N_3906);
or U4008 (N_4008,N_3924,N_3965);
nor U4009 (N_4009,N_3933,N_3941);
xnor U4010 (N_4010,N_3917,N_3972);
nor U4011 (N_4011,N_3992,N_3919);
nand U4012 (N_4012,N_3912,N_3993);
xor U4013 (N_4013,N_3935,N_3959);
or U4014 (N_4014,N_3998,N_3934);
nor U4015 (N_4015,N_3925,N_3905);
or U4016 (N_4016,N_3978,N_3980);
nor U4017 (N_4017,N_3928,N_3951);
nand U4018 (N_4018,N_3915,N_3920);
and U4019 (N_4019,N_3945,N_3979);
nand U4020 (N_4020,N_3967,N_3916);
xnor U4021 (N_4021,N_3984,N_3942);
and U4022 (N_4022,N_3921,N_3968);
nor U4023 (N_4023,N_3903,N_3948);
and U4024 (N_4024,N_3955,N_3987);
xnor U4025 (N_4025,N_3909,N_3908);
nor U4026 (N_4026,N_3943,N_3902);
xnor U4027 (N_4027,N_3952,N_3956);
nand U4028 (N_4028,N_3989,N_3926);
nand U4029 (N_4029,N_3991,N_3938);
nor U4030 (N_4030,N_3957,N_3910);
or U4031 (N_4031,N_3981,N_3913);
or U4032 (N_4032,N_3990,N_3961);
nand U4033 (N_4033,N_3986,N_3944);
xnor U4034 (N_4034,N_3932,N_3947);
and U4035 (N_4035,N_3954,N_3922);
and U4036 (N_4036,N_3966,N_3994);
xor U4037 (N_4037,N_3988,N_3946);
and U4038 (N_4038,N_3982,N_3983);
nand U4039 (N_4039,N_3985,N_3901);
xnor U4040 (N_4040,N_3918,N_3971);
nor U4041 (N_4041,N_3995,N_3940);
and U4042 (N_4042,N_3911,N_3969);
or U4043 (N_4043,N_3977,N_3964);
nand U4044 (N_4044,N_3953,N_3960);
or U4045 (N_4045,N_3997,N_3931);
nor U4046 (N_4046,N_3936,N_3949);
or U4047 (N_4047,N_3963,N_3939);
nand U4048 (N_4048,N_3937,N_3929);
and U4049 (N_4049,N_3996,N_3999);
nor U4050 (N_4050,N_3944,N_3966);
nor U4051 (N_4051,N_3965,N_3960);
and U4052 (N_4052,N_3909,N_3931);
and U4053 (N_4053,N_3956,N_3995);
nand U4054 (N_4054,N_3942,N_3901);
and U4055 (N_4055,N_3911,N_3929);
and U4056 (N_4056,N_3994,N_3913);
and U4057 (N_4057,N_3951,N_3916);
nor U4058 (N_4058,N_3963,N_3999);
nor U4059 (N_4059,N_3990,N_3974);
or U4060 (N_4060,N_3948,N_3931);
nand U4061 (N_4061,N_3906,N_3933);
or U4062 (N_4062,N_3929,N_3987);
and U4063 (N_4063,N_3990,N_3976);
nand U4064 (N_4064,N_3900,N_3955);
or U4065 (N_4065,N_3958,N_3938);
or U4066 (N_4066,N_3973,N_3944);
xor U4067 (N_4067,N_3986,N_3938);
nand U4068 (N_4068,N_3996,N_3941);
and U4069 (N_4069,N_3965,N_3934);
nand U4070 (N_4070,N_3902,N_3977);
xor U4071 (N_4071,N_3973,N_3923);
nand U4072 (N_4072,N_3940,N_3926);
and U4073 (N_4073,N_3909,N_3942);
nand U4074 (N_4074,N_3945,N_3912);
nand U4075 (N_4075,N_3935,N_3972);
or U4076 (N_4076,N_3981,N_3959);
nor U4077 (N_4077,N_3906,N_3912);
and U4078 (N_4078,N_3984,N_3990);
xor U4079 (N_4079,N_3982,N_3957);
or U4080 (N_4080,N_3917,N_3971);
or U4081 (N_4081,N_3960,N_3934);
xor U4082 (N_4082,N_3986,N_3977);
and U4083 (N_4083,N_3970,N_3939);
nor U4084 (N_4084,N_3909,N_3900);
xor U4085 (N_4085,N_3932,N_3965);
or U4086 (N_4086,N_3961,N_3985);
and U4087 (N_4087,N_3907,N_3933);
or U4088 (N_4088,N_3999,N_3991);
nor U4089 (N_4089,N_3991,N_3929);
nand U4090 (N_4090,N_3931,N_3913);
nor U4091 (N_4091,N_3911,N_3928);
or U4092 (N_4092,N_3975,N_3932);
or U4093 (N_4093,N_3955,N_3994);
and U4094 (N_4094,N_3972,N_3986);
and U4095 (N_4095,N_3932,N_3959);
and U4096 (N_4096,N_3944,N_3901);
xnor U4097 (N_4097,N_3911,N_3903);
nand U4098 (N_4098,N_3901,N_3978);
or U4099 (N_4099,N_3962,N_3998);
xor U4100 (N_4100,N_4046,N_4090);
nand U4101 (N_4101,N_4028,N_4018);
or U4102 (N_4102,N_4013,N_4052);
nor U4103 (N_4103,N_4086,N_4032);
nand U4104 (N_4104,N_4008,N_4036);
and U4105 (N_4105,N_4085,N_4055);
nor U4106 (N_4106,N_4014,N_4084);
nand U4107 (N_4107,N_4095,N_4062);
and U4108 (N_4108,N_4026,N_4057);
and U4109 (N_4109,N_4082,N_4031);
xor U4110 (N_4110,N_4078,N_4045);
and U4111 (N_4111,N_4049,N_4060);
nor U4112 (N_4112,N_4071,N_4012);
xnor U4113 (N_4113,N_4048,N_4068);
or U4114 (N_4114,N_4065,N_4038);
xor U4115 (N_4115,N_4081,N_4043);
nor U4116 (N_4116,N_4005,N_4030);
or U4117 (N_4117,N_4088,N_4070);
nor U4118 (N_4118,N_4039,N_4025);
or U4119 (N_4119,N_4000,N_4044);
nor U4120 (N_4120,N_4067,N_4047);
or U4121 (N_4121,N_4034,N_4075);
and U4122 (N_4122,N_4011,N_4015);
nor U4123 (N_4123,N_4042,N_4007);
xor U4124 (N_4124,N_4053,N_4041);
nand U4125 (N_4125,N_4072,N_4097);
nand U4126 (N_4126,N_4077,N_4096);
or U4127 (N_4127,N_4058,N_4087);
or U4128 (N_4128,N_4017,N_4033);
nand U4129 (N_4129,N_4069,N_4054);
nand U4130 (N_4130,N_4092,N_4024);
or U4131 (N_4131,N_4091,N_4021);
nand U4132 (N_4132,N_4073,N_4094);
and U4133 (N_4133,N_4037,N_4083);
and U4134 (N_4134,N_4051,N_4050);
nor U4135 (N_4135,N_4035,N_4020);
xnor U4136 (N_4136,N_4040,N_4001);
xor U4137 (N_4137,N_4006,N_4029);
and U4138 (N_4138,N_4009,N_4063);
nand U4139 (N_4139,N_4064,N_4059);
xnor U4140 (N_4140,N_4019,N_4002);
xor U4141 (N_4141,N_4004,N_4093);
xor U4142 (N_4142,N_4061,N_4016);
nor U4143 (N_4143,N_4099,N_4056);
nand U4144 (N_4144,N_4080,N_4022);
nand U4145 (N_4145,N_4023,N_4027);
and U4146 (N_4146,N_4076,N_4066);
and U4147 (N_4147,N_4010,N_4003);
and U4148 (N_4148,N_4079,N_4074);
and U4149 (N_4149,N_4098,N_4089);
nor U4150 (N_4150,N_4050,N_4034);
xnor U4151 (N_4151,N_4097,N_4073);
and U4152 (N_4152,N_4092,N_4002);
xnor U4153 (N_4153,N_4079,N_4093);
nand U4154 (N_4154,N_4078,N_4038);
xor U4155 (N_4155,N_4033,N_4042);
xor U4156 (N_4156,N_4056,N_4015);
and U4157 (N_4157,N_4014,N_4015);
xnor U4158 (N_4158,N_4071,N_4059);
and U4159 (N_4159,N_4038,N_4020);
nand U4160 (N_4160,N_4060,N_4008);
nand U4161 (N_4161,N_4062,N_4082);
xnor U4162 (N_4162,N_4047,N_4001);
xnor U4163 (N_4163,N_4000,N_4095);
and U4164 (N_4164,N_4039,N_4070);
and U4165 (N_4165,N_4028,N_4040);
nand U4166 (N_4166,N_4080,N_4049);
nand U4167 (N_4167,N_4022,N_4026);
xor U4168 (N_4168,N_4038,N_4058);
nor U4169 (N_4169,N_4091,N_4006);
nand U4170 (N_4170,N_4036,N_4010);
nor U4171 (N_4171,N_4061,N_4095);
or U4172 (N_4172,N_4077,N_4055);
xor U4173 (N_4173,N_4051,N_4048);
or U4174 (N_4174,N_4000,N_4066);
xor U4175 (N_4175,N_4015,N_4090);
nor U4176 (N_4176,N_4056,N_4022);
or U4177 (N_4177,N_4066,N_4014);
xnor U4178 (N_4178,N_4033,N_4044);
or U4179 (N_4179,N_4030,N_4056);
and U4180 (N_4180,N_4058,N_4085);
nor U4181 (N_4181,N_4092,N_4093);
or U4182 (N_4182,N_4051,N_4040);
or U4183 (N_4183,N_4037,N_4023);
or U4184 (N_4184,N_4066,N_4018);
and U4185 (N_4185,N_4004,N_4094);
and U4186 (N_4186,N_4080,N_4027);
nor U4187 (N_4187,N_4041,N_4025);
nand U4188 (N_4188,N_4070,N_4085);
xnor U4189 (N_4189,N_4033,N_4074);
nand U4190 (N_4190,N_4076,N_4024);
and U4191 (N_4191,N_4068,N_4003);
xor U4192 (N_4192,N_4016,N_4022);
nor U4193 (N_4193,N_4018,N_4059);
xnor U4194 (N_4194,N_4072,N_4044);
nand U4195 (N_4195,N_4008,N_4028);
xnor U4196 (N_4196,N_4021,N_4037);
xnor U4197 (N_4197,N_4090,N_4076);
nand U4198 (N_4198,N_4040,N_4067);
xor U4199 (N_4199,N_4054,N_4055);
or U4200 (N_4200,N_4109,N_4120);
xor U4201 (N_4201,N_4124,N_4149);
and U4202 (N_4202,N_4178,N_4165);
or U4203 (N_4203,N_4188,N_4127);
or U4204 (N_4204,N_4183,N_4162);
nand U4205 (N_4205,N_4155,N_4131);
nor U4206 (N_4206,N_4139,N_4176);
nand U4207 (N_4207,N_4170,N_4153);
and U4208 (N_4208,N_4186,N_4159);
xnor U4209 (N_4209,N_4108,N_4166);
xor U4210 (N_4210,N_4100,N_4177);
or U4211 (N_4211,N_4194,N_4154);
nand U4212 (N_4212,N_4101,N_4156);
xor U4213 (N_4213,N_4195,N_4163);
xor U4214 (N_4214,N_4110,N_4142);
and U4215 (N_4215,N_4121,N_4116);
and U4216 (N_4216,N_4168,N_4160);
nand U4217 (N_4217,N_4126,N_4191);
xnor U4218 (N_4218,N_4129,N_4118);
xor U4219 (N_4219,N_4128,N_4196);
and U4220 (N_4220,N_4179,N_4117);
nor U4221 (N_4221,N_4187,N_4190);
or U4222 (N_4222,N_4173,N_4122);
and U4223 (N_4223,N_4140,N_4198);
or U4224 (N_4224,N_4134,N_4161);
nand U4225 (N_4225,N_4169,N_4180);
or U4226 (N_4226,N_4146,N_4112);
xor U4227 (N_4227,N_4103,N_4147);
or U4228 (N_4228,N_4123,N_4184);
or U4229 (N_4229,N_4164,N_4137);
and U4230 (N_4230,N_4125,N_4175);
xnor U4231 (N_4231,N_4152,N_4114);
xor U4232 (N_4232,N_4182,N_4148);
nand U4233 (N_4233,N_4141,N_4158);
nor U4234 (N_4234,N_4130,N_4133);
and U4235 (N_4235,N_4171,N_4105);
nor U4236 (N_4236,N_4150,N_4151);
and U4237 (N_4237,N_4157,N_4115);
nor U4238 (N_4238,N_4104,N_4143);
or U4239 (N_4239,N_4138,N_4181);
and U4240 (N_4240,N_4192,N_4135);
nand U4241 (N_4241,N_4102,N_4193);
nor U4242 (N_4242,N_4197,N_4174);
xor U4243 (N_4243,N_4106,N_4199);
nand U4244 (N_4244,N_4144,N_4107);
xnor U4245 (N_4245,N_4119,N_4113);
xnor U4246 (N_4246,N_4185,N_4111);
and U4247 (N_4247,N_4189,N_4172);
xor U4248 (N_4248,N_4136,N_4167);
nand U4249 (N_4249,N_4145,N_4132);
nand U4250 (N_4250,N_4106,N_4115);
and U4251 (N_4251,N_4195,N_4118);
or U4252 (N_4252,N_4143,N_4137);
nand U4253 (N_4253,N_4108,N_4146);
xor U4254 (N_4254,N_4174,N_4159);
or U4255 (N_4255,N_4154,N_4177);
nand U4256 (N_4256,N_4180,N_4136);
or U4257 (N_4257,N_4151,N_4125);
xnor U4258 (N_4258,N_4101,N_4181);
xnor U4259 (N_4259,N_4146,N_4145);
nand U4260 (N_4260,N_4131,N_4122);
or U4261 (N_4261,N_4117,N_4183);
or U4262 (N_4262,N_4188,N_4153);
xor U4263 (N_4263,N_4134,N_4190);
xnor U4264 (N_4264,N_4164,N_4161);
or U4265 (N_4265,N_4143,N_4187);
or U4266 (N_4266,N_4161,N_4120);
and U4267 (N_4267,N_4109,N_4171);
nand U4268 (N_4268,N_4170,N_4119);
nor U4269 (N_4269,N_4154,N_4196);
nand U4270 (N_4270,N_4107,N_4170);
xor U4271 (N_4271,N_4167,N_4117);
or U4272 (N_4272,N_4147,N_4144);
nor U4273 (N_4273,N_4129,N_4148);
nand U4274 (N_4274,N_4196,N_4116);
nand U4275 (N_4275,N_4106,N_4114);
nand U4276 (N_4276,N_4185,N_4136);
nand U4277 (N_4277,N_4130,N_4160);
nor U4278 (N_4278,N_4189,N_4166);
nor U4279 (N_4279,N_4162,N_4170);
xnor U4280 (N_4280,N_4168,N_4173);
nand U4281 (N_4281,N_4121,N_4162);
nor U4282 (N_4282,N_4139,N_4180);
xnor U4283 (N_4283,N_4175,N_4118);
and U4284 (N_4284,N_4192,N_4179);
or U4285 (N_4285,N_4194,N_4117);
nor U4286 (N_4286,N_4117,N_4168);
and U4287 (N_4287,N_4140,N_4163);
nor U4288 (N_4288,N_4197,N_4156);
and U4289 (N_4289,N_4109,N_4189);
xnor U4290 (N_4290,N_4196,N_4195);
and U4291 (N_4291,N_4108,N_4132);
xor U4292 (N_4292,N_4123,N_4110);
and U4293 (N_4293,N_4112,N_4159);
nand U4294 (N_4294,N_4153,N_4115);
nand U4295 (N_4295,N_4123,N_4162);
nand U4296 (N_4296,N_4129,N_4177);
or U4297 (N_4297,N_4134,N_4126);
nand U4298 (N_4298,N_4164,N_4132);
or U4299 (N_4299,N_4107,N_4199);
xnor U4300 (N_4300,N_4221,N_4206);
nor U4301 (N_4301,N_4226,N_4248);
nor U4302 (N_4302,N_4294,N_4210);
nor U4303 (N_4303,N_4266,N_4202);
xor U4304 (N_4304,N_4219,N_4235);
nor U4305 (N_4305,N_4233,N_4203);
and U4306 (N_4306,N_4220,N_4222);
nor U4307 (N_4307,N_4262,N_4258);
nor U4308 (N_4308,N_4291,N_4256);
xor U4309 (N_4309,N_4289,N_4265);
and U4310 (N_4310,N_4243,N_4251);
or U4311 (N_4311,N_4255,N_4298);
xor U4312 (N_4312,N_4282,N_4295);
and U4313 (N_4313,N_4259,N_4254);
xnor U4314 (N_4314,N_4275,N_4253);
xnor U4315 (N_4315,N_4238,N_4237);
and U4316 (N_4316,N_4250,N_4272);
xor U4317 (N_4317,N_4276,N_4216);
or U4318 (N_4318,N_4278,N_4269);
or U4319 (N_4319,N_4234,N_4242);
and U4320 (N_4320,N_4299,N_4244);
and U4321 (N_4321,N_4209,N_4252);
nand U4322 (N_4322,N_4261,N_4270);
or U4323 (N_4323,N_4285,N_4231);
nor U4324 (N_4324,N_4263,N_4200);
nand U4325 (N_4325,N_4207,N_4229);
xnor U4326 (N_4326,N_4287,N_4230);
or U4327 (N_4327,N_4296,N_4271);
nor U4328 (N_4328,N_4267,N_4260);
nor U4329 (N_4329,N_4236,N_4218);
xor U4330 (N_4330,N_4212,N_4264);
nand U4331 (N_4331,N_4293,N_4249);
and U4332 (N_4332,N_4292,N_4224);
and U4333 (N_4333,N_4227,N_4273);
nor U4334 (N_4334,N_4257,N_4247);
nand U4335 (N_4335,N_4201,N_4217);
xor U4336 (N_4336,N_4239,N_4240);
or U4337 (N_4337,N_4245,N_4277);
nor U4338 (N_4338,N_4283,N_4225);
or U4339 (N_4339,N_4241,N_4215);
nor U4340 (N_4340,N_4204,N_4290);
and U4341 (N_4341,N_4213,N_4284);
nor U4342 (N_4342,N_4281,N_4205);
or U4343 (N_4343,N_4214,N_4232);
nor U4344 (N_4344,N_4274,N_4288);
and U4345 (N_4345,N_4286,N_4223);
nand U4346 (N_4346,N_4211,N_4280);
xnor U4347 (N_4347,N_4268,N_4246);
and U4348 (N_4348,N_4208,N_4297);
xor U4349 (N_4349,N_4228,N_4279);
xnor U4350 (N_4350,N_4224,N_4211);
nand U4351 (N_4351,N_4290,N_4285);
or U4352 (N_4352,N_4255,N_4256);
nor U4353 (N_4353,N_4205,N_4285);
and U4354 (N_4354,N_4270,N_4259);
or U4355 (N_4355,N_4264,N_4200);
or U4356 (N_4356,N_4290,N_4263);
nand U4357 (N_4357,N_4296,N_4259);
nand U4358 (N_4358,N_4274,N_4294);
nand U4359 (N_4359,N_4201,N_4279);
xnor U4360 (N_4360,N_4204,N_4264);
xnor U4361 (N_4361,N_4298,N_4280);
xnor U4362 (N_4362,N_4252,N_4278);
xnor U4363 (N_4363,N_4233,N_4216);
nand U4364 (N_4364,N_4223,N_4290);
xnor U4365 (N_4365,N_4250,N_4211);
nor U4366 (N_4366,N_4291,N_4257);
or U4367 (N_4367,N_4208,N_4293);
xnor U4368 (N_4368,N_4258,N_4239);
and U4369 (N_4369,N_4218,N_4245);
or U4370 (N_4370,N_4249,N_4226);
nand U4371 (N_4371,N_4299,N_4256);
xnor U4372 (N_4372,N_4212,N_4238);
and U4373 (N_4373,N_4289,N_4261);
nor U4374 (N_4374,N_4244,N_4213);
nor U4375 (N_4375,N_4229,N_4230);
and U4376 (N_4376,N_4246,N_4260);
nor U4377 (N_4377,N_4228,N_4217);
or U4378 (N_4378,N_4263,N_4213);
or U4379 (N_4379,N_4286,N_4299);
or U4380 (N_4380,N_4259,N_4220);
nand U4381 (N_4381,N_4204,N_4223);
nand U4382 (N_4382,N_4206,N_4286);
xor U4383 (N_4383,N_4243,N_4212);
and U4384 (N_4384,N_4280,N_4228);
xnor U4385 (N_4385,N_4249,N_4254);
xnor U4386 (N_4386,N_4235,N_4262);
xor U4387 (N_4387,N_4208,N_4214);
xor U4388 (N_4388,N_4294,N_4284);
nor U4389 (N_4389,N_4236,N_4234);
xnor U4390 (N_4390,N_4228,N_4273);
and U4391 (N_4391,N_4205,N_4223);
nand U4392 (N_4392,N_4275,N_4248);
nand U4393 (N_4393,N_4297,N_4292);
xnor U4394 (N_4394,N_4286,N_4215);
or U4395 (N_4395,N_4274,N_4271);
and U4396 (N_4396,N_4219,N_4244);
nand U4397 (N_4397,N_4220,N_4243);
nand U4398 (N_4398,N_4291,N_4263);
or U4399 (N_4399,N_4271,N_4248);
or U4400 (N_4400,N_4396,N_4321);
or U4401 (N_4401,N_4311,N_4309);
nand U4402 (N_4402,N_4350,N_4338);
or U4403 (N_4403,N_4331,N_4381);
nor U4404 (N_4404,N_4335,N_4319);
nand U4405 (N_4405,N_4384,N_4365);
nor U4406 (N_4406,N_4351,N_4395);
xnor U4407 (N_4407,N_4370,N_4306);
nor U4408 (N_4408,N_4393,N_4379);
or U4409 (N_4409,N_4383,N_4356);
xnor U4410 (N_4410,N_4367,N_4334);
and U4411 (N_4411,N_4374,N_4312);
nor U4412 (N_4412,N_4389,N_4394);
nor U4413 (N_4413,N_4308,N_4387);
and U4414 (N_4414,N_4346,N_4352);
nor U4415 (N_4415,N_4324,N_4382);
or U4416 (N_4416,N_4300,N_4342);
and U4417 (N_4417,N_4398,N_4375);
xnor U4418 (N_4418,N_4315,N_4337);
or U4419 (N_4419,N_4327,N_4318);
or U4420 (N_4420,N_4307,N_4361);
nor U4421 (N_4421,N_4316,N_4380);
xor U4422 (N_4422,N_4397,N_4344);
or U4423 (N_4423,N_4371,N_4386);
nand U4424 (N_4424,N_4343,N_4364);
or U4425 (N_4425,N_4330,N_4328);
nor U4426 (N_4426,N_4303,N_4388);
or U4427 (N_4427,N_4317,N_4329);
nand U4428 (N_4428,N_4368,N_4349);
nor U4429 (N_4429,N_4310,N_4376);
or U4430 (N_4430,N_4341,N_4326);
nor U4431 (N_4431,N_4348,N_4345);
xor U4432 (N_4432,N_4304,N_4392);
nor U4433 (N_4433,N_4357,N_4360);
nand U4434 (N_4434,N_4372,N_4320);
xor U4435 (N_4435,N_4391,N_4333);
xnor U4436 (N_4436,N_4377,N_4313);
or U4437 (N_4437,N_4323,N_4325);
or U4438 (N_4438,N_4390,N_4358);
and U4439 (N_4439,N_4332,N_4362);
nor U4440 (N_4440,N_4339,N_4359);
nor U4441 (N_4441,N_4353,N_4347);
and U4442 (N_4442,N_4354,N_4369);
nor U4443 (N_4443,N_4355,N_4363);
xnor U4444 (N_4444,N_4385,N_4366);
nand U4445 (N_4445,N_4302,N_4340);
and U4446 (N_4446,N_4373,N_4378);
nor U4447 (N_4447,N_4305,N_4399);
nand U4448 (N_4448,N_4314,N_4301);
nor U4449 (N_4449,N_4322,N_4336);
nor U4450 (N_4450,N_4315,N_4303);
and U4451 (N_4451,N_4326,N_4353);
or U4452 (N_4452,N_4334,N_4375);
nand U4453 (N_4453,N_4353,N_4349);
xnor U4454 (N_4454,N_4302,N_4338);
nand U4455 (N_4455,N_4396,N_4380);
or U4456 (N_4456,N_4377,N_4370);
and U4457 (N_4457,N_4309,N_4332);
xor U4458 (N_4458,N_4322,N_4341);
or U4459 (N_4459,N_4359,N_4390);
or U4460 (N_4460,N_4363,N_4319);
nor U4461 (N_4461,N_4321,N_4367);
or U4462 (N_4462,N_4339,N_4374);
or U4463 (N_4463,N_4394,N_4323);
xor U4464 (N_4464,N_4341,N_4354);
xnor U4465 (N_4465,N_4382,N_4339);
or U4466 (N_4466,N_4326,N_4398);
or U4467 (N_4467,N_4388,N_4395);
nand U4468 (N_4468,N_4307,N_4304);
xor U4469 (N_4469,N_4380,N_4381);
nor U4470 (N_4470,N_4378,N_4300);
nor U4471 (N_4471,N_4343,N_4362);
nor U4472 (N_4472,N_4347,N_4373);
nand U4473 (N_4473,N_4359,N_4371);
and U4474 (N_4474,N_4329,N_4343);
nand U4475 (N_4475,N_4333,N_4394);
nand U4476 (N_4476,N_4327,N_4361);
or U4477 (N_4477,N_4304,N_4341);
nor U4478 (N_4478,N_4326,N_4376);
xor U4479 (N_4479,N_4391,N_4376);
xor U4480 (N_4480,N_4382,N_4327);
nor U4481 (N_4481,N_4384,N_4380);
and U4482 (N_4482,N_4388,N_4309);
nor U4483 (N_4483,N_4389,N_4309);
xnor U4484 (N_4484,N_4350,N_4342);
and U4485 (N_4485,N_4367,N_4370);
xnor U4486 (N_4486,N_4347,N_4374);
or U4487 (N_4487,N_4385,N_4356);
and U4488 (N_4488,N_4313,N_4330);
or U4489 (N_4489,N_4365,N_4305);
nor U4490 (N_4490,N_4393,N_4314);
or U4491 (N_4491,N_4394,N_4352);
nand U4492 (N_4492,N_4351,N_4325);
or U4493 (N_4493,N_4348,N_4306);
or U4494 (N_4494,N_4370,N_4371);
or U4495 (N_4495,N_4371,N_4383);
or U4496 (N_4496,N_4332,N_4325);
nand U4497 (N_4497,N_4335,N_4314);
nor U4498 (N_4498,N_4320,N_4361);
nor U4499 (N_4499,N_4327,N_4354);
nor U4500 (N_4500,N_4419,N_4470);
xnor U4501 (N_4501,N_4446,N_4437);
or U4502 (N_4502,N_4469,N_4456);
and U4503 (N_4503,N_4421,N_4402);
or U4504 (N_4504,N_4452,N_4435);
xor U4505 (N_4505,N_4492,N_4494);
or U4506 (N_4506,N_4490,N_4480);
nor U4507 (N_4507,N_4409,N_4444);
and U4508 (N_4508,N_4415,N_4481);
nand U4509 (N_4509,N_4491,N_4445);
and U4510 (N_4510,N_4476,N_4432);
or U4511 (N_4511,N_4431,N_4475);
nand U4512 (N_4512,N_4451,N_4403);
or U4513 (N_4513,N_4493,N_4464);
xor U4514 (N_4514,N_4457,N_4441);
nor U4515 (N_4515,N_4420,N_4448);
or U4516 (N_4516,N_4449,N_4414);
or U4517 (N_4517,N_4404,N_4473);
or U4518 (N_4518,N_4425,N_4472);
and U4519 (N_4519,N_4474,N_4416);
xor U4520 (N_4520,N_4422,N_4427);
or U4521 (N_4521,N_4467,N_4401);
xor U4522 (N_4522,N_4486,N_4488);
nor U4523 (N_4523,N_4466,N_4418);
or U4524 (N_4524,N_4482,N_4462);
nor U4525 (N_4525,N_4450,N_4417);
xnor U4526 (N_4526,N_4413,N_4436);
nand U4527 (N_4527,N_4430,N_4463);
xor U4528 (N_4528,N_4405,N_4406);
xnor U4529 (N_4529,N_4411,N_4447);
or U4530 (N_4530,N_4438,N_4489);
or U4531 (N_4531,N_4433,N_4455);
nand U4532 (N_4532,N_4407,N_4408);
and U4533 (N_4533,N_4412,N_4468);
xnor U4534 (N_4534,N_4483,N_4428);
xnor U4535 (N_4535,N_4495,N_4498);
and U4536 (N_4536,N_4461,N_4477);
nor U4537 (N_4537,N_4423,N_4479);
or U4538 (N_4538,N_4460,N_4429);
nor U4539 (N_4539,N_4484,N_4442);
nor U4540 (N_4540,N_4496,N_4426);
or U4541 (N_4541,N_4497,N_4453);
nand U4542 (N_4542,N_4439,N_4485);
nor U4543 (N_4543,N_4454,N_4440);
xnor U4544 (N_4544,N_4487,N_4458);
nor U4545 (N_4545,N_4400,N_4465);
nand U4546 (N_4546,N_4424,N_4471);
nand U4547 (N_4547,N_4499,N_4478);
nand U4548 (N_4548,N_4459,N_4434);
nand U4549 (N_4549,N_4443,N_4410);
xnor U4550 (N_4550,N_4450,N_4478);
nor U4551 (N_4551,N_4456,N_4425);
nor U4552 (N_4552,N_4455,N_4447);
or U4553 (N_4553,N_4458,N_4431);
nand U4554 (N_4554,N_4471,N_4485);
and U4555 (N_4555,N_4439,N_4492);
nand U4556 (N_4556,N_4489,N_4499);
nor U4557 (N_4557,N_4434,N_4452);
nor U4558 (N_4558,N_4456,N_4415);
xor U4559 (N_4559,N_4472,N_4428);
nor U4560 (N_4560,N_4459,N_4467);
nand U4561 (N_4561,N_4482,N_4449);
xor U4562 (N_4562,N_4482,N_4489);
nand U4563 (N_4563,N_4444,N_4428);
xnor U4564 (N_4564,N_4413,N_4402);
and U4565 (N_4565,N_4477,N_4493);
and U4566 (N_4566,N_4441,N_4481);
xnor U4567 (N_4567,N_4468,N_4422);
nand U4568 (N_4568,N_4495,N_4475);
nand U4569 (N_4569,N_4403,N_4475);
xnor U4570 (N_4570,N_4467,N_4447);
nor U4571 (N_4571,N_4442,N_4497);
nand U4572 (N_4572,N_4481,N_4430);
nor U4573 (N_4573,N_4454,N_4410);
xor U4574 (N_4574,N_4426,N_4473);
xnor U4575 (N_4575,N_4422,N_4451);
nand U4576 (N_4576,N_4421,N_4468);
xnor U4577 (N_4577,N_4443,N_4447);
or U4578 (N_4578,N_4415,N_4492);
xnor U4579 (N_4579,N_4482,N_4444);
xor U4580 (N_4580,N_4476,N_4496);
nand U4581 (N_4581,N_4457,N_4469);
and U4582 (N_4582,N_4492,N_4436);
nor U4583 (N_4583,N_4439,N_4483);
and U4584 (N_4584,N_4485,N_4450);
nand U4585 (N_4585,N_4407,N_4418);
and U4586 (N_4586,N_4490,N_4410);
or U4587 (N_4587,N_4402,N_4415);
xnor U4588 (N_4588,N_4443,N_4409);
nand U4589 (N_4589,N_4435,N_4432);
nor U4590 (N_4590,N_4405,N_4441);
or U4591 (N_4591,N_4447,N_4489);
xor U4592 (N_4592,N_4400,N_4479);
nand U4593 (N_4593,N_4440,N_4407);
and U4594 (N_4594,N_4458,N_4473);
xor U4595 (N_4595,N_4423,N_4486);
and U4596 (N_4596,N_4440,N_4474);
and U4597 (N_4597,N_4495,N_4425);
xnor U4598 (N_4598,N_4488,N_4423);
xnor U4599 (N_4599,N_4424,N_4485);
or U4600 (N_4600,N_4577,N_4598);
xor U4601 (N_4601,N_4560,N_4515);
nand U4602 (N_4602,N_4591,N_4562);
and U4603 (N_4603,N_4569,N_4536);
and U4604 (N_4604,N_4584,N_4595);
and U4605 (N_4605,N_4578,N_4558);
nor U4606 (N_4606,N_4544,N_4583);
nand U4607 (N_4607,N_4561,N_4573);
and U4608 (N_4608,N_4597,N_4537);
nor U4609 (N_4609,N_4514,N_4535);
nand U4610 (N_4610,N_4543,N_4516);
or U4611 (N_4611,N_4522,N_4590);
xnor U4612 (N_4612,N_4545,N_4556);
or U4613 (N_4613,N_4581,N_4593);
and U4614 (N_4614,N_4504,N_4576);
xnor U4615 (N_4615,N_4534,N_4575);
or U4616 (N_4616,N_4570,N_4566);
and U4617 (N_4617,N_4518,N_4507);
xnor U4618 (N_4618,N_4555,N_4553);
xnor U4619 (N_4619,N_4525,N_4547);
and U4620 (N_4620,N_4502,N_4513);
nor U4621 (N_4621,N_4559,N_4585);
nand U4622 (N_4622,N_4511,N_4509);
nor U4623 (N_4623,N_4557,N_4538);
xnor U4624 (N_4624,N_4524,N_4550);
xnor U4625 (N_4625,N_4568,N_4512);
xor U4626 (N_4626,N_4526,N_4529);
xor U4627 (N_4627,N_4554,N_4542);
xor U4628 (N_4628,N_4564,N_4549);
nor U4629 (N_4629,N_4588,N_4563);
nor U4630 (N_4630,N_4586,N_4589);
nor U4631 (N_4631,N_4587,N_4527);
nand U4632 (N_4632,N_4596,N_4531);
or U4633 (N_4633,N_4539,N_4533);
nand U4634 (N_4634,N_4551,N_4520);
or U4635 (N_4635,N_4506,N_4574);
and U4636 (N_4636,N_4517,N_4508);
and U4637 (N_4637,N_4565,N_4572);
or U4638 (N_4638,N_4532,N_4580);
xor U4639 (N_4639,N_4503,N_4530);
and U4640 (N_4640,N_4528,N_4552);
and U4641 (N_4641,N_4519,N_4505);
and U4642 (N_4642,N_4582,N_4541);
xor U4643 (N_4643,N_4523,N_4500);
and U4644 (N_4644,N_4592,N_4599);
nand U4645 (N_4645,N_4521,N_4594);
nor U4646 (N_4646,N_4567,N_4510);
xor U4647 (N_4647,N_4501,N_4548);
xor U4648 (N_4648,N_4546,N_4540);
nand U4649 (N_4649,N_4579,N_4571);
and U4650 (N_4650,N_4558,N_4512);
xor U4651 (N_4651,N_4510,N_4562);
xor U4652 (N_4652,N_4551,N_4584);
xor U4653 (N_4653,N_4563,N_4566);
or U4654 (N_4654,N_4501,N_4520);
nand U4655 (N_4655,N_4534,N_4512);
nor U4656 (N_4656,N_4564,N_4521);
and U4657 (N_4657,N_4574,N_4535);
nand U4658 (N_4658,N_4584,N_4581);
xnor U4659 (N_4659,N_4533,N_4516);
xor U4660 (N_4660,N_4599,N_4559);
or U4661 (N_4661,N_4589,N_4564);
nand U4662 (N_4662,N_4514,N_4529);
xor U4663 (N_4663,N_4569,N_4592);
and U4664 (N_4664,N_4542,N_4516);
and U4665 (N_4665,N_4558,N_4568);
xnor U4666 (N_4666,N_4567,N_4555);
nor U4667 (N_4667,N_4576,N_4510);
or U4668 (N_4668,N_4561,N_4532);
or U4669 (N_4669,N_4539,N_4538);
nand U4670 (N_4670,N_4575,N_4580);
and U4671 (N_4671,N_4577,N_4546);
xnor U4672 (N_4672,N_4599,N_4525);
nor U4673 (N_4673,N_4538,N_4544);
and U4674 (N_4674,N_4589,N_4585);
xor U4675 (N_4675,N_4535,N_4517);
and U4676 (N_4676,N_4550,N_4569);
nand U4677 (N_4677,N_4549,N_4557);
and U4678 (N_4678,N_4549,N_4595);
xnor U4679 (N_4679,N_4519,N_4522);
and U4680 (N_4680,N_4576,N_4596);
nor U4681 (N_4681,N_4508,N_4574);
nand U4682 (N_4682,N_4540,N_4579);
nor U4683 (N_4683,N_4519,N_4558);
and U4684 (N_4684,N_4521,N_4584);
or U4685 (N_4685,N_4557,N_4579);
or U4686 (N_4686,N_4546,N_4508);
nand U4687 (N_4687,N_4515,N_4503);
nor U4688 (N_4688,N_4569,N_4546);
and U4689 (N_4689,N_4557,N_4531);
nor U4690 (N_4690,N_4599,N_4560);
and U4691 (N_4691,N_4539,N_4514);
nor U4692 (N_4692,N_4558,N_4505);
or U4693 (N_4693,N_4561,N_4520);
and U4694 (N_4694,N_4533,N_4528);
and U4695 (N_4695,N_4585,N_4512);
or U4696 (N_4696,N_4577,N_4557);
and U4697 (N_4697,N_4500,N_4576);
nand U4698 (N_4698,N_4555,N_4575);
and U4699 (N_4699,N_4543,N_4526);
and U4700 (N_4700,N_4690,N_4627);
or U4701 (N_4701,N_4671,N_4635);
or U4702 (N_4702,N_4644,N_4674);
xnor U4703 (N_4703,N_4633,N_4666);
and U4704 (N_4704,N_4626,N_4613);
nand U4705 (N_4705,N_4637,N_4602);
and U4706 (N_4706,N_4614,N_4618);
or U4707 (N_4707,N_4696,N_4632);
xnor U4708 (N_4708,N_4649,N_4663);
or U4709 (N_4709,N_4641,N_4628);
nand U4710 (N_4710,N_4651,N_4697);
or U4711 (N_4711,N_4642,N_4630);
xnor U4712 (N_4712,N_4678,N_4662);
or U4713 (N_4713,N_4619,N_4694);
or U4714 (N_4714,N_4673,N_4668);
nand U4715 (N_4715,N_4615,N_4681);
and U4716 (N_4716,N_4600,N_4616);
nor U4717 (N_4717,N_4617,N_4634);
or U4718 (N_4718,N_4623,N_4654);
or U4719 (N_4719,N_4604,N_4687);
nand U4720 (N_4720,N_4689,N_4609);
nand U4721 (N_4721,N_4698,N_4661);
and U4722 (N_4722,N_4640,N_4659);
and U4723 (N_4723,N_4670,N_4647);
xnor U4724 (N_4724,N_4691,N_4682);
xnor U4725 (N_4725,N_4692,N_4629);
nor U4726 (N_4726,N_4639,N_4605);
xnor U4727 (N_4727,N_4652,N_4675);
nor U4728 (N_4728,N_4610,N_4693);
and U4729 (N_4729,N_4669,N_4636);
or U4730 (N_4730,N_4665,N_4672);
and U4731 (N_4731,N_4631,N_4608);
xor U4732 (N_4732,N_4603,N_4664);
or U4733 (N_4733,N_4601,N_4653);
xor U4734 (N_4734,N_4685,N_4650);
and U4735 (N_4735,N_4680,N_4622);
or U4736 (N_4736,N_4679,N_4658);
xor U4737 (N_4737,N_4612,N_4677);
or U4738 (N_4738,N_4646,N_4621);
nor U4739 (N_4739,N_4638,N_4660);
nor U4740 (N_4740,N_4656,N_4645);
and U4741 (N_4741,N_4686,N_4657);
or U4742 (N_4742,N_4676,N_4625);
xor U4743 (N_4743,N_4607,N_4620);
nor U4744 (N_4744,N_4667,N_4606);
nor U4745 (N_4745,N_4648,N_4684);
xor U4746 (N_4746,N_4624,N_4611);
xor U4747 (N_4747,N_4695,N_4683);
nor U4748 (N_4748,N_4655,N_4699);
nor U4749 (N_4749,N_4643,N_4688);
xor U4750 (N_4750,N_4662,N_4644);
nand U4751 (N_4751,N_4698,N_4647);
or U4752 (N_4752,N_4659,N_4674);
and U4753 (N_4753,N_4675,N_4665);
or U4754 (N_4754,N_4622,N_4631);
xnor U4755 (N_4755,N_4671,N_4689);
nor U4756 (N_4756,N_4669,N_4691);
nand U4757 (N_4757,N_4603,N_4656);
nor U4758 (N_4758,N_4696,N_4681);
and U4759 (N_4759,N_4658,N_4669);
nor U4760 (N_4760,N_4638,N_4662);
nand U4761 (N_4761,N_4635,N_4615);
xnor U4762 (N_4762,N_4634,N_4683);
nand U4763 (N_4763,N_4669,N_4629);
nand U4764 (N_4764,N_4667,N_4631);
nor U4765 (N_4765,N_4666,N_4604);
and U4766 (N_4766,N_4635,N_4672);
and U4767 (N_4767,N_4681,N_4640);
xor U4768 (N_4768,N_4696,N_4692);
or U4769 (N_4769,N_4658,N_4639);
xor U4770 (N_4770,N_4621,N_4678);
xor U4771 (N_4771,N_4686,N_4663);
xor U4772 (N_4772,N_4668,N_4623);
nor U4773 (N_4773,N_4660,N_4699);
or U4774 (N_4774,N_4669,N_4676);
nor U4775 (N_4775,N_4600,N_4641);
xnor U4776 (N_4776,N_4638,N_4686);
xor U4777 (N_4777,N_4692,N_4680);
xor U4778 (N_4778,N_4679,N_4696);
or U4779 (N_4779,N_4680,N_4631);
or U4780 (N_4780,N_4694,N_4689);
or U4781 (N_4781,N_4627,N_4623);
or U4782 (N_4782,N_4645,N_4630);
nand U4783 (N_4783,N_4697,N_4696);
nor U4784 (N_4784,N_4676,N_4610);
nor U4785 (N_4785,N_4608,N_4696);
nand U4786 (N_4786,N_4683,N_4652);
and U4787 (N_4787,N_4677,N_4638);
and U4788 (N_4788,N_4631,N_4690);
nand U4789 (N_4789,N_4674,N_4645);
nor U4790 (N_4790,N_4683,N_4664);
or U4791 (N_4791,N_4646,N_4644);
nor U4792 (N_4792,N_4689,N_4605);
nor U4793 (N_4793,N_4611,N_4674);
xor U4794 (N_4794,N_4630,N_4655);
nand U4795 (N_4795,N_4625,N_4623);
or U4796 (N_4796,N_4627,N_4666);
or U4797 (N_4797,N_4610,N_4604);
nor U4798 (N_4798,N_4641,N_4674);
nand U4799 (N_4799,N_4626,N_4690);
or U4800 (N_4800,N_4765,N_4724);
nand U4801 (N_4801,N_4796,N_4755);
nor U4802 (N_4802,N_4710,N_4759);
xnor U4803 (N_4803,N_4795,N_4794);
xnor U4804 (N_4804,N_4718,N_4706);
or U4805 (N_4805,N_4732,N_4771);
nor U4806 (N_4806,N_4752,N_4712);
nand U4807 (N_4807,N_4701,N_4729);
xnor U4808 (N_4808,N_4749,N_4700);
and U4809 (N_4809,N_4761,N_4757);
or U4810 (N_4810,N_4722,N_4780);
nand U4811 (N_4811,N_4743,N_4721);
xor U4812 (N_4812,N_4747,N_4717);
xor U4813 (N_4813,N_4719,N_4772);
nor U4814 (N_4814,N_4769,N_4753);
xor U4815 (N_4815,N_4770,N_4704);
nor U4816 (N_4816,N_4709,N_4754);
nor U4817 (N_4817,N_4737,N_4787);
and U4818 (N_4818,N_4702,N_4748);
and U4819 (N_4819,N_4707,N_4725);
or U4820 (N_4820,N_4745,N_4708);
or U4821 (N_4821,N_4756,N_4733);
and U4822 (N_4822,N_4791,N_4720);
nand U4823 (N_4823,N_4740,N_4742);
nand U4824 (N_4824,N_4763,N_4741);
nand U4825 (N_4825,N_4797,N_4764);
and U4826 (N_4826,N_4731,N_4714);
xnor U4827 (N_4827,N_4775,N_4773);
xnor U4828 (N_4828,N_4776,N_4766);
or U4829 (N_4829,N_4777,N_4751);
xor U4830 (N_4830,N_4738,N_4768);
nand U4831 (N_4831,N_4792,N_4788);
nor U4832 (N_4832,N_4779,N_4723);
and U4833 (N_4833,N_4790,N_4716);
nor U4834 (N_4834,N_4782,N_4750);
and U4835 (N_4835,N_4711,N_4767);
and U4836 (N_4836,N_4736,N_4734);
xnor U4837 (N_4837,N_4705,N_4713);
and U4838 (N_4838,N_4735,N_4746);
xnor U4839 (N_4839,N_4727,N_4728);
nand U4840 (N_4840,N_4744,N_4703);
and U4841 (N_4841,N_4715,N_4785);
and U4842 (N_4842,N_4778,N_4783);
xor U4843 (N_4843,N_4730,N_4781);
and U4844 (N_4844,N_4774,N_4798);
nand U4845 (N_4845,N_4760,N_4739);
nand U4846 (N_4846,N_4784,N_4793);
or U4847 (N_4847,N_4789,N_4762);
and U4848 (N_4848,N_4799,N_4726);
nor U4849 (N_4849,N_4758,N_4786);
and U4850 (N_4850,N_4732,N_4777);
or U4851 (N_4851,N_4742,N_4796);
nor U4852 (N_4852,N_4707,N_4791);
xnor U4853 (N_4853,N_4744,N_4751);
nand U4854 (N_4854,N_4777,N_4747);
or U4855 (N_4855,N_4783,N_4776);
xor U4856 (N_4856,N_4737,N_4721);
and U4857 (N_4857,N_4712,N_4709);
xor U4858 (N_4858,N_4782,N_4715);
nor U4859 (N_4859,N_4748,N_4738);
and U4860 (N_4860,N_4722,N_4768);
and U4861 (N_4861,N_4774,N_4710);
and U4862 (N_4862,N_4780,N_4791);
nand U4863 (N_4863,N_4711,N_4739);
and U4864 (N_4864,N_4719,N_4755);
nor U4865 (N_4865,N_4791,N_4752);
nor U4866 (N_4866,N_4730,N_4711);
nand U4867 (N_4867,N_4729,N_4720);
xnor U4868 (N_4868,N_4739,N_4714);
and U4869 (N_4869,N_4742,N_4715);
xnor U4870 (N_4870,N_4703,N_4720);
nand U4871 (N_4871,N_4729,N_4757);
and U4872 (N_4872,N_4757,N_4760);
and U4873 (N_4873,N_4716,N_4711);
nand U4874 (N_4874,N_4748,N_4722);
nand U4875 (N_4875,N_4704,N_4746);
nor U4876 (N_4876,N_4776,N_4758);
or U4877 (N_4877,N_4773,N_4730);
nand U4878 (N_4878,N_4786,N_4727);
and U4879 (N_4879,N_4746,N_4723);
and U4880 (N_4880,N_4738,N_4713);
or U4881 (N_4881,N_4782,N_4738);
xnor U4882 (N_4882,N_4747,N_4793);
or U4883 (N_4883,N_4755,N_4718);
nor U4884 (N_4884,N_4713,N_4736);
or U4885 (N_4885,N_4730,N_4701);
and U4886 (N_4886,N_4758,N_4733);
xor U4887 (N_4887,N_4726,N_4721);
nor U4888 (N_4888,N_4728,N_4778);
xnor U4889 (N_4889,N_4711,N_4765);
and U4890 (N_4890,N_4706,N_4791);
nand U4891 (N_4891,N_4774,N_4700);
or U4892 (N_4892,N_4730,N_4746);
or U4893 (N_4893,N_4771,N_4769);
xnor U4894 (N_4894,N_4710,N_4705);
and U4895 (N_4895,N_4724,N_4759);
xnor U4896 (N_4896,N_4706,N_4738);
and U4897 (N_4897,N_4788,N_4783);
nand U4898 (N_4898,N_4750,N_4798);
nor U4899 (N_4899,N_4725,N_4732);
and U4900 (N_4900,N_4897,N_4861);
xnor U4901 (N_4901,N_4816,N_4873);
nand U4902 (N_4902,N_4869,N_4813);
nand U4903 (N_4903,N_4856,N_4898);
and U4904 (N_4904,N_4818,N_4839);
or U4905 (N_4905,N_4823,N_4831);
and U4906 (N_4906,N_4833,N_4871);
or U4907 (N_4907,N_4815,N_4899);
nand U4908 (N_4908,N_4874,N_4820);
or U4909 (N_4909,N_4838,N_4892);
nor U4910 (N_4910,N_4819,N_4886);
nor U4911 (N_4911,N_4868,N_4835);
and U4912 (N_4912,N_4883,N_4844);
or U4913 (N_4913,N_4875,N_4829);
or U4914 (N_4914,N_4832,N_4889);
and U4915 (N_4915,N_4852,N_4849);
or U4916 (N_4916,N_4811,N_4885);
or U4917 (N_4917,N_4836,N_4864);
nor U4918 (N_4918,N_4850,N_4804);
and U4919 (N_4919,N_4841,N_4806);
xnor U4920 (N_4920,N_4877,N_4876);
xor U4921 (N_4921,N_4888,N_4845);
nor U4922 (N_4922,N_4812,N_4830);
or U4923 (N_4923,N_4867,N_4872);
and U4924 (N_4924,N_4807,N_4808);
nand U4925 (N_4925,N_4847,N_4893);
or U4926 (N_4926,N_4846,N_4870);
or U4927 (N_4927,N_4805,N_4860);
nor U4928 (N_4928,N_4824,N_4810);
nand U4929 (N_4929,N_4859,N_4866);
xor U4930 (N_4930,N_4891,N_4801);
xor U4931 (N_4931,N_4843,N_4837);
nor U4932 (N_4932,N_4825,N_4821);
or U4933 (N_4933,N_4895,N_4822);
nand U4934 (N_4934,N_4809,N_4887);
xnor U4935 (N_4935,N_4840,N_4828);
xor U4936 (N_4936,N_4858,N_4865);
nor U4937 (N_4937,N_4851,N_4855);
nor U4938 (N_4938,N_4882,N_4857);
nand U4939 (N_4939,N_4884,N_4881);
and U4940 (N_4940,N_4800,N_4803);
and U4941 (N_4941,N_4894,N_4826);
nor U4942 (N_4942,N_4862,N_4827);
nand U4943 (N_4943,N_4834,N_4878);
xor U4944 (N_4944,N_4853,N_4880);
and U4945 (N_4945,N_4802,N_4848);
or U4946 (N_4946,N_4817,N_4842);
nor U4947 (N_4947,N_4896,N_4854);
and U4948 (N_4948,N_4879,N_4814);
or U4949 (N_4949,N_4863,N_4890);
nand U4950 (N_4950,N_4858,N_4883);
nand U4951 (N_4951,N_4808,N_4883);
or U4952 (N_4952,N_4869,N_4803);
nor U4953 (N_4953,N_4801,N_4856);
nand U4954 (N_4954,N_4829,N_4878);
and U4955 (N_4955,N_4858,N_4850);
nand U4956 (N_4956,N_4802,N_4827);
nand U4957 (N_4957,N_4810,N_4831);
and U4958 (N_4958,N_4869,N_4879);
nor U4959 (N_4959,N_4814,N_4829);
nor U4960 (N_4960,N_4804,N_4874);
xor U4961 (N_4961,N_4853,N_4893);
or U4962 (N_4962,N_4892,N_4807);
nand U4963 (N_4963,N_4865,N_4807);
nor U4964 (N_4964,N_4885,N_4836);
or U4965 (N_4965,N_4806,N_4885);
or U4966 (N_4966,N_4848,N_4807);
xor U4967 (N_4967,N_4802,N_4821);
nand U4968 (N_4968,N_4824,N_4895);
or U4969 (N_4969,N_4847,N_4850);
or U4970 (N_4970,N_4859,N_4894);
nand U4971 (N_4971,N_4814,N_4802);
xnor U4972 (N_4972,N_4883,N_4887);
nand U4973 (N_4973,N_4874,N_4863);
or U4974 (N_4974,N_4886,N_4810);
and U4975 (N_4975,N_4871,N_4853);
and U4976 (N_4976,N_4820,N_4817);
and U4977 (N_4977,N_4835,N_4871);
or U4978 (N_4978,N_4886,N_4897);
xnor U4979 (N_4979,N_4881,N_4897);
xor U4980 (N_4980,N_4812,N_4851);
nand U4981 (N_4981,N_4829,N_4869);
or U4982 (N_4982,N_4874,N_4851);
nand U4983 (N_4983,N_4894,N_4864);
or U4984 (N_4984,N_4871,N_4847);
and U4985 (N_4985,N_4887,N_4837);
nor U4986 (N_4986,N_4854,N_4820);
and U4987 (N_4987,N_4851,N_4802);
or U4988 (N_4988,N_4846,N_4873);
and U4989 (N_4989,N_4841,N_4888);
and U4990 (N_4990,N_4835,N_4828);
nor U4991 (N_4991,N_4824,N_4817);
xnor U4992 (N_4992,N_4886,N_4811);
xor U4993 (N_4993,N_4868,N_4845);
nand U4994 (N_4994,N_4881,N_4824);
or U4995 (N_4995,N_4828,N_4802);
nor U4996 (N_4996,N_4859,N_4855);
xnor U4997 (N_4997,N_4855,N_4884);
nor U4998 (N_4998,N_4810,N_4874);
or U4999 (N_4999,N_4862,N_4869);
or UO_0 (O_0,N_4999,N_4945);
nand UO_1 (O_1,N_4962,N_4944);
or UO_2 (O_2,N_4994,N_4925);
xor UO_3 (O_3,N_4991,N_4961);
nor UO_4 (O_4,N_4904,N_4918);
and UO_5 (O_5,N_4973,N_4969);
and UO_6 (O_6,N_4958,N_4957);
and UO_7 (O_7,N_4972,N_4976);
nand UO_8 (O_8,N_4966,N_4978);
and UO_9 (O_9,N_4967,N_4953);
or UO_10 (O_10,N_4990,N_4998);
xnor UO_11 (O_11,N_4981,N_4905);
xnor UO_12 (O_12,N_4983,N_4956);
xor UO_13 (O_13,N_4909,N_4993);
nand UO_14 (O_14,N_4921,N_4927);
nor UO_15 (O_15,N_4934,N_4922);
nor UO_16 (O_16,N_4926,N_4954);
and UO_17 (O_17,N_4907,N_4917);
and UO_18 (O_18,N_4968,N_4986);
or UO_19 (O_19,N_4911,N_4938);
or UO_20 (O_20,N_4955,N_4914);
xnor UO_21 (O_21,N_4935,N_4988);
and UO_22 (O_22,N_4908,N_4974);
and UO_23 (O_23,N_4947,N_4941);
nand UO_24 (O_24,N_4901,N_4924);
and UO_25 (O_25,N_4965,N_4971);
or UO_26 (O_26,N_4975,N_4929);
or UO_27 (O_27,N_4939,N_4950);
xor UO_28 (O_28,N_4979,N_4933);
nand UO_29 (O_29,N_4951,N_4946);
nor UO_30 (O_30,N_4902,N_4903);
and UO_31 (O_31,N_4985,N_4940);
xor UO_32 (O_32,N_4970,N_4936);
xnor UO_33 (O_33,N_4930,N_4995);
or UO_34 (O_34,N_4987,N_4984);
xor UO_35 (O_35,N_4977,N_4928);
or UO_36 (O_36,N_4920,N_4982);
nor UO_37 (O_37,N_4959,N_4960);
xnor UO_38 (O_38,N_4964,N_4906);
xnor UO_39 (O_39,N_4943,N_4932);
and UO_40 (O_40,N_4923,N_4937);
or UO_41 (O_41,N_4989,N_4996);
nand UO_42 (O_42,N_4916,N_4919);
and UO_43 (O_43,N_4952,N_4949);
nor UO_44 (O_44,N_4913,N_4900);
nand UO_45 (O_45,N_4910,N_4912);
xnor UO_46 (O_46,N_4992,N_4963);
xnor UO_47 (O_47,N_4948,N_4980);
nand UO_48 (O_48,N_4997,N_4915);
or UO_49 (O_49,N_4931,N_4942);
and UO_50 (O_50,N_4996,N_4921);
nor UO_51 (O_51,N_4987,N_4926);
xor UO_52 (O_52,N_4925,N_4939);
or UO_53 (O_53,N_4957,N_4986);
nor UO_54 (O_54,N_4934,N_4925);
xnor UO_55 (O_55,N_4917,N_4921);
nor UO_56 (O_56,N_4914,N_4962);
nor UO_57 (O_57,N_4978,N_4955);
or UO_58 (O_58,N_4934,N_4966);
nand UO_59 (O_59,N_4937,N_4970);
nor UO_60 (O_60,N_4959,N_4987);
and UO_61 (O_61,N_4971,N_4932);
nor UO_62 (O_62,N_4975,N_4976);
nor UO_63 (O_63,N_4991,N_4927);
nor UO_64 (O_64,N_4982,N_4986);
nand UO_65 (O_65,N_4973,N_4936);
nand UO_66 (O_66,N_4939,N_4905);
nand UO_67 (O_67,N_4906,N_4936);
nand UO_68 (O_68,N_4990,N_4969);
and UO_69 (O_69,N_4979,N_4925);
and UO_70 (O_70,N_4951,N_4995);
and UO_71 (O_71,N_4949,N_4948);
nand UO_72 (O_72,N_4959,N_4934);
nand UO_73 (O_73,N_4986,N_4951);
nor UO_74 (O_74,N_4907,N_4945);
or UO_75 (O_75,N_4922,N_4961);
or UO_76 (O_76,N_4913,N_4966);
nor UO_77 (O_77,N_4919,N_4988);
nor UO_78 (O_78,N_4964,N_4996);
nor UO_79 (O_79,N_4900,N_4902);
xor UO_80 (O_80,N_4959,N_4910);
nor UO_81 (O_81,N_4980,N_4931);
xor UO_82 (O_82,N_4947,N_4970);
and UO_83 (O_83,N_4997,N_4904);
xnor UO_84 (O_84,N_4997,N_4980);
nand UO_85 (O_85,N_4949,N_4995);
xor UO_86 (O_86,N_4912,N_4989);
xor UO_87 (O_87,N_4983,N_4984);
and UO_88 (O_88,N_4992,N_4900);
and UO_89 (O_89,N_4997,N_4918);
xor UO_90 (O_90,N_4946,N_4910);
nor UO_91 (O_91,N_4946,N_4969);
or UO_92 (O_92,N_4903,N_4964);
xnor UO_93 (O_93,N_4934,N_4996);
or UO_94 (O_94,N_4928,N_4971);
nand UO_95 (O_95,N_4977,N_4955);
nor UO_96 (O_96,N_4961,N_4968);
nand UO_97 (O_97,N_4975,N_4980);
nand UO_98 (O_98,N_4996,N_4968);
nor UO_99 (O_99,N_4990,N_4921);
and UO_100 (O_100,N_4937,N_4973);
xnor UO_101 (O_101,N_4916,N_4950);
xor UO_102 (O_102,N_4999,N_4912);
xnor UO_103 (O_103,N_4965,N_4976);
nor UO_104 (O_104,N_4935,N_4973);
nand UO_105 (O_105,N_4919,N_4902);
or UO_106 (O_106,N_4995,N_4954);
or UO_107 (O_107,N_4938,N_4959);
xnor UO_108 (O_108,N_4979,N_4935);
nand UO_109 (O_109,N_4915,N_4952);
nor UO_110 (O_110,N_4977,N_4939);
and UO_111 (O_111,N_4998,N_4996);
and UO_112 (O_112,N_4917,N_4920);
nand UO_113 (O_113,N_4959,N_4962);
or UO_114 (O_114,N_4952,N_4943);
or UO_115 (O_115,N_4936,N_4954);
or UO_116 (O_116,N_4922,N_4900);
nor UO_117 (O_117,N_4959,N_4973);
nand UO_118 (O_118,N_4907,N_4975);
nor UO_119 (O_119,N_4964,N_4917);
xor UO_120 (O_120,N_4910,N_4909);
nand UO_121 (O_121,N_4913,N_4908);
or UO_122 (O_122,N_4980,N_4900);
or UO_123 (O_123,N_4989,N_4923);
and UO_124 (O_124,N_4937,N_4963);
nor UO_125 (O_125,N_4914,N_4998);
xnor UO_126 (O_126,N_4916,N_4952);
nor UO_127 (O_127,N_4940,N_4955);
nor UO_128 (O_128,N_4965,N_4983);
nand UO_129 (O_129,N_4923,N_4966);
nor UO_130 (O_130,N_4949,N_4997);
nor UO_131 (O_131,N_4994,N_4929);
nand UO_132 (O_132,N_4942,N_4932);
xor UO_133 (O_133,N_4972,N_4921);
or UO_134 (O_134,N_4910,N_4999);
nand UO_135 (O_135,N_4914,N_4921);
or UO_136 (O_136,N_4931,N_4977);
and UO_137 (O_137,N_4949,N_4919);
or UO_138 (O_138,N_4968,N_4976);
nand UO_139 (O_139,N_4905,N_4995);
nor UO_140 (O_140,N_4958,N_4948);
nand UO_141 (O_141,N_4997,N_4975);
xor UO_142 (O_142,N_4990,N_4944);
nor UO_143 (O_143,N_4955,N_4949);
nand UO_144 (O_144,N_4991,N_4941);
xor UO_145 (O_145,N_4915,N_4966);
xnor UO_146 (O_146,N_4962,N_4941);
and UO_147 (O_147,N_4987,N_4953);
nor UO_148 (O_148,N_4966,N_4949);
or UO_149 (O_149,N_4928,N_4949);
xor UO_150 (O_150,N_4951,N_4936);
xnor UO_151 (O_151,N_4916,N_4957);
xor UO_152 (O_152,N_4948,N_4965);
nand UO_153 (O_153,N_4987,N_4957);
xnor UO_154 (O_154,N_4963,N_4933);
nand UO_155 (O_155,N_4906,N_4987);
and UO_156 (O_156,N_4902,N_4942);
or UO_157 (O_157,N_4996,N_4957);
xor UO_158 (O_158,N_4936,N_4940);
xnor UO_159 (O_159,N_4947,N_4966);
nor UO_160 (O_160,N_4950,N_4932);
xor UO_161 (O_161,N_4920,N_4953);
nor UO_162 (O_162,N_4918,N_4941);
nand UO_163 (O_163,N_4988,N_4952);
nand UO_164 (O_164,N_4937,N_4914);
xnor UO_165 (O_165,N_4934,N_4951);
and UO_166 (O_166,N_4932,N_4975);
or UO_167 (O_167,N_4965,N_4955);
or UO_168 (O_168,N_4969,N_4965);
nor UO_169 (O_169,N_4950,N_4999);
nand UO_170 (O_170,N_4982,N_4925);
nor UO_171 (O_171,N_4981,N_4994);
xor UO_172 (O_172,N_4946,N_4995);
nand UO_173 (O_173,N_4997,N_4983);
nor UO_174 (O_174,N_4929,N_4923);
nor UO_175 (O_175,N_4908,N_4941);
nand UO_176 (O_176,N_4939,N_4954);
and UO_177 (O_177,N_4927,N_4924);
nor UO_178 (O_178,N_4989,N_4993);
nand UO_179 (O_179,N_4914,N_4999);
or UO_180 (O_180,N_4950,N_4944);
nor UO_181 (O_181,N_4916,N_4995);
nand UO_182 (O_182,N_4976,N_4920);
nor UO_183 (O_183,N_4981,N_4991);
or UO_184 (O_184,N_4970,N_4924);
or UO_185 (O_185,N_4984,N_4985);
xor UO_186 (O_186,N_4939,N_4926);
or UO_187 (O_187,N_4917,N_4991);
xnor UO_188 (O_188,N_4923,N_4998);
and UO_189 (O_189,N_4940,N_4913);
xnor UO_190 (O_190,N_4997,N_4912);
nand UO_191 (O_191,N_4956,N_4966);
xnor UO_192 (O_192,N_4903,N_4924);
nor UO_193 (O_193,N_4986,N_4927);
and UO_194 (O_194,N_4905,N_4912);
nand UO_195 (O_195,N_4943,N_4985);
nor UO_196 (O_196,N_4990,N_4959);
nand UO_197 (O_197,N_4930,N_4937);
xnor UO_198 (O_198,N_4910,N_4972);
and UO_199 (O_199,N_4946,N_4905);
nand UO_200 (O_200,N_4910,N_4983);
nand UO_201 (O_201,N_4924,N_4908);
and UO_202 (O_202,N_4997,N_4922);
nand UO_203 (O_203,N_4918,N_4917);
or UO_204 (O_204,N_4917,N_4956);
xnor UO_205 (O_205,N_4920,N_4916);
and UO_206 (O_206,N_4921,N_4977);
or UO_207 (O_207,N_4971,N_4986);
xnor UO_208 (O_208,N_4914,N_4920);
or UO_209 (O_209,N_4978,N_4976);
nor UO_210 (O_210,N_4902,N_4926);
nor UO_211 (O_211,N_4932,N_4901);
or UO_212 (O_212,N_4984,N_4986);
nand UO_213 (O_213,N_4947,N_4977);
nor UO_214 (O_214,N_4970,N_4952);
and UO_215 (O_215,N_4921,N_4991);
or UO_216 (O_216,N_4967,N_4936);
or UO_217 (O_217,N_4967,N_4941);
nand UO_218 (O_218,N_4905,N_4907);
xor UO_219 (O_219,N_4908,N_4927);
and UO_220 (O_220,N_4905,N_4960);
nand UO_221 (O_221,N_4978,N_4918);
nor UO_222 (O_222,N_4983,N_4940);
xnor UO_223 (O_223,N_4942,N_4978);
xnor UO_224 (O_224,N_4905,N_4947);
or UO_225 (O_225,N_4977,N_4905);
xnor UO_226 (O_226,N_4943,N_4953);
or UO_227 (O_227,N_4906,N_4926);
nor UO_228 (O_228,N_4910,N_4971);
nand UO_229 (O_229,N_4963,N_4945);
or UO_230 (O_230,N_4908,N_4906);
nor UO_231 (O_231,N_4921,N_4976);
and UO_232 (O_232,N_4965,N_4942);
and UO_233 (O_233,N_4927,N_4946);
nand UO_234 (O_234,N_4951,N_4950);
and UO_235 (O_235,N_4924,N_4986);
or UO_236 (O_236,N_4994,N_4931);
nand UO_237 (O_237,N_4972,N_4992);
nor UO_238 (O_238,N_4912,N_4991);
nor UO_239 (O_239,N_4996,N_4972);
nor UO_240 (O_240,N_4952,N_4933);
and UO_241 (O_241,N_4997,N_4954);
nand UO_242 (O_242,N_4915,N_4967);
xor UO_243 (O_243,N_4921,N_4983);
nand UO_244 (O_244,N_4961,N_4965);
and UO_245 (O_245,N_4988,N_4982);
or UO_246 (O_246,N_4970,N_4905);
nand UO_247 (O_247,N_4983,N_4900);
nand UO_248 (O_248,N_4949,N_4960);
xor UO_249 (O_249,N_4948,N_4989);
nand UO_250 (O_250,N_4947,N_4974);
nand UO_251 (O_251,N_4958,N_4970);
and UO_252 (O_252,N_4903,N_4953);
nor UO_253 (O_253,N_4934,N_4958);
or UO_254 (O_254,N_4969,N_4902);
or UO_255 (O_255,N_4905,N_4964);
nand UO_256 (O_256,N_4982,N_4981);
and UO_257 (O_257,N_4936,N_4968);
nor UO_258 (O_258,N_4974,N_4984);
or UO_259 (O_259,N_4925,N_4997);
nand UO_260 (O_260,N_4981,N_4980);
nand UO_261 (O_261,N_4963,N_4971);
or UO_262 (O_262,N_4904,N_4964);
nor UO_263 (O_263,N_4942,N_4994);
or UO_264 (O_264,N_4994,N_4989);
nand UO_265 (O_265,N_4953,N_4934);
and UO_266 (O_266,N_4960,N_4955);
xnor UO_267 (O_267,N_4948,N_4983);
xnor UO_268 (O_268,N_4988,N_4924);
xnor UO_269 (O_269,N_4903,N_4970);
or UO_270 (O_270,N_4916,N_4990);
nand UO_271 (O_271,N_4912,N_4961);
and UO_272 (O_272,N_4991,N_4995);
nand UO_273 (O_273,N_4909,N_4979);
nand UO_274 (O_274,N_4995,N_4955);
nor UO_275 (O_275,N_4985,N_4915);
nand UO_276 (O_276,N_4991,N_4945);
and UO_277 (O_277,N_4968,N_4966);
nor UO_278 (O_278,N_4934,N_4950);
or UO_279 (O_279,N_4990,N_4919);
and UO_280 (O_280,N_4907,N_4959);
xor UO_281 (O_281,N_4903,N_4909);
and UO_282 (O_282,N_4964,N_4947);
nand UO_283 (O_283,N_4920,N_4926);
nor UO_284 (O_284,N_4947,N_4910);
xor UO_285 (O_285,N_4939,N_4969);
and UO_286 (O_286,N_4922,N_4968);
nor UO_287 (O_287,N_4939,N_4963);
and UO_288 (O_288,N_4968,N_4967);
nor UO_289 (O_289,N_4924,N_4904);
nand UO_290 (O_290,N_4920,N_4966);
nor UO_291 (O_291,N_4992,N_4957);
or UO_292 (O_292,N_4999,N_4943);
xor UO_293 (O_293,N_4979,N_4938);
or UO_294 (O_294,N_4904,N_4905);
xnor UO_295 (O_295,N_4977,N_4986);
xnor UO_296 (O_296,N_4946,N_4955);
nand UO_297 (O_297,N_4950,N_4982);
nor UO_298 (O_298,N_4911,N_4902);
or UO_299 (O_299,N_4988,N_4945);
and UO_300 (O_300,N_4964,N_4952);
or UO_301 (O_301,N_4907,N_4908);
nand UO_302 (O_302,N_4979,N_4936);
and UO_303 (O_303,N_4910,N_4965);
and UO_304 (O_304,N_4956,N_4923);
xnor UO_305 (O_305,N_4931,N_4926);
xnor UO_306 (O_306,N_4957,N_4946);
nand UO_307 (O_307,N_4914,N_4918);
xnor UO_308 (O_308,N_4920,N_4948);
xnor UO_309 (O_309,N_4964,N_4968);
nor UO_310 (O_310,N_4905,N_4997);
xnor UO_311 (O_311,N_4931,N_4947);
and UO_312 (O_312,N_4908,N_4912);
nor UO_313 (O_313,N_4963,N_4966);
or UO_314 (O_314,N_4931,N_4940);
nor UO_315 (O_315,N_4929,N_4980);
nor UO_316 (O_316,N_4960,N_4904);
nor UO_317 (O_317,N_4913,N_4964);
nor UO_318 (O_318,N_4962,N_4979);
xnor UO_319 (O_319,N_4924,N_4961);
or UO_320 (O_320,N_4944,N_4903);
or UO_321 (O_321,N_4922,N_4951);
and UO_322 (O_322,N_4910,N_4920);
xnor UO_323 (O_323,N_4919,N_4976);
xor UO_324 (O_324,N_4950,N_4998);
nor UO_325 (O_325,N_4951,N_4930);
nor UO_326 (O_326,N_4977,N_4943);
nand UO_327 (O_327,N_4903,N_4930);
nand UO_328 (O_328,N_4910,N_4930);
nor UO_329 (O_329,N_4939,N_4978);
or UO_330 (O_330,N_4929,N_4932);
xor UO_331 (O_331,N_4974,N_4928);
or UO_332 (O_332,N_4902,N_4972);
and UO_333 (O_333,N_4940,N_4946);
or UO_334 (O_334,N_4901,N_4903);
nor UO_335 (O_335,N_4929,N_4917);
xnor UO_336 (O_336,N_4992,N_4969);
nor UO_337 (O_337,N_4942,N_4993);
nor UO_338 (O_338,N_4927,N_4996);
nor UO_339 (O_339,N_4976,N_4952);
or UO_340 (O_340,N_4956,N_4979);
xnor UO_341 (O_341,N_4921,N_4902);
and UO_342 (O_342,N_4950,N_4993);
nand UO_343 (O_343,N_4951,N_4942);
xor UO_344 (O_344,N_4927,N_4959);
or UO_345 (O_345,N_4915,N_4950);
nor UO_346 (O_346,N_4982,N_4999);
or UO_347 (O_347,N_4934,N_4928);
nand UO_348 (O_348,N_4912,N_4915);
nand UO_349 (O_349,N_4915,N_4916);
nor UO_350 (O_350,N_4939,N_4947);
nor UO_351 (O_351,N_4929,N_4955);
nor UO_352 (O_352,N_4976,N_4944);
or UO_353 (O_353,N_4963,N_4990);
nor UO_354 (O_354,N_4944,N_4924);
or UO_355 (O_355,N_4975,N_4943);
and UO_356 (O_356,N_4924,N_4956);
nand UO_357 (O_357,N_4902,N_4982);
or UO_358 (O_358,N_4950,N_4957);
and UO_359 (O_359,N_4902,N_4975);
and UO_360 (O_360,N_4986,N_4939);
nor UO_361 (O_361,N_4960,N_4909);
nor UO_362 (O_362,N_4916,N_4987);
xor UO_363 (O_363,N_4990,N_4991);
xnor UO_364 (O_364,N_4924,N_4935);
nand UO_365 (O_365,N_4961,N_4946);
nand UO_366 (O_366,N_4949,N_4910);
nand UO_367 (O_367,N_4943,N_4980);
xnor UO_368 (O_368,N_4964,N_4961);
xnor UO_369 (O_369,N_4985,N_4974);
or UO_370 (O_370,N_4940,N_4998);
nand UO_371 (O_371,N_4970,N_4983);
nand UO_372 (O_372,N_4938,N_4995);
nand UO_373 (O_373,N_4922,N_4973);
xnor UO_374 (O_374,N_4948,N_4978);
and UO_375 (O_375,N_4969,N_4949);
nand UO_376 (O_376,N_4907,N_4958);
nor UO_377 (O_377,N_4951,N_4918);
xnor UO_378 (O_378,N_4926,N_4948);
xnor UO_379 (O_379,N_4954,N_4998);
or UO_380 (O_380,N_4981,N_4996);
xnor UO_381 (O_381,N_4996,N_4932);
and UO_382 (O_382,N_4973,N_4912);
nand UO_383 (O_383,N_4923,N_4915);
or UO_384 (O_384,N_4968,N_4990);
and UO_385 (O_385,N_4984,N_4902);
xnor UO_386 (O_386,N_4993,N_4979);
and UO_387 (O_387,N_4907,N_4995);
and UO_388 (O_388,N_4971,N_4940);
nand UO_389 (O_389,N_4941,N_4943);
xor UO_390 (O_390,N_4958,N_4927);
nor UO_391 (O_391,N_4969,N_4982);
nor UO_392 (O_392,N_4922,N_4917);
xor UO_393 (O_393,N_4907,N_4936);
xnor UO_394 (O_394,N_4905,N_4943);
and UO_395 (O_395,N_4942,N_4971);
and UO_396 (O_396,N_4957,N_4945);
nor UO_397 (O_397,N_4952,N_4998);
nand UO_398 (O_398,N_4969,N_4997);
xor UO_399 (O_399,N_4940,N_4908);
or UO_400 (O_400,N_4987,N_4933);
nor UO_401 (O_401,N_4975,N_4905);
xor UO_402 (O_402,N_4911,N_4932);
nor UO_403 (O_403,N_4987,N_4919);
nand UO_404 (O_404,N_4922,N_4972);
xor UO_405 (O_405,N_4965,N_4931);
or UO_406 (O_406,N_4971,N_4920);
nand UO_407 (O_407,N_4982,N_4918);
nand UO_408 (O_408,N_4943,N_4930);
nor UO_409 (O_409,N_4937,N_4913);
nand UO_410 (O_410,N_4996,N_4938);
nand UO_411 (O_411,N_4987,N_4907);
nand UO_412 (O_412,N_4935,N_4911);
or UO_413 (O_413,N_4980,N_4903);
nand UO_414 (O_414,N_4906,N_4927);
or UO_415 (O_415,N_4918,N_4934);
and UO_416 (O_416,N_4913,N_4903);
or UO_417 (O_417,N_4917,N_4969);
nand UO_418 (O_418,N_4926,N_4915);
xnor UO_419 (O_419,N_4904,N_4984);
or UO_420 (O_420,N_4922,N_4946);
and UO_421 (O_421,N_4990,N_4918);
and UO_422 (O_422,N_4930,N_4969);
nand UO_423 (O_423,N_4920,N_4990);
nor UO_424 (O_424,N_4995,N_4964);
nand UO_425 (O_425,N_4953,N_4990);
and UO_426 (O_426,N_4963,N_4973);
and UO_427 (O_427,N_4964,N_4967);
nor UO_428 (O_428,N_4950,N_4969);
nand UO_429 (O_429,N_4994,N_4977);
nor UO_430 (O_430,N_4969,N_4901);
nand UO_431 (O_431,N_4921,N_4904);
xor UO_432 (O_432,N_4973,N_4951);
or UO_433 (O_433,N_4943,N_4993);
nor UO_434 (O_434,N_4958,N_4962);
xor UO_435 (O_435,N_4912,N_4958);
xnor UO_436 (O_436,N_4945,N_4956);
and UO_437 (O_437,N_4934,N_4911);
nand UO_438 (O_438,N_4992,N_4974);
xnor UO_439 (O_439,N_4995,N_4944);
and UO_440 (O_440,N_4934,N_4939);
and UO_441 (O_441,N_4903,N_4957);
or UO_442 (O_442,N_4904,N_4914);
or UO_443 (O_443,N_4938,N_4918);
nor UO_444 (O_444,N_4969,N_4941);
nand UO_445 (O_445,N_4980,N_4950);
or UO_446 (O_446,N_4975,N_4950);
nand UO_447 (O_447,N_4911,N_4987);
xnor UO_448 (O_448,N_4991,N_4950);
or UO_449 (O_449,N_4967,N_4957);
nor UO_450 (O_450,N_4930,N_4977);
nand UO_451 (O_451,N_4959,N_4954);
xnor UO_452 (O_452,N_4982,N_4931);
or UO_453 (O_453,N_4962,N_4904);
nor UO_454 (O_454,N_4912,N_4936);
and UO_455 (O_455,N_4963,N_4948);
or UO_456 (O_456,N_4904,N_4907);
nor UO_457 (O_457,N_4994,N_4980);
nand UO_458 (O_458,N_4960,N_4914);
or UO_459 (O_459,N_4996,N_4997);
and UO_460 (O_460,N_4913,N_4904);
and UO_461 (O_461,N_4901,N_4939);
or UO_462 (O_462,N_4922,N_4908);
nand UO_463 (O_463,N_4908,N_4973);
or UO_464 (O_464,N_4940,N_4917);
or UO_465 (O_465,N_4987,N_4981);
nor UO_466 (O_466,N_4905,N_4945);
nor UO_467 (O_467,N_4978,N_4970);
and UO_468 (O_468,N_4906,N_4970);
nor UO_469 (O_469,N_4965,N_4934);
nor UO_470 (O_470,N_4950,N_4925);
or UO_471 (O_471,N_4926,N_4972);
xnor UO_472 (O_472,N_4975,N_4909);
xor UO_473 (O_473,N_4931,N_4988);
nand UO_474 (O_474,N_4983,N_4943);
and UO_475 (O_475,N_4971,N_4926);
nor UO_476 (O_476,N_4948,N_4913);
or UO_477 (O_477,N_4928,N_4946);
nor UO_478 (O_478,N_4958,N_4903);
xor UO_479 (O_479,N_4908,N_4958);
nor UO_480 (O_480,N_4915,N_4959);
xnor UO_481 (O_481,N_4999,N_4951);
nand UO_482 (O_482,N_4996,N_4990);
nand UO_483 (O_483,N_4967,N_4992);
xor UO_484 (O_484,N_4910,N_4961);
and UO_485 (O_485,N_4956,N_4965);
or UO_486 (O_486,N_4991,N_4908);
and UO_487 (O_487,N_4969,N_4916);
xnor UO_488 (O_488,N_4904,N_4961);
or UO_489 (O_489,N_4916,N_4974);
or UO_490 (O_490,N_4915,N_4905);
or UO_491 (O_491,N_4992,N_4998);
xor UO_492 (O_492,N_4955,N_4968);
and UO_493 (O_493,N_4958,N_4938);
nor UO_494 (O_494,N_4943,N_4992);
xor UO_495 (O_495,N_4950,N_4958);
or UO_496 (O_496,N_4964,N_4912);
nor UO_497 (O_497,N_4928,N_4986);
nor UO_498 (O_498,N_4948,N_4909);
or UO_499 (O_499,N_4944,N_4925);
or UO_500 (O_500,N_4900,N_4999);
and UO_501 (O_501,N_4977,N_4944);
xor UO_502 (O_502,N_4910,N_4956);
nor UO_503 (O_503,N_4904,N_4945);
or UO_504 (O_504,N_4979,N_4900);
or UO_505 (O_505,N_4912,N_4966);
nor UO_506 (O_506,N_4909,N_4921);
and UO_507 (O_507,N_4951,N_4966);
nand UO_508 (O_508,N_4912,N_4987);
or UO_509 (O_509,N_4991,N_4940);
or UO_510 (O_510,N_4974,N_4904);
nand UO_511 (O_511,N_4953,N_4992);
nand UO_512 (O_512,N_4995,N_4959);
nand UO_513 (O_513,N_4916,N_4921);
nor UO_514 (O_514,N_4976,N_4936);
nor UO_515 (O_515,N_4914,N_4971);
nand UO_516 (O_516,N_4993,N_4973);
nand UO_517 (O_517,N_4945,N_4969);
nor UO_518 (O_518,N_4956,N_4905);
nor UO_519 (O_519,N_4950,N_4923);
nand UO_520 (O_520,N_4967,N_4939);
nor UO_521 (O_521,N_4914,N_4978);
nand UO_522 (O_522,N_4914,N_4980);
xor UO_523 (O_523,N_4960,N_4943);
xor UO_524 (O_524,N_4927,N_4915);
or UO_525 (O_525,N_4959,N_4917);
and UO_526 (O_526,N_4951,N_4976);
and UO_527 (O_527,N_4992,N_4924);
nand UO_528 (O_528,N_4997,N_4902);
xnor UO_529 (O_529,N_4958,N_4902);
nor UO_530 (O_530,N_4954,N_4900);
nor UO_531 (O_531,N_4949,N_4920);
or UO_532 (O_532,N_4990,N_4901);
and UO_533 (O_533,N_4923,N_4970);
nor UO_534 (O_534,N_4960,N_4923);
nand UO_535 (O_535,N_4919,N_4937);
or UO_536 (O_536,N_4923,N_4994);
or UO_537 (O_537,N_4907,N_4946);
nor UO_538 (O_538,N_4910,N_4964);
or UO_539 (O_539,N_4996,N_4903);
nand UO_540 (O_540,N_4993,N_4982);
and UO_541 (O_541,N_4967,N_4972);
and UO_542 (O_542,N_4925,N_4986);
nor UO_543 (O_543,N_4934,N_4924);
nor UO_544 (O_544,N_4923,N_4991);
and UO_545 (O_545,N_4968,N_4947);
or UO_546 (O_546,N_4952,N_4931);
or UO_547 (O_547,N_4946,N_4991);
or UO_548 (O_548,N_4916,N_4953);
or UO_549 (O_549,N_4904,N_4926);
nand UO_550 (O_550,N_4978,N_4937);
xnor UO_551 (O_551,N_4909,N_4943);
nand UO_552 (O_552,N_4974,N_4929);
or UO_553 (O_553,N_4929,N_4952);
or UO_554 (O_554,N_4930,N_4914);
nand UO_555 (O_555,N_4995,N_4988);
xor UO_556 (O_556,N_4986,N_4949);
and UO_557 (O_557,N_4990,N_4910);
xnor UO_558 (O_558,N_4931,N_4993);
nor UO_559 (O_559,N_4916,N_4956);
or UO_560 (O_560,N_4995,N_4912);
xor UO_561 (O_561,N_4931,N_4975);
nand UO_562 (O_562,N_4948,N_4925);
nor UO_563 (O_563,N_4940,N_4965);
nor UO_564 (O_564,N_4937,N_4956);
nor UO_565 (O_565,N_4914,N_4941);
nand UO_566 (O_566,N_4998,N_4931);
and UO_567 (O_567,N_4919,N_4913);
nor UO_568 (O_568,N_4951,N_4972);
nor UO_569 (O_569,N_4994,N_4976);
or UO_570 (O_570,N_4963,N_4983);
nand UO_571 (O_571,N_4948,N_4916);
or UO_572 (O_572,N_4979,N_4975);
and UO_573 (O_573,N_4962,N_4942);
or UO_574 (O_574,N_4952,N_4905);
nor UO_575 (O_575,N_4945,N_4921);
nand UO_576 (O_576,N_4955,N_4910);
xor UO_577 (O_577,N_4908,N_4993);
nand UO_578 (O_578,N_4900,N_4950);
nand UO_579 (O_579,N_4923,N_4968);
nand UO_580 (O_580,N_4991,N_4934);
xnor UO_581 (O_581,N_4944,N_4959);
nand UO_582 (O_582,N_4918,N_4905);
nor UO_583 (O_583,N_4902,N_4968);
and UO_584 (O_584,N_4979,N_4914);
nand UO_585 (O_585,N_4923,N_4992);
or UO_586 (O_586,N_4952,N_4986);
nor UO_587 (O_587,N_4986,N_4909);
or UO_588 (O_588,N_4918,N_4940);
and UO_589 (O_589,N_4903,N_4976);
xnor UO_590 (O_590,N_4906,N_4920);
or UO_591 (O_591,N_4968,N_4991);
or UO_592 (O_592,N_4945,N_4976);
nand UO_593 (O_593,N_4979,N_4959);
xor UO_594 (O_594,N_4902,N_4915);
xnor UO_595 (O_595,N_4927,N_4932);
or UO_596 (O_596,N_4918,N_4963);
nand UO_597 (O_597,N_4912,N_4993);
and UO_598 (O_598,N_4925,N_4928);
xnor UO_599 (O_599,N_4944,N_4980);
nand UO_600 (O_600,N_4981,N_4989);
xor UO_601 (O_601,N_4978,N_4900);
and UO_602 (O_602,N_4987,N_4910);
nor UO_603 (O_603,N_4971,N_4912);
xnor UO_604 (O_604,N_4950,N_4931);
nand UO_605 (O_605,N_4968,N_4959);
and UO_606 (O_606,N_4910,N_4904);
nor UO_607 (O_607,N_4939,N_4949);
xnor UO_608 (O_608,N_4946,N_4934);
and UO_609 (O_609,N_4953,N_4983);
or UO_610 (O_610,N_4995,N_4921);
xor UO_611 (O_611,N_4980,N_4922);
nor UO_612 (O_612,N_4979,N_4911);
or UO_613 (O_613,N_4985,N_4957);
or UO_614 (O_614,N_4932,N_4947);
nor UO_615 (O_615,N_4996,N_4942);
nor UO_616 (O_616,N_4977,N_4911);
nand UO_617 (O_617,N_4928,N_4966);
nor UO_618 (O_618,N_4917,N_4958);
nor UO_619 (O_619,N_4931,N_4996);
nor UO_620 (O_620,N_4980,N_4930);
and UO_621 (O_621,N_4940,N_4993);
or UO_622 (O_622,N_4977,N_4981);
and UO_623 (O_623,N_4971,N_4969);
nand UO_624 (O_624,N_4969,N_4991);
and UO_625 (O_625,N_4970,N_4928);
xor UO_626 (O_626,N_4970,N_4911);
or UO_627 (O_627,N_4913,N_4986);
nor UO_628 (O_628,N_4914,N_4996);
or UO_629 (O_629,N_4932,N_4945);
or UO_630 (O_630,N_4995,N_4975);
nor UO_631 (O_631,N_4906,N_4980);
nor UO_632 (O_632,N_4979,N_4985);
or UO_633 (O_633,N_4929,N_4965);
and UO_634 (O_634,N_4960,N_4983);
and UO_635 (O_635,N_4935,N_4927);
nor UO_636 (O_636,N_4960,N_4935);
or UO_637 (O_637,N_4932,N_4969);
or UO_638 (O_638,N_4919,N_4961);
or UO_639 (O_639,N_4948,N_4914);
nor UO_640 (O_640,N_4967,N_4912);
xor UO_641 (O_641,N_4937,N_4910);
nand UO_642 (O_642,N_4920,N_4905);
and UO_643 (O_643,N_4956,N_4975);
nor UO_644 (O_644,N_4902,N_4963);
xnor UO_645 (O_645,N_4955,N_4930);
nor UO_646 (O_646,N_4914,N_4952);
and UO_647 (O_647,N_4998,N_4970);
nor UO_648 (O_648,N_4951,N_4993);
and UO_649 (O_649,N_4980,N_4925);
nand UO_650 (O_650,N_4911,N_4992);
nor UO_651 (O_651,N_4982,N_4961);
nor UO_652 (O_652,N_4989,N_4924);
nand UO_653 (O_653,N_4922,N_4993);
and UO_654 (O_654,N_4941,N_4961);
nor UO_655 (O_655,N_4948,N_4976);
xor UO_656 (O_656,N_4936,N_4950);
or UO_657 (O_657,N_4945,N_4955);
nor UO_658 (O_658,N_4964,N_4939);
and UO_659 (O_659,N_4957,N_4962);
and UO_660 (O_660,N_4976,N_4983);
xnor UO_661 (O_661,N_4967,N_4988);
or UO_662 (O_662,N_4913,N_4954);
and UO_663 (O_663,N_4959,N_4967);
or UO_664 (O_664,N_4934,N_4963);
and UO_665 (O_665,N_4944,N_4902);
xnor UO_666 (O_666,N_4911,N_4904);
or UO_667 (O_667,N_4923,N_4933);
nor UO_668 (O_668,N_4961,N_4934);
nand UO_669 (O_669,N_4932,N_4944);
nand UO_670 (O_670,N_4980,N_4901);
and UO_671 (O_671,N_4969,N_4958);
and UO_672 (O_672,N_4948,N_4904);
xor UO_673 (O_673,N_4909,N_4953);
xor UO_674 (O_674,N_4994,N_4927);
and UO_675 (O_675,N_4901,N_4961);
nor UO_676 (O_676,N_4958,N_4968);
and UO_677 (O_677,N_4930,N_4908);
xnor UO_678 (O_678,N_4935,N_4915);
nand UO_679 (O_679,N_4916,N_4942);
nor UO_680 (O_680,N_4935,N_4989);
nand UO_681 (O_681,N_4953,N_4988);
nand UO_682 (O_682,N_4976,N_4932);
nand UO_683 (O_683,N_4920,N_4924);
xor UO_684 (O_684,N_4936,N_4982);
xnor UO_685 (O_685,N_4981,N_4918);
or UO_686 (O_686,N_4975,N_4953);
xnor UO_687 (O_687,N_4971,N_4984);
and UO_688 (O_688,N_4904,N_4992);
nand UO_689 (O_689,N_4944,N_4989);
nand UO_690 (O_690,N_4948,N_4941);
xnor UO_691 (O_691,N_4965,N_4918);
nand UO_692 (O_692,N_4910,N_4938);
xor UO_693 (O_693,N_4916,N_4923);
xor UO_694 (O_694,N_4977,N_4923);
nand UO_695 (O_695,N_4900,N_4927);
and UO_696 (O_696,N_4900,N_4948);
or UO_697 (O_697,N_4923,N_4997);
nor UO_698 (O_698,N_4963,N_4904);
nor UO_699 (O_699,N_4991,N_4980);
or UO_700 (O_700,N_4933,N_4961);
or UO_701 (O_701,N_4903,N_4931);
nor UO_702 (O_702,N_4963,N_4998);
nor UO_703 (O_703,N_4946,N_4925);
nand UO_704 (O_704,N_4946,N_4915);
xnor UO_705 (O_705,N_4985,N_4960);
nor UO_706 (O_706,N_4901,N_4933);
and UO_707 (O_707,N_4986,N_4999);
or UO_708 (O_708,N_4961,N_4976);
or UO_709 (O_709,N_4971,N_4916);
nor UO_710 (O_710,N_4945,N_4935);
or UO_711 (O_711,N_4913,N_4992);
xor UO_712 (O_712,N_4921,N_4929);
nor UO_713 (O_713,N_4920,N_4944);
nand UO_714 (O_714,N_4902,N_4914);
and UO_715 (O_715,N_4912,N_4930);
nor UO_716 (O_716,N_4921,N_4913);
nor UO_717 (O_717,N_4990,N_4958);
xnor UO_718 (O_718,N_4902,N_4983);
and UO_719 (O_719,N_4974,N_4932);
or UO_720 (O_720,N_4958,N_4982);
and UO_721 (O_721,N_4973,N_4989);
nand UO_722 (O_722,N_4990,N_4966);
xnor UO_723 (O_723,N_4907,N_4913);
and UO_724 (O_724,N_4922,N_4969);
or UO_725 (O_725,N_4925,N_4915);
nand UO_726 (O_726,N_4921,N_4998);
nand UO_727 (O_727,N_4923,N_4984);
nor UO_728 (O_728,N_4915,N_4913);
nor UO_729 (O_729,N_4975,N_4970);
and UO_730 (O_730,N_4914,N_4946);
xor UO_731 (O_731,N_4949,N_4954);
nor UO_732 (O_732,N_4999,N_4916);
nand UO_733 (O_733,N_4974,N_4905);
or UO_734 (O_734,N_4975,N_4966);
xor UO_735 (O_735,N_4976,N_4967);
or UO_736 (O_736,N_4949,N_4946);
and UO_737 (O_737,N_4980,N_4973);
nand UO_738 (O_738,N_4975,N_4919);
nor UO_739 (O_739,N_4988,N_4955);
xnor UO_740 (O_740,N_4978,N_4961);
or UO_741 (O_741,N_4923,N_4925);
xor UO_742 (O_742,N_4991,N_4905);
xor UO_743 (O_743,N_4971,N_4925);
nor UO_744 (O_744,N_4901,N_4965);
and UO_745 (O_745,N_4924,N_4906);
nor UO_746 (O_746,N_4965,N_4967);
or UO_747 (O_747,N_4955,N_4900);
xnor UO_748 (O_748,N_4911,N_4915);
and UO_749 (O_749,N_4949,N_4904);
nor UO_750 (O_750,N_4911,N_4985);
nand UO_751 (O_751,N_4918,N_4919);
nor UO_752 (O_752,N_4932,N_4949);
nor UO_753 (O_753,N_4902,N_4950);
xnor UO_754 (O_754,N_4916,N_4926);
nand UO_755 (O_755,N_4917,N_4979);
xnor UO_756 (O_756,N_4904,N_4993);
nor UO_757 (O_757,N_4944,N_4958);
nand UO_758 (O_758,N_4999,N_4917);
nor UO_759 (O_759,N_4985,N_4962);
or UO_760 (O_760,N_4983,N_4947);
nor UO_761 (O_761,N_4933,N_4950);
nor UO_762 (O_762,N_4931,N_4945);
or UO_763 (O_763,N_4947,N_4961);
xor UO_764 (O_764,N_4912,N_4956);
nor UO_765 (O_765,N_4943,N_4956);
and UO_766 (O_766,N_4921,N_4992);
or UO_767 (O_767,N_4963,N_4915);
xor UO_768 (O_768,N_4902,N_4906);
and UO_769 (O_769,N_4934,N_4949);
nand UO_770 (O_770,N_4931,N_4939);
xnor UO_771 (O_771,N_4974,N_4982);
xor UO_772 (O_772,N_4936,N_4924);
nor UO_773 (O_773,N_4926,N_4984);
or UO_774 (O_774,N_4923,N_4922);
xor UO_775 (O_775,N_4958,N_4942);
and UO_776 (O_776,N_4971,N_4938);
xnor UO_777 (O_777,N_4907,N_4924);
xnor UO_778 (O_778,N_4917,N_4937);
nand UO_779 (O_779,N_4986,N_4920);
and UO_780 (O_780,N_4933,N_4941);
and UO_781 (O_781,N_4904,N_4989);
xor UO_782 (O_782,N_4941,N_4978);
nor UO_783 (O_783,N_4908,N_4919);
nand UO_784 (O_784,N_4962,N_4981);
nor UO_785 (O_785,N_4942,N_4995);
xor UO_786 (O_786,N_4982,N_4985);
xnor UO_787 (O_787,N_4969,N_4942);
or UO_788 (O_788,N_4955,N_4934);
and UO_789 (O_789,N_4961,N_4942);
nand UO_790 (O_790,N_4919,N_4923);
xor UO_791 (O_791,N_4903,N_4984);
nor UO_792 (O_792,N_4984,N_4970);
or UO_793 (O_793,N_4903,N_4949);
or UO_794 (O_794,N_4943,N_4965);
or UO_795 (O_795,N_4948,N_4935);
nor UO_796 (O_796,N_4992,N_4997);
nand UO_797 (O_797,N_4982,N_4971);
nor UO_798 (O_798,N_4967,N_4929);
nand UO_799 (O_799,N_4918,N_4983);
nand UO_800 (O_800,N_4996,N_4982);
nand UO_801 (O_801,N_4962,N_4902);
nor UO_802 (O_802,N_4928,N_4952);
and UO_803 (O_803,N_4996,N_4907);
xor UO_804 (O_804,N_4946,N_4982);
nand UO_805 (O_805,N_4903,N_4905);
or UO_806 (O_806,N_4975,N_4913);
or UO_807 (O_807,N_4989,N_4929);
and UO_808 (O_808,N_4989,N_4985);
and UO_809 (O_809,N_4912,N_4962);
xnor UO_810 (O_810,N_4980,N_4919);
nand UO_811 (O_811,N_4908,N_4984);
xnor UO_812 (O_812,N_4985,N_4932);
nand UO_813 (O_813,N_4950,N_4907);
nand UO_814 (O_814,N_4995,N_4999);
nor UO_815 (O_815,N_4961,N_4936);
or UO_816 (O_816,N_4915,N_4943);
xor UO_817 (O_817,N_4994,N_4998);
nor UO_818 (O_818,N_4980,N_4902);
xnor UO_819 (O_819,N_4931,N_4934);
or UO_820 (O_820,N_4930,N_4944);
nand UO_821 (O_821,N_4963,N_4931);
nor UO_822 (O_822,N_4938,N_4921);
xor UO_823 (O_823,N_4952,N_4999);
nor UO_824 (O_824,N_4975,N_4923);
nor UO_825 (O_825,N_4970,N_4957);
nor UO_826 (O_826,N_4975,N_4963);
and UO_827 (O_827,N_4910,N_4902);
xnor UO_828 (O_828,N_4989,N_4970);
nand UO_829 (O_829,N_4928,N_4933);
or UO_830 (O_830,N_4903,N_4985);
and UO_831 (O_831,N_4902,N_4949);
and UO_832 (O_832,N_4962,N_4946);
and UO_833 (O_833,N_4919,N_4900);
nand UO_834 (O_834,N_4904,N_4951);
nand UO_835 (O_835,N_4955,N_4931);
nor UO_836 (O_836,N_4968,N_4912);
and UO_837 (O_837,N_4952,N_4901);
nand UO_838 (O_838,N_4940,N_4980);
nand UO_839 (O_839,N_4956,N_4990);
and UO_840 (O_840,N_4925,N_4914);
xor UO_841 (O_841,N_4949,N_4967);
and UO_842 (O_842,N_4901,N_4992);
nor UO_843 (O_843,N_4967,N_4938);
nand UO_844 (O_844,N_4901,N_4983);
and UO_845 (O_845,N_4941,N_4929);
or UO_846 (O_846,N_4938,N_4906);
xnor UO_847 (O_847,N_4910,N_4970);
and UO_848 (O_848,N_4933,N_4948);
xor UO_849 (O_849,N_4946,N_4956);
nor UO_850 (O_850,N_4943,N_4957);
xor UO_851 (O_851,N_4905,N_4906);
xnor UO_852 (O_852,N_4933,N_4953);
and UO_853 (O_853,N_4989,N_4910);
and UO_854 (O_854,N_4924,N_4997);
and UO_855 (O_855,N_4962,N_4928);
xor UO_856 (O_856,N_4932,N_4990);
or UO_857 (O_857,N_4983,N_4949);
nand UO_858 (O_858,N_4914,N_4919);
nor UO_859 (O_859,N_4918,N_4945);
or UO_860 (O_860,N_4947,N_4906);
or UO_861 (O_861,N_4907,N_4912);
nand UO_862 (O_862,N_4937,N_4950);
and UO_863 (O_863,N_4906,N_4946);
nor UO_864 (O_864,N_4988,N_4978);
nor UO_865 (O_865,N_4994,N_4946);
xnor UO_866 (O_866,N_4945,N_4910);
nand UO_867 (O_867,N_4924,N_4999);
nor UO_868 (O_868,N_4914,N_4995);
or UO_869 (O_869,N_4915,N_4972);
and UO_870 (O_870,N_4950,N_4924);
or UO_871 (O_871,N_4945,N_4979);
nor UO_872 (O_872,N_4901,N_4900);
nand UO_873 (O_873,N_4984,N_4980);
or UO_874 (O_874,N_4934,N_4942);
or UO_875 (O_875,N_4933,N_4909);
nor UO_876 (O_876,N_4985,N_4944);
nand UO_877 (O_877,N_4954,N_4921);
nand UO_878 (O_878,N_4995,N_4980);
or UO_879 (O_879,N_4904,N_4940);
or UO_880 (O_880,N_4956,N_4935);
and UO_881 (O_881,N_4905,N_4971);
or UO_882 (O_882,N_4999,N_4965);
and UO_883 (O_883,N_4989,N_4916);
nand UO_884 (O_884,N_4913,N_4951);
nand UO_885 (O_885,N_4989,N_4952);
nand UO_886 (O_886,N_4926,N_4942);
xor UO_887 (O_887,N_4920,N_4945);
xnor UO_888 (O_888,N_4978,N_4933);
or UO_889 (O_889,N_4976,N_4923);
and UO_890 (O_890,N_4915,N_4975);
nand UO_891 (O_891,N_4992,N_4905);
xor UO_892 (O_892,N_4947,N_4993);
and UO_893 (O_893,N_4972,N_4945);
xor UO_894 (O_894,N_4946,N_4972);
nor UO_895 (O_895,N_4978,N_4932);
nand UO_896 (O_896,N_4994,N_4951);
nor UO_897 (O_897,N_4994,N_4973);
nand UO_898 (O_898,N_4998,N_4988);
nand UO_899 (O_899,N_4951,N_4900);
nand UO_900 (O_900,N_4991,N_4948);
nand UO_901 (O_901,N_4936,N_4932);
nor UO_902 (O_902,N_4974,N_4938);
xor UO_903 (O_903,N_4989,N_4945);
or UO_904 (O_904,N_4969,N_4994);
nor UO_905 (O_905,N_4930,N_4962);
xnor UO_906 (O_906,N_4953,N_4938);
nand UO_907 (O_907,N_4931,N_4958);
nand UO_908 (O_908,N_4980,N_4927);
and UO_909 (O_909,N_4910,N_4944);
and UO_910 (O_910,N_4925,N_4940);
nor UO_911 (O_911,N_4918,N_4947);
nor UO_912 (O_912,N_4926,N_4933);
nor UO_913 (O_913,N_4959,N_4992);
nand UO_914 (O_914,N_4928,N_4956);
and UO_915 (O_915,N_4930,N_4939);
or UO_916 (O_916,N_4978,N_4910);
nor UO_917 (O_917,N_4948,N_4903);
nor UO_918 (O_918,N_4905,N_4934);
nand UO_919 (O_919,N_4913,N_4970);
or UO_920 (O_920,N_4986,N_4933);
nor UO_921 (O_921,N_4908,N_4935);
nor UO_922 (O_922,N_4943,N_4913);
nor UO_923 (O_923,N_4934,N_4999);
nor UO_924 (O_924,N_4921,N_4942);
nor UO_925 (O_925,N_4900,N_4925);
nor UO_926 (O_926,N_4956,N_4921);
nor UO_927 (O_927,N_4929,N_4984);
and UO_928 (O_928,N_4998,N_4925);
nand UO_929 (O_929,N_4957,N_4921);
nor UO_930 (O_930,N_4992,N_4909);
nor UO_931 (O_931,N_4942,N_4966);
or UO_932 (O_932,N_4925,N_4936);
nand UO_933 (O_933,N_4911,N_4947);
nor UO_934 (O_934,N_4985,N_4945);
nand UO_935 (O_935,N_4960,N_4915);
nand UO_936 (O_936,N_4945,N_4950);
nand UO_937 (O_937,N_4969,N_4903);
or UO_938 (O_938,N_4983,N_4922);
and UO_939 (O_939,N_4931,N_4904);
nand UO_940 (O_940,N_4979,N_4992);
or UO_941 (O_941,N_4987,N_4952);
and UO_942 (O_942,N_4954,N_4947);
nor UO_943 (O_943,N_4969,N_4928);
or UO_944 (O_944,N_4924,N_4949);
nand UO_945 (O_945,N_4919,N_4929);
and UO_946 (O_946,N_4954,N_4951);
and UO_947 (O_947,N_4981,N_4920);
xnor UO_948 (O_948,N_4931,N_4984);
xor UO_949 (O_949,N_4925,N_4905);
or UO_950 (O_950,N_4901,N_4942);
nor UO_951 (O_951,N_4935,N_4950);
nand UO_952 (O_952,N_4975,N_4920);
and UO_953 (O_953,N_4999,N_4976);
nor UO_954 (O_954,N_4907,N_4994);
or UO_955 (O_955,N_4930,N_4932);
and UO_956 (O_956,N_4942,N_4922);
nand UO_957 (O_957,N_4956,N_4944);
or UO_958 (O_958,N_4943,N_4925);
or UO_959 (O_959,N_4900,N_4936);
nor UO_960 (O_960,N_4923,N_4965);
nor UO_961 (O_961,N_4978,N_4959);
nand UO_962 (O_962,N_4909,N_4998);
xnor UO_963 (O_963,N_4931,N_4979);
xor UO_964 (O_964,N_4902,N_4930);
or UO_965 (O_965,N_4948,N_4919);
nand UO_966 (O_966,N_4991,N_4983);
and UO_967 (O_967,N_4955,N_4950);
or UO_968 (O_968,N_4904,N_4975);
xor UO_969 (O_969,N_4984,N_4988);
or UO_970 (O_970,N_4965,N_4914);
xor UO_971 (O_971,N_4939,N_4975);
nand UO_972 (O_972,N_4967,N_4920);
nor UO_973 (O_973,N_4903,N_4919);
nand UO_974 (O_974,N_4999,N_4969);
xor UO_975 (O_975,N_4987,N_4968);
nor UO_976 (O_976,N_4919,N_4984);
nor UO_977 (O_977,N_4980,N_4961);
nor UO_978 (O_978,N_4900,N_4976);
or UO_979 (O_979,N_4908,N_4904);
or UO_980 (O_980,N_4939,N_4929);
or UO_981 (O_981,N_4925,N_4902);
nor UO_982 (O_982,N_4940,N_4982);
nand UO_983 (O_983,N_4971,N_4993);
nand UO_984 (O_984,N_4914,N_4975);
and UO_985 (O_985,N_4914,N_4988);
nand UO_986 (O_986,N_4963,N_4970);
nand UO_987 (O_987,N_4986,N_4970);
or UO_988 (O_988,N_4962,N_4975);
nor UO_989 (O_989,N_4915,N_4920);
nor UO_990 (O_990,N_4927,N_4972);
nor UO_991 (O_991,N_4990,N_4922);
nor UO_992 (O_992,N_4992,N_4995);
xnor UO_993 (O_993,N_4942,N_4941);
nand UO_994 (O_994,N_4938,N_4902);
and UO_995 (O_995,N_4952,N_4957);
and UO_996 (O_996,N_4942,N_4935);
xnor UO_997 (O_997,N_4955,N_4959);
or UO_998 (O_998,N_4958,N_4910);
or UO_999 (O_999,N_4923,N_4902);
endmodule