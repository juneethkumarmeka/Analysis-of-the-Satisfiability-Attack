module basic_1000_10000_1500_4_levels_2xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
and U0 (N_0,In_428,In_547);
and U1 (N_1,In_85,In_631);
or U2 (N_2,In_921,In_431);
nor U3 (N_3,In_460,In_79);
or U4 (N_4,In_105,In_379);
and U5 (N_5,In_31,In_71);
nor U6 (N_6,In_552,In_92);
and U7 (N_7,In_99,In_157);
and U8 (N_8,In_228,In_935);
or U9 (N_9,In_665,In_809);
or U10 (N_10,In_793,In_322);
or U11 (N_11,In_898,In_108);
nor U12 (N_12,In_590,In_207);
or U13 (N_13,In_347,In_404);
nand U14 (N_14,In_393,In_224);
nor U15 (N_15,In_610,In_883);
or U16 (N_16,In_421,In_253);
and U17 (N_17,In_786,In_450);
or U18 (N_18,In_54,In_971);
and U19 (N_19,In_83,In_959);
nor U20 (N_20,In_981,In_977);
nand U21 (N_21,In_62,In_113);
and U22 (N_22,In_842,In_748);
nor U23 (N_23,In_938,In_510);
or U24 (N_24,In_504,In_409);
nand U25 (N_25,In_463,In_373);
nor U26 (N_26,In_558,In_693);
nor U27 (N_27,In_260,In_823);
nor U28 (N_28,In_104,In_465);
nand U29 (N_29,In_616,In_335);
nand U30 (N_30,In_964,In_109);
nor U31 (N_31,In_613,In_803);
and U32 (N_32,In_1,In_565);
or U33 (N_33,In_423,In_426);
or U34 (N_34,In_61,In_515);
nor U35 (N_35,In_129,In_226);
nand U36 (N_36,In_199,In_97);
nand U37 (N_37,In_672,In_682);
and U38 (N_38,In_169,In_917);
nand U39 (N_39,In_433,In_554);
or U40 (N_40,In_294,In_663);
and U41 (N_41,In_182,In_572);
nor U42 (N_42,In_239,In_644);
nor U43 (N_43,In_652,In_768);
nand U44 (N_44,In_332,In_960);
or U45 (N_45,In_988,In_100);
nand U46 (N_46,In_592,In_601);
nor U47 (N_47,In_167,In_117);
nor U48 (N_48,In_930,In_91);
nand U49 (N_49,In_598,In_309);
and U50 (N_50,In_843,In_493);
nor U51 (N_51,In_544,In_600);
and U52 (N_52,In_406,In_405);
nand U53 (N_53,In_384,In_185);
and U54 (N_54,In_424,In_51);
or U55 (N_55,In_700,In_87);
or U56 (N_56,In_95,In_524);
nor U57 (N_57,In_623,In_779);
or U58 (N_58,In_760,In_640);
or U59 (N_59,In_408,In_999);
or U60 (N_60,In_850,In_762);
and U61 (N_61,In_688,In_902);
or U62 (N_62,In_788,In_120);
or U63 (N_63,In_470,In_881);
and U64 (N_64,In_103,In_683);
and U65 (N_65,In_48,In_269);
xor U66 (N_66,In_86,In_634);
and U67 (N_67,In_675,In_249);
and U68 (N_68,In_98,In_969);
or U69 (N_69,In_326,In_794);
and U70 (N_70,In_934,In_65);
nor U71 (N_71,In_284,In_516);
nand U72 (N_72,In_940,In_501);
and U73 (N_73,In_948,In_630);
and U74 (N_74,In_18,In_336);
or U75 (N_75,In_666,In_102);
or U76 (N_76,In_627,In_751);
or U77 (N_77,In_606,In_929);
and U78 (N_78,In_17,In_522);
xor U79 (N_79,In_179,In_24);
nand U80 (N_80,In_770,In_952);
or U81 (N_81,In_134,In_804);
nand U82 (N_82,In_885,In_538);
or U83 (N_83,In_435,In_746);
nand U84 (N_84,In_314,In_456);
and U85 (N_85,In_965,In_7);
xor U86 (N_86,In_202,In_247);
nand U87 (N_87,In_986,In_142);
and U88 (N_88,In_532,In_642);
and U89 (N_89,In_25,In_670);
and U90 (N_90,In_840,In_234);
and U91 (N_91,In_81,In_101);
nor U92 (N_92,In_434,In_28);
or U93 (N_93,In_39,In_615);
nand U94 (N_94,In_646,In_268);
nand U95 (N_95,In_353,In_714);
nand U96 (N_96,In_947,In_481);
nand U97 (N_97,In_798,In_726);
and U98 (N_98,In_55,In_681);
nand U99 (N_99,In_724,In_928);
or U100 (N_100,In_829,In_818);
and U101 (N_101,In_484,In_933);
or U102 (N_102,In_359,In_776);
nand U103 (N_103,In_469,In_351);
xnor U104 (N_104,In_953,In_696);
nand U105 (N_105,In_784,In_584);
and U106 (N_106,In_360,In_651);
nor U107 (N_107,In_356,In_411);
nor U108 (N_108,In_853,In_432);
nor U109 (N_109,In_58,In_846);
nor U110 (N_110,In_227,In_647);
nand U111 (N_111,In_140,In_759);
nand U112 (N_112,In_989,In_240);
or U113 (N_113,In_719,In_82);
and U114 (N_114,In_325,In_168);
nand U115 (N_115,In_483,In_250);
or U116 (N_116,In_876,In_317);
nand U117 (N_117,In_46,In_440);
nand U118 (N_118,In_566,In_187);
nor U119 (N_119,In_814,In_706);
or U120 (N_120,In_212,In_523);
and U121 (N_121,In_713,In_67);
and U122 (N_122,In_232,In_63);
and U123 (N_123,In_604,In_855);
nand U124 (N_124,In_507,In_715);
nor U125 (N_125,In_632,In_43);
and U126 (N_126,In_758,In_645);
or U127 (N_127,In_531,In_488);
or U128 (N_128,In_560,In_414);
nand U129 (N_129,In_936,In_744);
nor U130 (N_130,In_128,In_860);
or U131 (N_131,In_884,In_236);
or U132 (N_132,In_267,In_443);
nor U133 (N_133,In_164,In_529);
and U134 (N_134,In_910,In_252);
and U135 (N_135,In_299,In_684);
or U136 (N_136,In_661,In_42);
or U137 (N_137,In_304,In_190);
nand U138 (N_138,In_453,In_607);
nor U139 (N_139,In_455,In_19);
or U140 (N_140,In_973,In_705);
nand U141 (N_141,In_820,In_416);
nor U142 (N_142,In_491,In_594);
nor U143 (N_143,In_887,In_135);
and U144 (N_144,In_278,In_72);
nor U145 (N_145,In_474,In_279);
and U146 (N_146,In_192,In_21);
nor U147 (N_147,In_303,In_703);
nor U148 (N_148,In_919,In_815);
and U149 (N_149,In_992,In_293);
nand U150 (N_150,In_14,In_70);
or U151 (N_151,In_892,In_344);
or U152 (N_152,In_525,In_852);
nand U153 (N_153,In_564,In_781);
nand U154 (N_154,In_849,In_478);
and U155 (N_155,In_127,In_545);
nand U156 (N_156,In_352,In_479);
nand U157 (N_157,In_559,In_16);
or U158 (N_158,In_330,In_75);
nand U159 (N_159,In_217,In_595);
and U160 (N_160,In_60,In_276);
or U161 (N_161,In_444,In_126);
xor U162 (N_162,In_660,In_500);
nand U163 (N_163,In_649,In_984);
and U164 (N_164,In_805,In_797);
and U165 (N_165,In_394,In_94);
nor U166 (N_166,In_707,In_738);
nor U167 (N_167,In_257,In_802);
and U168 (N_168,In_913,In_327);
nor U169 (N_169,In_150,In_578);
nand U170 (N_170,In_861,In_462);
xnor U171 (N_171,In_115,In_368);
and U172 (N_172,In_76,In_301);
nand U173 (N_173,In_783,In_889);
nand U174 (N_174,In_34,In_648);
and U175 (N_175,In_580,In_720);
xor U176 (N_176,In_755,In_637);
and U177 (N_177,In_621,In_445);
and U178 (N_178,In_882,In_878);
nand U179 (N_179,In_297,In_401);
nor U180 (N_180,In_331,In_731);
nor U181 (N_181,In_599,In_376);
or U182 (N_182,In_3,In_341);
and U183 (N_183,In_425,In_5);
nand U184 (N_184,In_619,In_691);
nand U185 (N_185,In_742,In_374);
nor U186 (N_186,In_785,In_446);
or U187 (N_187,In_163,In_614);
nand U188 (N_188,In_717,In_879);
nand U189 (N_189,In_740,In_154);
nor U190 (N_190,In_526,In_896);
and U191 (N_191,In_308,In_982);
nor U192 (N_192,In_305,In_518);
or U193 (N_193,In_396,In_904);
and U194 (N_194,In_337,In_451);
and U195 (N_195,In_570,In_967);
nor U196 (N_196,In_12,In_266);
nor U197 (N_197,In_66,In_877);
or U198 (N_198,In_378,In_10);
and U199 (N_199,In_361,In_605);
nor U200 (N_200,In_817,In_867);
nor U201 (N_201,In_402,In_533);
and U202 (N_202,In_589,In_441);
nand U203 (N_203,In_386,In_514);
nand U204 (N_204,In_442,In_668);
and U205 (N_205,In_124,In_870);
or U206 (N_206,In_50,In_213);
and U207 (N_207,In_395,In_505);
nor U208 (N_208,In_674,In_966);
nand U209 (N_209,In_697,In_836);
or U210 (N_210,In_281,In_641);
nand U211 (N_211,In_362,In_245);
xnor U212 (N_212,In_59,In_517);
nand U213 (N_213,In_657,In_84);
nand U214 (N_214,In_761,In_618);
nor U215 (N_215,In_155,In_941);
or U216 (N_216,In_363,In_40);
and U217 (N_217,In_73,In_871);
or U218 (N_218,In_272,In_698);
or U219 (N_219,In_459,In_868);
and U220 (N_220,In_711,In_689);
or U221 (N_221,In_729,In_958);
or U222 (N_222,In_873,In_521);
and U223 (N_223,In_153,In_949);
or U224 (N_224,In_628,In_208);
or U225 (N_225,In_574,In_901);
nor U226 (N_226,In_174,In_807);
nand U227 (N_227,In_201,In_835);
and U228 (N_228,In_975,In_375);
nor U229 (N_229,In_220,In_172);
and U230 (N_230,In_822,In_310);
nand U231 (N_231,In_264,In_890);
and U232 (N_232,In_482,In_158);
nor U233 (N_233,In_561,In_311);
nor U234 (N_234,In_962,In_171);
nand U235 (N_235,In_716,In_26);
and U236 (N_236,In_677,In_944);
nand U237 (N_237,In_68,In_447);
and U238 (N_238,In_712,In_778);
or U239 (N_239,In_143,In_312);
nand U240 (N_240,In_782,In_149);
and U241 (N_241,In_20,In_333);
and U242 (N_242,In_29,In_241);
and U243 (N_243,In_539,In_27);
nor U244 (N_244,In_195,In_38);
nor U245 (N_245,In_695,In_502);
and U246 (N_246,In_288,In_857);
or U247 (N_247,In_439,In_905);
nor U248 (N_248,In_290,In_49);
or U249 (N_249,In_221,In_256);
or U250 (N_250,In_562,In_957);
nor U251 (N_251,In_418,In_242);
nand U252 (N_252,In_816,In_246);
nand U253 (N_253,In_367,In_197);
nor U254 (N_254,In_943,In_160);
nand U255 (N_255,In_650,In_854);
nand U256 (N_256,In_790,In_702);
xor U257 (N_257,In_968,In_830);
nor U258 (N_258,In_792,In_747);
and U259 (N_259,In_80,In_15);
and U260 (N_260,In_215,In_739);
nor U261 (N_261,In_254,In_987);
nor U262 (N_262,In_448,In_391);
or U263 (N_263,In_321,In_139);
nor U264 (N_264,In_951,In_110);
nor U265 (N_265,In_555,In_692);
and U266 (N_266,In_285,In_495);
or U267 (N_267,In_436,In_398);
nand U268 (N_268,In_579,In_370);
nor U269 (N_269,In_800,In_397);
and U270 (N_270,In_122,In_856);
nand U271 (N_271,In_924,In_834);
or U272 (N_272,In_263,In_315);
nand U273 (N_273,In_289,In_399);
nand U274 (N_274,In_571,In_382);
nor U275 (N_275,In_146,In_654);
nor U276 (N_276,In_230,In_513);
nand U277 (N_277,In_419,In_136);
or U278 (N_278,In_8,In_490);
or U279 (N_279,In_198,In_736);
or U280 (N_280,In_653,In_780);
nand U281 (N_281,In_313,In_458);
nor U282 (N_282,In_292,In_93);
and U283 (N_283,In_184,In_506);
or U284 (N_284,In_546,In_235);
xor U285 (N_285,In_990,In_673);
nor U286 (N_286,In_983,In_400);
nand U287 (N_287,In_243,In_549);
nand U288 (N_288,In_833,In_258);
or U289 (N_289,In_123,In_955);
nor U290 (N_290,In_111,In_819);
or U291 (N_291,In_911,In_851);
or U292 (N_292,In_78,In_231);
or U293 (N_293,In_978,In_357);
nand U294 (N_294,In_914,In_69);
nand U295 (N_295,In_22,In_218);
or U296 (N_296,In_183,In_348);
or U297 (N_297,In_669,In_638);
and U298 (N_298,In_723,In_186);
or U299 (N_299,In_56,In_548);
nor U300 (N_300,In_946,In_214);
nand U301 (N_301,In_550,In_741);
or U302 (N_302,In_690,In_725);
or U303 (N_303,In_274,In_461);
or U304 (N_304,In_537,In_286);
nor U305 (N_305,In_365,In_925);
and U306 (N_306,In_827,In_567);
or U307 (N_307,In_372,In_903);
or U308 (N_308,In_90,In_541);
and U309 (N_309,In_534,In_512);
and U310 (N_310,In_118,In_656);
nor U311 (N_311,In_388,In_542);
or U312 (N_312,In_635,In_175);
nor U313 (N_313,In_497,In_177);
nor U314 (N_314,In_324,In_710);
nor U315 (N_315,In_757,In_956);
nand U316 (N_316,In_141,In_338);
or U317 (N_317,In_316,In_480);
or U318 (N_318,In_845,In_2);
or U319 (N_319,In_342,In_583);
and U320 (N_320,In_789,In_858);
nor U321 (N_321,In_166,In_872);
or U322 (N_322,In_528,In_639);
and U323 (N_323,In_733,In_473);
nand U324 (N_324,In_407,In_808);
xor U325 (N_325,In_277,In_282);
nor U326 (N_326,In_131,In_275);
or U327 (N_327,In_976,In_492);
nor U328 (N_328,In_233,In_223);
or U329 (N_329,In_909,In_107);
or U330 (N_330,In_721,In_162);
or U331 (N_331,In_125,In_622);
and U332 (N_332,In_64,In_991);
nor U333 (N_333,In_467,In_886);
or U334 (N_334,In_159,In_307);
and U335 (N_335,In_866,In_509);
and U336 (N_336,In_520,In_6);
and U337 (N_337,In_908,In_568);
nor U338 (N_338,In_259,In_553);
nor U339 (N_339,In_148,In_170);
and U340 (N_340,In_385,In_403);
and U341 (N_341,In_676,In_323);
or U342 (N_342,In_718,In_477);
and U343 (N_343,In_161,In_210);
and U344 (N_344,In_728,In_828);
nand U345 (N_345,In_659,In_611);
or U346 (N_346,In_380,In_735);
nor U347 (N_347,In_620,In_392);
or U348 (N_348,In_180,In_602);
nand U349 (N_349,In_291,In_466);
nand U350 (N_350,In_994,In_273);
and U351 (N_351,In_189,In_457);
xor U352 (N_352,In_270,In_265);
or U353 (N_353,In_918,In_454);
and U354 (N_354,In_147,In_563);
and U355 (N_355,In_114,In_888);
and U356 (N_356,In_222,In_205);
nand U357 (N_357,In_764,In_387);
nor U358 (N_358,In_897,In_121);
or U359 (N_359,In_152,In_848);
nor U360 (N_360,In_907,In_503);
nand U361 (N_361,In_826,In_138);
and U362 (N_362,In_900,In_334);
or U363 (N_363,In_53,In_306);
and U364 (N_364,In_899,In_191);
and U365 (N_365,In_597,In_699);
or U366 (N_366,In_350,In_519);
nand U367 (N_367,In_194,In_730);
or U368 (N_368,In_841,In_181);
nor U369 (N_369,In_612,In_633);
nand U370 (N_370,In_35,In_775);
or U371 (N_371,In_727,In_824);
or U372 (N_372,In_687,In_979);
or U373 (N_373,In_427,In_543);
xor U374 (N_374,In_496,In_133);
nand U375 (N_375,In_116,In_475);
or U376 (N_376,In_251,In_664);
nand U377 (N_377,In_880,In_329);
nand U378 (N_378,In_844,In_722);
nand U379 (N_379,In_796,In_617);
or U380 (N_380,In_864,In_769);
or U381 (N_381,In_643,In_280);
nor U382 (N_382,In_132,In_203);
nand U383 (N_383,In_464,In_993);
or U384 (N_384,In_874,In_678);
and U385 (N_385,In_176,In_756);
and U386 (N_386,In_57,In_821);
and U387 (N_387,In_963,In_206);
nor U388 (N_388,In_23,In_112);
and U389 (N_389,In_799,In_995);
nand U390 (N_390,In_449,In_211);
or U391 (N_391,In_271,In_832);
and U392 (N_392,In_998,In_489);
and U393 (N_393,In_296,In_787);
nor U394 (N_394,In_145,In_45);
nand U395 (N_395,In_972,In_662);
xor U396 (N_396,In_486,In_767);
nand U397 (N_397,In_931,In_345);
and U398 (N_398,In_863,In_319);
or U399 (N_399,In_298,In_302);
nor U400 (N_400,In_499,In_577);
nor U401 (N_401,In_950,In_320);
or U402 (N_402,In_283,In_551);
and U403 (N_403,In_766,In_9);
nand U404 (N_404,In_295,In_916);
nand U405 (N_405,In_923,In_765);
nand U406 (N_406,In_358,In_763);
or U407 (N_407,In_355,In_685);
nand U408 (N_408,In_130,In_997);
nand U409 (N_409,In_178,In_996);
nand U410 (N_410,In_261,In_680);
nand U411 (N_411,In_922,In_985);
xnor U412 (N_412,In_527,In_77);
nand U413 (N_413,In_608,In_945);
and U414 (N_414,In_390,In_237);
nor U415 (N_415,In_188,In_36);
nor U416 (N_416,In_626,In_737);
or U417 (N_417,In_701,In_593);
nand U418 (N_418,In_749,In_586);
xor U419 (N_419,In_318,In_813);
nor U420 (N_420,In_937,In_915);
and U421 (N_421,In_225,In_591);
nor U422 (N_422,In_413,In_216);
and U423 (N_423,In_0,In_151);
nand U424 (N_424,In_912,In_340);
nand U425 (N_425,In_472,In_772);
and U426 (N_426,In_920,In_629);
nor U427 (N_427,In_974,In_89);
or U428 (N_428,In_540,In_745);
and U429 (N_429,In_839,In_364);
or U430 (N_430,In_13,In_33);
nand U431 (N_431,In_193,In_354);
nand U432 (N_432,In_865,In_229);
nand U433 (N_433,In_468,In_573);
or U434 (N_434,In_422,In_238);
xor U435 (N_435,In_204,In_437);
and U436 (N_436,In_825,In_575);
or U437 (N_437,In_417,In_895);
nor U438 (N_438,In_576,In_961);
and U439 (N_439,In_452,In_954);
nor U440 (N_440,In_862,In_556);
xor U441 (N_441,In_349,In_754);
and U442 (N_442,In_636,In_377);
nand U443 (N_443,In_927,In_811);
xnor U444 (N_444,In_893,In_812);
nor U445 (N_445,In_511,In_4);
nand U446 (N_446,In_655,In_603);
nor U447 (N_447,In_906,In_859);
or U448 (N_448,In_262,In_389);
nor U449 (N_449,In_743,In_679);
nand U450 (N_450,In_734,In_686);
and U451 (N_451,In_875,In_791);
nand U452 (N_452,In_200,In_588);
nor U453 (N_453,In_535,In_381);
or U454 (N_454,In_536,In_137);
nor U455 (N_455,In_926,In_777);
nor U456 (N_456,In_287,In_106);
or U457 (N_457,In_587,In_165);
xnor U458 (N_458,In_582,In_476);
and U459 (N_459,In_801,In_430);
nor U460 (N_460,In_96,In_810);
and U461 (N_461,In_156,In_383);
nand U462 (N_462,In_52,In_709);
nor U463 (N_463,In_248,In_869);
nand U464 (N_464,In_346,In_410);
or U465 (N_465,In_667,In_485);
or U466 (N_466,In_752,In_694);
and U467 (N_467,In_658,In_771);
nor U468 (N_468,In_32,In_41);
and U469 (N_469,In_847,In_806);
and U470 (N_470,In_569,In_343);
nor U471 (N_471,In_369,In_932);
and U472 (N_472,In_471,In_30);
nand U473 (N_473,In_894,In_173);
nor U474 (N_474,In_508,In_196);
nand U475 (N_475,In_438,In_144);
nor U476 (N_476,In_557,In_339);
and U477 (N_477,In_581,In_750);
nand U478 (N_478,In_609,In_795);
nand U479 (N_479,In_415,In_980);
nor U480 (N_480,In_74,In_119);
and U481 (N_481,In_371,In_596);
nand U482 (N_482,In_420,In_366);
nand U483 (N_483,In_708,In_209);
and U484 (N_484,In_412,In_773);
nor U485 (N_485,In_704,In_837);
nor U486 (N_486,In_47,In_328);
and U487 (N_487,In_11,In_88);
and U488 (N_488,In_244,In_219);
nand U489 (N_489,In_37,In_625);
nand U490 (N_490,In_774,In_891);
and U491 (N_491,In_753,In_624);
or U492 (N_492,In_494,In_831);
nor U493 (N_493,In_300,In_585);
and U494 (N_494,In_942,In_970);
nor U495 (N_495,In_255,In_487);
nor U496 (N_496,In_429,In_530);
nand U497 (N_497,In_671,In_838);
or U498 (N_498,In_44,In_732);
nand U499 (N_499,In_498,In_939);
or U500 (N_500,In_979,In_579);
and U501 (N_501,In_466,In_499);
or U502 (N_502,In_739,In_531);
nor U503 (N_503,In_842,In_521);
or U504 (N_504,In_187,In_542);
nand U505 (N_505,In_518,In_364);
or U506 (N_506,In_173,In_542);
nand U507 (N_507,In_629,In_35);
nand U508 (N_508,In_202,In_851);
and U509 (N_509,In_677,In_441);
nand U510 (N_510,In_797,In_81);
and U511 (N_511,In_827,In_811);
or U512 (N_512,In_136,In_443);
and U513 (N_513,In_894,In_360);
xor U514 (N_514,In_794,In_994);
and U515 (N_515,In_117,In_435);
nor U516 (N_516,In_321,In_447);
and U517 (N_517,In_860,In_193);
and U518 (N_518,In_57,In_589);
nand U519 (N_519,In_275,In_98);
and U520 (N_520,In_698,In_498);
nor U521 (N_521,In_523,In_909);
or U522 (N_522,In_36,In_881);
nor U523 (N_523,In_851,In_362);
nand U524 (N_524,In_888,In_861);
and U525 (N_525,In_541,In_66);
and U526 (N_526,In_861,In_284);
nand U527 (N_527,In_343,In_692);
and U528 (N_528,In_803,In_382);
and U529 (N_529,In_835,In_725);
or U530 (N_530,In_784,In_521);
and U531 (N_531,In_189,In_867);
or U532 (N_532,In_209,In_726);
or U533 (N_533,In_690,In_522);
nand U534 (N_534,In_274,In_315);
nor U535 (N_535,In_623,In_671);
nor U536 (N_536,In_806,In_166);
or U537 (N_537,In_985,In_425);
or U538 (N_538,In_146,In_330);
or U539 (N_539,In_86,In_278);
nand U540 (N_540,In_905,In_482);
and U541 (N_541,In_433,In_961);
and U542 (N_542,In_668,In_722);
or U543 (N_543,In_330,In_166);
nor U544 (N_544,In_765,In_990);
and U545 (N_545,In_41,In_39);
and U546 (N_546,In_889,In_589);
nor U547 (N_547,In_458,In_110);
xor U548 (N_548,In_672,In_60);
nor U549 (N_549,In_632,In_630);
nor U550 (N_550,In_658,In_468);
or U551 (N_551,In_41,In_980);
and U552 (N_552,In_110,In_107);
and U553 (N_553,In_919,In_42);
nor U554 (N_554,In_151,In_817);
nor U555 (N_555,In_873,In_673);
or U556 (N_556,In_331,In_740);
and U557 (N_557,In_490,In_134);
xor U558 (N_558,In_910,In_854);
nand U559 (N_559,In_243,In_166);
nand U560 (N_560,In_366,In_80);
or U561 (N_561,In_646,In_660);
and U562 (N_562,In_685,In_187);
or U563 (N_563,In_64,In_177);
or U564 (N_564,In_571,In_747);
or U565 (N_565,In_339,In_922);
xnor U566 (N_566,In_723,In_714);
and U567 (N_567,In_620,In_193);
nor U568 (N_568,In_766,In_82);
or U569 (N_569,In_47,In_473);
nor U570 (N_570,In_115,In_794);
nand U571 (N_571,In_396,In_353);
nand U572 (N_572,In_328,In_884);
nor U573 (N_573,In_508,In_279);
nand U574 (N_574,In_609,In_180);
and U575 (N_575,In_534,In_842);
nor U576 (N_576,In_55,In_167);
nand U577 (N_577,In_576,In_32);
or U578 (N_578,In_416,In_226);
nor U579 (N_579,In_312,In_289);
nand U580 (N_580,In_441,In_946);
nand U581 (N_581,In_516,In_620);
and U582 (N_582,In_68,In_759);
and U583 (N_583,In_364,In_689);
nand U584 (N_584,In_534,In_60);
xor U585 (N_585,In_25,In_253);
and U586 (N_586,In_262,In_659);
xor U587 (N_587,In_889,In_581);
or U588 (N_588,In_869,In_227);
xor U589 (N_589,In_211,In_483);
or U590 (N_590,In_252,In_877);
and U591 (N_591,In_152,In_409);
nand U592 (N_592,In_269,In_817);
or U593 (N_593,In_38,In_522);
or U594 (N_594,In_517,In_296);
nand U595 (N_595,In_862,In_563);
nand U596 (N_596,In_903,In_400);
nand U597 (N_597,In_772,In_771);
or U598 (N_598,In_500,In_191);
nand U599 (N_599,In_168,In_633);
or U600 (N_600,In_746,In_21);
nand U601 (N_601,In_827,In_277);
nand U602 (N_602,In_820,In_784);
nor U603 (N_603,In_209,In_318);
or U604 (N_604,In_656,In_134);
and U605 (N_605,In_789,In_451);
or U606 (N_606,In_799,In_724);
nor U607 (N_607,In_305,In_785);
nand U608 (N_608,In_314,In_197);
nor U609 (N_609,In_292,In_409);
nand U610 (N_610,In_544,In_330);
nor U611 (N_611,In_368,In_338);
and U612 (N_612,In_480,In_672);
xor U613 (N_613,In_658,In_580);
nor U614 (N_614,In_135,In_514);
or U615 (N_615,In_308,In_382);
or U616 (N_616,In_772,In_141);
nand U617 (N_617,In_793,In_145);
and U618 (N_618,In_0,In_26);
nand U619 (N_619,In_621,In_989);
or U620 (N_620,In_196,In_143);
and U621 (N_621,In_871,In_192);
nand U622 (N_622,In_503,In_110);
and U623 (N_623,In_730,In_388);
and U624 (N_624,In_539,In_383);
and U625 (N_625,In_885,In_137);
nor U626 (N_626,In_519,In_220);
nand U627 (N_627,In_589,In_332);
or U628 (N_628,In_405,In_42);
or U629 (N_629,In_22,In_943);
or U630 (N_630,In_787,In_601);
and U631 (N_631,In_918,In_302);
or U632 (N_632,In_295,In_228);
and U633 (N_633,In_226,In_394);
nor U634 (N_634,In_330,In_260);
or U635 (N_635,In_374,In_735);
nand U636 (N_636,In_432,In_764);
nand U637 (N_637,In_47,In_714);
nand U638 (N_638,In_770,In_139);
or U639 (N_639,In_417,In_479);
nor U640 (N_640,In_34,In_587);
nor U641 (N_641,In_367,In_74);
nor U642 (N_642,In_120,In_411);
nand U643 (N_643,In_246,In_13);
nor U644 (N_644,In_550,In_433);
nor U645 (N_645,In_388,In_512);
nor U646 (N_646,In_929,In_510);
nor U647 (N_647,In_505,In_625);
nand U648 (N_648,In_977,In_914);
or U649 (N_649,In_301,In_826);
and U650 (N_650,In_838,In_63);
or U651 (N_651,In_424,In_829);
nor U652 (N_652,In_772,In_750);
or U653 (N_653,In_202,In_665);
nor U654 (N_654,In_270,In_902);
nand U655 (N_655,In_650,In_531);
nor U656 (N_656,In_222,In_643);
and U657 (N_657,In_387,In_506);
nand U658 (N_658,In_164,In_581);
and U659 (N_659,In_461,In_932);
nand U660 (N_660,In_272,In_686);
xnor U661 (N_661,In_562,In_225);
nor U662 (N_662,In_164,In_437);
or U663 (N_663,In_598,In_503);
or U664 (N_664,In_782,In_294);
nor U665 (N_665,In_193,In_23);
nor U666 (N_666,In_64,In_579);
or U667 (N_667,In_712,In_18);
nand U668 (N_668,In_898,In_899);
nor U669 (N_669,In_829,In_307);
and U670 (N_670,In_340,In_480);
and U671 (N_671,In_998,In_237);
nand U672 (N_672,In_258,In_281);
or U673 (N_673,In_535,In_554);
or U674 (N_674,In_786,In_248);
or U675 (N_675,In_911,In_307);
nor U676 (N_676,In_764,In_398);
nor U677 (N_677,In_789,In_282);
nand U678 (N_678,In_48,In_542);
and U679 (N_679,In_472,In_522);
nand U680 (N_680,In_914,In_855);
nand U681 (N_681,In_772,In_743);
and U682 (N_682,In_637,In_238);
nor U683 (N_683,In_272,In_3);
nor U684 (N_684,In_612,In_571);
nand U685 (N_685,In_974,In_941);
or U686 (N_686,In_92,In_667);
nand U687 (N_687,In_684,In_155);
and U688 (N_688,In_182,In_983);
nand U689 (N_689,In_995,In_440);
or U690 (N_690,In_544,In_725);
nor U691 (N_691,In_788,In_423);
or U692 (N_692,In_194,In_918);
and U693 (N_693,In_273,In_882);
nand U694 (N_694,In_279,In_481);
nor U695 (N_695,In_774,In_945);
and U696 (N_696,In_763,In_898);
and U697 (N_697,In_240,In_275);
and U698 (N_698,In_788,In_703);
or U699 (N_699,In_51,In_905);
xor U700 (N_700,In_45,In_152);
and U701 (N_701,In_170,In_517);
nand U702 (N_702,In_357,In_617);
nand U703 (N_703,In_451,In_460);
nor U704 (N_704,In_201,In_110);
and U705 (N_705,In_240,In_290);
and U706 (N_706,In_525,In_873);
nor U707 (N_707,In_255,In_193);
or U708 (N_708,In_513,In_254);
nor U709 (N_709,In_21,In_245);
and U710 (N_710,In_9,In_316);
nor U711 (N_711,In_829,In_279);
or U712 (N_712,In_74,In_66);
nand U713 (N_713,In_188,In_990);
nor U714 (N_714,In_177,In_284);
nor U715 (N_715,In_80,In_573);
and U716 (N_716,In_764,In_533);
nand U717 (N_717,In_625,In_286);
or U718 (N_718,In_333,In_2);
and U719 (N_719,In_35,In_86);
nor U720 (N_720,In_93,In_323);
or U721 (N_721,In_734,In_861);
and U722 (N_722,In_621,In_150);
or U723 (N_723,In_349,In_294);
and U724 (N_724,In_237,In_987);
or U725 (N_725,In_325,In_99);
and U726 (N_726,In_723,In_866);
or U727 (N_727,In_504,In_157);
and U728 (N_728,In_465,In_780);
and U729 (N_729,In_911,In_37);
and U730 (N_730,In_350,In_966);
xnor U731 (N_731,In_521,In_688);
nand U732 (N_732,In_167,In_506);
or U733 (N_733,In_990,In_352);
or U734 (N_734,In_811,In_775);
xnor U735 (N_735,In_360,In_429);
or U736 (N_736,In_753,In_920);
or U737 (N_737,In_320,In_827);
and U738 (N_738,In_567,In_688);
nor U739 (N_739,In_221,In_261);
nor U740 (N_740,In_968,In_200);
and U741 (N_741,In_242,In_842);
or U742 (N_742,In_749,In_21);
or U743 (N_743,In_285,In_277);
xor U744 (N_744,In_329,In_901);
nand U745 (N_745,In_836,In_81);
and U746 (N_746,In_23,In_669);
and U747 (N_747,In_305,In_559);
or U748 (N_748,In_184,In_259);
nand U749 (N_749,In_458,In_146);
nor U750 (N_750,In_355,In_535);
nand U751 (N_751,In_283,In_317);
nand U752 (N_752,In_880,In_953);
and U753 (N_753,In_30,In_745);
nor U754 (N_754,In_974,In_399);
nor U755 (N_755,In_510,In_755);
nor U756 (N_756,In_478,In_243);
and U757 (N_757,In_856,In_900);
nor U758 (N_758,In_162,In_591);
or U759 (N_759,In_352,In_558);
nor U760 (N_760,In_543,In_659);
nand U761 (N_761,In_994,In_597);
nand U762 (N_762,In_544,In_646);
and U763 (N_763,In_498,In_509);
nand U764 (N_764,In_575,In_387);
nor U765 (N_765,In_97,In_177);
and U766 (N_766,In_928,In_466);
xor U767 (N_767,In_584,In_480);
or U768 (N_768,In_650,In_300);
or U769 (N_769,In_174,In_281);
or U770 (N_770,In_470,In_275);
nand U771 (N_771,In_272,In_171);
xnor U772 (N_772,In_229,In_907);
nor U773 (N_773,In_784,In_905);
nand U774 (N_774,In_109,In_658);
or U775 (N_775,In_609,In_287);
nor U776 (N_776,In_709,In_661);
nand U777 (N_777,In_275,In_899);
nand U778 (N_778,In_670,In_764);
nor U779 (N_779,In_194,In_421);
nor U780 (N_780,In_827,In_553);
or U781 (N_781,In_129,In_131);
nand U782 (N_782,In_53,In_584);
or U783 (N_783,In_624,In_172);
nand U784 (N_784,In_785,In_878);
and U785 (N_785,In_104,In_930);
nor U786 (N_786,In_496,In_978);
and U787 (N_787,In_7,In_729);
and U788 (N_788,In_125,In_83);
and U789 (N_789,In_68,In_484);
or U790 (N_790,In_437,In_433);
or U791 (N_791,In_433,In_696);
and U792 (N_792,In_820,In_487);
and U793 (N_793,In_204,In_308);
and U794 (N_794,In_480,In_110);
or U795 (N_795,In_304,In_260);
and U796 (N_796,In_998,In_880);
nor U797 (N_797,In_929,In_686);
or U798 (N_798,In_160,In_287);
nand U799 (N_799,In_770,In_457);
nand U800 (N_800,In_285,In_484);
or U801 (N_801,In_702,In_487);
nor U802 (N_802,In_630,In_326);
nor U803 (N_803,In_822,In_914);
nand U804 (N_804,In_959,In_259);
nor U805 (N_805,In_520,In_244);
nor U806 (N_806,In_128,In_863);
and U807 (N_807,In_290,In_352);
nor U808 (N_808,In_392,In_337);
nand U809 (N_809,In_855,In_267);
and U810 (N_810,In_518,In_177);
nand U811 (N_811,In_296,In_17);
nor U812 (N_812,In_468,In_559);
or U813 (N_813,In_980,In_198);
or U814 (N_814,In_31,In_630);
and U815 (N_815,In_725,In_194);
nand U816 (N_816,In_426,In_691);
and U817 (N_817,In_592,In_704);
or U818 (N_818,In_596,In_34);
and U819 (N_819,In_530,In_151);
and U820 (N_820,In_313,In_6);
or U821 (N_821,In_188,In_746);
or U822 (N_822,In_13,In_984);
or U823 (N_823,In_900,In_682);
nand U824 (N_824,In_484,In_4);
and U825 (N_825,In_414,In_124);
or U826 (N_826,In_297,In_555);
or U827 (N_827,In_5,In_339);
nand U828 (N_828,In_819,In_927);
or U829 (N_829,In_712,In_786);
nor U830 (N_830,In_835,In_331);
nand U831 (N_831,In_426,In_291);
nand U832 (N_832,In_950,In_612);
nor U833 (N_833,In_809,In_129);
or U834 (N_834,In_518,In_839);
and U835 (N_835,In_2,In_557);
and U836 (N_836,In_215,In_868);
nand U837 (N_837,In_33,In_134);
or U838 (N_838,In_577,In_261);
nand U839 (N_839,In_802,In_278);
nand U840 (N_840,In_665,In_215);
nor U841 (N_841,In_660,In_80);
nand U842 (N_842,In_48,In_431);
nor U843 (N_843,In_866,In_591);
or U844 (N_844,In_485,In_723);
xnor U845 (N_845,In_553,In_20);
nand U846 (N_846,In_209,In_917);
and U847 (N_847,In_327,In_706);
nand U848 (N_848,In_636,In_175);
nand U849 (N_849,In_0,In_76);
or U850 (N_850,In_967,In_174);
xnor U851 (N_851,In_190,In_744);
nand U852 (N_852,In_243,In_182);
and U853 (N_853,In_618,In_645);
nand U854 (N_854,In_377,In_284);
nand U855 (N_855,In_133,In_695);
nand U856 (N_856,In_897,In_550);
and U857 (N_857,In_289,In_515);
and U858 (N_858,In_78,In_492);
nor U859 (N_859,In_124,In_103);
nor U860 (N_860,In_306,In_547);
nor U861 (N_861,In_919,In_429);
or U862 (N_862,In_163,In_63);
and U863 (N_863,In_862,In_90);
nor U864 (N_864,In_223,In_492);
or U865 (N_865,In_617,In_943);
nand U866 (N_866,In_134,In_759);
and U867 (N_867,In_251,In_723);
xor U868 (N_868,In_437,In_840);
nor U869 (N_869,In_616,In_267);
and U870 (N_870,In_136,In_333);
nand U871 (N_871,In_643,In_144);
nand U872 (N_872,In_556,In_413);
xor U873 (N_873,In_472,In_671);
nand U874 (N_874,In_950,In_899);
nand U875 (N_875,In_403,In_212);
nor U876 (N_876,In_494,In_940);
and U877 (N_877,In_673,In_17);
nor U878 (N_878,In_212,In_492);
or U879 (N_879,In_165,In_595);
nor U880 (N_880,In_606,In_88);
nor U881 (N_881,In_338,In_179);
nand U882 (N_882,In_718,In_243);
nand U883 (N_883,In_104,In_530);
or U884 (N_884,In_658,In_788);
and U885 (N_885,In_196,In_426);
nor U886 (N_886,In_521,In_388);
xor U887 (N_887,In_786,In_862);
nor U888 (N_888,In_87,In_688);
or U889 (N_889,In_668,In_243);
nand U890 (N_890,In_890,In_642);
nor U891 (N_891,In_101,In_264);
and U892 (N_892,In_704,In_667);
nor U893 (N_893,In_175,In_649);
nand U894 (N_894,In_648,In_897);
nand U895 (N_895,In_831,In_898);
nor U896 (N_896,In_939,In_429);
and U897 (N_897,In_266,In_122);
and U898 (N_898,In_404,In_249);
nand U899 (N_899,In_488,In_908);
nor U900 (N_900,In_58,In_252);
or U901 (N_901,In_345,In_541);
or U902 (N_902,In_256,In_12);
nand U903 (N_903,In_909,In_898);
nor U904 (N_904,In_270,In_926);
and U905 (N_905,In_856,In_225);
nor U906 (N_906,In_772,In_641);
or U907 (N_907,In_21,In_305);
and U908 (N_908,In_393,In_974);
or U909 (N_909,In_978,In_264);
nand U910 (N_910,In_310,In_762);
nand U911 (N_911,In_202,In_43);
nand U912 (N_912,In_735,In_199);
nor U913 (N_913,In_388,In_938);
nand U914 (N_914,In_114,In_386);
or U915 (N_915,In_718,In_480);
or U916 (N_916,In_809,In_752);
and U917 (N_917,In_330,In_862);
and U918 (N_918,In_997,In_251);
and U919 (N_919,In_981,In_828);
nor U920 (N_920,In_369,In_262);
and U921 (N_921,In_720,In_514);
nor U922 (N_922,In_91,In_470);
nand U923 (N_923,In_160,In_138);
nand U924 (N_924,In_539,In_407);
nand U925 (N_925,In_449,In_509);
and U926 (N_926,In_928,In_334);
and U927 (N_927,In_975,In_33);
nor U928 (N_928,In_447,In_638);
nand U929 (N_929,In_884,In_694);
and U930 (N_930,In_288,In_616);
or U931 (N_931,In_815,In_185);
or U932 (N_932,In_787,In_606);
or U933 (N_933,In_2,In_466);
or U934 (N_934,In_121,In_199);
nor U935 (N_935,In_512,In_958);
nor U936 (N_936,In_724,In_529);
or U937 (N_937,In_795,In_515);
or U938 (N_938,In_685,In_148);
nor U939 (N_939,In_859,In_111);
nor U940 (N_940,In_617,In_240);
or U941 (N_941,In_175,In_145);
or U942 (N_942,In_59,In_744);
and U943 (N_943,In_888,In_77);
nor U944 (N_944,In_954,In_937);
nand U945 (N_945,In_871,In_782);
nor U946 (N_946,In_989,In_726);
or U947 (N_947,In_57,In_960);
nand U948 (N_948,In_331,In_255);
and U949 (N_949,In_109,In_676);
or U950 (N_950,In_691,In_971);
nor U951 (N_951,In_653,In_447);
and U952 (N_952,In_6,In_596);
and U953 (N_953,In_616,In_380);
nor U954 (N_954,In_633,In_602);
or U955 (N_955,In_228,In_34);
nor U956 (N_956,In_791,In_449);
and U957 (N_957,In_842,In_775);
nand U958 (N_958,In_73,In_906);
nand U959 (N_959,In_16,In_547);
and U960 (N_960,In_959,In_930);
and U961 (N_961,In_705,In_330);
nand U962 (N_962,In_472,In_632);
and U963 (N_963,In_590,In_140);
or U964 (N_964,In_391,In_879);
or U965 (N_965,In_234,In_568);
nor U966 (N_966,In_699,In_171);
xnor U967 (N_967,In_453,In_777);
or U968 (N_968,In_33,In_577);
and U969 (N_969,In_268,In_159);
and U970 (N_970,In_131,In_744);
or U971 (N_971,In_229,In_41);
nor U972 (N_972,In_803,In_492);
xnor U973 (N_973,In_22,In_469);
nor U974 (N_974,In_490,In_611);
or U975 (N_975,In_165,In_644);
nand U976 (N_976,In_827,In_380);
xor U977 (N_977,In_817,In_245);
or U978 (N_978,In_664,In_222);
xor U979 (N_979,In_561,In_730);
or U980 (N_980,In_347,In_721);
and U981 (N_981,In_204,In_402);
or U982 (N_982,In_58,In_197);
nand U983 (N_983,In_261,In_511);
xnor U984 (N_984,In_131,In_166);
and U985 (N_985,In_219,In_187);
nor U986 (N_986,In_373,In_68);
or U987 (N_987,In_618,In_530);
nand U988 (N_988,In_979,In_747);
nand U989 (N_989,In_943,In_889);
or U990 (N_990,In_279,In_410);
or U991 (N_991,In_720,In_791);
nand U992 (N_992,In_703,In_660);
or U993 (N_993,In_160,In_563);
or U994 (N_994,In_69,In_357);
nand U995 (N_995,In_166,In_699);
nor U996 (N_996,In_896,In_271);
or U997 (N_997,In_720,In_574);
xor U998 (N_998,In_732,In_144);
or U999 (N_999,In_489,In_555);
xnor U1000 (N_1000,In_110,In_510);
xnor U1001 (N_1001,In_461,In_256);
nand U1002 (N_1002,In_930,In_637);
nor U1003 (N_1003,In_458,In_310);
xor U1004 (N_1004,In_89,In_423);
or U1005 (N_1005,In_597,In_945);
nor U1006 (N_1006,In_839,In_128);
and U1007 (N_1007,In_665,In_424);
nand U1008 (N_1008,In_862,In_720);
and U1009 (N_1009,In_696,In_914);
and U1010 (N_1010,In_547,In_344);
and U1011 (N_1011,In_329,In_241);
nor U1012 (N_1012,In_115,In_516);
nor U1013 (N_1013,In_285,In_553);
xnor U1014 (N_1014,In_749,In_105);
or U1015 (N_1015,In_854,In_200);
nor U1016 (N_1016,In_879,In_191);
nand U1017 (N_1017,In_567,In_12);
or U1018 (N_1018,In_284,In_281);
and U1019 (N_1019,In_822,In_238);
nand U1020 (N_1020,In_412,In_364);
nor U1021 (N_1021,In_188,In_550);
nor U1022 (N_1022,In_439,In_263);
or U1023 (N_1023,In_607,In_568);
and U1024 (N_1024,In_920,In_487);
or U1025 (N_1025,In_403,In_309);
nand U1026 (N_1026,In_574,In_823);
and U1027 (N_1027,In_840,In_87);
or U1028 (N_1028,In_89,In_848);
nand U1029 (N_1029,In_79,In_304);
xnor U1030 (N_1030,In_627,In_278);
or U1031 (N_1031,In_334,In_563);
xnor U1032 (N_1032,In_950,In_369);
nor U1033 (N_1033,In_118,In_497);
or U1034 (N_1034,In_960,In_885);
or U1035 (N_1035,In_368,In_957);
and U1036 (N_1036,In_46,In_479);
nand U1037 (N_1037,In_686,In_318);
and U1038 (N_1038,In_531,In_687);
nand U1039 (N_1039,In_899,In_893);
and U1040 (N_1040,In_621,In_940);
xor U1041 (N_1041,In_599,In_561);
or U1042 (N_1042,In_134,In_629);
nand U1043 (N_1043,In_595,In_716);
xnor U1044 (N_1044,In_835,In_819);
nand U1045 (N_1045,In_832,In_681);
nand U1046 (N_1046,In_677,In_945);
and U1047 (N_1047,In_421,In_883);
and U1048 (N_1048,In_453,In_472);
nor U1049 (N_1049,In_727,In_642);
and U1050 (N_1050,In_960,In_726);
nand U1051 (N_1051,In_476,In_133);
nor U1052 (N_1052,In_409,In_416);
or U1053 (N_1053,In_29,In_538);
nand U1054 (N_1054,In_746,In_264);
and U1055 (N_1055,In_988,In_333);
nand U1056 (N_1056,In_263,In_535);
nor U1057 (N_1057,In_227,In_612);
nand U1058 (N_1058,In_547,In_475);
nand U1059 (N_1059,In_785,In_285);
nand U1060 (N_1060,In_822,In_258);
and U1061 (N_1061,In_843,In_831);
and U1062 (N_1062,In_706,In_452);
and U1063 (N_1063,In_903,In_403);
nand U1064 (N_1064,In_969,In_822);
and U1065 (N_1065,In_681,In_321);
nand U1066 (N_1066,In_176,In_260);
nor U1067 (N_1067,In_781,In_313);
nor U1068 (N_1068,In_369,In_212);
nand U1069 (N_1069,In_699,In_554);
or U1070 (N_1070,In_244,In_924);
or U1071 (N_1071,In_636,In_296);
nor U1072 (N_1072,In_596,In_721);
nor U1073 (N_1073,In_574,In_122);
nand U1074 (N_1074,In_817,In_71);
nor U1075 (N_1075,In_962,In_366);
and U1076 (N_1076,In_663,In_762);
and U1077 (N_1077,In_665,In_329);
nand U1078 (N_1078,In_866,In_469);
nand U1079 (N_1079,In_992,In_623);
and U1080 (N_1080,In_328,In_40);
nand U1081 (N_1081,In_748,In_711);
nand U1082 (N_1082,In_281,In_563);
or U1083 (N_1083,In_436,In_670);
nor U1084 (N_1084,In_467,In_88);
nor U1085 (N_1085,In_776,In_755);
nand U1086 (N_1086,In_522,In_434);
and U1087 (N_1087,In_376,In_53);
xnor U1088 (N_1088,In_303,In_131);
or U1089 (N_1089,In_820,In_121);
nand U1090 (N_1090,In_201,In_192);
or U1091 (N_1091,In_924,In_392);
nor U1092 (N_1092,In_339,In_880);
and U1093 (N_1093,In_15,In_171);
or U1094 (N_1094,In_512,In_909);
and U1095 (N_1095,In_172,In_647);
nor U1096 (N_1096,In_242,In_796);
nand U1097 (N_1097,In_76,In_972);
nor U1098 (N_1098,In_647,In_461);
nand U1099 (N_1099,In_771,In_19);
xor U1100 (N_1100,In_139,In_407);
or U1101 (N_1101,In_829,In_134);
and U1102 (N_1102,In_911,In_584);
or U1103 (N_1103,In_886,In_60);
nand U1104 (N_1104,In_275,In_144);
nor U1105 (N_1105,In_861,In_695);
nand U1106 (N_1106,In_272,In_151);
or U1107 (N_1107,In_999,In_713);
and U1108 (N_1108,In_314,In_123);
nand U1109 (N_1109,In_446,In_175);
nor U1110 (N_1110,In_358,In_473);
and U1111 (N_1111,In_972,In_864);
and U1112 (N_1112,In_455,In_144);
or U1113 (N_1113,In_931,In_493);
nor U1114 (N_1114,In_455,In_573);
nand U1115 (N_1115,In_393,In_798);
nor U1116 (N_1116,In_759,In_711);
or U1117 (N_1117,In_711,In_702);
nor U1118 (N_1118,In_988,In_973);
nand U1119 (N_1119,In_596,In_451);
nand U1120 (N_1120,In_87,In_325);
or U1121 (N_1121,In_645,In_29);
and U1122 (N_1122,In_791,In_910);
or U1123 (N_1123,In_712,In_980);
nor U1124 (N_1124,In_223,In_97);
nor U1125 (N_1125,In_158,In_148);
and U1126 (N_1126,In_673,In_951);
nor U1127 (N_1127,In_67,In_649);
nand U1128 (N_1128,In_13,In_393);
nand U1129 (N_1129,In_870,In_444);
nand U1130 (N_1130,In_390,In_527);
and U1131 (N_1131,In_590,In_107);
nor U1132 (N_1132,In_786,In_553);
xor U1133 (N_1133,In_771,In_466);
and U1134 (N_1134,In_426,In_693);
and U1135 (N_1135,In_843,In_70);
or U1136 (N_1136,In_227,In_289);
or U1137 (N_1137,In_520,In_765);
nor U1138 (N_1138,In_135,In_919);
and U1139 (N_1139,In_624,In_380);
nand U1140 (N_1140,In_481,In_390);
or U1141 (N_1141,In_538,In_194);
nand U1142 (N_1142,In_178,In_918);
or U1143 (N_1143,In_42,In_416);
nor U1144 (N_1144,In_399,In_841);
and U1145 (N_1145,In_535,In_159);
nand U1146 (N_1146,In_664,In_700);
nand U1147 (N_1147,In_596,In_696);
nor U1148 (N_1148,In_279,In_927);
and U1149 (N_1149,In_305,In_784);
or U1150 (N_1150,In_511,In_723);
nor U1151 (N_1151,In_420,In_680);
nor U1152 (N_1152,In_852,In_801);
nor U1153 (N_1153,In_732,In_804);
nand U1154 (N_1154,In_261,In_34);
and U1155 (N_1155,In_893,In_540);
nand U1156 (N_1156,In_432,In_458);
nor U1157 (N_1157,In_975,In_571);
and U1158 (N_1158,In_444,In_858);
and U1159 (N_1159,In_991,In_895);
nand U1160 (N_1160,In_523,In_460);
or U1161 (N_1161,In_1,In_317);
or U1162 (N_1162,In_126,In_250);
nor U1163 (N_1163,In_154,In_209);
or U1164 (N_1164,In_40,In_60);
nor U1165 (N_1165,In_51,In_342);
nor U1166 (N_1166,In_629,In_345);
nand U1167 (N_1167,In_556,In_26);
xnor U1168 (N_1168,In_751,In_807);
nand U1169 (N_1169,In_852,In_991);
and U1170 (N_1170,In_923,In_114);
or U1171 (N_1171,In_579,In_308);
nor U1172 (N_1172,In_228,In_923);
or U1173 (N_1173,In_128,In_724);
nor U1174 (N_1174,In_472,In_12);
nand U1175 (N_1175,In_655,In_66);
and U1176 (N_1176,In_709,In_369);
nand U1177 (N_1177,In_752,In_505);
and U1178 (N_1178,In_974,In_724);
or U1179 (N_1179,In_688,In_255);
nor U1180 (N_1180,In_471,In_777);
or U1181 (N_1181,In_286,In_674);
nand U1182 (N_1182,In_636,In_951);
or U1183 (N_1183,In_686,In_183);
or U1184 (N_1184,In_872,In_505);
nand U1185 (N_1185,In_937,In_73);
nor U1186 (N_1186,In_498,In_849);
or U1187 (N_1187,In_638,In_542);
and U1188 (N_1188,In_476,In_580);
or U1189 (N_1189,In_568,In_434);
or U1190 (N_1190,In_373,In_909);
nor U1191 (N_1191,In_471,In_749);
and U1192 (N_1192,In_316,In_665);
and U1193 (N_1193,In_32,In_214);
or U1194 (N_1194,In_838,In_158);
and U1195 (N_1195,In_780,In_783);
and U1196 (N_1196,In_349,In_869);
or U1197 (N_1197,In_424,In_93);
and U1198 (N_1198,In_834,In_535);
and U1199 (N_1199,In_769,In_85);
nor U1200 (N_1200,In_474,In_735);
nor U1201 (N_1201,In_574,In_851);
nor U1202 (N_1202,In_830,In_484);
and U1203 (N_1203,In_485,In_978);
and U1204 (N_1204,In_961,In_57);
nand U1205 (N_1205,In_369,In_618);
and U1206 (N_1206,In_761,In_513);
and U1207 (N_1207,In_168,In_164);
xor U1208 (N_1208,In_798,In_863);
nand U1209 (N_1209,In_184,In_218);
nand U1210 (N_1210,In_197,In_400);
and U1211 (N_1211,In_465,In_183);
nor U1212 (N_1212,In_941,In_642);
nand U1213 (N_1213,In_294,In_552);
and U1214 (N_1214,In_85,In_706);
or U1215 (N_1215,In_940,In_270);
or U1216 (N_1216,In_335,In_910);
nand U1217 (N_1217,In_518,In_589);
nand U1218 (N_1218,In_0,In_627);
nor U1219 (N_1219,In_76,In_173);
nor U1220 (N_1220,In_710,In_218);
nor U1221 (N_1221,In_19,In_618);
nor U1222 (N_1222,In_402,In_790);
nor U1223 (N_1223,In_66,In_248);
nor U1224 (N_1224,In_81,In_200);
and U1225 (N_1225,In_929,In_186);
nor U1226 (N_1226,In_309,In_234);
nand U1227 (N_1227,In_656,In_755);
nand U1228 (N_1228,In_669,In_379);
nor U1229 (N_1229,In_742,In_154);
or U1230 (N_1230,In_204,In_225);
nand U1231 (N_1231,In_754,In_734);
or U1232 (N_1232,In_868,In_272);
or U1233 (N_1233,In_264,In_474);
and U1234 (N_1234,In_982,In_531);
nand U1235 (N_1235,In_917,In_644);
nor U1236 (N_1236,In_876,In_543);
nor U1237 (N_1237,In_25,In_201);
nand U1238 (N_1238,In_470,In_183);
or U1239 (N_1239,In_997,In_990);
nor U1240 (N_1240,In_22,In_891);
nor U1241 (N_1241,In_752,In_923);
nor U1242 (N_1242,In_83,In_372);
nor U1243 (N_1243,In_787,In_503);
and U1244 (N_1244,In_550,In_72);
nor U1245 (N_1245,In_791,In_123);
nor U1246 (N_1246,In_864,In_179);
or U1247 (N_1247,In_761,In_631);
and U1248 (N_1248,In_199,In_502);
xor U1249 (N_1249,In_410,In_16);
xnor U1250 (N_1250,In_971,In_126);
nor U1251 (N_1251,In_320,In_391);
nor U1252 (N_1252,In_771,In_335);
and U1253 (N_1253,In_535,In_498);
or U1254 (N_1254,In_239,In_309);
nor U1255 (N_1255,In_68,In_376);
or U1256 (N_1256,In_801,In_83);
nor U1257 (N_1257,In_272,In_400);
nand U1258 (N_1258,In_209,In_176);
nand U1259 (N_1259,In_494,In_276);
and U1260 (N_1260,In_717,In_396);
or U1261 (N_1261,In_746,In_793);
nand U1262 (N_1262,In_154,In_217);
or U1263 (N_1263,In_364,In_307);
nand U1264 (N_1264,In_921,In_497);
nor U1265 (N_1265,In_319,In_50);
nand U1266 (N_1266,In_38,In_467);
nor U1267 (N_1267,In_860,In_525);
nor U1268 (N_1268,In_363,In_268);
nand U1269 (N_1269,In_729,In_596);
and U1270 (N_1270,In_171,In_676);
or U1271 (N_1271,In_989,In_541);
nand U1272 (N_1272,In_275,In_496);
nor U1273 (N_1273,In_331,In_744);
and U1274 (N_1274,In_30,In_539);
and U1275 (N_1275,In_997,In_957);
and U1276 (N_1276,In_49,In_193);
and U1277 (N_1277,In_639,In_11);
nor U1278 (N_1278,In_213,In_896);
nor U1279 (N_1279,In_985,In_363);
nor U1280 (N_1280,In_289,In_161);
and U1281 (N_1281,In_976,In_646);
nand U1282 (N_1282,In_256,In_413);
and U1283 (N_1283,In_20,In_794);
nand U1284 (N_1284,In_97,In_13);
or U1285 (N_1285,In_189,In_849);
xor U1286 (N_1286,In_462,In_784);
nand U1287 (N_1287,In_699,In_366);
nand U1288 (N_1288,In_51,In_434);
nand U1289 (N_1289,In_514,In_483);
or U1290 (N_1290,In_983,In_599);
nand U1291 (N_1291,In_389,In_923);
or U1292 (N_1292,In_28,In_564);
nor U1293 (N_1293,In_360,In_17);
and U1294 (N_1294,In_867,In_610);
or U1295 (N_1295,In_387,In_608);
nand U1296 (N_1296,In_565,In_22);
nand U1297 (N_1297,In_644,In_329);
nand U1298 (N_1298,In_614,In_139);
and U1299 (N_1299,In_266,In_995);
and U1300 (N_1300,In_695,In_730);
nand U1301 (N_1301,In_677,In_273);
nand U1302 (N_1302,In_37,In_117);
or U1303 (N_1303,In_822,In_621);
nand U1304 (N_1304,In_414,In_873);
nor U1305 (N_1305,In_826,In_36);
and U1306 (N_1306,In_938,In_519);
nand U1307 (N_1307,In_434,In_310);
nand U1308 (N_1308,In_736,In_523);
or U1309 (N_1309,In_412,In_334);
or U1310 (N_1310,In_89,In_432);
and U1311 (N_1311,In_630,In_751);
nand U1312 (N_1312,In_551,In_353);
xnor U1313 (N_1313,In_882,In_60);
and U1314 (N_1314,In_253,In_17);
nand U1315 (N_1315,In_960,In_194);
and U1316 (N_1316,In_870,In_510);
or U1317 (N_1317,In_368,In_475);
nand U1318 (N_1318,In_310,In_513);
nand U1319 (N_1319,In_98,In_470);
or U1320 (N_1320,In_507,In_587);
nand U1321 (N_1321,In_296,In_654);
nand U1322 (N_1322,In_505,In_271);
nand U1323 (N_1323,In_616,In_512);
nand U1324 (N_1324,In_727,In_226);
or U1325 (N_1325,In_200,In_392);
nor U1326 (N_1326,In_112,In_422);
and U1327 (N_1327,In_704,In_625);
and U1328 (N_1328,In_774,In_918);
or U1329 (N_1329,In_803,In_226);
nand U1330 (N_1330,In_96,In_235);
and U1331 (N_1331,In_992,In_105);
or U1332 (N_1332,In_798,In_114);
nor U1333 (N_1333,In_963,In_47);
nor U1334 (N_1334,In_419,In_492);
xor U1335 (N_1335,In_874,In_468);
nor U1336 (N_1336,In_211,In_747);
nand U1337 (N_1337,In_511,In_664);
and U1338 (N_1338,In_608,In_485);
and U1339 (N_1339,In_614,In_769);
nor U1340 (N_1340,In_787,In_202);
and U1341 (N_1341,In_338,In_538);
or U1342 (N_1342,In_761,In_122);
and U1343 (N_1343,In_970,In_932);
or U1344 (N_1344,In_622,In_670);
nand U1345 (N_1345,In_540,In_8);
or U1346 (N_1346,In_462,In_166);
nand U1347 (N_1347,In_819,In_315);
and U1348 (N_1348,In_612,In_223);
nand U1349 (N_1349,In_766,In_722);
and U1350 (N_1350,In_106,In_998);
and U1351 (N_1351,In_632,In_361);
and U1352 (N_1352,In_797,In_544);
and U1353 (N_1353,In_399,In_692);
and U1354 (N_1354,In_126,In_811);
or U1355 (N_1355,In_779,In_158);
or U1356 (N_1356,In_681,In_805);
xor U1357 (N_1357,In_282,In_452);
and U1358 (N_1358,In_216,In_338);
and U1359 (N_1359,In_815,In_757);
nand U1360 (N_1360,In_339,In_238);
or U1361 (N_1361,In_463,In_335);
and U1362 (N_1362,In_819,In_528);
and U1363 (N_1363,In_306,In_208);
and U1364 (N_1364,In_623,In_646);
or U1365 (N_1365,In_105,In_561);
nand U1366 (N_1366,In_676,In_196);
nand U1367 (N_1367,In_164,In_414);
nand U1368 (N_1368,In_291,In_899);
or U1369 (N_1369,In_35,In_223);
nor U1370 (N_1370,In_492,In_353);
or U1371 (N_1371,In_25,In_409);
nor U1372 (N_1372,In_688,In_15);
nand U1373 (N_1373,In_506,In_491);
or U1374 (N_1374,In_504,In_887);
nand U1375 (N_1375,In_38,In_457);
xnor U1376 (N_1376,In_28,In_98);
nand U1377 (N_1377,In_610,In_928);
nand U1378 (N_1378,In_684,In_63);
nand U1379 (N_1379,In_413,In_682);
nand U1380 (N_1380,In_896,In_385);
and U1381 (N_1381,In_748,In_107);
nand U1382 (N_1382,In_343,In_104);
nor U1383 (N_1383,In_252,In_632);
and U1384 (N_1384,In_501,In_409);
or U1385 (N_1385,In_819,In_884);
nor U1386 (N_1386,In_1,In_404);
nor U1387 (N_1387,In_854,In_864);
nor U1388 (N_1388,In_102,In_250);
or U1389 (N_1389,In_217,In_882);
or U1390 (N_1390,In_818,In_399);
nand U1391 (N_1391,In_318,In_666);
nor U1392 (N_1392,In_489,In_572);
nand U1393 (N_1393,In_222,In_69);
and U1394 (N_1394,In_314,In_235);
or U1395 (N_1395,In_688,In_151);
nor U1396 (N_1396,In_128,In_980);
nand U1397 (N_1397,In_135,In_589);
and U1398 (N_1398,In_590,In_116);
and U1399 (N_1399,In_389,In_631);
nand U1400 (N_1400,In_919,In_669);
nor U1401 (N_1401,In_290,In_384);
or U1402 (N_1402,In_913,In_468);
nor U1403 (N_1403,In_416,In_591);
nand U1404 (N_1404,In_928,In_300);
nand U1405 (N_1405,In_570,In_912);
nor U1406 (N_1406,In_218,In_479);
and U1407 (N_1407,In_446,In_706);
and U1408 (N_1408,In_805,In_854);
and U1409 (N_1409,In_66,In_588);
or U1410 (N_1410,In_890,In_690);
and U1411 (N_1411,In_909,In_968);
or U1412 (N_1412,In_22,In_324);
nand U1413 (N_1413,In_915,In_311);
nand U1414 (N_1414,In_952,In_139);
and U1415 (N_1415,In_466,In_772);
nand U1416 (N_1416,In_198,In_824);
nand U1417 (N_1417,In_489,In_113);
and U1418 (N_1418,In_613,In_953);
or U1419 (N_1419,In_294,In_795);
nor U1420 (N_1420,In_344,In_943);
nor U1421 (N_1421,In_85,In_886);
and U1422 (N_1422,In_348,In_512);
nand U1423 (N_1423,In_843,In_227);
and U1424 (N_1424,In_906,In_278);
and U1425 (N_1425,In_66,In_612);
and U1426 (N_1426,In_972,In_931);
and U1427 (N_1427,In_82,In_691);
nor U1428 (N_1428,In_861,In_646);
or U1429 (N_1429,In_934,In_173);
and U1430 (N_1430,In_509,In_538);
nand U1431 (N_1431,In_639,In_149);
and U1432 (N_1432,In_188,In_398);
nand U1433 (N_1433,In_492,In_883);
and U1434 (N_1434,In_967,In_39);
nand U1435 (N_1435,In_374,In_519);
or U1436 (N_1436,In_350,In_746);
nand U1437 (N_1437,In_246,In_532);
and U1438 (N_1438,In_546,In_169);
or U1439 (N_1439,In_182,In_132);
or U1440 (N_1440,In_648,In_227);
and U1441 (N_1441,In_408,In_391);
and U1442 (N_1442,In_806,In_543);
or U1443 (N_1443,In_3,In_566);
and U1444 (N_1444,In_370,In_871);
xnor U1445 (N_1445,In_997,In_386);
and U1446 (N_1446,In_374,In_942);
nand U1447 (N_1447,In_826,In_354);
nor U1448 (N_1448,In_542,In_988);
nor U1449 (N_1449,In_527,In_257);
and U1450 (N_1450,In_419,In_284);
or U1451 (N_1451,In_296,In_561);
and U1452 (N_1452,In_735,In_583);
nor U1453 (N_1453,In_542,In_444);
nand U1454 (N_1454,In_786,In_649);
nor U1455 (N_1455,In_370,In_836);
and U1456 (N_1456,In_470,In_754);
and U1457 (N_1457,In_344,In_134);
nand U1458 (N_1458,In_36,In_251);
or U1459 (N_1459,In_885,In_378);
nor U1460 (N_1460,In_136,In_341);
or U1461 (N_1461,In_952,In_349);
nor U1462 (N_1462,In_337,In_425);
nand U1463 (N_1463,In_843,In_92);
or U1464 (N_1464,In_376,In_970);
and U1465 (N_1465,In_721,In_414);
nand U1466 (N_1466,In_212,In_990);
or U1467 (N_1467,In_244,In_81);
nand U1468 (N_1468,In_448,In_392);
nand U1469 (N_1469,In_453,In_483);
and U1470 (N_1470,In_945,In_85);
nand U1471 (N_1471,In_333,In_189);
and U1472 (N_1472,In_307,In_683);
or U1473 (N_1473,In_182,In_694);
and U1474 (N_1474,In_286,In_496);
or U1475 (N_1475,In_829,In_174);
nor U1476 (N_1476,In_681,In_364);
or U1477 (N_1477,In_29,In_173);
nand U1478 (N_1478,In_341,In_143);
and U1479 (N_1479,In_630,In_282);
or U1480 (N_1480,In_368,In_566);
and U1481 (N_1481,In_389,In_465);
and U1482 (N_1482,In_738,In_661);
nor U1483 (N_1483,In_226,In_74);
nand U1484 (N_1484,In_716,In_899);
nand U1485 (N_1485,In_109,In_916);
nand U1486 (N_1486,In_819,In_157);
or U1487 (N_1487,In_426,In_344);
and U1488 (N_1488,In_637,In_24);
nand U1489 (N_1489,In_490,In_418);
and U1490 (N_1490,In_351,In_206);
nand U1491 (N_1491,In_576,In_676);
and U1492 (N_1492,In_18,In_256);
or U1493 (N_1493,In_520,In_42);
and U1494 (N_1494,In_489,In_410);
nand U1495 (N_1495,In_38,In_965);
and U1496 (N_1496,In_156,In_912);
or U1497 (N_1497,In_214,In_928);
nand U1498 (N_1498,In_271,In_852);
or U1499 (N_1499,In_223,In_722);
nand U1500 (N_1500,In_612,In_879);
nor U1501 (N_1501,In_547,In_159);
or U1502 (N_1502,In_133,In_234);
nor U1503 (N_1503,In_947,In_151);
nand U1504 (N_1504,In_630,In_695);
or U1505 (N_1505,In_54,In_272);
or U1506 (N_1506,In_795,In_228);
nand U1507 (N_1507,In_610,In_312);
or U1508 (N_1508,In_658,In_948);
nand U1509 (N_1509,In_188,In_769);
and U1510 (N_1510,In_400,In_381);
nand U1511 (N_1511,In_162,In_754);
or U1512 (N_1512,In_830,In_482);
nor U1513 (N_1513,In_549,In_699);
nor U1514 (N_1514,In_681,In_460);
nor U1515 (N_1515,In_908,In_145);
or U1516 (N_1516,In_985,In_386);
or U1517 (N_1517,In_875,In_917);
and U1518 (N_1518,In_726,In_377);
and U1519 (N_1519,In_237,In_260);
nor U1520 (N_1520,In_156,In_836);
nand U1521 (N_1521,In_462,In_790);
nand U1522 (N_1522,In_712,In_831);
or U1523 (N_1523,In_595,In_698);
and U1524 (N_1524,In_988,In_452);
or U1525 (N_1525,In_50,In_269);
nor U1526 (N_1526,In_751,In_46);
or U1527 (N_1527,In_323,In_325);
nor U1528 (N_1528,In_810,In_832);
or U1529 (N_1529,In_971,In_266);
or U1530 (N_1530,In_652,In_482);
nand U1531 (N_1531,In_813,In_448);
nand U1532 (N_1532,In_682,In_437);
and U1533 (N_1533,In_680,In_436);
or U1534 (N_1534,In_531,In_35);
or U1535 (N_1535,In_107,In_131);
or U1536 (N_1536,In_161,In_836);
or U1537 (N_1537,In_427,In_677);
nand U1538 (N_1538,In_638,In_593);
or U1539 (N_1539,In_333,In_230);
nor U1540 (N_1540,In_236,In_274);
nor U1541 (N_1541,In_875,In_148);
and U1542 (N_1542,In_135,In_749);
and U1543 (N_1543,In_607,In_713);
and U1544 (N_1544,In_819,In_765);
nor U1545 (N_1545,In_881,In_337);
nand U1546 (N_1546,In_595,In_418);
and U1547 (N_1547,In_343,In_228);
nor U1548 (N_1548,In_244,In_779);
and U1549 (N_1549,In_93,In_418);
and U1550 (N_1550,In_421,In_396);
and U1551 (N_1551,In_274,In_406);
nor U1552 (N_1552,In_997,In_367);
nor U1553 (N_1553,In_983,In_593);
nor U1554 (N_1554,In_241,In_448);
nor U1555 (N_1555,In_381,In_181);
nand U1556 (N_1556,In_119,In_947);
nor U1557 (N_1557,In_114,In_512);
nor U1558 (N_1558,In_114,In_440);
xor U1559 (N_1559,In_678,In_18);
nand U1560 (N_1560,In_681,In_875);
or U1561 (N_1561,In_744,In_534);
or U1562 (N_1562,In_291,In_514);
or U1563 (N_1563,In_845,In_668);
or U1564 (N_1564,In_898,In_233);
nand U1565 (N_1565,In_402,In_846);
nand U1566 (N_1566,In_45,In_871);
nand U1567 (N_1567,In_21,In_352);
or U1568 (N_1568,In_481,In_813);
nor U1569 (N_1569,In_305,In_190);
nand U1570 (N_1570,In_40,In_512);
nor U1571 (N_1571,In_689,In_185);
nand U1572 (N_1572,In_493,In_115);
nand U1573 (N_1573,In_310,In_719);
or U1574 (N_1574,In_25,In_369);
nor U1575 (N_1575,In_674,In_842);
and U1576 (N_1576,In_190,In_439);
and U1577 (N_1577,In_920,In_260);
or U1578 (N_1578,In_708,In_963);
nand U1579 (N_1579,In_578,In_52);
nor U1580 (N_1580,In_416,In_753);
and U1581 (N_1581,In_539,In_748);
or U1582 (N_1582,In_119,In_888);
and U1583 (N_1583,In_698,In_847);
and U1584 (N_1584,In_174,In_339);
and U1585 (N_1585,In_678,In_883);
and U1586 (N_1586,In_826,In_503);
nor U1587 (N_1587,In_968,In_23);
or U1588 (N_1588,In_647,In_351);
and U1589 (N_1589,In_883,In_752);
nand U1590 (N_1590,In_962,In_705);
or U1591 (N_1591,In_912,In_957);
nand U1592 (N_1592,In_232,In_795);
or U1593 (N_1593,In_902,In_428);
nor U1594 (N_1594,In_196,In_974);
and U1595 (N_1595,In_903,In_92);
or U1596 (N_1596,In_352,In_796);
nand U1597 (N_1597,In_597,In_14);
nand U1598 (N_1598,In_149,In_301);
or U1599 (N_1599,In_207,In_293);
and U1600 (N_1600,In_928,In_818);
and U1601 (N_1601,In_102,In_971);
and U1602 (N_1602,In_664,In_499);
and U1603 (N_1603,In_834,In_769);
and U1604 (N_1604,In_330,In_223);
nand U1605 (N_1605,In_228,In_171);
nand U1606 (N_1606,In_821,In_875);
or U1607 (N_1607,In_539,In_144);
nand U1608 (N_1608,In_792,In_41);
nor U1609 (N_1609,In_762,In_389);
nor U1610 (N_1610,In_281,In_787);
and U1611 (N_1611,In_928,In_620);
nor U1612 (N_1612,In_721,In_51);
xnor U1613 (N_1613,In_168,In_257);
nor U1614 (N_1614,In_237,In_774);
and U1615 (N_1615,In_329,In_163);
and U1616 (N_1616,In_692,In_749);
or U1617 (N_1617,In_666,In_352);
or U1618 (N_1618,In_21,In_644);
nand U1619 (N_1619,In_936,In_211);
and U1620 (N_1620,In_828,In_405);
or U1621 (N_1621,In_975,In_773);
nand U1622 (N_1622,In_691,In_289);
nor U1623 (N_1623,In_80,In_969);
nor U1624 (N_1624,In_473,In_547);
nor U1625 (N_1625,In_248,In_363);
or U1626 (N_1626,In_173,In_924);
nor U1627 (N_1627,In_990,In_110);
nand U1628 (N_1628,In_3,In_643);
and U1629 (N_1629,In_588,In_914);
nor U1630 (N_1630,In_430,In_380);
and U1631 (N_1631,In_215,In_124);
and U1632 (N_1632,In_173,In_417);
nor U1633 (N_1633,In_426,In_965);
xnor U1634 (N_1634,In_918,In_413);
nor U1635 (N_1635,In_410,In_996);
nor U1636 (N_1636,In_423,In_333);
nand U1637 (N_1637,In_134,In_565);
nor U1638 (N_1638,In_417,In_632);
or U1639 (N_1639,In_182,In_865);
and U1640 (N_1640,In_936,In_467);
nor U1641 (N_1641,In_360,In_540);
nor U1642 (N_1642,In_657,In_113);
xnor U1643 (N_1643,In_17,In_367);
or U1644 (N_1644,In_783,In_561);
and U1645 (N_1645,In_541,In_28);
and U1646 (N_1646,In_112,In_884);
or U1647 (N_1647,In_862,In_181);
or U1648 (N_1648,In_163,In_348);
or U1649 (N_1649,In_854,In_580);
or U1650 (N_1650,In_401,In_935);
and U1651 (N_1651,In_453,In_78);
nor U1652 (N_1652,In_989,In_133);
xnor U1653 (N_1653,In_608,In_952);
nor U1654 (N_1654,In_859,In_355);
or U1655 (N_1655,In_551,In_155);
nor U1656 (N_1656,In_719,In_818);
nand U1657 (N_1657,In_43,In_214);
and U1658 (N_1658,In_264,In_108);
nor U1659 (N_1659,In_336,In_206);
nor U1660 (N_1660,In_617,In_119);
nor U1661 (N_1661,In_593,In_935);
and U1662 (N_1662,In_164,In_866);
and U1663 (N_1663,In_85,In_847);
and U1664 (N_1664,In_636,In_680);
nand U1665 (N_1665,In_155,In_277);
nand U1666 (N_1666,In_757,In_184);
nor U1667 (N_1667,In_806,In_867);
and U1668 (N_1668,In_722,In_532);
nor U1669 (N_1669,In_901,In_13);
nor U1670 (N_1670,In_637,In_119);
or U1671 (N_1671,In_526,In_173);
and U1672 (N_1672,In_100,In_379);
nand U1673 (N_1673,In_72,In_157);
or U1674 (N_1674,In_693,In_368);
or U1675 (N_1675,In_483,In_323);
nor U1676 (N_1676,In_77,In_659);
nor U1677 (N_1677,In_239,In_132);
nand U1678 (N_1678,In_587,In_811);
nor U1679 (N_1679,In_112,In_845);
or U1680 (N_1680,In_476,In_629);
nor U1681 (N_1681,In_845,In_367);
nor U1682 (N_1682,In_134,In_352);
and U1683 (N_1683,In_890,In_320);
nor U1684 (N_1684,In_256,In_805);
or U1685 (N_1685,In_126,In_388);
and U1686 (N_1686,In_622,In_843);
nor U1687 (N_1687,In_705,In_577);
xnor U1688 (N_1688,In_915,In_177);
or U1689 (N_1689,In_171,In_651);
and U1690 (N_1690,In_993,In_875);
or U1691 (N_1691,In_805,In_361);
nand U1692 (N_1692,In_111,In_955);
or U1693 (N_1693,In_528,In_689);
nand U1694 (N_1694,In_250,In_267);
and U1695 (N_1695,In_62,In_997);
nand U1696 (N_1696,In_627,In_434);
and U1697 (N_1697,In_399,In_292);
and U1698 (N_1698,In_905,In_461);
nor U1699 (N_1699,In_227,In_935);
or U1700 (N_1700,In_230,In_670);
nand U1701 (N_1701,In_497,In_181);
and U1702 (N_1702,In_123,In_417);
nor U1703 (N_1703,In_298,In_826);
nand U1704 (N_1704,In_766,In_821);
nor U1705 (N_1705,In_224,In_595);
and U1706 (N_1706,In_455,In_51);
or U1707 (N_1707,In_72,In_441);
or U1708 (N_1708,In_836,In_194);
or U1709 (N_1709,In_446,In_159);
and U1710 (N_1710,In_767,In_773);
nand U1711 (N_1711,In_525,In_601);
xnor U1712 (N_1712,In_476,In_490);
nand U1713 (N_1713,In_194,In_668);
or U1714 (N_1714,In_688,In_637);
or U1715 (N_1715,In_737,In_799);
nor U1716 (N_1716,In_409,In_672);
and U1717 (N_1717,In_6,In_307);
or U1718 (N_1718,In_516,In_153);
and U1719 (N_1719,In_827,In_483);
and U1720 (N_1720,In_543,In_852);
nor U1721 (N_1721,In_299,In_559);
or U1722 (N_1722,In_589,In_261);
or U1723 (N_1723,In_586,In_795);
nand U1724 (N_1724,In_508,In_156);
nand U1725 (N_1725,In_830,In_86);
and U1726 (N_1726,In_969,In_338);
nor U1727 (N_1727,In_313,In_428);
nand U1728 (N_1728,In_504,In_758);
nand U1729 (N_1729,In_824,In_934);
xnor U1730 (N_1730,In_486,In_552);
or U1731 (N_1731,In_959,In_186);
or U1732 (N_1732,In_627,In_494);
nand U1733 (N_1733,In_43,In_811);
xnor U1734 (N_1734,In_303,In_355);
or U1735 (N_1735,In_338,In_394);
or U1736 (N_1736,In_317,In_76);
nor U1737 (N_1737,In_137,In_920);
or U1738 (N_1738,In_6,In_813);
and U1739 (N_1739,In_42,In_943);
nand U1740 (N_1740,In_226,In_785);
nor U1741 (N_1741,In_245,In_158);
or U1742 (N_1742,In_670,In_656);
nor U1743 (N_1743,In_339,In_338);
nor U1744 (N_1744,In_444,In_826);
nor U1745 (N_1745,In_793,In_135);
nor U1746 (N_1746,In_562,In_510);
nand U1747 (N_1747,In_991,In_487);
and U1748 (N_1748,In_228,In_726);
xnor U1749 (N_1749,In_35,In_613);
nand U1750 (N_1750,In_617,In_246);
or U1751 (N_1751,In_825,In_460);
nand U1752 (N_1752,In_921,In_551);
and U1753 (N_1753,In_517,In_615);
and U1754 (N_1754,In_93,In_286);
and U1755 (N_1755,In_753,In_226);
or U1756 (N_1756,In_614,In_124);
nand U1757 (N_1757,In_118,In_70);
or U1758 (N_1758,In_408,In_576);
nor U1759 (N_1759,In_667,In_21);
nand U1760 (N_1760,In_351,In_205);
or U1761 (N_1761,In_329,In_139);
and U1762 (N_1762,In_210,In_29);
nand U1763 (N_1763,In_790,In_567);
and U1764 (N_1764,In_122,In_895);
or U1765 (N_1765,In_362,In_738);
xnor U1766 (N_1766,In_826,In_234);
nand U1767 (N_1767,In_551,In_191);
and U1768 (N_1768,In_191,In_347);
and U1769 (N_1769,In_793,In_525);
xor U1770 (N_1770,In_608,In_292);
nand U1771 (N_1771,In_437,In_351);
or U1772 (N_1772,In_111,In_730);
nor U1773 (N_1773,In_30,In_340);
nor U1774 (N_1774,In_333,In_39);
or U1775 (N_1775,In_982,In_970);
or U1776 (N_1776,In_761,In_10);
or U1777 (N_1777,In_719,In_152);
nand U1778 (N_1778,In_646,In_248);
nand U1779 (N_1779,In_715,In_904);
and U1780 (N_1780,In_938,In_515);
and U1781 (N_1781,In_330,In_773);
and U1782 (N_1782,In_575,In_272);
or U1783 (N_1783,In_534,In_295);
nand U1784 (N_1784,In_41,In_830);
nor U1785 (N_1785,In_720,In_42);
nor U1786 (N_1786,In_28,In_611);
or U1787 (N_1787,In_647,In_865);
nand U1788 (N_1788,In_228,In_624);
and U1789 (N_1789,In_302,In_117);
and U1790 (N_1790,In_176,In_326);
or U1791 (N_1791,In_816,In_141);
and U1792 (N_1792,In_291,In_975);
or U1793 (N_1793,In_685,In_268);
nand U1794 (N_1794,In_390,In_588);
nand U1795 (N_1795,In_648,In_559);
and U1796 (N_1796,In_425,In_848);
and U1797 (N_1797,In_433,In_752);
and U1798 (N_1798,In_78,In_423);
or U1799 (N_1799,In_471,In_266);
or U1800 (N_1800,In_562,In_786);
nand U1801 (N_1801,In_640,In_643);
and U1802 (N_1802,In_648,In_797);
nor U1803 (N_1803,In_442,In_838);
and U1804 (N_1804,In_694,In_487);
nor U1805 (N_1805,In_959,In_533);
nor U1806 (N_1806,In_168,In_542);
nand U1807 (N_1807,In_908,In_320);
nand U1808 (N_1808,In_609,In_880);
or U1809 (N_1809,In_761,In_882);
or U1810 (N_1810,In_2,In_660);
nand U1811 (N_1811,In_654,In_669);
or U1812 (N_1812,In_741,In_551);
and U1813 (N_1813,In_882,In_774);
nand U1814 (N_1814,In_467,In_723);
and U1815 (N_1815,In_167,In_758);
or U1816 (N_1816,In_931,In_866);
or U1817 (N_1817,In_529,In_199);
and U1818 (N_1818,In_42,In_141);
or U1819 (N_1819,In_397,In_793);
xor U1820 (N_1820,In_983,In_960);
nor U1821 (N_1821,In_489,In_119);
nand U1822 (N_1822,In_258,In_651);
and U1823 (N_1823,In_361,In_552);
and U1824 (N_1824,In_392,In_358);
nand U1825 (N_1825,In_854,In_529);
nand U1826 (N_1826,In_598,In_824);
and U1827 (N_1827,In_606,In_62);
nand U1828 (N_1828,In_396,In_990);
nand U1829 (N_1829,In_55,In_410);
nor U1830 (N_1830,In_214,In_336);
or U1831 (N_1831,In_726,In_672);
nand U1832 (N_1832,In_831,In_978);
nand U1833 (N_1833,In_900,In_395);
xnor U1834 (N_1834,In_46,In_404);
xnor U1835 (N_1835,In_469,In_132);
nor U1836 (N_1836,In_984,In_995);
and U1837 (N_1837,In_924,In_910);
nand U1838 (N_1838,In_939,In_399);
nor U1839 (N_1839,In_606,In_782);
nor U1840 (N_1840,In_578,In_551);
nand U1841 (N_1841,In_773,In_103);
and U1842 (N_1842,In_795,In_566);
or U1843 (N_1843,In_224,In_402);
nand U1844 (N_1844,In_573,In_200);
nor U1845 (N_1845,In_164,In_338);
nor U1846 (N_1846,In_952,In_647);
nand U1847 (N_1847,In_744,In_946);
nand U1848 (N_1848,In_191,In_650);
nor U1849 (N_1849,In_635,In_836);
nand U1850 (N_1850,In_187,In_291);
nor U1851 (N_1851,In_177,In_522);
nor U1852 (N_1852,In_593,In_585);
nand U1853 (N_1853,In_794,In_236);
or U1854 (N_1854,In_296,In_490);
nand U1855 (N_1855,In_606,In_582);
or U1856 (N_1856,In_595,In_115);
nor U1857 (N_1857,In_216,In_314);
nand U1858 (N_1858,In_57,In_994);
and U1859 (N_1859,In_850,In_147);
nor U1860 (N_1860,In_568,In_356);
or U1861 (N_1861,In_746,In_694);
and U1862 (N_1862,In_353,In_634);
and U1863 (N_1863,In_824,In_470);
or U1864 (N_1864,In_999,In_986);
nand U1865 (N_1865,In_69,In_815);
nand U1866 (N_1866,In_715,In_506);
and U1867 (N_1867,In_659,In_301);
nand U1868 (N_1868,In_529,In_213);
nor U1869 (N_1869,In_937,In_456);
nor U1870 (N_1870,In_797,In_903);
xnor U1871 (N_1871,In_861,In_159);
nand U1872 (N_1872,In_769,In_949);
nand U1873 (N_1873,In_143,In_573);
nor U1874 (N_1874,In_163,In_176);
nand U1875 (N_1875,In_681,In_483);
nor U1876 (N_1876,In_968,In_351);
and U1877 (N_1877,In_118,In_714);
nand U1878 (N_1878,In_243,In_501);
and U1879 (N_1879,In_488,In_78);
or U1880 (N_1880,In_42,In_173);
and U1881 (N_1881,In_399,In_653);
and U1882 (N_1882,In_552,In_478);
or U1883 (N_1883,In_812,In_983);
and U1884 (N_1884,In_486,In_948);
or U1885 (N_1885,In_138,In_422);
or U1886 (N_1886,In_635,In_618);
nand U1887 (N_1887,In_633,In_879);
or U1888 (N_1888,In_635,In_672);
or U1889 (N_1889,In_827,In_960);
nand U1890 (N_1890,In_296,In_789);
and U1891 (N_1891,In_752,In_519);
or U1892 (N_1892,In_357,In_861);
nor U1893 (N_1893,In_59,In_574);
or U1894 (N_1894,In_681,In_997);
nand U1895 (N_1895,In_308,In_21);
nor U1896 (N_1896,In_478,In_22);
and U1897 (N_1897,In_938,In_797);
nand U1898 (N_1898,In_725,In_167);
nand U1899 (N_1899,In_222,In_743);
and U1900 (N_1900,In_671,In_423);
and U1901 (N_1901,In_734,In_432);
or U1902 (N_1902,In_432,In_841);
and U1903 (N_1903,In_42,In_851);
nor U1904 (N_1904,In_664,In_888);
nand U1905 (N_1905,In_502,In_895);
or U1906 (N_1906,In_281,In_441);
or U1907 (N_1907,In_759,In_316);
nor U1908 (N_1908,In_863,In_482);
and U1909 (N_1909,In_841,In_638);
or U1910 (N_1910,In_460,In_194);
or U1911 (N_1911,In_759,In_2);
or U1912 (N_1912,In_258,In_403);
nor U1913 (N_1913,In_109,In_780);
or U1914 (N_1914,In_194,In_702);
or U1915 (N_1915,In_598,In_405);
or U1916 (N_1916,In_81,In_553);
and U1917 (N_1917,In_281,In_683);
nand U1918 (N_1918,In_405,In_865);
and U1919 (N_1919,In_489,In_217);
nand U1920 (N_1920,In_537,In_455);
nor U1921 (N_1921,In_872,In_111);
nand U1922 (N_1922,In_394,In_611);
and U1923 (N_1923,In_257,In_227);
and U1924 (N_1924,In_889,In_857);
or U1925 (N_1925,In_195,In_830);
and U1926 (N_1926,In_319,In_209);
nor U1927 (N_1927,In_60,In_177);
and U1928 (N_1928,In_973,In_154);
nor U1929 (N_1929,In_926,In_855);
and U1930 (N_1930,In_467,In_795);
nor U1931 (N_1931,In_918,In_166);
nand U1932 (N_1932,In_624,In_126);
nor U1933 (N_1933,In_952,In_380);
or U1934 (N_1934,In_638,In_547);
nor U1935 (N_1935,In_659,In_709);
and U1936 (N_1936,In_660,In_874);
and U1937 (N_1937,In_430,In_71);
or U1938 (N_1938,In_419,In_511);
or U1939 (N_1939,In_434,In_720);
nand U1940 (N_1940,In_118,In_988);
xnor U1941 (N_1941,In_872,In_627);
nand U1942 (N_1942,In_41,In_521);
nor U1943 (N_1943,In_139,In_602);
nor U1944 (N_1944,In_850,In_842);
nor U1945 (N_1945,In_723,In_683);
and U1946 (N_1946,In_439,In_513);
and U1947 (N_1947,In_561,In_35);
and U1948 (N_1948,In_185,In_115);
or U1949 (N_1949,In_211,In_498);
or U1950 (N_1950,In_883,In_326);
xnor U1951 (N_1951,In_263,In_594);
nor U1952 (N_1952,In_37,In_997);
or U1953 (N_1953,In_106,In_492);
nor U1954 (N_1954,In_208,In_219);
or U1955 (N_1955,In_856,In_830);
nor U1956 (N_1956,In_392,In_920);
or U1957 (N_1957,In_799,In_971);
and U1958 (N_1958,In_347,In_26);
nor U1959 (N_1959,In_166,In_734);
and U1960 (N_1960,In_204,In_956);
or U1961 (N_1961,In_442,In_706);
or U1962 (N_1962,In_378,In_723);
nor U1963 (N_1963,In_163,In_733);
or U1964 (N_1964,In_431,In_546);
nand U1965 (N_1965,In_445,In_105);
nor U1966 (N_1966,In_284,In_625);
and U1967 (N_1967,In_669,In_703);
nor U1968 (N_1968,In_867,In_76);
xnor U1969 (N_1969,In_568,In_430);
or U1970 (N_1970,In_818,In_784);
or U1971 (N_1971,In_817,In_394);
xnor U1972 (N_1972,In_979,In_388);
nor U1973 (N_1973,In_44,In_411);
nand U1974 (N_1974,In_288,In_642);
nor U1975 (N_1975,In_787,In_744);
or U1976 (N_1976,In_76,In_168);
or U1977 (N_1977,In_848,In_807);
nand U1978 (N_1978,In_65,In_965);
and U1979 (N_1979,In_208,In_648);
nand U1980 (N_1980,In_951,In_348);
or U1981 (N_1981,In_901,In_163);
and U1982 (N_1982,In_496,In_662);
or U1983 (N_1983,In_421,In_527);
nor U1984 (N_1984,In_607,In_690);
nand U1985 (N_1985,In_323,In_803);
nor U1986 (N_1986,In_299,In_546);
or U1987 (N_1987,In_930,In_252);
nor U1988 (N_1988,In_413,In_617);
and U1989 (N_1989,In_35,In_305);
and U1990 (N_1990,In_513,In_235);
nand U1991 (N_1991,In_387,In_100);
and U1992 (N_1992,In_354,In_87);
nand U1993 (N_1993,In_397,In_186);
and U1994 (N_1994,In_957,In_261);
xnor U1995 (N_1995,In_551,In_509);
nand U1996 (N_1996,In_594,In_607);
nor U1997 (N_1997,In_622,In_218);
and U1998 (N_1998,In_396,In_257);
nand U1999 (N_1999,In_120,In_372);
nor U2000 (N_2000,In_938,In_362);
nand U2001 (N_2001,In_820,In_790);
nor U2002 (N_2002,In_873,In_380);
nor U2003 (N_2003,In_498,In_756);
and U2004 (N_2004,In_540,In_968);
nand U2005 (N_2005,In_472,In_591);
xor U2006 (N_2006,In_63,In_336);
nand U2007 (N_2007,In_76,In_751);
xor U2008 (N_2008,In_909,In_279);
or U2009 (N_2009,In_72,In_582);
nor U2010 (N_2010,In_853,In_758);
or U2011 (N_2011,In_515,In_430);
nand U2012 (N_2012,In_891,In_846);
and U2013 (N_2013,In_971,In_455);
xor U2014 (N_2014,In_101,In_720);
or U2015 (N_2015,In_731,In_185);
or U2016 (N_2016,In_573,In_864);
nand U2017 (N_2017,In_88,In_918);
or U2018 (N_2018,In_906,In_272);
and U2019 (N_2019,In_835,In_249);
nor U2020 (N_2020,In_653,In_617);
or U2021 (N_2021,In_487,In_550);
or U2022 (N_2022,In_2,In_962);
xnor U2023 (N_2023,In_154,In_361);
nor U2024 (N_2024,In_936,In_351);
nand U2025 (N_2025,In_695,In_522);
or U2026 (N_2026,In_205,In_476);
or U2027 (N_2027,In_928,In_660);
and U2028 (N_2028,In_434,In_343);
nand U2029 (N_2029,In_924,In_638);
and U2030 (N_2030,In_469,In_743);
and U2031 (N_2031,In_250,In_537);
and U2032 (N_2032,In_118,In_315);
nand U2033 (N_2033,In_382,In_302);
nand U2034 (N_2034,In_571,In_703);
and U2035 (N_2035,In_549,In_934);
nand U2036 (N_2036,In_177,In_376);
nor U2037 (N_2037,In_258,In_140);
and U2038 (N_2038,In_593,In_722);
nand U2039 (N_2039,In_197,In_671);
and U2040 (N_2040,In_354,In_875);
or U2041 (N_2041,In_803,In_733);
nand U2042 (N_2042,In_363,In_480);
nor U2043 (N_2043,In_610,In_474);
nor U2044 (N_2044,In_971,In_55);
or U2045 (N_2045,In_204,In_858);
nor U2046 (N_2046,In_142,In_884);
nand U2047 (N_2047,In_61,In_248);
and U2048 (N_2048,In_300,In_691);
and U2049 (N_2049,In_660,In_499);
or U2050 (N_2050,In_961,In_631);
xor U2051 (N_2051,In_847,In_190);
or U2052 (N_2052,In_446,In_299);
or U2053 (N_2053,In_652,In_299);
nand U2054 (N_2054,In_906,In_249);
nand U2055 (N_2055,In_251,In_364);
and U2056 (N_2056,In_207,In_433);
nor U2057 (N_2057,In_450,In_77);
nand U2058 (N_2058,In_679,In_172);
nand U2059 (N_2059,In_833,In_55);
and U2060 (N_2060,In_616,In_902);
and U2061 (N_2061,In_502,In_563);
and U2062 (N_2062,In_227,In_841);
nand U2063 (N_2063,In_837,In_978);
nor U2064 (N_2064,In_818,In_304);
nand U2065 (N_2065,In_78,In_794);
or U2066 (N_2066,In_693,In_431);
nand U2067 (N_2067,In_341,In_493);
nand U2068 (N_2068,In_627,In_31);
nand U2069 (N_2069,In_452,In_376);
or U2070 (N_2070,In_30,In_756);
nand U2071 (N_2071,In_285,In_647);
nor U2072 (N_2072,In_151,In_302);
and U2073 (N_2073,In_307,In_339);
and U2074 (N_2074,In_95,In_285);
and U2075 (N_2075,In_803,In_282);
nand U2076 (N_2076,In_47,In_852);
and U2077 (N_2077,In_424,In_286);
nand U2078 (N_2078,In_442,In_147);
nand U2079 (N_2079,In_912,In_692);
nand U2080 (N_2080,In_853,In_623);
nand U2081 (N_2081,In_548,In_150);
and U2082 (N_2082,In_969,In_295);
nand U2083 (N_2083,In_25,In_693);
or U2084 (N_2084,In_380,In_313);
xor U2085 (N_2085,In_473,In_892);
nor U2086 (N_2086,In_553,In_557);
and U2087 (N_2087,In_695,In_154);
and U2088 (N_2088,In_421,In_358);
nor U2089 (N_2089,In_717,In_387);
nand U2090 (N_2090,In_822,In_507);
nor U2091 (N_2091,In_406,In_707);
or U2092 (N_2092,In_61,In_449);
and U2093 (N_2093,In_676,In_283);
nor U2094 (N_2094,In_405,In_638);
nand U2095 (N_2095,In_240,In_446);
nor U2096 (N_2096,In_291,In_372);
and U2097 (N_2097,In_414,In_332);
nor U2098 (N_2098,In_765,In_331);
nor U2099 (N_2099,In_530,In_752);
and U2100 (N_2100,In_838,In_866);
and U2101 (N_2101,In_65,In_626);
and U2102 (N_2102,In_568,In_706);
nor U2103 (N_2103,In_406,In_418);
and U2104 (N_2104,In_367,In_834);
nor U2105 (N_2105,In_173,In_429);
or U2106 (N_2106,In_800,In_832);
or U2107 (N_2107,In_472,In_944);
or U2108 (N_2108,In_997,In_880);
and U2109 (N_2109,In_619,In_40);
and U2110 (N_2110,In_80,In_765);
and U2111 (N_2111,In_347,In_847);
and U2112 (N_2112,In_559,In_282);
or U2113 (N_2113,In_927,In_410);
and U2114 (N_2114,In_282,In_804);
nand U2115 (N_2115,In_194,In_838);
and U2116 (N_2116,In_788,In_631);
nor U2117 (N_2117,In_44,In_42);
or U2118 (N_2118,In_536,In_520);
and U2119 (N_2119,In_909,In_659);
xnor U2120 (N_2120,In_476,In_291);
nor U2121 (N_2121,In_553,In_699);
nor U2122 (N_2122,In_108,In_663);
and U2123 (N_2123,In_211,In_312);
nor U2124 (N_2124,In_953,In_419);
and U2125 (N_2125,In_634,In_536);
nand U2126 (N_2126,In_708,In_278);
nand U2127 (N_2127,In_705,In_952);
and U2128 (N_2128,In_949,In_656);
and U2129 (N_2129,In_432,In_872);
nand U2130 (N_2130,In_317,In_971);
nor U2131 (N_2131,In_201,In_682);
nand U2132 (N_2132,In_808,In_120);
or U2133 (N_2133,In_28,In_85);
or U2134 (N_2134,In_465,In_117);
nand U2135 (N_2135,In_418,In_458);
nand U2136 (N_2136,In_747,In_853);
nand U2137 (N_2137,In_529,In_47);
and U2138 (N_2138,In_573,In_65);
nand U2139 (N_2139,In_275,In_860);
and U2140 (N_2140,In_360,In_510);
or U2141 (N_2141,In_821,In_515);
and U2142 (N_2142,In_346,In_258);
nor U2143 (N_2143,In_552,In_200);
xnor U2144 (N_2144,In_317,In_88);
or U2145 (N_2145,In_815,In_954);
and U2146 (N_2146,In_96,In_894);
and U2147 (N_2147,In_478,In_553);
nor U2148 (N_2148,In_408,In_238);
or U2149 (N_2149,In_905,In_825);
nor U2150 (N_2150,In_420,In_286);
nand U2151 (N_2151,In_56,In_932);
and U2152 (N_2152,In_293,In_697);
and U2153 (N_2153,In_537,In_935);
nor U2154 (N_2154,In_631,In_609);
or U2155 (N_2155,In_176,In_511);
nand U2156 (N_2156,In_841,In_822);
or U2157 (N_2157,In_61,In_331);
nand U2158 (N_2158,In_254,In_190);
and U2159 (N_2159,In_990,In_85);
nand U2160 (N_2160,In_606,In_70);
nand U2161 (N_2161,In_111,In_21);
nor U2162 (N_2162,In_97,In_36);
nor U2163 (N_2163,In_734,In_76);
or U2164 (N_2164,In_597,In_582);
or U2165 (N_2165,In_490,In_488);
and U2166 (N_2166,In_599,In_803);
or U2167 (N_2167,In_500,In_956);
nor U2168 (N_2168,In_309,In_638);
nand U2169 (N_2169,In_727,In_488);
or U2170 (N_2170,In_421,In_919);
or U2171 (N_2171,In_929,In_672);
and U2172 (N_2172,In_976,In_810);
or U2173 (N_2173,In_832,In_928);
and U2174 (N_2174,In_10,In_959);
and U2175 (N_2175,In_223,In_357);
nand U2176 (N_2176,In_422,In_811);
or U2177 (N_2177,In_473,In_411);
or U2178 (N_2178,In_314,In_591);
and U2179 (N_2179,In_969,In_900);
or U2180 (N_2180,In_718,In_561);
nand U2181 (N_2181,In_892,In_998);
nor U2182 (N_2182,In_307,In_503);
nor U2183 (N_2183,In_941,In_541);
nor U2184 (N_2184,In_377,In_182);
nor U2185 (N_2185,In_57,In_748);
nor U2186 (N_2186,In_788,In_687);
nand U2187 (N_2187,In_931,In_910);
nor U2188 (N_2188,In_272,In_485);
nor U2189 (N_2189,In_489,In_631);
nand U2190 (N_2190,In_796,In_394);
nor U2191 (N_2191,In_21,In_98);
or U2192 (N_2192,In_520,In_425);
nand U2193 (N_2193,In_881,In_418);
and U2194 (N_2194,In_603,In_847);
and U2195 (N_2195,In_775,In_890);
or U2196 (N_2196,In_615,In_193);
or U2197 (N_2197,In_265,In_160);
and U2198 (N_2198,In_525,In_981);
nor U2199 (N_2199,In_550,In_994);
nand U2200 (N_2200,In_823,In_983);
or U2201 (N_2201,In_694,In_95);
and U2202 (N_2202,In_347,In_392);
nor U2203 (N_2203,In_279,In_370);
or U2204 (N_2204,In_811,In_859);
or U2205 (N_2205,In_857,In_820);
and U2206 (N_2206,In_86,In_929);
or U2207 (N_2207,In_438,In_216);
nor U2208 (N_2208,In_373,In_205);
nand U2209 (N_2209,In_198,In_850);
xnor U2210 (N_2210,In_688,In_38);
nand U2211 (N_2211,In_211,In_517);
or U2212 (N_2212,In_83,In_719);
or U2213 (N_2213,In_654,In_205);
nand U2214 (N_2214,In_342,In_62);
and U2215 (N_2215,In_315,In_271);
and U2216 (N_2216,In_835,In_14);
nor U2217 (N_2217,In_543,In_506);
and U2218 (N_2218,In_576,In_872);
nand U2219 (N_2219,In_547,In_790);
nand U2220 (N_2220,In_237,In_156);
and U2221 (N_2221,In_296,In_676);
nand U2222 (N_2222,In_98,In_537);
nand U2223 (N_2223,In_41,In_105);
or U2224 (N_2224,In_254,In_874);
nor U2225 (N_2225,In_587,In_543);
nand U2226 (N_2226,In_477,In_663);
nor U2227 (N_2227,In_311,In_142);
nor U2228 (N_2228,In_250,In_232);
xor U2229 (N_2229,In_218,In_991);
or U2230 (N_2230,In_484,In_911);
or U2231 (N_2231,In_516,In_169);
or U2232 (N_2232,In_278,In_367);
or U2233 (N_2233,In_381,In_277);
and U2234 (N_2234,In_681,In_293);
nor U2235 (N_2235,In_54,In_206);
nor U2236 (N_2236,In_95,In_296);
nand U2237 (N_2237,In_572,In_799);
or U2238 (N_2238,In_524,In_517);
nor U2239 (N_2239,In_725,In_391);
and U2240 (N_2240,In_287,In_300);
and U2241 (N_2241,In_508,In_656);
and U2242 (N_2242,In_437,In_159);
or U2243 (N_2243,In_680,In_517);
nor U2244 (N_2244,In_41,In_607);
and U2245 (N_2245,In_691,In_481);
and U2246 (N_2246,In_91,In_604);
nor U2247 (N_2247,In_830,In_609);
nor U2248 (N_2248,In_769,In_916);
nand U2249 (N_2249,In_972,In_974);
nor U2250 (N_2250,In_511,In_130);
nor U2251 (N_2251,In_235,In_939);
nor U2252 (N_2252,In_505,In_39);
nand U2253 (N_2253,In_959,In_736);
nand U2254 (N_2254,In_440,In_709);
nor U2255 (N_2255,In_756,In_628);
nor U2256 (N_2256,In_688,In_163);
xnor U2257 (N_2257,In_43,In_117);
nor U2258 (N_2258,In_412,In_320);
nand U2259 (N_2259,In_905,In_539);
and U2260 (N_2260,In_555,In_776);
nand U2261 (N_2261,In_383,In_967);
nor U2262 (N_2262,In_554,In_384);
and U2263 (N_2263,In_691,In_458);
nor U2264 (N_2264,In_605,In_242);
and U2265 (N_2265,In_472,In_513);
or U2266 (N_2266,In_25,In_926);
nand U2267 (N_2267,In_644,In_74);
nand U2268 (N_2268,In_684,In_498);
xnor U2269 (N_2269,In_114,In_964);
xor U2270 (N_2270,In_142,In_399);
nor U2271 (N_2271,In_915,In_416);
nor U2272 (N_2272,In_832,In_755);
and U2273 (N_2273,In_991,In_100);
or U2274 (N_2274,In_502,In_850);
or U2275 (N_2275,In_643,In_233);
nor U2276 (N_2276,In_335,In_672);
nand U2277 (N_2277,In_170,In_455);
or U2278 (N_2278,In_259,In_442);
nor U2279 (N_2279,In_566,In_798);
or U2280 (N_2280,In_39,In_600);
or U2281 (N_2281,In_277,In_56);
nand U2282 (N_2282,In_842,In_401);
nand U2283 (N_2283,In_711,In_276);
nor U2284 (N_2284,In_271,In_684);
nand U2285 (N_2285,In_605,In_131);
or U2286 (N_2286,In_470,In_168);
and U2287 (N_2287,In_997,In_361);
and U2288 (N_2288,In_578,In_605);
or U2289 (N_2289,In_309,In_787);
nand U2290 (N_2290,In_245,In_454);
nand U2291 (N_2291,In_846,In_727);
and U2292 (N_2292,In_818,In_722);
and U2293 (N_2293,In_302,In_808);
nor U2294 (N_2294,In_953,In_222);
or U2295 (N_2295,In_413,In_50);
nor U2296 (N_2296,In_798,In_727);
and U2297 (N_2297,In_127,In_866);
or U2298 (N_2298,In_707,In_903);
or U2299 (N_2299,In_29,In_45);
nand U2300 (N_2300,In_51,In_973);
or U2301 (N_2301,In_936,In_382);
nand U2302 (N_2302,In_684,In_266);
nor U2303 (N_2303,In_85,In_924);
nor U2304 (N_2304,In_266,In_809);
xnor U2305 (N_2305,In_784,In_666);
or U2306 (N_2306,In_588,In_668);
nand U2307 (N_2307,In_929,In_432);
and U2308 (N_2308,In_509,In_230);
or U2309 (N_2309,In_799,In_328);
nand U2310 (N_2310,In_745,In_863);
or U2311 (N_2311,In_210,In_966);
nor U2312 (N_2312,In_231,In_618);
and U2313 (N_2313,In_656,In_982);
and U2314 (N_2314,In_543,In_966);
and U2315 (N_2315,In_730,In_649);
or U2316 (N_2316,In_380,In_759);
nand U2317 (N_2317,In_813,In_486);
nand U2318 (N_2318,In_128,In_378);
nand U2319 (N_2319,In_597,In_3);
nand U2320 (N_2320,In_217,In_570);
nor U2321 (N_2321,In_196,In_130);
and U2322 (N_2322,In_613,In_385);
xor U2323 (N_2323,In_697,In_246);
nand U2324 (N_2324,In_794,In_516);
nor U2325 (N_2325,In_504,In_212);
xnor U2326 (N_2326,In_477,In_868);
and U2327 (N_2327,In_828,In_517);
or U2328 (N_2328,In_237,In_128);
or U2329 (N_2329,In_171,In_540);
nand U2330 (N_2330,In_393,In_985);
or U2331 (N_2331,In_703,In_44);
or U2332 (N_2332,In_926,In_248);
nor U2333 (N_2333,In_602,In_616);
nand U2334 (N_2334,In_148,In_447);
nand U2335 (N_2335,In_440,In_604);
nand U2336 (N_2336,In_818,In_627);
nand U2337 (N_2337,In_842,In_458);
or U2338 (N_2338,In_828,In_939);
nor U2339 (N_2339,In_93,In_993);
and U2340 (N_2340,In_913,In_743);
nor U2341 (N_2341,In_143,In_592);
nor U2342 (N_2342,In_47,In_938);
nor U2343 (N_2343,In_982,In_600);
nor U2344 (N_2344,In_406,In_766);
nor U2345 (N_2345,In_331,In_687);
and U2346 (N_2346,In_102,In_97);
xnor U2347 (N_2347,In_272,In_594);
nor U2348 (N_2348,In_749,In_332);
nand U2349 (N_2349,In_524,In_440);
and U2350 (N_2350,In_211,In_476);
xor U2351 (N_2351,In_464,In_679);
or U2352 (N_2352,In_141,In_155);
nor U2353 (N_2353,In_466,In_870);
or U2354 (N_2354,In_274,In_50);
and U2355 (N_2355,In_415,In_133);
nor U2356 (N_2356,In_479,In_108);
or U2357 (N_2357,In_812,In_555);
nor U2358 (N_2358,In_246,In_503);
nor U2359 (N_2359,In_324,In_735);
nand U2360 (N_2360,In_566,In_831);
or U2361 (N_2361,In_540,In_960);
and U2362 (N_2362,In_185,In_376);
nor U2363 (N_2363,In_794,In_208);
and U2364 (N_2364,In_904,In_63);
and U2365 (N_2365,In_696,In_105);
or U2366 (N_2366,In_13,In_968);
or U2367 (N_2367,In_451,In_534);
nor U2368 (N_2368,In_701,In_914);
nand U2369 (N_2369,In_534,In_458);
or U2370 (N_2370,In_561,In_792);
nand U2371 (N_2371,In_763,In_97);
or U2372 (N_2372,In_296,In_137);
and U2373 (N_2373,In_451,In_503);
and U2374 (N_2374,In_132,In_473);
or U2375 (N_2375,In_38,In_587);
and U2376 (N_2376,In_256,In_425);
nor U2377 (N_2377,In_122,In_351);
and U2378 (N_2378,In_563,In_457);
and U2379 (N_2379,In_228,In_42);
or U2380 (N_2380,In_897,In_691);
nor U2381 (N_2381,In_710,In_799);
nor U2382 (N_2382,In_544,In_470);
nor U2383 (N_2383,In_54,In_699);
nor U2384 (N_2384,In_239,In_805);
or U2385 (N_2385,In_993,In_974);
nor U2386 (N_2386,In_698,In_508);
and U2387 (N_2387,In_755,In_496);
or U2388 (N_2388,In_150,In_367);
or U2389 (N_2389,In_515,In_553);
and U2390 (N_2390,In_45,In_12);
or U2391 (N_2391,In_469,In_752);
and U2392 (N_2392,In_574,In_89);
and U2393 (N_2393,In_523,In_899);
nand U2394 (N_2394,In_149,In_488);
or U2395 (N_2395,In_811,In_771);
nor U2396 (N_2396,In_206,In_209);
nor U2397 (N_2397,In_727,In_134);
nor U2398 (N_2398,In_134,In_639);
and U2399 (N_2399,In_4,In_166);
and U2400 (N_2400,In_499,In_69);
xor U2401 (N_2401,In_130,In_790);
nor U2402 (N_2402,In_30,In_282);
nand U2403 (N_2403,In_629,In_209);
and U2404 (N_2404,In_110,In_735);
and U2405 (N_2405,In_478,In_5);
or U2406 (N_2406,In_995,In_284);
nor U2407 (N_2407,In_586,In_298);
nand U2408 (N_2408,In_261,In_817);
nand U2409 (N_2409,In_94,In_391);
or U2410 (N_2410,In_678,In_629);
and U2411 (N_2411,In_492,In_411);
and U2412 (N_2412,In_211,In_358);
or U2413 (N_2413,In_746,In_27);
or U2414 (N_2414,In_542,In_274);
or U2415 (N_2415,In_286,In_64);
nor U2416 (N_2416,In_253,In_671);
nor U2417 (N_2417,In_927,In_366);
or U2418 (N_2418,In_57,In_923);
and U2419 (N_2419,In_945,In_987);
or U2420 (N_2420,In_295,In_118);
nor U2421 (N_2421,In_707,In_351);
nor U2422 (N_2422,In_650,In_964);
nor U2423 (N_2423,In_364,In_284);
nor U2424 (N_2424,In_345,In_946);
nand U2425 (N_2425,In_481,In_516);
nand U2426 (N_2426,In_544,In_119);
or U2427 (N_2427,In_726,In_490);
or U2428 (N_2428,In_689,In_272);
nor U2429 (N_2429,In_52,In_776);
nor U2430 (N_2430,In_12,In_17);
nor U2431 (N_2431,In_916,In_417);
or U2432 (N_2432,In_312,In_608);
nand U2433 (N_2433,In_19,In_110);
nand U2434 (N_2434,In_999,In_761);
or U2435 (N_2435,In_775,In_926);
or U2436 (N_2436,In_933,In_781);
nor U2437 (N_2437,In_866,In_683);
and U2438 (N_2438,In_422,In_535);
xnor U2439 (N_2439,In_686,In_924);
or U2440 (N_2440,In_468,In_752);
or U2441 (N_2441,In_292,In_441);
or U2442 (N_2442,In_237,In_106);
and U2443 (N_2443,In_391,In_480);
or U2444 (N_2444,In_187,In_465);
nor U2445 (N_2445,In_941,In_652);
nand U2446 (N_2446,In_986,In_67);
and U2447 (N_2447,In_857,In_32);
nor U2448 (N_2448,In_990,In_920);
nand U2449 (N_2449,In_770,In_241);
nor U2450 (N_2450,In_372,In_416);
xor U2451 (N_2451,In_666,In_168);
or U2452 (N_2452,In_722,In_505);
nand U2453 (N_2453,In_98,In_511);
or U2454 (N_2454,In_683,In_358);
and U2455 (N_2455,In_641,In_69);
nor U2456 (N_2456,In_112,In_42);
or U2457 (N_2457,In_533,In_397);
nand U2458 (N_2458,In_875,In_724);
nor U2459 (N_2459,In_291,In_731);
nor U2460 (N_2460,In_643,In_522);
nand U2461 (N_2461,In_345,In_794);
and U2462 (N_2462,In_976,In_755);
nand U2463 (N_2463,In_397,In_337);
nor U2464 (N_2464,In_153,In_787);
or U2465 (N_2465,In_43,In_952);
nor U2466 (N_2466,In_655,In_285);
and U2467 (N_2467,In_569,In_535);
nor U2468 (N_2468,In_800,In_280);
or U2469 (N_2469,In_402,In_963);
nor U2470 (N_2470,In_91,In_518);
or U2471 (N_2471,In_733,In_716);
xor U2472 (N_2472,In_158,In_991);
and U2473 (N_2473,In_895,In_582);
nand U2474 (N_2474,In_257,In_999);
xnor U2475 (N_2475,In_673,In_535);
nor U2476 (N_2476,In_263,In_597);
or U2477 (N_2477,In_613,In_594);
nand U2478 (N_2478,In_403,In_332);
and U2479 (N_2479,In_63,In_168);
and U2480 (N_2480,In_956,In_709);
nand U2481 (N_2481,In_952,In_475);
nand U2482 (N_2482,In_943,In_482);
or U2483 (N_2483,In_307,In_170);
nand U2484 (N_2484,In_296,In_880);
and U2485 (N_2485,In_933,In_617);
and U2486 (N_2486,In_673,In_308);
nand U2487 (N_2487,In_545,In_15);
and U2488 (N_2488,In_591,In_694);
nor U2489 (N_2489,In_379,In_453);
nand U2490 (N_2490,In_604,In_597);
and U2491 (N_2491,In_720,In_771);
nand U2492 (N_2492,In_16,In_901);
nor U2493 (N_2493,In_447,In_433);
or U2494 (N_2494,In_253,In_157);
nor U2495 (N_2495,In_267,In_451);
nor U2496 (N_2496,In_742,In_726);
nand U2497 (N_2497,In_974,In_325);
nand U2498 (N_2498,In_282,In_594);
and U2499 (N_2499,In_20,In_972);
or U2500 (N_2500,N_2081,N_134);
or U2501 (N_2501,N_2160,N_874);
or U2502 (N_2502,N_450,N_2021);
nor U2503 (N_2503,N_491,N_1962);
nand U2504 (N_2504,N_866,N_541);
nand U2505 (N_2505,N_2079,N_27);
or U2506 (N_2506,N_72,N_324);
nor U2507 (N_2507,N_945,N_965);
and U2508 (N_2508,N_1036,N_2307);
nor U2509 (N_2509,N_1181,N_1875);
and U2510 (N_2510,N_2284,N_1415);
or U2511 (N_2511,N_22,N_829);
nand U2512 (N_2512,N_519,N_219);
nand U2513 (N_2513,N_103,N_1747);
nand U2514 (N_2514,N_327,N_1932);
or U2515 (N_2515,N_2147,N_173);
or U2516 (N_2516,N_1558,N_1233);
or U2517 (N_2517,N_2106,N_2302);
nor U2518 (N_2518,N_1766,N_280);
nor U2519 (N_2519,N_851,N_675);
nor U2520 (N_2520,N_162,N_1318);
or U2521 (N_2521,N_1987,N_959);
nand U2522 (N_2522,N_1300,N_983);
nand U2523 (N_2523,N_1539,N_1907);
and U2524 (N_2524,N_941,N_662);
nor U2525 (N_2525,N_1629,N_687);
and U2526 (N_2526,N_2199,N_585);
nor U2527 (N_2527,N_1247,N_1693);
or U2528 (N_2528,N_2159,N_427);
nor U2529 (N_2529,N_465,N_2188);
or U2530 (N_2530,N_1941,N_644);
or U2531 (N_2531,N_1441,N_270);
and U2532 (N_2532,N_839,N_1966);
or U2533 (N_2533,N_1027,N_1787);
and U2534 (N_2534,N_2367,N_78);
or U2535 (N_2535,N_1072,N_1597);
and U2536 (N_2536,N_1136,N_57);
or U2537 (N_2537,N_216,N_2185);
and U2538 (N_2538,N_735,N_1492);
or U2539 (N_2539,N_2399,N_2195);
or U2540 (N_2540,N_323,N_489);
nor U2541 (N_2541,N_1807,N_770);
nor U2542 (N_2542,N_272,N_1420);
nor U2543 (N_2543,N_1196,N_1778);
nor U2544 (N_2544,N_249,N_1288);
or U2545 (N_2545,N_1674,N_2049);
nor U2546 (N_2546,N_2155,N_651);
or U2547 (N_2547,N_1719,N_157);
nand U2548 (N_2548,N_1982,N_811);
and U2549 (N_2549,N_1725,N_133);
or U2550 (N_2550,N_437,N_440);
or U2551 (N_2551,N_1600,N_830);
nor U2552 (N_2552,N_1582,N_1180);
nand U2553 (N_2553,N_321,N_1283);
and U2554 (N_2554,N_2388,N_316);
nor U2555 (N_2555,N_2067,N_1240);
nor U2556 (N_2556,N_1595,N_1699);
nand U2557 (N_2557,N_747,N_2212);
nand U2558 (N_2558,N_1642,N_1955);
or U2559 (N_2559,N_225,N_915);
nor U2560 (N_2560,N_1411,N_867);
and U2561 (N_2561,N_412,N_118);
and U2562 (N_2562,N_181,N_1089);
nand U2563 (N_2563,N_24,N_1111);
or U2564 (N_2564,N_1248,N_643);
and U2565 (N_2565,N_2259,N_198);
xnor U2566 (N_2566,N_862,N_1447);
nand U2567 (N_2567,N_424,N_1227);
and U2568 (N_2568,N_661,N_1236);
nor U2569 (N_2569,N_574,N_2277);
nand U2570 (N_2570,N_387,N_766);
or U2571 (N_2571,N_2347,N_325);
and U2572 (N_2572,N_1826,N_533);
or U2573 (N_2573,N_2036,N_1745);
and U2574 (N_2574,N_371,N_2357);
or U2575 (N_2575,N_1351,N_1495);
or U2576 (N_2576,N_158,N_711);
or U2577 (N_2577,N_375,N_479);
nor U2578 (N_2578,N_1781,N_1533);
nor U2579 (N_2579,N_749,N_2055);
or U2580 (N_2580,N_1664,N_2436);
and U2581 (N_2581,N_1880,N_632);
and U2582 (N_2582,N_1093,N_968);
nand U2583 (N_2583,N_495,N_2132);
nor U2584 (N_2584,N_396,N_1366);
nand U2585 (N_2585,N_2197,N_1692);
or U2586 (N_2586,N_1127,N_2270);
nor U2587 (N_2587,N_1849,N_425);
nand U2588 (N_2588,N_691,N_456);
nor U2589 (N_2589,N_2348,N_123);
nand U2590 (N_2590,N_1617,N_1273);
and U2591 (N_2591,N_2070,N_1919);
or U2592 (N_2592,N_799,N_302);
and U2593 (N_2593,N_842,N_1296);
nor U2594 (N_2594,N_765,N_1520);
and U2595 (N_2595,N_1491,N_403);
nand U2596 (N_2596,N_1455,N_1347);
nor U2597 (N_2597,N_1147,N_508);
or U2598 (N_2598,N_1293,N_580);
nand U2599 (N_2599,N_1626,N_2017);
and U2600 (N_2600,N_2107,N_716);
xor U2601 (N_2601,N_1678,N_531);
nand U2602 (N_2602,N_459,N_995);
nor U2603 (N_2603,N_909,N_1334);
nand U2604 (N_2604,N_1834,N_1446);
and U2605 (N_2605,N_1910,N_1731);
or U2606 (N_2606,N_806,N_934);
or U2607 (N_2607,N_50,N_1365);
or U2608 (N_2608,N_2114,N_628);
or U2609 (N_2609,N_2222,N_721);
nand U2610 (N_2610,N_2464,N_1663);
or U2611 (N_2611,N_53,N_534);
nor U2612 (N_2612,N_1020,N_2254);
nor U2613 (N_2613,N_1398,N_1412);
nand U2614 (N_2614,N_1499,N_51);
and U2615 (N_2615,N_1439,N_415);
nor U2616 (N_2616,N_1771,N_989);
nand U2617 (N_2617,N_1490,N_2450);
nor U2618 (N_2618,N_1425,N_1218);
and U2619 (N_2619,N_1454,N_523);
nand U2620 (N_2620,N_1906,N_816);
nand U2621 (N_2621,N_2475,N_1418);
and U2622 (N_2622,N_448,N_1339);
and U2623 (N_2623,N_512,N_1200);
or U2624 (N_2624,N_1104,N_1079);
and U2625 (N_2625,N_468,N_75);
nand U2626 (N_2626,N_1717,N_226);
or U2627 (N_2627,N_596,N_1610);
and U2628 (N_2628,N_2085,N_414);
or U2629 (N_2629,N_1637,N_761);
nand U2630 (N_2630,N_2310,N_2059);
nor U2631 (N_2631,N_1917,N_366);
or U2632 (N_2632,N_802,N_1060);
nor U2633 (N_2633,N_733,N_1805);
and U2634 (N_2634,N_926,N_429);
or U2635 (N_2635,N_602,N_1094);
nand U2636 (N_2636,N_573,N_294);
nand U2637 (N_2637,N_1523,N_1677);
or U2638 (N_2638,N_167,N_201);
or U2639 (N_2639,N_358,N_621);
and U2640 (N_2640,N_681,N_992);
nand U2641 (N_2641,N_1464,N_1914);
nor U2642 (N_2642,N_449,N_99);
nor U2643 (N_2643,N_2193,N_1574);
or U2644 (N_2644,N_1676,N_266);
nand U2645 (N_2645,N_1791,N_762);
or U2646 (N_2646,N_738,N_790);
and U2647 (N_2647,N_284,N_2335);
and U2648 (N_2648,N_1067,N_1080);
and U2649 (N_2649,N_406,N_2285);
or U2650 (N_2650,N_115,N_1225);
or U2651 (N_2651,N_2172,N_2022);
or U2652 (N_2652,N_2250,N_564);
and U2653 (N_2653,N_1668,N_312);
and U2654 (N_2654,N_1115,N_2040);
nor U2655 (N_2655,N_530,N_946);
nor U2656 (N_2656,N_1018,N_125);
or U2657 (N_2657,N_1945,N_767);
nand U2658 (N_2658,N_1947,N_692);
and U2659 (N_2659,N_1278,N_1728);
nor U2660 (N_2660,N_402,N_341);
and U2661 (N_2661,N_273,N_1666);
or U2662 (N_2662,N_795,N_49);
nand U2663 (N_2663,N_2192,N_1623);
nand U2664 (N_2664,N_2170,N_1249);
nor U2665 (N_2665,N_943,N_746);
nor U2666 (N_2666,N_1265,N_1484);
or U2667 (N_2667,N_1475,N_559);
and U2668 (N_2668,N_1011,N_2390);
or U2669 (N_2669,N_433,N_1156);
and U2670 (N_2670,N_224,N_2334);
or U2671 (N_2671,N_2297,N_1546);
and U2672 (N_2672,N_346,N_475);
or U2673 (N_2673,N_1948,N_2306);
nand U2674 (N_2674,N_993,N_1815);
and U2675 (N_2675,N_1723,N_1860);
or U2676 (N_2676,N_2374,N_2445);
and U2677 (N_2677,N_26,N_870);
or U2678 (N_2678,N_146,N_2029);
or U2679 (N_2679,N_430,N_2455);
and U2680 (N_2680,N_84,N_357);
and U2681 (N_2681,N_2123,N_1665);
nor U2682 (N_2682,N_595,N_1496);
nor U2683 (N_2683,N_1762,N_901);
nor U2684 (N_2684,N_760,N_947);
nand U2685 (N_2685,N_885,N_1209);
nor U2686 (N_2686,N_1368,N_1197);
and U2687 (N_2687,N_1607,N_1034);
and U2688 (N_2688,N_2339,N_1129);
nor U2689 (N_2689,N_2099,N_546);
or U2690 (N_2690,N_1633,N_1592);
xnor U2691 (N_2691,N_1126,N_895);
and U2692 (N_2692,N_2331,N_1062);
or U2693 (N_2693,N_1952,N_1133);
and U2694 (N_2694,N_554,N_82);
and U2695 (N_2695,N_1980,N_1088);
nor U2696 (N_2696,N_2325,N_1243);
nor U2697 (N_2697,N_659,N_929);
and U2698 (N_2698,N_251,N_2109);
nor U2699 (N_2699,N_111,N_1853);
and U2700 (N_2700,N_2257,N_834);
or U2701 (N_2701,N_859,N_1501);
nand U2702 (N_2702,N_382,N_44);
and U2703 (N_2703,N_177,N_789);
nor U2704 (N_2704,N_652,N_1322);
nor U2705 (N_2705,N_473,N_488);
nand U2706 (N_2706,N_1304,N_2171);
or U2707 (N_2707,N_259,N_2377);
nand U2708 (N_2708,N_431,N_2373);
nor U2709 (N_2709,N_1896,N_1868);
nor U2710 (N_2710,N_306,N_278);
xnor U2711 (N_2711,N_863,N_1114);
and U2712 (N_2712,N_1700,N_1065);
nor U2713 (N_2713,N_1410,N_1904);
and U2714 (N_2714,N_2096,N_229);
nand U2715 (N_2715,N_2312,N_883);
nor U2716 (N_2716,N_1383,N_1989);
or U2717 (N_2717,N_1172,N_1949);
nand U2718 (N_2718,N_2174,N_2002);
or U2719 (N_2719,N_1306,N_10);
xnor U2720 (N_2720,N_887,N_973);
nand U2721 (N_2721,N_1810,N_630);
or U2722 (N_2722,N_2318,N_1075);
or U2723 (N_2723,N_209,N_2336);
or U2724 (N_2724,N_258,N_2379);
nand U2725 (N_2725,N_2164,N_1557);
and U2726 (N_2726,N_2191,N_1603);
nor U2727 (N_2727,N_61,N_1330);
nand U2728 (N_2728,N_309,N_138);
and U2729 (N_2729,N_1930,N_742);
or U2730 (N_2730,N_187,N_2416);
or U2731 (N_2731,N_361,N_1754);
nand U2732 (N_2732,N_1797,N_2411);
or U2733 (N_2733,N_360,N_218);
nand U2734 (N_2734,N_2052,N_2382);
or U2735 (N_2735,N_1310,N_2088);
nand U2736 (N_2736,N_2241,N_2104);
and U2737 (N_2737,N_1489,N_496);
or U2738 (N_2738,N_108,N_2208);
and U2739 (N_2739,N_1695,N_389);
or U2740 (N_2740,N_1924,N_2095);
nand U2741 (N_2741,N_2414,N_1673);
nor U2742 (N_2742,N_1046,N_1097);
nand U2743 (N_2743,N_2053,N_1482);
or U2744 (N_2744,N_2442,N_961);
or U2745 (N_2745,N_1809,N_1513);
nand U2746 (N_2746,N_1006,N_1528);
nand U2747 (N_2747,N_1052,N_1636);
nor U2748 (N_2748,N_670,N_707);
and U2749 (N_2749,N_2082,N_1162);
and U2750 (N_2750,N_1378,N_744);
nand U2751 (N_2751,N_1445,N_855);
nor U2752 (N_2752,N_1979,N_2056);
or U2753 (N_2753,N_2314,N_117);
xor U2754 (N_2754,N_1843,N_1159);
xor U2755 (N_2755,N_757,N_1993);
and U2756 (N_2756,N_1871,N_1393);
and U2757 (N_2757,N_1427,N_1707);
nor U2758 (N_2758,N_1995,N_2326);
and U2759 (N_2759,N_1239,N_2295);
nand U2760 (N_2760,N_900,N_2069);
and U2761 (N_2761,N_2043,N_1083);
nand U2762 (N_2762,N_422,N_1171);
or U2763 (N_2763,N_1685,N_680);
or U2764 (N_2764,N_977,N_2409);
or U2765 (N_2765,N_568,N_168);
or U2766 (N_2766,N_121,N_1294);
nor U2767 (N_2767,N_679,N_367);
and U2768 (N_2768,N_369,N_1505);
xor U2769 (N_2769,N_555,N_128);
nor U2770 (N_2770,N_2299,N_763);
and U2771 (N_2771,N_2395,N_1892);
or U2772 (N_2772,N_1658,N_2420);
or U2773 (N_2773,N_1784,N_1231);
nor U2774 (N_2774,N_1158,N_1887);
and U2775 (N_2775,N_798,N_2240);
nand U2776 (N_2776,N_764,N_2216);
or U2777 (N_2777,N_1481,N_1184);
nand U2778 (N_2778,N_1937,N_1399);
nor U2779 (N_2779,N_2189,N_2173);
nor U2780 (N_2780,N_1929,N_166);
or U2781 (N_2781,N_1369,N_1063);
or U2782 (N_2782,N_1132,N_337);
and U2783 (N_2783,N_288,N_524);
or U2784 (N_2784,N_516,N_1836);
nand U2785 (N_2785,N_2473,N_1656);
and U2786 (N_2786,N_1169,N_2417);
and U2787 (N_2787,N_1396,N_1748);
nor U2788 (N_2788,N_1806,N_1045);
and U2789 (N_2789,N_363,N_1788);
nor U2790 (N_2790,N_1370,N_2272);
nand U2791 (N_2791,N_729,N_1584);
and U2792 (N_2792,N_2231,N_624);
and U2793 (N_2793,N_1462,N_2032);
or U2794 (N_2794,N_1654,N_996);
and U2795 (N_2795,N_188,N_1869);
or U2796 (N_2796,N_1028,N_570);
nor U2797 (N_2797,N_186,N_731);
or U2798 (N_2798,N_1206,N_2480);
nand U2799 (N_2799,N_2322,N_2349);
nor U2800 (N_2800,N_1422,N_598);
nand U2801 (N_2801,N_2204,N_2457);
nor U2802 (N_2802,N_322,N_876);
nor U2803 (N_2803,N_2202,N_654);
nand U2804 (N_2804,N_1486,N_974);
or U2805 (N_2805,N_1031,N_1992);
and U2806 (N_2806,N_2156,N_328);
and U2807 (N_2807,N_776,N_2038);
nor U2808 (N_2808,N_1732,N_809);
and U2809 (N_2809,N_77,N_840);
and U2810 (N_2810,N_1235,N_1715);
or U2811 (N_2811,N_476,N_1389);
nand U2812 (N_2812,N_285,N_2361);
and U2813 (N_2813,N_107,N_1615);
nor U2814 (N_2814,N_1388,N_206);
nand U2815 (N_2815,N_2364,N_2075);
nor U2816 (N_2816,N_690,N_1532);
nor U2817 (N_2817,N_11,N_1145);
nand U2818 (N_2818,N_2316,N_1795);
nor U2819 (N_2819,N_447,N_1360);
and U2820 (N_2820,N_2383,N_1219);
and U2821 (N_2821,N_2265,N_812);
nand U2822 (N_2822,N_635,N_2003);
and U2823 (N_2823,N_149,N_2482);
xor U2824 (N_2824,N_2111,N_263);
or U2825 (N_2825,N_395,N_2186);
or U2826 (N_2826,N_2352,N_33);
nand U2827 (N_2827,N_21,N_1276);
nor U2828 (N_2828,N_2267,N_1825);
nand U2829 (N_2829,N_2140,N_1988);
nor U2830 (N_2830,N_2015,N_2167);
nor U2831 (N_2831,N_1244,N_1085);
and U2832 (N_2832,N_241,N_1405);
nand U2833 (N_2833,N_669,N_308);
nand U2834 (N_2834,N_1400,N_1324);
or U2835 (N_2835,N_2091,N_804);
or U2836 (N_2836,N_2498,N_1440);
and U2837 (N_2837,N_1477,N_2320);
nand U2838 (N_2838,N_469,N_478);
nand U2839 (N_2839,N_1182,N_1024);
nor U2840 (N_2840,N_1845,N_1530);
nand U2841 (N_2841,N_1912,N_1165);
nor U2842 (N_2842,N_1572,N_693);
or U2843 (N_2843,N_674,N_1119);
nor U2844 (N_2844,N_1261,N_2253);
nand U2845 (N_2845,N_1652,N_212);
and U2846 (N_2846,N_1434,N_65);
nand U2847 (N_2847,N_36,N_1599);
or U2848 (N_2848,N_301,N_1620);
and U2849 (N_2849,N_1585,N_1918);
nand U2850 (N_2850,N_1155,N_1721);
or U2851 (N_2851,N_1217,N_317);
nor U2852 (N_2852,N_1752,N_1632);
nand U2853 (N_2853,N_1022,N_163);
and U2854 (N_2854,N_1109,N_1385);
nor U2855 (N_2855,N_2486,N_1429);
and U2856 (N_2856,N_1886,N_1312);
nand U2857 (N_2857,N_754,N_1936);
nor U2858 (N_2858,N_66,N_2403);
and U2859 (N_2859,N_2175,N_2404);
or U2860 (N_2860,N_2050,N_247);
or U2861 (N_2861,N_676,N_820);
nor U2862 (N_2862,N_647,N_2115);
nand U2863 (N_2863,N_1569,N_2385);
nor U2864 (N_2864,N_420,N_1140);
and U2865 (N_2865,N_2093,N_927);
or U2866 (N_2866,N_2415,N_688);
or U2867 (N_2867,N_882,N_1804);
nor U2868 (N_2868,N_1280,N_1812);
or U2869 (N_2869,N_1472,N_1355);
and U2870 (N_2870,N_1307,N_1198);
nor U2871 (N_2871,N_7,N_877);
and U2872 (N_2872,N_2440,N_1091);
or U2873 (N_2873,N_1163,N_550);
nand U2874 (N_2874,N_2145,N_792);
or U2875 (N_2875,N_1551,N_1271);
nor U2876 (N_2876,N_979,N_1559);
nand U2877 (N_2877,N_265,N_1047);
nand U2878 (N_2878,N_2426,N_1984);
nand U2879 (N_2879,N_1401,N_1905);
or U2880 (N_2880,N_1879,N_1576);
or U2881 (N_2881,N_1716,N_383);
or U2882 (N_2882,N_769,N_626);
and U2883 (N_2883,N_1769,N_2124);
or U2884 (N_2884,N_2278,N_1562);
nand U2885 (N_2885,N_1195,N_58);
nor U2886 (N_2886,N_1641,N_1059);
nor U2887 (N_2887,N_1627,N_1598);
nand U2888 (N_2888,N_319,N_141);
nand U2889 (N_2889,N_1759,N_1961);
and U2890 (N_2890,N_405,N_1403);
nor U2891 (N_2891,N_233,N_994);
nand U2892 (N_2892,N_2378,N_2101);
nand U2893 (N_2893,N_1702,N_2087);
or U2894 (N_2894,N_932,N_1618);
nand U2895 (N_2895,N_2353,N_345);
or U2896 (N_2896,N_1733,N_230);
and U2897 (N_2897,N_718,N_794);
nor U2898 (N_2898,N_730,N_1529);
nand U2899 (N_2899,N_828,N_1511);
or U2900 (N_2900,N_1096,N_728);
or U2901 (N_2901,N_1210,N_813);
and U2902 (N_2902,N_1026,N_503);
or U2903 (N_2903,N_1359,N_339);
or U2904 (N_2904,N_1755,N_9);
nor U2905 (N_2905,N_1095,N_2100);
nor U2906 (N_2906,N_2494,N_1473);
and U2907 (N_2907,N_1015,N_1257);
or U2908 (N_2908,N_83,N_782);
or U2909 (N_2909,N_919,N_2294);
nand U2910 (N_2910,N_1534,N_411);
xnor U2911 (N_2911,N_826,N_2230);
nand U2912 (N_2912,N_147,N_1286);
or U2913 (N_2913,N_89,N_2176);
nor U2914 (N_2914,N_2271,N_1579);
nor U2915 (N_2915,N_1916,N_2435);
and U2916 (N_2916,N_982,N_904);
nor U2917 (N_2917,N_1451,N_151);
or U2918 (N_2918,N_1686,N_1819);
nand U2919 (N_2919,N_666,N_140);
or U2920 (N_2920,N_315,N_1524);
and U2921 (N_2921,N_1864,N_74);
and U2922 (N_2922,N_527,N_608);
nor U2923 (N_2923,N_1313,N_116);
or U2924 (N_2924,N_714,N_1134);
nor U2925 (N_2925,N_629,N_737);
or U2926 (N_2926,N_2177,N_801);
and U2927 (N_2927,N_1138,N_1170);
nand U2928 (N_2928,N_889,N_775);
nor U2929 (N_2929,N_2005,N_706);
nand U2930 (N_2930,N_255,N_376);
nor U2931 (N_2931,N_1263,N_1120);
nand U2932 (N_2932,N_1541,N_633);
nor U2933 (N_2933,N_607,N_1311);
or U2934 (N_2934,N_1841,N_254);
nor U2935 (N_2935,N_1229,N_13);
nand U2936 (N_2936,N_2439,N_131);
nand U2937 (N_2937,N_1975,N_1190);
or U2938 (N_2938,N_567,N_76);
and U2939 (N_2939,N_1474,N_1714);
nand U2940 (N_2940,N_858,N_1480);
or U2941 (N_2941,N_1648,N_2255);
and U2942 (N_2942,N_1554,N_1765);
or U2943 (N_2943,N_1643,N_645);
and U2944 (N_2944,N_190,N_1631);
and U2945 (N_2945,N_2371,N_1670);
or U2946 (N_2946,N_1019,N_2086);
nor U2947 (N_2947,N_2350,N_1824);
xor U2948 (N_2948,N_2419,N_195);
nor U2949 (N_2949,N_785,N_379);
nand U2950 (N_2950,N_2000,N_1012);
nand U2951 (N_2951,N_1688,N_1354);
or U2952 (N_2952,N_2218,N_1958);
nor U2953 (N_2953,N_726,N_204);
nand U2954 (N_2954,N_443,N_2468);
nor U2955 (N_2955,N_1395,N_935);
nand U2956 (N_2956,N_368,N_719);
nand U2957 (N_2957,N_1646,N_1284);
xnor U2958 (N_2958,N_665,N_1578);
and U2959 (N_2959,N_1611,N_2476);
nor U2960 (N_2960,N_2045,N_222);
and U2961 (N_2961,N_2180,N_2402);
and U2962 (N_2962,N_1146,N_1909);
nor U2963 (N_2963,N_786,N_2019);
nand U2964 (N_2964,N_2009,N_1588);
nor U2965 (N_2965,N_2219,N_1459);
nand U2966 (N_2966,N_2276,N_1667);
and U2967 (N_2967,N_1266,N_1269);
nor U2968 (N_2968,N_634,N_612);
and U2969 (N_2969,N_724,N_522);
or U2970 (N_2970,N_2452,N_1606);
nor U2971 (N_2971,N_939,N_1816);
or U2972 (N_2972,N_1743,N_435);
or U2973 (N_2973,N_1051,N_1895);
or U2974 (N_2974,N_1177,N_1660);
nor U2975 (N_2975,N_2024,N_2449);
and U2976 (N_2976,N_2337,N_2042);
and U2977 (N_2977,N_511,N_484);
or U2978 (N_2978,N_532,N_1568);
or U2979 (N_2979,N_1423,N_2023);
or U2980 (N_2980,N_2181,N_391);
and U2981 (N_2981,N_884,N_2233);
and U2982 (N_2982,N_940,N_1303);
nor U2983 (N_2983,N_1463,N_2342);
nand U2984 (N_2984,N_1100,N_1202);
and U2985 (N_2985,N_1394,N_2247);
nand U2986 (N_2986,N_1790,N_1057);
nand U2987 (N_2987,N_1927,N_184);
or U2988 (N_2988,N_1763,N_305);
and U2989 (N_2989,N_2293,N_1587);
nor U2990 (N_2990,N_2369,N_1174);
nand U2991 (N_2991,N_2097,N_1976);
or U2992 (N_2992,N_2287,N_2333);
nand U2993 (N_2993,N_23,N_1192);
nand U2994 (N_2994,N_1384,N_525);
nand U2995 (N_2995,N_891,N_1135);
or U2996 (N_2996,N_373,N_899);
or U2997 (N_2997,N_1884,N_1794);
or U2998 (N_2998,N_214,N_2149);
or U2999 (N_2999,N_239,N_2190);
nand U3000 (N_3000,N_1242,N_727);
and U3001 (N_3001,N_144,N_171);
or U3002 (N_3002,N_2472,N_2194);
and U3003 (N_3003,N_599,N_1090);
nand U3004 (N_3004,N_1840,N_446);
nor U3005 (N_3005,N_1008,N_1935);
or U3006 (N_3006,N_2443,N_1553);
nor U3007 (N_3007,N_231,N_793);
or U3008 (N_3008,N_2227,N_1435);
nor U3009 (N_3009,N_2201,N_1536);
nor U3010 (N_3010,N_1013,N_2063);
nor U3011 (N_3011,N_1328,N_521);
nor U3012 (N_3012,N_59,N_2215);
nor U3013 (N_3013,N_2074,N_1703);
or U3014 (N_3014,N_986,N_988);
nor U3015 (N_3015,N_656,N_182);
nand U3016 (N_3016,N_1148,N_457);
nand U3017 (N_3017,N_817,N_1542);
or U3018 (N_3018,N_603,N_1122);
nor U3019 (N_3019,N_1761,N_1846);
and U3020 (N_3020,N_1314,N_2366);
or U3021 (N_3021,N_2290,N_952);
nor U3022 (N_3022,N_1801,N_1635);
and U3023 (N_3023,N_1792,N_587);
and U3024 (N_3024,N_69,N_2329);
or U3025 (N_3025,N_1054,N_2134);
or U3026 (N_3026,N_1839,N_2249);
nand U3027 (N_3027,N_617,N_1736);
nand U3028 (N_3028,N_1332,N_2422);
nor U3029 (N_3029,N_408,N_1444);
nor U3030 (N_3030,N_1010,N_287);
or U3031 (N_3031,N_1035,N_1074);
xnor U3032 (N_3032,N_1738,N_1437);
nor U3033 (N_3033,N_1921,N_912);
nor U3034 (N_3034,N_461,N_2076);
nand U3035 (N_3035,N_1223,N_1386);
or U3036 (N_3036,N_998,N_936);
and U3037 (N_3037,N_55,N_2451);
or U3038 (N_3038,N_1275,N_781);
and U3039 (N_3039,N_1070,N_313);
nand U3040 (N_3040,N_1713,N_417);
or U3041 (N_3041,N_1751,N_1850);
and U3042 (N_3042,N_1295,N_636);
nand U3043 (N_3043,N_2041,N_581);
or U3044 (N_3044,N_1888,N_1589);
or U3045 (N_3045,N_1833,N_985);
and U3046 (N_3046,N_2116,N_1720);
xor U3047 (N_3047,N_455,N_1709);
and U3048 (N_3048,N_185,N_745);
nand U3049 (N_3049,N_606,N_963);
or U3050 (N_3050,N_1376,N_558);
nand U3051 (N_3051,N_390,N_1902);
nand U3052 (N_3052,N_931,N_822);
nor U3053 (N_3053,N_1402,N_20);
or U3054 (N_3054,N_1352,N_2251);
or U3055 (N_3055,N_380,N_2397);
nand U3056 (N_3056,N_827,N_614);
and U3057 (N_3057,N_1903,N_161);
nand U3058 (N_3058,N_464,N_622);
and U3059 (N_3059,N_803,N_1029);
or U3060 (N_3060,N_1331,N_1042);
nand U3061 (N_3061,N_894,N_689);
or U3062 (N_3062,N_1327,N_1344);
nor U3063 (N_3063,N_1662,N_646);
or U3064 (N_3064,N_486,N_642);
or U3065 (N_3065,N_1289,N_336);
nand U3066 (N_3066,N_653,N_311);
nor U3067 (N_3067,N_2221,N_1548);
and U3068 (N_3068,N_2483,N_1299);
xnor U3069 (N_3069,N_1838,N_2039);
nor U3070 (N_3070,N_2235,N_600);
nand U3071 (N_3071,N_1827,N_400);
nor U3072 (N_3072,N_1450,N_112);
and U3073 (N_3073,N_205,N_303);
nor U3074 (N_3074,N_1877,N_199);
or U3075 (N_3075,N_1021,N_1466);
and U3076 (N_3076,N_458,N_398);
or U3077 (N_3077,N_492,N_275);
and U3078 (N_3078,N_562,N_897);
nor U3079 (N_3079,N_572,N_2330);
nor U3080 (N_3080,N_668,N_1005);
or U3081 (N_3081,N_2263,N_2495);
nand U3082 (N_3082,N_342,N_394);
nor U3083 (N_3083,N_1270,N_1873);
nand U3084 (N_3084,N_1940,N_1981);
nor U3085 (N_3085,N_2359,N_441);
nor U3086 (N_3086,N_1102,N_1820);
nand U3087 (N_3087,N_836,N_1829);
or U3088 (N_3088,N_2054,N_1854);
or U3089 (N_3089,N_1504,N_658);
and U3090 (N_3090,N_1596,N_2077);
and U3091 (N_3091,N_377,N_2154);
and U3092 (N_3092,N_215,N_1793);
and U3093 (N_3093,N_1684,N_578);
nor U3094 (N_3094,N_56,N_1201);
nor U3095 (N_3095,N_1292,N_1001);
nor U3096 (N_3096,N_507,N_416);
and U3097 (N_3097,N_1954,N_752);
nor U3098 (N_3098,N_1796,N_920);
nand U3099 (N_3099,N_1946,N_756);
and U3100 (N_3100,N_2158,N_1397);
nor U3101 (N_3101,N_2376,N_1977);
and U3102 (N_3102,N_1566,N_1290);
nor U3103 (N_3103,N_165,N_1340);
nand U3104 (N_3104,N_2437,N_1601);
xnor U3105 (N_3105,N_2065,N_649);
nor U3106 (N_3106,N_217,N_1221);
nor U3107 (N_3107,N_2469,N_349);
nor U3108 (N_3108,N_833,N_1931);
nor U3109 (N_3109,N_903,N_329);
and U3110 (N_3110,N_2405,N_584);
and U3111 (N_3111,N_1237,N_1204);
or U3112 (N_3112,N_1356,N_1897);
or U3113 (N_3113,N_1681,N_2358);
and U3114 (N_3114,N_1956,N_684);
and U3115 (N_3115,N_41,N_338);
or U3116 (N_3116,N_477,N_207);
nand U3117 (N_3117,N_2217,N_1003);
nor U3118 (N_3118,N_1972,N_179);
nand U3119 (N_3119,N_2135,N_2324);
nand U3120 (N_3120,N_232,N_1990);
and U3121 (N_3121,N_152,N_552);
nor U3122 (N_3122,N_1272,N_1187);
or U3123 (N_3123,N_1253,N_509);
nor U3124 (N_3124,N_1624,N_1342);
nand U3125 (N_3125,N_2343,N_404);
nand U3126 (N_3126,N_1507,N_1343);
nand U3127 (N_3127,N_980,N_1082);
nand U3128 (N_3128,N_2004,N_970);
or U3129 (N_3129,N_2423,N_240);
nand U3130 (N_3130,N_1724,N_2232);
nor U3131 (N_3131,N_2001,N_1);
or U3132 (N_3132,N_639,N_80);
nand U3133 (N_3133,N_709,N_1942);
and U3134 (N_3134,N_1465,N_1260);
and U3135 (N_3135,N_1580,N_1866);
and U3136 (N_3136,N_924,N_1991);
nand U3137 (N_3137,N_2220,N_958);
nand U3138 (N_3138,N_30,N_2026);
nor U3139 (N_3139,N_2068,N_1960);
or U3140 (N_3140,N_1124,N_1609);
nor U3141 (N_3141,N_2356,N_1281);
and U3142 (N_3142,N_698,N_392);
and U3143 (N_3143,N_2126,N_2489);
nor U3144 (N_3144,N_286,N_778);
xnor U3145 (N_3145,N_1112,N_2275);
or U3146 (N_3146,N_605,N_1205);
and U3147 (N_3147,N_650,N_1164);
nor U3148 (N_3148,N_710,N_236);
and U3149 (N_3149,N_264,N_1438);
or U3150 (N_3150,N_388,N_1149);
or U3151 (N_3151,N_2011,N_1009);
and U3152 (N_3152,N_2394,N_238);
or U3153 (N_3153,N_260,N_2128);
and U3154 (N_3154,N_741,N_956);
xnor U3155 (N_3155,N_1349,N_1161);
and U3156 (N_3156,N_1044,N_2141);
and U3157 (N_3157,N_528,N_2033);
and U3158 (N_3158,N_70,N_1527);
nor U3159 (N_3159,N_98,N_1783);
and U3160 (N_3160,N_740,N_1178);
nand U3161 (N_3161,N_594,N_2345);
and U3162 (N_3162,N_1372,N_589);
or U3163 (N_3163,N_2210,N_2122);
and U3164 (N_3164,N_1073,N_2444);
or U3165 (N_3165,N_1680,N_2338);
xnor U3166 (N_3166,N_1348,N_1640);
nor U3167 (N_3167,N_1154,N_576);
nor U3168 (N_3168,N_1739,N_1682);
or U3169 (N_3169,N_223,N_625);
nand U3170 (N_3170,N_2044,N_2429);
or U3171 (N_3171,N_1099,N_1957);
nand U3172 (N_3172,N_1000,N_335);
and U3173 (N_3173,N_2094,N_1563);
xnor U3174 (N_3174,N_410,N_124);
xor U3175 (N_3175,N_969,N_1922);
nor U3176 (N_3176,N_2016,N_1722);
or U3177 (N_3177,N_1215,N_1594);
xor U3178 (N_3178,N_397,N_1855);
or U3179 (N_3179,N_1923,N_1407);
and U3180 (N_3180,N_1226,N_2301);
nand U3181 (N_3181,N_282,N_1457);
and U3182 (N_3182,N_1882,N_2252);
nand U3183 (N_3183,N_544,N_352);
nand U3184 (N_3184,N_3,N_1848);
nand U3185 (N_3185,N_575,N_1655);
or U3186 (N_3186,N_1470,N_1785);
nand U3187 (N_3187,N_172,N_237);
and U3188 (N_3188,N_569,N_34);
or U3189 (N_3189,N_604,N_1775);
or U3190 (N_3190,N_1683,N_758);
and U3191 (N_3191,N_777,N_85);
nand U3192 (N_3192,N_592,N_2118);
nor U3193 (N_3193,N_2470,N_122);
and U3194 (N_3194,N_2424,N_2467);
nand U3195 (N_3195,N_2090,N_753);
nor U3196 (N_3196,N_1077,N_1433);
or U3197 (N_3197,N_409,N_972);
xor U3198 (N_3198,N_1379,N_854);
or U3199 (N_3199,N_462,N_2071);
or U3200 (N_3200,N_2206,N_295);
nand U3201 (N_3201,N_1185,N_18);
or U3202 (N_3202,N_1690,N_1774);
and U3203 (N_3203,N_500,N_2328);
nor U3204 (N_3204,N_1424,N_1802);
and U3205 (N_3205,N_1959,N_2428);
and U3206 (N_3206,N_1211,N_857);
nor U3207 (N_3207,N_1881,N_1254);
nor U3208 (N_3208,N_787,N_911);
nand U3209 (N_3209,N_2034,N_557);
nor U3210 (N_3210,N_898,N_343);
and U3211 (N_3211,N_1821,N_2137);
nand U3212 (N_3212,N_751,N_1967);
nand U3213 (N_3213,N_2148,N_1166);
or U3214 (N_3214,N_384,N_2478);
nand U3215 (N_3215,N_620,N_590);
or U3216 (N_3216,N_837,N_2305);
xor U3217 (N_3217,N_743,N_281);
xor U3218 (N_3218,N_246,N_615);
nand U3219 (N_3219,N_1064,N_548);
or U3220 (N_3220,N_1503,N_1053);
nand U3221 (N_3221,N_2484,N_1419);
nand U3222 (N_3222,N_1830,N_1228);
nor U3223 (N_3223,N_29,N_1799);
xnor U3224 (N_3224,N_561,N_2225);
or U3225 (N_3225,N_333,N_1591);
and U3226 (N_3226,N_2340,N_143);
and U3227 (N_3227,N_2286,N_244);
or U3228 (N_3228,N_838,N_824);
or U3229 (N_3229,N_1391,N_220);
xor U3230 (N_3230,N_1153,N_2308);
nor U3231 (N_3231,N_1634,N_1213);
nor U3232 (N_3232,N_180,N_1125);
nand U3233 (N_3233,N_1345,N_1087);
and U3234 (N_3234,N_2139,N_1487);
nand U3235 (N_3235,N_2400,N_2205);
nor U3236 (N_3236,N_703,N_1039);
and U3237 (N_3237,N_42,N_846);
and U3238 (N_3238,N_1878,N_1426);
and U3239 (N_3239,N_835,N_566);
and U3240 (N_3240,N_1750,N_1298);
nand U3241 (N_3241,N_1194,N_1512);
or U3242 (N_3242,N_2465,N_1130);
and U3243 (N_3243,N_1224,N_921);
xor U3244 (N_3244,N_1377,N_583);
and U3245 (N_3245,N_8,N_1199);
or U3246 (N_3246,N_2153,N_2381);
nand U3247 (N_3247,N_2161,N_563);
nor U3248 (N_3248,N_292,N_289);
nand U3249 (N_3249,N_1564,N_2162);
nand U3250 (N_3250,N_1837,N_923);
and U3251 (N_3251,N_588,N_1297);
and U3252 (N_3252,N_821,N_1004);
or U3253 (N_3253,N_1443,N_768);
and U3254 (N_3254,N_1776,N_860);
nor U3255 (N_3255,N_677,N_1078);
nor U3256 (N_3256,N_110,N_914);
or U3257 (N_3257,N_1777,N_783);
nand U3258 (N_3258,N_537,N_880);
or U3259 (N_3259,N_1144,N_1891);
or U3260 (N_3260,N_1113,N_1502);
nor U3261 (N_3261,N_933,N_1066);
nor U3262 (N_3262,N_1460,N_818);
or U3263 (N_3263,N_2183,N_779);
nor U3264 (N_3264,N_1608,N_2430);
and U3265 (N_3265,N_2288,N_2228);
or U3266 (N_3266,N_1540,N_861);
nand U3267 (N_3267,N_2246,N_1143);
or U3268 (N_3268,N_1605,N_150);
or U3269 (N_3269,N_1262,N_1048);
or U3270 (N_3270,N_136,N_485);
nor U3271 (N_3271,N_873,N_2481);
nor U3272 (N_3272,N_1506,N_470);
nand U3273 (N_3273,N_2317,N_1461);
and U3274 (N_3274,N_159,N_702);
nand U3275 (N_3275,N_393,N_1358);
xor U3276 (N_3276,N_290,N_1844);
nand U3277 (N_3277,N_1002,N_879);
nand U3278 (N_3278,N_2237,N_2057);
or U3279 (N_3279,N_849,N_1404);
nor U3280 (N_3280,N_291,N_1151);
and U3281 (N_3281,N_1168,N_1023);
or U3282 (N_3282,N_1550,N_454);
nand U3283 (N_3283,N_1212,N_1971);
nor U3284 (N_3284,N_2080,N_2447);
and U3285 (N_3285,N_354,N_105);
nor U3286 (N_3286,N_2238,N_1560);
xor U3287 (N_3287,N_1639,N_467);
and U3288 (N_3288,N_1374,N_1740);
or U3289 (N_3289,N_832,N_1387);
or U3290 (N_3290,N_1773,N_2010);
nand U3291 (N_3291,N_2266,N_271);
nand U3292 (N_3292,N_1277,N_543);
or U3293 (N_3293,N_1337,N_1561);
nand U3294 (N_3294,N_2136,N_540);
nor U3295 (N_3295,N_1485,N_2061);
and U3296 (N_3296,N_1076,N_955);
or U3297 (N_3297,N_2456,N_2073);
nand U3298 (N_3298,N_1650,N_1963);
and U3299 (N_3299,N_1619,N_978);
and U3300 (N_3300,N_1953,N_1017);
nor U3301 (N_3301,N_1556,N_481);
nand U3302 (N_3302,N_1428,N_2089);
nor U3303 (N_3303,N_1390,N_705);
nor U3304 (N_3304,N_648,N_1583);
nand U3305 (N_3305,N_148,N_506);
and U3306 (N_3306,N_850,N_1951);
and U3307 (N_3307,N_1669,N_153);
nor U3308 (N_3308,N_501,N_991);
and U3309 (N_3309,N_2393,N_261);
and U3310 (N_3310,N_1814,N_2006);
nand U3311 (N_3311,N_1835,N_2213);
nand U3312 (N_3312,N_2281,N_1782);
or U3313 (N_3313,N_268,N_175);
nor U3314 (N_3314,N_631,N_418);
or U3315 (N_3315,N_1256,N_351);
nand U3316 (N_3316,N_1899,N_536);
nor U3317 (N_3317,N_399,N_267);
or U3318 (N_3318,N_1575,N_1985);
and U3319 (N_3319,N_611,N_1628);
nor U3320 (N_3320,N_1350,N_487);
and U3321 (N_3321,N_203,N_252);
nor U3322 (N_3322,N_31,N_32);
nand U3323 (N_3323,N_2163,N_62);
xor U3324 (N_3324,N_2152,N_1780);
or U3325 (N_3325,N_967,N_547);
nor U3326 (N_3326,N_2184,N_2459);
nor U3327 (N_3327,N_2315,N_2471);
or U3328 (N_3328,N_2387,N_807);
nand U3329 (N_3329,N_1861,N_1406);
nand U3330 (N_3330,N_2418,N_299);
and U3331 (N_3331,N_2283,N_597);
or U3332 (N_3332,N_499,N_1430);
nand U3333 (N_3333,N_1121,N_421);
or U3334 (N_3334,N_1493,N_52);
or U3335 (N_3335,N_1118,N_1208);
and U3336 (N_3336,N_845,N_1653);
nor U3337 (N_3337,N_2360,N_1479);
nand U3338 (N_3338,N_682,N_129);
nor U3339 (N_3339,N_2401,N_2037);
nand U3340 (N_3340,N_2406,N_627);
and U3341 (N_3341,N_1317,N_2466);
nand U3342 (N_3342,N_655,N_407);
nor U3343 (N_3343,N_176,N_913);
and U3344 (N_3344,N_526,N_942);
nand U3345 (N_3345,N_2370,N_1901);
or U3346 (N_3346,N_1856,N_174);
xnor U3347 (N_3347,N_1268,N_1943);
and U3348 (N_3348,N_1251,N_1939);
nor U3349 (N_3349,N_1965,N_1571);
nand U3350 (N_3350,N_2463,N_243);
and U3351 (N_3351,N_197,N_893);
and U3352 (N_3352,N_1338,N_2150);
nor U3353 (N_3353,N_1167,N_2407);
and U3354 (N_3354,N_1117,N_2121);
and U3355 (N_3355,N_2060,N_825);
nand U3356 (N_3356,N_1857,N_2182);
nand U3357 (N_3357,N_2078,N_1442);
nand U3358 (N_3358,N_618,N_1416);
and U3359 (N_3359,N_331,N_748);
nor U3360 (N_3360,N_619,N_385);
nand U3361 (N_3361,N_2321,N_2098);
or U3362 (N_3362,N_92,N_2166);
and U3363 (N_3363,N_609,N_88);
nor U3364 (N_3364,N_1061,N_1128);
nand U3365 (N_3365,N_37,N_1320);
nor U3366 (N_3366,N_4,N_990);
and U3367 (N_3367,N_471,N_1586);
and U3368 (N_3368,N_1103,N_966);
nand U3369 (N_3369,N_1086,N_119);
nor U3370 (N_3370,N_1432,N_2479);
nand U3371 (N_3371,N_332,N_1694);
or U3372 (N_3372,N_1543,N_1508);
or U3373 (N_3373,N_1689,N_1726);
nor U3374 (N_3374,N_46,N_957);
or U3375 (N_3375,N_780,N_16);
nand U3376 (N_3376,N_38,N_2007);
nor U3377 (N_3377,N_739,N_2487);
and U3378 (N_3378,N_178,N_169);
and U3379 (N_3379,N_320,N_886);
nor U3380 (N_3380,N_2365,N_1996);
xor U3381 (N_3381,N_819,N_1828);
and U3382 (N_3382,N_1757,N_39);
and U3383 (N_3383,N_2113,N_1758);
nand U3384 (N_3384,N_2214,N_1651);
nor U3385 (N_3385,N_1708,N_344);
nor U3386 (N_3386,N_1570,N_1659);
nand U3387 (N_3387,N_1329,N_2304);
and U3388 (N_3388,N_699,N_2279);
or U3389 (N_3389,N_623,N_881);
or U3390 (N_3390,N_355,N_1214);
or U3391 (N_3391,N_1274,N_318);
nor U3392 (N_3392,N_1913,N_1116);
nor U3393 (N_3393,N_1876,N_372);
nand U3394 (N_3394,N_1625,N_2391);
nand U3395 (N_3395,N_1498,N_93);
and U3396 (N_3396,N_810,N_47);
and U3397 (N_3397,N_276,N_1375);
nand U3398 (N_3398,N_1517,N_2273);
nand U3399 (N_3399,N_678,N_423);
nor U3400 (N_3400,N_2289,N_1746);
and U3401 (N_3401,N_1915,N_347);
nor U3402 (N_3402,N_1285,N_1865);
nand U3403 (N_3403,N_1364,N_510);
nand U3404 (N_3404,N_1526,N_242);
or U3405 (N_3405,N_1139,N_191);
or U3406 (N_3406,N_772,N_538);
nand U3407 (N_3407,N_2048,N_2485);
or U3408 (N_3408,N_304,N_1363);
nor U3409 (N_3409,N_1456,N_1545);
or U3410 (N_3410,N_1687,N_953);
nand U3411 (N_3411,N_917,N_137);
and U3412 (N_3412,N_1730,N_2260);
nor U3413 (N_3413,N_1823,N_2421);
nand U3414 (N_3414,N_910,N_1335);
nor U3415 (N_3415,N_1084,N_2224);
nand U3416 (N_3416,N_517,N_683);
nand U3417 (N_3417,N_1803,N_950);
and U3418 (N_3418,N_14,N_497);
or U3419 (N_3419,N_1101,N_784);
nand U3420 (N_3420,N_520,N_800);
nor U3421 (N_3421,N_104,N_1179);
and U3422 (N_3422,N_2386,N_1373);
nand U3423 (N_3423,N_908,N_364);
nor U3424 (N_3424,N_1973,N_381);
nand U3425 (N_3425,N_2269,N_2355);
and U3426 (N_3426,N_1056,N_831);
nand U3427 (N_3427,N_586,N_2363);
and U3428 (N_3428,N_1742,N_2256);
nand U3429 (N_3429,N_2300,N_2282);
and U3430 (N_3430,N_256,N_2244);
or U3431 (N_3431,N_954,N_1357);
nand U3432 (N_3432,N_663,N_1998);
nor U3433 (N_3433,N_386,N_2207);
and U3434 (N_3434,N_2203,N_2309);
nand U3435 (N_3435,N_2229,N_2242);
and U3436 (N_3436,N_2311,N_571);
and U3437 (N_3437,N_145,N_1282);
and U3438 (N_3438,N_2200,N_1710);
and U3439 (N_3439,N_1367,N_498);
nand U3440 (N_3440,N_213,N_2223);
and U3441 (N_3441,N_2453,N_2274);
or U3442 (N_3442,N_2258,N_2196);
nor U3443 (N_3443,N_1152,N_1645);
nor U3444 (N_3444,N_732,N_1735);
and U3445 (N_3445,N_2117,N_17);
nand U3446 (N_3446,N_515,N_949);
or U3447 (N_3447,N_1250,N_2462);
or U3448 (N_3448,N_1222,N_1944);
or U3449 (N_3449,N_1500,N_326);
or U3450 (N_3450,N_43,N_81);
nand U3451 (N_3451,N_556,N_210);
nor U3452 (N_3452,N_2127,N_1644);
nand U3453 (N_3453,N_2120,N_1938);
nor U3454 (N_3454,N_1336,N_2146);
and U3455 (N_3455,N_843,N_637);
or U3456 (N_3456,N_513,N_1590);
and U3457 (N_3457,N_1315,N_2248);
nor U3458 (N_3458,N_1193,N_0);
or U3459 (N_3459,N_2108,N_164);
or U3460 (N_3460,N_200,N_221);
nor U3461 (N_3461,N_2035,N_100);
nand U3462 (N_3462,N_1567,N_432);
and U3463 (N_3463,N_2280,N_1188);
nand U3464 (N_3464,N_1847,N_2030);
nor U3465 (N_3465,N_1071,N_1381);
nor U3466 (N_3466,N_228,N_1537);
nor U3467 (N_3467,N_2245,N_330);
nand U3468 (N_3468,N_2384,N_1131);
or U3469 (N_3469,N_1408,N_1767);
nand U3470 (N_3470,N_35,N_1691);
nand U3471 (N_3471,N_856,N_1301);
nor U3472 (N_3472,N_193,N_815);
and U3473 (N_3473,N_109,N_1436);
nand U3474 (N_3474,N_1509,N_755);
nand U3475 (N_3475,N_2084,N_1414);
or U3476 (N_3476,N_1671,N_1497);
or U3477 (N_3477,N_878,N_183);
and U3478 (N_3478,N_2346,N_1870);
nand U3479 (N_3479,N_1514,N_25);
nand U3480 (N_3480,N_1786,N_593);
nor U3481 (N_3481,N_2380,N_2168);
nor U3482 (N_3482,N_2092,N_1055);
or U3483 (N_3483,N_235,N_1382);
and U3484 (N_3484,N_1216,N_1908);
and U3485 (N_3485,N_1267,N_759);
nand U3486 (N_3486,N_1741,N_2008);
or U3487 (N_3487,N_1050,N_2410);
or U3488 (N_3488,N_91,N_1727);
nor U3489 (N_3489,N_1453,N_539);
and U3490 (N_3490,N_717,N_307);
nand U3491 (N_3491,N_359,N_482);
nand U3492 (N_3492,N_896,N_1175);
or U3493 (N_3493,N_704,N_2474);
or U3494 (N_3494,N_1614,N_101);
xnor U3495 (N_3495,N_1043,N_1346);
or U3496 (N_3496,N_1478,N_2292);
or U3497 (N_3497,N_1203,N_12);
nand U3498 (N_3498,N_667,N_1898);
or U3499 (N_3499,N_1538,N_120);
nor U3500 (N_3500,N_253,N_350);
nand U3501 (N_3501,N_156,N_937);
nand U3502 (N_3502,N_2375,N_370);
or U3503 (N_3503,N_725,N_2262);
nand U3504 (N_3504,N_1183,N_1852);
nor U3505 (N_3505,N_701,N_298);
and U3506 (N_3506,N_2313,N_2446);
nand U3507 (N_3507,N_791,N_334);
and U3508 (N_3508,N_712,N_2129);
nand U3509 (N_3509,N_1858,N_1110);
nor U3510 (N_3510,N_1555,N_2047);
nor U3511 (N_3511,N_453,N_1037);
or U3512 (N_3512,N_2458,N_1007);
nor U3513 (N_3513,N_2209,N_1831);
or U3514 (N_3514,N_374,N_474);
and U3515 (N_3515,N_60,N_2372);
nand U3516 (N_3516,N_1040,N_1744);
nand U3517 (N_3517,N_2013,N_2438);
or U3518 (N_3518,N_1525,N_944);
or U3519 (N_3519,N_2110,N_2130);
and U3520 (N_3520,N_2072,N_113);
nand U3521 (N_3521,N_2433,N_2413);
or U3522 (N_3522,N_64,N_2131);
nor U3523 (N_3523,N_700,N_1970);
nor U3524 (N_3524,N_1531,N_2239);
nand U3525 (N_3525,N_723,N_975);
nor U3526 (N_3526,N_269,N_2102);
nand U3527 (N_3527,N_1842,N_1325);
or U3528 (N_3528,N_610,N_1353);
and U3529 (N_3529,N_1734,N_928);
nand U3530 (N_3530,N_378,N_1789);
or U3531 (N_3531,N_549,N_1469);
nor U3532 (N_3532,N_2298,N_1934);
or U3533 (N_3533,N_1032,N_1928);
or U3534 (N_3534,N_419,N_672);
nand U3535 (N_3535,N_1862,N_1705);
or U3536 (N_3536,N_1808,N_1049);
and U3537 (N_3537,N_2492,N_19);
nand U3538 (N_3538,N_1255,N_2028);
and U3539 (N_3539,N_67,N_697);
xor U3540 (N_3540,N_1894,N_211);
nand U3541 (N_3541,N_1510,N_964);
and U3542 (N_3542,N_1622,N_1291);
and U3543 (N_3543,N_999,N_208);
nand U3544 (N_3544,N_948,N_300);
or U3545 (N_3545,N_1483,N_79);
nand U3546 (N_3546,N_296,N_1279);
nand U3547 (N_3547,N_1893,N_1081);
nand U3548 (N_3548,N_553,N_1672);
or U3549 (N_3549,N_1068,N_1371);
nand U3550 (N_3550,N_1316,N_869);
and U3551 (N_3551,N_97,N_2105);
nand U3552 (N_3552,N_1016,N_1549);
nand U3553 (N_3553,N_2151,N_2490);
or U3554 (N_3554,N_997,N_73);
and U3555 (N_3555,N_1986,N_1417);
nor U3556 (N_3556,N_96,N_90);
nand U3557 (N_3557,N_505,N_1264);
nand U3558 (N_3558,N_1872,N_1245);
or U3559 (N_3559,N_283,N_494);
and U3560 (N_3560,N_713,N_1092);
and U3561 (N_3561,N_814,N_1729);
nand U3562 (N_3562,N_971,N_132);
and U3563 (N_3563,N_890,N_1515);
nand U3564 (N_3564,N_582,N_227);
and U3565 (N_3565,N_1768,N_1999);
nor U3566 (N_3566,N_514,N_2432);
or U3567 (N_3567,N_1704,N_160);
and U3568 (N_3568,N_45,N_1033);
and U3569 (N_3569,N_696,N_6);
or U3570 (N_3570,N_2425,N_591);
and U3571 (N_3571,N_918,N_356);
or U3572 (N_3572,N_1593,N_1997);
nor U3573 (N_3573,N_641,N_2198);
or U3574 (N_3574,N_1920,N_823);
and U3575 (N_3575,N_1817,N_2268);
nor U3576 (N_3576,N_466,N_192);
nor U3577 (N_3577,N_984,N_1696);
xnor U3578 (N_3578,N_1014,N_1259);
nand U3579 (N_3579,N_852,N_1661);
nor U3580 (N_3580,N_194,N_808);
or U3581 (N_3581,N_1380,N_1577);
nand U3582 (N_3582,N_551,N_1173);
nand U3583 (N_3583,N_2066,N_2014);
and U3584 (N_3584,N_279,N_875);
nand U3585 (N_3585,N_1883,N_601);
or U3586 (N_3586,N_1994,N_1341);
nor U3587 (N_3587,N_1926,N_545);
xor U3588 (N_3588,N_722,N_444);
nand U3589 (N_3589,N_1241,N_1176);
or U3590 (N_3590,N_1431,N_2368);
and U3591 (N_3591,N_2303,N_170);
or U3592 (N_3592,N_1230,N_1252);
nor U3593 (N_3593,N_922,N_1207);
nor U3594 (N_3594,N_1604,N_2291);
nor U3595 (N_3595,N_2460,N_353);
nand U3596 (N_3596,N_1105,N_2157);
and U3597 (N_3597,N_1760,N_796);
or U3598 (N_3598,N_1361,N_490);
nand U3599 (N_3599,N_2051,N_1613);
and U3600 (N_3600,N_981,N_1287);
or U3601 (N_3601,N_2493,N_1142);
xnor U3602 (N_3602,N_542,N_434);
nor U3603 (N_3603,N_616,N_1621);
and U3604 (N_3604,N_2012,N_734);
and U3605 (N_3605,N_2389,N_1933);
and U3606 (N_3606,N_930,N_40);
or U3607 (N_3607,N_1544,N_1409);
nand U3608 (N_3608,N_872,N_483);
and U3609 (N_3609,N_463,N_1753);
or U3610 (N_3610,N_841,N_1421);
or U3611 (N_3611,N_1911,N_257);
nor U3612 (N_3612,N_245,N_1779);
and U3613 (N_3613,N_1238,N_436);
or U3614 (N_3614,N_1616,N_960);
nand U3615 (N_3615,N_1890,N_2179);
nand U3616 (N_3616,N_2243,N_1900);
and U3617 (N_3617,N_771,N_871);
nor U3618 (N_3618,N_2144,N_1885);
nand U3619 (N_3619,N_413,N_673);
nand U3620 (N_3620,N_773,N_925);
nor U3621 (N_3621,N_686,N_127);
or U3622 (N_3622,N_2,N_1649);
nand U3623 (N_3623,N_2354,N_297);
and U3624 (N_3624,N_1647,N_2027);
and U3625 (N_3625,N_1030,N_1476);
nor U3626 (N_3626,N_695,N_365);
nor U3627 (N_3627,N_1978,N_472);
nor U3628 (N_3628,N_439,N_987);
nand U3629 (N_3629,N_1535,N_1950);
nor U3630 (N_3630,N_2448,N_1025);
and U3631 (N_3631,N_1449,N_2412);
xnor U3632 (N_3632,N_1925,N_1157);
nand U3633 (N_3633,N_95,N_480);
and U3634 (N_3634,N_2332,N_1519);
xor U3635 (N_3635,N_1679,N_2119);
or U3636 (N_3636,N_640,N_1573);
nor U3637 (N_3637,N_1968,N_451);
and U3638 (N_3638,N_2499,N_130);
nor U3639 (N_3639,N_2398,N_2211);
or U3640 (N_3640,N_1889,N_1521);
or U3641 (N_3641,N_579,N_864);
or U3642 (N_3642,N_529,N_1772);
nor U3643 (N_3643,N_1058,N_1038);
or U3644 (N_3644,N_314,N_2064);
and U3645 (N_3645,N_126,N_1107);
xnor U3646 (N_3646,N_54,N_63);
or U3647 (N_3647,N_94,N_114);
nand U3648 (N_3648,N_87,N_2392);
nand U3649 (N_3649,N_708,N_1706);
nand U3650 (N_3650,N_1969,N_962);
nand U3651 (N_3651,N_1471,N_750);
or U3652 (N_3652,N_1675,N_493);
nand U3653 (N_3653,N_1863,N_671);
nand U3654 (N_3654,N_844,N_2165);
or U3655 (N_3655,N_736,N_2431);
nand U3656 (N_3656,N_1413,N_1309);
xnor U3657 (N_3657,N_310,N_774);
and U3658 (N_3658,N_853,N_142);
and U3659 (N_3659,N_1701,N_1697);
nor U3660 (N_3660,N_685,N_2103);
nor U3661 (N_3661,N_2441,N_2351);
or U3662 (N_3662,N_847,N_2341);
nor U3663 (N_3663,N_154,N_1160);
nor U3664 (N_3664,N_2234,N_1756);
or U3665 (N_3665,N_906,N_1818);
and U3666 (N_3666,N_71,N_1718);
and U3667 (N_3667,N_664,N_189);
nand U3668 (N_3668,N_1302,N_48);
and U3669 (N_3669,N_1983,N_28);
and U3670 (N_3670,N_1867,N_460);
nand U3671 (N_3671,N_2454,N_2497);
and U3672 (N_3672,N_401,N_907);
and U3673 (N_3673,N_1488,N_248);
and U3674 (N_3674,N_2362,N_428);
nor U3675 (N_3675,N_577,N_976);
and U3676 (N_3676,N_1448,N_1258);
or U3677 (N_3677,N_2046,N_518);
and U3678 (N_3678,N_139,N_888);
xnor U3679 (N_3679,N_1452,N_1516);
and U3680 (N_3680,N_2062,N_15);
or U3681 (N_3681,N_613,N_788);
and U3682 (N_3682,N_1698,N_1467);
and U3683 (N_3683,N_1106,N_1813);
and U3684 (N_3684,N_1874,N_1552);
xnor U3685 (N_3685,N_1974,N_1798);
and U3686 (N_3686,N_1602,N_848);
nand U3687 (N_3687,N_1494,N_1612);
and U3688 (N_3688,N_2296,N_1638);
or U3689 (N_3689,N_902,N_1308);
and U3690 (N_3690,N_1326,N_2112);
nand U3691 (N_3691,N_426,N_565);
nand U3692 (N_3692,N_2138,N_2025);
and U3693 (N_3693,N_797,N_1234);
and U3694 (N_3694,N_2461,N_2264);
nor U3695 (N_3695,N_1518,N_720);
nand U3696 (N_3696,N_1137,N_362);
nor U3697 (N_3697,N_250,N_2133);
or U3698 (N_3698,N_1333,N_1565);
nor U3699 (N_3699,N_86,N_2020);
or U3700 (N_3700,N_805,N_1770);
nor U3701 (N_3701,N_1123,N_638);
or U3702 (N_3702,N_2491,N_2344);
and U3703 (N_3703,N_1547,N_502);
and U3704 (N_3704,N_2327,N_715);
or U3705 (N_3705,N_452,N_1657);
nand U3706 (N_3706,N_2496,N_2427);
nand U3707 (N_3707,N_657,N_1749);
nor U3708 (N_3708,N_660,N_1581);
or U3709 (N_3709,N_938,N_2187);
and U3710 (N_3710,N_1098,N_865);
nand U3711 (N_3711,N_1737,N_2319);
nor U3712 (N_3712,N_1859,N_2018);
or U3713 (N_3713,N_2488,N_868);
nand U3714 (N_3714,N_2396,N_234);
nor U3715 (N_3715,N_1323,N_68);
nor U3716 (N_3716,N_1822,N_445);
nor U3717 (N_3717,N_1220,N_2477);
nand U3718 (N_3718,N_1800,N_1811);
nand U3719 (N_3719,N_2142,N_1319);
and U3720 (N_3720,N_155,N_1468);
nand U3721 (N_3721,N_1186,N_293);
and U3722 (N_3722,N_2434,N_1362);
and U3723 (N_3723,N_1964,N_1321);
or U3724 (N_3724,N_905,N_102);
nor U3725 (N_3725,N_2058,N_1246);
nand U3726 (N_3726,N_2261,N_560);
and U3727 (N_3727,N_2408,N_2083);
nand U3728 (N_3728,N_892,N_1712);
and U3729 (N_3729,N_135,N_916);
nand U3730 (N_3730,N_2323,N_2178);
nand U3731 (N_3731,N_348,N_1041);
or U3732 (N_3732,N_442,N_2031);
nor U3733 (N_3733,N_1191,N_1832);
nor U3734 (N_3734,N_2236,N_1764);
nor U3735 (N_3735,N_504,N_1458);
and U3736 (N_3736,N_196,N_1108);
nor U3737 (N_3737,N_1711,N_1141);
nor U3738 (N_3738,N_1522,N_106);
and U3739 (N_3739,N_5,N_2143);
or U3740 (N_3740,N_535,N_274);
and U3741 (N_3741,N_2169,N_1232);
nand U3742 (N_3742,N_1150,N_1305);
nor U3743 (N_3743,N_438,N_1392);
nand U3744 (N_3744,N_202,N_340);
nor U3745 (N_3745,N_694,N_1851);
or U3746 (N_3746,N_951,N_2226);
nand U3747 (N_3747,N_1630,N_1189);
nor U3748 (N_3748,N_262,N_277);
and U3749 (N_3749,N_2125,N_1069);
or U3750 (N_3750,N_1514,N_1101);
nor U3751 (N_3751,N_502,N_743);
nand U3752 (N_3752,N_503,N_545);
nand U3753 (N_3753,N_2056,N_377);
and U3754 (N_3754,N_1391,N_2463);
nand U3755 (N_3755,N_979,N_42);
or U3756 (N_3756,N_1836,N_4);
nor U3757 (N_3757,N_225,N_858);
or U3758 (N_3758,N_924,N_2113);
and U3759 (N_3759,N_1363,N_111);
or U3760 (N_3760,N_1287,N_1554);
nor U3761 (N_3761,N_115,N_1252);
and U3762 (N_3762,N_1599,N_1216);
and U3763 (N_3763,N_1832,N_2240);
and U3764 (N_3764,N_902,N_1903);
nand U3765 (N_3765,N_126,N_63);
nor U3766 (N_3766,N_2012,N_64);
or U3767 (N_3767,N_13,N_711);
nand U3768 (N_3768,N_1392,N_2203);
nand U3769 (N_3769,N_1645,N_1193);
and U3770 (N_3770,N_1870,N_403);
or U3771 (N_3771,N_2339,N_1329);
nand U3772 (N_3772,N_1543,N_861);
and U3773 (N_3773,N_709,N_2384);
nor U3774 (N_3774,N_953,N_180);
and U3775 (N_3775,N_143,N_1131);
and U3776 (N_3776,N_1299,N_2412);
nor U3777 (N_3777,N_635,N_2157);
and U3778 (N_3778,N_2498,N_258);
nand U3779 (N_3779,N_687,N_810);
and U3780 (N_3780,N_1194,N_143);
nand U3781 (N_3781,N_196,N_966);
or U3782 (N_3782,N_1937,N_819);
or U3783 (N_3783,N_867,N_1864);
and U3784 (N_3784,N_1632,N_187);
nor U3785 (N_3785,N_1187,N_1851);
and U3786 (N_3786,N_2441,N_1962);
and U3787 (N_3787,N_1798,N_116);
nand U3788 (N_3788,N_442,N_2374);
and U3789 (N_3789,N_2297,N_1623);
or U3790 (N_3790,N_2470,N_2322);
nor U3791 (N_3791,N_1394,N_681);
nor U3792 (N_3792,N_1314,N_556);
and U3793 (N_3793,N_1409,N_2124);
and U3794 (N_3794,N_1504,N_2303);
and U3795 (N_3795,N_1401,N_310);
or U3796 (N_3796,N_1128,N_1638);
xnor U3797 (N_3797,N_1146,N_2176);
and U3798 (N_3798,N_488,N_2455);
nor U3799 (N_3799,N_1474,N_1077);
or U3800 (N_3800,N_2027,N_168);
and U3801 (N_3801,N_200,N_1983);
nand U3802 (N_3802,N_1680,N_1487);
and U3803 (N_3803,N_1952,N_99);
or U3804 (N_3804,N_66,N_2046);
and U3805 (N_3805,N_182,N_412);
nor U3806 (N_3806,N_891,N_1694);
or U3807 (N_3807,N_680,N_924);
or U3808 (N_3808,N_1971,N_1602);
or U3809 (N_3809,N_1126,N_1597);
and U3810 (N_3810,N_1796,N_848);
nand U3811 (N_3811,N_628,N_37);
nor U3812 (N_3812,N_2120,N_1024);
nor U3813 (N_3813,N_601,N_483);
nor U3814 (N_3814,N_2186,N_1928);
nand U3815 (N_3815,N_1227,N_1725);
or U3816 (N_3816,N_1339,N_740);
and U3817 (N_3817,N_691,N_550);
nand U3818 (N_3818,N_1639,N_229);
xor U3819 (N_3819,N_1116,N_1080);
and U3820 (N_3820,N_2085,N_183);
and U3821 (N_3821,N_2374,N_800);
nand U3822 (N_3822,N_1891,N_1734);
nor U3823 (N_3823,N_2316,N_2123);
nand U3824 (N_3824,N_337,N_2427);
nand U3825 (N_3825,N_938,N_2447);
xor U3826 (N_3826,N_2126,N_2294);
nor U3827 (N_3827,N_837,N_1511);
and U3828 (N_3828,N_1920,N_898);
or U3829 (N_3829,N_1404,N_415);
or U3830 (N_3830,N_883,N_1888);
nor U3831 (N_3831,N_930,N_1157);
nor U3832 (N_3832,N_538,N_1799);
nor U3833 (N_3833,N_110,N_1195);
nand U3834 (N_3834,N_1514,N_427);
nand U3835 (N_3835,N_737,N_589);
or U3836 (N_3836,N_1638,N_1578);
nor U3837 (N_3837,N_164,N_274);
nand U3838 (N_3838,N_2323,N_605);
nand U3839 (N_3839,N_56,N_462);
nor U3840 (N_3840,N_601,N_2053);
nor U3841 (N_3841,N_894,N_577);
xnor U3842 (N_3842,N_1573,N_769);
nor U3843 (N_3843,N_780,N_71);
nor U3844 (N_3844,N_1996,N_2081);
nor U3845 (N_3845,N_1002,N_1260);
nor U3846 (N_3846,N_793,N_2474);
nand U3847 (N_3847,N_1919,N_80);
nor U3848 (N_3848,N_1104,N_990);
and U3849 (N_3849,N_950,N_1207);
or U3850 (N_3850,N_1679,N_930);
xnor U3851 (N_3851,N_2430,N_972);
nand U3852 (N_3852,N_1720,N_360);
or U3853 (N_3853,N_2206,N_1834);
and U3854 (N_3854,N_2484,N_880);
nor U3855 (N_3855,N_95,N_270);
and U3856 (N_3856,N_1338,N_2126);
nand U3857 (N_3857,N_200,N_2081);
or U3858 (N_3858,N_391,N_1902);
nor U3859 (N_3859,N_1572,N_1215);
nor U3860 (N_3860,N_2456,N_833);
nor U3861 (N_3861,N_1912,N_1355);
or U3862 (N_3862,N_1704,N_2379);
and U3863 (N_3863,N_1698,N_1307);
nand U3864 (N_3864,N_1274,N_919);
nand U3865 (N_3865,N_941,N_267);
or U3866 (N_3866,N_571,N_2410);
nor U3867 (N_3867,N_1059,N_2208);
nand U3868 (N_3868,N_741,N_332);
nand U3869 (N_3869,N_1478,N_90);
and U3870 (N_3870,N_2479,N_340);
or U3871 (N_3871,N_936,N_720);
nand U3872 (N_3872,N_1262,N_2057);
nor U3873 (N_3873,N_2239,N_2002);
nand U3874 (N_3874,N_1924,N_336);
or U3875 (N_3875,N_2231,N_320);
and U3876 (N_3876,N_1030,N_397);
or U3877 (N_3877,N_871,N_2085);
or U3878 (N_3878,N_122,N_745);
or U3879 (N_3879,N_1120,N_217);
and U3880 (N_3880,N_2499,N_1864);
or U3881 (N_3881,N_1335,N_1197);
and U3882 (N_3882,N_801,N_1602);
nand U3883 (N_3883,N_1920,N_563);
and U3884 (N_3884,N_2398,N_490);
nor U3885 (N_3885,N_8,N_1336);
nand U3886 (N_3886,N_545,N_356);
and U3887 (N_3887,N_374,N_916);
nor U3888 (N_3888,N_1027,N_2262);
nand U3889 (N_3889,N_1055,N_721);
xor U3890 (N_3890,N_1647,N_2298);
nand U3891 (N_3891,N_2040,N_165);
and U3892 (N_3892,N_1880,N_1193);
nor U3893 (N_3893,N_800,N_2248);
nor U3894 (N_3894,N_1385,N_978);
or U3895 (N_3895,N_266,N_686);
nor U3896 (N_3896,N_1805,N_8);
and U3897 (N_3897,N_518,N_42);
nor U3898 (N_3898,N_695,N_822);
or U3899 (N_3899,N_817,N_2475);
nor U3900 (N_3900,N_1860,N_597);
or U3901 (N_3901,N_1627,N_92);
nor U3902 (N_3902,N_1977,N_1425);
nand U3903 (N_3903,N_1023,N_610);
and U3904 (N_3904,N_44,N_2062);
nand U3905 (N_3905,N_1646,N_1225);
and U3906 (N_3906,N_398,N_1346);
nand U3907 (N_3907,N_1192,N_1660);
and U3908 (N_3908,N_1665,N_1272);
or U3909 (N_3909,N_1960,N_2105);
nand U3910 (N_3910,N_1275,N_190);
nor U3911 (N_3911,N_1248,N_2156);
and U3912 (N_3912,N_1302,N_835);
or U3913 (N_3913,N_674,N_2437);
nor U3914 (N_3914,N_19,N_1485);
nand U3915 (N_3915,N_1297,N_2077);
nand U3916 (N_3916,N_2008,N_1095);
and U3917 (N_3917,N_1617,N_1767);
nor U3918 (N_3918,N_1151,N_2391);
and U3919 (N_3919,N_1585,N_256);
and U3920 (N_3920,N_2051,N_2497);
or U3921 (N_3921,N_1726,N_1906);
and U3922 (N_3922,N_1617,N_573);
nor U3923 (N_3923,N_980,N_2443);
or U3924 (N_3924,N_241,N_2223);
nand U3925 (N_3925,N_1459,N_607);
nand U3926 (N_3926,N_2286,N_771);
and U3927 (N_3927,N_378,N_665);
nor U3928 (N_3928,N_1164,N_1432);
nand U3929 (N_3929,N_1032,N_1348);
or U3930 (N_3930,N_2005,N_1241);
or U3931 (N_3931,N_2451,N_285);
or U3932 (N_3932,N_638,N_49);
nor U3933 (N_3933,N_448,N_621);
nor U3934 (N_3934,N_1413,N_943);
nor U3935 (N_3935,N_1166,N_929);
and U3936 (N_3936,N_1083,N_1141);
or U3937 (N_3937,N_963,N_447);
nand U3938 (N_3938,N_759,N_746);
and U3939 (N_3939,N_1487,N_1109);
nand U3940 (N_3940,N_1188,N_636);
or U3941 (N_3941,N_117,N_1876);
nand U3942 (N_3942,N_2400,N_1645);
or U3943 (N_3943,N_613,N_1721);
nor U3944 (N_3944,N_455,N_408);
or U3945 (N_3945,N_1885,N_1181);
and U3946 (N_3946,N_1960,N_2225);
xnor U3947 (N_3947,N_699,N_1679);
nand U3948 (N_3948,N_86,N_2463);
nand U3949 (N_3949,N_1784,N_686);
and U3950 (N_3950,N_1218,N_1929);
or U3951 (N_3951,N_2442,N_1821);
nor U3952 (N_3952,N_756,N_1445);
and U3953 (N_3953,N_2134,N_465);
or U3954 (N_3954,N_2166,N_397);
nor U3955 (N_3955,N_2183,N_2040);
nor U3956 (N_3956,N_1892,N_1086);
nand U3957 (N_3957,N_18,N_686);
and U3958 (N_3958,N_244,N_131);
or U3959 (N_3959,N_815,N_1532);
nor U3960 (N_3960,N_1877,N_499);
nor U3961 (N_3961,N_1507,N_978);
and U3962 (N_3962,N_1352,N_1049);
nand U3963 (N_3963,N_2169,N_447);
and U3964 (N_3964,N_2277,N_594);
nand U3965 (N_3965,N_2435,N_352);
or U3966 (N_3966,N_5,N_2242);
and U3967 (N_3967,N_1039,N_919);
and U3968 (N_3968,N_2073,N_673);
nand U3969 (N_3969,N_1700,N_1304);
and U3970 (N_3970,N_1539,N_1514);
nand U3971 (N_3971,N_2037,N_2087);
nand U3972 (N_3972,N_450,N_367);
nand U3973 (N_3973,N_901,N_25);
nand U3974 (N_3974,N_1732,N_283);
nand U3975 (N_3975,N_1320,N_2158);
and U3976 (N_3976,N_658,N_1434);
or U3977 (N_3977,N_2104,N_2306);
nor U3978 (N_3978,N_1224,N_356);
and U3979 (N_3979,N_2334,N_827);
nor U3980 (N_3980,N_1742,N_554);
and U3981 (N_3981,N_1225,N_2178);
or U3982 (N_3982,N_297,N_620);
nor U3983 (N_3983,N_1848,N_2418);
or U3984 (N_3984,N_1797,N_61);
and U3985 (N_3985,N_319,N_1400);
nor U3986 (N_3986,N_895,N_1019);
or U3987 (N_3987,N_1594,N_1114);
and U3988 (N_3988,N_1525,N_1051);
or U3989 (N_3989,N_2338,N_1844);
nand U3990 (N_3990,N_2469,N_1513);
nand U3991 (N_3991,N_1089,N_1696);
and U3992 (N_3992,N_2474,N_754);
and U3993 (N_3993,N_1391,N_2335);
nand U3994 (N_3994,N_2404,N_360);
nand U3995 (N_3995,N_352,N_2367);
and U3996 (N_3996,N_836,N_178);
nand U3997 (N_3997,N_2111,N_1142);
and U3998 (N_3998,N_1531,N_1355);
and U3999 (N_3999,N_15,N_652);
and U4000 (N_4000,N_542,N_1369);
or U4001 (N_4001,N_1363,N_2367);
nand U4002 (N_4002,N_1353,N_1520);
or U4003 (N_4003,N_1428,N_1737);
or U4004 (N_4004,N_734,N_1453);
nor U4005 (N_4005,N_1901,N_1191);
nor U4006 (N_4006,N_130,N_126);
or U4007 (N_4007,N_1518,N_1678);
and U4008 (N_4008,N_1718,N_1673);
or U4009 (N_4009,N_384,N_1251);
nand U4010 (N_4010,N_1222,N_865);
and U4011 (N_4011,N_1541,N_1202);
nor U4012 (N_4012,N_148,N_1901);
and U4013 (N_4013,N_1295,N_1928);
nor U4014 (N_4014,N_184,N_374);
and U4015 (N_4015,N_1193,N_920);
nor U4016 (N_4016,N_1489,N_1717);
nor U4017 (N_4017,N_1984,N_1076);
nand U4018 (N_4018,N_1919,N_2337);
nor U4019 (N_4019,N_58,N_923);
nand U4020 (N_4020,N_2174,N_1088);
or U4021 (N_4021,N_2127,N_1336);
and U4022 (N_4022,N_1169,N_2328);
and U4023 (N_4023,N_1776,N_2056);
nand U4024 (N_4024,N_1038,N_1574);
nand U4025 (N_4025,N_2018,N_1335);
or U4026 (N_4026,N_1271,N_1408);
nor U4027 (N_4027,N_2008,N_1369);
nor U4028 (N_4028,N_677,N_1759);
or U4029 (N_4029,N_509,N_1439);
or U4030 (N_4030,N_153,N_101);
or U4031 (N_4031,N_402,N_852);
and U4032 (N_4032,N_773,N_175);
or U4033 (N_4033,N_827,N_252);
nor U4034 (N_4034,N_1513,N_1600);
nor U4035 (N_4035,N_1288,N_2456);
nor U4036 (N_4036,N_1011,N_1129);
nand U4037 (N_4037,N_1198,N_1655);
nor U4038 (N_4038,N_520,N_196);
nand U4039 (N_4039,N_684,N_350);
nor U4040 (N_4040,N_2092,N_2022);
nand U4041 (N_4041,N_354,N_2497);
nand U4042 (N_4042,N_180,N_424);
and U4043 (N_4043,N_1652,N_181);
nand U4044 (N_4044,N_525,N_973);
and U4045 (N_4045,N_363,N_491);
and U4046 (N_4046,N_2160,N_716);
nand U4047 (N_4047,N_1416,N_1693);
and U4048 (N_4048,N_6,N_65);
or U4049 (N_4049,N_2151,N_1737);
or U4050 (N_4050,N_883,N_717);
and U4051 (N_4051,N_2346,N_1461);
or U4052 (N_4052,N_1162,N_1423);
nor U4053 (N_4053,N_2372,N_573);
and U4054 (N_4054,N_2479,N_410);
or U4055 (N_4055,N_1352,N_1120);
nor U4056 (N_4056,N_485,N_1162);
or U4057 (N_4057,N_463,N_2376);
and U4058 (N_4058,N_316,N_2444);
or U4059 (N_4059,N_2082,N_216);
nor U4060 (N_4060,N_1845,N_2217);
or U4061 (N_4061,N_395,N_17);
nand U4062 (N_4062,N_1430,N_1271);
nor U4063 (N_4063,N_821,N_1817);
or U4064 (N_4064,N_611,N_1277);
nand U4065 (N_4065,N_492,N_2196);
or U4066 (N_4066,N_489,N_1962);
or U4067 (N_4067,N_2355,N_1855);
and U4068 (N_4068,N_798,N_2197);
or U4069 (N_4069,N_1019,N_312);
nand U4070 (N_4070,N_2350,N_1336);
and U4071 (N_4071,N_1989,N_1594);
or U4072 (N_4072,N_383,N_176);
and U4073 (N_4073,N_1370,N_54);
nor U4074 (N_4074,N_575,N_1675);
and U4075 (N_4075,N_153,N_604);
and U4076 (N_4076,N_1380,N_714);
xor U4077 (N_4077,N_1650,N_2462);
or U4078 (N_4078,N_960,N_474);
xor U4079 (N_4079,N_884,N_1185);
nor U4080 (N_4080,N_1501,N_282);
nor U4081 (N_4081,N_673,N_338);
nor U4082 (N_4082,N_1534,N_74);
nand U4083 (N_4083,N_260,N_797);
nor U4084 (N_4084,N_1282,N_1250);
nand U4085 (N_4085,N_770,N_392);
and U4086 (N_4086,N_1876,N_811);
nor U4087 (N_4087,N_1279,N_2094);
or U4088 (N_4088,N_5,N_778);
or U4089 (N_4089,N_841,N_438);
nand U4090 (N_4090,N_2312,N_2185);
nor U4091 (N_4091,N_288,N_792);
and U4092 (N_4092,N_160,N_1708);
nor U4093 (N_4093,N_364,N_561);
nor U4094 (N_4094,N_232,N_1380);
nor U4095 (N_4095,N_1315,N_1004);
and U4096 (N_4096,N_1826,N_1917);
nor U4097 (N_4097,N_587,N_429);
or U4098 (N_4098,N_1941,N_162);
or U4099 (N_4099,N_1142,N_495);
nand U4100 (N_4100,N_1697,N_502);
or U4101 (N_4101,N_2343,N_1846);
and U4102 (N_4102,N_1145,N_1765);
nor U4103 (N_4103,N_783,N_1811);
nand U4104 (N_4104,N_2396,N_336);
and U4105 (N_4105,N_929,N_1329);
nand U4106 (N_4106,N_1708,N_2083);
and U4107 (N_4107,N_2294,N_373);
or U4108 (N_4108,N_740,N_851);
and U4109 (N_4109,N_498,N_513);
nor U4110 (N_4110,N_174,N_1382);
or U4111 (N_4111,N_2340,N_2209);
nand U4112 (N_4112,N_2323,N_953);
xnor U4113 (N_4113,N_622,N_664);
and U4114 (N_4114,N_1881,N_2038);
xnor U4115 (N_4115,N_301,N_2129);
nor U4116 (N_4116,N_2017,N_597);
xor U4117 (N_4117,N_1180,N_2093);
nor U4118 (N_4118,N_571,N_324);
and U4119 (N_4119,N_1106,N_17);
nand U4120 (N_4120,N_2257,N_497);
nand U4121 (N_4121,N_2163,N_2266);
or U4122 (N_4122,N_1021,N_2114);
nor U4123 (N_4123,N_1438,N_1691);
nor U4124 (N_4124,N_163,N_684);
or U4125 (N_4125,N_551,N_1525);
nor U4126 (N_4126,N_2298,N_1967);
and U4127 (N_4127,N_970,N_2438);
and U4128 (N_4128,N_1500,N_1821);
nor U4129 (N_4129,N_782,N_2075);
xnor U4130 (N_4130,N_830,N_1552);
nand U4131 (N_4131,N_126,N_1903);
nor U4132 (N_4132,N_1072,N_600);
or U4133 (N_4133,N_419,N_1394);
and U4134 (N_4134,N_1368,N_969);
nor U4135 (N_4135,N_1948,N_651);
or U4136 (N_4136,N_818,N_1286);
or U4137 (N_4137,N_2406,N_1420);
nor U4138 (N_4138,N_1404,N_2467);
or U4139 (N_4139,N_1190,N_2446);
nor U4140 (N_4140,N_1414,N_1395);
and U4141 (N_4141,N_127,N_1452);
and U4142 (N_4142,N_289,N_1673);
or U4143 (N_4143,N_753,N_2349);
and U4144 (N_4144,N_1143,N_2174);
or U4145 (N_4145,N_1537,N_1003);
or U4146 (N_4146,N_498,N_475);
nand U4147 (N_4147,N_737,N_1091);
or U4148 (N_4148,N_845,N_1347);
or U4149 (N_4149,N_1232,N_475);
or U4150 (N_4150,N_368,N_806);
nand U4151 (N_4151,N_32,N_988);
or U4152 (N_4152,N_399,N_1084);
and U4153 (N_4153,N_534,N_1519);
nand U4154 (N_4154,N_659,N_307);
and U4155 (N_4155,N_2460,N_1214);
nor U4156 (N_4156,N_2320,N_2063);
nand U4157 (N_4157,N_2160,N_246);
nor U4158 (N_4158,N_1962,N_1663);
nor U4159 (N_4159,N_1789,N_629);
or U4160 (N_4160,N_2150,N_73);
nor U4161 (N_4161,N_388,N_1206);
and U4162 (N_4162,N_1969,N_957);
nand U4163 (N_4163,N_82,N_673);
nand U4164 (N_4164,N_1947,N_1489);
and U4165 (N_4165,N_466,N_2084);
nor U4166 (N_4166,N_539,N_1617);
nor U4167 (N_4167,N_2495,N_2036);
and U4168 (N_4168,N_2087,N_1857);
nand U4169 (N_4169,N_2062,N_196);
or U4170 (N_4170,N_2420,N_768);
nor U4171 (N_4171,N_207,N_152);
nor U4172 (N_4172,N_758,N_2075);
nor U4173 (N_4173,N_2408,N_538);
or U4174 (N_4174,N_457,N_1396);
nor U4175 (N_4175,N_60,N_1913);
or U4176 (N_4176,N_215,N_789);
and U4177 (N_4177,N_1437,N_1862);
and U4178 (N_4178,N_1388,N_137);
nor U4179 (N_4179,N_102,N_1935);
nand U4180 (N_4180,N_1450,N_2419);
nor U4181 (N_4181,N_2016,N_203);
and U4182 (N_4182,N_1949,N_800);
and U4183 (N_4183,N_484,N_657);
and U4184 (N_4184,N_1638,N_1117);
nor U4185 (N_4185,N_238,N_1853);
and U4186 (N_4186,N_1014,N_1418);
nand U4187 (N_4187,N_635,N_278);
nor U4188 (N_4188,N_420,N_2493);
and U4189 (N_4189,N_2179,N_1266);
xor U4190 (N_4190,N_994,N_37);
xnor U4191 (N_4191,N_536,N_1942);
nor U4192 (N_4192,N_1245,N_256);
and U4193 (N_4193,N_552,N_150);
or U4194 (N_4194,N_2152,N_2102);
nand U4195 (N_4195,N_1821,N_2301);
nand U4196 (N_4196,N_692,N_2085);
or U4197 (N_4197,N_679,N_65);
nor U4198 (N_4198,N_1756,N_1293);
nand U4199 (N_4199,N_1937,N_2497);
nand U4200 (N_4200,N_2328,N_355);
and U4201 (N_4201,N_570,N_646);
nor U4202 (N_4202,N_1469,N_1434);
nor U4203 (N_4203,N_2199,N_288);
nand U4204 (N_4204,N_1263,N_1642);
or U4205 (N_4205,N_59,N_760);
nor U4206 (N_4206,N_1037,N_2000);
nor U4207 (N_4207,N_4,N_390);
or U4208 (N_4208,N_2223,N_2449);
or U4209 (N_4209,N_1497,N_1129);
and U4210 (N_4210,N_2197,N_1866);
nor U4211 (N_4211,N_501,N_2212);
or U4212 (N_4212,N_2062,N_1720);
nand U4213 (N_4213,N_2090,N_2243);
and U4214 (N_4214,N_122,N_1055);
and U4215 (N_4215,N_945,N_2486);
and U4216 (N_4216,N_743,N_1413);
or U4217 (N_4217,N_358,N_463);
or U4218 (N_4218,N_333,N_1631);
and U4219 (N_4219,N_698,N_1095);
and U4220 (N_4220,N_180,N_27);
nor U4221 (N_4221,N_598,N_2130);
nor U4222 (N_4222,N_1107,N_2068);
and U4223 (N_4223,N_1994,N_152);
and U4224 (N_4224,N_1079,N_1685);
or U4225 (N_4225,N_2016,N_2440);
nand U4226 (N_4226,N_841,N_2361);
nor U4227 (N_4227,N_1832,N_1740);
or U4228 (N_4228,N_807,N_1522);
nand U4229 (N_4229,N_2215,N_1002);
or U4230 (N_4230,N_1663,N_1458);
and U4231 (N_4231,N_303,N_1290);
nand U4232 (N_4232,N_2437,N_1060);
and U4233 (N_4233,N_355,N_498);
or U4234 (N_4234,N_330,N_2285);
or U4235 (N_4235,N_1163,N_2423);
nand U4236 (N_4236,N_335,N_2289);
or U4237 (N_4237,N_1635,N_2136);
or U4238 (N_4238,N_1194,N_1832);
nor U4239 (N_4239,N_1121,N_821);
or U4240 (N_4240,N_29,N_515);
or U4241 (N_4241,N_1578,N_986);
nor U4242 (N_4242,N_1280,N_2021);
nand U4243 (N_4243,N_863,N_169);
xnor U4244 (N_4244,N_771,N_2200);
and U4245 (N_4245,N_583,N_985);
or U4246 (N_4246,N_1125,N_812);
nand U4247 (N_4247,N_222,N_1840);
nor U4248 (N_4248,N_770,N_329);
or U4249 (N_4249,N_1386,N_1789);
nor U4250 (N_4250,N_1982,N_580);
nand U4251 (N_4251,N_1446,N_970);
and U4252 (N_4252,N_464,N_1427);
and U4253 (N_4253,N_918,N_1290);
xnor U4254 (N_4254,N_1763,N_2444);
nand U4255 (N_4255,N_2331,N_553);
nor U4256 (N_4256,N_2121,N_1274);
nand U4257 (N_4257,N_642,N_318);
nand U4258 (N_4258,N_1273,N_2134);
or U4259 (N_4259,N_570,N_762);
nand U4260 (N_4260,N_2218,N_920);
nor U4261 (N_4261,N_766,N_188);
nand U4262 (N_4262,N_120,N_215);
nor U4263 (N_4263,N_1541,N_1413);
nand U4264 (N_4264,N_1896,N_318);
xor U4265 (N_4265,N_2076,N_970);
nor U4266 (N_4266,N_2005,N_1479);
nand U4267 (N_4267,N_1807,N_558);
nand U4268 (N_4268,N_1497,N_2378);
nand U4269 (N_4269,N_1990,N_202);
and U4270 (N_4270,N_2166,N_23);
or U4271 (N_4271,N_1716,N_413);
nor U4272 (N_4272,N_736,N_412);
nand U4273 (N_4273,N_2413,N_1882);
nand U4274 (N_4274,N_1159,N_1882);
or U4275 (N_4275,N_2222,N_2220);
and U4276 (N_4276,N_1282,N_1443);
nand U4277 (N_4277,N_2364,N_1073);
nand U4278 (N_4278,N_1395,N_964);
nor U4279 (N_4279,N_1639,N_726);
nor U4280 (N_4280,N_2283,N_2231);
nor U4281 (N_4281,N_1353,N_1384);
and U4282 (N_4282,N_419,N_772);
or U4283 (N_4283,N_1076,N_1580);
nand U4284 (N_4284,N_1349,N_975);
nand U4285 (N_4285,N_1355,N_278);
and U4286 (N_4286,N_961,N_1267);
nor U4287 (N_4287,N_2391,N_1023);
nand U4288 (N_4288,N_793,N_1674);
nor U4289 (N_4289,N_1085,N_485);
or U4290 (N_4290,N_1416,N_1948);
nor U4291 (N_4291,N_153,N_1638);
nor U4292 (N_4292,N_1264,N_2131);
and U4293 (N_4293,N_118,N_1482);
and U4294 (N_4294,N_620,N_1911);
and U4295 (N_4295,N_201,N_91);
and U4296 (N_4296,N_761,N_2174);
nor U4297 (N_4297,N_467,N_1151);
or U4298 (N_4298,N_899,N_2395);
nand U4299 (N_4299,N_362,N_1965);
nor U4300 (N_4300,N_2144,N_17);
nand U4301 (N_4301,N_2178,N_1894);
nor U4302 (N_4302,N_1816,N_1978);
and U4303 (N_4303,N_1495,N_557);
nand U4304 (N_4304,N_2214,N_286);
nand U4305 (N_4305,N_795,N_536);
and U4306 (N_4306,N_152,N_1097);
and U4307 (N_4307,N_1309,N_1008);
nand U4308 (N_4308,N_40,N_683);
and U4309 (N_4309,N_783,N_1075);
nor U4310 (N_4310,N_180,N_1310);
xnor U4311 (N_4311,N_2199,N_992);
nor U4312 (N_4312,N_2026,N_453);
or U4313 (N_4313,N_2437,N_1080);
nand U4314 (N_4314,N_1873,N_400);
or U4315 (N_4315,N_583,N_1292);
or U4316 (N_4316,N_1653,N_741);
or U4317 (N_4317,N_1531,N_1019);
and U4318 (N_4318,N_229,N_1126);
nand U4319 (N_4319,N_326,N_2261);
nand U4320 (N_4320,N_1649,N_1018);
and U4321 (N_4321,N_59,N_1438);
nand U4322 (N_4322,N_272,N_751);
and U4323 (N_4323,N_682,N_2298);
and U4324 (N_4324,N_1811,N_379);
nor U4325 (N_4325,N_1628,N_1092);
and U4326 (N_4326,N_2286,N_532);
and U4327 (N_4327,N_2479,N_1505);
nor U4328 (N_4328,N_1181,N_1801);
or U4329 (N_4329,N_1636,N_19);
or U4330 (N_4330,N_1844,N_2458);
and U4331 (N_4331,N_700,N_1356);
and U4332 (N_4332,N_862,N_2288);
and U4333 (N_4333,N_1479,N_1601);
nor U4334 (N_4334,N_1549,N_1093);
nand U4335 (N_4335,N_1401,N_2257);
nor U4336 (N_4336,N_2111,N_1684);
nand U4337 (N_4337,N_2117,N_1769);
and U4338 (N_4338,N_2139,N_2201);
nand U4339 (N_4339,N_2149,N_1478);
nor U4340 (N_4340,N_1230,N_2262);
nand U4341 (N_4341,N_14,N_949);
or U4342 (N_4342,N_278,N_856);
and U4343 (N_4343,N_2117,N_1462);
nor U4344 (N_4344,N_1999,N_1523);
xnor U4345 (N_4345,N_2182,N_1509);
nand U4346 (N_4346,N_1878,N_2261);
and U4347 (N_4347,N_985,N_1260);
or U4348 (N_4348,N_708,N_150);
nor U4349 (N_4349,N_2393,N_431);
nor U4350 (N_4350,N_2457,N_2491);
and U4351 (N_4351,N_985,N_1724);
or U4352 (N_4352,N_561,N_2285);
nand U4353 (N_4353,N_1797,N_1958);
or U4354 (N_4354,N_1062,N_205);
nand U4355 (N_4355,N_1468,N_2472);
nor U4356 (N_4356,N_1786,N_1073);
or U4357 (N_4357,N_1751,N_1944);
or U4358 (N_4358,N_1829,N_731);
and U4359 (N_4359,N_100,N_1632);
nor U4360 (N_4360,N_971,N_2376);
nand U4361 (N_4361,N_1916,N_2496);
nand U4362 (N_4362,N_314,N_1189);
nor U4363 (N_4363,N_464,N_2164);
nor U4364 (N_4364,N_2458,N_2111);
nor U4365 (N_4365,N_1775,N_170);
and U4366 (N_4366,N_2223,N_439);
nand U4367 (N_4367,N_1968,N_893);
nand U4368 (N_4368,N_2109,N_1121);
xor U4369 (N_4369,N_457,N_371);
nand U4370 (N_4370,N_289,N_1653);
nor U4371 (N_4371,N_2493,N_968);
or U4372 (N_4372,N_1545,N_1903);
or U4373 (N_4373,N_1364,N_1967);
and U4374 (N_4374,N_810,N_335);
and U4375 (N_4375,N_2483,N_1302);
nand U4376 (N_4376,N_2167,N_1379);
and U4377 (N_4377,N_2021,N_1994);
or U4378 (N_4378,N_2353,N_264);
nor U4379 (N_4379,N_1325,N_1727);
nor U4380 (N_4380,N_1441,N_1372);
or U4381 (N_4381,N_906,N_755);
nor U4382 (N_4382,N_984,N_1585);
nor U4383 (N_4383,N_2285,N_1807);
nor U4384 (N_4384,N_20,N_45);
nor U4385 (N_4385,N_52,N_585);
or U4386 (N_4386,N_1174,N_2368);
or U4387 (N_4387,N_531,N_2343);
nor U4388 (N_4388,N_1912,N_982);
and U4389 (N_4389,N_453,N_1569);
or U4390 (N_4390,N_2215,N_2276);
nor U4391 (N_4391,N_676,N_2359);
and U4392 (N_4392,N_244,N_662);
and U4393 (N_4393,N_377,N_1275);
or U4394 (N_4394,N_397,N_287);
nand U4395 (N_4395,N_2455,N_566);
or U4396 (N_4396,N_1694,N_929);
nand U4397 (N_4397,N_940,N_755);
nor U4398 (N_4398,N_1673,N_720);
nand U4399 (N_4399,N_825,N_839);
nand U4400 (N_4400,N_2494,N_2026);
nor U4401 (N_4401,N_1651,N_1289);
or U4402 (N_4402,N_1851,N_649);
nand U4403 (N_4403,N_33,N_2258);
nor U4404 (N_4404,N_1677,N_306);
nor U4405 (N_4405,N_1855,N_856);
and U4406 (N_4406,N_1312,N_1904);
nor U4407 (N_4407,N_1708,N_2175);
or U4408 (N_4408,N_918,N_90);
nor U4409 (N_4409,N_1603,N_940);
nand U4410 (N_4410,N_211,N_2372);
and U4411 (N_4411,N_2040,N_705);
nor U4412 (N_4412,N_2383,N_2176);
and U4413 (N_4413,N_1020,N_1170);
and U4414 (N_4414,N_650,N_1644);
or U4415 (N_4415,N_2310,N_492);
or U4416 (N_4416,N_246,N_408);
nand U4417 (N_4417,N_683,N_543);
nand U4418 (N_4418,N_2112,N_622);
nor U4419 (N_4419,N_1821,N_844);
or U4420 (N_4420,N_256,N_116);
nand U4421 (N_4421,N_931,N_1286);
nor U4422 (N_4422,N_1588,N_494);
nor U4423 (N_4423,N_1489,N_924);
nand U4424 (N_4424,N_1107,N_856);
and U4425 (N_4425,N_2255,N_2317);
or U4426 (N_4426,N_438,N_1820);
or U4427 (N_4427,N_7,N_1946);
nor U4428 (N_4428,N_1464,N_2438);
nand U4429 (N_4429,N_1496,N_2024);
and U4430 (N_4430,N_2021,N_799);
and U4431 (N_4431,N_820,N_2255);
nand U4432 (N_4432,N_1179,N_2340);
nand U4433 (N_4433,N_2263,N_2405);
or U4434 (N_4434,N_687,N_1519);
nand U4435 (N_4435,N_225,N_1523);
or U4436 (N_4436,N_2454,N_1397);
nand U4437 (N_4437,N_1103,N_1284);
nor U4438 (N_4438,N_2354,N_2120);
and U4439 (N_4439,N_2427,N_2416);
nor U4440 (N_4440,N_255,N_2173);
nor U4441 (N_4441,N_265,N_2322);
nand U4442 (N_4442,N_1139,N_396);
nor U4443 (N_4443,N_1895,N_1894);
and U4444 (N_4444,N_177,N_948);
nand U4445 (N_4445,N_1499,N_1564);
or U4446 (N_4446,N_2098,N_1499);
and U4447 (N_4447,N_797,N_2179);
or U4448 (N_4448,N_1375,N_1549);
or U4449 (N_4449,N_43,N_1782);
nor U4450 (N_4450,N_268,N_1452);
nor U4451 (N_4451,N_713,N_1172);
and U4452 (N_4452,N_2407,N_1892);
or U4453 (N_4453,N_1231,N_1232);
nor U4454 (N_4454,N_581,N_1881);
nor U4455 (N_4455,N_83,N_80);
nor U4456 (N_4456,N_1229,N_651);
and U4457 (N_4457,N_553,N_129);
nand U4458 (N_4458,N_257,N_759);
or U4459 (N_4459,N_819,N_1497);
nor U4460 (N_4460,N_57,N_2438);
nor U4461 (N_4461,N_1855,N_1240);
nand U4462 (N_4462,N_1900,N_229);
nand U4463 (N_4463,N_845,N_589);
and U4464 (N_4464,N_1293,N_1347);
or U4465 (N_4465,N_2194,N_802);
and U4466 (N_4466,N_1106,N_1709);
and U4467 (N_4467,N_597,N_479);
nor U4468 (N_4468,N_1979,N_1137);
or U4469 (N_4469,N_2324,N_258);
or U4470 (N_4470,N_1107,N_1334);
nand U4471 (N_4471,N_1000,N_418);
nor U4472 (N_4472,N_1075,N_1293);
nor U4473 (N_4473,N_2079,N_455);
nor U4474 (N_4474,N_2454,N_2158);
nor U4475 (N_4475,N_683,N_553);
nor U4476 (N_4476,N_776,N_1944);
and U4477 (N_4477,N_236,N_937);
nand U4478 (N_4478,N_724,N_1073);
nor U4479 (N_4479,N_885,N_2190);
nor U4480 (N_4480,N_70,N_1675);
and U4481 (N_4481,N_1316,N_1785);
nor U4482 (N_4482,N_251,N_574);
xnor U4483 (N_4483,N_293,N_481);
nand U4484 (N_4484,N_681,N_902);
nor U4485 (N_4485,N_1587,N_1330);
nor U4486 (N_4486,N_128,N_705);
nand U4487 (N_4487,N_342,N_1159);
nand U4488 (N_4488,N_153,N_571);
nor U4489 (N_4489,N_313,N_769);
or U4490 (N_4490,N_268,N_1613);
or U4491 (N_4491,N_2022,N_520);
nor U4492 (N_4492,N_968,N_390);
or U4493 (N_4493,N_1446,N_147);
or U4494 (N_4494,N_1898,N_1761);
nor U4495 (N_4495,N_1055,N_1200);
nor U4496 (N_4496,N_647,N_975);
and U4497 (N_4497,N_485,N_1979);
nor U4498 (N_4498,N_460,N_2407);
nand U4499 (N_4499,N_321,N_2488);
and U4500 (N_4500,N_2432,N_1664);
xnor U4501 (N_4501,N_1343,N_886);
and U4502 (N_4502,N_2453,N_1687);
or U4503 (N_4503,N_1139,N_2468);
and U4504 (N_4504,N_2217,N_698);
nand U4505 (N_4505,N_572,N_1909);
or U4506 (N_4506,N_1603,N_430);
xnor U4507 (N_4507,N_2358,N_134);
or U4508 (N_4508,N_732,N_2348);
or U4509 (N_4509,N_1077,N_511);
or U4510 (N_4510,N_792,N_198);
and U4511 (N_4511,N_2224,N_1529);
or U4512 (N_4512,N_1155,N_178);
and U4513 (N_4513,N_1103,N_2155);
and U4514 (N_4514,N_1734,N_1176);
nor U4515 (N_4515,N_343,N_749);
or U4516 (N_4516,N_1602,N_274);
or U4517 (N_4517,N_1639,N_236);
nor U4518 (N_4518,N_958,N_1774);
and U4519 (N_4519,N_1566,N_1651);
nor U4520 (N_4520,N_2453,N_1557);
or U4521 (N_4521,N_331,N_196);
nand U4522 (N_4522,N_2250,N_91);
nand U4523 (N_4523,N_2055,N_1091);
nand U4524 (N_4524,N_1288,N_1708);
and U4525 (N_4525,N_910,N_400);
and U4526 (N_4526,N_2067,N_820);
and U4527 (N_4527,N_1876,N_1616);
nand U4528 (N_4528,N_174,N_1182);
nor U4529 (N_4529,N_800,N_1336);
or U4530 (N_4530,N_616,N_662);
and U4531 (N_4531,N_1651,N_1530);
or U4532 (N_4532,N_2232,N_1258);
or U4533 (N_4533,N_1188,N_980);
and U4534 (N_4534,N_2074,N_329);
nand U4535 (N_4535,N_1853,N_940);
nor U4536 (N_4536,N_2131,N_1347);
nor U4537 (N_4537,N_762,N_1052);
and U4538 (N_4538,N_1234,N_1420);
or U4539 (N_4539,N_280,N_600);
nand U4540 (N_4540,N_1636,N_1235);
nand U4541 (N_4541,N_139,N_1332);
or U4542 (N_4542,N_1392,N_941);
nor U4543 (N_4543,N_679,N_1605);
or U4544 (N_4544,N_974,N_1844);
nand U4545 (N_4545,N_2424,N_2373);
nand U4546 (N_4546,N_2259,N_467);
and U4547 (N_4547,N_286,N_1243);
and U4548 (N_4548,N_2090,N_1042);
nor U4549 (N_4549,N_254,N_2497);
and U4550 (N_4550,N_1553,N_602);
nand U4551 (N_4551,N_2117,N_1377);
nand U4552 (N_4552,N_1738,N_1359);
or U4553 (N_4553,N_2228,N_2018);
nor U4554 (N_4554,N_192,N_2202);
and U4555 (N_4555,N_305,N_1088);
nor U4556 (N_4556,N_861,N_777);
nand U4557 (N_4557,N_1359,N_419);
nand U4558 (N_4558,N_425,N_127);
nor U4559 (N_4559,N_1248,N_1711);
or U4560 (N_4560,N_942,N_1518);
nand U4561 (N_4561,N_275,N_867);
nand U4562 (N_4562,N_1962,N_2194);
nor U4563 (N_4563,N_103,N_2232);
nor U4564 (N_4564,N_387,N_1635);
nand U4565 (N_4565,N_1156,N_522);
or U4566 (N_4566,N_1675,N_1666);
and U4567 (N_4567,N_1511,N_2455);
nand U4568 (N_4568,N_2447,N_1703);
nand U4569 (N_4569,N_2498,N_1638);
nor U4570 (N_4570,N_1287,N_991);
xor U4571 (N_4571,N_1814,N_22);
and U4572 (N_4572,N_2001,N_799);
nand U4573 (N_4573,N_1613,N_2346);
xor U4574 (N_4574,N_1926,N_210);
and U4575 (N_4575,N_1661,N_1043);
and U4576 (N_4576,N_1189,N_955);
nand U4577 (N_4577,N_10,N_1807);
or U4578 (N_4578,N_1597,N_1896);
or U4579 (N_4579,N_587,N_206);
nor U4580 (N_4580,N_2343,N_2061);
or U4581 (N_4581,N_1572,N_1132);
and U4582 (N_4582,N_942,N_899);
nor U4583 (N_4583,N_1561,N_502);
nor U4584 (N_4584,N_2442,N_1724);
nand U4585 (N_4585,N_2025,N_883);
and U4586 (N_4586,N_693,N_1219);
and U4587 (N_4587,N_1929,N_1736);
and U4588 (N_4588,N_2368,N_2149);
and U4589 (N_4589,N_35,N_2172);
and U4590 (N_4590,N_163,N_1702);
or U4591 (N_4591,N_807,N_1251);
nand U4592 (N_4592,N_850,N_447);
or U4593 (N_4593,N_1603,N_1932);
and U4594 (N_4594,N_1904,N_1211);
and U4595 (N_4595,N_1672,N_203);
or U4596 (N_4596,N_202,N_1483);
or U4597 (N_4597,N_691,N_1323);
nand U4598 (N_4598,N_724,N_1795);
nor U4599 (N_4599,N_1705,N_1380);
nor U4600 (N_4600,N_399,N_2272);
or U4601 (N_4601,N_2338,N_776);
nor U4602 (N_4602,N_509,N_231);
nand U4603 (N_4603,N_1020,N_2234);
and U4604 (N_4604,N_101,N_1459);
nand U4605 (N_4605,N_1382,N_2271);
nor U4606 (N_4606,N_1720,N_939);
and U4607 (N_4607,N_679,N_1598);
nand U4608 (N_4608,N_757,N_1104);
nand U4609 (N_4609,N_412,N_14);
and U4610 (N_4610,N_1726,N_2081);
or U4611 (N_4611,N_2457,N_539);
nor U4612 (N_4612,N_1605,N_1750);
and U4613 (N_4613,N_1119,N_1685);
xnor U4614 (N_4614,N_1582,N_2371);
and U4615 (N_4615,N_369,N_81);
nor U4616 (N_4616,N_1897,N_1896);
and U4617 (N_4617,N_191,N_1036);
and U4618 (N_4618,N_615,N_903);
and U4619 (N_4619,N_1562,N_1672);
nor U4620 (N_4620,N_1531,N_723);
nor U4621 (N_4621,N_1856,N_48);
nor U4622 (N_4622,N_1641,N_103);
and U4623 (N_4623,N_1573,N_677);
nand U4624 (N_4624,N_2117,N_2115);
nand U4625 (N_4625,N_539,N_143);
nand U4626 (N_4626,N_1875,N_1644);
xnor U4627 (N_4627,N_773,N_2099);
or U4628 (N_4628,N_35,N_894);
nand U4629 (N_4629,N_308,N_1666);
or U4630 (N_4630,N_2137,N_1948);
nor U4631 (N_4631,N_1287,N_2429);
and U4632 (N_4632,N_1571,N_1064);
and U4633 (N_4633,N_714,N_2437);
nor U4634 (N_4634,N_581,N_1429);
nand U4635 (N_4635,N_1969,N_1379);
xnor U4636 (N_4636,N_2437,N_148);
nand U4637 (N_4637,N_1336,N_639);
nor U4638 (N_4638,N_1541,N_2277);
and U4639 (N_4639,N_2060,N_1997);
or U4640 (N_4640,N_475,N_1633);
or U4641 (N_4641,N_2477,N_1185);
and U4642 (N_4642,N_180,N_2206);
and U4643 (N_4643,N_1040,N_1111);
and U4644 (N_4644,N_974,N_223);
or U4645 (N_4645,N_2121,N_2255);
xnor U4646 (N_4646,N_1092,N_1498);
nor U4647 (N_4647,N_2364,N_382);
nor U4648 (N_4648,N_923,N_241);
nand U4649 (N_4649,N_1727,N_1210);
and U4650 (N_4650,N_134,N_2496);
nor U4651 (N_4651,N_138,N_2384);
nor U4652 (N_4652,N_1363,N_1482);
or U4653 (N_4653,N_502,N_2009);
nor U4654 (N_4654,N_308,N_1539);
nand U4655 (N_4655,N_1107,N_57);
nor U4656 (N_4656,N_2411,N_1548);
and U4657 (N_4657,N_1225,N_778);
and U4658 (N_4658,N_1834,N_2456);
nand U4659 (N_4659,N_1662,N_381);
or U4660 (N_4660,N_2260,N_349);
or U4661 (N_4661,N_884,N_719);
and U4662 (N_4662,N_462,N_1569);
and U4663 (N_4663,N_2438,N_1928);
nand U4664 (N_4664,N_568,N_1147);
nand U4665 (N_4665,N_1372,N_1173);
nor U4666 (N_4666,N_1152,N_2378);
nor U4667 (N_4667,N_1647,N_201);
nor U4668 (N_4668,N_1950,N_1136);
and U4669 (N_4669,N_1127,N_1651);
nor U4670 (N_4670,N_2224,N_1200);
nand U4671 (N_4671,N_1409,N_1309);
and U4672 (N_4672,N_2382,N_2083);
nand U4673 (N_4673,N_358,N_907);
and U4674 (N_4674,N_1617,N_2463);
nor U4675 (N_4675,N_494,N_2193);
and U4676 (N_4676,N_2369,N_506);
or U4677 (N_4677,N_2483,N_884);
nor U4678 (N_4678,N_2498,N_19);
nand U4679 (N_4679,N_529,N_1984);
xnor U4680 (N_4680,N_1073,N_577);
and U4681 (N_4681,N_200,N_1343);
xor U4682 (N_4682,N_1569,N_1269);
or U4683 (N_4683,N_988,N_1707);
nor U4684 (N_4684,N_1197,N_2272);
or U4685 (N_4685,N_1596,N_1683);
and U4686 (N_4686,N_409,N_783);
or U4687 (N_4687,N_946,N_2341);
nand U4688 (N_4688,N_606,N_1762);
or U4689 (N_4689,N_658,N_1001);
or U4690 (N_4690,N_741,N_895);
nor U4691 (N_4691,N_1582,N_65);
nor U4692 (N_4692,N_2449,N_1009);
nand U4693 (N_4693,N_27,N_1783);
nand U4694 (N_4694,N_1597,N_1586);
or U4695 (N_4695,N_18,N_1742);
nor U4696 (N_4696,N_1755,N_1006);
or U4697 (N_4697,N_2442,N_2096);
nand U4698 (N_4698,N_364,N_1366);
and U4699 (N_4699,N_1512,N_507);
or U4700 (N_4700,N_1618,N_1299);
and U4701 (N_4701,N_2102,N_1498);
or U4702 (N_4702,N_2419,N_1862);
nor U4703 (N_4703,N_111,N_820);
and U4704 (N_4704,N_2179,N_2176);
and U4705 (N_4705,N_2431,N_1066);
nor U4706 (N_4706,N_897,N_1750);
xor U4707 (N_4707,N_789,N_1323);
nor U4708 (N_4708,N_1666,N_1926);
and U4709 (N_4709,N_1939,N_2091);
or U4710 (N_4710,N_361,N_233);
or U4711 (N_4711,N_8,N_2328);
and U4712 (N_4712,N_2210,N_675);
or U4713 (N_4713,N_924,N_2203);
nand U4714 (N_4714,N_72,N_2011);
and U4715 (N_4715,N_1164,N_850);
nand U4716 (N_4716,N_688,N_2441);
or U4717 (N_4717,N_2413,N_758);
nand U4718 (N_4718,N_1627,N_250);
nor U4719 (N_4719,N_1163,N_515);
xor U4720 (N_4720,N_1538,N_477);
xor U4721 (N_4721,N_1363,N_1418);
or U4722 (N_4722,N_77,N_2434);
or U4723 (N_4723,N_668,N_1202);
and U4724 (N_4724,N_1660,N_257);
or U4725 (N_4725,N_1871,N_1894);
nor U4726 (N_4726,N_291,N_354);
or U4727 (N_4727,N_1533,N_271);
xnor U4728 (N_4728,N_975,N_1240);
or U4729 (N_4729,N_1872,N_419);
nor U4730 (N_4730,N_864,N_1914);
and U4731 (N_4731,N_441,N_2481);
or U4732 (N_4732,N_1938,N_2278);
and U4733 (N_4733,N_1561,N_1230);
nor U4734 (N_4734,N_2171,N_578);
nor U4735 (N_4735,N_2298,N_1319);
nor U4736 (N_4736,N_1138,N_16);
or U4737 (N_4737,N_2309,N_2471);
nor U4738 (N_4738,N_156,N_1398);
and U4739 (N_4739,N_2009,N_2475);
nand U4740 (N_4740,N_1439,N_1681);
nor U4741 (N_4741,N_2066,N_605);
and U4742 (N_4742,N_1337,N_718);
or U4743 (N_4743,N_784,N_442);
or U4744 (N_4744,N_1107,N_794);
and U4745 (N_4745,N_1750,N_953);
nor U4746 (N_4746,N_2458,N_1833);
and U4747 (N_4747,N_2461,N_1157);
xor U4748 (N_4748,N_586,N_360);
xnor U4749 (N_4749,N_287,N_2002);
and U4750 (N_4750,N_947,N_1939);
and U4751 (N_4751,N_917,N_1779);
nor U4752 (N_4752,N_2297,N_2083);
and U4753 (N_4753,N_1595,N_1137);
and U4754 (N_4754,N_578,N_1214);
nand U4755 (N_4755,N_240,N_1498);
nand U4756 (N_4756,N_31,N_896);
nand U4757 (N_4757,N_1245,N_2465);
nand U4758 (N_4758,N_493,N_1119);
and U4759 (N_4759,N_1358,N_1952);
or U4760 (N_4760,N_2304,N_2278);
nor U4761 (N_4761,N_963,N_701);
nor U4762 (N_4762,N_1034,N_214);
xnor U4763 (N_4763,N_569,N_1317);
or U4764 (N_4764,N_1632,N_1570);
and U4765 (N_4765,N_54,N_2422);
or U4766 (N_4766,N_865,N_954);
or U4767 (N_4767,N_178,N_2394);
or U4768 (N_4768,N_2484,N_2212);
nand U4769 (N_4769,N_648,N_122);
or U4770 (N_4770,N_364,N_1556);
nor U4771 (N_4771,N_1626,N_234);
nor U4772 (N_4772,N_818,N_1999);
nor U4773 (N_4773,N_530,N_1551);
nor U4774 (N_4774,N_1186,N_543);
or U4775 (N_4775,N_798,N_1866);
and U4776 (N_4776,N_1355,N_1384);
nand U4777 (N_4777,N_23,N_1409);
nor U4778 (N_4778,N_1692,N_422);
nand U4779 (N_4779,N_1440,N_1875);
and U4780 (N_4780,N_1072,N_151);
nor U4781 (N_4781,N_832,N_2017);
and U4782 (N_4782,N_743,N_1027);
nor U4783 (N_4783,N_599,N_1553);
and U4784 (N_4784,N_2373,N_2007);
nand U4785 (N_4785,N_102,N_560);
or U4786 (N_4786,N_2007,N_1048);
nor U4787 (N_4787,N_955,N_1185);
or U4788 (N_4788,N_887,N_479);
nor U4789 (N_4789,N_993,N_725);
or U4790 (N_4790,N_2101,N_1664);
and U4791 (N_4791,N_1404,N_1417);
nand U4792 (N_4792,N_532,N_335);
xor U4793 (N_4793,N_305,N_1607);
nand U4794 (N_4794,N_729,N_2031);
xnor U4795 (N_4795,N_2008,N_2140);
xnor U4796 (N_4796,N_818,N_335);
and U4797 (N_4797,N_533,N_1831);
and U4798 (N_4798,N_1293,N_2354);
xor U4799 (N_4799,N_1100,N_271);
nor U4800 (N_4800,N_124,N_1748);
or U4801 (N_4801,N_1436,N_1754);
or U4802 (N_4802,N_1982,N_2342);
or U4803 (N_4803,N_867,N_2273);
and U4804 (N_4804,N_2281,N_2273);
nor U4805 (N_4805,N_1154,N_624);
and U4806 (N_4806,N_1694,N_2116);
or U4807 (N_4807,N_1358,N_134);
nor U4808 (N_4808,N_671,N_1796);
and U4809 (N_4809,N_1706,N_1345);
nand U4810 (N_4810,N_512,N_1178);
nand U4811 (N_4811,N_1920,N_1143);
nand U4812 (N_4812,N_1489,N_1174);
or U4813 (N_4813,N_2496,N_900);
and U4814 (N_4814,N_2245,N_2148);
nor U4815 (N_4815,N_1152,N_1666);
xnor U4816 (N_4816,N_2015,N_662);
nor U4817 (N_4817,N_503,N_2416);
nand U4818 (N_4818,N_154,N_151);
nor U4819 (N_4819,N_1674,N_574);
or U4820 (N_4820,N_129,N_1552);
and U4821 (N_4821,N_1151,N_136);
or U4822 (N_4822,N_666,N_2089);
and U4823 (N_4823,N_521,N_1088);
xor U4824 (N_4824,N_2465,N_1053);
nand U4825 (N_4825,N_1193,N_2130);
nor U4826 (N_4826,N_191,N_50);
or U4827 (N_4827,N_1077,N_559);
or U4828 (N_4828,N_1025,N_562);
nor U4829 (N_4829,N_332,N_1873);
nand U4830 (N_4830,N_322,N_2363);
or U4831 (N_4831,N_198,N_2230);
xor U4832 (N_4832,N_1354,N_1678);
nor U4833 (N_4833,N_1908,N_797);
and U4834 (N_4834,N_525,N_2113);
or U4835 (N_4835,N_2473,N_301);
nand U4836 (N_4836,N_379,N_816);
and U4837 (N_4837,N_693,N_385);
nor U4838 (N_4838,N_697,N_2198);
or U4839 (N_4839,N_774,N_852);
or U4840 (N_4840,N_1736,N_128);
nand U4841 (N_4841,N_217,N_1172);
and U4842 (N_4842,N_2421,N_2271);
nand U4843 (N_4843,N_259,N_1077);
nor U4844 (N_4844,N_2081,N_105);
or U4845 (N_4845,N_780,N_1895);
or U4846 (N_4846,N_890,N_1902);
nand U4847 (N_4847,N_1343,N_1966);
nor U4848 (N_4848,N_524,N_1987);
and U4849 (N_4849,N_79,N_1179);
nor U4850 (N_4850,N_1661,N_543);
and U4851 (N_4851,N_2145,N_562);
nand U4852 (N_4852,N_1950,N_195);
or U4853 (N_4853,N_1420,N_707);
or U4854 (N_4854,N_1254,N_944);
or U4855 (N_4855,N_1158,N_2226);
nand U4856 (N_4856,N_26,N_2093);
nor U4857 (N_4857,N_1830,N_185);
and U4858 (N_4858,N_1177,N_1778);
nand U4859 (N_4859,N_594,N_786);
nand U4860 (N_4860,N_1725,N_134);
and U4861 (N_4861,N_702,N_1285);
or U4862 (N_4862,N_692,N_487);
nor U4863 (N_4863,N_2218,N_1308);
or U4864 (N_4864,N_827,N_1488);
nand U4865 (N_4865,N_352,N_1989);
or U4866 (N_4866,N_1509,N_1364);
nor U4867 (N_4867,N_326,N_1018);
nor U4868 (N_4868,N_1891,N_647);
nor U4869 (N_4869,N_900,N_1288);
and U4870 (N_4870,N_93,N_2364);
and U4871 (N_4871,N_1700,N_380);
or U4872 (N_4872,N_1331,N_959);
nand U4873 (N_4873,N_662,N_198);
nor U4874 (N_4874,N_2300,N_689);
and U4875 (N_4875,N_1512,N_172);
nor U4876 (N_4876,N_1484,N_279);
and U4877 (N_4877,N_1252,N_1113);
or U4878 (N_4878,N_2249,N_1498);
and U4879 (N_4879,N_561,N_2499);
or U4880 (N_4880,N_1838,N_1946);
and U4881 (N_4881,N_1146,N_260);
and U4882 (N_4882,N_442,N_1859);
nor U4883 (N_4883,N_23,N_459);
and U4884 (N_4884,N_2487,N_2117);
and U4885 (N_4885,N_2233,N_1104);
and U4886 (N_4886,N_1719,N_692);
nand U4887 (N_4887,N_1903,N_783);
nor U4888 (N_4888,N_2393,N_558);
nor U4889 (N_4889,N_173,N_79);
and U4890 (N_4890,N_148,N_1059);
nand U4891 (N_4891,N_1147,N_221);
nor U4892 (N_4892,N_1255,N_861);
nand U4893 (N_4893,N_2269,N_445);
nand U4894 (N_4894,N_2270,N_2453);
or U4895 (N_4895,N_274,N_1621);
or U4896 (N_4896,N_69,N_1479);
and U4897 (N_4897,N_880,N_1879);
nor U4898 (N_4898,N_1557,N_1701);
and U4899 (N_4899,N_1130,N_2023);
nand U4900 (N_4900,N_1448,N_1124);
and U4901 (N_4901,N_2180,N_654);
nand U4902 (N_4902,N_6,N_2277);
nand U4903 (N_4903,N_1069,N_2247);
and U4904 (N_4904,N_1624,N_1417);
nor U4905 (N_4905,N_1799,N_1374);
nor U4906 (N_4906,N_1199,N_1863);
and U4907 (N_4907,N_55,N_1178);
and U4908 (N_4908,N_1571,N_2267);
or U4909 (N_4909,N_2406,N_1093);
or U4910 (N_4910,N_1607,N_1189);
or U4911 (N_4911,N_1646,N_2098);
and U4912 (N_4912,N_663,N_208);
or U4913 (N_4913,N_310,N_603);
nand U4914 (N_4914,N_1325,N_1847);
or U4915 (N_4915,N_1756,N_1635);
or U4916 (N_4916,N_2147,N_269);
nand U4917 (N_4917,N_885,N_869);
or U4918 (N_4918,N_1484,N_1947);
or U4919 (N_4919,N_341,N_87);
nor U4920 (N_4920,N_2032,N_950);
nand U4921 (N_4921,N_457,N_1067);
and U4922 (N_4922,N_831,N_2412);
or U4923 (N_4923,N_668,N_1033);
nand U4924 (N_4924,N_1021,N_2097);
or U4925 (N_4925,N_1361,N_4);
nor U4926 (N_4926,N_515,N_591);
nor U4927 (N_4927,N_119,N_1927);
and U4928 (N_4928,N_639,N_345);
nand U4929 (N_4929,N_2148,N_318);
and U4930 (N_4930,N_1141,N_1161);
and U4931 (N_4931,N_1474,N_2207);
nor U4932 (N_4932,N_2238,N_1416);
nand U4933 (N_4933,N_1374,N_310);
nand U4934 (N_4934,N_370,N_1532);
or U4935 (N_4935,N_2239,N_472);
or U4936 (N_4936,N_374,N_728);
and U4937 (N_4937,N_2228,N_2048);
nor U4938 (N_4938,N_1583,N_510);
and U4939 (N_4939,N_1331,N_968);
nor U4940 (N_4940,N_852,N_552);
nand U4941 (N_4941,N_1124,N_694);
or U4942 (N_4942,N_934,N_768);
or U4943 (N_4943,N_2124,N_194);
or U4944 (N_4944,N_506,N_286);
or U4945 (N_4945,N_1503,N_1114);
or U4946 (N_4946,N_756,N_106);
xnor U4947 (N_4947,N_1387,N_910);
and U4948 (N_4948,N_2456,N_205);
xnor U4949 (N_4949,N_424,N_2346);
and U4950 (N_4950,N_339,N_1560);
or U4951 (N_4951,N_1328,N_863);
or U4952 (N_4952,N_1906,N_1636);
nor U4953 (N_4953,N_2327,N_1666);
nor U4954 (N_4954,N_1307,N_469);
and U4955 (N_4955,N_463,N_403);
or U4956 (N_4956,N_2004,N_895);
nor U4957 (N_4957,N_1295,N_1799);
nor U4958 (N_4958,N_1783,N_2362);
nor U4959 (N_4959,N_1059,N_2123);
or U4960 (N_4960,N_2468,N_1332);
or U4961 (N_4961,N_321,N_2479);
nor U4962 (N_4962,N_82,N_32);
or U4963 (N_4963,N_1495,N_34);
nand U4964 (N_4964,N_295,N_2067);
nor U4965 (N_4965,N_514,N_1514);
and U4966 (N_4966,N_1463,N_469);
and U4967 (N_4967,N_1982,N_945);
nor U4968 (N_4968,N_2139,N_2007);
and U4969 (N_4969,N_1097,N_1297);
nand U4970 (N_4970,N_1103,N_1611);
or U4971 (N_4971,N_351,N_2255);
and U4972 (N_4972,N_1474,N_341);
or U4973 (N_4973,N_2137,N_1258);
nand U4974 (N_4974,N_2482,N_1698);
or U4975 (N_4975,N_2312,N_1910);
or U4976 (N_4976,N_1027,N_1225);
nand U4977 (N_4977,N_1596,N_1011);
nor U4978 (N_4978,N_22,N_2064);
and U4979 (N_4979,N_789,N_1140);
nor U4980 (N_4980,N_2069,N_2410);
and U4981 (N_4981,N_664,N_1335);
or U4982 (N_4982,N_2251,N_835);
nor U4983 (N_4983,N_1915,N_1676);
nor U4984 (N_4984,N_1488,N_1313);
nor U4985 (N_4985,N_2281,N_2000);
xnor U4986 (N_4986,N_2483,N_1732);
nand U4987 (N_4987,N_2446,N_2452);
nor U4988 (N_4988,N_1512,N_2338);
and U4989 (N_4989,N_1410,N_389);
and U4990 (N_4990,N_1888,N_615);
and U4991 (N_4991,N_1586,N_986);
nor U4992 (N_4992,N_2452,N_2065);
nand U4993 (N_4993,N_557,N_2426);
xnor U4994 (N_4994,N_1068,N_1367);
or U4995 (N_4995,N_2414,N_1265);
nand U4996 (N_4996,N_2307,N_2468);
nand U4997 (N_4997,N_462,N_948);
nand U4998 (N_4998,N_2181,N_368);
and U4999 (N_4999,N_2450,N_1162);
or U5000 (N_5000,N_4967,N_4261);
nand U5001 (N_5001,N_4505,N_4718);
and U5002 (N_5002,N_2779,N_3855);
nor U5003 (N_5003,N_4957,N_2694);
nor U5004 (N_5004,N_2579,N_3014);
or U5005 (N_5005,N_3270,N_4551);
nand U5006 (N_5006,N_3577,N_4041);
and U5007 (N_5007,N_2558,N_2555);
nand U5008 (N_5008,N_3903,N_4402);
nand U5009 (N_5009,N_2968,N_4230);
and U5010 (N_5010,N_3991,N_3022);
xnor U5011 (N_5011,N_4308,N_4013);
nor U5012 (N_5012,N_3243,N_3558);
nand U5013 (N_5013,N_3866,N_4382);
nor U5014 (N_5014,N_4777,N_4122);
or U5015 (N_5015,N_3478,N_3203);
nor U5016 (N_5016,N_3811,N_4012);
nand U5017 (N_5017,N_3027,N_3017);
nor U5018 (N_5018,N_3928,N_4866);
and U5019 (N_5019,N_2552,N_4670);
and U5020 (N_5020,N_3808,N_3926);
nor U5021 (N_5021,N_3396,N_2526);
and U5022 (N_5022,N_2587,N_4445);
and U5023 (N_5023,N_4702,N_3562);
and U5024 (N_5024,N_2812,N_2863);
and U5025 (N_5025,N_4606,N_3605);
or U5026 (N_5026,N_3216,N_3776);
xor U5027 (N_5027,N_4137,N_3366);
nor U5028 (N_5028,N_3629,N_4085);
nand U5029 (N_5029,N_3631,N_3563);
nand U5030 (N_5030,N_3876,N_2749);
nor U5031 (N_5031,N_4274,N_3362);
nand U5032 (N_5032,N_3600,N_4635);
or U5033 (N_5033,N_4193,N_4146);
nand U5034 (N_5034,N_3934,N_4808);
or U5035 (N_5035,N_2818,N_3601);
nand U5036 (N_5036,N_4864,N_2972);
and U5037 (N_5037,N_4961,N_4069);
nand U5038 (N_5038,N_2953,N_3268);
nor U5039 (N_5039,N_4185,N_3395);
and U5040 (N_5040,N_4344,N_3594);
and U5041 (N_5041,N_4253,N_4538);
or U5042 (N_5042,N_4731,N_2997);
nand U5043 (N_5043,N_3127,N_4802);
nor U5044 (N_5044,N_4296,N_4201);
and U5045 (N_5045,N_3158,N_3457);
or U5046 (N_5046,N_3319,N_4276);
nor U5047 (N_5047,N_3411,N_4541);
or U5048 (N_5048,N_4794,N_3382);
or U5049 (N_5049,N_4547,N_3625);
nor U5050 (N_5050,N_2529,N_4181);
and U5051 (N_5051,N_4269,N_2769);
nand U5052 (N_5052,N_3378,N_3497);
and U5053 (N_5053,N_3920,N_4713);
or U5054 (N_5054,N_3181,N_3691);
nor U5055 (N_5055,N_2831,N_2576);
nand U5056 (N_5056,N_3185,N_2640);
and U5057 (N_5057,N_2781,N_4785);
and U5058 (N_5058,N_3551,N_4485);
and U5059 (N_5059,N_3720,N_4873);
nand U5060 (N_5060,N_3039,N_3221);
or U5061 (N_5061,N_4807,N_2903);
nand U5062 (N_5062,N_2731,N_4047);
or U5063 (N_5063,N_2509,N_4717);
or U5064 (N_5064,N_4401,N_4599);
nor U5065 (N_5065,N_3169,N_3024);
nand U5066 (N_5066,N_2856,N_3211);
nor U5067 (N_5067,N_4951,N_4611);
and U5068 (N_5068,N_4224,N_4238);
nand U5069 (N_5069,N_3495,N_2837);
nand U5070 (N_5070,N_3503,N_4701);
or U5071 (N_5071,N_3980,N_4075);
nand U5072 (N_5072,N_3512,N_4558);
nor U5073 (N_5073,N_4818,N_4865);
nand U5074 (N_5074,N_3377,N_4275);
or U5075 (N_5075,N_4350,N_4149);
nor U5076 (N_5076,N_4716,N_2808);
nor U5077 (N_5077,N_3525,N_4755);
and U5078 (N_5078,N_4067,N_3687);
and U5079 (N_5079,N_2566,N_4175);
and U5080 (N_5080,N_4658,N_3363);
nand U5081 (N_5081,N_2852,N_4916);
nor U5082 (N_5082,N_3147,N_3170);
or U5083 (N_5083,N_4513,N_2686);
and U5084 (N_5084,N_4893,N_4992);
nor U5085 (N_5085,N_4407,N_3199);
nor U5086 (N_5086,N_2627,N_2581);
and U5087 (N_5087,N_2921,N_2667);
and U5088 (N_5088,N_3736,N_2613);
nor U5089 (N_5089,N_2884,N_2910);
xnor U5090 (N_5090,N_4791,N_2963);
and U5091 (N_5091,N_4301,N_3735);
or U5092 (N_5092,N_2680,N_4862);
nor U5093 (N_5093,N_2958,N_2950);
and U5094 (N_5094,N_4180,N_2524);
nor U5095 (N_5095,N_4753,N_4241);
or U5096 (N_5096,N_4489,N_3586);
and U5097 (N_5097,N_2805,N_3047);
and U5098 (N_5098,N_4434,N_4102);
nor U5099 (N_5099,N_2612,N_3642);
nand U5100 (N_5100,N_4176,N_4838);
or U5101 (N_5101,N_4897,N_4405);
nand U5102 (N_5102,N_3204,N_2766);
or U5103 (N_5103,N_4570,N_4194);
and U5104 (N_5104,N_4053,N_3316);
or U5105 (N_5105,N_3385,N_2821);
nand U5106 (N_5106,N_4955,N_4508);
or U5107 (N_5107,N_3435,N_3746);
nand U5108 (N_5108,N_4004,N_4303);
nor U5109 (N_5109,N_3544,N_3538);
nor U5110 (N_5110,N_2634,N_4414);
nand U5111 (N_5111,N_2711,N_2625);
nand U5112 (N_5112,N_4647,N_2696);
nand U5113 (N_5113,N_4934,N_4305);
nor U5114 (N_5114,N_4298,N_3037);
nor U5115 (N_5115,N_4686,N_2671);
or U5116 (N_5116,N_4142,N_3130);
nand U5117 (N_5117,N_3429,N_3781);
and U5118 (N_5118,N_2543,N_4913);
and U5119 (N_5119,N_4465,N_3419);
and U5120 (N_5120,N_2632,N_4619);
nand U5121 (N_5121,N_3452,N_4145);
and U5122 (N_5122,N_3422,N_4582);
or U5123 (N_5123,N_3985,N_3794);
or U5124 (N_5124,N_4498,N_3844);
nand U5125 (N_5125,N_2530,N_4923);
nor U5126 (N_5126,N_4363,N_4560);
nor U5127 (N_5127,N_2550,N_4097);
or U5128 (N_5128,N_4831,N_2836);
and U5129 (N_5129,N_3105,N_3099);
or U5130 (N_5130,N_2771,N_4025);
nor U5131 (N_5131,N_2752,N_3554);
and U5132 (N_5132,N_4958,N_3004);
nor U5133 (N_5133,N_2712,N_4747);
or U5134 (N_5134,N_2739,N_4861);
or U5135 (N_5135,N_4491,N_4826);
and U5136 (N_5136,N_2508,N_4054);
or U5137 (N_5137,N_4210,N_2853);
nand U5138 (N_5138,N_2652,N_4191);
nand U5139 (N_5139,N_4902,N_3884);
nand U5140 (N_5140,N_2924,N_4795);
nor U5141 (N_5141,N_2516,N_3662);
or U5142 (N_5142,N_3937,N_3798);
or U5143 (N_5143,N_3804,N_3230);
and U5144 (N_5144,N_4628,N_2518);
or U5145 (N_5145,N_4799,N_4250);
nand U5146 (N_5146,N_4484,N_4711);
and U5147 (N_5147,N_4815,N_3144);
nand U5148 (N_5148,N_4474,N_4788);
nand U5149 (N_5149,N_3982,N_3095);
nor U5150 (N_5150,N_2784,N_3548);
and U5151 (N_5151,N_2570,N_2879);
or U5152 (N_5152,N_3823,N_3400);
or U5153 (N_5153,N_2925,N_3897);
or U5154 (N_5154,N_3567,N_4131);
nand U5155 (N_5155,N_3228,N_3759);
and U5156 (N_5156,N_4256,N_3040);
xor U5157 (N_5157,N_3895,N_3682);
nand U5158 (N_5158,N_2504,N_3660);
nand U5159 (N_5159,N_4760,N_4273);
nor U5160 (N_5160,N_2964,N_4199);
or U5161 (N_5161,N_4302,N_2913);
nor U5162 (N_5162,N_2944,N_3123);
nand U5163 (N_5163,N_4983,N_2569);
nand U5164 (N_5164,N_3649,N_4700);
xnor U5165 (N_5165,N_3530,N_3549);
and U5166 (N_5166,N_4394,N_2607);
or U5167 (N_5167,N_3025,N_3570);
nor U5168 (N_5168,N_2567,N_2692);
nor U5169 (N_5169,N_3755,N_3151);
nand U5170 (N_5170,N_4036,N_2626);
nor U5171 (N_5171,N_4463,N_3420);
or U5172 (N_5172,N_4178,N_4659);
or U5173 (N_5173,N_3472,N_3241);
nand U5174 (N_5174,N_4362,N_4002);
nand U5175 (N_5175,N_4042,N_4315);
and U5176 (N_5176,N_3838,N_2773);
and U5177 (N_5177,N_2742,N_3486);
or U5178 (N_5178,N_4398,N_3878);
and U5179 (N_5179,N_4821,N_3796);
nand U5180 (N_5180,N_3775,N_4011);
nand U5181 (N_5181,N_2644,N_2770);
or U5182 (N_5182,N_3783,N_2843);
nor U5183 (N_5183,N_4268,N_2698);
or U5184 (N_5184,N_4767,N_3565);
nand U5185 (N_5185,N_3141,N_3580);
and U5186 (N_5186,N_3455,N_2936);
and U5187 (N_5187,N_2892,N_4429);
nor U5188 (N_5188,N_4566,N_4384);
nand U5189 (N_5189,N_3762,N_2734);
or U5190 (N_5190,N_3882,N_2973);
nand U5191 (N_5191,N_2719,N_4460);
and U5192 (N_5192,N_4390,N_4473);
or U5193 (N_5193,N_3664,N_2732);
and U5194 (N_5194,N_4410,N_3673);
nor U5195 (N_5195,N_2617,N_4446);
or U5196 (N_5196,N_3208,N_4827);
nor U5197 (N_5197,N_4741,N_4775);
nand U5198 (N_5198,N_3350,N_4855);
and U5199 (N_5199,N_3591,N_3871);
nand U5200 (N_5200,N_4493,N_3029);
and U5201 (N_5201,N_4286,N_2717);
nor U5202 (N_5202,N_3913,N_3957);
and U5203 (N_5203,N_4027,N_3252);
nor U5204 (N_5204,N_4117,N_4228);
nand U5205 (N_5205,N_2738,N_2583);
nand U5206 (N_5206,N_3653,N_3550);
nor U5207 (N_5207,N_4031,N_4721);
nand U5208 (N_5208,N_4453,N_2825);
and U5209 (N_5209,N_3621,N_3295);
or U5210 (N_5210,N_2592,N_3191);
nand U5211 (N_5211,N_4311,N_2914);
and U5212 (N_5212,N_2544,N_3930);
and U5213 (N_5213,N_4341,N_4735);
xor U5214 (N_5214,N_4642,N_3842);
and U5215 (N_5215,N_4352,N_2793);
or U5216 (N_5216,N_2867,N_4921);
nor U5217 (N_5217,N_3068,N_3715);
and U5218 (N_5218,N_4919,N_3259);
and U5219 (N_5219,N_3212,N_3134);
or U5220 (N_5220,N_2728,N_3639);
nor U5221 (N_5221,N_2556,N_3724);
nor U5222 (N_5222,N_3744,N_2685);
nor U5223 (N_5223,N_2540,N_2977);
or U5224 (N_5224,N_4615,N_2900);
or U5225 (N_5225,N_4545,N_3635);
and U5226 (N_5226,N_4602,N_2662);
or U5227 (N_5227,N_4532,N_2941);
nand U5228 (N_5228,N_3206,N_3557);
nand U5229 (N_5229,N_3949,N_2703);
or U5230 (N_5230,N_4070,N_4511);
nand U5231 (N_5231,N_3761,N_3137);
or U5232 (N_5232,N_4132,N_2896);
xor U5233 (N_5233,N_3482,N_4556);
and U5234 (N_5234,N_4395,N_4552);
nand U5235 (N_5235,N_4282,N_3006);
xor U5236 (N_5236,N_2737,N_3611);
nor U5237 (N_5237,N_3873,N_4739);
nor U5238 (N_5238,N_3771,N_2653);
nor U5239 (N_5239,N_3726,N_3041);
nor U5240 (N_5240,N_4078,N_2800);
or U5241 (N_5241,N_3089,N_4480);
nor U5242 (N_5242,N_2639,N_3942);
or U5243 (N_5243,N_4008,N_3166);
or U5244 (N_5244,N_3995,N_3877);
or U5245 (N_5245,N_4840,N_3469);
and U5246 (N_5246,N_3142,N_3303);
nor U5247 (N_5247,N_4317,N_4099);
nand U5248 (N_5248,N_4148,N_3159);
or U5249 (N_5249,N_3383,N_4306);
and U5250 (N_5250,N_3836,N_2503);
nor U5251 (N_5251,N_3829,N_3542);
nor U5252 (N_5252,N_4287,N_4147);
and U5253 (N_5253,N_4366,N_3915);
nand U5254 (N_5254,N_3533,N_3674);
nor U5255 (N_5255,N_4666,N_4839);
nor U5256 (N_5256,N_3659,N_3427);
nor U5257 (N_5257,N_4391,N_2594);
nand U5258 (N_5258,N_3731,N_4722);
or U5259 (N_5259,N_3136,N_3856);
or U5260 (N_5260,N_3623,N_4980);
or U5261 (N_5261,N_4910,N_4853);
nand U5262 (N_5262,N_3404,N_4165);
or U5263 (N_5263,N_3850,N_4884);
and U5264 (N_5264,N_3911,N_4533);
or U5265 (N_5265,N_3669,N_4066);
nand U5266 (N_5266,N_3793,N_4709);
and U5267 (N_5267,N_3729,N_3690);
and U5268 (N_5268,N_3833,N_3791);
nand U5269 (N_5269,N_3593,N_4470);
nand U5270 (N_5270,N_2995,N_3568);
and U5271 (N_5271,N_4968,N_4046);
and U5272 (N_5272,N_3925,N_4657);
nor U5273 (N_5273,N_3063,N_2889);
nand U5274 (N_5274,N_3663,N_4925);
and U5275 (N_5275,N_4805,N_2933);
and U5276 (N_5276,N_4631,N_4850);
and U5277 (N_5277,N_4417,N_4325);
nor U5278 (N_5278,N_4898,N_4613);
or U5279 (N_5279,N_4503,N_4639);
or U5280 (N_5280,N_4814,N_4842);
nand U5281 (N_5281,N_3408,N_2561);
xor U5282 (N_5282,N_4705,N_4320);
nand U5283 (N_5283,N_2762,N_3862);
nand U5284 (N_5284,N_4707,N_3706);
and U5285 (N_5285,N_2539,N_4490);
and U5286 (N_5286,N_4653,N_4291);
nor U5287 (N_5287,N_3604,N_4801);
and U5288 (N_5288,N_2693,N_4632);
and U5289 (N_5289,N_3656,N_4454);
and U5290 (N_5290,N_4107,N_4817);
and U5291 (N_5291,N_3526,N_4595);
nor U5292 (N_5292,N_4745,N_4096);
nand U5293 (N_5293,N_2733,N_4494);
or U5294 (N_5294,N_2674,N_2729);
xnor U5295 (N_5295,N_3943,N_2785);
nand U5296 (N_5296,N_4931,N_3092);
nand U5297 (N_5297,N_3225,N_4420);
and U5298 (N_5298,N_4901,N_3011);
nand U5299 (N_5299,N_4984,N_4051);
nand U5300 (N_5300,N_4048,N_3727);
nor U5301 (N_5301,N_4572,N_4123);
nor U5302 (N_5302,N_4664,N_4907);
or U5303 (N_5303,N_2931,N_3750);
and U5304 (N_5304,N_4157,N_3492);
or U5305 (N_5305,N_4962,N_4618);
nand U5306 (N_5306,N_3412,N_4918);
xnor U5307 (N_5307,N_2595,N_4086);
nor U5308 (N_5308,N_3242,N_4056);
or U5309 (N_5309,N_3666,N_3197);
xnor U5310 (N_5310,N_3962,N_4516);
or U5311 (N_5311,N_3959,N_3442);
or U5312 (N_5312,N_3116,N_4633);
nor U5313 (N_5313,N_2599,N_3232);
nand U5314 (N_5314,N_3299,N_4424);
nor U5315 (N_5315,N_4397,N_3509);
or U5316 (N_5316,N_2943,N_4988);
nor U5317 (N_5317,N_2983,N_3483);
nor U5318 (N_5318,N_3093,N_4612);
or U5319 (N_5319,N_2809,N_4675);
nor U5320 (N_5320,N_2735,N_4034);
nor U5321 (N_5321,N_3868,N_3624);
and U5322 (N_5322,N_3852,N_3531);
or U5323 (N_5323,N_3179,N_3956);
nor U5324 (N_5324,N_4010,N_4607);
and U5325 (N_5325,N_3254,N_2803);
nor U5326 (N_5326,N_4360,N_3325);
or U5327 (N_5327,N_4020,N_3756);
nor U5328 (N_5328,N_3900,N_4720);
nor U5329 (N_5329,N_4321,N_3450);
and U5330 (N_5330,N_2597,N_3880);
or U5331 (N_5331,N_4019,N_2624);
nand U5332 (N_5332,N_3692,N_2756);
or U5333 (N_5333,N_4527,N_4637);
nand U5334 (N_5334,N_3365,N_3370);
nand U5335 (N_5335,N_4579,N_4076);
or U5336 (N_5336,N_4662,N_4935);
nor U5337 (N_5337,N_3436,N_4906);
nor U5338 (N_5338,N_2513,N_4543);
and U5339 (N_5339,N_2591,N_3012);
or U5340 (N_5340,N_3261,N_3167);
and U5341 (N_5341,N_3425,N_4433);
nand U5342 (N_5342,N_4049,N_2507);
nor U5343 (N_5343,N_4982,N_4752);
and U5344 (N_5344,N_4385,N_3332);
nor U5345 (N_5345,N_3392,N_4003);
nand U5346 (N_5346,N_3818,N_2901);
nand U5347 (N_5347,N_3018,N_4787);
nor U5348 (N_5348,N_4243,N_3488);
nor U5349 (N_5349,N_2826,N_4186);
nand U5350 (N_5350,N_2954,N_3284);
nor U5351 (N_5351,N_2932,N_3806);
and U5352 (N_5352,N_2801,N_3080);
nor U5353 (N_5353,N_3263,N_3015);
or U5354 (N_5354,N_2861,N_3990);
and U5355 (N_5355,N_3875,N_3300);
nor U5356 (N_5356,N_2600,N_3367);
or U5357 (N_5357,N_3327,N_2527);
and U5358 (N_5358,N_4277,N_3313);
nor U5359 (N_5359,N_4316,N_4604);
nor U5360 (N_5360,N_3288,N_4173);
and U5361 (N_5361,N_3282,N_3894);
nand U5362 (N_5362,N_3599,N_3824);
and U5363 (N_5363,N_4835,N_3369);
nand U5364 (N_5364,N_2811,N_4509);
nand U5365 (N_5365,N_4355,N_3305);
nor U5366 (N_5366,N_3951,N_4155);
and U5367 (N_5367,N_4712,N_3700);
or U5368 (N_5368,N_3825,N_2895);
and U5369 (N_5369,N_4105,N_2955);
and U5370 (N_5370,N_3904,N_4023);
nor U5371 (N_5371,N_4009,N_2708);
nor U5372 (N_5372,N_4314,N_2962);
nor U5373 (N_5373,N_3391,N_3402);
nand U5374 (N_5374,N_2928,N_4259);
nor U5375 (N_5375,N_4342,N_3397);
nand U5376 (N_5376,N_2528,N_2730);
nor U5377 (N_5377,N_3657,N_3201);
and U5378 (N_5378,N_3444,N_4333);
nor U5379 (N_5379,N_3885,N_3924);
nor U5380 (N_5380,N_4515,N_2578);
or U5381 (N_5381,N_4945,N_3065);
or U5382 (N_5382,N_2888,N_4072);
or U5383 (N_5383,N_3036,N_3493);
xnor U5384 (N_5384,N_4285,N_4679);
or U5385 (N_5385,N_4144,N_4685);
and U5386 (N_5386,N_4134,N_2501);
nand U5387 (N_5387,N_2799,N_4156);
nor U5388 (N_5388,N_4636,N_4589);
and U5389 (N_5389,N_4338,N_3008);
nor U5390 (N_5390,N_4696,N_2782);
nor U5391 (N_5391,N_3869,N_4880);
nand U5392 (N_5392,N_2628,N_4265);
or U5393 (N_5393,N_3117,N_3893);
nand U5394 (N_5394,N_3845,N_4294);
nor U5395 (N_5395,N_3891,N_4202);
and U5396 (N_5396,N_4064,N_2618);
or U5397 (N_5397,N_3209,N_2870);
or U5398 (N_5398,N_4239,N_3789);
or U5399 (N_5399,N_4792,N_3222);
nor U5400 (N_5400,N_4264,N_3976);
nand U5401 (N_5401,N_3707,N_4488);
or U5402 (N_5402,N_4112,N_4284);
or U5403 (N_5403,N_2525,N_4396);
xnor U5404 (N_5404,N_4762,N_3342);
nand U5405 (N_5405,N_4954,N_4479);
xor U5406 (N_5406,N_2679,N_3172);
or U5407 (N_5407,N_4847,N_2827);
and U5408 (N_5408,N_3398,N_4029);
nand U5409 (N_5409,N_2606,N_3139);
nor U5410 (N_5410,N_3505,N_4649);
nand U5411 (N_5411,N_2650,N_3262);
and U5412 (N_5412,N_4368,N_3860);
or U5413 (N_5413,N_4403,N_2790);
or U5414 (N_5414,N_3401,N_3795);
and U5415 (N_5415,N_2796,N_3237);
nand U5416 (N_5416,N_2706,N_2621);
nor U5417 (N_5417,N_4793,N_3952);
or U5418 (N_5418,N_3267,N_4167);
and U5419 (N_5419,N_4914,N_2795);
or U5420 (N_5420,N_4236,N_3078);
nor U5421 (N_5421,N_2960,N_3210);
and U5422 (N_5422,N_3612,N_3536);
or U5423 (N_5423,N_3464,N_3413);
or U5424 (N_5424,N_4704,N_4677);
nor U5425 (N_5425,N_2683,N_2854);
and U5426 (N_5426,N_3758,N_4482);
nor U5427 (N_5427,N_3133,N_2786);
or U5428 (N_5428,N_2992,N_4654);
nand U5429 (N_5429,N_2596,N_3590);
nor U5430 (N_5430,N_4266,N_4601);
or U5431 (N_5431,N_4946,N_4377);
xnor U5432 (N_5432,N_3641,N_4136);
or U5433 (N_5433,N_3349,N_3932);
nor U5434 (N_5434,N_4040,N_4790);
nor U5435 (N_5435,N_4220,N_4889);
nor U5436 (N_5436,N_4229,N_4756);
nand U5437 (N_5437,N_4581,N_3043);
or U5438 (N_5438,N_3033,N_2834);
nor U5439 (N_5439,N_3922,N_4727);
nand U5440 (N_5440,N_3049,N_4692);
and U5441 (N_5441,N_4211,N_2601);
xor U5442 (N_5442,N_3532,N_4726);
and U5443 (N_5443,N_3311,N_3613);
and U5444 (N_5444,N_3713,N_3514);
nand U5445 (N_5445,N_4903,N_3596);
nand U5446 (N_5446,N_4358,N_3161);
and U5447 (N_5447,N_4523,N_4388);
nor U5448 (N_5448,N_3394,N_3372);
or U5449 (N_5449,N_2763,N_3010);
or U5450 (N_5450,N_3622,N_3966);
or U5451 (N_5451,N_4304,N_2912);
or U5452 (N_5452,N_3857,N_4213);
xnor U5453 (N_5453,N_4845,N_4870);
nand U5454 (N_5454,N_4118,N_4772);
and U5455 (N_5455,N_4339,N_2844);
nor U5456 (N_5456,N_3615,N_3091);
or U5457 (N_5457,N_4452,N_2982);
or U5458 (N_5458,N_2687,N_2658);
and U5459 (N_5459,N_3384,N_4006);
or U5460 (N_5460,N_3986,N_3338);
nand U5461 (N_5461,N_3847,N_3745);
or U5462 (N_5462,N_3689,N_4693);
nor U5463 (N_5463,N_3057,N_3048);
nand U5464 (N_5464,N_2929,N_3090);
nand U5465 (N_5465,N_4018,N_4977);
and U5466 (N_5466,N_3719,N_2542);
nand U5467 (N_5467,N_3646,N_3344);
and U5468 (N_5468,N_4715,N_2757);
nand U5469 (N_5469,N_4776,N_4087);
and U5470 (N_5470,N_3522,N_4697);
and U5471 (N_5471,N_3837,N_3907);
nand U5472 (N_5472,N_2598,N_2532);
nand U5473 (N_5473,N_3638,N_3619);
xnor U5474 (N_5474,N_2707,N_4719);
and U5475 (N_5475,N_4426,N_3023);
nand U5476 (N_5476,N_3410,N_3126);
nand U5477 (N_5477,N_4917,N_2715);
nand U5478 (N_5478,N_2819,N_3120);
and U5479 (N_5479,N_4904,N_3513);
or U5480 (N_5480,N_3009,N_4415);
or U5481 (N_5481,N_4400,N_2897);
and U5482 (N_5482,N_3220,N_3343);
and U5483 (N_5483,N_3165,N_4379);
nand U5484 (N_5484,N_4000,N_4499);
or U5485 (N_5485,N_3461,N_2688);
or U5486 (N_5486,N_2765,N_3407);
nand U5487 (N_5487,N_3406,N_4896);
nand U5488 (N_5488,N_3840,N_4800);
nor U5489 (N_5489,N_3358,N_2909);
nor U5490 (N_5490,N_4703,N_4583);
nor U5491 (N_5491,N_4640,N_2710);
and U5492 (N_5492,N_4214,N_3815);
or U5493 (N_5493,N_3138,N_4455);
or U5494 (N_5494,N_4439,N_4088);
and U5495 (N_5495,N_2871,N_3680);
or U5496 (N_5496,N_4723,N_4872);
and U5497 (N_5497,N_4179,N_2629);
or U5498 (N_5498,N_3712,N_3676);
or U5499 (N_5499,N_2838,N_3923);
nor U5500 (N_5500,N_3180,N_4383);
or U5501 (N_5501,N_4381,N_2575);
and U5502 (N_5502,N_4106,N_4376);
and U5503 (N_5503,N_3598,N_2672);
nor U5504 (N_5504,N_2622,N_2949);
nor U5505 (N_5505,N_4329,N_3552);
nand U5506 (N_5506,N_3571,N_3792);
or U5507 (N_5507,N_4517,N_3480);
nand U5508 (N_5508,N_3742,N_2969);
or U5509 (N_5509,N_3801,N_3709);
or U5510 (N_5510,N_2894,N_3569);
nand U5511 (N_5511,N_4367,N_3948);
nand U5512 (N_5512,N_2610,N_3087);
nand U5513 (N_5513,N_3696,N_3308);
and U5514 (N_5514,N_2651,N_4706);
nor U5515 (N_5515,N_4330,N_3826);
nor U5516 (N_5516,N_2723,N_4996);
nand U5517 (N_5517,N_4478,N_4153);
nand U5518 (N_5518,N_4413,N_2593);
nand U5519 (N_5519,N_2947,N_2887);
nand U5520 (N_5520,N_4596,N_3717);
or U5521 (N_5521,N_4820,N_4978);
nor U5522 (N_5522,N_4578,N_3684);
xor U5523 (N_5523,N_3634,N_4976);
nor U5524 (N_5524,N_3902,N_4504);
nand U5525 (N_5525,N_4169,N_3448);
or U5526 (N_5526,N_4151,N_3654);
nand U5527 (N_5527,N_3511,N_4279);
and U5528 (N_5528,N_4852,N_4183);
nor U5529 (N_5529,N_4714,N_2743);
and U5530 (N_5530,N_4399,N_3035);
and U5531 (N_5531,N_2859,N_4501);
or U5532 (N_5532,N_3207,N_3834);
nand U5533 (N_5533,N_4447,N_3938);
xnor U5534 (N_5534,N_4378,N_2750);
and U5535 (N_5535,N_2695,N_4518);
nand U5536 (N_5536,N_3465,N_4135);
nand U5537 (N_5537,N_4912,N_3058);
nor U5538 (N_5538,N_4467,N_3239);
xor U5539 (N_5539,N_2754,N_3380);
nand U5540 (N_5540,N_4140,N_2505);
and U5541 (N_5541,N_3906,N_4746);
and U5542 (N_5542,N_3438,N_2939);
and U5543 (N_5543,N_4158,N_2705);
nor U5544 (N_5544,N_2946,N_3357);
and U5545 (N_5545,N_4129,N_4028);
and U5546 (N_5546,N_2988,N_2971);
nor U5547 (N_5547,N_3921,N_4079);
or U5548 (N_5548,N_3636,N_3618);
nor U5549 (N_5549,N_4766,N_4240);
nor U5550 (N_5550,N_4114,N_3453);
and U5551 (N_5551,N_2656,N_4553);
nand U5552 (N_5552,N_3294,N_4882);
nor U5553 (N_5553,N_3044,N_2772);
and U5554 (N_5554,N_4584,N_3240);
or U5555 (N_5555,N_3104,N_3304);
nor U5556 (N_5556,N_3741,N_2893);
nand U5557 (N_5557,N_2828,N_4313);
nand U5558 (N_5558,N_3703,N_3782);
and U5559 (N_5559,N_3246,N_4035);
or U5560 (N_5560,N_2590,N_4895);
and U5561 (N_5561,N_2747,N_3280);
nor U5562 (N_5562,N_4380,N_4887);
nor U5563 (N_5563,N_3386,N_3864);
and U5564 (N_5564,N_3339,N_4590);
nand U5565 (N_5565,N_3335,N_4412);
nor U5566 (N_5566,N_4844,N_4044);
or U5567 (N_5567,N_4819,N_3097);
or U5568 (N_5568,N_4859,N_4953);
and U5569 (N_5569,N_3946,N_4254);
or U5570 (N_5570,N_4091,N_2882);
and U5571 (N_5571,N_3328,N_2713);
nor U5572 (N_5572,N_4749,N_4871);
nor U5573 (N_5573,N_4648,N_4477);
and U5574 (N_5574,N_4353,N_3835);
nor U5575 (N_5575,N_4319,N_4966);
or U5576 (N_5576,N_3146,N_4890);
nor U5577 (N_5577,N_3853,N_4233);
or U5578 (N_5578,N_2906,N_4652);
and U5579 (N_5579,N_2904,N_3079);
nand U5580 (N_5580,N_2744,N_3076);
or U5581 (N_5581,N_4408,N_3471);
nand U5582 (N_5582,N_4610,N_3255);
and U5583 (N_5583,N_3652,N_4856);
nor U5584 (N_5584,N_3321,N_3060);
or U5585 (N_5585,N_2930,N_3905);
or U5586 (N_5586,N_4782,N_3785);
nor U5587 (N_5587,N_4834,N_3389);
xor U5588 (N_5588,N_4765,N_4074);
and U5589 (N_5589,N_4371,N_3426);
nand U5590 (N_5590,N_4617,N_2572);
nor U5591 (N_5591,N_2676,N_3912);
nor U5592 (N_5592,N_2665,N_2993);
or U5593 (N_5593,N_4620,N_4540);
nand U5594 (N_5594,N_4824,N_3874);
and U5595 (N_5595,N_3094,N_2880);
nor U5596 (N_5596,N_3730,N_3725);
and U5597 (N_5597,N_4437,N_2534);
nor U5598 (N_5598,N_4773,N_4216);
or U5599 (N_5599,N_4849,N_4336);
or U5600 (N_5600,N_3975,N_2918);
or U5601 (N_5601,N_4226,N_2701);
and U5602 (N_5602,N_4081,N_4567);
or U5603 (N_5603,N_4128,N_3861);
or U5604 (N_5604,N_3589,N_2751);
or U5605 (N_5605,N_3799,N_4456);
or U5606 (N_5606,N_4592,N_2660);
and U5607 (N_5607,N_4964,N_3474);
nor U5608 (N_5608,N_4323,N_2519);
or U5609 (N_5609,N_3517,N_3190);
or U5610 (N_5610,N_3779,N_4038);
nor U5611 (N_5611,N_3588,N_3416);
nor U5612 (N_5612,N_3100,N_4963);
nand U5613 (N_5613,N_3387,N_2885);
and U5614 (N_5614,N_3988,N_4625);
nor U5615 (N_5615,N_3846,N_3272);
or U5616 (N_5616,N_3200,N_3916);
nor U5617 (N_5617,N_3289,N_3681);
nand U5618 (N_5618,N_3053,N_4139);
or U5619 (N_5619,N_2554,N_4271);
or U5620 (N_5620,N_2538,N_4249);
and U5621 (N_5621,N_4998,N_4113);
and U5622 (N_5622,N_3760,N_3888);
nand U5623 (N_5623,N_3193,N_3809);
or U5624 (N_5624,N_3188,N_2669);
and U5625 (N_5625,N_3989,N_2636);
nand U5626 (N_5626,N_3678,N_3066);
nor U5627 (N_5627,N_3315,N_3213);
and U5628 (N_5628,N_3038,N_2620);
and U5629 (N_5629,N_2546,N_2987);
and U5630 (N_5630,N_4440,N_4416);
and U5631 (N_5631,N_4528,N_3248);
or U5632 (N_5632,N_2881,N_4255);
nor U5633 (N_5633,N_3701,N_4080);
nor U5634 (N_5634,N_3774,N_4823);
nor U5635 (N_5635,N_3125,N_3340);
or U5636 (N_5636,N_3977,N_3476);
or U5637 (N_5637,N_4124,N_3184);
nand U5638 (N_5638,N_3899,N_4937);
nand U5639 (N_5639,N_4663,N_4328);
nor U5640 (N_5640,N_3883,N_2675);
nor U5641 (N_5641,N_3699,N_4660);
or U5642 (N_5642,N_4283,N_3364);
nor U5643 (N_5643,N_3056,N_4851);
nand U5644 (N_5644,N_3898,N_2824);
and U5645 (N_5645,N_2792,N_3573);
and U5646 (N_5646,N_4803,N_2614);
nand U5647 (N_5647,N_3843,N_2535);
nor U5648 (N_5648,N_3249,N_4130);
and U5649 (N_5649,N_4725,N_4492);
nor U5650 (N_5650,N_4212,N_4680);
nand U5651 (N_5651,N_3718,N_3279);
and U5652 (N_5652,N_4986,N_3437);
nor U5653 (N_5653,N_3595,N_3683);
nand U5654 (N_5654,N_3560,N_3747);
and U5655 (N_5655,N_2678,N_4472);
or U5656 (N_5656,N_2648,N_3434);
and U5657 (N_5657,N_3506,N_4205);
or U5658 (N_5658,N_3331,N_4495);
nor U5659 (N_5659,N_3941,N_3061);
or U5660 (N_5660,N_4340,N_4936);
and U5661 (N_5661,N_3148,N_3485);
nand U5662 (N_5662,N_3484,N_3494);
nor U5663 (N_5663,N_3075,N_2619);
nor U5664 (N_5664,N_4026,N_3984);
nor U5665 (N_5665,N_3523,N_4526);
nand U5666 (N_5666,N_4744,N_3168);
nor U5667 (N_5667,N_3784,N_4160);
nor U5668 (N_5668,N_4121,N_2974);
and U5669 (N_5669,N_4092,N_2689);
or U5670 (N_5670,N_3345,N_3566);
nand U5671 (N_5671,N_3154,N_3260);
or U5672 (N_5672,N_3217,N_4634);
or U5673 (N_5673,N_4476,N_4822);
or U5674 (N_5674,N_3238,N_4443);
nor U5675 (N_5675,N_3890,N_3999);
and U5676 (N_5676,N_3667,N_3953);
nand U5677 (N_5677,N_3460,N_4290);
and U5678 (N_5678,N_4846,N_4836);
nand U5679 (N_5679,N_4883,N_3393);
or U5680 (N_5680,N_3524,N_3143);
and U5681 (N_5681,N_2952,N_2646);
nor U5682 (N_5682,N_3302,N_4514);
and U5683 (N_5683,N_3320,N_2980);
and U5684 (N_5684,N_3346,N_3062);
nand U5685 (N_5685,N_4841,N_4292);
or U5686 (N_5686,N_3226,N_4555);
or U5687 (N_5687,N_2740,N_3772);
or U5688 (N_5688,N_3944,N_2515);
nand U5689 (N_5689,N_4886,N_2934);
and U5690 (N_5690,N_4736,N_4406);
and U5691 (N_5691,N_3050,N_3432);
or U5692 (N_5692,N_2965,N_3500);
nor U5693 (N_5693,N_3757,N_4163);
or U5694 (N_5694,N_2850,N_2580);
or U5695 (N_5695,N_4059,N_4939);
and U5696 (N_5696,N_4920,N_3851);
nor U5697 (N_5697,N_2807,N_4177);
and U5698 (N_5698,N_3352,N_3630);
xnor U5699 (N_5699,N_3155,N_3371);
or U5700 (N_5700,N_2681,N_2517);
or U5701 (N_5701,N_4554,N_4689);
nor U5702 (N_5702,N_3521,N_4970);
nor U5703 (N_5703,N_4374,N_3098);
or U5704 (N_5704,N_4187,N_3329);
nand U5705 (N_5705,N_3585,N_4990);
or U5706 (N_5706,N_2975,N_4585);
nand U5707 (N_5707,N_2682,N_4770);
nand U5708 (N_5708,N_3515,N_2873);
xnor U5709 (N_5709,N_4232,N_2978);
and U5710 (N_5710,N_3274,N_3247);
or U5711 (N_5711,N_3537,N_4138);
and U5712 (N_5712,N_4577,N_3318);
nor U5713 (N_5713,N_2531,N_4300);
and U5714 (N_5714,N_4152,N_3229);
nand U5715 (N_5715,N_3414,N_3301);
or U5716 (N_5716,N_3607,N_3695);
nor U5717 (N_5717,N_4780,N_3083);
nand U5718 (N_5718,N_3162,N_4119);
or U5719 (N_5719,N_3661,N_3812);
nor U5720 (N_5720,N_4295,N_4928);
or U5721 (N_5721,N_4364,N_3182);
nand U5722 (N_5722,N_3892,N_3348);
and U5723 (N_5723,N_3013,N_3128);
and U5724 (N_5724,N_3433,N_3616);
nor U5725 (N_5725,N_2858,N_4441);
and U5726 (N_5726,N_3617,N_4933);
or U5727 (N_5727,N_2638,N_3714);
nor U5728 (N_5728,N_3251,N_4534);
nand U5729 (N_5729,N_3983,N_4608);
nand U5730 (N_5730,N_3740,N_4869);
and U5731 (N_5731,N_2536,N_3918);
and U5732 (N_5732,N_4222,N_4586);
or U5733 (N_5733,N_4956,N_3074);
and U5734 (N_5734,N_3016,N_4428);
nand U5735 (N_5735,N_4562,N_2996);
nand U5736 (N_5736,N_2533,N_4324);
nand U5737 (N_5737,N_4068,N_3910);
or U5738 (N_5738,N_3361,N_2832);
nand U5739 (N_5739,N_4600,N_2902);
or U5740 (N_5740,N_2985,N_3914);
nor U5741 (N_5741,N_3849,N_4816);
or U5742 (N_5742,N_2886,N_3769);
nor U5743 (N_5743,N_4524,N_3996);
nor U5744 (N_5744,N_2907,N_4626);
nand U5745 (N_5745,N_3379,N_4603);
and U5746 (N_5746,N_3405,N_4104);
and U5747 (N_5747,N_3766,N_2916);
nor U5748 (N_5748,N_3931,N_4198);
or U5749 (N_5749,N_4924,N_3777);
nand U5750 (N_5750,N_4461,N_4569);
nor U5751 (N_5751,N_4127,N_2923);
nor U5752 (N_5752,N_4234,N_4940);
or U5753 (N_5753,N_4754,N_4184);
and U5754 (N_5754,N_3306,N_3264);
nor U5755 (N_5755,N_4404,N_4039);
or U5756 (N_5756,N_3753,N_3219);
xnor U5757 (N_5757,N_4574,N_3688);
or U5758 (N_5758,N_3119,N_3559);
xor U5759 (N_5759,N_4442,N_3608);
nor U5760 (N_5760,N_2898,N_3196);
or U5761 (N_5761,N_2761,N_3195);
nor U5762 (N_5762,N_3341,N_4166);
nand U5763 (N_5763,N_4806,N_3174);
nor U5764 (N_5764,N_4985,N_2608);
nand U5765 (N_5765,N_4975,N_3244);
nor U5766 (N_5766,N_4231,N_2510);
and U5767 (N_5767,N_4077,N_4459);
or U5768 (N_5768,N_2657,N_3529);
and U5769 (N_5769,N_4591,N_3929);
and U5770 (N_5770,N_3475,N_4651);
nor U5771 (N_5771,N_3708,N_3972);
and U5772 (N_5772,N_2979,N_3702);
or U5773 (N_5773,N_3754,N_2991);
nand U5774 (N_5774,N_3963,N_2851);
nand U5775 (N_5775,N_4671,N_3881);
and U5776 (N_5776,N_2810,N_4571);
or U5777 (N_5777,N_2700,N_2919);
xor U5778 (N_5778,N_4950,N_4262);
nor U5779 (N_5779,N_3581,N_2541);
nor U5780 (N_5780,N_4947,N_3997);
or U5781 (N_5781,N_4559,N_4347);
or U5782 (N_5782,N_4969,N_4309);
xor U5783 (N_5783,N_2605,N_3106);
nor U5784 (N_5784,N_4879,N_3998);
xnor U5785 (N_5785,N_4351,N_3909);
and U5786 (N_5786,N_4133,N_2522);
and U5787 (N_5787,N_3767,N_4257);
nor U5788 (N_5788,N_3131,N_3333);
and U5789 (N_5789,N_3620,N_3848);
nand U5790 (N_5790,N_3291,N_4297);
nand U5791 (N_5791,N_3122,N_3637);
xnor U5792 (N_5792,N_4537,N_2647);
or U5793 (N_5793,N_4742,N_4235);
nand U5794 (N_5794,N_3218,N_3643);
and U5795 (N_5795,N_3234,N_3644);
xor U5796 (N_5796,N_3751,N_4561);
or U5797 (N_5797,N_3353,N_4055);
xnor U5798 (N_5798,N_2780,N_3069);
nand U5799 (N_5799,N_3816,N_3665);
or U5800 (N_5800,N_4345,N_4743);
or U5801 (N_5801,N_4959,N_4941);
nand U5802 (N_5802,N_4288,N_4758);
and U5803 (N_5803,N_3787,N_3132);
and U5804 (N_5804,N_3610,N_4280);
nand U5805 (N_5805,N_4458,N_4449);
nand U5806 (N_5806,N_4359,N_4798);
nand U5807 (N_5807,N_3728,N_2745);
or U5808 (N_5808,N_3430,N_2664);
or U5809 (N_5809,N_3192,N_3648);
or U5810 (N_5810,N_4965,N_2564);
nor U5811 (N_5811,N_2736,N_4774);
and U5812 (N_5812,N_3748,N_3285);
or U5813 (N_5813,N_3424,N_4245);
nor U5814 (N_5814,N_3070,N_4926);
nor U5815 (N_5815,N_4519,N_4674);
nand U5816 (N_5816,N_2846,N_3449);
nand U5817 (N_5817,N_3820,N_4759);
or U5818 (N_5818,N_2927,N_3711);
or U5819 (N_5819,N_4888,N_3498);
nand U5820 (N_5820,N_3045,N_3113);
and U5821 (N_5821,N_4892,N_4858);
or U5822 (N_5822,N_4681,N_3231);
or U5823 (N_5823,N_3003,N_3463);
and U5824 (N_5824,N_3790,N_3286);
and U5825 (N_5825,N_3632,N_4605);
and U5826 (N_5826,N_4237,N_3153);
or U5827 (N_5827,N_3290,N_4337);
or U5828 (N_5828,N_4549,N_3431);
nand U5829 (N_5829,N_4083,N_3001);
nand U5830 (N_5830,N_4738,N_3749);
and U5831 (N_5831,N_4781,N_3415);
nand U5832 (N_5832,N_4307,N_3487);
and U5833 (N_5833,N_4260,N_4981);
or U5834 (N_5834,N_3390,N_4682);
or U5835 (N_5835,N_4991,N_3114);
and U5836 (N_5836,N_2956,N_4521);
or U5837 (N_5837,N_4457,N_4171);
nand U5838 (N_5838,N_4621,N_2957);
and U5839 (N_5839,N_4354,N_4927);
xnor U5840 (N_5840,N_3723,N_3479);
or U5841 (N_5841,N_3178,N_4073);
nand U5842 (N_5842,N_2998,N_4737);
nor U5843 (N_5843,N_2999,N_4375);
and U5844 (N_5844,N_4938,N_2970);
nand U5845 (N_5845,N_4708,N_3115);
nand U5846 (N_5846,N_2573,N_4357);
or U5847 (N_5847,N_3547,N_4084);
and U5848 (N_5848,N_2864,N_3032);
and U5849 (N_5849,N_3870,N_4695);
or U5850 (N_5850,N_2654,N_2691);
nor U5851 (N_5851,N_3149,N_3121);
nand U5852 (N_5852,N_3813,N_4530);
and U5853 (N_5853,N_3005,N_4761);
nand U5854 (N_5854,N_4419,N_3160);
xor U5855 (N_5855,N_4462,N_3704);
nand U5856 (N_5856,N_3293,N_3046);
or U5857 (N_5857,N_2899,N_3067);
nor U5858 (N_5858,N_4779,N_2523);
and U5859 (N_5859,N_3275,N_3827);
or U5860 (N_5860,N_2783,N_3283);
or U5861 (N_5861,N_4251,N_4911);
nand U5862 (N_5862,N_3403,N_3734);
nor U5863 (N_5863,N_3578,N_2951);
and U5864 (N_5864,N_2755,N_3323);
xor U5865 (N_5865,N_3467,N_4289);
xor U5866 (N_5866,N_4045,N_3867);
nand U5867 (N_5867,N_4863,N_2830);
and U5868 (N_5868,N_2545,N_2500);
and U5869 (N_5869,N_4189,N_4225);
or U5870 (N_5870,N_3694,N_3518);
or U5871 (N_5871,N_3510,N_4525);
nor U5872 (N_5872,N_4594,N_3428);
or U5873 (N_5873,N_4094,N_3101);
nor U5874 (N_5874,N_2817,N_4763);
or U5875 (N_5875,N_2915,N_4797);
nand U5876 (N_5876,N_4141,N_4071);
or U5877 (N_5877,N_2702,N_4546);
nand U5878 (N_5878,N_3235,N_3445);
nand U5879 (N_5879,N_4825,N_4694);
or U5880 (N_5880,N_3807,N_4900);
and U5881 (N_5881,N_4563,N_4597);
or U5882 (N_5882,N_4430,N_2875);
nor U5883 (N_5883,N_4669,N_2659);
nand U5884 (N_5884,N_4857,N_4204);
and U5885 (N_5885,N_2718,N_2990);
or U5886 (N_5886,N_3330,N_4170);
nor U5887 (N_5887,N_3421,N_2549);
and U5888 (N_5888,N_3954,N_3778);
nor U5889 (N_5889,N_4987,N_3839);
nand U5890 (N_5890,N_4973,N_3176);
nor U5891 (N_5891,N_4550,N_3609);
or U5892 (N_5892,N_4629,N_3227);
or U5893 (N_5893,N_4464,N_2720);
nor U5894 (N_5894,N_4221,N_3042);
nor U5895 (N_5895,N_4668,N_4500);
and U5896 (N_5896,N_4522,N_3626);
and U5897 (N_5897,N_4370,N_3614);
and U5898 (N_5898,N_3447,N_4813);
nor U5899 (N_5899,N_3451,N_2883);
and U5900 (N_5900,N_3215,N_4905);
nand U5901 (N_5901,N_4944,N_3102);
and U5902 (N_5902,N_2926,N_2582);
and U5903 (N_5903,N_4548,N_4771);
nor U5904 (N_5904,N_2981,N_2778);
and U5905 (N_5905,N_3919,N_3297);
nor U5906 (N_5906,N_3183,N_2868);
nor U5907 (N_5907,N_3064,N_3606);
or U5908 (N_5908,N_2794,N_3908);
nand U5909 (N_5909,N_3872,N_3958);
or U5910 (N_5910,N_4874,N_4673);
and U5911 (N_5911,N_3939,N_4203);
or U5912 (N_5912,N_3583,N_2604);
nand U5913 (N_5913,N_4310,N_3322);
nand U5914 (N_5914,N_2942,N_3527);
nand U5915 (N_5915,N_4829,N_4050);
nor U5916 (N_5916,N_4622,N_3111);
and U5917 (N_5917,N_4278,N_3356);
nor U5918 (N_5918,N_3296,N_3059);
and U5919 (N_5919,N_3555,N_4082);
and U5920 (N_5920,N_3693,N_3592);
and U5921 (N_5921,N_4676,N_4638);
and U5922 (N_5922,N_2753,N_4614);
or U5923 (N_5923,N_3677,N_3640);
or U5924 (N_5924,N_4327,N_3672);
xor U5925 (N_5925,N_2822,N_2789);
or U5926 (N_5926,N_3470,N_4751);
nand U5927 (N_5927,N_4520,N_4687);
nand U5928 (N_5928,N_3633,N_2855);
nor U5929 (N_5929,N_4270,N_4219);
nor U5930 (N_5930,N_4001,N_4387);
or U5931 (N_5931,N_3519,N_3520);
and U5932 (N_5932,N_3584,N_2989);
nand U5933 (N_5933,N_2661,N_4974);
nor U5934 (N_5934,N_4258,N_4365);
nand U5935 (N_5935,N_3508,N_3456);
xnor U5936 (N_5936,N_4999,N_3124);
or U5937 (N_5937,N_3458,N_3462);
or U5938 (N_5938,N_3164,N_2635);
or U5939 (N_5939,N_3175,N_4409);
nor U5940 (N_5940,N_3800,N_4778);
nand U5941 (N_5941,N_4789,N_4217);
nor U5942 (N_5942,N_3575,N_2842);
nor U5943 (N_5943,N_4860,N_4348);
nor U5944 (N_5944,N_2615,N_3546);
or U5945 (N_5945,N_2841,N_4101);
xnor U5946 (N_5946,N_3697,N_4728);
nand U5947 (N_5947,N_3841,N_4207);
or U5948 (N_5948,N_3651,N_4786);
or U5949 (N_5949,N_3171,N_4272);
nor U5950 (N_5950,N_4103,N_4724);
nand U5951 (N_5951,N_3650,N_4089);
and U5952 (N_5952,N_2551,N_3927);
nor U5953 (N_5953,N_4192,N_3945);
and U5954 (N_5954,N_2768,N_3969);
or U5955 (N_5955,N_2759,N_4223);
nor U5956 (N_5956,N_2722,N_4932);
nor U5957 (N_5957,N_4909,N_3376);
or U5958 (N_5958,N_4007,N_2802);
or U5959 (N_5959,N_3802,N_3088);
and U5960 (N_5960,N_3271,N_4043);
and U5961 (N_5961,N_2609,N_4110);
or U5962 (N_5962,N_2727,N_2940);
nand U5963 (N_5963,N_3491,N_4698);
or U5964 (N_5964,N_4769,N_3597);
and U5965 (N_5965,N_3355,N_3504);
nor U5966 (N_5966,N_4161,N_4188);
nand U5967 (N_5967,N_3886,N_2643);
nor U5968 (N_5968,N_4740,N_4557);
nor U5969 (N_5969,N_4536,N_2767);
or U5970 (N_5970,N_4014,N_4098);
and U5971 (N_5971,N_3317,N_2537);
nand U5972 (N_5972,N_4580,N_4242);
nand U5973 (N_5973,N_4878,N_3994);
and U5974 (N_5974,N_4154,N_4971);
and U5975 (N_5975,N_4326,N_3698);
or U5976 (N_5976,N_3324,N_3933);
or U5977 (N_5977,N_2917,N_4565);
or U5978 (N_5978,N_2829,N_3214);
or U5979 (N_5979,N_2813,N_3256);
nand U5980 (N_5980,N_4576,N_2869);
and U5981 (N_5981,N_2557,N_2804);
and U5982 (N_5982,N_3628,N_4750);
and U5983 (N_5983,N_3031,N_3780);
and U5984 (N_5984,N_4868,N_3096);
nor U5985 (N_5985,N_3764,N_3854);
nand U5986 (N_5986,N_2959,N_3177);
or U5987 (N_5987,N_2876,N_2777);
nor U5988 (N_5988,N_4281,N_4218);
and U5989 (N_5989,N_4812,N_4891);
and U5990 (N_5990,N_4466,N_2797);
and U5991 (N_5991,N_4372,N_4875);
or U5992 (N_5992,N_2994,N_3901);
nor U5993 (N_5993,N_3528,N_4373);
or U5994 (N_5994,N_3675,N_3961);
or U5995 (N_5995,N_3722,N_4248);
and U5996 (N_5996,N_2511,N_4299);
or U5997 (N_5997,N_4432,N_4115);
nor U5998 (N_5998,N_3935,N_3819);
nand U5999 (N_5999,N_2602,N_4448);
and U6000 (N_6000,N_2976,N_4063);
nor U6001 (N_6001,N_4624,N_3257);
xor U6002 (N_6002,N_2514,N_2585);
nand U6003 (N_6003,N_4672,N_4215);
nor U6004 (N_6004,N_4436,N_4174);
xor U6005 (N_6005,N_4247,N_3863);
xor U6006 (N_6006,N_4125,N_2588);
nor U6007 (N_6007,N_4172,N_3054);
nor U6008 (N_6008,N_3739,N_3236);
and U6009 (N_6009,N_4730,N_3489);
nor U6010 (N_6010,N_4877,N_2908);
and U6011 (N_6011,N_3705,N_2616);
nor U6012 (N_6012,N_4022,N_4322);
nand U6013 (N_6013,N_3086,N_4960);
and U6014 (N_6014,N_3810,N_3202);
and U6015 (N_6015,N_4116,N_3685);
or U6016 (N_6016,N_3443,N_4021);
and U6017 (N_6017,N_2603,N_3026);
nand U6018 (N_6018,N_4832,N_2666);
and U6019 (N_6019,N_3543,N_2560);
nand U6020 (N_6020,N_3974,N_2714);
nand U6021 (N_6021,N_3108,N_4120);
or U6022 (N_6022,N_3668,N_4510);
or U6023 (N_6023,N_3223,N_4421);
or U6024 (N_6024,N_3163,N_4486);
or U6025 (N_6025,N_3273,N_3716);
or U6026 (N_6026,N_2563,N_2791);
nand U6027 (N_6027,N_4361,N_3773);
and U6028 (N_6028,N_3020,N_3375);
nand U6029 (N_6029,N_2967,N_2586);
and U6030 (N_6030,N_3157,N_2839);
and U6031 (N_6031,N_4643,N_4469);
nor U6032 (N_6032,N_4318,N_4411);
nand U6033 (N_6033,N_3786,N_3417);
nor U6034 (N_6034,N_4108,N_3454);
nor U6035 (N_6035,N_4496,N_3499);
nand U6036 (N_6036,N_3788,N_4481);
nor U6037 (N_6037,N_2690,N_4768);
and U6038 (N_6038,N_4060,N_4810);
and U6039 (N_6039,N_3052,N_4732);
nor U6040 (N_6040,N_4616,N_4535);
or U6041 (N_6041,N_3152,N_3084);
nor U6042 (N_6042,N_3103,N_3964);
and U6043 (N_6043,N_4979,N_3859);
nand U6044 (N_6044,N_2502,N_2548);
nand U6045 (N_6045,N_4930,N_2704);
or U6046 (N_6046,N_3602,N_3887);
nand U6047 (N_6047,N_4468,N_4208);
or U6048 (N_6048,N_4037,N_3107);
and U6049 (N_6049,N_4030,N_2847);
or U6050 (N_6050,N_4573,N_4100);
and U6051 (N_6051,N_3770,N_4057);
and U6052 (N_6052,N_3979,N_3051);
and U6053 (N_6053,N_4422,N_4196);
nand U6054 (N_6054,N_4854,N_2668);
or U6055 (N_6055,N_4688,N_3821);
xnor U6056 (N_6056,N_3545,N_2637);
and U6057 (N_6057,N_3516,N_4483);
and U6058 (N_6058,N_4915,N_3109);
and U6059 (N_6059,N_3556,N_2553);
nand U6060 (N_6060,N_2589,N_4876);
nand U6061 (N_6061,N_4343,N_4531);
and U6062 (N_6062,N_4894,N_4899);
or U6063 (N_6063,N_3354,N_4994);
and U6064 (N_6064,N_3738,N_4644);
nand U6065 (N_6065,N_2814,N_3534);
and U6066 (N_6066,N_2677,N_3007);
nand U6067 (N_6067,N_2865,N_3981);
nand U6068 (N_6068,N_4126,N_3936);
xnor U6069 (N_6069,N_4867,N_4061);
nor U6070 (N_6070,N_3189,N_4588);
xnor U6071 (N_6071,N_2877,N_3490);
nand U6072 (N_6072,N_3381,N_4748);
and U6073 (N_6073,N_4168,N_3993);
nor U6074 (N_6074,N_3686,N_4952);
nand U6075 (N_6075,N_4593,N_3502);
nand U6076 (N_6076,N_4667,N_3960);
nand U6077 (N_6077,N_3535,N_4809);
and U6078 (N_6078,N_2641,N_4783);
or U6079 (N_6079,N_4837,N_4995);
and U6080 (N_6080,N_4162,N_4058);
and U6081 (N_6081,N_4471,N_4733);
and U6082 (N_6082,N_3310,N_2506);
nand U6083 (N_6083,N_3140,N_2815);
or U6084 (N_6084,N_4764,N_2724);
or U6085 (N_6085,N_4843,N_3269);
or U6086 (N_6086,N_2787,N_4997);
and U6087 (N_6087,N_2562,N_4929);
nor U6088 (N_6088,N_2520,N_2709);
nor U6089 (N_6089,N_2512,N_3679);
or U6090 (N_6090,N_4506,N_3828);
nor U6091 (N_6091,N_2849,N_3743);
nand U6092 (N_6092,N_4942,N_3737);
or U6093 (N_6093,N_3351,N_4444);
or U6094 (N_6094,N_3655,N_2862);
nand U6095 (N_6095,N_3307,N_4438);
nand U6096 (N_6096,N_4650,N_3145);
and U6097 (N_6097,N_4312,N_4502);
nand U6098 (N_6098,N_3572,N_3763);
and U6099 (N_6099,N_4710,N_4386);
and U6100 (N_6100,N_4095,N_4246);
and U6101 (N_6101,N_4683,N_3253);
and U6102 (N_6102,N_3797,N_4796);
nor U6103 (N_6103,N_2920,N_4757);
nor U6104 (N_6104,N_4111,N_2663);
xnor U6105 (N_6105,N_2966,N_4784);
and U6106 (N_6106,N_4209,N_4332);
nand U6107 (N_6107,N_3298,N_3459);
or U6108 (N_6108,N_3071,N_4609);
nand U6109 (N_6109,N_3733,N_3658);
or U6110 (N_6110,N_2820,N_2741);
and U6111 (N_6111,N_3540,N_2673);
nor U6112 (N_6112,N_2571,N_2670);
nand U6113 (N_6113,N_2937,N_2938);
and U6114 (N_6114,N_2630,N_2559);
and U6115 (N_6115,N_3627,N_4848);
nor U6116 (N_6116,N_2945,N_4389);
and U6117 (N_6117,N_3359,N_3278);
nor U6118 (N_6118,N_3968,N_3334);
or U6119 (N_6119,N_3822,N_4090);
or U6120 (N_6120,N_4734,N_3418);
nor U6121 (N_6121,N_4699,N_4356);
or U6122 (N_6122,N_3312,N_4331);
or U6123 (N_6123,N_2833,N_4182);
and U6124 (N_6124,N_4497,N_3831);
nor U6125 (N_6125,N_2776,N_2866);
nand U6126 (N_6126,N_4190,N_4830);
or U6127 (N_6127,N_3940,N_3085);
and U6128 (N_6128,N_3173,N_2649);
nor U6129 (N_6129,N_2611,N_3373);
and U6130 (N_6130,N_3987,N_2758);
or U6131 (N_6131,N_4512,N_4885);
and U6132 (N_6132,N_4568,N_3992);
or U6133 (N_6133,N_3287,N_3539);
nor U6134 (N_6134,N_4200,N_3732);
nor U6135 (N_6135,N_4016,N_3564);
and U6136 (N_6136,N_4544,N_4661);
nor U6137 (N_6137,N_3468,N_3314);
or U6138 (N_6138,N_3245,N_3082);
nand U6139 (N_6139,N_3266,N_3388);
nor U6140 (N_6140,N_3336,N_2984);
or U6141 (N_6141,N_4164,N_3034);
and U6142 (N_6142,N_2746,N_2986);
and U6143 (N_6143,N_3889,N_2655);
and U6144 (N_6144,N_4645,N_4922);
nand U6145 (N_6145,N_3768,N_2725);
nand U6146 (N_6146,N_3965,N_3194);
nor U6147 (N_6147,N_4159,N_3187);
nor U6148 (N_6148,N_2806,N_4033);
and U6149 (N_6149,N_3466,N_3118);
xnor U6150 (N_6150,N_2547,N_3879);
nor U6151 (N_6151,N_4665,N_3030);
nor U6152 (N_6152,N_3368,N_3156);
nor U6153 (N_6153,N_3072,N_3374);
and U6154 (N_6154,N_4691,N_4487);
or U6155 (N_6155,N_3198,N_2760);
nand U6156 (N_6156,N_4024,N_2697);
nand U6157 (N_6157,N_3970,N_2633);
or U6158 (N_6158,N_3496,N_4641);
nor U6159 (N_6159,N_3950,N_2577);
and U6160 (N_6160,N_4206,N_2890);
and U6161 (N_6161,N_4197,N_4227);
nor U6162 (N_6162,N_4195,N_2774);
and U6163 (N_6163,N_2905,N_3265);
and U6164 (N_6164,N_2716,N_4015);
or U6165 (N_6165,N_4908,N_3326);
nor U6166 (N_6166,N_3019,N_3481);
and U6167 (N_6167,N_4539,N_3110);
nor U6168 (N_6168,N_4587,N_4435);
nand U6169 (N_6169,N_3186,N_2521);
or U6170 (N_6170,N_3205,N_3501);
nor U6171 (N_6171,N_2835,N_3002);
or U6172 (N_6172,N_4335,N_4143);
and U6173 (N_6173,N_4267,N_4005);
and U6174 (N_6174,N_4564,N_4542);
and U6175 (N_6175,N_4052,N_4349);
or U6176 (N_6176,N_3670,N_4244);
and U6177 (N_6177,N_3973,N_4427);
and U6178 (N_6178,N_2948,N_2726);
and U6179 (N_6179,N_3000,N_3671);
or U6180 (N_6180,N_3803,N_3947);
nor U6181 (N_6181,N_4623,N_3233);
nor U6182 (N_6182,N_4804,N_4093);
nor U6183 (N_6183,N_4690,N_4684);
nor U6184 (N_6184,N_4972,N_4529);
nand U6185 (N_6185,N_3832,N_3579);
and U6186 (N_6186,N_3576,N_3710);
and U6187 (N_6187,N_3971,N_3409);
nand U6188 (N_6188,N_3752,N_4646);
or U6189 (N_6189,N_4369,N_4062);
nand U6190 (N_6190,N_3587,N_2584);
nand U6191 (N_6191,N_2845,N_2840);
and U6192 (N_6192,N_4993,N_2878);
nor U6193 (N_6193,N_3224,N_2823);
and U6194 (N_6194,N_3865,N_2848);
nand U6195 (N_6195,N_4475,N_2775);
nand U6196 (N_6196,N_3967,N_2922);
nor U6197 (N_6197,N_4989,N_3337);
nor U6198 (N_6198,N_4948,N_4833);
or U6199 (N_6199,N_3135,N_4949);
or U6200 (N_6200,N_3805,N_4263);
nand U6201 (N_6201,N_3129,N_2748);
nor U6202 (N_6202,N_3446,N_2565);
and U6203 (N_6203,N_3541,N_4943);
nor U6204 (N_6204,N_3081,N_3817);
and U6205 (N_6205,N_3858,N_3021);
nor U6206 (N_6206,N_3360,N_3423);
nor U6207 (N_6207,N_4575,N_4828);
xnor U6208 (N_6208,N_4334,N_3281);
and U6209 (N_6209,N_2642,N_4678);
nand U6210 (N_6210,N_4017,N_4811);
nor U6211 (N_6211,N_4598,N_3507);
nand U6212 (N_6212,N_2684,N_3603);
nor U6213 (N_6213,N_4346,N_3721);
nand U6214 (N_6214,N_4729,N_3473);
or U6215 (N_6215,N_4450,N_2574);
or U6216 (N_6216,N_3073,N_2935);
and U6217 (N_6217,N_3477,N_4418);
nor U6218 (N_6218,N_3645,N_3347);
nand U6219 (N_6219,N_4881,N_4392);
nand U6220 (N_6220,N_4655,N_3647);
or U6221 (N_6221,N_3277,N_3574);
nor U6222 (N_6222,N_3399,N_3814);
nor U6223 (N_6223,N_4393,N_4656);
nor U6224 (N_6224,N_2961,N_2874);
and U6225 (N_6225,N_2568,N_4252);
nand U6226 (N_6226,N_4293,N_3276);
and U6227 (N_6227,N_2764,N_2872);
nor U6228 (N_6228,N_4032,N_3055);
nand U6229 (N_6229,N_3440,N_4423);
or U6230 (N_6230,N_2891,N_3028);
nand U6231 (N_6231,N_4065,N_3250);
nand U6232 (N_6232,N_4150,N_3765);
or U6233 (N_6233,N_3112,N_3150);
nor U6234 (N_6234,N_3561,N_3553);
nand U6235 (N_6235,N_4630,N_3582);
nand U6236 (N_6236,N_3309,N_3917);
or U6237 (N_6237,N_4109,N_4627);
or U6238 (N_6238,N_3955,N_3077);
nor U6239 (N_6239,N_4507,N_3258);
and U6240 (N_6240,N_2721,N_2788);
and U6241 (N_6241,N_3439,N_3441);
nand U6242 (N_6242,N_3830,N_2857);
or U6243 (N_6243,N_2860,N_3978);
nand U6244 (N_6244,N_2798,N_2911);
and U6245 (N_6245,N_2699,N_2816);
nand U6246 (N_6246,N_4451,N_2623);
nor U6247 (N_6247,N_4425,N_3292);
or U6248 (N_6248,N_4431,N_3896);
and U6249 (N_6249,N_2645,N_2631);
nor U6250 (N_6250,N_4733,N_2593);
and U6251 (N_6251,N_2659,N_4349);
nor U6252 (N_6252,N_4690,N_3144);
xnor U6253 (N_6253,N_3990,N_4498);
and U6254 (N_6254,N_4154,N_4862);
nand U6255 (N_6255,N_3462,N_3183);
nand U6256 (N_6256,N_3712,N_4735);
nand U6257 (N_6257,N_4487,N_3952);
and U6258 (N_6258,N_3867,N_3903);
or U6259 (N_6259,N_4458,N_3119);
and U6260 (N_6260,N_3797,N_3035);
or U6261 (N_6261,N_4238,N_2739);
and U6262 (N_6262,N_4238,N_2735);
xor U6263 (N_6263,N_4751,N_2668);
nand U6264 (N_6264,N_4671,N_4964);
nand U6265 (N_6265,N_3269,N_3259);
and U6266 (N_6266,N_4054,N_3758);
nor U6267 (N_6267,N_2760,N_4388);
or U6268 (N_6268,N_4429,N_4525);
and U6269 (N_6269,N_4378,N_4345);
nand U6270 (N_6270,N_4746,N_4533);
or U6271 (N_6271,N_4612,N_4568);
nor U6272 (N_6272,N_3989,N_4521);
nand U6273 (N_6273,N_3911,N_4141);
xnor U6274 (N_6274,N_4493,N_3910);
and U6275 (N_6275,N_4200,N_3039);
nor U6276 (N_6276,N_3570,N_4491);
or U6277 (N_6277,N_3091,N_3903);
and U6278 (N_6278,N_2835,N_2627);
nor U6279 (N_6279,N_4104,N_4072);
nand U6280 (N_6280,N_4404,N_3128);
and U6281 (N_6281,N_3817,N_4599);
nand U6282 (N_6282,N_3986,N_4449);
and U6283 (N_6283,N_3100,N_2880);
nor U6284 (N_6284,N_4184,N_3242);
xor U6285 (N_6285,N_3836,N_3788);
nor U6286 (N_6286,N_4685,N_4219);
and U6287 (N_6287,N_4577,N_3998);
and U6288 (N_6288,N_2610,N_3697);
nand U6289 (N_6289,N_3927,N_2916);
or U6290 (N_6290,N_4110,N_4675);
and U6291 (N_6291,N_4323,N_3704);
or U6292 (N_6292,N_4888,N_4847);
nand U6293 (N_6293,N_2977,N_4392);
or U6294 (N_6294,N_3716,N_3252);
or U6295 (N_6295,N_3386,N_3199);
or U6296 (N_6296,N_4660,N_4676);
nand U6297 (N_6297,N_4556,N_2920);
and U6298 (N_6298,N_4120,N_3304);
nand U6299 (N_6299,N_3612,N_4393);
and U6300 (N_6300,N_4154,N_4630);
nand U6301 (N_6301,N_4182,N_4105);
nand U6302 (N_6302,N_2724,N_4433);
and U6303 (N_6303,N_3974,N_3223);
nor U6304 (N_6304,N_4663,N_3616);
or U6305 (N_6305,N_4039,N_3303);
and U6306 (N_6306,N_2770,N_3559);
nand U6307 (N_6307,N_3120,N_4438);
nor U6308 (N_6308,N_4206,N_4179);
nor U6309 (N_6309,N_2629,N_4680);
nand U6310 (N_6310,N_4021,N_3863);
and U6311 (N_6311,N_3508,N_3563);
and U6312 (N_6312,N_3520,N_4039);
or U6313 (N_6313,N_3201,N_4070);
nor U6314 (N_6314,N_2764,N_4026);
nor U6315 (N_6315,N_2663,N_4323);
or U6316 (N_6316,N_4107,N_4372);
or U6317 (N_6317,N_4140,N_3941);
or U6318 (N_6318,N_3263,N_4979);
xnor U6319 (N_6319,N_4525,N_4522);
nand U6320 (N_6320,N_2550,N_4881);
xor U6321 (N_6321,N_2850,N_3361);
or U6322 (N_6322,N_2609,N_3102);
and U6323 (N_6323,N_3337,N_2898);
and U6324 (N_6324,N_3637,N_3734);
or U6325 (N_6325,N_3572,N_3028);
or U6326 (N_6326,N_3275,N_2905);
or U6327 (N_6327,N_3153,N_3634);
and U6328 (N_6328,N_4798,N_4677);
nor U6329 (N_6329,N_2600,N_2559);
or U6330 (N_6330,N_4094,N_4321);
nand U6331 (N_6331,N_2792,N_3262);
or U6332 (N_6332,N_2921,N_3416);
or U6333 (N_6333,N_2716,N_4795);
or U6334 (N_6334,N_4441,N_4803);
and U6335 (N_6335,N_3938,N_3361);
nor U6336 (N_6336,N_4974,N_2982);
nor U6337 (N_6337,N_4558,N_2598);
and U6338 (N_6338,N_4869,N_4245);
nand U6339 (N_6339,N_4032,N_3538);
and U6340 (N_6340,N_2903,N_2707);
nand U6341 (N_6341,N_3842,N_3263);
nand U6342 (N_6342,N_2687,N_4360);
nand U6343 (N_6343,N_4463,N_3234);
and U6344 (N_6344,N_3064,N_3326);
or U6345 (N_6345,N_3803,N_4609);
and U6346 (N_6346,N_3464,N_4597);
nor U6347 (N_6347,N_3523,N_4935);
nor U6348 (N_6348,N_4291,N_2612);
nand U6349 (N_6349,N_4307,N_4211);
and U6350 (N_6350,N_3303,N_3811);
nand U6351 (N_6351,N_4222,N_4391);
nand U6352 (N_6352,N_3735,N_4005);
or U6353 (N_6353,N_2536,N_4204);
or U6354 (N_6354,N_4628,N_3033);
or U6355 (N_6355,N_4172,N_2952);
or U6356 (N_6356,N_4816,N_4647);
nand U6357 (N_6357,N_3541,N_3731);
nand U6358 (N_6358,N_4244,N_2570);
nand U6359 (N_6359,N_3511,N_2882);
or U6360 (N_6360,N_3495,N_4796);
nor U6361 (N_6361,N_4092,N_4618);
nor U6362 (N_6362,N_3573,N_4538);
nand U6363 (N_6363,N_4078,N_3445);
and U6364 (N_6364,N_3007,N_2928);
nor U6365 (N_6365,N_3495,N_3604);
or U6366 (N_6366,N_3555,N_2614);
nand U6367 (N_6367,N_2707,N_4648);
nor U6368 (N_6368,N_4170,N_4505);
nor U6369 (N_6369,N_3954,N_4481);
xnor U6370 (N_6370,N_2645,N_4674);
or U6371 (N_6371,N_2972,N_4036);
or U6372 (N_6372,N_3736,N_2701);
nor U6373 (N_6373,N_3904,N_2740);
or U6374 (N_6374,N_3904,N_3026);
or U6375 (N_6375,N_3553,N_4642);
or U6376 (N_6376,N_4430,N_3490);
nand U6377 (N_6377,N_4709,N_4799);
and U6378 (N_6378,N_3527,N_3886);
or U6379 (N_6379,N_4868,N_3126);
nand U6380 (N_6380,N_3986,N_3910);
nor U6381 (N_6381,N_3567,N_3773);
nand U6382 (N_6382,N_2930,N_4615);
nand U6383 (N_6383,N_4030,N_4523);
nand U6384 (N_6384,N_2971,N_4112);
nand U6385 (N_6385,N_4115,N_4331);
or U6386 (N_6386,N_4286,N_4910);
nor U6387 (N_6387,N_3849,N_2801);
or U6388 (N_6388,N_3989,N_3012);
and U6389 (N_6389,N_4397,N_4008);
or U6390 (N_6390,N_4015,N_3155);
nand U6391 (N_6391,N_3445,N_4182);
nor U6392 (N_6392,N_3338,N_4261);
or U6393 (N_6393,N_3498,N_3575);
nor U6394 (N_6394,N_3874,N_3122);
xor U6395 (N_6395,N_2575,N_3198);
nand U6396 (N_6396,N_2892,N_3691);
nand U6397 (N_6397,N_2629,N_3674);
and U6398 (N_6398,N_3237,N_3359);
or U6399 (N_6399,N_3138,N_4309);
or U6400 (N_6400,N_3935,N_3644);
nor U6401 (N_6401,N_2616,N_4943);
or U6402 (N_6402,N_4751,N_2998);
nand U6403 (N_6403,N_4294,N_4662);
nand U6404 (N_6404,N_3805,N_4664);
or U6405 (N_6405,N_4222,N_2732);
nand U6406 (N_6406,N_2886,N_4399);
and U6407 (N_6407,N_2757,N_3095);
nand U6408 (N_6408,N_4874,N_4386);
nor U6409 (N_6409,N_4734,N_3185);
or U6410 (N_6410,N_2800,N_4972);
or U6411 (N_6411,N_3427,N_3036);
or U6412 (N_6412,N_2994,N_2582);
nand U6413 (N_6413,N_4583,N_2947);
xnor U6414 (N_6414,N_4708,N_3535);
nand U6415 (N_6415,N_4692,N_3175);
or U6416 (N_6416,N_4265,N_4537);
or U6417 (N_6417,N_3808,N_4556);
or U6418 (N_6418,N_2919,N_4259);
nor U6419 (N_6419,N_4283,N_4541);
nor U6420 (N_6420,N_3316,N_2925);
nor U6421 (N_6421,N_4828,N_4467);
and U6422 (N_6422,N_3782,N_4158);
nor U6423 (N_6423,N_3218,N_4432);
or U6424 (N_6424,N_3772,N_3474);
nor U6425 (N_6425,N_3604,N_2831);
nand U6426 (N_6426,N_4183,N_3051);
or U6427 (N_6427,N_2679,N_4273);
or U6428 (N_6428,N_4501,N_3511);
nand U6429 (N_6429,N_3511,N_2943);
or U6430 (N_6430,N_4720,N_2995);
and U6431 (N_6431,N_4073,N_4205);
or U6432 (N_6432,N_4730,N_2684);
nand U6433 (N_6433,N_4423,N_4891);
xnor U6434 (N_6434,N_3997,N_3168);
or U6435 (N_6435,N_2576,N_3780);
and U6436 (N_6436,N_4291,N_2735);
or U6437 (N_6437,N_2884,N_4618);
nor U6438 (N_6438,N_3386,N_3914);
nand U6439 (N_6439,N_4219,N_4591);
and U6440 (N_6440,N_3368,N_3483);
and U6441 (N_6441,N_2546,N_3897);
or U6442 (N_6442,N_4560,N_2949);
and U6443 (N_6443,N_4143,N_3953);
or U6444 (N_6444,N_2926,N_3185);
and U6445 (N_6445,N_4350,N_4255);
nor U6446 (N_6446,N_3036,N_3745);
nor U6447 (N_6447,N_3288,N_3914);
or U6448 (N_6448,N_4459,N_3304);
and U6449 (N_6449,N_3423,N_3126);
and U6450 (N_6450,N_2573,N_4990);
xnor U6451 (N_6451,N_4751,N_3297);
or U6452 (N_6452,N_4059,N_3393);
and U6453 (N_6453,N_3415,N_3368);
or U6454 (N_6454,N_3617,N_3901);
nor U6455 (N_6455,N_3162,N_4098);
nand U6456 (N_6456,N_4901,N_2980);
and U6457 (N_6457,N_3086,N_2925);
nand U6458 (N_6458,N_2829,N_4195);
and U6459 (N_6459,N_4612,N_4065);
nand U6460 (N_6460,N_3003,N_3095);
nor U6461 (N_6461,N_2882,N_4697);
and U6462 (N_6462,N_2808,N_3639);
nand U6463 (N_6463,N_3853,N_4787);
and U6464 (N_6464,N_2618,N_2535);
nand U6465 (N_6465,N_4429,N_2810);
nor U6466 (N_6466,N_4803,N_4329);
xor U6467 (N_6467,N_3760,N_2803);
nor U6468 (N_6468,N_4946,N_3548);
or U6469 (N_6469,N_2840,N_3105);
and U6470 (N_6470,N_3853,N_3332);
and U6471 (N_6471,N_4376,N_3927);
and U6472 (N_6472,N_4893,N_4037);
nor U6473 (N_6473,N_2638,N_4352);
nand U6474 (N_6474,N_4108,N_4245);
nand U6475 (N_6475,N_4549,N_3050);
nand U6476 (N_6476,N_3175,N_2562);
or U6477 (N_6477,N_3016,N_2597);
or U6478 (N_6478,N_4069,N_3377);
nand U6479 (N_6479,N_3340,N_3553);
nor U6480 (N_6480,N_4430,N_3180);
xor U6481 (N_6481,N_4124,N_3877);
or U6482 (N_6482,N_4108,N_4201);
nand U6483 (N_6483,N_2898,N_3653);
nor U6484 (N_6484,N_4286,N_4654);
nor U6485 (N_6485,N_2935,N_4033);
or U6486 (N_6486,N_3992,N_4874);
nand U6487 (N_6487,N_2921,N_2607);
nor U6488 (N_6488,N_3365,N_4504);
or U6489 (N_6489,N_3362,N_4912);
nor U6490 (N_6490,N_3290,N_2707);
nor U6491 (N_6491,N_2992,N_3393);
or U6492 (N_6492,N_4703,N_2544);
nand U6493 (N_6493,N_3594,N_4264);
nand U6494 (N_6494,N_3032,N_4110);
nand U6495 (N_6495,N_4916,N_2636);
and U6496 (N_6496,N_4333,N_3308);
nand U6497 (N_6497,N_3194,N_4430);
nand U6498 (N_6498,N_3877,N_4423);
nand U6499 (N_6499,N_4427,N_3286);
and U6500 (N_6500,N_3869,N_4174);
and U6501 (N_6501,N_2770,N_4675);
or U6502 (N_6502,N_4599,N_4576);
nand U6503 (N_6503,N_4774,N_3612);
nor U6504 (N_6504,N_2752,N_2950);
nor U6505 (N_6505,N_3317,N_3819);
or U6506 (N_6506,N_4539,N_4648);
nor U6507 (N_6507,N_4965,N_4325);
or U6508 (N_6508,N_3260,N_4061);
nand U6509 (N_6509,N_4228,N_4190);
or U6510 (N_6510,N_4934,N_3017);
or U6511 (N_6511,N_3093,N_4310);
nor U6512 (N_6512,N_3009,N_4675);
or U6513 (N_6513,N_3457,N_3875);
nor U6514 (N_6514,N_3899,N_2599);
nand U6515 (N_6515,N_2533,N_4287);
nor U6516 (N_6516,N_4351,N_4985);
nand U6517 (N_6517,N_3815,N_4856);
nor U6518 (N_6518,N_3427,N_4575);
or U6519 (N_6519,N_3418,N_3350);
or U6520 (N_6520,N_3055,N_2732);
nand U6521 (N_6521,N_4174,N_3850);
nand U6522 (N_6522,N_3714,N_2571);
xnor U6523 (N_6523,N_2525,N_2777);
and U6524 (N_6524,N_2848,N_4140);
nand U6525 (N_6525,N_3632,N_4320);
or U6526 (N_6526,N_2821,N_2599);
nor U6527 (N_6527,N_2568,N_4723);
and U6528 (N_6528,N_2749,N_2568);
nand U6529 (N_6529,N_3888,N_2860);
and U6530 (N_6530,N_4720,N_4264);
nand U6531 (N_6531,N_3753,N_4929);
and U6532 (N_6532,N_3050,N_4629);
or U6533 (N_6533,N_3772,N_3451);
nor U6534 (N_6534,N_3234,N_2674);
and U6535 (N_6535,N_2883,N_3555);
or U6536 (N_6536,N_2748,N_3653);
nand U6537 (N_6537,N_4298,N_3373);
nand U6538 (N_6538,N_2948,N_3292);
nor U6539 (N_6539,N_3717,N_3318);
or U6540 (N_6540,N_3726,N_3017);
nor U6541 (N_6541,N_4099,N_2901);
or U6542 (N_6542,N_4722,N_3122);
and U6543 (N_6543,N_3217,N_3706);
nor U6544 (N_6544,N_3614,N_3547);
nor U6545 (N_6545,N_3207,N_3833);
or U6546 (N_6546,N_4071,N_2704);
nor U6547 (N_6547,N_3511,N_3481);
nor U6548 (N_6548,N_4033,N_3606);
or U6549 (N_6549,N_4545,N_2690);
nor U6550 (N_6550,N_4713,N_3424);
or U6551 (N_6551,N_4028,N_3482);
nand U6552 (N_6552,N_4557,N_4425);
nand U6553 (N_6553,N_3520,N_3199);
or U6554 (N_6554,N_3952,N_2975);
nor U6555 (N_6555,N_2907,N_4534);
or U6556 (N_6556,N_4690,N_4361);
nand U6557 (N_6557,N_3994,N_4232);
and U6558 (N_6558,N_4054,N_2813);
nand U6559 (N_6559,N_2564,N_3848);
xnor U6560 (N_6560,N_3702,N_4559);
and U6561 (N_6561,N_3171,N_3060);
nand U6562 (N_6562,N_3286,N_4719);
nor U6563 (N_6563,N_4244,N_2703);
nor U6564 (N_6564,N_4839,N_4101);
nand U6565 (N_6565,N_4189,N_4913);
or U6566 (N_6566,N_2604,N_4326);
nor U6567 (N_6567,N_4325,N_4566);
or U6568 (N_6568,N_4205,N_4804);
and U6569 (N_6569,N_2647,N_3378);
xnor U6570 (N_6570,N_3284,N_2735);
or U6571 (N_6571,N_3898,N_2694);
or U6572 (N_6572,N_3417,N_3331);
and U6573 (N_6573,N_3778,N_2581);
or U6574 (N_6574,N_2961,N_2843);
or U6575 (N_6575,N_3015,N_4916);
or U6576 (N_6576,N_4835,N_2742);
and U6577 (N_6577,N_3182,N_4793);
nand U6578 (N_6578,N_2674,N_4053);
nand U6579 (N_6579,N_4603,N_4360);
or U6580 (N_6580,N_3726,N_3070);
nand U6581 (N_6581,N_2934,N_3640);
nand U6582 (N_6582,N_4450,N_4031);
and U6583 (N_6583,N_2708,N_4904);
nor U6584 (N_6584,N_3662,N_3136);
nand U6585 (N_6585,N_4516,N_4566);
nor U6586 (N_6586,N_2574,N_4430);
nor U6587 (N_6587,N_3364,N_3518);
nand U6588 (N_6588,N_4495,N_3293);
nor U6589 (N_6589,N_4270,N_4746);
nor U6590 (N_6590,N_2920,N_2583);
and U6591 (N_6591,N_4442,N_2672);
and U6592 (N_6592,N_4617,N_4057);
or U6593 (N_6593,N_4550,N_3740);
or U6594 (N_6594,N_2912,N_3389);
nor U6595 (N_6595,N_3151,N_3101);
or U6596 (N_6596,N_3418,N_2709);
and U6597 (N_6597,N_4695,N_3800);
and U6598 (N_6598,N_3321,N_4577);
xor U6599 (N_6599,N_4240,N_4156);
nor U6600 (N_6600,N_2793,N_3079);
nand U6601 (N_6601,N_2994,N_3192);
nor U6602 (N_6602,N_3977,N_4205);
nor U6603 (N_6603,N_4523,N_4202);
nor U6604 (N_6604,N_2568,N_4266);
nand U6605 (N_6605,N_4967,N_3858);
or U6606 (N_6606,N_2683,N_4010);
nand U6607 (N_6607,N_3096,N_4754);
and U6608 (N_6608,N_3210,N_3156);
or U6609 (N_6609,N_4434,N_3069);
and U6610 (N_6610,N_4818,N_3059);
and U6611 (N_6611,N_2782,N_4721);
nor U6612 (N_6612,N_4130,N_4136);
or U6613 (N_6613,N_2640,N_3119);
nor U6614 (N_6614,N_2885,N_3785);
xnor U6615 (N_6615,N_4465,N_3531);
nand U6616 (N_6616,N_3423,N_4391);
nand U6617 (N_6617,N_2562,N_4138);
or U6618 (N_6618,N_3661,N_3318);
and U6619 (N_6619,N_4112,N_3332);
and U6620 (N_6620,N_3766,N_4193);
and U6621 (N_6621,N_2519,N_3770);
and U6622 (N_6622,N_3878,N_3710);
or U6623 (N_6623,N_2996,N_4943);
nor U6624 (N_6624,N_4284,N_3423);
nand U6625 (N_6625,N_3110,N_2517);
or U6626 (N_6626,N_4624,N_4636);
or U6627 (N_6627,N_3018,N_3789);
or U6628 (N_6628,N_3044,N_3225);
nand U6629 (N_6629,N_3686,N_2717);
or U6630 (N_6630,N_2684,N_4837);
or U6631 (N_6631,N_3535,N_4544);
nor U6632 (N_6632,N_4415,N_3315);
and U6633 (N_6633,N_4441,N_4320);
nand U6634 (N_6634,N_2710,N_4945);
or U6635 (N_6635,N_3076,N_2785);
nor U6636 (N_6636,N_2574,N_2782);
or U6637 (N_6637,N_3514,N_4806);
and U6638 (N_6638,N_3314,N_4388);
nor U6639 (N_6639,N_4987,N_4245);
and U6640 (N_6640,N_3423,N_3745);
nor U6641 (N_6641,N_2843,N_3641);
nand U6642 (N_6642,N_3669,N_4593);
or U6643 (N_6643,N_2807,N_4392);
or U6644 (N_6644,N_4147,N_3048);
and U6645 (N_6645,N_4445,N_4168);
and U6646 (N_6646,N_4849,N_4932);
nand U6647 (N_6647,N_4959,N_3133);
or U6648 (N_6648,N_4783,N_3085);
and U6649 (N_6649,N_3167,N_3663);
or U6650 (N_6650,N_2671,N_4662);
xnor U6651 (N_6651,N_3175,N_4488);
nor U6652 (N_6652,N_2813,N_4148);
or U6653 (N_6653,N_2808,N_3192);
or U6654 (N_6654,N_3682,N_4853);
and U6655 (N_6655,N_3476,N_4097);
nand U6656 (N_6656,N_3624,N_3687);
nor U6657 (N_6657,N_4415,N_3911);
nor U6658 (N_6658,N_4397,N_4514);
or U6659 (N_6659,N_2978,N_2704);
nor U6660 (N_6660,N_3241,N_4709);
nor U6661 (N_6661,N_4213,N_2962);
and U6662 (N_6662,N_4251,N_4814);
nor U6663 (N_6663,N_2659,N_3979);
and U6664 (N_6664,N_3102,N_4660);
or U6665 (N_6665,N_3698,N_2955);
and U6666 (N_6666,N_2809,N_4359);
and U6667 (N_6667,N_3285,N_4743);
and U6668 (N_6668,N_4895,N_4502);
or U6669 (N_6669,N_2725,N_2810);
nand U6670 (N_6670,N_4604,N_2657);
and U6671 (N_6671,N_2691,N_4740);
or U6672 (N_6672,N_3978,N_4645);
and U6673 (N_6673,N_4430,N_3188);
or U6674 (N_6674,N_2592,N_3793);
nand U6675 (N_6675,N_4844,N_3837);
or U6676 (N_6676,N_3340,N_4126);
and U6677 (N_6677,N_4278,N_2746);
nand U6678 (N_6678,N_3573,N_3699);
or U6679 (N_6679,N_4872,N_4428);
or U6680 (N_6680,N_2654,N_4468);
or U6681 (N_6681,N_2605,N_3670);
nand U6682 (N_6682,N_4523,N_3512);
nand U6683 (N_6683,N_4566,N_2725);
nor U6684 (N_6684,N_4407,N_2589);
or U6685 (N_6685,N_2910,N_3734);
xor U6686 (N_6686,N_4471,N_2910);
nor U6687 (N_6687,N_3213,N_4897);
and U6688 (N_6688,N_3770,N_3098);
nor U6689 (N_6689,N_3099,N_4906);
nor U6690 (N_6690,N_3148,N_3249);
nor U6691 (N_6691,N_2810,N_2684);
or U6692 (N_6692,N_3745,N_4084);
xor U6693 (N_6693,N_3464,N_3514);
nand U6694 (N_6694,N_3532,N_3649);
xor U6695 (N_6695,N_3436,N_2862);
or U6696 (N_6696,N_3648,N_2945);
and U6697 (N_6697,N_2790,N_4431);
or U6698 (N_6698,N_2509,N_3684);
nand U6699 (N_6699,N_4330,N_4547);
nor U6700 (N_6700,N_4048,N_4317);
nor U6701 (N_6701,N_4950,N_3169);
or U6702 (N_6702,N_3124,N_3103);
xor U6703 (N_6703,N_4748,N_4602);
nor U6704 (N_6704,N_4936,N_3075);
or U6705 (N_6705,N_2657,N_2677);
nand U6706 (N_6706,N_2639,N_3996);
or U6707 (N_6707,N_3214,N_2556);
and U6708 (N_6708,N_2876,N_4348);
nor U6709 (N_6709,N_4607,N_3136);
or U6710 (N_6710,N_3538,N_4847);
or U6711 (N_6711,N_3767,N_2598);
nand U6712 (N_6712,N_4160,N_3004);
nand U6713 (N_6713,N_4439,N_2872);
or U6714 (N_6714,N_2630,N_3769);
nand U6715 (N_6715,N_2873,N_3569);
and U6716 (N_6716,N_2552,N_4634);
nor U6717 (N_6717,N_4055,N_3417);
nor U6718 (N_6718,N_2672,N_2710);
nor U6719 (N_6719,N_4586,N_4053);
nor U6720 (N_6720,N_4556,N_3108);
nor U6721 (N_6721,N_3299,N_3963);
or U6722 (N_6722,N_4408,N_4935);
nor U6723 (N_6723,N_2881,N_3164);
or U6724 (N_6724,N_2682,N_4819);
nand U6725 (N_6725,N_4967,N_4624);
and U6726 (N_6726,N_2865,N_2509);
or U6727 (N_6727,N_4765,N_4607);
nand U6728 (N_6728,N_3840,N_2967);
nor U6729 (N_6729,N_3045,N_4568);
or U6730 (N_6730,N_3735,N_3388);
and U6731 (N_6731,N_3362,N_2835);
and U6732 (N_6732,N_3356,N_4899);
nor U6733 (N_6733,N_3488,N_3156);
nor U6734 (N_6734,N_3458,N_3442);
nor U6735 (N_6735,N_4294,N_2911);
and U6736 (N_6736,N_2994,N_3471);
nor U6737 (N_6737,N_3949,N_3320);
nand U6738 (N_6738,N_4932,N_4540);
and U6739 (N_6739,N_3303,N_4377);
and U6740 (N_6740,N_4967,N_2738);
nand U6741 (N_6741,N_3011,N_3038);
xor U6742 (N_6742,N_2653,N_3773);
nand U6743 (N_6743,N_2859,N_3131);
and U6744 (N_6744,N_4068,N_4436);
or U6745 (N_6745,N_4010,N_4167);
nor U6746 (N_6746,N_3432,N_4966);
nand U6747 (N_6747,N_4597,N_3508);
nand U6748 (N_6748,N_4359,N_4927);
or U6749 (N_6749,N_2869,N_4679);
and U6750 (N_6750,N_3157,N_3631);
nor U6751 (N_6751,N_3229,N_4879);
nor U6752 (N_6752,N_4248,N_2988);
nand U6753 (N_6753,N_3661,N_3907);
nand U6754 (N_6754,N_2667,N_2622);
and U6755 (N_6755,N_3157,N_4037);
nor U6756 (N_6756,N_3953,N_2831);
nor U6757 (N_6757,N_3521,N_4410);
and U6758 (N_6758,N_4919,N_3108);
nor U6759 (N_6759,N_2851,N_4217);
nor U6760 (N_6760,N_3473,N_4403);
nand U6761 (N_6761,N_2778,N_3577);
or U6762 (N_6762,N_4770,N_3066);
or U6763 (N_6763,N_4789,N_3695);
nor U6764 (N_6764,N_4163,N_4566);
nand U6765 (N_6765,N_3419,N_4445);
and U6766 (N_6766,N_4906,N_2527);
nor U6767 (N_6767,N_3491,N_4509);
nand U6768 (N_6768,N_3602,N_4704);
or U6769 (N_6769,N_4633,N_4062);
nand U6770 (N_6770,N_3773,N_3996);
nor U6771 (N_6771,N_3085,N_3575);
and U6772 (N_6772,N_3367,N_3669);
nand U6773 (N_6773,N_3414,N_4807);
or U6774 (N_6774,N_3557,N_3293);
nor U6775 (N_6775,N_3606,N_2508);
nor U6776 (N_6776,N_4066,N_4080);
nand U6777 (N_6777,N_4570,N_4322);
or U6778 (N_6778,N_4404,N_2640);
nand U6779 (N_6779,N_3278,N_4619);
nor U6780 (N_6780,N_3631,N_4546);
nor U6781 (N_6781,N_3733,N_3695);
or U6782 (N_6782,N_4154,N_3479);
and U6783 (N_6783,N_4741,N_2542);
and U6784 (N_6784,N_4680,N_4051);
and U6785 (N_6785,N_2654,N_2694);
or U6786 (N_6786,N_2966,N_4199);
nand U6787 (N_6787,N_4121,N_4512);
or U6788 (N_6788,N_3704,N_4855);
and U6789 (N_6789,N_4046,N_3987);
or U6790 (N_6790,N_4598,N_4869);
and U6791 (N_6791,N_3132,N_3962);
xnor U6792 (N_6792,N_3555,N_4233);
nand U6793 (N_6793,N_4683,N_4021);
nor U6794 (N_6794,N_3293,N_2590);
or U6795 (N_6795,N_3551,N_3654);
nor U6796 (N_6796,N_3050,N_2635);
or U6797 (N_6797,N_4839,N_4853);
nand U6798 (N_6798,N_2602,N_3342);
or U6799 (N_6799,N_3440,N_4054);
or U6800 (N_6800,N_3311,N_4088);
and U6801 (N_6801,N_4972,N_4574);
nand U6802 (N_6802,N_4518,N_3712);
or U6803 (N_6803,N_3827,N_4053);
nand U6804 (N_6804,N_3447,N_3561);
nor U6805 (N_6805,N_3766,N_4665);
nor U6806 (N_6806,N_3426,N_4434);
and U6807 (N_6807,N_4184,N_4000);
nor U6808 (N_6808,N_3415,N_3487);
and U6809 (N_6809,N_3017,N_3997);
or U6810 (N_6810,N_3405,N_3512);
or U6811 (N_6811,N_4873,N_2783);
or U6812 (N_6812,N_4296,N_4628);
nor U6813 (N_6813,N_4946,N_3638);
or U6814 (N_6814,N_3673,N_3289);
and U6815 (N_6815,N_4186,N_3532);
and U6816 (N_6816,N_4209,N_3668);
and U6817 (N_6817,N_2642,N_4650);
or U6818 (N_6818,N_3408,N_2962);
nor U6819 (N_6819,N_4669,N_4943);
or U6820 (N_6820,N_4178,N_3550);
nor U6821 (N_6821,N_4509,N_4261);
or U6822 (N_6822,N_3295,N_4733);
nor U6823 (N_6823,N_3222,N_4994);
or U6824 (N_6824,N_3346,N_3909);
nor U6825 (N_6825,N_4354,N_4946);
and U6826 (N_6826,N_2657,N_2830);
nor U6827 (N_6827,N_3229,N_4164);
nand U6828 (N_6828,N_4746,N_4555);
nor U6829 (N_6829,N_3697,N_3255);
or U6830 (N_6830,N_2704,N_3109);
nor U6831 (N_6831,N_3434,N_2536);
or U6832 (N_6832,N_4197,N_3951);
nand U6833 (N_6833,N_4381,N_2881);
and U6834 (N_6834,N_3249,N_4768);
nand U6835 (N_6835,N_2801,N_4199);
nor U6836 (N_6836,N_2553,N_4644);
or U6837 (N_6837,N_4688,N_4896);
xor U6838 (N_6838,N_2770,N_4736);
nand U6839 (N_6839,N_4936,N_4354);
and U6840 (N_6840,N_4030,N_4941);
and U6841 (N_6841,N_2831,N_2932);
and U6842 (N_6842,N_4361,N_2732);
nor U6843 (N_6843,N_3272,N_2966);
and U6844 (N_6844,N_4787,N_4473);
nand U6845 (N_6845,N_4012,N_3230);
nor U6846 (N_6846,N_3131,N_4947);
nand U6847 (N_6847,N_4628,N_2657);
nand U6848 (N_6848,N_3231,N_4564);
and U6849 (N_6849,N_3929,N_2837);
nand U6850 (N_6850,N_4348,N_4068);
or U6851 (N_6851,N_3748,N_3349);
or U6852 (N_6852,N_4761,N_3375);
nor U6853 (N_6853,N_4307,N_4584);
or U6854 (N_6854,N_4444,N_2576);
or U6855 (N_6855,N_3909,N_4842);
or U6856 (N_6856,N_4949,N_3187);
and U6857 (N_6857,N_3234,N_2634);
nor U6858 (N_6858,N_4772,N_2946);
and U6859 (N_6859,N_3551,N_4703);
xnor U6860 (N_6860,N_4536,N_3365);
nor U6861 (N_6861,N_3026,N_2847);
and U6862 (N_6862,N_2875,N_3902);
nor U6863 (N_6863,N_3834,N_3002);
or U6864 (N_6864,N_4860,N_4569);
nand U6865 (N_6865,N_4465,N_4025);
and U6866 (N_6866,N_3930,N_4477);
nand U6867 (N_6867,N_2950,N_3799);
nor U6868 (N_6868,N_2663,N_4514);
nor U6869 (N_6869,N_4898,N_2624);
and U6870 (N_6870,N_3070,N_3405);
or U6871 (N_6871,N_4203,N_3341);
or U6872 (N_6872,N_4825,N_3621);
nor U6873 (N_6873,N_4286,N_4249);
nor U6874 (N_6874,N_3965,N_2523);
and U6875 (N_6875,N_3455,N_4807);
nand U6876 (N_6876,N_4292,N_3074);
or U6877 (N_6877,N_2656,N_3495);
nor U6878 (N_6878,N_4091,N_4440);
nor U6879 (N_6879,N_2654,N_3667);
nand U6880 (N_6880,N_4316,N_4996);
nor U6881 (N_6881,N_4836,N_4233);
or U6882 (N_6882,N_4267,N_3066);
and U6883 (N_6883,N_4837,N_2705);
or U6884 (N_6884,N_4648,N_3630);
nand U6885 (N_6885,N_4975,N_4836);
xor U6886 (N_6886,N_3083,N_4214);
and U6887 (N_6887,N_3512,N_3751);
nor U6888 (N_6888,N_3320,N_4877);
and U6889 (N_6889,N_2602,N_4151);
and U6890 (N_6890,N_4724,N_4106);
nand U6891 (N_6891,N_2891,N_4167);
or U6892 (N_6892,N_3990,N_2546);
or U6893 (N_6893,N_4219,N_3872);
or U6894 (N_6894,N_3566,N_3883);
nor U6895 (N_6895,N_2851,N_4559);
and U6896 (N_6896,N_3923,N_3594);
nand U6897 (N_6897,N_3739,N_4545);
and U6898 (N_6898,N_2915,N_3986);
nand U6899 (N_6899,N_2575,N_4700);
or U6900 (N_6900,N_3412,N_3313);
nor U6901 (N_6901,N_3213,N_3861);
nor U6902 (N_6902,N_2954,N_2561);
nor U6903 (N_6903,N_3454,N_2962);
and U6904 (N_6904,N_3266,N_3605);
or U6905 (N_6905,N_3121,N_4589);
nor U6906 (N_6906,N_2824,N_4129);
or U6907 (N_6907,N_3013,N_4426);
nand U6908 (N_6908,N_2688,N_4294);
and U6909 (N_6909,N_4727,N_4910);
or U6910 (N_6910,N_4371,N_3041);
nand U6911 (N_6911,N_4911,N_4714);
and U6912 (N_6912,N_4763,N_2940);
nor U6913 (N_6913,N_2738,N_2900);
nor U6914 (N_6914,N_2663,N_4896);
or U6915 (N_6915,N_3412,N_4245);
and U6916 (N_6916,N_4585,N_3275);
or U6917 (N_6917,N_3822,N_4805);
nand U6918 (N_6918,N_3273,N_4867);
and U6919 (N_6919,N_4344,N_3678);
nor U6920 (N_6920,N_4946,N_4809);
and U6921 (N_6921,N_3290,N_3523);
or U6922 (N_6922,N_2644,N_2725);
nor U6923 (N_6923,N_4554,N_3451);
and U6924 (N_6924,N_2874,N_4821);
nand U6925 (N_6925,N_4583,N_2578);
and U6926 (N_6926,N_2560,N_4816);
nand U6927 (N_6927,N_4198,N_4024);
nand U6928 (N_6928,N_4469,N_3082);
or U6929 (N_6929,N_3510,N_3764);
nor U6930 (N_6930,N_2791,N_4247);
nand U6931 (N_6931,N_3500,N_4984);
xnor U6932 (N_6932,N_3854,N_2846);
nand U6933 (N_6933,N_2879,N_3997);
xnor U6934 (N_6934,N_3414,N_4484);
nand U6935 (N_6935,N_4465,N_4434);
and U6936 (N_6936,N_2503,N_3940);
nor U6937 (N_6937,N_3576,N_3588);
or U6938 (N_6938,N_3214,N_4753);
nand U6939 (N_6939,N_3779,N_3260);
nor U6940 (N_6940,N_3093,N_3386);
nand U6941 (N_6941,N_3352,N_3870);
nand U6942 (N_6942,N_3970,N_3710);
or U6943 (N_6943,N_3997,N_4838);
xor U6944 (N_6944,N_3858,N_2650);
and U6945 (N_6945,N_2997,N_3316);
or U6946 (N_6946,N_4662,N_2537);
or U6947 (N_6947,N_4648,N_4756);
nand U6948 (N_6948,N_3610,N_4580);
nor U6949 (N_6949,N_3700,N_4837);
or U6950 (N_6950,N_3404,N_3201);
nand U6951 (N_6951,N_4097,N_4948);
nor U6952 (N_6952,N_3964,N_3374);
or U6953 (N_6953,N_2845,N_4133);
nor U6954 (N_6954,N_4185,N_3029);
nor U6955 (N_6955,N_2617,N_2904);
nor U6956 (N_6956,N_4826,N_3574);
or U6957 (N_6957,N_3682,N_3967);
or U6958 (N_6958,N_3373,N_3147);
nand U6959 (N_6959,N_4386,N_4699);
and U6960 (N_6960,N_3674,N_4104);
or U6961 (N_6961,N_4937,N_2806);
or U6962 (N_6962,N_2560,N_3919);
nand U6963 (N_6963,N_3222,N_4647);
nand U6964 (N_6964,N_3659,N_3466);
and U6965 (N_6965,N_3159,N_3285);
or U6966 (N_6966,N_2710,N_4671);
or U6967 (N_6967,N_4391,N_2965);
and U6968 (N_6968,N_4094,N_2912);
xnor U6969 (N_6969,N_3961,N_4849);
nand U6970 (N_6970,N_3651,N_2774);
or U6971 (N_6971,N_3346,N_3640);
or U6972 (N_6972,N_2625,N_3898);
or U6973 (N_6973,N_4347,N_2977);
xor U6974 (N_6974,N_4333,N_4986);
or U6975 (N_6975,N_3770,N_2510);
or U6976 (N_6976,N_3332,N_4032);
nand U6977 (N_6977,N_3373,N_3648);
or U6978 (N_6978,N_3734,N_2562);
nor U6979 (N_6979,N_4961,N_2747);
or U6980 (N_6980,N_3039,N_2980);
nand U6981 (N_6981,N_2910,N_2699);
and U6982 (N_6982,N_3226,N_2731);
nor U6983 (N_6983,N_4622,N_4253);
and U6984 (N_6984,N_2779,N_3260);
nor U6985 (N_6985,N_4109,N_4626);
nor U6986 (N_6986,N_2525,N_2977);
or U6987 (N_6987,N_2687,N_4238);
nand U6988 (N_6988,N_4934,N_3980);
nor U6989 (N_6989,N_3333,N_2917);
nor U6990 (N_6990,N_3104,N_2519);
and U6991 (N_6991,N_2908,N_2844);
nand U6992 (N_6992,N_2879,N_2635);
nand U6993 (N_6993,N_4949,N_2702);
nand U6994 (N_6994,N_4127,N_4119);
or U6995 (N_6995,N_2800,N_3703);
or U6996 (N_6996,N_4868,N_2697);
nand U6997 (N_6997,N_4091,N_3877);
nor U6998 (N_6998,N_4908,N_3006);
xnor U6999 (N_6999,N_4198,N_4987);
or U7000 (N_7000,N_2864,N_4422);
nor U7001 (N_7001,N_4336,N_4824);
or U7002 (N_7002,N_2972,N_3712);
nand U7003 (N_7003,N_2957,N_3245);
and U7004 (N_7004,N_4114,N_2826);
and U7005 (N_7005,N_3658,N_4309);
nand U7006 (N_7006,N_3013,N_2583);
nor U7007 (N_7007,N_3967,N_4917);
nor U7008 (N_7008,N_3802,N_2514);
and U7009 (N_7009,N_4245,N_3432);
nor U7010 (N_7010,N_3475,N_3301);
xnor U7011 (N_7011,N_3227,N_4451);
nand U7012 (N_7012,N_3085,N_3057);
and U7013 (N_7013,N_4153,N_3712);
nor U7014 (N_7014,N_4665,N_4248);
nand U7015 (N_7015,N_3214,N_3428);
nand U7016 (N_7016,N_4704,N_4270);
nand U7017 (N_7017,N_4320,N_3724);
xor U7018 (N_7018,N_3085,N_3686);
or U7019 (N_7019,N_4693,N_4724);
and U7020 (N_7020,N_4731,N_4086);
and U7021 (N_7021,N_2884,N_4544);
and U7022 (N_7022,N_3607,N_2696);
or U7023 (N_7023,N_3364,N_2534);
nor U7024 (N_7024,N_4244,N_3379);
and U7025 (N_7025,N_3973,N_3554);
nor U7026 (N_7026,N_2588,N_4673);
nor U7027 (N_7027,N_4089,N_2876);
nand U7028 (N_7028,N_2575,N_4141);
nor U7029 (N_7029,N_4792,N_2569);
and U7030 (N_7030,N_3638,N_4548);
and U7031 (N_7031,N_4489,N_4285);
or U7032 (N_7032,N_3028,N_4091);
or U7033 (N_7033,N_4942,N_4258);
or U7034 (N_7034,N_2537,N_3510);
nor U7035 (N_7035,N_3781,N_3091);
or U7036 (N_7036,N_4915,N_4232);
and U7037 (N_7037,N_4731,N_2977);
nor U7038 (N_7038,N_3533,N_2638);
nand U7039 (N_7039,N_4116,N_4859);
nand U7040 (N_7040,N_2569,N_3478);
or U7041 (N_7041,N_3835,N_2780);
nor U7042 (N_7042,N_2957,N_3835);
and U7043 (N_7043,N_4083,N_4281);
and U7044 (N_7044,N_3397,N_4064);
and U7045 (N_7045,N_3311,N_4871);
nor U7046 (N_7046,N_4633,N_4420);
and U7047 (N_7047,N_4018,N_2955);
nand U7048 (N_7048,N_4366,N_4785);
or U7049 (N_7049,N_4610,N_2713);
and U7050 (N_7050,N_3769,N_4090);
or U7051 (N_7051,N_4055,N_4069);
nand U7052 (N_7052,N_4748,N_3645);
or U7053 (N_7053,N_2841,N_3128);
nand U7054 (N_7054,N_2684,N_3763);
nand U7055 (N_7055,N_3674,N_4685);
and U7056 (N_7056,N_4591,N_3168);
or U7057 (N_7057,N_3449,N_3477);
and U7058 (N_7058,N_3463,N_4001);
and U7059 (N_7059,N_4989,N_2703);
nor U7060 (N_7060,N_2991,N_4169);
and U7061 (N_7061,N_3724,N_3734);
nor U7062 (N_7062,N_3635,N_4745);
and U7063 (N_7063,N_2644,N_4402);
or U7064 (N_7064,N_3626,N_2664);
and U7065 (N_7065,N_4434,N_4600);
xor U7066 (N_7066,N_3281,N_3718);
nor U7067 (N_7067,N_3749,N_4649);
nand U7068 (N_7068,N_3636,N_4464);
nor U7069 (N_7069,N_2784,N_4528);
nand U7070 (N_7070,N_3534,N_3301);
nand U7071 (N_7071,N_3781,N_3256);
nand U7072 (N_7072,N_4088,N_2977);
and U7073 (N_7073,N_2839,N_3300);
and U7074 (N_7074,N_4869,N_3362);
or U7075 (N_7075,N_2996,N_4595);
nor U7076 (N_7076,N_4886,N_4854);
nor U7077 (N_7077,N_4556,N_3284);
nand U7078 (N_7078,N_4519,N_4587);
nand U7079 (N_7079,N_4876,N_2794);
nor U7080 (N_7080,N_2516,N_3495);
nand U7081 (N_7081,N_4962,N_4456);
or U7082 (N_7082,N_3275,N_4228);
nand U7083 (N_7083,N_2676,N_4785);
nand U7084 (N_7084,N_2937,N_4295);
nand U7085 (N_7085,N_3829,N_3193);
nor U7086 (N_7086,N_4801,N_3714);
nor U7087 (N_7087,N_3370,N_2804);
and U7088 (N_7088,N_3179,N_3682);
nor U7089 (N_7089,N_3809,N_3141);
and U7090 (N_7090,N_4217,N_2623);
nor U7091 (N_7091,N_4745,N_4393);
and U7092 (N_7092,N_4749,N_3367);
nor U7093 (N_7093,N_3628,N_2699);
xnor U7094 (N_7094,N_4484,N_3557);
nor U7095 (N_7095,N_3067,N_4185);
or U7096 (N_7096,N_4410,N_3977);
and U7097 (N_7097,N_2803,N_4003);
or U7098 (N_7098,N_4659,N_2587);
or U7099 (N_7099,N_3521,N_2961);
or U7100 (N_7100,N_3159,N_3791);
nor U7101 (N_7101,N_3467,N_4072);
nand U7102 (N_7102,N_3119,N_4277);
and U7103 (N_7103,N_3249,N_4645);
nand U7104 (N_7104,N_3823,N_3304);
xnor U7105 (N_7105,N_4568,N_4552);
or U7106 (N_7106,N_2873,N_2693);
or U7107 (N_7107,N_4300,N_4621);
or U7108 (N_7108,N_3665,N_3614);
nor U7109 (N_7109,N_3405,N_3667);
or U7110 (N_7110,N_4741,N_3472);
or U7111 (N_7111,N_4674,N_3033);
or U7112 (N_7112,N_2914,N_3605);
or U7113 (N_7113,N_3039,N_4380);
or U7114 (N_7114,N_4136,N_4274);
nor U7115 (N_7115,N_4906,N_4657);
and U7116 (N_7116,N_3840,N_3165);
nand U7117 (N_7117,N_4959,N_3958);
nand U7118 (N_7118,N_3587,N_3304);
nor U7119 (N_7119,N_4810,N_3270);
nor U7120 (N_7120,N_4360,N_3507);
nand U7121 (N_7121,N_4340,N_4832);
and U7122 (N_7122,N_3504,N_3723);
or U7123 (N_7123,N_4053,N_3179);
nor U7124 (N_7124,N_3673,N_2936);
and U7125 (N_7125,N_4077,N_3645);
or U7126 (N_7126,N_4776,N_3162);
or U7127 (N_7127,N_3188,N_3276);
xor U7128 (N_7128,N_4058,N_4375);
and U7129 (N_7129,N_2826,N_3249);
nor U7130 (N_7130,N_4460,N_2505);
nor U7131 (N_7131,N_4232,N_3209);
or U7132 (N_7132,N_4258,N_3741);
and U7133 (N_7133,N_2552,N_3417);
nand U7134 (N_7134,N_2870,N_3129);
nor U7135 (N_7135,N_3044,N_2567);
and U7136 (N_7136,N_4439,N_3965);
nand U7137 (N_7137,N_4000,N_4450);
nor U7138 (N_7138,N_4054,N_2991);
nor U7139 (N_7139,N_2792,N_2781);
or U7140 (N_7140,N_3710,N_4511);
and U7141 (N_7141,N_3434,N_3209);
and U7142 (N_7142,N_3264,N_3178);
or U7143 (N_7143,N_3611,N_3953);
or U7144 (N_7144,N_4881,N_3515);
nor U7145 (N_7145,N_3216,N_3896);
nor U7146 (N_7146,N_3738,N_3306);
nor U7147 (N_7147,N_2587,N_3969);
and U7148 (N_7148,N_4293,N_2952);
and U7149 (N_7149,N_3359,N_2616);
nand U7150 (N_7150,N_4278,N_3641);
and U7151 (N_7151,N_3164,N_2920);
and U7152 (N_7152,N_4184,N_4516);
nand U7153 (N_7153,N_3187,N_4169);
nand U7154 (N_7154,N_3791,N_4237);
nor U7155 (N_7155,N_4263,N_2802);
xor U7156 (N_7156,N_3853,N_3574);
or U7157 (N_7157,N_4937,N_3682);
and U7158 (N_7158,N_4446,N_2737);
or U7159 (N_7159,N_4467,N_4270);
and U7160 (N_7160,N_4767,N_4918);
and U7161 (N_7161,N_3514,N_3531);
nand U7162 (N_7162,N_4559,N_3953);
or U7163 (N_7163,N_4444,N_3921);
nor U7164 (N_7164,N_3526,N_3034);
nor U7165 (N_7165,N_4609,N_4735);
nand U7166 (N_7166,N_4286,N_2736);
or U7167 (N_7167,N_4092,N_3705);
or U7168 (N_7168,N_2984,N_3656);
nor U7169 (N_7169,N_3472,N_4145);
and U7170 (N_7170,N_2670,N_4328);
or U7171 (N_7171,N_3730,N_3285);
and U7172 (N_7172,N_2776,N_3371);
nand U7173 (N_7173,N_3159,N_4243);
and U7174 (N_7174,N_4698,N_3030);
nand U7175 (N_7175,N_2786,N_2905);
nand U7176 (N_7176,N_4715,N_4738);
and U7177 (N_7177,N_4675,N_4481);
nand U7178 (N_7178,N_3408,N_2794);
or U7179 (N_7179,N_3505,N_4468);
nand U7180 (N_7180,N_4472,N_2804);
nor U7181 (N_7181,N_2564,N_3695);
or U7182 (N_7182,N_2521,N_3805);
or U7183 (N_7183,N_3444,N_4025);
nand U7184 (N_7184,N_2923,N_4852);
and U7185 (N_7185,N_3701,N_2532);
and U7186 (N_7186,N_3019,N_2618);
nand U7187 (N_7187,N_3730,N_4121);
nand U7188 (N_7188,N_3320,N_4148);
or U7189 (N_7189,N_4234,N_3615);
or U7190 (N_7190,N_3045,N_2839);
or U7191 (N_7191,N_4624,N_3558);
and U7192 (N_7192,N_4085,N_2865);
and U7193 (N_7193,N_3526,N_4713);
nand U7194 (N_7194,N_3414,N_4133);
nand U7195 (N_7195,N_4371,N_4448);
or U7196 (N_7196,N_4113,N_3370);
nor U7197 (N_7197,N_2888,N_2756);
and U7198 (N_7198,N_4654,N_3836);
nor U7199 (N_7199,N_2711,N_3378);
nand U7200 (N_7200,N_3042,N_4515);
nand U7201 (N_7201,N_3433,N_2517);
and U7202 (N_7202,N_3302,N_2562);
and U7203 (N_7203,N_4955,N_3373);
or U7204 (N_7204,N_3704,N_4445);
and U7205 (N_7205,N_3877,N_4544);
nand U7206 (N_7206,N_2935,N_3281);
nor U7207 (N_7207,N_3376,N_3259);
nand U7208 (N_7208,N_4732,N_3181);
or U7209 (N_7209,N_3412,N_3480);
nor U7210 (N_7210,N_4190,N_3868);
or U7211 (N_7211,N_2913,N_4099);
nand U7212 (N_7212,N_4912,N_4604);
and U7213 (N_7213,N_3730,N_3337);
and U7214 (N_7214,N_4898,N_3758);
nor U7215 (N_7215,N_3914,N_3108);
xor U7216 (N_7216,N_3997,N_4561);
nand U7217 (N_7217,N_2610,N_3807);
nand U7218 (N_7218,N_3627,N_3267);
nor U7219 (N_7219,N_2877,N_3832);
nor U7220 (N_7220,N_4040,N_2600);
nand U7221 (N_7221,N_4803,N_4168);
and U7222 (N_7222,N_4254,N_2881);
xor U7223 (N_7223,N_3562,N_3189);
and U7224 (N_7224,N_2806,N_4251);
nor U7225 (N_7225,N_3939,N_4988);
nor U7226 (N_7226,N_3666,N_4261);
or U7227 (N_7227,N_4721,N_3570);
nand U7228 (N_7228,N_4315,N_2740);
and U7229 (N_7229,N_3103,N_4546);
or U7230 (N_7230,N_3151,N_4148);
or U7231 (N_7231,N_4969,N_3779);
nor U7232 (N_7232,N_3847,N_4674);
or U7233 (N_7233,N_2677,N_4214);
nand U7234 (N_7234,N_3844,N_3984);
or U7235 (N_7235,N_3948,N_3536);
nor U7236 (N_7236,N_3514,N_4423);
and U7237 (N_7237,N_4208,N_4840);
xor U7238 (N_7238,N_3537,N_3545);
and U7239 (N_7239,N_3109,N_4429);
nor U7240 (N_7240,N_4577,N_4474);
xnor U7241 (N_7241,N_2945,N_3445);
and U7242 (N_7242,N_2910,N_4217);
nand U7243 (N_7243,N_2863,N_3191);
or U7244 (N_7244,N_4671,N_2759);
nand U7245 (N_7245,N_4293,N_3000);
and U7246 (N_7246,N_2600,N_4658);
nand U7247 (N_7247,N_3801,N_4341);
and U7248 (N_7248,N_4827,N_4044);
and U7249 (N_7249,N_4049,N_3386);
nand U7250 (N_7250,N_2573,N_3362);
or U7251 (N_7251,N_3968,N_3318);
nand U7252 (N_7252,N_4031,N_2558);
or U7253 (N_7253,N_3986,N_4436);
nor U7254 (N_7254,N_4638,N_2720);
or U7255 (N_7255,N_3714,N_4371);
nand U7256 (N_7256,N_4958,N_3464);
and U7257 (N_7257,N_2799,N_2584);
or U7258 (N_7258,N_3826,N_4438);
and U7259 (N_7259,N_4470,N_2505);
or U7260 (N_7260,N_4933,N_2523);
nor U7261 (N_7261,N_2976,N_4983);
and U7262 (N_7262,N_4126,N_4313);
and U7263 (N_7263,N_2748,N_3114);
nor U7264 (N_7264,N_2871,N_4782);
nor U7265 (N_7265,N_4834,N_3882);
or U7266 (N_7266,N_4459,N_3850);
nand U7267 (N_7267,N_4625,N_4026);
and U7268 (N_7268,N_3202,N_2584);
nand U7269 (N_7269,N_3015,N_4010);
nand U7270 (N_7270,N_2653,N_4904);
nor U7271 (N_7271,N_4722,N_2963);
nor U7272 (N_7272,N_3516,N_2859);
and U7273 (N_7273,N_3171,N_3042);
nor U7274 (N_7274,N_4836,N_3150);
nand U7275 (N_7275,N_3555,N_4825);
and U7276 (N_7276,N_3036,N_3553);
nand U7277 (N_7277,N_3190,N_3014);
nand U7278 (N_7278,N_4409,N_3157);
nor U7279 (N_7279,N_4375,N_4305);
or U7280 (N_7280,N_2788,N_3132);
nor U7281 (N_7281,N_4988,N_4768);
nor U7282 (N_7282,N_3817,N_2995);
or U7283 (N_7283,N_2849,N_4044);
nand U7284 (N_7284,N_3822,N_4625);
nor U7285 (N_7285,N_4216,N_3052);
nor U7286 (N_7286,N_3026,N_4940);
and U7287 (N_7287,N_4387,N_3917);
nand U7288 (N_7288,N_3326,N_4792);
or U7289 (N_7289,N_4947,N_4116);
nand U7290 (N_7290,N_3270,N_4630);
or U7291 (N_7291,N_3136,N_4935);
or U7292 (N_7292,N_3352,N_4373);
and U7293 (N_7293,N_3266,N_3322);
and U7294 (N_7294,N_3359,N_2733);
nor U7295 (N_7295,N_3164,N_4991);
xor U7296 (N_7296,N_3377,N_3514);
and U7297 (N_7297,N_2898,N_2658);
or U7298 (N_7298,N_4211,N_3379);
nand U7299 (N_7299,N_3148,N_2529);
and U7300 (N_7300,N_4727,N_3716);
nor U7301 (N_7301,N_3358,N_4821);
xor U7302 (N_7302,N_3548,N_3160);
or U7303 (N_7303,N_3198,N_2981);
and U7304 (N_7304,N_2990,N_3469);
or U7305 (N_7305,N_4008,N_2649);
or U7306 (N_7306,N_3888,N_3083);
or U7307 (N_7307,N_2974,N_3213);
nand U7308 (N_7308,N_4651,N_4418);
nor U7309 (N_7309,N_3926,N_3273);
nor U7310 (N_7310,N_4870,N_4757);
or U7311 (N_7311,N_4633,N_2999);
or U7312 (N_7312,N_4867,N_3692);
nand U7313 (N_7313,N_3895,N_2959);
nor U7314 (N_7314,N_3039,N_4378);
nand U7315 (N_7315,N_3269,N_4867);
nor U7316 (N_7316,N_4125,N_2535);
and U7317 (N_7317,N_3769,N_4731);
nand U7318 (N_7318,N_4740,N_2839);
or U7319 (N_7319,N_2535,N_4002);
nor U7320 (N_7320,N_3331,N_4525);
or U7321 (N_7321,N_3140,N_3428);
or U7322 (N_7322,N_4548,N_4830);
and U7323 (N_7323,N_2974,N_4739);
and U7324 (N_7324,N_4348,N_4006);
nor U7325 (N_7325,N_4687,N_2861);
and U7326 (N_7326,N_3902,N_4801);
nor U7327 (N_7327,N_4339,N_4575);
nor U7328 (N_7328,N_2598,N_4602);
nor U7329 (N_7329,N_3831,N_3773);
and U7330 (N_7330,N_4073,N_3208);
and U7331 (N_7331,N_4679,N_3568);
nor U7332 (N_7332,N_3364,N_4387);
and U7333 (N_7333,N_3667,N_2903);
or U7334 (N_7334,N_3813,N_2507);
and U7335 (N_7335,N_4294,N_3002);
or U7336 (N_7336,N_4467,N_3128);
or U7337 (N_7337,N_4418,N_4010);
nor U7338 (N_7338,N_3671,N_4832);
or U7339 (N_7339,N_2802,N_3601);
and U7340 (N_7340,N_4132,N_3986);
nand U7341 (N_7341,N_3752,N_3484);
nor U7342 (N_7342,N_3444,N_4987);
nand U7343 (N_7343,N_3609,N_4689);
nand U7344 (N_7344,N_3367,N_2977);
nand U7345 (N_7345,N_3003,N_2995);
and U7346 (N_7346,N_4471,N_2637);
nor U7347 (N_7347,N_3237,N_3040);
and U7348 (N_7348,N_4824,N_3531);
nand U7349 (N_7349,N_2849,N_4759);
and U7350 (N_7350,N_2807,N_3638);
or U7351 (N_7351,N_3592,N_3974);
nor U7352 (N_7352,N_3053,N_4909);
nor U7353 (N_7353,N_2607,N_3715);
nor U7354 (N_7354,N_3470,N_4955);
nand U7355 (N_7355,N_3220,N_3147);
and U7356 (N_7356,N_3902,N_4877);
nor U7357 (N_7357,N_3810,N_4334);
and U7358 (N_7358,N_4378,N_4947);
nand U7359 (N_7359,N_2579,N_4015);
nor U7360 (N_7360,N_4290,N_3830);
nor U7361 (N_7361,N_3215,N_4421);
or U7362 (N_7362,N_3453,N_2668);
nor U7363 (N_7363,N_4038,N_4789);
nor U7364 (N_7364,N_3906,N_2779);
nand U7365 (N_7365,N_2676,N_4465);
and U7366 (N_7366,N_4431,N_4615);
nand U7367 (N_7367,N_4009,N_3319);
and U7368 (N_7368,N_2628,N_4788);
or U7369 (N_7369,N_3300,N_4911);
nor U7370 (N_7370,N_3514,N_4669);
or U7371 (N_7371,N_3529,N_4632);
and U7372 (N_7372,N_3931,N_4311);
xnor U7373 (N_7373,N_3904,N_2971);
nor U7374 (N_7374,N_2711,N_3158);
or U7375 (N_7375,N_4926,N_4463);
and U7376 (N_7376,N_2964,N_2825);
or U7377 (N_7377,N_2539,N_3911);
nand U7378 (N_7378,N_4077,N_3826);
nor U7379 (N_7379,N_4723,N_4664);
nand U7380 (N_7380,N_2746,N_4269);
nand U7381 (N_7381,N_4612,N_4911);
and U7382 (N_7382,N_4050,N_3000);
nand U7383 (N_7383,N_3572,N_3926);
xor U7384 (N_7384,N_4753,N_4257);
and U7385 (N_7385,N_3332,N_4726);
xor U7386 (N_7386,N_3719,N_3180);
and U7387 (N_7387,N_4902,N_2811);
nor U7388 (N_7388,N_3602,N_3516);
nor U7389 (N_7389,N_2714,N_4111);
nor U7390 (N_7390,N_2934,N_2501);
nor U7391 (N_7391,N_3729,N_2545);
nand U7392 (N_7392,N_3053,N_3879);
nor U7393 (N_7393,N_3534,N_2633);
or U7394 (N_7394,N_4412,N_4797);
or U7395 (N_7395,N_3016,N_4434);
and U7396 (N_7396,N_3788,N_3938);
and U7397 (N_7397,N_4150,N_2837);
nand U7398 (N_7398,N_3619,N_3140);
and U7399 (N_7399,N_4431,N_4952);
or U7400 (N_7400,N_2758,N_4095);
or U7401 (N_7401,N_4007,N_3520);
and U7402 (N_7402,N_4484,N_4302);
or U7403 (N_7403,N_3539,N_3589);
nor U7404 (N_7404,N_4603,N_2896);
and U7405 (N_7405,N_4762,N_2574);
or U7406 (N_7406,N_3387,N_2794);
nand U7407 (N_7407,N_4105,N_2543);
or U7408 (N_7408,N_4737,N_4854);
and U7409 (N_7409,N_3189,N_3873);
or U7410 (N_7410,N_2581,N_3851);
or U7411 (N_7411,N_3646,N_3315);
and U7412 (N_7412,N_3737,N_3450);
xor U7413 (N_7413,N_2815,N_3587);
nand U7414 (N_7414,N_2877,N_3417);
and U7415 (N_7415,N_4161,N_3440);
nand U7416 (N_7416,N_4868,N_4635);
nand U7417 (N_7417,N_4602,N_4319);
nor U7418 (N_7418,N_4471,N_4697);
nand U7419 (N_7419,N_4201,N_3756);
nor U7420 (N_7420,N_3076,N_2970);
nand U7421 (N_7421,N_3628,N_3844);
and U7422 (N_7422,N_3137,N_3051);
nand U7423 (N_7423,N_2887,N_3485);
nand U7424 (N_7424,N_4231,N_4844);
nor U7425 (N_7425,N_2564,N_3520);
or U7426 (N_7426,N_2580,N_3176);
or U7427 (N_7427,N_3834,N_4909);
nor U7428 (N_7428,N_4170,N_4556);
and U7429 (N_7429,N_4983,N_4755);
and U7430 (N_7430,N_4188,N_4245);
or U7431 (N_7431,N_4060,N_4533);
nand U7432 (N_7432,N_4146,N_2623);
nor U7433 (N_7433,N_3937,N_4396);
and U7434 (N_7434,N_3878,N_4020);
and U7435 (N_7435,N_4441,N_4077);
and U7436 (N_7436,N_4181,N_2720);
nand U7437 (N_7437,N_2951,N_3775);
nand U7438 (N_7438,N_2744,N_4615);
or U7439 (N_7439,N_2617,N_4591);
xnor U7440 (N_7440,N_4843,N_2904);
and U7441 (N_7441,N_3364,N_3615);
nor U7442 (N_7442,N_3015,N_4791);
or U7443 (N_7443,N_3001,N_2748);
nor U7444 (N_7444,N_2989,N_4314);
nor U7445 (N_7445,N_2652,N_3765);
and U7446 (N_7446,N_4672,N_4360);
and U7447 (N_7447,N_4317,N_4734);
nor U7448 (N_7448,N_3087,N_4966);
nand U7449 (N_7449,N_3923,N_2538);
nand U7450 (N_7450,N_3734,N_2523);
nor U7451 (N_7451,N_4607,N_4369);
nand U7452 (N_7452,N_4177,N_4441);
nor U7453 (N_7453,N_3968,N_2597);
nand U7454 (N_7454,N_4657,N_3276);
or U7455 (N_7455,N_3800,N_3926);
or U7456 (N_7456,N_4918,N_4385);
nor U7457 (N_7457,N_4033,N_3530);
nand U7458 (N_7458,N_2599,N_3802);
nand U7459 (N_7459,N_4013,N_4204);
nand U7460 (N_7460,N_2950,N_4718);
nor U7461 (N_7461,N_4932,N_2926);
nand U7462 (N_7462,N_3989,N_2878);
nor U7463 (N_7463,N_4666,N_3487);
nor U7464 (N_7464,N_4012,N_3633);
and U7465 (N_7465,N_4115,N_2587);
and U7466 (N_7466,N_4100,N_2629);
and U7467 (N_7467,N_3803,N_4791);
xnor U7468 (N_7468,N_2631,N_3948);
nor U7469 (N_7469,N_4270,N_4477);
nor U7470 (N_7470,N_3724,N_2870);
and U7471 (N_7471,N_4485,N_4254);
nand U7472 (N_7472,N_3704,N_3088);
or U7473 (N_7473,N_3069,N_2808);
nor U7474 (N_7474,N_3480,N_4226);
or U7475 (N_7475,N_4242,N_2784);
or U7476 (N_7476,N_4347,N_3103);
nand U7477 (N_7477,N_3722,N_2731);
nor U7478 (N_7478,N_3853,N_2712);
nor U7479 (N_7479,N_4383,N_3557);
nor U7480 (N_7480,N_4070,N_4535);
nor U7481 (N_7481,N_4035,N_3819);
nor U7482 (N_7482,N_3255,N_3946);
and U7483 (N_7483,N_4928,N_4088);
nand U7484 (N_7484,N_4079,N_3250);
or U7485 (N_7485,N_4989,N_4836);
nor U7486 (N_7486,N_2721,N_4797);
and U7487 (N_7487,N_4413,N_2676);
and U7488 (N_7488,N_4411,N_3089);
and U7489 (N_7489,N_3653,N_4506);
nand U7490 (N_7490,N_4906,N_4695);
or U7491 (N_7491,N_2944,N_3529);
or U7492 (N_7492,N_4410,N_4242);
nor U7493 (N_7493,N_2725,N_2852);
and U7494 (N_7494,N_3958,N_2932);
nor U7495 (N_7495,N_3689,N_2965);
nor U7496 (N_7496,N_3301,N_3847);
nor U7497 (N_7497,N_4820,N_2948);
or U7498 (N_7498,N_3582,N_3237);
nand U7499 (N_7499,N_4388,N_4076);
nor U7500 (N_7500,N_6979,N_6550);
or U7501 (N_7501,N_6398,N_7077);
or U7502 (N_7502,N_5190,N_6909);
nor U7503 (N_7503,N_6506,N_5181);
and U7504 (N_7504,N_5819,N_6004);
and U7505 (N_7505,N_6110,N_5132);
nor U7506 (N_7506,N_7371,N_6719);
and U7507 (N_7507,N_5827,N_6799);
or U7508 (N_7508,N_7280,N_6540);
nor U7509 (N_7509,N_6793,N_5216);
or U7510 (N_7510,N_6744,N_7224);
nor U7511 (N_7511,N_6235,N_5406);
nor U7512 (N_7512,N_5022,N_6310);
nand U7513 (N_7513,N_7347,N_5995);
xor U7514 (N_7514,N_5336,N_5062);
nor U7515 (N_7515,N_5722,N_7042);
and U7516 (N_7516,N_6162,N_6094);
or U7517 (N_7517,N_6949,N_6479);
nand U7518 (N_7518,N_6671,N_7311);
or U7519 (N_7519,N_6127,N_5385);
nor U7520 (N_7520,N_5854,N_7226);
or U7521 (N_7521,N_6493,N_6111);
and U7522 (N_7522,N_6301,N_6902);
nor U7523 (N_7523,N_5294,N_5528);
nor U7524 (N_7524,N_6866,N_5665);
or U7525 (N_7525,N_7382,N_7205);
nand U7526 (N_7526,N_6495,N_7143);
and U7527 (N_7527,N_5456,N_5471);
nor U7528 (N_7528,N_7272,N_6831);
or U7529 (N_7529,N_6581,N_5851);
nor U7530 (N_7530,N_6203,N_6698);
and U7531 (N_7531,N_5772,N_6922);
nor U7532 (N_7532,N_5979,N_5400);
or U7533 (N_7533,N_6832,N_6354);
or U7534 (N_7534,N_7370,N_7207);
and U7535 (N_7535,N_6780,N_6429);
or U7536 (N_7536,N_6346,N_7297);
or U7537 (N_7537,N_5185,N_6112);
nor U7538 (N_7538,N_5726,N_6234);
or U7539 (N_7539,N_6473,N_5978);
and U7540 (N_7540,N_7255,N_6408);
or U7541 (N_7541,N_6779,N_6239);
nor U7542 (N_7542,N_5554,N_6841);
nand U7543 (N_7543,N_6500,N_5694);
and U7544 (N_7544,N_5501,N_5170);
or U7545 (N_7545,N_6747,N_6328);
nor U7546 (N_7546,N_5041,N_5834);
nor U7547 (N_7547,N_5291,N_6659);
or U7548 (N_7548,N_5455,N_5850);
nand U7549 (N_7549,N_7088,N_5478);
nand U7550 (N_7550,N_7283,N_6789);
nor U7551 (N_7551,N_6341,N_6131);
nand U7552 (N_7552,N_7436,N_5201);
nor U7553 (N_7553,N_6851,N_7173);
nor U7554 (N_7554,N_6293,N_5522);
nor U7555 (N_7555,N_6017,N_5929);
or U7556 (N_7556,N_6694,N_5713);
or U7557 (N_7557,N_6674,N_5133);
or U7558 (N_7558,N_5167,N_7444);
and U7559 (N_7559,N_5441,N_6802);
or U7560 (N_7560,N_5561,N_5240);
nor U7561 (N_7561,N_7117,N_6236);
or U7562 (N_7562,N_6844,N_6058);
nand U7563 (N_7563,N_7355,N_7149);
nand U7564 (N_7564,N_7246,N_7467);
nand U7565 (N_7565,N_5731,N_7136);
or U7566 (N_7566,N_6191,N_5231);
and U7567 (N_7567,N_5050,N_5865);
nor U7568 (N_7568,N_7217,N_5923);
or U7569 (N_7569,N_6396,N_7485);
or U7570 (N_7570,N_6304,N_7235);
and U7571 (N_7571,N_6758,N_6374);
nand U7572 (N_7572,N_6284,N_5119);
or U7573 (N_7573,N_6483,N_7102);
nand U7574 (N_7574,N_6032,N_6044);
or U7575 (N_7575,N_7164,N_6957);
or U7576 (N_7576,N_5335,N_6726);
and U7577 (N_7577,N_7270,N_5176);
nor U7578 (N_7578,N_5241,N_6942);
nand U7579 (N_7579,N_6040,N_6247);
and U7580 (N_7580,N_7429,N_6880);
and U7581 (N_7581,N_5072,N_6063);
or U7582 (N_7582,N_5435,N_6580);
nand U7583 (N_7583,N_5810,N_5540);
nand U7584 (N_7584,N_5826,N_5272);
and U7585 (N_7585,N_5005,N_6045);
xnor U7586 (N_7586,N_6418,N_5642);
nor U7587 (N_7587,N_6097,N_7031);
or U7588 (N_7588,N_7144,N_6065);
nand U7589 (N_7589,N_5958,N_5303);
nand U7590 (N_7590,N_6353,N_5996);
nor U7591 (N_7591,N_5402,N_5392);
and U7592 (N_7592,N_6382,N_6811);
nand U7593 (N_7593,N_5314,N_6220);
nor U7594 (N_7594,N_6404,N_7397);
nand U7595 (N_7595,N_5643,N_5331);
nor U7596 (N_7596,N_5483,N_6583);
or U7597 (N_7597,N_7212,N_7016);
or U7598 (N_7598,N_6924,N_5001);
and U7599 (N_7599,N_6734,N_6271);
and U7600 (N_7600,N_6971,N_6068);
nor U7601 (N_7601,N_5110,N_5484);
and U7602 (N_7602,N_5841,N_5422);
and U7603 (N_7603,N_6283,N_6255);
nor U7604 (N_7604,N_6120,N_5567);
and U7605 (N_7605,N_5755,N_6945);
and U7606 (N_7606,N_5019,N_5289);
or U7607 (N_7607,N_5320,N_6998);
nand U7608 (N_7608,N_5386,N_7121);
and U7609 (N_7609,N_6415,N_5434);
nor U7610 (N_7610,N_5604,N_5662);
nor U7611 (N_7611,N_5683,N_5278);
nand U7612 (N_7612,N_7021,N_5117);
nor U7613 (N_7613,N_5063,N_6082);
nor U7614 (N_7614,N_5756,N_6960);
nor U7615 (N_7615,N_7474,N_5437);
nand U7616 (N_7616,N_6208,N_7253);
nor U7617 (N_7617,N_5248,N_5079);
and U7618 (N_7618,N_6069,N_6891);
nand U7619 (N_7619,N_7067,N_7400);
and U7620 (N_7620,N_6848,N_5036);
or U7621 (N_7621,N_5616,N_6502);
nor U7622 (N_7622,N_5893,N_5427);
nor U7623 (N_7623,N_5130,N_6253);
or U7624 (N_7624,N_5382,N_6072);
or U7625 (N_7625,N_5351,N_6656);
nor U7626 (N_7626,N_7048,N_6009);
nor U7627 (N_7627,N_5803,N_7247);
nor U7628 (N_7628,N_6826,N_7101);
nand U7629 (N_7629,N_7464,N_5171);
xnor U7630 (N_7630,N_6707,N_7484);
nand U7631 (N_7631,N_5947,N_7133);
nor U7632 (N_7632,N_6636,N_6148);
nor U7633 (N_7633,N_6287,N_6225);
nand U7634 (N_7634,N_5405,N_7038);
nand U7635 (N_7635,N_5749,N_5640);
nor U7636 (N_7636,N_6416,N_7074);
nor U7637 (N_7637,N_6512,N_6307);
and U7638 (N_7638,N_5828,N_6556);
nor U7639 (N_7639,N_7083,N_6198);
or U7640 (N_7640,N_5730,N_6951);
xor U7641 (N_7641,N_7028,N_5074);
nor U7642 (N_7642,N_5966,N_5154);
or U7643 (N_7643,N_7183,N_5907);
and U7644 (N_7644,N_7043,N_7369);
nor U7645 (N_7645,N_7058,N_7229);
nand U7646 (N_7646,N_6143,N_5083);
xnor U7647 (N_7647,N_7137,N_5476);
or U7648 (N_7648,N_5071,N_7119);
and U7649 (N_7649,N_5105,N_5602);
or U7650 (N_7650,N_5225,N_5806);
or U7651 (N_7651,N_5621,N_5428);
nor U7652 (N_7652,N_5473,N_7262);
and U7653 (N_7653,N_7189,N_6917);
or U7654 (N_7654,N_6447,N_7415);
or U7655 (N_7655,N_6970,N_7391);
and U7656 (N_7656,N_7155,N_6845);
or U7657 (N_7657,N_7265,N_7291);
and U7658 (N_7658,N_5268,N_5959);
and U7659 (N_7659,N_7448,N_6913);
nand U7660 (N_7660,N_5757,N_7104);
nor U7661 (N_7661,N_7366,N_6996);
and U7662 (N_7662,N_5077,N_6978);
nand U7663 (N_7663,N_6921,N_5046);
nand U7664 (N_7664,N_5507,N_5477);
nor U7665 (N_7665,N_7326,N_5511);
and U7666 (N_7666,N_6509,N_7378);
nor U7667 (N_7667,N_6810,N_6083);
or U7668 (N_7668,N_6485,N_6003);
nor U7669 (N_7669,N_6625,N_5908);
and U7670 (N_7670,N_6684,N_6272);
nand U7671 (N_7671,N_5932,N_5160);
xnor U7672 (N_7672,N_7336,N_5301);
nor U7673 (N_7673,N_6829,N_6440);
and U7674 (N_7674,N_6603,N_5560);
xor U7675 (N_7675,N_6850,N_7339);
nand U7676 (N_7676,N_5205,N_7142);
nand U7677 (N_7677,N_6592,N_6529);
nor U7678 (N_7678,N_7139,N_7047);
xor U7679 (N_7679,N_6291,N_7196);
and U7680 (N_7680,N_6189,N_5153);
nand U7681 (N_7681,N_7232,N_5344);
nor U7682 (N_7682,N_5358,N_6461);
or U7683 (N_7683,N_5312,N_6676);
nand U7684 (N_7684,N_5080,N_5052);
nand U7685 (N_7685,N_7060,N_6691);
or U7686 (N_7686,N_6815,N_5964);
nand U7687 (N_7687,N_5902,N_6798);
nor U7688 (N_7688,N_6375,N_6643);
nand U7689 (N_7689,N_5054,N_6155);
nand U7690 (N_7690,N_5710,N_5784);
nor U7691 (N_7691,N_7124,N_5218);
nor U7692 (N_7692,N_6977,N_5580);
or U7693 (N_7693,N_5396,N_5124);
and U7694 (N_7694,N_6449,N_7284);
and U7695 (N_7695,N_6167,N_7496);
nand U7696 (N_7696,N_5342,N_6391);
nand U7697 (N_7697,N_6520,N_7040);
or U7698 (N_7698,N_5552,N_5924);
nor U7699 (N_7699,N_5156,N_5967);
nand U7700 (N_7700,N_6916,N_5699);
nor U7701 (N_7701,N_5702,N_6233);
and U7702 (N_7702,N_6202,N_5372);
or U7703 (N_7703,N_7234,N_6890);
nand U7704 (N_7704,N_6649,N_6761);
nor U7705 (N_7705,N_6884,N_7399);
nand U7706 (N_7706,N_5655,N_7440);
nand U7707 (N_7707,N_6149,N_6195);
nor U7708 (N_7708,N_7179,N_6248);
or U7709 (N_7709,N_6604,N_5539);
nand U7710 (N_7710,N_7398,N_7242);
nor U7711 (N_7711,N_5013,N_6788);
nor U7712 (N_7712,N_5686,N_6825);
nand U7713 (N_7713,N_5720,N_5420);
nor U7714 (N_7714,N_6064,N_5692);
nand U7715 (N_7715,N_6268,N_6286);
or U7716 (N_7716,N_7276,N_5585);
and U7717 (N_7717,N_6790,N_5261);
nor U7718 (N_7718,N_5697,N_7071);
or U7719 (N_7719,N_6665,N_5524);
or U7720 (N_7720,N_5273,N_5355);
or U7721 (N_7721,N_7428,N_6941);
or U7722 (N_7722,N_5945,N_6946);
or U7723 (N_7723,N_5230,N_5636);
nor U7724 (N_7724,N_5368,N_6348);
and U7725 (N_7725,N_5251,N_6392);
nand U7726 (N_7726,N_7360,N_6563);
nand U7727 (N_7727,N_6070,N_5998);
nor U7728 (N_7728,N_7432,N_6801);
or U7729 (N_7729,N_5488,N_7035);
nand U7730 (N_7730,N_5039,N_6492);
and U7731 (N_7731,N_5209,N_5546);
and U7732 (N_7732,N_5674,N_5413);
and U7733 (N_7733,N_6709,N_7070);
nor U7734 (N_7734,N_7017,N_6026);
or U7735 (N_7735,N_5265,N_6387);
nand U7736 (N_7736,N_6976,N_7044);
and U7737 (N_7737,N_7446,N_5813);
and U7738 (N_7738,N_5003,N_6530);
nand U7739 (N_7739,N_7037,N_5766);
nor U7740 (N_7740,N_7050,N_6768);
nor U7741 (N_7741,N_7472,N_5974);
nand U7742 (N_7742,N_6480,N_6591);
and U7743 (N_7743,N_6194,N_7252);
nor U7744 (N_7744,N_5418,N_5453);
and U7745 (N_7745,N_5461,N_6096);
or U7746 (N_7746,N_6329,N_6338);
and U7747 (N_7747,N_5364,N_5333);
nand U7748 (N_7748,N_5061,N_6187);
xor U7749 (N_7749,N_7294,N_6538);
or U7750 (N_7750,N_5242,N_7080);
nand U7751 (N_7751,N_5898,N_6190);
or U7752 (N_7752,N_7105,N_6994);
and U7753 (N_7753,N_7129,N_6666);
nand U7754 (N_7754,N_7480,N_6251);
or U7755 (N_7755,N_6242,N_6369);
or U7756 (N_7756,N_7277,N_5513);
nand U7757 (N_7757,N_5419,N_5649);
and U7758 (N_7758,N_6664,N_6489);
nand U7759 (N_7759,N_5693,N_7055);
nand U7760 (N_7760,N_7019,N_6231);
and U7761 (N_7761,N_7064,N_5379);
nand U7762 (N_7762,N_7458,N_6828);
nor U7763 (N_7763,N_5549,N_6739);
nor U7764 (N_7764,N_6836,N_5792);
xor U7765 (N_7765,N_5458,N_5021);
nand U7766 (N_7766,N_6748,N_5323);
nand U7767 (N_7767,N_5147,N_6918);
nand U7768 (N_7768,N_6138,N_5239);
and U7769 (N_7769,N_6200,N_5373);
nand U7770 (N_7770,N_6778,N_6962);
nand U7771 (N_7771,N_6765,N_6224);
nor U7772 (N_7772,N_6572,N_5092);
nor U7773 (N_7773,N_5523,N_5651);
and U7774 (N_7774,N_6337,N_6885);
and U7775 (N_7775,N_6743,N_5660);
or U7776 (N_7776,N_7275,N_5056);
or U7777 (N_7777,N_5421,N_7337);
and U7778 (N_7778,N_5873,N_7309);
or U7779 (N_7779,N_6290,N_7163);
nand U7780 (N_7780,N_5107,N_5903);
xor U7781 (N_7781,N_6751,N_6652);
nor U7782 (N_7782,N_5076,N_5353);
and U7783 (N_7783,N_6372,N_6067);
nor U7784 (N_7784,N_7490,N_6627);
nand U7785 (N_7785,N_5647,N_6335);
and U7786 (N_7786,N_5187,N_7010);
or U7787 (N_7787,N_5040,N_5531);
or U7788 (N_7788,N_6561,N_5360);
nor U7789 (N_7789,N_5606,N_7402);
nor U7790 (N_7790,N_5543,N_5296);
nand U7791 (N_7791,N_6539,N_6088);
nand U7792 (N_7792,N_7271,N_6634);
nor U7793 (N_7793,N_7166,N_7216);
nand U7794 (N_7794,N_5804,N_5768);
and U7795 (N_7795,N_6366,N_7357);
nand U7796 (N_7796,N_6056,N_6370);
nand U7797 (N_7797,N_5569,N_6471);
or U7798 (N_7798,N_5222,N_5744);
nor U7799 (N_7799,N_7195,N_6688);
nand U7800 (N_7800,N_5809,N_6725);
nor U7801 (N_7801,N_5948,N_5397);
or U7802 (N_7802,N_5238,N_5760);
and U7803 (N_7803,N_7286,N_5563);
nand U7804 (N_7804,N_5214,N_5442);
and U7805 (N_7805,N_6077,N_5440);
nor U7806 (N_7806,N_5093,N_5696);
or U7807 (N_7807,N_5479,N_6711);
or U7808 (N_7808,N_5404,N_5029);
nor U7809 (N_7809,N_5310,N_5460);
or U7810 (N_7810,N_5790,N_6029);
nand U7811 (N_7811,N_6002,N_5118);
nor U7812 (N_7812,N_6042,N_6582);
nor U7813 (N_7813,N_6930,N_5260);
nor U7814 (N_7814,N_5078,N_6318);
nand U7815 (N_7815,N_5431,N_6967);
nand U7816 (N_7816,N_7111,N_6767);
and U7817 (N_7817,N_7424,N_6617);
or U7818 (N_7818,N_6755,N_7061);
or U7819 (N_7819,N_6873,N_5994);
nor U7820 (N_7820,N_5391,N_6481);
nand U7821 (N_7821,N_6632,N_5700);
and U7822 (N_7822,N_6608,N_7085);
and U7823 (N_7823,N_7220,N_7239);
nor U7824 (N_7824,N_5858,N_6669);
and U7825 (N_7825,N_6423,N_5591);
or U7826 (N_7826,N_6470,N_7175);
nor U7827 (N_7827,N_6727,N_6730);
nor U7828 (N_7828,N_6847,N_7045);
nand U7829 (N_7829,N_6452,N_7123);
xor U7830 (N_7830,N_5394,N_6785);
nand U7831 (N_7831,N_6223,N_5055);
and U7832 (N_7832,N_5250,N_6215);
or U7833 (N_7833,N_6651,N_5367);
or U7834 (N_7834,N_7443,N_6319);
or U7835 (N_7835,N_6153,N_6313);
nand U7836 (N_7836,N_6935,N_6543);
and U7837 (N_7837,N_7498,N_6007);
and U7838 (N_7838,N_7321,N_5459);
or U7839 (N_7839,N_7346,N_7052);
nor U7840 (N_7840,N_6555,N_6670);
nor U7841 (N_7841,N_5904,N_5123);
or U7842 (N_7842,N_6079,N_5840);
and U7843 (N_7843,N_5375,N_6618);
nand U7844 (N_7844,N_5166,N_6264);
and U7845 (N_7845,N_7245,N_5293);
or U7846 (N_7846,N_6459,N_6358);
nor U7847 (N_7847,N_6380,N_6330);
and U7848 (N_7848,N_5877,N_5545);
and U7849 (N_7849,N_6451,N_5457);
nor U7850 (N_7850,N_6275,N_5691);
and U7851 (N_7851,N_7118,N_6180);
nand U7852 (N_7852,N_6438,N_5112);
nand U7853 (N_7853,N_7086,N_5617);
and U7854 (N_7854,N_6516,N_6701);
nand U7855 (N_7855,N_5255,N_6588);
nand U7856 (N_7856,N_5253,N_5941);
nand U7857 (N_7857,N_5783,N_5298);
or U7858 (N_7858,N_5551,N_6134);
nand U7859 (N_7859,N_6124,N_6457);
nor U7860 (N_7860,N_5416,N_6812);
and U7861 (N_7861,N_7034,N_6428);
nand U7862 (N_7862,N_5952,N_5263);
or U7863 (N_7863,N_7026,N_6433);
nand U7864 (N_7864,N_7109,N_5014);
nand U7865 (N_7865,N_5605,N_5277);
nand U7866 (N_7866,N_6532,N_6658);
and U7867 (N_7867,N_6560,N_6524);
nand U7868 (N_7868,N_6679,N_6322);
nand U7869 (N_7869,N_6278,N_6724);
or U7870 (N_7870,N_5829,N_7332);
nor U7871 (N_7871,N_5085,N_7076);
nand U7872 (N_7872,N_5403,N_5856);
or U7873 (N_7873,N_5454,N_5279);
nand U7874 (N_7874,N_7329,N_6037);
or U7875 (N_7875,N_6590,N_6997);
and U7876 (N_7876,N_6795,N_7385);
and U7877 (N_7877,N_7230,N_5109);
nor U7878 (N_7878,N_6175,N_5191);
nor U7879 (N_7879,N_5347,N_5499);
nor U7880 (N_7880,N_7204,N_7198);
nor U7881 (N_7881,N_6872,N_5000);
nor U7882 (N_7882,N_6887,N_6259);
nor U7883 (N_7883,N_5064,N_6963);
and U7884 (N_7884,N_5571,N_5350);
nand U7885 (N_7885,N_6490,N_7174);
nor U7886 (N_7886,N_6075,N_5818);
and U7887 (N_7887,N_5960,N_6186);
or U7888 (N_7888,N_5969,N_5228);
nand U7889 (N_7889,N_5598,N_5884);
or U7890 (N_7890,N_5175,N_6548);
or U7891 (N_7891,N_6397,N_6171);
nor U7892 (N_7892,N_6549,N_5433);
or U7893 (N_7893,N_7159,N_5704);
or U7894 (N_7894,N_7301,N_6606);
or U7895 (N_7895,N_5550,N_6061);
nor U7896 (N_7896,N_5234,N_5808);
and U7897 (N_7897,N_7184,N_6388);
nor U7898 (N_7898,N_5653,N_5822);
and U7899 (N_7899,N_6274,N_7299);
and U7900 (N_7900,N_7348,N_6105);
nor U7901 (N_7901,N_6914,N_7338);
nand U7902 (N_7902,N_5800,N_6702);
nand U7903 (N_7903,N_5305,N_6434);
and U7904 (N_7904,N_6518,N_5915);
nor U7905 (N_7905,N_6868,N_6568);
or U7906 (N_7906,N_5938,N_6325);
or U7907 (N_7907,N_6905,N_7425);
nor U7908 (N_7908,N_6972,N_6262);
nand U7909 (N_7909,N_5346,N_6653);
nor U7910 (N_7910,N_5680,N_5716);
or U7911 (N_7911,N_6115,N_7219);
nor U7912 (N_7912,N_6280,N_6787);
or U7913 (N_7913,N_6491,N_7463);
nor U7914 (N_7914,N_6376,N_6409);
or U7915 (N_7915,N_5538,N_5006);
nand U7916 (N_7916,N_5180,N_5332);
or U7917 (N_7917,N_6958,N_5395);
nand U7918 (N_7918,N_7053,N_5786);
nand U7919 (N_7919,N_5163,N_5579);
and U7920 (N_7920,N_7006,N_6093);
nor U7921 (N_7921,N_6939,N_5113);
nand U7922 (N_7922,N_6542,N_6720);
nand U7923 (N_7923,N_5410,N_6320);
or U7924 (N_7924,N_6620,N_5556);
nand U7925 (N_7925,N_5380,N_6059);
or U7926 (N_7926,N_5832,N_5774);
and U7927 (N_7927,N_6877,N_6952);
and U7928 (N_7928,N_6109,N_6897);
nor U7929 (N_7929,N_6655,N_5399);
and U7930 (N_7930,N_7192,N_5762);
nor U7931 (N_7931,N_5087,N_7389);
nand U7932 (N_7932,N_5735,N_5334);
and U7933 (N_7933,N_5432,N_6742);
nand U7934 (N_7934,N_5148,N_6689);
nor U7935 (N_7935,N_7110,N_6456);
and U7936 (N_7936,N_6327,N_6733);
or U7937 (N_7937,N_6896,N_7494);
or U7938 (N_7938,N_5562,N_7353);
nor U7939 (N_7939,N_7007,N_5140);
and U7940 (N_7940,N_6732,N_5688);
nor U7941 (N_7941,N_6152,N_5490);
and U7942 (N_7942,N_6950,N_5515);
and U7943 (N_7943,N_6682,N_5145);
and U7944 (N_7944,N_5512,N_5297);
and U7945 (N_7945,N_7441,N_5207);
nand U7946 (N_7946,N_6207,N_7203);
and U7947 (N_7947,N_6401,N_6595);
nor U7948 (N_7948,N_6984,N_6631);
and U7949 (N_7949,N_6156,N_7354);
nor U7950 (N_7950,N_7112,N_7116);
nand U7951 (N_7951,N_5770,N_6296);
or U7952 (N_7952,N_6439,N_6911);
or U7953 (N_7953,N_6853,N_7363);
and U7954 (N_7954,N_7132,N_7487);
nand U7955 (N_7955,N_6087,N_6526);
nand U7956 (N_7956,N_6308,N_6182);
nand U7957 (N_7957,N_5775,N_6311);
nor U7958 (N_7958,N_5196,N_6119);
and U7959 (N_7959,N_5984,N_7249);
nand U7960 (N_7960,N_7029,N_5282);
or U7961 (N_7961,N_6903,N_6600);
and U7962 (N_7962,N_5910,N_7373);
nand U7963 (N_7963,N_7206,N_6647);
and U7964 (N_7964,N_5573,N_5949);
nor U7965 (N_7965,N_7427,N_6673);
and U7966 (N_7966,N_5503,N_5835);
or U7967 (N_7967,N_5861,N_7289);
or U7968 (N_7968,N_5576,N_6908);
and U7969 (N_7969,N_6057,N_6558);
nor U7970 (N_7970,N_6226,N_5370);
nor U7971 (N_7971,N_6460,N_6822);
or U7972 (N_7972,N_5597,N_7421);
or U7973 (N_7973,N_6258,N_6051);
nand U7974 (N_7974,N_5313,N_5487);
or U7975 (N_7975,N_5509,N_7200);
nor U7976 (N_7976,N_6635,N_6756);
or U7977 (N_7977,N_5918,N_5226);
nand U7978 (N_7978,N_5971,N_6562);
nand U7979 (N_7979,N_5256,N_5769);
or U7980 (N_7980,N_5204,N_6806);
and U7981 (N_7981,N_6422,N_5438);
nand U7982 (N_7982,N_5848,N_5137);
nand U7983 (N_7983,N_6464,N_7256);
nand U7984 (N_7984,N_5065,N_6813);
nand U7985 (N_7985,N_5776,N_7036);
nor U7986 (N_7986,N_5237,N_5254);
nand U7987 (N_7987,N_6165,N_5603);
and U7988 (N_7988,N_6199,N_5359);
nor U7989 (N_7989,N_6298,N_5703);
and U7990 (N_7990,N_5798,N_5658);
nor U7991 (N_7991,N_7154,N_6197);
nor U7992 (N_7992,N_6597,N_6270);
nor U7993 (N_7993,N_6578,N_5281);
or U7994 (N_7994,N_5849,N_5780);
and U7995 (N_7995,N_6876,N_5659);
or U7996 (N_7996,N_5219,N_6710);
or U7997 (N_7997,N_6125,N_6760);
nand U7998 (N_7998,N_6379,N_6020);
nand U7999 (N_7999,N_5761,N_6613);
nand U8000 (N_8000,N_7218,N_6106);
nor U8001 (N_8001,N_6467,N_7075);
or U8002 (N_8002,N_5102,N_5824);
nor U8003 (N_8003,N_6638,N_5613);
nand U8004 (N_8004,N_6299,N_6472);
nor U8005 (N_8005,N_5623,N_6151);
nand U8006 (N_8006,N_5245,N_7201);
or U8007 (N_8007,N_6721,N_5566);
and U8008 (N_8008,N_6277,N_5988);
xor U8009 (N_8009,N_5729,N_6888);
or U8010 (N_8010,N_5677,N_5134);
and U8011 (N_8011,N_5208,N_7303);
or U8012 (N_8012,N_7279,N_6269);
and U8013 (N_8013,N_6394,N_5814);
nor U8014 (N_8014,N_6886,N_5142);
and U8015 (N_8015,N_5596,N_7213);
or U8016 (N_8016,N_5189,N_5247);
and U8017 (N_8017,N_7098,N_5541);
or U8018 (N_8018,N_5099,N_7422);
nand U8019 (N_8019,N_5504,N_7295);
nand U8020 (N_8020,N_7158,N_7096);
nand U8021 (N_8021,N_7170,N_7138);
nand U8022 (N_8022,N_6927,N_6584);
nor U8023 (N_8023,N_7057,N_7008);
nor U8024 (N_8024,N_5876,N_7456);
nor U8025 (N_8025,N_5695,N_5887);
nor U8026 (N_8026,N_7250,N_5151);
and U8027 (N_8027,N_7359,N_5091);
and U8028 (N_8028,N_6660,N_6589);
or U8029 (N_8029,N_7435,N_7344);
or U8030 (N_8030,N_5894,N_5362);
and U8031 (N_8031,N_5266,N_5981);
nand U8032 (N_8032,N_6808,N_5508);
or U8033 (N_8033,N_7318,N_5330);
nor U8034 (N_8034,N_6161,N_7125);
or U8035 (N_8035,N_6983,N_6944);
nand U8036 (N_8036,N_6895,N_5179);
xnor U8037 (N_8037,N_5721,N_6117);
nand U8038 (N_8038,N_5936,N_6864);
nor U8039 (N_8039,N_7089,N_5644);
and U8040 (N_8040,N_6610,N_5341);
nor U8041 (N_8041,N_7412,N_7447);
and U8042 (N_8042,N_7477,N_6499);
or U8043 (N_8043,N_5131,N_6693);
nor U8044 (N_8044,N_5257,N_5863);
nor U8045 (N_8045,N_5466,N_5869);
or U8046 (N_8046,N_5927,N_7014);
nor U8047 (N_8047,N_7131,N_5526);
and U8048 (N_8048,N_6123,N_6014);
nand U8049 (N_8049,N_6964,N_6221);
and U8050 (N_8050,N_7418,N_6443);
or U8051 (N_8051,N_7406,N_5747);
and U8052 (N_8052,N_5047,N_7380);
nor U8053 (N_8053,N_5751,N_6678);
nor U8054 (N_8054,N_7325,N_6623);
and U8055 (N_8055,N_6144,N_6544);
nor U8056 (N_8056,N_6497,N_7300);
nor U8057 (N_8057,N_7190,N_7488);
or U8058 (N_8058,N_5470,N_6263);
or U8059 (N_8059,N_6536,N_7030);
and U8060 (N_8060,N_7315,N_6085);
and U8061 (N_8061,N_5557,N_6784);
or U8062 (N_8062,N_5578,N_5295);
or U8063 (N_8063,N_6496,N_5880);
or U8064 (N_8064,N_5831,N_5188);
nand U8065 (N_8065,N_7261,N_5141);
nand U8066 (N_8066,N_7020,N_7130);
nor U8067 (N_8067,N_5215,N_7223);
xor U8068 (N_8068,N_6368,N_6466);
nor U8069 (N_8069,N_5901,N_5101);
nand U8070 (N_8070,N_7082,N_6893);
nor U8071 (N_8071,N_5639,N_7257);
nor U8072 (N_8072,N_6750,N_5590);
and U8073 (N_8073,N_7365,N_5027);
nand U8074 (N_8074,N_5244,N_6132);
nor U8075 (N_8075,N_5987,N_6240);
nand U8076 (N_8076,N_6968,N_6586);
or U8077 (N_8077,N_6185,N_5787);
nand U8078 (N_8078,N_5363,N_5727);
and U8079 (N_8079,N_7268,N_6437);
xor U8080 (N_8080,N_5685,N_5985);
and U8081 (N_8081,N_6027,N_6599);
or U8082 (N_8082,N_6141,N_5049);
or U8083 (N_8083,N_5495,N_5489);
nor U8084 (N_8084,N_5719,N_6113);
and U8085 (N_8085,N_6333,N_5280);
or U8086 (N_8086,N_5174,N_5011);
or U8087 (N_8087,N_6039,N_5897);
nand U8088 (N_8088,N_5555,N_5318);
and U8089 (N_8089,N_5018,N_7092);
or U8090 (N_8090,N_6458,N_6931);
nor U8091 (N_8091,N_5144,N_6222);
or U8092 (N_8092,N_6881,N_5592);
nor U8093 (N_8093,N_6519,N_5627);
and U8094 (N_8094,N_7140,N_6552);
nor U8095 (N_8095,N_7469,N_7386);
or U8096 (N_8096,N_5095,N_5899);
or U8097 (N_8097,N_6206,N_5090);
or U8098 (N_8098,N_6773,N_6008);
or U8099 (N_8099,N_7167,N_5227);
nand U8100 (N_8100,N_5687,N_6450);
or U8101 (N_8101,N_5035,N_6928);
nor U8102 (N_8102,N_5671,N_6629);
nor U8103 (N_8103,N_5672,N_5802);
nand U8104 (N_8104,N_7238,N_7100);
or U8105 (N_8105,N_5108,N_6446);
and U8106 (N_8106,N_7307,N_5905);
nor U8107 (N_8107,N_6243,N_7430);
xnor U8108 (N_8108,N_6169,N_5701);
nor U8109 (N_8109,N_6052,N_7087);
or U8110 (N_8110,N_5378,N_7046);
nor U8111 (N_8111,N_5081,N_6342);
nor U8112 (N_8112,N_6792,N_7146);
nor U8113 (N_8113,N_5600,N_5274);
or U8114 (N_8114,N_5892,N_5168);
or U8115 (N_8115,N_7478,N_5339);
or U8116 (N_8116,N_6230,N_7298);
or U8117 (N_8117,N_5575,N_5626);
or U8118 (N_8118,N_7202,N_5564);
nor U8119 (N_8119,N_5717,N_7407);
nand U8120 (N_8120,N_6351,N_7375);
and U8121 (N_8121,N_7475,N_6022);
or U8122 (N_8122,N_7004,N_6662);
and U8123 (N_8123,N_6513,N_6114);
nand U8124 (N_8124,N_6882,N_5069);
nor U8125 (N_8125,N_5525,N_6504);
nand U8126 (N_8126,N_7068,N_5374);
or U8127 (N_8127,N_6803,N_5485);
nand U8128 (N_8128,N_6863,N_6431);
nor U8129 (N_8129,N_5890,N_7264);
or U8130 (N_8130,N_5321,N_5094);
nor U8131 (N_8131,N_7408,N_5480);
nand U8132 (N_8132,N_5506,N_6514);
nor U8133 (N_8133,N_7160,N_6426);
and U8134 (N_8134,N_6177,N_5837);
and U8135 (N_8135,N_5271,N_5620);
and U8136 (N_8136,N_7025,N_5922);
and U8137 (N_8137,N_5114,N_7377);
or U8138 (N_8138,N_6740,N_5612);
nor U8139 (N_8139,N_5067,N_6515);
nor U8140 (N_8140,N_6925,N_7486);
nor U8141 (N_8141,N_5340,N_7334);
or U8142 (N_8142,N_6442,N_6136);
xor U8143 (N_8143,N_5911,N_5388);
nor U8144 (N_8144,N_5111,N_6421);
nand U8145 (N_8145,N_5024,N_5464);
nand U8146 (N_8146,N_6763,N_5805);
nand U8147 (N_8147,N_7493,N_5327);
and U8148 (N_8148,N_5881,N_7466);
nor U8149 (N_8149,N_6455,N_5909);
nor U8150 (N_8150,N_6400,N_5199);
nand U8151 (N_8151,N_6912,N_6420);
nor U8152 (N_8152,N_7221,N_7093);
nand U8153 (N_8153,N_6041,N_6644);
nor U8154 (N_8154,N_6076,N_6937);
nor U8155 (N_8155,N_6741,N_7450);
and U8156 (N_8156,N_5633,N_6349);
nor U8157 (N_8157,N_6071,N_5916);
nor U8158 (N_8158,N_7352,N_7081);
nor U8159 (N_8159,N_5883,N_7065);
nor U8160 (N_8160,N_5896,N_6098);
and U8161 (N_8161,N_5521,N_6804);
or U8162 (N_8162,N_6817,N_6510);
or U8163 (N_8163,N_6861,N_5968);
nor U8164 (N_8164,N_7103,N_5365);
and U8165 (N_8165,N_5917,N_5750);
or U8166 (N_8166,N_6874,N_5625);
and U8167 (N_8167,N_6989,N_6315);
and U8168 (N_8168,N_6140,N_7312);
nand U8169 (N_8169,N_5570,N_5162);
and U8170 (N_8170,N_6534,N_6066);
or U8171 (N_8171,N_7263,N_5951);
and U8172 (N_8172,N_6350,N_7376);
or U8173 (N_8173,N_5870,N_5963);
nand U8174 (N_8174,N_6477,N_7278);
nand U8175 (N_8175,N_5839,N_6862);
nand U8176 (N_8176,N_6192,N_6661);
and U8177 (N_8177,N_5150,N_5300);
and U8178 (N_8178,N_6783,N_7331);
nor U8179 (N_8179,N_6501,N_6859);
and U8180 (N_8180,N_7368,N_6444);
or U8181 (N_8181,N_6402,N_5048);
and U8182 (N_8182,N_7032,N_7244);
nand U8183 (N_8183,N_6091,N_5926);
and U8184 (N_8184,N_5286,N_6860);
nand U8185 (N_8185,N_5630,N_6362);
or U8186 (N_8186,N_5739,N_6282);
or U8187 (N_8187,N_6774,N_7364);
and U8188 (N_8188,N_7361,N_6019);
and U8189 (N_8189,N_5711,N_5548);
and U8190 (N_8190,N_5308,N_5830);
nand U8191 (N_8191,N_7191,N_6934);
nand U8192 (N_8192,N_7147,N_6628);
nor U8193 (N_8193,N_5675,N_7012);
or U8194 (N_8194,N_5491,N_7228);
and U8195 (N_8195,N_6395,N_6889);
nor U8196 (N_8196,N_6680,N_5742);
nand U8197 (N_8197,N_7151,N_6505);
and U8198 (N_8198,N_6046,N_7481);
nor U8199 (N_8199,N_6697,N_6559);
or U8200 (N_8200,N_6196,N_7274);
nor U8201 (N_8201,N_5641,N_7182);
nor U8202 (N_8202,N_5976,N_7168);
nor U8203 (N_8203,N_6672,N_7384);
nor U8204 (N_8204,N_5991,N_7156);
nor U8205 (N_8205,N_6646,N_5622);
xor U8206 (N_8206,N_5010,N_5681);
or U8207 (N_8207,N_7358,N_5986);
nor U8208 (N_8208,N_5472,N_5931);
nor U8209 (N_8209,N_6062,N_7465);
nor U8210 (N_8210,N_7180,N_7290);
and U8211 (N_8211,N_6932,N_5990);
nand U8212 (N_8212,N_7327,N_6378);
or U8213 (N_8213,N_5276,N_5859);
nor U8214 (N_8214,N_5492,N_6569);
nand U8215 (N_8215,N_5089,N_5875);
and U8216 (N_8216,N_6172,N_6344);
nand U8217 (N_8217,N_6522,N_6469);
nor U8218 (N_8218,N_6145,N_6754);
nand U8219 (N_8219,N_5594,N_7296);
nor U8220 (N_8220,N_7003,N_6982);
or U8221 (N_8221,N_5846,N_6241);
nand U8222 (N_8222,N_7241,N_7162);
nand U8223 (N_8223,N_6715,N_5384);
or U8224 (N_8224,N_7345,N_6827);
and U8225 (N_8225,N_5690,N_7335);
xnor U8226 (N_8226,N_6947,N_5232);
xnor U8227 (N_8227,N_5423,N_5212);
nand U8228 (N_8228,N_7106,N_6705);
or U8229 (N_8229,N_7141,N_5955);
or U8230 (N_8230,N_7248,N_5057);
or U8231 (N_8231,N_7193,N_7499);
nand U8232 (N_8232,N_6176,N_5587);
or U8233 (N_8233,N_6712,N_6133);
and U8234 (N_8234,N_7462,N_5601);
nor U8235 (N_8235,N_6816,N_5664);
nor U8236 (N_8236,N_7367,N_6718);
nand U8237 (N_8237,N_6706,N_5519);
or U8238 (N_8238,N_5939,N_6188);
and U8239 (N_8239,N_7383,N_5044);
nand U8240 (N_8240,N_5816,N_7009);
nand U8241 (N_8241,N_7404,N_6011);
or U8242 (N_8242,N_5942,N_7011);
and U8243 (N_8243,N_5264,N_6468);
and U8244 (N_8244,N_7099,N_5267);
nor U8245 (N_8245,N_5534,N_5407);
nand U8246 (N_8246,N_6630,N_7419);
or U8247 (N_8247,N_5864,N_6566);
nand U8248 (N_8248,N_6005,N_7282);
and U8249 (N_8249,N_5753,N_7330);
nor U8250 (N_8250,N_5059,N_5275);
xnor U8251 (N_8251,N_6839,N_5794);
nor U8252 (N_8252,N_6080,N_6273);
nor U8253 (N_8253,N_7152,N_5354);
nor U8254 (N_8254,N_6535,N_5614);
nor U8255 (N_8255,N_5610,N_6648);
nor U8256 (N_8256,N_6546,N_6695);
and U8257 (N_8257,N_5782,N_5481);
nor U8258 (N_8258,N_6987,N_5450);
nand U8259 (N_8259,N_7476,N_6517);
nor U8260 (N_8260,N_5608,N_6432);
or U8261 (N_8261,N_6995,N_6474);
nand U8262 (N_8262,N_7054,N_5152);
nand U8263 (N_8263,N_6878,N_6279);
or U8264 (N_8264,N_5900,N_5383);
nand U8265 (N_8265,N_5825,N_6900);
nor U8266 (N_8266,N_5738,N_6818);
and U8267 (N_8267,N_5319,N_6365);
and U8268 (N_8268,N_5066,N_6834);
nand U8269 (N_8269,N_5970,N_6814);
nand U8270 (N_8270,N_6541,N_7362);
or U8271 (N_8271,N_5120,N_6667);
nand U8272 (N_8272,N_5326,N_6614);
nand U8273 (N_8273,N_5983,N_6340);
or U8274 (N_8274,N_5872,N_6321);
or U8275 (N_8275,N_6842,N_6184);
nor U8276 (N_8276,N_5705,N_7056);
and U8277 (N_8277,N_6178,N_6800);
and U8278 (N_8278,N_5429,N_5652);
and U8279 (N_8279,N_5098,N_6683);
nor U8280 (N_8280,N_5352,N_6103);
xor U8281 (N_8281,N_7122,N_5913);
or U8282 (N_8282,N_5668,N_6245);
nor U8283 (N_8283,N_6419,N_6527);
and U8284 (N_8284,N_5965,N_6641);
and U8285 (N_8285,N_6181,N_7459);
nand U8286 (N_8286,N_5514,N_5707);
and U8287 (N_8287,N_5127,N_6507);
nand U8288 (N_8288,N_5486,N_6384);
and U8289 (N_8289,N_6324,N_7236);
and U8290 (N_8290,N_7471,N_7320);
nor U8291 (N_8291,N_5611,N_5844);
nand U8292 (N_8292,N_6749,N_6959);
and U8293 (N_8293,N_5430,N_6139);
nor U8294 (N_8294,N_6687,N_5930);
nor U8295 (N_8295,N_5183,N_5533);
and U8296 (N_8296,N_6227,N_6033);
nand U8297 (N_8297,N_7273,N_6010);
or U8298 (N_8298,N_6488,N_5527);
nor U8299 (N_8299,N_6685,N_6794);
and U8300 (N_8300,N_5051,N_6585);
or U8301 (N_8301,N_5518,N_7063);
or U8302 (N_8302,N_6975,N_5957);
nor U8303 (N_8303,N_6023,N_6533);
nand U8304 (N_8304,N_6015,N_5992);
nor U8305 (N_8305,N_5443,N_7439);
nor U8306 (N_8306,N_6306,N_5763);
nor U8307 (N_8307,N_5914,N_5012);
or U8308 (N_8308,N_5053,N_5635);
or U8309 (N_8309,N_5304,N_6487);
or U8310 (N_8310,N_5670,N_5125);
nor U8311 (N_8311,N_5654,N_6309);
nand U8312 (N_8312,N_5736,N_5008);
or U8313 (N_8313,N_5748,N_5542);
and U8314 (N_8314,N_5426,N_6593);
nor U8315 (N_8315,N_6448,N_5624);
nor U8316 (N_8316,N_6692,N_5698);
and U8317 (N_8317,N_7095,N_6940);
nand U8318 (N_8318,N_7097,N_7410);
and U8319 (N_8319,N_5676,N_5415);
and U8320 (N_8320,N_5417,N_5868);
nor U8321 (N_8321,N_5262,N_6846);
nand U8322 (N_8322,N_6137,N_6357);
nor U8323 (N_8323,N_6411,N_6135);
and U8324 (N_8324,N_6174,N_6722);
nor U8325 (N_8325,N_6612,N_6577);
nand U8326 (N_8326,N_6753,N_6018);
nor U8327 (N_8327,N_5975,N_5637);
and U8328 (N_8328,N_5116,N_6121);
or U8329 (N_8329,N_6302,N_5821);
or U8330 (N_8330,N_6677,N_6146);
and U8331 (N_8331,N_6923,N_5634);
nor U8332 (N_8332,N_6465,N_6173);
or U8333 (N_8333,N_5164,N_7108);
or U8334 (N_8334,N_6048,N_6772);
or U8335 (N_8335,N_5577,N_6576);
or U8336 (N_8336,N_6128,N_5186);
or U8337 (N_8337,N_6050,N_5788);
nand U8338 (N_8338,N_5412,N_5638);
nand U8339 (N_8339,N_5270,N_7023);
xnor U8340 (N_8340,N_6326,N_6289);
and U8341 (N_8341,N_6147,N_6390);
or U8342 (N_8342,N_7254,N_7197);
nand U8343 (N_8343,N_6573,N_6209);
nand U8344 (N_8344,N_7306,N_7316);
nand U8345 (N_8345,N_6213,N_6371);
nand U8346 (N_8346,N_7308,N_6430);
nor U8347 (N_8347,N_6406,N_5366);
and U8348 (N_8348,N_5891,N_7409);
nor U8349 (N_8349,N_7292,N_7438);
and U8350 (N_8350,N_6104,N_6095);
nand U8351 (N_8351,N_7079,N_6303);
xor U8352 (N_8352,N_6001,N_6024);
and U8353 (N_8353,N_6331,N_6266);
or U8354 (N_8354,N_5371,N_6000);
nor U8355 (N_8355,N_7134,N_6427);
nor U8356 (N_8356,N_5852,N_5866);
nand U8357 (N_8357,N_6988,N_6639);
and U8358 (N_8358,N_5338,N_5424);
nor U8359 (N_8359,N_7374,N_6663);
and U8360 (N_8360,N_5935,N_7416);
nor U8361 (N_8361,N_7310,N_6602);
and U8362 (N_8362,N_6478,N_5853);
or U8363 (N_8363,N_6163,N_6511);
and U8364 (N_8364,N_5337,N_6991);
and U8365 (N_8365,N_5532,N_6168);
and U8366 (N_8366,N_6288,N_6907);
and U8367 (N_8367,N_5871,N_7455);
or U8368 (N_8368,N_6571,N_6738);
nor U8369 (N_8369,N_5867,N_7251);
or U8370 (N_8370,N_6150,N_5009);
and U8371 (N_8371,N_5584,N_7222);
nor U8372 (N_8372,N_5159,N_6334);
nor U8373 (N_8373,N_5467,N_7266);
or U8374 (N_8374,N_6179,N_6910);
nor U8375 (N_8375,N_7094,N_6906);
nor U8376 (N_8376,N_6055,N_6867);
nor U8377 (N_8377,N_6899,N_5045);
and U8378 (N_8378,N_6373,N_5789);
nand U8379 (N_8379,N_7022,N_6990);
nor U8380 (N_8380,N_7405,N_6980);
or U8381 (N_8381,N_7328,N_5989);
nor U8382 (N_8382,N_5895,N_5322);
or U8383 (N_8383,N_5236,N_7392);
nand U8384 (N_8384,N_5999,N_7333);
or U8385 (N_8385,N_6054,N_7150);
nand U8386 (N_8386,N_5656,N_5648);
nand U8387 (N_8387,N_5104,N_5678);
nor U8388 (N_8388,N_7452,N_5284);
or U8389 (N_8389,N_5785,N_5553);
nand U8390 (N_8390,N_6668,N_7288);
and U8391 (N_8391,N_7171,N_6244);
nand U8392 (N_8392,N_6901,N_5933);
nor U8393 (N_8393,N_6229,N_7039);
nor U8394 (N_8394,N_5252,N_6089);
or U8395 (N_8395,N_6170,N_5494);
or U8396 (N_8396,N_5444,N_5807);
nand U8397 (N_8397,N_5462,N_7169);
or U8398 (N_8398,N_5497,N_5855);
nand U8399 (N_8399,N_5885,N_5206);
and U8400 (N_8400,N_7314,N_6919);
and U8401 (N_8401,N_7072,N_6100);
and U8402 (N_8402,N_5202,N_5414);
and U8403 (N_8403,N_5192,N_6699);
or U8404 (N_8404,N_5944,N_6840);
or U8405 (N_8405,N_5158,N_5015);
nand U8406 (N_8406,N_6986,N_5812);
and U8407 (N_8407,N_5249,N_6553);
and U8408 (N_8408,N_5033,N_6714);
or U8409 (N_8409,N_5547,N_6102);
or U8410 (N_8410,N_5709,N_6116);
or U8411 (N_8411,N_5182,N_5505);
nand U8412 (N_8412,N_7215,N_7483);
nor U8413 (N_8413,N_6276,N_6650);
nor U8414 (N_8414,N_5997,N_6265);
and U8415 (N_8415,N_6126,N_5758);
nand U8416 (N_8416,N_5743,N_6622);
nand U8417 (N_8417,N_6232,N_5843);
or U8418 (N_8418,N_7027,N_5096);
and U8419 (N_8419,N_7148,N_6183);
nor U8420 (N_8420,N_5589,N_5389);
nand U8421 (N_8421,N_6030,N_7153);
nor U8422 (N_8422,N_7231,N_6214);
or U8423 (N_8423,N_7324,N_6254);
nor U8424 (N_8424,N_6154,N_5879);
and U8425 (N_8425,N_6615,N_5465);
and U8426 (N_8426,N_5862,N_6217);
nor U8427 (N_8427,N_5445,N_5724);
or U8428 (N_8428,N_5934,N_7041);
or U8429 (N_8429,N_6219,N_5258);
nand U8430 (N_8430,N_6955,N_5356);
and U8431 (N_8431,N_6462,N_5502);
and U8432 (N_8432,N_5615,N_5714);
nand U8433 (N_8433,N_5128,N_7317);
and U8434 (N_8434,N_6377,N_7379);
or U8435 (N_8435,N_6086,N_5285);
nor U8436 (N_8436,N_5020,N_5169);
nor U8437 (N_8437,N_7176,N_5026);
and U8438 (N_8438,N_6021,N_5842);
nand U8439 (N_8439,N_5377,N_6616);
nor U8440 (N_8440,N_5223,N_5343);
nor U8441 (N_8441,N_7393,N_6414);
nand U8442 (N_8442,N_7240,N_6107);
and U8443 (N_8443,N_5138,N_6294);
xor U8444 (N_8444,N_5200,N_5568);
or U8445 (N_8445,N_6681,N_6904);
nor U8446 (N_8446,N_6587,N_6713);
or U8447 (N_8447,N_6969,N_7482);
or U8448 (N_8448,N_6961,N_6645);
nor U8449 (N_8449,N_5235,N_7340);
nor U8450 (N_8450,N_5535,N_7414);
nor U8451 (N_8451,N_6974,N_6723);
and U8452 (N_8452,N_5582,N_5220);
or U8453 (N_8453,N_6441,N_5954);
and U8454 (N_8454,N_5741,N_6601);
or U8455 (N_8455,N_5599,N_6547);
and U8456 (N_8456,N_6805,N_5689);
nand U8457 (N_8457,N_5791,N_5559);
nor U8458 (N_8458,N_6300,N_6929);
nor U8459 (N_8459,N_5058,N_6486);
and U8460 (N_8460,N_6898,N_5084);
or U8461 (N_8461,N_7491,N_6654);
nand U8462 (N_8462,N_6393,N_5993);
or U8463 (N_8463,N_6508,N_7281);
or U8464 (N_8464,N_7473,N_6985);
or U8465 (N_8465,N_7437,N_6201);
or U8466 (N_8466,N_5082,N_5043);
nor U8467 (N_8467,N_5361,N_6892);
and U8468 (N_8468,N_6212,N_6746);
or U8469 (N_8469,N_5146,N_7194);
nand U8470 (N_8470,N_6028,N_6410);
nor U8471 (N_8471,N_5401,N_6345);
nor U8472 (N_8472,N_6981,N_6954);
or U8473 (N_8473,N_5646,N_5962);
and U8474 (N_8474,N_6256,N_5221);
nor U8475 (N_8475,N_6865,N_5070);
nor U8476 (N_8476,N_6870,N_6238);
and U8477 (N_8477,N_5536,N_7426);
and U8478 (N_8478,N_6999,N_5977);
or U8479 (N_8479,N_6696,N_7059);
nor U8480 (N_8480,N_6626,N_7024);
and U8481 (N_8481,N_5325,N_5004);
and U8482 (N_8482,N_5411,N_7417);
nor U8483 (N_8483,N_5292,N_6703);
or U8484 (N_8484,N_6092,N_6281);
and U8485 (N_8485,N_5193,N_7049);
and U8486 (N_8486,N_5106,N_6364);
and U8487 (N_8487,N_7433,N_6837);
or U8488 (N_8488,N_6412,N_6417);
or U8489 (N_8489,N_6854,N_6637);
and U8490 (N_8490,N_5517,N_5754);
nor U8491 (N_8491,N_7495,N_6484);
or U8492 (N_8492,N_5980,N_6006);
nor U8493 (N_8493,N_5259,N_7172);
nor U8494 (N_8494,N_5211,N_7411);
nor U8495 (N_8495,N_6871,N_5068);
nor U8496 (N_8496,N_6363,N_5468);
and U8497 (N_8497,N_5565,N_6567);
nor U8498 (N_8498,N_6717,N_5921);
nand U8499 (N_8499,N_5165,N_7350);
nand U8500 (N_8500,N_5874,N_5631);
or U8501 (N_8501,N_7394,N_6736);
nand U8502 (N_8502,N_5097,N_6926);
nand U8503 (N_8503,N_5906,N_7423);
nand U8504 (N_8504,N_7497,N_6843);
and U8505 (N_8505,N_7069,N_5425);
and U8506 (N_8506,N_6352,N_5387);
xnor U8507 (N_8507,N_6686,N_5771);
nor U8508 (N_8508,N_5593,N_6633);
nand U8509 (N_8509,N_6596,N_6210);
xnor U8510 (N_8510,N_5103,N_5628);
or U8511 (N_8511,N_7066,N_6657);
and U8512 (N_8512,N_6791,N_6830);
and U8513 (N_8513,N_7233,N_6122);
and U8514 (N_8514,N_5537,N_6475);
nor U8515 (N_8515,N_5708,N_6193);
nand U8516 (N_8516,N_7002,N_6204);
and U8517 (N_8517,N_5712,N_7342);
nand U8518 (N_8518,N_5799,N_7453);
nand U8519 (N_8519,N_7177,N_6869);
xor U8520 (N_8520,N_6920,N_5956);
or U8521 (N_8521,N_5734,N_7302);
nor U8522 (N_8522,N_7323,N_5666);
and U8523 (N_8523,N_6036,N_5348);
or U8524 (N_8524,N_5482,N_6084);
nand U8525 (N_8525,N_6781,N_7051);
and U8526 (N_8526,N_5682,N_6875);
or U8527 (N_8527,N_5817,N_6775);
and U8528 (N_8528,N_6938,N_7341);
and U8529 (N_8529,N_6554,N_5213);
nand U8530 (N_8530,N_6797,N_7000);
or U8531 (N_8531,N_5498,N_6728);
nand U8532 (N_8532,N_7243,N_6305);
and U8533 (N_8533,N_5733,N_5583);
nor U8534 (N_8534,N_6453,N_6551);
nor U8535 (N_8535,N_6966,N_5728);
and U8536 (N_8536,N_5878,N_6012);
nor U8537 (N_8537,N_5448,N_5195);
nor U8538 (N_8538,N_5073,N_5595);
nor U8539 (N_8539,N_5833,N_6043);
nand U8540 (N_8540,N_5773,N_5889);
and U8541 (N_8541,N_5447,N_7209);
nor U8542 (N_8542,N_5496,N_6494);
nand U8543 (N_8543,N_7178,N_6833);
or U8544 (N_8544,N_5510,N_5928);
or U8545 (N_8545,N_5815,N_5645);
nor U8546 (N_8546,N_5161,N_6454);
or U8547 (N_8547,N_6074,N_6716);
nand U8548 (N_8548,N_6777,N_5667);
xor U8549 (N_8549,N_6570,N_6312);
nor U8550 (N_8550,N_6476,N_6260);
nor U8551 (N_8551,N_5075,N_6574);
and U8552 (N_8552,N_6609,N_5224);
nand U8553 (N_8553,N_5737,N_6565);
and U8554 (N_8554,N_7062,N_6158);
nor U8555 (N_8555,N_6407,N_6820);
or U8556 (N_8556,N_6708,N_6731);
nor U8557 (N_8557,N_7451,N_5203);
and U8558 (N_8558,N_6129,N_6856);
nand U8559 (N_8559,N_7431,N_6619);
nand U8560 (N_8560,N_6413,N_6381);
and U8561 (N_8561,N_5316,N_5474);
or U8562 (N_8562,N_7214,N_6108);
nand U8563 (N_8563,N_7114,N_6557);
and U8564 (N_8564,N_6249,N_5243);
nand U8565 (N_8565,N_6992,N_7287);
nor U8566 (N_8566,N_5307,N_6482);
nor U8567 (N_8567,N_5529,N_5393);
or U8568 (N_8568,N_6118,N_5857);
or U8569 (N_8569,N_5037,N_6332);
nor U8570 (N_8570,N_7128,N_5229);
and U8571 (N_8571,N_5618,N_5972);
and U8572 (N_8572,N_5122,N_7381);
nor U8573 (N_8573,N_7460,N_5925);
nand U8574 (N_8574,N_6356,N_6745);
nand U8575 (N_8575,N_7434,N_7161);
nor U8576 (N_8576,N_5157,N_5663);
and U8577 (N_8577,N_7356,N_5516);
and U8578 (N_8578,N_5882,N_6852);
nor U8579 (N_8579,N_5178,N_7461);
and U8580 (N_8580,N_6640,N_6360);
nand U8581 (N_8581,N_5475,N_5017);
nor U8582 (N_8582,N_5381,N_6764);
or U8583 (N_8583,N_6537,N_6735);
or U8584 (N_8584,N_6605,N_6246);
nand U8585 (N_8585,N_5088,N_7401);
or U8586 (N_8586,N_7145,N_5302);
nand U8587 (N_8587,N_5328,N_6047);
or U8588 (N_8588,N_6016,N_6403);
or U8589 (N_8589,N_7390,N_6973);
xor U8590 (N_8590,N_6445,N_7033);
or U8591 (N_8591,N_6771,N_5718);
nand U8592 (N_8592,N_6425,N_6250);
and U8593 (N_8593,N_6993,N_5793);
nor U8594 (N_8594,N_6463,N_7305);
or U8595 (N_8595,N_6336,N_5136);
nand U8596 (N_8596,N_5607,N_5439);
nand U8597 (N_8597,N_7187,N_6295);
or U8598 (N_8598,N_7127,N_6786);
and U8599 (N_8599,N_6948,N_5795);
nand U8600 (N_8600,N_7225,N_5586);
or U8601 (N_8601,N_6211,N_6752);
nor U8602 (N_8602,N_6166,N_5767);
and U8603 (N_8603,N_5469,N_6025);
or U8604 (N_8604,N_5796,N_6953);
and U8605 (N_8605,N_6521,N_6101);
or U8606 (N_8606,N_5838,N_6367);
nor U8607 (N_8607,N_5725,N_6849);
nor U8608 (N_8608,N_5115,N_6621);
or U8609 (N_8609,N_5801,N_6607);
or U8610 (N_8610,N_6594,N_6164);
and U8611 (N_8611,N_6424,N_7403);
and U8612 (N_8612,N_7454,N_5912);
nand U8613 (N_8613,N_6297,N_5669);
nor U8614 (N_8614,N_6386,N_5940);
nand U8615 (N_8615,N_6252,N_7388);
and U8616 (N_8616,N_6762,N_5581);
or U8617 (N_8617,N_7013,N_5173);
nand U8618 (N_8618,N_6205,N_7395);
or U8619 (N_8619,N_5194,N_7211);
or U8620 (N_8620,N_5500,N_6858);
nand U8621 (N_8621,N_6700,N_6757);
nor U8622 (N_8622,N_6575,N_6675);
and U8623 (N_8623,N_5408,N_6809);
or U8624 (N_8624,N_5463,N_7492);
nand U8625 (N_8625,N_5779,N_7078);
and U8626 (N_8626,N_6729,N_6642);
nor U8627 (N_8627,N_6216,N_5315);
nand U8628 (N_8628,N_5446,N_5632);
nor U8629 (N_8629,N_5390,N_6237);
nand U8630 (N_8630,N_5764,N_5324);
nor U8631 (N_8631,N_5287,N_6157);
nand U8632 (N_8632,N_5349,N_7208);
or U8633 (N_8633,N_5451,N_6879);
nor U8634 (N_8634,N_7479,N_5657);
nor U8635 (N_8635,N_7185,N_5002);
nand U8636 (N_8636,N_6598,N_5520);
nand U8637 (N_8637,N_7343,N_6218);
and U8638 (N_8638,N_5025,N_6261);
or U8639 (N_8639,N_5860,N_5023);
nor U8640 (N_8640,N_5886,N_7322);
or U8641 (N_8641,N_7018,N_7259);
nand U8642 (N_8642,N_6038,N_6704);
or U8643 (N_8643,N_7442,N_6049);
nor U8644 (N_8644,N_6355,N_5920);
nor U8645 (N_8645,N_7084,N_6257);
nor U8646 (N_8646,N_6528,N_6690);
nand U8647 (N_8647,N_7237,N_5684);
nor U8648 (N_8648,N_5060,N_7449);
nor U8649 (N_8649,N_6498,N_7349);
nand U8650 (N_8650,N_6292,N_5679);
nor U8651 (N_8651,N_6824,N_5031);
nand U8652 (N_8652,N_5574,N_6523);
nor U8653 (N_8653,N_6766,N_7107);
nand U8654 (N_8654,N_5034,N_5086);
or U8655 (N_8655,N_7126,N_6160);
and U8656 (N_8656,N_6013,N_6525);
nor U8657 (N_8657,N_7269,N_6737);
nor U8658 (N_8658,N_5745,N_5100);
or U8659 (N_8659,N_6579,N_5823);
and U8660 (N_8660,N_5765,N_7120);
nor U8661 (N_8661,N_5283,N_7470);
nand U8662 (N_8662,N_5609,N_6819);
and U8663 (N_8663,N_5016,N_6857);
nor U8664 (N_8664,N_5032,N_6130);
and U8665 (N_8665,N_7489,N_5797);
or U8666 (N_8666,N_5919,N_5269);
nand U8667 (N_8667,N_6883,N_7457);
xor U8668 (N_8668,N_5650,N_5149);
nor U8669 (N_8669,N_6316,N_6347);
nand U8670 (N_8670,N_7005,N_5398);
or U8671 (N_8671,N_6838,N_5740);
nand U8672 (N_8672,N_6823,N_6835);
and U8673 (N_8673,N_6361,N_6031);
xor U8674 (N_8674,N_7073,N_5953);
and U8675 (N_8675,N_6385,N_5376);
and U8676 (N_8676,N_5943,N_6399);
nor U8677 (N_8677,N_6936,N_5246);
or U8678 (N_8678,N_5210,N_5950);
and U8679 (N_8679,N_5759,N_7420);
nand U8680 (N_8680,N_6073,N_5847);
and U8681 (N_8681,N_6503,N_7468);
or U8682 (N_8682,N_6855,N_5409);
nand U8683 (N_8683,N_6035,N_6956);
nor U8684 (N_8684,N_7260,N_6099);
or U8685 (N_8685,N_5028,N_5752);
nor U8686 (N_8686,N_5135,N_6915);
and U8687 (N_8687,N_5946,N_6965);
nand U8688 (N_8688,N_6034,N_5436);
or U8689 (N_8689,N_6435,N_6053);
nand U8690 (N_8690,N_5778,N_5619);
nand U8691 (N_8691,N_5888,N_7199);
nand U8692 (N_8692,N_5198,N_6383);
nor U8693 (N_8693,N_7188,N_5558);
and U8694 (N_8694,N_6531,N_5197);
nor U8695 (N_8695,N_5177,N_6624);
nand U8696 (N_8696,N_6759,N_6776);
nand U8697 (N_8697,N_6317,N_7396);
and U8698 (N_8698,N_5184,N_5982);
or U8699 (N_8699,N_5937,N_5781);
and U8700 (N_8700,N_5126,N_5530);
and U8701 (N_8701,N_5452,N_5007);
or U8702 (N_8702,N_5673,N_6933);
and U8703 (N_8703,N_5143,N_5345);
xnor U8704 (N_8704,N_7181,N_6142);
nor U8705 (N_8705,N_6821,N_6090);
nand U8706 (N_8706,N_6343,N_7372);
nor U8707 (N_8707,N_7258,N_5820);
nor U8708 (N_8708,N_7186,N_6545);
or U8709 (N_8709,N_7015,N_6770);
or U8710 (N_8710,N_6285,N_5317);
xnor U8711 (N_8711,N_7304,N_7285);
and U8712 (N_8712,N_5121,N_6405);
or U8713 (N_8713,N_5661,N_7157);
or U8714 (N_8714,N_7090,N_5746);
nand U8715 (N_8715,N_5030,N_6228);
or U8716 (N_8716,N_5129,N_7113);
and U8717 (N_8717,N_5309,N_6389);
or U8718 (N_8718,N_5217,N_5288);
and U8719 (N_8719,N_6267,N_5845);
nor U8720 (N_8720,N_5629,N_5299);
xor U8721 (N_8721,N_5139,N_7091);
and U8722 (N_8722,N_5306,N_5038);
nand U8723 (N_8723,N_5572,N_5449);
nand U8724 (N_8724,N_5777,N_5723);
nor U8725 (N_8725,N_7267,N_5311);
nor U8726 (N_8726,N_5493,N_5155);
nor U8727 (N_8727,N_5172,N_6339);
or U8728 (N_8728,N_7115,N_6436);
and U8729 (N_8729,N_7319,N_6314);
nand U8730 (N_8730,N_6894,N_6564);
nor U8731 (N_8731,N_5836,N_5329);
and U8732 (N_8732,N_7387,N_6060);
or U8733 (N_8733,N_5357,N_5588);
nand U8734 (N_8734,N_7227,N_7210);
and U8735 (N_8735,N_6769,N_5811);
nor U8736 (N_8736,N_5369,N_6782);
nand U8737 (N_8737,N_7445,N_7313);
xnor U8738 (N_8738,N_6323,N_5961);
or U8739 (N_8739,N_5973,N_7293);
and U8740 (N_8740,N_7135,N_7165);
nand U8741 (N_8741,N_6611,N_6943);
and U8742 (N_8742,N_5233,N_6359);
nand U8743 (N_8743,N_6796,N_5715);
nor U8744 (N_8744,N_7001,N_5732);
nand U8745 (N_8745,N_5706,N_5544);
and U8746 (N_8746,N_6807,N_7351);
or U8747 (N_8747,N_6081,N_6159);
nand U8748 (N_8748,N_6078,N_5290);
nor U8749 (N_8749,N_5042,N_7413);
and U8750 (N_8750,N_6785,N_6385);
nand U8751 (N_8751,N_6525,N_6140);
nand U8752 (N_8752,N_7196,N_5819);
and U8753 (N_8753,N_7008,N_6141);
or U8754 (N_8754,N_7440,N_6405);
nand U8755 (N_8755,N_5130,N_6682);
nor U8756 (N_8756,N_6089,N_6857);
nor U8757 (N_8757,N_5885,N_5797);
nand U8758 (N_8758,N_6658,N_6679);
nand U8759 (N_8759,N_6251,N_5002);
nor U8760 (N_8760,N_7446,N_6724);
or U8761 (N_8761,N_5709,N_7217);
and U8762 (N_8762,N_6249,N_5460);
nor U8763 (N_8763,N_6296,N_6183);
nor U8764 (N_8764,N_5377,N_6546);
and U8765 (N_8765,N_5570,N_5179);
nor U8766 (N_8766,N_5302,N_6684);
nand U8767 (N_8767,N_5682,N_7214);
or U8768 (N_8768,N_6966,N_6654);
or U8769 (N_8769,N_6581,N_5558);
nor U8770 (N_8770,N_5583,N_6433);
and U8771 (N_8771,N_5355,N_5685);
and U8772 (N_8772,N_5188,N_7383);
nand U8773 (N_8773,N_5762,N_5884);
xnor U8774 (N_8774,N_6440,N_6433);
nand U8775 (N_8775,N_5785,N_5450);
nand U8776 (N_8776,N_5567,N_6795);
and U8777 (N_8777,N_6001,N_5317);
nand U8778 (N_8778,N_5493,N_6855);
nor U8779 (N_8779,N_5045,N_6159);
nand U8780 (N_8780,N_5403,N_6339);
nor U8781 (N_8781,N_6083,N_7213);
nand U8782 (N_8782,N_5710,N_6859);
nand U8783 (N_8783,N_7490,N_6700);
nor U8784 (N_8784,N_5306,N_6367);
and U8785 (N_8785,N_7094,N_6136);
nand U8786 (N_8786,N_6300,N_6004);
or U8787 (N_8787,N_5729,N_5083);
xor U8788 (N_8788,N_6742,N_5196);
nor U8789 (N_8789,N_6700,N_7208);
xor U8790 (N_8790,N_6627,N_5153);
nor U8791 (N_8791,N_7498,N_6041);
nand U8792 (N_8792,N_6279,N_5758);
nand U8793 (N_8793,N_6321,N_6593);
xor U8794 (N_8794,N_5512,N_6145);
or U8795 (N_8795,N_6180,N_7281);
and U8796 (N_8796,N_6850,N_7172);
or U8797 (N_8797,N_7280,N_7486);
or U8798 (N_8798,N_6627,N_7486);
and U8799 (N_8799,N_5128,N_5337);
or U8800 (N_8800,N_5511,N_6573);
or U8801 (N_8801,N_6499,N_5064);
xor U8802 (N_8802,N_5381,N_5550);
and U8803 (N_8803,N_6083,N_5849);
nor U8804 (N_8804,N_7413,N_5260);
and U8805 (N_8805,N_5020,N_6106);
and U8806 (N_8806,N_5915,N_6685);
nor U8807 (N_8807,N_6739,N_6460);
and U8808 (N_8808,N_6572,N_6801);
nand U8809 (N_8809,N_5878,N_5670);
nor U8810 (N_8810,N_7323,N_6491);
or U8811 (N_8811,N_7237,N_6351);
nand U8812 (N_8812,N_6024,N_7386);
nor U8813 (N_8813,N_6841,N_5522);
nand U8814 (N_8814,N_6373,N_6358);
or U8815 (N_8815,N_6352,N_7199);
or U8816 (N_8816,N_5520,N_6522);
nand U8817 (N_8817,N_7399,N_6412);
nor U8818 (N_8818,N_7191,N_7424);
xnor U8819 (N_8819,N_6646,N_5109);
nor U8820 (N_8820,N_6694,N_5190);
nand U8821 (N_8821,N_5428,N_6396);
nand U8822 (N_8822,N_5621,N_6325);
nand U8823 (N_8823,N_7278,N_6293);
or U8824 (N_8824,N_5385,N_7260);
and U8825 (N_8825,N_7230,N_7051);
nor U8826 (N_8826,N_5760,N_5776);
nor U8827 (N_8827,N_6270,N_7382);
nand U8828 (N_8828,N_6945,N_6960);
nor U8829 (N_8829,N_5732,N_5972);
xor U8830 (N_8830,N_5644,N_7306);
or U8831 (N_8831,N_5853,N_6307);
and U8832 (N_8832,N_7201,N_6742);
and U8833 (N_8833,N_5224,N_7303);
nand U8834 (N_8834,N_5185,N_7490);
or U8835 (N_8835,N_6970,N_6955);
nand U8836 (N_8836,N_5549,N_6625);
or U8837 (N_8837,N_6816,N_5119);
nor U8838 (N_8838,N_5530,N_5304);
nor U8839 (N_8839,N_5184,N_6303);
or U8840 (N_8840,N_6240,N_7472);
or U8841 (N_8841,N_5597,N_5909);
and U8842 (N_8842,N_7255,N_5327);
nor U8843 (N_8843,N_6750,N_5584);
or U8844 (N_8844,N_6629,N_5804);
and U8845 (N_8845,N_7148,N_5043);
nor U8846 (N_8846,N_5276,N_7483);
and U8847 (N_8847,N_6457,N_7126);
and U8848 (N_8848,N_5415,N_6907);
nand U8849 (N_8849,N_6031,N_6727);
and U8850 (N_8850,N_5972,N_5843);
nor U8851 (N_8851,N_5857,N_6977);
and U8852 (N_8852,N_6445,N_6264);
nand U8853 (N_8853,N_6548,N_6417);
nor U8854 (N_8854,N_5617,N_7242);
or U8855 (N_8855,N_6152,N_5045);
and U8856 (N_8856,N_6882,N_5382);
nor U8857 (N_8857,N_5331,N_5474);
nor U8858 (N_8858,N_6814,N_5935);
nor U8859 (N_8859,N_6683,N_5084);
and U8860 (N_8860,N_7208,N_5756);
or U8861 (N_8861,N_6067,N_5729);
and U8862 (N_8862,N_5881,N_5156);
nor U8863 (N_8863,N_5989,N_5371);
nand U8864 (N_8864,N_7111,N_6591);
and U8865 (N_8865,N_7083,N_6447);
and U8866 (N_8866,N_6192,N_6325);
or U8867 (N_8867,N_5152,N_6419);
nor U8868 (N_8868,N_6093,N_6400);
or U8869 (N_8869,N_7020,N_7450);
nor U8870 (N_8870,N_6289,N_6637);
or U8871 (N_8871,N_7193,N_7164);
nand U8872 (N_8872,N_6723,N_5068);
or U8873 (N_8873,N_5728,N_7164);
nor U8874 (N_8874,N_6233,N_5642);
or U8875 (N_8875,N_6677,N_5844);
nor U8876 (N_8876,N_7499,N_5039);
and U8877 (N_8877,N_5788,N_5076);
and U8878 (N_8878,N_7269,N_6844);
xnor U8879 (N_8879,N_6617,N_5297);
nor U8880 (N_8880,N_7094,N_7271);
and U8881 (N_8881,N_6027,N_6537);
and U8882 (N_8882,N_5250,N_7297);
nand U8883 (N_8883,N_5377,N_5654);
nand U8884 (N_8884,N_5920,N_7008);
nor U8885 (N_8885,N_6472,N_6150);
and U8886 (N_8886,N_5832,N_6355);
and U8887 (N_8887,N_5209,N_5255);
nor U8888 (N_8888,N_7375,N_5907);
and U8889 (N_8889,N_6366,N_5007);
nor U8890 (N_8890,N_7145,N_7368);
or U8891 (N_8891,N_5023,N_6181);
nand U8892 (N_8892,N_6430,N_6191);
nand U8893 (N_8893,N_5174,N_7066);
nor U8894 (N_8894,N_5776,N_6420);
nor U8895 (N_8895,N_5406,N_7234);
nand U8896 (N_8896,N_7074,N_6823);
nand U8897 (N_8897,N_5799,N_6617);
or U8898 (N_8898,N_6010,N_6949);
nor U8899 (N_8899,N_5612,N_6560);
and U8900 (N_8900,N_6458,N_6314);
and U8901 (N_8901,N_7305,N_5386);
or U8902 (N_8902,N_5249,N_5975);
nor U8903 (N_8903,N_6804,N_5166);
and U8904 (N_8904,N_5951,N_7234);
and U8905 (N_8905,N_6827,N_5640);
or U8906 (N_8906,N_5730,N_5297);
or U8907 (N_8907,N_6839,N_7303);
or U8908 (N_8908,N_5520,N_7254);
and U8909 (N_8909,N_5870,N_6465);
nand U8910 (N_8910,N_6921,N_5789);
nand U8911 (N_8911,N_6235,N_5719);
and U8912 (N_8912,N_6741,N_6392);
and U8913 (N_8913,N_6091,N_7357);
and U8914 (N_8914,N_6117,N_6650);
and U8915 (N_8915,N_5533,N_7440);
nand U8916 (N_8916,N_7173,N_6083);
or U8917 (N_8917,N_5360,N_7450);
or U8918 (N_8918,N_6721,N_6747);
nand U8919 (N_8919,N_5059,N_6270);
and U8920 (N_8920,N_7207,N_6650);
nor U8921 (N_8921,N_5453,N_7312);
nor U8922 (N_8922,N_6404,N_5688);
or U8923 (N_8923,N_5544,N_6620);
and U8924 (N_8924,N_7109,N_5697);
or U8925 (N_8925,N_5655,N_7328);
or U8926 (N_8926,N_6247,N_6781);
nor U8927 (N_8927,N_6496,N_6475);
nor U8928 (N_8928,N_5419,N_6900);
nor U8929 (N_8929,N_6510,N_5353);
nor U8930 (N_8930,N_7113,N_5194);
nor U8931 (N_8931,N_7134,N_7145);
nor U8932 (N_8932,N_5115,N_5281);
or U8933 (N_8933,N_7217,N_6562);
xnor U8934 (N_8934,N_5977,N_5204);
nor U8935 (N_8935,N_5150,N_6421);
and U8936 (N_8936,N_6187,N_6570);
nor U8937 (N_8937,N_6871,N_5623);
xor U8938 (N_8938,N_6743,N_5965);
or U8939 (N_8939,N_5095,N_5804);
nand U8940 (N_8940,N_5937,N_6024);
nor U8941 (N_8941,N_7071,N_6437);
nand U8942 (N_8942,N_6978,N_6710);
and U8943 (N_8943,N_7476,N_5419);
nand U8944 (N_8944,N_7040,N_6152);
or U8945 (N_8945,N_5999,N_6366);
or U8946 (N_8946,N_6439,N_6681);
nand U8947 (N_8947,N_6753,N_7046);
and U8948 (N_8948,N_5887,N_7367);
nand U8949 (N_8949,N_5521,N_5689);
and U8950 (N_8950,N_6536,N_7150);
nand U8951 (N_8951,N_5346,N_7010);
nor U8952 (N_8952,N_6191,N_6442);
nor U8953 (N_8953,N_5053,N_6635);
and U8954 (N_8954,N_6505,N_7091);
or U8955 (N_8955,N_6725,N_5181);
nor U8956 (N_8956,N_5182,N_6500);
nor U8957 (N_8957,N_7017,N_6381);
and U8958 (N_8958,N_5513,N_7331);
and U8959 (N_8959,N_6577,N_6007);
nor U8960 (N_8960,N_5523,N_5476);
and U8961 (N_8961,N_5345,N_6469);
and U8962 (N_8962,N_6287,N_6158);
or U8963 (N_8963,N_5482,N_6583);
or U8964 (N_8964,N_5318,N_5733);
and U8965 (N_8965,N_6802,N_6696);
nand U8966 (N_8966,N_7355,N_6217);
or U8967 (N_8967,N_5083,N_5932);
nor U8968 (N_8968,N_5129,N_6823);
or U8969 (N_8969,N_6540,N_5737);
nand U8970 (N_8970,N_6094,N_6702);
or U8971 (N_8971,N_7216,N_6167);
or U8972 (N_8972,N_7128,N_7302);
nor U8973 (N_8973,N_6599,N_6232);
nand U8974 (N_8974,N_7005,N_5121);
and U8975 (N_8975,N_6428,N_5149);
and U8976 (N_8976,N_7245,N_5847);
nand U8977 (N_8977,N_7353,N_5269);
and U8978 (N_8978,N_6334,N_6267);
nand U8979 (N_8979,N_6873,N_5504);
nand U8980 (N_8980,N_5379,N_6622);
and U8981 (N_8981,N_6399,N_7312);
or U8982 (N_8982,N_5254,N_6524);
nand U8983 (N_8983,N_5682,N_5476);
nor U8984 (N_8984,N_7212,N_7063);
nand U8985 (N_8985,N_5274,N_6229);
or U8986 (N_8986,N_6430,N_5000);
nor U8987 (N_8987,N_5736,N_6665);
and U8988 (N_8988,N_5828,N_5360);
nor U8989 (N_8989,N_5437,N_6447);
nor U8990 (N_8990,N_6644,N_6086);
nand U8991 (N_8991,N_6046,N_5050);
nor U8992 (N_8992,N_5268,N_6906);
nor U8993 (N_8993,N_7259,N_7016);
nand U8994 (N_8994,N_6328,N_5014);
or U8995 (N_8995,N_6171,N_7058);
nand U8996 (N_8996,N_6849,N_6303);
nand U8997 (N_8997,N_6286,N_5394);
xor U8998 (N_8998,N_6951,N_6670);
nor U8999 (N_8999,N_7248,N_5219);
or U9000 (N_9000,N_7022,N_5473);
and U9001 (N_9001,N_6472,N_5321);
and U9002 (N_9002,N_5099,N_7486);
or U9003 (N_9003,N_5632,N_7366);
nand U9004 (N_9004,N_5167,N_6851);
nand U9005 (N_9005,N_6407,N_5750);
and U9006 (N_9006,N_5896,N_5808);
nand U9007 (N_9007,N_6417,N_6757);
nor U9008 (N_9008,N_6008,N_5826);
and U9009 (N_9009,N_6531,N_5187);
and U9010 (N_9010,N_6027,N_6181);
nor U9011 (N_9011,N_5592,N_6453);
or U9012 (N_9012,N_6526,N_5004);
nor U9013 (N_9013,N_5598,N_5066);
nand U9014 (N_9014,N_5661,N_5547);
or U9015 (N_9015,N_5999,N_6682);
nor U9016 (N_9016,N_6905,N_6312);
and U9017 (N_9017,N_5960,N_6050);
nand U9018 (N_9018,N_6476,N_5043);
nand U9019 (N_9019,N_5098,N_6582);
and U9020 (N_9020,N_5064,N_6046);
nand U9021 (N_9021,N_6625,N_6168);
and U9022 (N_9022,N_6942,N_6658);
and U9023 (N_9023,N_6257,N_5461);
nand U9024 (N_9024,N_5523,N_5120);
nor U9025 (N_9025,N_5307,N_6718);
xor U9026 (N_9026,N_6038,N_6360);
nand U9027 (N_9027,N_5605,N_5495);
nor U9028 (N_9028,N_5087,N_6365);
and U9029 (N_9029,N_6039,N_7060);
nand U9030 (N_9030,N_6161,N_5876);
and U9031 (N_9031,N_7354,N_5311);
xor U9032 (N_9032,N_5663,N_5414);
and U9033 (N_9033,N_6815,N_6969);
or U9034 (N_9034,N_5275,N_7476);
nor U9035 (N_9035,N_6971,N_6816);
nand U9036 (N_9036,N_5539,N_7367);
xnor U9037 (N_9037,N_6878,N_7431);
or U9038 (N_9038,N_5783,N_5913);
or U9039 (N_9039,N_6079,N_6316);
and U9040 (N_9040,N_6430,N_6937);
and U9041 (N_9041,N_7227,N_6783);
xor U9042 (N_9042,N_7231,N_5319);
and U9043 (N_9043,N_6944,N_7285);
or U9044 (N_9044,N_7068,N_6806);
or U9045 (N_9045,N_6512,N_6599);
and U9046 (N_9046,N_6122,N_6890);
nor U9047 (N_9047,N_5495,N_5164);
nand U9048 (N_9048,N_5069,N_7380);
or U9049 (N_9049,N_6296,N_7140);
nand U9050 (N_9050,N_5126,N_6449);
or U9051 (N_9051,N_5724,N_5053);
nand U9052 (N_9052,N_5227,N_6358);
and U9053 (N_9053,N_6691,N_6654);
or U9054 (N_9054,N_6756,N_7400);
nand U9055 (N_9055,N_6211,N_5856);
nor U9056 (N_9056,N_7135,N_7179);
or U9057 (N_9057,N_5934,N_6576);
nor U9058 (N_9058,N_5726,N_6787);
nand U9059 (N_9059,N_6429,N_6679);
nand U9060 (N_9060,N_6059,N_6126);
nand U9061 (N_9061,N_6318,N_6124);
and U9062 (N_9062,N_6040,N_6129);
nor U9063 (N_9063,N_5048,N_6540);
or U9064 (N_9064,N_7455,N_6824);
nand U9065 (N_9065,N_6935,N_6122);
nor U9066 (N_9066,N_5960,N_5202);
nor U9067 (N_9067,N_6446,N_6226);
nor U9068 (N_9068,N_7325,N_7482);
nand U9069 (N_9069,N_5291,N_5638);
or U9070 (N_9070,N_5192,N_5607);
and U9071 (N_9071,N_5101,N_5695);
or U9072 (N_9072,N_5474,N_6791);
or U9073 (N_9073,N_6884,N_6144);
xor U9074 (N_9074,N_5640,N_7164);
nand U9075 (N_9075,N_6466,N_7137);
or U9076 (N_9076,N_5581,N_6733);
nand U9077 (N_9077,N_5556,N_5395);
nor U9078 (N_9078,N_7176,N_7276);
nand U9079 (N_9079,N_5615,N_6291);
and U9080 (N_9080,N_5693,N_5549);
nor U9081 (N_9081,N_5563,N_5417);
nor U9082 (N_9082,N_6093,N_6854);
nand U9083 (N_9083,N_7174,N_5799);
xnor U9084 (N_9084,N_6251,N_5578);
nand U9085 (N_9085,N_5361,N_7368);
xnor U9086 (N_9086,N_6810,N_5744);
and U9087 (N_9087,N_5170,N_5572);
nand U9088 (N_9088,N_5475,N_6743);
or U9089 (N_9089,N_6637,N_7320);
and U9090 (N_9090,N_5101,N_5357);
or U9091 (N_9091,N_7470,N_6758);
or U9092 (N_9092,N_5044,N_6695);
and U9093 (N_9093,N_6188,N_5167);
and U9094 (N_9094,N_6744,N_7219);
nor U9095 (N_9095,N_6304,N_5279);
or U9096 (N_9096,N_7131,N_6317);
and U9097 (N_9097,N_6404,N_7233);
nand U9098 (N_9098,N_5901,N_5051);
nand U9099 (N_9099,N_6068,N_5543);
nor U9100 (N_9100,N_6574,N_6760);
nor U9101 (N_9101,N_5797,N_6436);
nor U9102 (N_9102,N_5436,N_5328);
nor U9103 (N_9103,N_6385,N_5272);
and U9104 (N_9104,N_6931,N_6219);
xnor U9105 (N_9105,N_6907,N_7220);
or U9106 (N_9106,N_5372,N_5978);
and U9107 (N_9107,N_5073,N_7306);
nand U9108 (N_9108,N_7057,N_5407);
or U9109 (N_9109,N_6605,N_6129);
nand U9110 (N_9110,N_5705,N_7421);
or U9111 (N_9111,N_5426,N_6769);
or U9112 (N_9112,N_5492,N_5223);
nor U9113 (N_9113,N_6439,N_5838);
or U9114 (N_9114,N_6978,N_6006);
and U9115 (N_9115,N_5767,N_5858);
or U9116 (N_9116,N_6086,N_6223);
and U9117 (N_9117,N_5231,N_6666);
nor U9118 (N_9118,N_6567,N_6587);
nand U9119 (N_9119,N_6075,N_5402);
or U9120 (N_9120,N_6018,N_6887);
nand U9121 (N_9121,N_5997,N_5884);
nor U9122 (N_9122,N_7362,N_6067);
and U9123 (N_9123,N_5007,N_6998);
or U9124 (N_9124,N_5029,N_6960);
nand U9125 (N_9125,N_6090,N_7001);
and U9126 (N_9126,N_6279,N_5521);
nor U9127 (N_9127,N_7089,N_7211);
nand U9128 (N_9128,N_6828,N_5766);
nand U9129 (N_9129,N_6350,N_5266);
nor U9130 (N_9130,N_6919,N_7167);
and U9131 (N_9131,N_7313,N_6118);
xor U9132 (N_9132,N_6453,N_6488);
or U9133 (N_9133,N_5411,N_6671);
nor U9134 (N_9134,N_5622,N_6187);
nand U9135 (N_9135,N_5591,N_5311);
nand U9136 (N_9136,N_5445,N_7423);
nor U9137 (N_9137,N_6735,N_5584);
nand U9138 (N_9138,N_5574,N_5397);
or U9139 (N_9139,N_6581,N_6664);
nor U9140 (N_9140,N_6748,N_6998);
nand U9141 (N_9141,N_6295,N_5276);
nand U9142 (N_9142,N_6840,N_6101);
nor U9143 (N_9143,N_5565,N_7037);
nand U9144 (N_9144,N_6077,N_5351);
or U9145 (N_9145,N_5887,N_6938);
nand U9146 (N_9146,N_5103,N_5715);
or U9147 (N_9147,N_5761,N_6225);
nand U9148 (N_9148,N_5168,N_5718);
nand U9149 (N_9149,N_6158,N_6855);
and U9150 (N_9150,N_5631,N_5702);
nand U9151 (N_9151,N_6823,N_6963);
nand U9152 (N_9152,N_7435,N_5026);
nor U9153 (N_9153,N_6297,N_6172);
nand U9154 (N_9154,N_6426,N_6249);
nand U9155 (N_9155,N_6414,N_5971);
nor U9156 (N_9156,N_5545,N_5954);
nor U9157 (N_9157,N_6529,N_6426);
or U9158 (N_9158,N_6257,N_5652);
nor U9159 (N_9159,N_5276,N_5597);
and U9160 (N_9160,N_5349,N_6811);
nand U9161 (N_9161,N_6561,N_5870);
nand U9162 (N_9162,N_5847,N_6327);
or U9163 (N_9163,N_6794,N_5256);
and U9164 (N_9164,N_5716,N_6373);
or U9165 (N_9165,N_5218,N_6226);
nor U9166 (N_9166,N_5251,N_5959);
xnor U9167 (N_9167,N_5097,N_6599);
nor U9168 (N_9168,N_7066,N_6344);
nand U9169 (N_9169,N_6414,N_5011);
or U9170 (N_9170,N_6058,N_7193);
nor U9171 (N_9171,N_6035,N_5237);
nor U9172 (N_9172,N_6017,N_5940);
nand U9173 (N_9173,N_5919,N_6823);
nand U9174 (N_9174,N_6190,N_5552);
or U9175 (N_9175,N_5106,N_6713);
and U9176 (N_9176,N_6683,N_5123);
and U9177 (N_9177,N_5415,N_7189);
and U9178 (N_9178,N_5165,N_6122);
or U9179 (N_9179,N_6063,N_5572);
or U9180 (N_9180,N_7010,N_5273);
and U9181 (N_9181,N_6588,N_5094);
or U9182 (N_9182,N_5084,N_5939);
nor U9183 (N_9183,N_6439,N_5182);
and U9184 (N_9184,N_5656,N_6802);
or U9185 (N_9185,N_5237,N_6031);
nand U9186 (N_9186,N_6883,N_5974);
nor U9187 (N_9187,N_7037,N_6050);
nand U9188 (N_9188,N_7173,N_7351);
nor U9189 (N_9189,N_5160,N_7035);
and U9190 (N_9190,N_5110,N_7284);
and U9191 (N_9191,N_7434,N_6893);
or U9192 (N_9192,N_6182,N_6767);
nor U9193 (N_9193,N_6768,N_6336);
or U9194 (N_9194,N_6607,N_7215);
nand U9195 (N_9195,N_7043,N_7099);
nand U9196 (N_9196,N_7318,N_5632);
nand U9197 (N_9197,N_5551,N_5853);
nor U9198 (N_9198,N_6356,N_5192);
or U9199 (N_9199,N_6548,N_6152);
or U9200 (N_9200,N_6566,N_6510);
nor U9201 (N_9201,N_6205,N_7252);
nand U9202 (N_9202,N_5505,N_5012);
and U9203 (N_9203,N_6114,N_5291);
nor U9204 (N_9204,N_5881,N_7320);
or U9205 (N_9205,N_6103,N_7215);
or U9206 (N_9206,N_6541,N_6636);
or U9207 (N_9207,N_6706,N_7480);
nor U9208 (N_9208,N_7047,N_6233);
or U9209 (N_9209,N_5577,N_6856);
nor U9210 (N_9210,N_5226,N_5701);
nor U9211 (N_9211,N_5714,N_7268);
nand U9212 (N_9212,N_5615,N_6153);
or U9213 (N_9213,N_7456,N_5044);
nor U9214 (N_9214,N_7094,N_6239);
and U9215 (N_9215,N_6155,N_7346);
nor U9216 (N_9216,N_5931,N_5528);
or U9217 (N_9217,N_5274,N_6097);
nor U9218 (N_9218,N_6104,N_6937);
nand U9219 (N_9219,N_5857,N_5703);
nand U9220 (N_9220,N_5375,N_5708);
nand U9221 (N_9221,N_5157,N_5419);
nand U9222 (N_9222,N_7047,N_5108);
nand U9223 (N_9223,N_5849,N_5513);
and U9224 (N_9224,N_5773,N_6678);
nor U9225 (N_9225,N_6260,N_6039);
and U9226 (N_9226,N_5891,N_6847);
and U9227 (N_9227,N_5673,N_7347);
nor U9228 (N_9228,N_6277,N_6134);
xnor U9229 (N_9229,N_6714,N_7426);
nand U9230 (N_9230,N_6006,N_6493);
or U9231 (N_9231,N_5041,N_6714);
nand U9232 (N_9232,N_7452,N_5816);
and U9233 (N_9233,N_5832,N_5830);
or U9234 (N_9234,N_7122,N_5236);
nor U9235 (N_9235,N_7092,N_5455);
nand U9236 (N_9236,N_6085,N_6629);
or U9237 (N_9237,N_7180,N_6955);
nor U9238 (N_9238,N_6018,N_6948);
or U9239 (N_9239,N_5154,N_6381);
or U9240 (N_9240,N_5245,N_6420);
nor U9241 (N_9241,N_5188,N_6185);
xnor U9242 (N_9242,N_7167,N_6184);
and U9243 (N_9243,N_5633,N_5201);
and U9244 (N_9244,N_7033,N_5296);
and U9245 (N_9245,N_6467,N_5472);
nor U9246 (N_9246,N_6451,N_5395);
and U9247 (N_9247,N_6992,N_5599);
or U9248 (N_9248,N_5785,N_6628);
nor U9249 (N_9249,N_5487,N_6342);
nand U9250 (N_9250,N_5122,N_5213);
and U9251 (N_9251,N_5360,N_7001);
and U9252 (N_9252,N_6592,N_6102);
nor U9253 (N_9253,N_6881,N_6377);
nor U9254 (N_9254,N_5315,N_6147);
and U9255 (N_9255,N_5398,N_6296);
or U9256 (N_9256,N_5707,N_6258);
and U9257 (N_9257,N_6222,N_5190);
or U9258 (N_9258,N_7073,N_6322);
and U9259 (N_9259,N_7275,N_6554);
and U9260 (N_9260,N_5051,N_5483);
or U9261 (N_9261,N_6239,N_5523);
or U9262 (N_9262,N_5781,N_6626);
and U9263 (N_9263,N_7063,N_7240);
or U9264 (N_9264,N_5896,N_7363);
nor U9265 (N_9265,N_6844,N_6859);
nand U9266 (N_9266,N_6459,N_5795);
and U9267 (N_9267,N_5167,N_6686);
and U9268 (N_9268,N_5199,N_5509);
nor U9269 (N_9269,N_5470,N_5323);
and U9270 (N_9270,N_6319,N_5047);
and U9271 (N_9271,N_5175,N_6416);
or U9272 (N_9272,N_5250,N_6133);
and U9273 (N_9273,N_7242,N_6162);
nand U9274 (N_9274,N_5994,N_5013);
or U9275 (N_9275,N_5594,N_5264);
and U9276 (N_9276,N_6792,N_5594);
and U9277 (N_9277,N_7163,N_6353);
or U9278 (N_9278,N_6854,N_5940);
nor U9279 (N_9279,N_5325,N_5972);
xor U9280 (N_9280,N_5087,N_5825);
and U9281 (N_9281,N_6700,N_5473);
and U9282 (N_9282,N_6246,N_7158);
or U9283 (N_9283,N_7115,N_7368);
nand U9284 (N_9284,N_5689,N_6726);
or U9285 (N_9285,N_7367,N_5946);
nand U9286 (N_9286,N_6107,N_5465);
nand U9287 (N_9287,N_7456,N_6899);
or U9288 (N_9288,N_6358,N_6317);
nor U9289 (N_9289,N_6761,N_7058);
and U9290 (N_9290,N_5936,N_6248);
or U9291 (N_9291,N_5841,N_5272);
or U9292 (N_9292,N_5215,N_7004);
nand U9293 (N_9293,N_7120,N_6569);
nand U9294 (N_9294,N_7337,N_7442);
nor U9295 (N_9295,N_6169,N_5221);
and U9296 (N_9296,N_5571,N_5117);
and U9297 (N_9297,N_5976,N_6684);
or U9298 (N_9298,N_5184,N_6571);
and U9299 (N_9299,N_5187,N_6812);
and U9300 (N_9300,N_5945,N_5870);
and U9301 (N_9301,N_6513,N_6568);
or U9302 (N_9302,N_5975,N_5237);
nor U9303 (N_9303,N_6094,N_5677);
or U9304 (N_9304,N_7241,N_7369);
nor U9305 (N_9305,N_7020,N_6821);
nand U9306 (N_9306,N_5143,N_5902);
nor U9307 (N_9307,N_5507,N_5114);
nand U9308 (N_9308,N_7260,N_5883);
nand U9309 (N_9309,N_7485,N_6445);
xor U9310 (N_9310,N_6101,N_7030);
nor U9311 (N_9311,N_6665,N_6842);
xor U9312 (N_9312,N_6150,N_7382);
nor U9313 (N_9313,N_5547,N_7348);
nor U9314 (N_9314,N_5204,N_7470);
or U9315 (N_9315,N_5428,N_5582);
and U9316 (N_9316,N_6347,N_6784);
or U9317 (N_9317,N_7278,N_7230);
nand U9318 (N_9318,N_6703,N_6166);
nand U9319 (N_9319,N_5403,N_5221);
or U9320 (N_9320,N_6622,N_6787);
nand U9321 (N_9321,N_5470,N_6335);
nor U9322 (N_9322,N_7360,N_5445);
and U9323 (N_9323,N_6091,N_5731);
nor U9324 (N_9324,N_6341,N_6500);
nand U9325 (N_9325,N_5686,N_5639);
or U9326 (N_9326,N_6357,N_5487);
nor U9327 (N_9327,N_7242,N_6572);
and U9328 (N_9328,N_6040,N_5433);
nor U9329 (N_9329,N_6431,N_7064);
or U9330 (N_9330,N_7137,N_6636);
nor U9331 (N_9331,N_7108,N_6471);
nor U9332 (N_9332,N_6736,N_6273);
nor U9333 (N_9333,N_6477,N_6803);
nand U9334 (N_9334,N_7172,N_7229);
nand U9335 (N_9335,N_5935,N_5805);
and U9336 (N_9336,N_7024,N_6844);
and U9337 (N_9337,N_6323,N_5889);
or U9338 (N_9338,N_7022,N_7237);
or U9339 (N_9339,N_6900,N_7165);
and U9340 (N_9340,N_7446,N_5974);
and U9341 (N_9341,N_5242,N_7003);
or U9342 (N_9342,N_7378,N_6467);
and U9343 (N_9343,N_5849,N_5843);
nor U9344 (N_9344,N_5865,N_6964);
and U9345 (N_9345,N_7375,N_7216);
or U9346 (N_9346,N_6588,N_7218);
xnor U9347 (N_9347,N_6679,N_6910);
nor U9348 (N_9348,N_5799,N_5567);
xor U9349 (N_9349,N_6055,N_5090);
nand U9350 (N_9350,N_5518,N_6044);
nor U9351 (N_9351,N_6869,N_7227);
and U9352 (N_9352,N_7210,N_5288);
and U9353 (N_9353,N_5924,N_6581);
nor U9354 (N_9354,N_5315,N_6474);
or U9355 (N_9355,N_5999,N_5436);
or U9356 (N_9356,N_6394,N_6921);
or U9357 (N_9357,N_7291,N_6265);
nor U9358 (N_9358,N_5396,N_5382);
nor U9359 (N_9359,N_5913,N_7209);
nor U9360 (N_9360,N_5852,N_6833);
and U9361 (N_9361,N_6609,N_5515);
and U9362 (N_9362,N_5333,N_5797);
nor U9363 (N_9363,N_5096,N_7170);
and U9364 (N_9364,N_7038,N_5727);
nor U9365 (N_9365,N_5573,N_5659);
xor U9366 (N_9366,N_5354,N_5473);
nand U9367 (N_9367,N_7143,N_5584);
or U9368 (N_9368,N_5609,N_5464);
nor U9369 (N_9369,N_7483,N_7337);
nor U9370 (N_9370,N_5271,N_5478);
nand U9371 (N_9371,N_6832,N_5073);
or U9372 (N_9372,N_7040,N_7288);
and U9373 (N_9373,N_5052,N_7281);
nor U9374 (N_9374,N_5609,N_5057);
nand U9375 (N_9375,N_5538,N_5456);
or U9376 (N_9376,N_6252,N_6278);
or U9377 (N_9377,N_5911,N_6328);
and U9378 (N_9378,N_6537,N_6938);
and U9379 (N_9379,N_5048,N_5996);
or U9380 (N_9380,N_6960,N_6984);
or U9381 (N_9381,N_5551,N_5979);
and U9382 (N_9382,N_6411,N_5978);
or U9383 (N_9383,N_6694,N_7172);
nor U9384 (N_9384,N_7480,N_5063);
and U9385 (N_9385,N_6763,N_5812);
nor U9386 (N_9386,N_7327,N_6208);
and U9387 (N_9387,N_6183,N_6420);
or U9388 (N_9388,N_5385,N_6634);
and U9389 (N_9389,N_6611,N_6658);
nand U9390 (N_9390,N_6272,N_6153);
nand U9391 (N_9391,N_5899,N_7439);
and U9392 (N_9392,N_5764,N_5228);
or U9393 (N_9393,N_6227,N_7026);
or U9394 (N_9394,N_5393,N_5078);
nor U9395 (N_9395,N_6154,N_5116);
and U9396 (N_9396,N_6537,N_6146);
nor U9397 (N_9397,N_5849,N_6447);
xor U9398 (N_9398,N_6401,N_6683);
or U9399 (N_9399,N_6509,N_5874);
nor U9400 (N_9400,N_6361,N_5279);
xnor U9401 (N_9401,N_6311,N_7321);
and U9402 (N_9402,N_5321,N_5989);
or U9403 (N_9403,N_6272,N_5280);
nand U9404 (N_9404,N_6311,N_6320);
and U9405 (N_9405,N_6685,N_5201);
nor U9406 (N_9406,N_6603,N_5354);
nand U9407 (N_9407,N_6463,N_6732);
and U9408 (N_9408,N_6954,N_5913);
and U9409 (N_9409,N_6103,N_5647);
or U9410 (N_9410,N_6503,N_6559);
or U9411 (N_9411,N_5899,N_6267);
and U9412 (N_9412,N_6967,N_6844);
or U9413 (N_9413,N_5089,N_7343);
or U9414 (N_9414,N_7473,N_6411);
and U9415 (N_9415,N_6150,N_6494);
nand U9416 (N_9416,N_5991,N_5282);
and U9417 (N_9417,N_6502,N_6187);
nand U9418 (N_9418,N_6269,N_6510);
or U9419 (N_9419,N_6629,N_5200);
nand U9420 (N_9420,N_6797,N_6317);
and U9421 (N_9421,N_5568,N_5673);
and U9422 (N_9422,N_6942,N_6003);
and U9423 (N_9423,N_6786,N_5465);
nor U9424 (N_9424,N_5250,N_5732);
or U9425 (N_9425,N_7232,N_5576);
and U9426 (N_9426,N_6916,N_6045);
nand U9427 (N_9427,N_6041,N_6595);
or U9428 (N_9428,N_6356,N_6647);
nor U9429 (N_9429,N_5593,N_5878);
or U9430 (N_9430,N_7040,N_5946);
nand U9431 (N_9431,N_6914,N_6280);
and U9432 (N_9432,N_7130,N_5769);
and U9433 (N_9433,N_5169,N_6500);
nand U9434 (N_9434,N_5661,N_5851);
or U9435 (N_9435,N_6154,N_6129);
or U9436 (N_9436,N_5999,N_7198);
nand U9437 (N_9437,N_6946,N_5089);
or U9438 (N_9438,N_6893,N_7366);
nor U9439 (N_9439,N_5352,N_6617);
or U9440 (N_9440,N_6792,N_6032);
nor U9441 (N_9441,N_5691,N_7287);
and U9442 (N_9442,N_5259,N_6049);
and U9443 (N_9443,N_5666,N_6146);
nand U9444 (N_9444,N_7422,N_5146);
and U9445 (N_9445,N_5543,N_5358);
nor U9446 (N_9446,N_5547,N_6249);
nand U9447 (N_9447,N_5840,N_5611);
nand U9448 (N_9448,N_6467,N_6115);
and U9449 (N_9449,N_5210,N_7119);
or U9450 (N_9450,N_5514,N_5400);
and U9451 (N_9451,N_6977,N_7435);
nand U9452 (N_9452,N_5163,N_5653);
or U9453 (N_9453,N_6374,N_6146);
nor U9454 (N_9454,N_5351,N_5977);
nor U9455 (N_9455,N_6902,N_5202);
nor U9456 (N_9456,N_7232,N_5072);
and U9457 (N_9457,N_5859,N_6937);
xnor U9458 (N_9458,N_7205,N_6855);
nand U9459 (N_9459,N_5282,N_6563);
nor U9460 (N_9460,N_6266,N_6169);
nor U9461 (N_9461,N_6182,N_7408);
nor U9462 (N_9462,N_6263,N_6370);
nor U9463 (N_9463,N_5770,N_7376);
or U9464 (N_9464,N_6586,N_6078);
or U9465 (N_9465,N_5764,N_6933);
nor U9466 (N_9466,N_5478,N_6973);
xor U9467 (N_9467,N_6135,N_5701);
nor U9468 (N_9468,N_7198,N_5114);
nand U9469 (N_9469,N_5665,N_5367);
nand U9470 (N_9470,N_6656,N_6403);
and U9471 (N_9471,N_7474,N_5644);
and U9472 (N_9472,N_6931,N_6528);
and U9473 (N_9473,N_6972,N_6195);
or U9474 (N_9474,N_5871,N_5563);
or U9475 (N_9475,N_7362,N_5728);
nand U9476 (N_9476,N_6979,N_7414);
or U9477 (N_9477,N_7011,N_5413);
or U9478 (N_9478,N_7087,N_6320);
nor U9479 (N_9479,N_7304,N_5645);
and U9480 (N_9480,N_5585,N_7461);
or U9481 (N_9481,N_5233,N_6818);
and U9482 (N_9482,N_5626,N_5556);
nor U9483 (N_9483,N_5376,N_5272);
or U9484 (N_9484,N_7136,N_5146);
and U9485 (N_9485,N_6698,N_6593);
or U9486 (N_9486,N_5101,N_6144);
nor U9487 (N_9487,N_7431,N_6559);
xor U9488 (N_9488,N_7151,N_5260);
nor U9489 (N_9489,N_7024,N_6069);
and U9490 (N_9490,N_6515,N_5851);
nand U9491 (N_9491,N_6859,N_5433);
and U9492 (N_9492,N_5216,N_5226);
or U9493 (N_9493,N_6585,N_6743);
nor U9494 (N_9494,N_7139,N_6386);
nand U9495 (N_9495,N_7208,N_6818);
nor U9496 (N_9496,N_7178,N_5794);
and U9497 (N_9497,N_7278,N_5450);
xor U9498 (N_9498,N_5691,N_7297);
nor U9499 (N_9499,N_7460,N_5510);
and U9500 (N_9500,N_6347,N_5529);
nand U9501 (N_9501,N_6468,N_5319);
and U9502 (N_9502,N_7462,N_5731);
nand U9503 (N_9503,N_6032,N_7124);
and U9504 (N_9504,N_7476,N_5894);
and U9505 (N_9505,N_5713,N_6854);
nor U9506 (N_9506,N_5582,N_6857);
nand U9507 (N_9507,N_6875,N_6591);
and U9508 (N_9508,N_5992,N_5758);
nand U9509 (N_9509,N_6594,N_5999);
and U9510 (N_9510,N_6896,N_5157);
nand U9511 (N_9511,N_5008,N_7461);
nand U9512 (N_9512,N_7494,N_5567);
or U9513 (N_9513,N_5542,N_7398);
or U9514 (N_9514,N_5468,N_5027);
nand U9515 (N_9515,N_5471,N_5514);
or U9516 (N_9516,N_5897,N_6493);
or U9517 (N_9517,N_6538,N_6897);
or U9518 (N_9518,N_6673,N_5170);
nand U9519 (N_9519,N_7081,N_6445);
and U9520 (N_9520,N_7013,N_6947);
and U9521 (N_9521,N_5311,N_6364);
or U9522 (N_9522,N_7460,N_6280);
and U9523 (N_9523,N_7216,N_5389);
nor U9524 (N_9524,N_6495,N_6991);
nor U9525 (N_9525,N_5832,N_5290);
and U9526 (N_9526,N_6872,N_5544);
nor U9527 (N_9527,N_7490,N_6809);
nand U9528 (N_9528,N_5040,N_6458);
nor U9529 (N_9529,N_5561,N_5980);
nor U9530 (N_9530,N_5270,N_6674);
or U9531 (N_9531,N_7234,N_7315);
or U9532 (N_9532,N_6372,N_6957);
and U9533 (N_9533,N_7010,N_5325);
nor U9534 (N_9534,N_7098,N_7041);
and U9535 (N_9535,N_6209,N_7360);
and U9536 (N_9536,N_5734,N_6499);
and U9537 (N_9537,N_6461,N_6393);
or U9538 (N_9538,N_5227,N_7226);
and U9539 (N_9539,N_6364,N_5865);
or U9540 (N_9540,N_5127,N_6935);
and U9541 (N_9541,N_6566,N_7340);
nor U9542 (N_9542,N_6753,N_6516);
nor U9543 (N_9543,N_5287,N_7188);
or U9544 (N_9544,N_6435,N_5877);
nand U9545 (N_9545,N_5853,N_6412);
and U9546 (N_9546,N_6651,N_5689);
nor U9547 (N_9547,N_5600,N_7044);
or U9548 (N_9548,N_7026,N_6902);
nor U9549 (N_9549,N_5970,N_5644);
or U9550 (N_9550,N_5534,N_5014);
and U9551 (N_9551,N_6529,N_5092);
nand U9552 (N_9552,N_6043,N_5965);
nand U9553 (N_9553,N_5708,N_5829);
or U9554 (N_9554,N_6043,N_5598);
or U9555 (N_9555,N_5776,N_6258);
and U9556 (N_9556,N_5588,N_5101);
or U9557 (N_9557,N_6417,N_5491);
and U9558 (N_9558,N_6841,N_6344);
nand U9559 (N_9559,N_5146,N_6136);
or U9560 (N_9560,N_7229,N_5727);
nor U9561 (N_9561,N_5106,N_6317);
nand U9562 (N_9562,N_6012,N_6152);
and U9563 (N_9563,N_5250,N_7063);
and U9564 (N_9564,N_5528,N_6615);
and U9565 (N_9565,N_7126,N_5152);
nor U9566 (N_9566,N_5746,N_7340);
and U9567 (N_9567,N_7128,N_7106);
or U9568 (N_9568,N_7095,N_7072);
nand U9569 (N_9569,N_7460,N_6454);
xor U9570 (N_9570,N_6984,N_5375);
nor U9571 (N_9571,N_6087,N_6126);
or U9572 (N_9572,N_5215,N_7042);
nand U9573 (N_9573,N_7314,N_5467);
and U9574 (N_9574,N_6993,N_5108);
or U9575 (N_9575,N_5774,N_7485);
or U9576 (N_9576,N_5388,N_6217);
nor U9577 (N_9577,N_7078,N_7147);
or U9578 (N_9578,N_6727,N_6398);
nand U9579 (N_9579,N_6442,N_5889);
nand U9580 (N_9580,N_6332,N_7433);
or U9581 (N_9581,N_5427,N_6826);
xor U9582 (N_9582,N_6902,N_6090);
xor U9583 (N_9583,N_5655,N_6495);
or U9584 (N_9584,N_6606,N_7338);
xor U9585 (N_9585,N_5834,N_5104);
or U9586 (N_9586,N_6206,N_7435);
and U9587 (N_9587,N_6434,N_6144);
nor U9588 (N_9588,N_6717,N_5093);
nand U9589 (N_9589,N_5987,N_6643);
nor U9590 (N_9590,N_7106,N_6862);
and U9591 (N_9591,N_7205,N_6892);
and U9592 (N_9592,N_5363,N_5941);
nor U9593 (N_9593,N_6171,N_5622);
or U9594 (N_9594,N_7338,N_6515);
nor U9595 (N_9595,N_5263,N_6966);
or U9596 (N_9596,N_5988,N_6458);
nand U9597 (N_9597,N_6141,N_6967);
or U9598 (N_9598,N_6408,N_6383);
xnor U9599 (N_9599,N_5516,N_7248);
or U9600 (N_9600,N_5426,N_5820);
nor U9601 (N_9601,N_7451,N_7181);
nor U9602 (N_9602,N_5114,N_5522);
or U9603 (N_9603,N_6160,N_5197);
nand U9604 (N_9604,N_7268,N_6026);
nand U9605 (N_9605,N_6199,N_6529);
nor U9606 (N_9606,N_5314,N_5904);
nand U9607 (N_9607,N_5275,N_7111);
and U9608 (N_9608,N_5574,N_6245);
nor U9609 (N_9609,N_7429,N_7360);
nand U9610 (N_9610,N_5734,N_5309);
nand U9611 (N_9611,N_6448,N_6437);
or U9612 (N_9612,N_7041,N_7181);
and U9613 (N_9613,N_5410,N_6233);
and U9614 (N_9614,N_5719,N_6494);
nand U9615 (N_9615,N_6939,N_5597);
and U9616 (N_9616,N_5637,N_6328);
nor U9617 (N_9617,N_6888,N_5098);
nor U9618 (N_9618,N_6006,N_7409);
or U9619 (N_9619,N_5585,N_7013);
nand U9620 (N_9620,N_6008,N_6616);
or U9621 (N_9621,N_6763,N_6485);
nand U9622 (N_9622,N_5717,N_7022);
nor U9623 (N_9623,N_7206,N_5157);
xor U9624 (N_9624,N_6117,N_6929);
nor U9625 (N_9625,N_5225,N_5434);
and U9626 (N_9626,N_6610,N_5144);
nand U9627 (N_9627,N_5178,N_5618);
or U9628 (N_9628,N_5059,N_5705);
nor U9629 (N_9629,N_6755,N_5116);
nand U9630 (N_9630,N_6045,N_7457);
and U9631 (N_9631,N_5446,N_6539);
or U9632 (N_9632,N_7072,N_5750);
nand U9633 (N_9633,N_6394,N_6856);
and U9634 (N_9634,N_7236,N_5553);
xnor U9635 (N_9635,N_6199,N_6834);
and U9636 (N_9636,N_7372,N_5422);
and U9637 (N_9637,N_5772,N_5700);
and U9638 (N_9638,N_6401,N_6200);
and U9639 (N_9639,N_6001,N_7310);
and U9640 (N_9640,N_7163,N_6336);
nand U9641 (N_9641,N_5287,N_5730);
nor U9642 (N_9642,N_6124,N_6830);
or U9643 (N_9643,N_5829,N_7401);
and U9644 (N_9644,N_6356,N_6104);
xnor U9645 (N_9645,N_7365,N_7232);
nor U9646 (N_9646,N_5017,N_6188);
or U9647 (N_9647,N_5764,N_5936);
or U9648 (N_9648,N_5639,N_5934);
nand U9649 (N_9649,N_6291,N_6040);
nand U9650 (N_9650,N_5121,N_6478);
xor U9651 (N_9651,N_6645,N_7376);
nor U9652 (N_9652,N_6615,N_6084);
nor U9653 (N_9653,N_5000,N_5939);
nor U9654 (N_9654,N_6190,N_6772);
and U9655 (N_9655,N_5294,N_5406);
or U9656 (N_9656,N_5553,N_6538);
nor U9657 (N_9657,N_6378,N_5736);
nand U9658 (N_9658,N_6955,N_6587);
nor U9659 (N_9659,N_6137,N_5116);
and U9660 (N_9660,N_5302,N_6061);
and U9661 (N_9661,N_7209,N_6881);
nor U9662 (N_9662,N_5782,N_5899);
nand U9663 (N_9663,N_5331,N_6634);
nand U9664 (N_9664,N_6941,N_6948);
or U9665 (N_9665,N_6268,N_6055);
nand U9666 (N_9666,N_5634,N_7009);
and U9667 (N_9667,N_6796,N_6398);
nand U9668 (N_9668,N_7467,N_7148);
nand U9669 (N_9669,N_7115,N_6938);
and U9670 (N_9670,N_7143,N_5999);
nor U9671 (N_9671,N_7277,N_6983);
nor U9672 (N_9672,N_6655,N_5332);
nand U9673 (N_9673,N_5293,N_6917);
nand U9674 (N_9674,N_6184,N_6042);
nand U9675 (N_9675,N_6870,N_7215);
and U9676 (N_9676,N_5394,N_6894);
and U9677 (N_9677,N_5430,N_6149);
nand U9678 (N_9678,N_5175,N_7358);
and U9679 (N_9679,N_6870,N_7026);
nor U9680 (N_9680,N_6256,N_6999);
nand U9681 (N_9681,N_5460,N_7279);
xor U9682 (N_9682,N_5615,N_5297);
nand U9683 (N_9683,N_6269,N_7284);
nand U9684 (N_9684,N_6523,N_6054);
nor U9685 (N_9685,N_5114,N_6569);
nor U9686 (N_9686,N_5119,N_6028);
or U9687 (N_9687,N_6638,N_7168);
and U9688 (N_9688,N_5706,N_6879);
nor U9689 (N_9689,N_7420,N_5631);
and U9690 (N_9690,N_7295,N_5380);
or U9691 (N_9691,N_7015,N_5593);
xnor U9692 (N_9692,N_5441,N_5051);
or U9693 (N_9693,N_6401,N_5411);
nand U9694 (N_9694,N_7288,N_5143);
nand U9695 (N_9695,N_5566,N_6478);
xnor U9696 (N_9696,N_7197,N_6793);
and U9697 (N_9697,N_5829,N_7015);
and U9698 (N_9698,N_6156,N_5105);
nand U9699 (N_9699,N_5049,N_6181);
nor U9700 (N_9700,N_7481,N_6028);
and U9701 (N_9701,N_5882,N_5584);
and U9702 (N_9702,N_6686,N_7356);
or U9703 (N_9703,N_6093,N_6300);
nor U9704 (N_9704,N_5891,N_7285);
nor U9705 (N_9705,N_6055,N_6331);
nor U9706 (N_9706,N_5983,N_5992);
nor U9707 (N_9707,N_7158,N_5562);
nand U9708 (N_9708,N_7276,N_5404);
or U9709 (N_9709,N_7088,N_5680);
or U9710 (N_9710,N_5037,N_6407);
and U9711 (N_9711,N_6350,N_5407);
or U9712 (N_9712,N_5687,N_5782);
nor U9713 (N_9713,N_5836,N_6137);
nor U9714 (N_9714,N_7479,N_6698);
nor U9715 (N_9715,N_5255,N_5706);
and U9716 (N_9716,N_6883,N_6733);
nor U9717 (N_9717,N_7033,N_5138);
or U9718 (N_9718,N_7101,N_6167);
nand U9719 (N_9719,N_6417,N_7291);
nor U9720 (N_9720,N_5642,N_7422);
and U9721 (N_9721,N_5733,N_6096);
and U9722 (N_9722,N_6830,N_6130);
or U9723 (N_9723,N_6328,N_5536);
or U9724 (N_9724,N_5632,N_5740);
and U9725 (N_9725,N_7418,N_6024);
or U9726 (N_9726,N_5846,N_7367);
and U9727 (N_9727,N_6186,N_7117);
nor U9728 (N_9728,N_5192,N_6211);
and U9729 (N_9729,N_6089,N_6889);
nand U9730 (N_9730,N_7444,N_7442);
or U9731 (N_9731,N_5595,N_6023);
xor U9732 (N_9732,N_5134,N_7418);
nor U9733 (N_9733,N_6466,N_6505);
nand U9734 (N_9734,N_6855,N_5504);
nor U9735 (N_9735,N_6557,N_7120);
xnor U9736 (N_9736,N_7006,N_7255);
and U9737 (N_9737,N_5912,N_5313);
nand U9738 (N_9738,N_5237,N_6203);
and U9739 (N_9739,N_5285,N_6018);
or U9740 (N_9740,N_6347,N_5998);
or U9741 (N_9741,N_6929,N_6347);
nor U9742 (N_9742,N_6338,N_7006);
and U9743 (N_9743,N_7239,N_6476);
or U9744 (N_9744,N_5267,N_6519);
nor U9745 (N_9745,N_5069,N_5731);
nand U9746 (N_9746,N_7068,N_6985);
nor U9747 (N_9747,N_6952,N_5588);
or U9748 (N_9748,N_6578,N_5650);
nor U9749 (N_9749,N_6175,N_7334);
or U9750 (N_9750,N_6644,N_6089);
nor U9751 (N_9751,N_7226,N_5916);
and U9752 (N_9752,N_6470,N_6085);
or U9753 (N_9753,N_6836,N_7152);
nand U9754 (N_9754,N_5040,N_5537);
xnor U9755 (N_9755,N_6955,N_5816);
and U9756 (N_9756,N_5144,N_7335);
or U9757 (N_9757,N_5149,N_6220);
or U9758 (N_9758,N_5102,N_5945);
nand U9759 (N_9759,N_5535,N_5519);
or U9760 (N_9760,N_7120,N_6185);
nor U9761 (N_9761,N_5233,N_5679);
xnor U9762 (N_9762,N_6777,N_5791);
xor U9763 (N_9763,N_7125,N_5592);
nor U9764 (N_9764,N_5197,N_5302);
and U9765 (N_9765,N_6335,N_5768);
nor U9766 (N_9766,N_5006,N_7407);
or U9767 (N_9767,N_5742,N_6414);
nor U9768 (N_9768,N_7204,N_6791);
nor U9769 (N_9769,N_6913,N_5120);
and U9770 (N_9770,N_6414,N_5749);
nor U9771 (N_9771,N_5814,N_6734);
and U9772 (N_9772,N_5467,N_6957);
and U9773 (N_9773,N_6216,N_6541);
or U9774 (N_9774,N_5734,N_6420);
or U9775 (N_9775,N_7427,N_6762);
nand U9776 (N_9776,N_5540,N_6596);
and U9777 (N_9777,N_5610,N_7326);
nor U9778 (N_9778,N_6822,N_6465);
nor U9779 (N_9779,N_7023,N_5623);
nor U9780 (N_9780,N_6082,N_5071);
or U9781 (N_9781,N_5708,N_5659);
nand U9782 (N_9782,N_6655,N_7459);
nand U9783 (N_9783,N_5774,N_6159);
or U9784 (N_9784,N_5105,N_7032);
nor U9785 (N_9785,N_6914,N_5081);
nand U9786 (N_9786,N_5585,N_6852);
nand U9787 (N_9787,N_7234,N_6444);
and U9788 (N_9788,N_6816,N_6399);
and U9789 (N_9789,N_6668,N_5388);
and U9790 (N_9790,N_6286,N_5048);
nand U9791 (N_9791,N_6053,N_7088);
and U9792 (N_9792,N_6832,N_5918);
nor U9793 (N_9793,N_5062,N_5373);
or U9794 (N_9794,N_6252,N_6240);
and U9795 (N_9795,N_6730,N_7394);
nand U9796 (N_9796,N_5670,N_5538);
and U9797 (N_9797,N_5269,N_5197);
nand U9798 (N_9798,N_6429,N_5280);
and U9799 (N_9799,N_7452,N_6306);
and U9800 (N_9800,N_6871,N_5490);
nand U9801 (N_9801,N_6440,N_6330);
xnor U9802 (N_9802,N_6287,N_7017);
nand U9803 (N_9803,N_5373,N_6262);
nor U9804 (N_9804,N_5801,N_5309);
xor U9805 (N_9805,N_7405,N_6776);
nand U9806 (N_9806,N_7058,N_7242);
and U9807 (N_9807,N_6344,N_7348);
nor U9808 (N_9808,N_5055,N_5989);
nor U9809 (N_9809,N_5536,N_6057);
nor U9810 (N_9810,N_5026,N_5480);
or U9811 (N_9811,N_6438,N_5057);
or U9812 (N_9812,N_6842,N_5699);
nor U9813 (N_9813,N_7282,N_7038);
and U9814 (N_9814,N_6124,N_5893);
or U9815 (N_9815,N_7425,N_7060);
nor U9816 (N_9816,N_6737,N_5261);
and U9817 (N_9817,N_7466,N_6115);
and U9818 (N_9818,N_6587,N_5623);
nor U9819 (N_9819,N_6312,N_5399);
and U9820 (N_9820,N_6359,N_5926);
xor U9821 (N_9821,N_7117,N_7482);
nand U9822 (N_9822,N_6400,N_5383);
or U9823 (N_9823,N_5425,N_6045);
nor U9824 (N_9824,N_6255,N_5903);
or U9825 (N_9825,N_6417,N_5616);
or U9826 (N_9826,N_6307,N_6148);
and U9827 (N_9827,N_6494,N_7264);
nor U9828 (N_9828,N_7158,N_7153);
and U9829 (N_9829,N_6548,N_5611);
nand U9830 (N_9830,N_6673,N_6844);
or U9831 (N_9831,N_5331,N_5463);
nor U9832 (N_9832,N_5226,N_6910);
or U9833 (N_9833,N_6754,N_5561);
nand U9834 (N_9834,N_5028,N_5353);
nand U9835 (N_9835,N_7423,N_5845);
nand U9836 (N_9836,N_6513,N_5813);
nor U9837 (N_9837,N_7185,N_5342);
nand U9838 (N_9838,N_7047,N_6165);
or U9839 (N_9839,N_7119,N_5208);
nand U9840 (N_9840,N_6956,N_6996);
or U9841 (N_9841,N_5945,N_5984);
nor U9842 (N_9842,N_5449,N_5863);
and U9843 (N_9843,N_5885,N_6657);
or U9844 (N_9844,N_7433,N_7468);
or U9845 (N_9845,N_6344,N_6430);
nand U9846 (N_9846,N_5157,N_5026);
nand U9847 (N_9847,N_5151,N_5202);
or U9848 (N_9848,N_5970,N_6896);
and U9849 (N_9849,N_5228,N_5939);
and U9850 (N_9850,N_5912,N_5259);
nand U9851 (N_9851,N_5707,N_7138);
nor U9852 (N_9852,N_7482,N_5912);
nor U9853 (N_9853,N_6109,N_6249);
and U9854 (N_9854,N_7057,N_5787);
or U9855 (N_9855,N_6061,N_6002);
and U9856 (N_9856,N_7226,N_5642);
or U9857 (N_9857,N_5084,N_6047);
xnor U9858 (N_9858,N_5285,N_5718);
nand U9859 (N_9859,N_5142,N_6630);
or U9860 (N_9860,N_5989,N_5741);
nor U9861 (N_9861,N_6446,N_7356);
nor U9862 (N_9862,N_5021,N_7413);
nand U9863 (N_9863,N_5123,N_6826);
and U9864 (N_9864,N_6967,N_5124);
and U9865 (N_9865,N_6455,N_5054);
or U9866 (N_9866,N_6255,N_5468);
nand U9867 (N_9867,N_5550,N_5677);
or U9868 (N_9868,N_5233,N_6111);
nor U9869 (N_9869,N_6881,N_6409);
and U9870 (N_9870,N_5764,N_5534);
nand U9871 (N_9871,N_6436,N_5963);
and U9872 (N_9872,N_5623,N_6307);
and U9873 (N_9873,N_5012,N_6393);
and U9874 (N_9874,N_6384,N_6341);
nor U9875 (N_9875,N_6243,N_5802);
nor U9876 (N_9876,N_5553,N_6651);
or U9877 (N_9877,N_5006,N_5718);
or U9878 (N_9878,N_5870,N_5141);
nand U9879 (N_9879,N_5602,N_7335);
nor U9880 (N_9880,N_7186,N_7382);
or U9881 (N_9881,N_5074,N_6499);
nor U9882 (N_9882,N_6509,N_5002);
nand U9883 (N_9883,N_5469,N_7439);
and U9884 (N_9884,N_6538,N_6689);
nor U9885 (N_9885,N_7369,N_6003);
nor U9886 (N_9886,N_6997,N_5484);
and U9887 (N_9887,N_6770,N_5866);
and U9888 (N_9888,N_6469,N_5692);
and U9889 (N_9889,N_7254,N_5925);
nor U9890 (N_9890,N_6242,N_6310);
nand U9891 (N_9891,N_5659,N_5837);
nor U9892 (N_9892,N_6189,N_6611);
nand U9893 (N_9893,N_6616,N_7152);
or U9894 (N_9894,N_5138,N_5860);
and U9895 (N_9895,N_5003,N_6582);
nand U9896 (N_9896,N_6788,N_7486);
and U9897 (N_9897,N_7218,N_6986);
nor U9898 (N_9898,N_6363,N_6855);
nor U9899 (N_9899,N_6575,N_6659);
nand U9900 (N_9900,N_7206,N_5632);
nor U9901 (N_9901,N_7319,N_7342);
or U9902 (N_9902,N_6647,N_6965);
nor U9903 (N_9903,N_7058,N_5235);
and U9904 (N_9904,N_5518,N_6393);
nor U9905 (N_9905,N_5331,N_7245);
nor U9906 (N_9906,N_5401,N_7200);
or U9907 (N_9907,N_7398,N_6866);
nor U9908 (N_9908,N_7010,N_6498);
or U9909 (N_9909,N_5957,N_5916);
nand U9910 (N_9910,N_5393,N_6043);
and U9911 (N_9911,N_7266,N_5580);
xnor U9912 (N_9912,N_5137,N_7128);
nand U9913 (N_9913,N_6886,N_6579);
nand U9914 (N_9914,N_7084,N_5071);
or U9915 (N_9915,N_5832,N_7491);
nor U9916 (N_9916,N_6911,N_5788);
or U9917 (N_9917,N_5452,N_5282);
nand U9918 (N_9918,N_6686,N_5636);
nand U9919 (N_9919,N_7062,N_5213);
and U9920 (N_9920,N_5082,N_6811);
nor U9921 (N_9921,N_5570,N_7337);
nor U9922 (N_9922,N_5135,N_5115);
nand U9923 (N_9923,N_6696,N_5395);
and U9924 (N_9924,N_7092,N_5099);
and U9925 (N_9925,N_5670,N_5522);
and U9926 (N_9926,N_6609,N_6321);
nand U9927 (N_9927,N_7040,N_5530);
and U9928 (N_9928,N_6351,N_6826);
nor U9929 (N_9929,N_7490,N_6232);
or U9930 (N_9930,N_7372,N_6447);
and U9931 (N_9931,N_5083,N_6198);
and U9932 (N_9932,N_5729,N_6878);
xor U9933 (N_9933,N_7120,N_5035);
nor U9934 (N_9934,N_7420,N_6712);
or U9935 (N_9935,N_5818,N_5972);
nand U9936 (N_9936,N_6262,N_5076);
and U9937 (N_9937,N_5718,N_6003);
or U9938 (N_9938,N_5374,N_5476);
or U9939 (N_9939,N_6181,N_5869);
nor U9940 (N_9940,N_5240,N_6469);
xnor U9941 (N_9941,N_5743,N_5199);
or U9942 (N_9942,N_6480,N_5088);
nor U9943 (N_9943,N_6721,N_6299);
nor U9944 (N_9944,N_5617,N_5942);
nand U9945 (N_9945,N_7000,N_6464);
nor U9946 (N_9946,N_5207,N_6951);
nand U9947 (N_9947,N_6223,N_7171);
nor U9948 (N_9948,N_6029,N_6416);
or U9949 (N_9949,N_5225,N_7490);
or U9950 (N_9950,N_7054,N_5958);
or U9951 (N_9951,N_6998,N_7440);
nor U9952 (N_9952,N_7341,N_5027);
nor U9953 (N_9953,N_5955,N_7054);
and U9954 (N_9954,N_5807,N_6244);
nor U9955 (N_9955,N_7130,N_6000);
or U9956 (N_9956,N_5714,N_6882);
or U9957 (N_9957,N_6983,N_5277);
or U9958 (N_9958,N_6635,N_6897);
nand U9959 (N_9959,N_7269,N_6411);
nand U9960 (N_9960,N_5444,N_6286);
and U9961 (N_9961,N_6384,N_6262);
nand U9962 (N_9962,N_6669,N_6888);
or U9963 (N_9963,N_5438,N_6733);
nand U9964 (N_9964,N_5591,N_7249);
and U9965 (N_9965,N_6724,N_6619);
or U9966 (N_9966,N_6471,N_5020);
or U9967 (N_9967,N_7411,N_6701);
and U9968 (N_9968,N_5752,N_5898);
or U9969 (N_9969,N_6721,N_6491);
nand U9970 (N_9970,N_5563,N_7079);
nor U9971 (N_9971,N_6759,N_5759);
nor U9972 (N_9972,N_5629,N_6105);
and U9973 (N_9973,N_6392,N_5248);
nand U9974 (N_9974,N_6611,N_5493);
or U9975 (N_9975,N_5351,N_7099);
and U9976 (N_9976,N_5621,N_6812);
or U9977 (N_9977,N_6684,N_7159);
or U9978 (N_9978,N_6353,N_6633);
nand U9979 (N_9979,N_5190,N_5926);
nor U9980 (N_9980,N_5323,N_7340);
or U9981 (N_9981,N_6052,N_5614);
nor U9982 (N_9982,N_5016,N_6354);
nor U9983 (N_9983,N_5684,N_7122);
nor U9984 (N_9984,N_6173,N_7275);
nand U9985 (N_9985,N_6902,N_7413);
nor U9986 (N_9986,N_6898,N_5006);
nor U9987 (N_9987,N_7383,N_7409);
and U9988 (N_9988,N_5456,N_6983);
nand U9989 (N_9989,N_6015,N_6798);
or U9990 (N_9990,N_5766,N_7212);
nand U9991 (N_9991,N_7372,N_6026);
nand U9992 (N_9992,N_5259,N_5058);
nor U9993 (N_9993,N_5599,N_5161);
nor U9994 (N_9994,N_5884,N_5699);
nand U9995 (N_9995,N_6077,N_6360);
or U9996 (N_9996,N_5631,N_5275);
nor U9997 (N_9997,N_6637,N_6207);
or U9998 (N_9998,N_6633,N_6722);
nor U9999 (N_9999,N_5894,N_7016);
and UO_0 (O_0,N_9379,N_8505);
and UO_1 (O_1,N_9268,N_8297);
and UO_2 (O_2,N_7656,N_8471);
nand UO_3 (O_3,N_7724,N_8462);
or UO_4 (O_4,N_9093,N_8424);
and UO_5 (O_5,N_8710,N_8705);
or UO_6 (O_6,N_7616,N_8496);
and UO_7 (O_7,N_9127,N_8659);
nor UO_8 (O_8,N_9369,N_7844);
and UO_9 (O_9,N_8727,N_8841);
nand UO_10 (O_10,N_8794,N_7636);
nor UO_11 (O_11,N_8222,N_9508);
nand UO_12 (O_12,N_9538,N_9961);
and UO_13 (O_13,N_8316,N_7903);
or UO_14 (O_14,N_8272,N_8388);
nand UO_15 (O_15,N_7852,N_8582);
nand UO_16 (O_16,N_9677,N_8457);
or UO_17 (O_17,N_9329,N_7750);
and UO_18 (O_18,N_8153,N_8818);
nand UO_19 (O_19,N_8939,N_7605);
or UO_20 (O_20,N_9852,N_9381);
nand UO_21 (O_21,N_8867,N_8121);
nor UO_22 (O_22,N_8674,N_8355);
and UO_23 (O_23,N_9750,N_9260);
and UO_24 (O_24,N_7836,N_8732);
nand UO_25 (O_25,N_8797,N_8994);
nand UO_26 (O_26,N_9294,N_9086);
and UO_27 (O_27,N_9546,N_8651);
nor UO_28 (O_28,N_8545,N_9194);
nand UO_29 (O_29,N_8429,N_8661);
and UO_30 (O_30,N_8416,N_7709);
and UO_31 (O_31,N_8100,N_7807);
nand UO_32 (O_32,N_9461,N_9905);
nand UO_33 (O_33,N_9278,N_8967);
nor UO_34 (O_34,N_8996,N_8176);
nor UO_35 (O_35,N_8893,N_8826);
and UO_36 (O_36,N_8790,N_7869);
or UO_37 (O_37,N_9238,N_8615);
nor UO_38 (O_38,N_8387,N_8850);
nand UO_39 (O_39,N_8979,N_7774);
xnor UO_40 (O_40,N_9046,N_9516);
or UO_41 (O_41,N_8108,N_9535);
nand UO_42 (O_42,N_9228,N_8959);
or UO_43 (O_43,N_8601,N_8626);
or UO_44 (O_44,N_8037,N_8776);
or UO_45 (O_45,N_8948,N_8629);
or UO_46 (O_46,N_7984,N_9235);
and UO_47 (O_47,N_8420,N_8354);
or UO_48 (O_48,N_9080,N_8603);
and UO_49 (O_49,N_9200,N_9050);
nor UO_50 (O_50,N_7883,N_9747);
and UO_51 (O_51,N_9533,N_9934);
or UO_52 (O_52,N_9201,N_7940);
or UO_53 (O_53,N_9659,N_9562);
and UO_54 (O_54,N_9174,N_7973);
nand UO_55 (O_55,N_7783,N_9156);
xnor UO_56 (O_56,N_9146,N_9366);
or UO_57 (O_57,N_7968,N_9950);
nor UO_58 (O_58,N_8038,N_8785);
nand UO_59 (O_59,N_8061,N_9143);
and UO_60 (O_60,N_7592,N_8366);
nor UO_61 (O_61,N_7582,N_8908);
and UO_62 (O_62,N_8623,N_9343);
xor UO_63 (O_63,N_9918,N_7812);
or UO_64 (O_64,N_9488,N_7822);
and UO_65 (O_65,N_8305,N_8887);
nor UO_66 (O_66,N_9577,N_9920);
or UO_67 (O_67,N_9894,N_9887);
and UO_68 (O_68,N_9339,N_9024);
nor UO_69 (O_69,N_8021,N_9341);
nand UO_70 (O_70,N_8289,N_9797);
or UO_71 (O_71,N_8955,N_9888);
or UO_72 (O_72,N_9741,N_8288);
or UO_73 (O_73,N_8528,N_8567);
and UO_74 (O_74,N_8124,N_8902);
nor UO_75 (O_75,N_9970,N_7632);
or UO_76 (O_76,N_7639,N_9303);
or UO_77 (O_77,N_7865,N_8164);
nand UO_78 (O_78,N_8800,N_9353);
and UO_79 (O_79,N_9752,N_9927);
nand UO_80 (O_80,N_7544,N_8283);
nor UO_81 (O_81,N_8183,N_9053);
nand UO_82 (O_82,N_9135,N_7568);
and UO_83 (O_83,N_8750,N_9338);
and UO_84 (O_84,N_9181,N_9385);
and UO_85 (O_85,N_9237,N_8123);
nand UO_86 (O_86,N_9394,N_8443);
nor UO_87 (O_87,N_7536,N_7957);
nand UO_88 (O_88,N_9580,N_9791);
and UO_89 (O_89,N_9250,N_9030);
nor UO_90 (O_90,N_8533,N_9881);
or UO_91 (O_91,N_8331,N_7813);
or UO_92 (O_92,N_7522,N_8071);
or UO_93 (O_93,N_8386,N_9510);
nand UO_94 (O_94,N_7675,N_7601);
nand UO_95 (O_95,N_7557,N_7612);
or UO_96 (O_96,N_9273,N_8763);
nand UO_97 (O_97,N_8287,N_8357);
nor UO_98 (O_98,N_7771,N_9781);
nand UO_99 (O_99,N_7864,N_9568);
nand UO_100 (O_100,N_9660,N_8811);
xnor UO_101 (O_101,N_7727,N_8001);
or UO_102 (O_102,N_9634,N_8918);
and UO_103 (O_103,N_8261,N_7546);
nand UO_104 (O_104,N_7631,N_8595);
nor UO_105 (O_105,N_7885,N_8521);
nand UO_106 (O_106,N_8873,N_8799);
nand UO_107 (O_107,N_9414,N_9555);
or UO_108 (O_108,N_8620,N_8039);
or UO_109 (O_109,N_8680,N_7517);
nor UO_110 (O_110,N_9993,N_7983);
or UO_111 (O_111,N_8053,N_7654);
and UO_112 (O_112,N_9316,N_9081);
nor UO_113 (O_113,N_9012,N_7897);
nand UO_114 (O_114,N_9236,N_8900);
nor UO_115 (O_115,N_8360,N_7628);
and UO_116 (O_116,N_8648,N_8532);
nand UO_117 (O_117,N_8824,N_7689);
nand UO_118 (O_118,N_7737,N_9331);
nor UO_119 (O_119,N_7593,N_9551);
nor UO_120 (O_120,N_8094,N_7978);
nand UO_121 (O_121,N_8141,N_8281);
nand UO_122 (O_122,N_8655,N_7846);
or UO_123 (O_123,N_8260,N_8976);
nand UO_124 (O_124,N_9779,N_8768);
nor UO_125 (O_125,N_7746,N_9091);
nand UO_126 (O_126,N_8993,N_7784);
and UO_127 (O_127,N_9256,N_8547);
xnor UO_128 (O_128,N_9554,N_8158);
nor UO_129 (O_129,N_9732,N_9966);
or UO_130 (O_130,N_9479,N_7567);
nand UO_131 (O_131,N_7573,N_9532);
nor UO_132 (O_132,N_9189,N_9854);
xor UO_133 (O_133,N_7788,N_7624);
nor UO_134 (O_134,N_9429,N_8554);
nand UO_135 (O_135,N_8250,N_9988);
or UO_136 (O_136,N_9020,N_9528);
and UO_137 (O_137,N_8947,N_8014);
nand UO_138 (O_138,N_9664,N_8495);
or UO_139 (O_139,N_7979,N_8453);
nor UO_140 (O_140,N_9842,N_7898);
and UO_141 (O_141,N_8235,N_9957);
or UO_142 (O_142,N_9611,N_8734);
or UO_143 (O_143,N_7986,N_8971);
nand UO_144 (O_144,N_9929,N_9088);
nand UO_145 (O_145,N_9573,N_9018);
nor UO_146 (O_146,N_9272,N_9460);
or UO_147 (O_147,N_9217,N_7977);
nor UO_148 (O_148,N_9214,N_9262);
nor UO_149 (O_149,N_9754,N_9398);
or UO_150 (O_150,N_8546,N_9507);
or UO_151 (O_151,N_8147,N_7694);
and UO_152 (O_152,N_9424,N_8929);
nand UO_153 (O_153,N_8975,N_7611);
and UO_154 (O_154,N_8173,N_8374);
and UO_155 (O_155,N_8390,N_8458);
nand UO_156 (O_156,N_9641,N_9847);
nand UO_157 (O_157,N_8980,N_8307);
and UO_158 (O_158,N_8432,N_9282);
and UO_159 (O_159,N_9128,N_8407);
nand UO_160 (O_160,N_9982,N_9198);
or UO_161 (O_161,N_9065,N_9219);
xnor UO_162 (O_162,N_9359,N_9959);
nor UO_163 (O_163,N_9963,N_9351);
or UO_164 (O_164,N_9814,N_8990);
or UO_165 (O_165,N_9073,N_8512);
or UO_166 (O_166,N_8275,N_8499);
and UO_167 (O_167,N_9407,N_9221);
nor UO_168 (O_168,N_7534,N_9861);
or UO_169 (O_169,N_8593,N_8258);
nor UO_170 (O_170,N_9945,N_8191);
nand UO_171 (O_171,N_9231,N_9734);
nor UO_172 (O_172,N_8408,N_7699);
nor UO_173 (O_173,N_8560,N_9983);
nand UO_174 (O_174,N_9816,N_8842);
or UO_175 (O_175,N_8237,N_8912);
nor UO_176 (O_176,N_8490,N_9491);
nor UO_177 (O_177,N_8318,N_8397);
or UO_178 (O_178,N_8154,N_8782);
nor UO_179 (O_179,N_8540,N_8217);
and UO_180 (O_180,N_7946,N_9824);
nor UO_181 (O_181,N_8069,N_7733);
and UO_182 (O_182,N_8212,N_8923);
nor UO_183 (O_183,N_8704,N_9013);
or UO_184 (O_184,N_8373,N_8810);
nand UO_185 (O_185,N_8911,N_8840);
nand UO_186 (O_186,N_9283,N_9432);
nand UO_187 (O_187,N_9788,N_8330);
or UO_188 (O_188,N_8379,N_8519);
or UO_189 (O_189,N_8203,N_9731);
nor UO_190 (O_190,N_9939,N_8145);
or UO_191 (O_191,N_8774,N_9179);
nor UO_192 (O_192,N_8688,N_8338);
and UO_193 (O_193,N_8803,N_9378);
and UO_194 (O_194,N_8370,N_9994);
nor UO_195 (O_195,N_7795,N_9737);
or UO_196 (O_196,N_9897,N_9293);
nand UO_197 (O_197,N_9114,N_7829);
or UO_198 (O_198,N_9632,N_8451);
and UO_199 (O_199,N_8625,N_9936);
nand UO_200 (O_200,N_9785,N_8433);
or UO_201 (O_201,N_8962,N_7687);
or UO_202 (O_202,N_8199,N_8454);
and UO_203 (O_203,N_8413,N_9315);
nand UO_204 (O_204,N_7893,N_9416);
and UO_205 (O_205,N_9800,N_8737);
xor UO_206 (O_206,N_7981,N_8111);
or UO_207 (O_207,N_8713,N_7756);
or UO_208 (O_208,N_8755,N_9248);
and UO_209 (O_209,N_8116,N_9213);
xor UO_210 (O_210,N_8589,N_7778);
nor UO_211 (O_211,N_9365,N_9396);
and UO_212 (O_212,N_9220,N_7518);
xor UO_213 (O_213,N_8707,N_7598);
and UO_214 (O_214,N_9813,N_8205);
and UO_215 (O_215,N_9622,N_9155);
nor UO_216 (O_216,N_8468,N_9669);
nand UO_217 (O_217,N_9387,N_9765);
and UO_218 (O_218,N_7899,N_9952);
nor UO_219 (O_219,N_7594,N_8204);
and UO_220 (O_220,N_9287,N_7591);
nor UO_221 (O_221,N_8162,N_9074);
and UO_222 (O_222,N_8293,N_9834);
nor UO_223 (O_223,N_9638,N_9404);
nand UO_224 (O_224,N_8575,N_7740);
nor UO_225 (O_225,N_9399,N_8874);
nand UO_226 (O_226,N_8114,N_9848);
nor UO_227 (O_227,N_9629,N_8034);
or UO_228 (O_228,N_7511,N_7831);
or UO_229 (O_229,N_8741,N_8228);
or UO_230 (O_230,N_8482,N_9601);
and UO_231 (O_231,N_9623,N_9523);
xor UO_232 (O_232,N_7692,N_9827);
xor UO_233 (O_233,N_7585,N_7571);
and UO_234 (O_234,N_8711,N_7637);
and UO_235 (O_235,N_9613,N_8571);
and UO_236 (O_236,N_9149,N_9830);
nor UO_237 (O_237,N_8229,N_8876);
nand UO_238 (O_238,N_9410,N_9599);
nand UO_239 (O_239,N_8525,N_8752);
nand UO_240 (O_240,N_8983,N_7682);
or UO_241 (O_241,N_8999,N_8029);
or UO_242 (O_242,N_7630,N_8278);
or UO_243 (O_243,N_8050,N_8957);
nand UO_244 (O_244,N_8871,N_9537);
and UO_245 (O_245,N_8155,N_7589);
and UO_246 (O_246,N_7886,N_7558);
or UO_247 (O_247,N_9166,N_9954);
nor UO_248 (O_248,N_7857,N_8328);
or UO_249 (O_249,N_7866,N_8159);
nor UO_250 (O_250,N_9776,N_9152);
nand UO_251 (O_251,N_8831,N_8273);
or UO_252 (O_252,N_9140,N_7933);
nor UO_253 (O_253,N_8766,N_9518);
or UO_254 (O_254,N_8078,N_9932);
nor UO_255 (O_255,N_7608,N_7712);
nand UO_256 (O_256,N_9631,N_9045);
nand UO_257 (O_257,N_9987,N_9645);
nor UO_258 (O_258,N_9326,N_8368);
and UO_259 (O_259,N_8643,N_8455);
and UO_260 (O_260,N_9126,N_8506);
xor UO_261 (O_261,N_9984,N_7583);
and UO_262 (O_262,N_9105,N_9471);
nor UO_263 (O_263,N_9862,N_9676);
or UO_264 (O_264,N_8066,N_7906);
nand UO_265 (O_265,N_8269,N_9259);
xor UO_266 (O_266,N_9775,N_7599);
nor UO_267 (O_267,N_7707,N_9478);
nand UO_268 (O_268,N_8500,N_8665);
nor UO_269 (O_269,N_8296,N_9131);
and UO_270 (O_270,N_8700,N_7781);
xor UO_271 (O_271,N_8684,N_9475);
xnor UO_272 (O_272,N_8294,N_7776);
nor UO_273 (O_273,N_9098,N_9517);
and UO_274 (O_274,N_9112,N_8290);
xnor UO_275 (O_275,N_8234,N_7919);
or UO_276 (O_276,N_8182,N_9176);
nand UO_277 (O_277,N_9992,N_9600);
nor UO_278 (O_278,N_7786,N_8343);
and UO_279 (O_279,N_9699,N_9560);
nor UO_280 (O_280,N_9072,N_7703);
nand UO_281 (O_281,N_9519,N_9925);
nor UO_282 (O_282,N_8781,N_9609);
and UO_283 (O_283,N_8862,N_9484);
nand UO_284 (O_284,N_7650,N_9142);
or UO_285 (O_285,N_9962,N_8138);
nand UO_286 (O_286,N_9969,N_7805);
nand UO_287 (O_287,N_8697,N_7993);
xor UO_288 (O_288,N_7763,N_8808);
xnor UO_289 (O_289,N_8177,N_9043);
or UO_290 (O_290,N_9704,N_9868);
or UO_291 (O_291,N_7758,N_8714);
or UO_292 (O_292,N_9245,N_9034);
and UO_293 (O_293,N_7980,N_9647);
or UO_294 (O_294,N_8364,N_7790);
or UO_295 (O_295,N_9646,N_9505);
nand UO_296 (O_296,N_9102,N_9810);
or UO_297 (O_297,N_8435,N_8724);
nand UO_298 (O_298,N_8475,N_8965);
nor UO_299 (O_299,N_9055,N_9464);
xor UO_300 (O_300,N_9735,N_8534);
nor UO_301 (O_301,N_8098,N_9292);
or UO_302 (O_302,N_7876,N_8622);
nand UO_303 (O_303,N_9335,N_9358);
or UO_304 (O_304,N_8812,N_8042);
and UO_305 (O_305,N_8464,N_8645);
and UO_306 (O_306,N_9085,N_8543);
nand UO_307 (O_307,N_7739,N_8779);
nor UO_308 (O_308,N_9130,N_9291);
nor UO_309 (O_309,N_7798,N_7691);
nor UO_310 (O_310,N_9572,N_9559);
xor UO_311 (O_311,N_8646,N_8847);
nor UO_312 (O_312,N_9923,N_7814);
and UO_313 (O_313,N_7658,N_8195);
nor UO_314 (O_314,N_7747,N_8002);
nand UO_315 (O_315,N_8516,N_8012);
and UO_316 (O_316,N_9990,N_9199);
or UO_317 (O_317,N_8469,N_9186);
and UO_318 (O_318,N_9047,N_7997);
and UO_319 (O_319,N_7730,N_8246);
nand UO_320 (O_320,N_9270,N_8356);
nor UO_321 (O_321,N_9336,N_7974);
nor UO_322 (O_322,N_8376,N_7958);
nor UO_323 (O_323,N_9406,N_8857);
nand UO_324 (O_324,N_7705,N_9314);
nand UO_325 (O_325,N_9783,N_8339);
or UO_326 (O_326,N_9500,N_8522);
and UO_327 (O_327,N_7762,N_9652);
nor UO_328 (O_328,N_9493,N_8712);
nor UO_329 (O_329,N_8075,N_7913);
and UO_330 (O_330,N_8074,N_9007);
nor UO_331 (O_331,N_9721,N_9408);
or UO_332 (O_332,N_8101,N_7540);
and UO_333 (O_333,N_8485,N_7570);
xor UO_334 (O_334,N_8604,N_8438);
or UO_335 (O_335,N_8349,N_9026);
nand UO_336 (O_336,N_8562,N_7500);
nand UO_337 (O_337,N_9882,N_8216);
or UO_338 (O_338,N_9360,N_8610);
nand UO_339 (O_339,N_9692,N_8897);
nand UO_340 (O_340,N_9960,N_8148);
nand UO_341 (O_341,N_9892,N_8987);
nand UO_342 (O_342,N_8285,N_8441);
and UO_343 (O_343,N_8647,N_8206);
nand UO_344 (O_344,N_9222,N_8491);
and UO_345 (O_345,N_9789,N_7872);
nor UO_346 (O_346,N_9107,N_7751);
or UO_347 (O_347,N_9477,N_7519);
or UO_348 (O_348,N_8970,N_9879);
nand UO_349 (O_349,N_9758,N_8227);
and UO_350 (O_350,N_7515,N_9017);
or UO_351 (O_351,N_9210,N_8215);
and UO_352 (O_352,N_7738,N_8641);
and UO_353 (O_353,N_8313,N_9150);
and UO_354 (O_354,N_7863,N_8207);
and UO_355 (O_355,N_8686,N_7904);
nor UO_356 (O_356,N_9736,N_8334);
nor UO_357 (O_357,N_7734,N_9548);
or UO_358 (O_358,N_8118,N_9440);
or UO_359 (O_359,N_8557,N_8346);
and UO_360 (O_360,N_8030,N_8056);
and UO_361 (O_361,N_8673,N_8232);
nand UO_362 (O_362,N_8907,N_8813);
nand UO_363 (O_363,N_9252,N_7665);
nor UO_364 (O_364,N_8966,N_9768);
nor UO_365 (O_365,N_8925,N_9106);
nand UO_366 (O_366,N_7950,N_7888);
nor UO_367 (O_367,N_9831,N_9565);
or UO_368 (O_368,N_9856,N_7701);
nand UO_369 (O_369,N_8927,N_8105);
nor UO_370 (O_370,N_8583,N_9042);
or UO_371 (O_371,N_9031,N_8406);
nand UO_372 (O_372,N_9151,N_8309);
and UO_373 (O_373,N_8662,N_8514);
and UO_374 (O_374,N_7547,N_9713);
nand UO_375 (O_375,N_9172,N_7532);
or UO_376 (O_376,N_8504,N_7706);
nand UO_377 (O_377,N_8063,N_7635);
nor UO_378 (O_378,N_8517,N_9743);
and UO_379 (O_379,N_9465,N_8398);
nand UO_380 (O_380,N_9938,N_8559);
nor UO_381 (O_381,N_8426,N_7741);
or UO_382 (O_382,N_7660,N_8624);
and UO_383 (O_383,N_9100,N_8650);
nand UO_384 (O_384,N_9267,N_8302);
nand UO_385 (O_385,N_8669,N_9742);
or UO_386 (O_386,N_9610,N_7556);
nor UO_387 (O_387,N_9707,N_7900);
and UO_388 (O_388,N_9684,N_8565);
and UO_389 (O_389,N_8992,N_7538);
nand UO_390 (O_390,N_9832,N_9288);
nand UO_391 (O_391,N_7604,N_7504);
nor UO_392 (O_392,N_9701,N_8563);
nor UO_393 (O_393,N_9027,N_7620);
or UO_394 (O_394,N_9639,N_8577);
and UO_395 (O_395,N_8561,N_9371);
and UO_396 (O_396,N_9340,N_8825);
xnor UO_397 (O_397,N_7816,N_8152);
or UO_398 (O_398,N_8961,N_9921);
nor UO_399 (O_399,N_8898,N_9853);
nor UO_400 (O_400,N_8915,N_9224);
and UO_401 (O_401,N_9968,N_8007);
and UO_402 (O_402,N_8938,N_8047);
xnor UO_403 (O_403,N_7901,N_9913);
nand UO_404 (O_404,N_8544,N_7673);
nor UO_405 (O_405,N_7760,N_8502);
nor UO_406 (O_406,N_9986,N_9719);
nor UO_407 (O_407,N_8423,N_8245);
nand UO_408 (O_408,N_9441,N_8715);
and UO_409 (O_409,N_9873,N_9474);
and UO_410 (O_410,N_8174,N_8744);
nand UO_411 (O_411,N_8299,N_9612);
nor UO_412 (O_412,N_9304,N_8421);
and UO_413 (O_413,N_9108,N_8187);
or UO_414 (O_414,N_8006,N_9354);
or UO_415 (O_415,N_9694,N_9476);
nand UO_416 (O_416,N_7525,N_8401);
and UO_417 (O_417,N_7808,N_9139);
nand UO_418 (O_418,N_9242,N_8783);
xnor UO_419 (O_419,N_8949,N_7552);
and UO_420 (O_420,N_9383,N_9490);
or UO_421 (O_421,N_9625,N_9413);
nor UO_422 (O_422,N_9722,N_8165);
nor UO_423 (O_423,N_9207,N_8564);
nand UO_424 (O_424,N_9616,N_7633);
nor UO_425 (O_425,N_7773,N_9307);
and UO_426 (O_426,N_7819,N_8459);
nor UO_427 (O_427,N_9885,N_8045);
or UO_428 (O_428,N_9971,N_7939);
and UO_429 (O_429,N_9356,N_9972);
and UO_430 (O_430,N_9313,N_8969);
nand UO_431 (O_431,N_7891,N_8144);
and UO_432 (O_432,N_7956,N_9253);
and UO_433 (O_433,N_9730,N_7775);
nand UO_434 (O_434,N_8951,N_9635);
or UO_435 (O_435,N_8102,N_8868);
nand UO_436 (O_436,N_9522,N_9361);
nand UO_437 (O_437,N_8638,N_8478);
nor UO_438 (O_438,N_7642,N_8016);
and UO_439 (O_439,N_8329,N_9261);
and UO_440 (O_440,N_9956,N_7543);
nand UO_441 (O_441,N_9912,N_9003);
or UO_442 (O_442,N_9060,N_8640);
nand UO_443 (O_443,N_7649,N_8498);
or UO_444 (O_444,N_9317,N_9666);
nand UO_445 (O_445,N_9431,N_7595);
and UO_446 (O_446,N_8427,N_9372);
or UO_447 (O_447,N_8706,N_9321);
nand UO_448 (O_448,N_8815,N_9605);
and UO_449 (O_449,N_7840,N_7791);
or UO_450 (O_450,N_9680,N_8717);
or UO_451 (O_451,N_8851,N_8526);
or UO_452 (O_452,N_7996,N_9521);
or UO_453 (O_453,N_9591,N_8201);
and UO_454 (O_454,N_9393,N_9534);
or UO_455 (O_455,N_8383,N_9583);
and UO_456 (O_456,N_9193,N_7729);
and UO_457 (O_457,N_8991,N_7584);
nand UO_458 (O_458,N_7938,N_8308);
or UO_459 (O_459,N_8657,N_8391);
nand UO_460 (O_460,N_9667,N_9458);
nand UO_461 (O_461,N_7607,N_9643);
nand UO_462 (O_462,N_9101,N_9376);
or UO_463 (O_463,N_7723,N_9298);
and UO_464 (O_464,N_9422,N_7923);
nor UO_465 (O_465,N_8146,N_9553);
nand UO_466 (O_466,N_8086,N_8209);
or UO_467 (O_467,N_8168,N_7721);
nor UO_468 (O_468,N_7680,N_7847);
nor UO_469 (O_469,N_9900,N_8160);
and UO_470 (O_470,N_8586,N_7693);
nor UO_471 (O_471,N_8409,N_7926);
nor UO_472 (O_472,N_8696,N_7810);
xnor UO_473 (O_473,N_8835,N_9289);
or UO_474 (O_474,N_7622,N_8150);
nand UO_475 (O_475,N_8026,N_9801);
nand UO_476 (O_476,N_8266,N_7686);
nand UO_477 (O_477,N_9545,N_7672);
or UO_478 (O_478,N_9125,N_9295);
and UO_479 (O_479,N_8865,N_9305);
or UO_480 (O_480,N_9450,N_9374);
and UO_481 (O_481,N_8493,N_9835);
and UO_482 (O_482,N_8262,N_9071);
nor UO_483 (O_483,N_8248,N_9312);
and UO_484 (O_484,N_8186,N_8916);
nand UO_485 (O_485,N_9628,N_9447);
nor UO_486 (O_486,N_9782,N_7875);
nor UO_487 (O_487,N_8972,N_9296);
or UO_488 (O_488,N_9197,N_8973);
nor UO_489 (O_489,N_8530,N_9244);
nand UO_490 (O_490,N_7731,N_7768);
nand UO_491 (O_491,N_9482,N_9168);
and UO_492 (O_492,N_8351,N_9849);
nand UO_493 (O_493,N_9651,N_7566);
nor UO_494 (O_494,N_7569,N_9136);
nand UO_495 (O_495,N_9865,N_7647);
and UO_496 (O_496,N_7815,N_9526);
nand UO_497 (O_497,N_7964,N_9541);
nand UO_498 (O_498,N_9826,N_9454);
or UO_499 (O_499,N_9035,N_7580);
nor UO_500 (O_500,N_9025,N_8581);
nand UO_501 (O_501,N_7728,N_8369);
and UO_502 (O_502,N_7735,N_7625);
or UO_503 (O_503,N_9837,N_9530);
nand UO_504 (O_504,N_9792,N_8292);
or UO_505 (O_505,N_9710,N_9095);
or UO_506 (O_506,N_9615,N_8621);
or UO_507 (O_507,N_8910,N_7767);
or UO_508 (O_508,N_8085,N_8068);
and UO_509 (O_509,N_9756,N_9588);
nand UO_510 (O_510,N_9495,N_8837);
and UO_511 (O_511,N_8933,N_8080);
and UO_512 (O_512,N_8137,N_7972);
nand UO_513 (O_513,N_7999,N_9761);
nor UO_514 (O_514,N_7529,N_7696);
or UO_515 (O_515,N_8214,N_7530);
or UO_516 (O_516,N_9434,N_8632);
nand UO_517 (O_517,N_8833,N_9089);
and UO_518 (O_518,N_8894,N_7765);
nor UO_519 (O_519,N_8089,N_9344);
and UO_520 (O_520,N_7925,N_7742);
xor UO_521 (O_521,N_7826,N_9512);
nand UO_522 (O_522,N_9808,N_7676);
nor UO_523 (O_523,N_9594,N_9485);
nand UO_524 (O_524,N_8855,N_7718);
nand UO_525 (O_525,N_7748,N_8310);
or UO_526 (O_526,N_8848,N_9010);
nand UO_527 (O_527,N_9582,N_7945);
nor UO_528 (O_528,N_7982,N_8072);
nor UO_529 (O_529,N_9506,N_9606);
and UO_530 (O_530,N_9996,N_9229);
and UO_531 (O_531,N_8425,N_9698);
or UO_532 (O_532,N_9182,N_9056);
nor UO_533 (O_533,N_9603,N_8465);
nor UO_534 (O_534,N_7975,N_9400);
and UO_535 (O_535,N_9196,N_8440);
and UO_536 (O_536,N_9636,N_7877);
nand UO_537 (O_537,N_7514,N_9536);
and UO_538 (O_538,N_9334,N_8960);
and UO_539 (O_539,N_8058,N_9247);
nand UO_540 (O_540,N_9790,N_7664);
and UO_541 (O_541,N_9708,N_8885);
or UO_542 (O_542,N_7685,N_8762);
and UO_543 (O_543,N_9794,N_9766);
or UO_544 (O_544,N_9068,N_9593);
nor UO_545 (O_545,N_9979,N_9818);
nor UO_546 (O_546,N_7678,N_9604);
nand UO_547 (O_547,N_9877,N_8479);
and UO_548 (O_548,N_9998,N_9943);
or UO_549 (O_549,N_8494,N_7581);
nand UO_550 (O_550,N_8342,N_9608);
or UO_551 (O_551,N_9211,N_9486);
and UO_552 (O_552,N_9702,N_9215);
or UO_553 (O_553,N_9755,N_8566);
nand UO_554 (O_554,N_9578,N_9891);
or UO_555 (O_555,N_7955,N_8109);
and UO_556 (O_556,N_8904,N_9700);
nand UO_557 (O_557,N_9753,N_8185);
and UO_558 (O_558,N_9350,N_7934);
and UO_559 (O_559,N_9965,N_8377);
nand UO_560 (O_560,N_8558,N_7817);
nand UO_561 (O_561,N_8236,N_8314);
or UO_562 (O_562,N_8198,N_8181);
or UO_563 (O_563,N_9621,N_8473);
or UO_564 (O_564,N_9899,N_9595);
or UO_565 (O_565,N_8040,N_7861);
nand UO_566 (O_566,N_9663,N_8325);
and UO_567 (O_567,N_7521,N_9596);
xor UO_568 (O_568,N_7614,N_7590);
or UO_569 (O_569,N_7634,N_8890);
or UO_570 (O_570,N_9675,N_9981);
xnor UO_571 (O_571,N_7834,N_8036);
nand UO_572 (O_572,N_8190,N_7531);
and UO_573 (O_573,N_7868,N_8130);
nand UO_574 (O_574,N_8765,N_9120);
or UO_575 (O_575,N_8213,N_8798);
nand UO_576 (O_576,N_9318,N_8428);
and UO_577 (O_577,N_8754,N_7732);
nand UO_578 (O_578,N_8693,N_9346);
nor UO_579 (O_579,N_9037,N_9391);
and UO_580 (O_580,N_9820,N_9254);
and UO_581 (O_581,N_7505,N_7821);
and UO_582 (O_582,N_7526,N_9036);
nand UO_583 (O_583,N_9084,N_9430);
nand UO_584 (O_584,N_9592,N_7651);
xnor UO_585 (O_585,N_7561,N_9403);
nor UO_586 (O_586,N_8612,N_9607);
or UO_587 (O_587,N_8431,N_7769);
and UO_588 (O_588,N_9570,N_8054);
and UO_589 (O_589,N_8541,N_9880);
and UO_590 (O_590,N_9911,N_8161);
nor UO_591 (O_591,N_8303,N_8096);
nand UO_592 (O_592,N_7848,N_7961);
nor UO_593 (O_593,N_8097,N_9524);
or UO_594 (O_594,N_9137,N_8448);
and UO_595 (O_595,N_9860,N_9347);
nand UO_596 (O_596,N_8508,N_8817);
nor UO_597 (O_597,N_7627,N_9798);
xnor UO_598 (O_598,N_8172,N_9421);
nand UO_599 (O_599,N_9342,N_9838);
or UO_600 (O_600,N_9529,N_9087);
nand UO_601 (O_601,N_7715,N_9953);
nand UO_602 (O_602,N_9218,N_8652);
and UO_603 (O_603,N_7550,N_9822);
or UO_604 (O_604,N_8913,N_7736);
and UO_605 (O_605,N_7711,N_9274);
nand UO_606 (O_606,N_7683,N_7600);
nand UO_607 (O_607,N_8503,N_9076);
nor UO_608 (O_608,N_8675,N_9703);
nor UO_609 (O_609,N_7914,N_9901);
and UO_610 (O_610,N_9212,N_8928);
or UO_611 (O_611,N_7623,N_7969);
nor UO_612 (O_612,N_9681,N_9863);
and UO_613 (O_613,N_8689,N_7867);
and UO_614 (O_614,N_7804,N_8211);
nand UO_615 (O_615,N_9438,N_9062);
nor UO_616 (O_616,N_7613,N_7827);
or UO_617 (O_617,N_9241,N_7907);
and UO_618 (O_618,N_8764,N_9670);
nor UO_619 (O_619,N_8613,N_8654);
or UO_620 (O_620,N_7912,N_9499);
or UO_621 (O_621,N_8359,N_8467);
nand UO_622 (O_622,N_8125,N_9038);
nand UO_623 (O_623,N_9094,N_8319);
nand UO_624 (O_624,N_9738,N_9169);
nor UO_625 (O_625,N_7998,N_7792);
nand UO_626 (O_626,N_7725,N_8122);
nand UO_627 (O_627,N_7757,N_8139);
or UO_628 (O_628,N_8549,N_8194);
or UO_629 (O_629,N_8119,N_9330);
nand UO_630 (O_630,N_9175,N_9271);
or UO_631 (O_631,N_8527,N_8456);
and UO_632 (O_632,N_9771,N_7779);
or UO_633 (O_633,N_8282,N_9620);
nand UO_634 (O_634,N_9928,N_8796);
nor UO_635 (O_635,N_8019,N_8834);
nor UO_636 (O_636,N_7895,N_9581);
nand UO_637 (O_637,N_9557,N_8930);
or UO_638 (O_638,N_9451,N_8832);
and UO_639 (O_639,N_8179,N_8450);
and UO_640 (O_640,N_8742,N_8412);
nor UO_641 (O_641,N_8677,N_7843);
or UO_642 (O_642,N_7555,N_9930);
and UO_643 (O_643,N_9415,N_9352);
nand UO_644 (O_644,N_7917,N_7794);
nor UO_645 (O_645,N_8598,N_9205);
nor UO_646 (O_646,N_9805,N_7743);
and UO_647 (O_647,N_7818,N_8341);
and UO_648 (O_648,N_8520,N_9672);
nand UO_649 (O_649,N_9696,N_8027);
nand UO_650 (O_650,N_9144,N_7873);
and UO_651 (O_651,N_8816,N_9370);
nand UO_652 (O_652,N_9948,N_8396);
nand UO_653 (O_653,N_7811,N_7761);
nor UO_654 (O_654,N_9774,N_8415);
nor UO_655 (O_655,N_8515,N_9226);
nor UO_656 (O_656,N_8974,N_8434);
and UO_657 (O_657,N_9656,N_7782);
xor UO_658 (O_658,N_7645,N_8257);
and UO_659 (O_659,N_9974,N_9846);
nor UO_660 (O_660,N_7971,N_9748);
nor UO_661 (O_661,N_9784,N_8032);
nor UO_662 (O_662,N_9841,N_7941);
nor UO_663 (O_663,N_9263,N_7542);
nand UO_664 (O_664,N_9297,N_8208);
and UO_665 (O_665,N_9000,N_9185);
nor UO_666 (O_666,N_8015,N_8668);
nand UO_667 (O_667,N_8786,N_7507);
and UO_668 (O_668,N_7690,N_9893);
nor UO_669 (O_669,N_7659,N_9955);
xor UO_670 (O_670,N_9552,N_8010);
or UO_671 (O_671,N_8430,N_8748);
or UO_672 (O_672,N_8311,N_9724);
nor UO_673 (O_673,N_8671,N_9281);
xor UO_674 (O_674,N_7874,N_7657);
nand UO_675 (O_675,N_7588,N_8889);
or UO_676 (O_676,N_8753,N_8133);
or UO_677 (O_677,N_8239,N_7516);
nor UO_678 (O_678,N_9417,N_8322);
and UO_679 (O_679,N_9067,N_8025);
nor UO_680 (O_680,N_9437,N_8404);
nor UO_681 (O_681,N_8585,N_8989);
or UO_682 (O_682,N_8393,N_9022);
nor UO_683 (O_683,N_8941,N_7745);
or UO_684 (O_684,N_9803,N_7789);
and UO_685 (O_685,N_8363,N_8474);
xor UO_686 (O_686,N_9951,N_9129);
or UO_687 (O_687,N_9843,N_9069);
nor UO_688 (O_688,N_9368,N_8131);
nand UO_689 (O_689,N_9695,N_8320);
nand UO_690 (O_690,N_9118,N_8631);
nor UO_691 (O_691,N_8510,N_8606);
or UO_692 (O_692,N_7970,N_8576);
and UO_693 (O_693,N_8555,N_8088);
and UO_694 (O_694,N_8087,N_9531);
or UO_695 (O_695,N_7860,N_8863);
and UO_696 (O_696,N_8156,N_7508);
and UO_697 (O_697,N_9051,N_8590);
nand UO_698 (O_698,N_8127,N_7545);
or UO_699 (O_699,N_7677,N_9871);
or UO_700 (O_700,N_9673,N_9423);
nor UO_701 (O_701,N_8304,N_8954);
and UO_702 (O_702,N_9693,N_8226);
nand UO_703 (O_703,N_8169,N_8247);
xnor UO_704 (O_704,N_8681,N_9558);
nor UO_705 (O_705,N_8568,N_7749);
nor UO_706 (O_706,N_9944,N_9858);
and UO_707 (O_707,N_9160,N_9712);
and UO_708 (O_708,N_9011,N_8791);
nor UO_709 (O_709,N_8197,N_7992);
nand UO_710 (O_710,N_8616,N_8252);
and UO_711 (O_711,N_8830,N_9280);
nor UO_712 (O_712,N_9373,N_8104);
and UO_713 (O_713,N_8667,N_8129);
or UO_714 (O_714,N_9306,N_9549);
or UO_715 (O_715,N_8241,N_8740);
nand UO_716 (O_716,N_9171,N_8703);
nor UO_717 (O_717,N_8958,N_7881);
or UO_718 (O_718,N_8805,N_7839);
nor UO_719 (O_719,N_7951,N_9671);
or UO_720 (O_720,N_8013,N_9501);
and UO_721 (O_721,N_9566,N_7838);
and UO_722 (O_722,N_9799,N_9749);
and UO_723 (O_723,N_9527,N_9898);
and UO_724 (O_724,N_8090,N_9919);
nand UO_725 (O_725,N_7988,N_8708);
nor UO_726 (O_726,N_8905,N_9349);
or UO_727 (O_727,N_9989,N_8998);
nand UO_728 (O_728,N_8690,N_8009);
nor UO_729 (O_729,N_8128,N_9469);
or UO_730 (O_730,N_8718,N_8858);
or UO_731 (O_731,N_9153,N_9855);
and UO_732 (O_732,N_9054,N_8348);
or UO_733 (O_733,N_7770,N_8823);
nand UO_734 (O_734,N_7793,N_8084);
or UO_735 (O_735,N_8920,N_8518);
xor UO_736 (O_736,N_9890,N_8759);
nand UO_737 (O_737,N_8749,N_9999);
nand UO_738 (O_738,N_8410,N_8804);
or UO_739 (O_739,N_8679,N_9494);
nor UO_740 (O_740,N_9682,N_9392);
and UO_741 (O_741,N_9324,N_8402);
or UO_742 (O_742,N_8634,N_8188);
nand UO_743 (O_743,N_9462,N_8489);
or UO_744 (O_744,N_7937,N_8225);
nor UO_745 (O_745,N_9048,N_9683);
and UO_746 (O_746,N_7908,N_7890);
nor UO_747 (O_747,N_9367,N_8277);
or UO_748 (O_748,N_8306,N_8044);
nand UO_749 (O_749,N_9780,N_9985);
nand UO_750 (O_750,N_8300,N_9567);
nand UO_751 (O_751,N_8035,N_8249);
nand UO_752 (O_752,N_8483,N_9191);
and UO_753 (O_753,N_8184,N_8264);
or UO_754 (O_754,N_8760,N_8117);
and UO_755 (O_755,N_8611,N_8446);
nor UO_756 (O_756,N_9561,N_8166);
and UO_757 (O_757,N_8419,N_9489);
or UO_758 (O_758,N_7916,N_9389);
and UO_759 (O_759,N_9812,N_9579);
nor UO_760 (O_760,N_9225,N_9204);
xnor UO_761 (O_761,N_8268,N_9503);
and UO_762 (O_762,N_9234,N_9109);
and UO_763 (O_763,N_7533,N_8210);
nand UO_764 (O_764,N_8952,N_7603);
or UO_765 (O_765,N_8956,N_9246);
and UO_766 (O_766,N_9688,N_9285);
or UO_767 (O_767,N_9302,N_9362);
or UO_768 (O_768,N_7952,N_8347);
nand UO_769 (O_769,N_8103,N_7841);
or UO_770 (O_770,N_9070,N_9311);
and UO_771 (O_771,N_7856,N_9864);
nand UO_772 (O_772,N_8827,N_8223);
nand UO_773 (O_773,N_9511,N_8552);
and UO_774 (O_774,N_9819,N_9427);
and UO_775 (O_775,N_9795,N_7506);
or UO_776 (O_776,N_9914,N_9903);
nor UO_777 (O_777,N_8607,N_9266);
nand UO_778 (O_778,N_8636,N_9239);
nand UO_779 (O_779,N_9844,N_8253);
nor UO_780 (O_780,N_8600,N_8644);
nor UO_781 (O_781,N_8859,N_7910);
nor UO_782 (O_782,N_9916,N_8051);
nor UO_783 (O_783,N_8787,N_8924);
nand UO_784 (O_784,N_9976,N_8591);
nand UO_785 (O_785,N_9733,N_8224);
nand UO_786 (O_786,N_8372,N_8535);
and UO_787 (O_787,N_7921,N_9886);
xor UO_788 (O_788,N_9975,N_8073);
nand UO_789 (O_789,N_7976,N_8676);
and UO_790 (O_790,N_8822,N_8332);
and UO_791 (O_791,N_9323,N_8460);
and UO_792 (O_792,N_8361,N_9472);
and UO_793 (O_793,N_9487,N_9804);
nor UO_794 (O_794,N_7859,N_9866);
and UO_795 (O_795,N_9991,N_8536);
nor UO_796 (O_796,N_8584,N_8112);
and UO_797 (O_797,N_8821,N_7991);
or UO_798 (O_798,N_9802,N_9760);
nor UO_799 (O_799,N_9064,N_8445);
nand UO_800 (O_800,N_8619,N_8064);
and UO_801 (O_801,N_7764,N_8943);
nand UO_802 (O_802,N_8829,N_9290);
or UO_803 (O_803,N_8937,N_9926);
or UO_804 (O_804,N_9815,N_7960);
and UO_805 (O_805,N_9412,N_9332);
or UO_806 (O_806,N_9420,N_7575);
and UO_807 (O_807,N_9809,N_9159);
nor UO_808 (O_808,N_9924,N_8321);
nor UO_809 (O_809,N_7671,N_8592);
and UO_810 (O_810,N_8442,N_8337);
nor UO_811 (O_811,N_8653,N_8470);
and UO_812 (O_812,N_9158,N_8022);
nand UO_813 (O_813,N_7889,N_9833);
or UO_814 (O_814,N_7799,N_8411);
or UO_815 (O_815,N_8860,N_8739);
and UO_816 (O_816,N_7909,N_9173);
and UO_817 (O_817,N_8614,N_9170);
nor UO_818 (O_818,N_7803,N_7714);
nand UO_819 (O_819,N_8853,N_7854);
and UO_820 (O_820,N_9678,N_8694);
and UO_821 (O_821,N_8157,N_7943);
nor UO_822 (O_822,N_9497,N_9057);
nand UO_823 (O_823,N_8509,N_9082);
or UO_824 (O_824,N_9269,N_8375);
or UO_825 (O_825,N_9299,N_8231);
nor UO_826 (O_826,N_7985,N_9584);
or UO_827 (O_827,N_9909,N_7564);
or UO_828 (O_828,N_7503,N_8843);
nor UO_829 (O_829,N_8336,N_8418);
nor UO_830 (O_830,N_9746,N_8852);
nand UO_831 (O_831,N_8323,N_9767);
nor UO_832 (O_832,N_8167,N_9111);
nand UO_833 (O_833,N_9585,N_7935);
or UO_834 (O_834,N_9277,N_9264);
nor UO_835 (O_835,N_9723,N_8795);
and UO_836 (O_836,N_9188,N_8507);
nor UO_837 (O_837,N_9147,N_7641);
or UO_838 (O_838,N_9874,N_9840);
or UO_839 (O_839,N_9384,N_9377);
nand UO_840 (O_840,N_7609,N_8597);
nor UO_841 (O_841,N_9598,N_9119);
or UO_842 (O_842,N_9845,N_7597);
nand UO_843 (O_843,N_9778,N_9395);
nor UO_844 (O_844,N_7722,N_7576);
or UO_845 (O_845,N_9857,N_8767);
nor UO_846 (O_846,N_7990,N_9015);
nor UO_847 (O_847,N_7963,N_9980);
or UO_848 (O_848,N_8335,N_7579);
nand UO_849 (O_849,N_7994,N_8240);
and UO_850 (O_850,N_8984,N_9910);
and UO_851 (O_851,N_9883,N_9902);
nor UO_852 (O_852,N_7510,N_9870);
nor UO_853 (O_853,N_9772,N_7560);
nand UO_854 (O_854,N_9397,N_8513);
and UO_855 (O_855,N_8219,N_7502);
nand UO_856 (O_856,N_9121,N_9569);
nand UO_857 (O_857,N_9851,N_9028);
nand UO_858 (O_858,N_7704,N_8772);
nor UO_859 (O_859,N_7894,N_7549);
and UO_860 (O_860,N_8274,N_8270);
or UO_861 (O_861,N_8466,N_9658);
or UO_862 (O_862,N_9544,N_8886);
nand UO_863 (O_863,N_9626,N_7527);
and UO_864 (O_864,N_9255,N_8439);
or UO_865 (O_865,N_9439,N_9044);
or UO_866 (O_866,N_8524,N_9964);
nand UO_867 (O_867,N_9077,N_8789);
nor UO_868 (O_868,N_8807,N_8609);
xor UO_869 (O_869,N_8149,N_9904);
and UO_870 (O_870,N_7824,N_8020);
or UO_871 (O_871,N_8775,N_7833);
nor UO_872 (O_872,N_8580,N_9203);
and UO_873 (O_873,N_8218,N_8276);
or UO_874 (O_874,N_8687,N_9745);
and UO_875 (O_875,N_8371,N_7942);
nand UO_876 (O_876,N_7574,N_8758);
or UO_877 (O_877,N_7936,N_8942);
and UO_878 (O_878,N_9807,N_7615);
or UO_879 (O_879,N_9947,N_8175);
and UO_880 (O_880,N_8382,N_9550);
and UO_881 (O_881,N_7572,N_9504);
nor UO_882 (O_882,N_9637,N_8921);
nand UO_883 (O_883,N_8171,N_9463);
and UO_884 (O_884,N_9040,N_8033);
and UO_885 (O_885,N_8556,N_9436);
nor UO_886 (O_886,N_9382,N_7924);
nor UO_887 (O_887,N_7610,N_7911);
or UO_888 (O_888,N_7902,N_8579);
nand UO_889 (O_889,N_9751,N_8344);
xnor UO_890 (O_890,N_8381,N_9099);
and UO_891 (O_891,N_9576,N_9828);
nand UO_892 (O_892,N_8284,N_8914);
and UO_893 (O_893,N_8950,N_7708);
nor UO_894 (O_894,N_9167,N_9426);
or UO_895 (O_895,N_7920,N_8745);
and UO_896 (O_896,N_8809,N_8076);
nor UO_897 (O_897,N_7626,N_8692);
nor UO_898 (O_898,N_9301,N_9941);
or UO_899 (O_899,N_8537,N_8618);
or UO_900 (O_900,N_9141,N_8899);
nand UO_901 (O_901,N_8553,N_8220);
nor UO_902 (O_902,N_7959,N_8082);
and UO_903 (O_903,N_8041,N_8698);
nor UO_904 (O_904,N_8389,N_9648);
or UO_905 (O_905,N_7619,N_9726);
or UO_906 (O_906,N_9061,N_9279);
nor UO_907 (O_907,N_9455,N_9540);
or UO_908 (O_908,N_8751,N_7666);
or UO_909 (O_909,N_8070,N_8539);
xor UO_910 (O_910,N_8005,N_7655);
nand UO_911 (O_911,N_8107,N_9445);
and UO_912 (O_912,N_8892,N_7915);
nand UO_913 (O_913,N_7717,N_8931);
nor UO_914 (O_914,N_9208,N_9777);
nor UO_915 (O_915,N_8801,N_8771);
nand UO_916 (O_916,N_8353,N_8488);
and UO_917 (O_917,N_8836,N_8747);
nor UO_918 (O_918,N_8221,N_9869);
nor UO_919 (O_919,N_7880,N_9029);
or UO_920 (O_920,N_8757,N_7845);
and UO_921 (O_921,N_9978,N_8477);
nor UO_922 (O_922,N_9322,N_8024);
nand UO_923 (O_923,N_9908,N_9668);
and UO_924 (O_924,N_8633,N_9161);
or UO_925 (O_925,N_7953,N_8664);
nor UO_926 (O_926,N_9542,N_9275);
and UO_927 (O_927,N_9258,N_9496);
or UO_928 (O_928,N_8945,N_9364);
or UO_929 (O_929,N_9649,N_9515);
nand UO_930 (O_930,N_7553,N_9618);
or UO_931 (O_931,N_7577,N_8617);
or UO_932 (O_932,N_8678,N_8770);
or UO_933 (O_933,N_9032,N_8922);
or UO_934 (O_934,N_8981,N_8746);
and UO_935 (O_935,N_8151,N_8891);
or UO_936 (O_936,N_9895,N_9190);
nand UO_937 (O_937,N_8656,N_9206);
nor UO_938 (O_938,N_9345,N_8701);
xor UO_939 (O_939,N_7931,N_8437);
nor UO_940 (O_940,N_8365,N_9575);
and UO_941 (O_941,N_8642,N_9564);
nand UO_942 (O_942,N_8896,N_9492);
or UO_943 (O_943,N_8254,N_8849);
nand UO_944 (O_944,N_8721,N_9442);
or UO_945 (O_945,N_8839,N_8878);
nand UO_946 (O_946,N_9706,N_8378);
and UO_947 (O_947,N_9456,N_8099);
nor UO_948 (O_948,N_9148,N_9728);
or UO_949 (O_949,N_8736,N_8903);
nor UO_950 (O_950,N_8846,N_8399);
nand UO_951 (O_951,N_9162,N_7855);
nor UO_952 (O_952,N_8301,N_7695);
or UO_953 (O_953,N_8523,N_9498);
or UO_954 (O_954,N_9744,N_8630);
nand UO_955 (O_955,N_7578,N_8492);
nand UO_956 (O_956,N_8472,N_8926);
and UO_957 (O_957,N_8735,N_9764);
or UO_958 (O_958,N_9829,N_9079);
nor UO_959 (O_959,N_9655,N_8594);
nor UO_960 (O_960,N_8004,N_7720);
nand UO_961 (O_961,N_9850,N_9058);
nand UO_962 (O_962,N_8092,N_9627);
nor UO_963 (O_963,N_8985,N_8777);
and UO_964 (O_964,N_8106,N_9714);
nor UO_965 (O_965,N_8877,N_9375);
or UO_966 (O_966,N_7850,N_7879);
and UO_967 (O_967,N_7513,N_9661);
nor UO_968 (O_968,N_8178,N_8997);
nand UO_969 (O_969,N_8599,N_8649);
xnor UO_970 (O_970,N_8233,N_9769);
nand UO_971 (O_971,N_7541,N_7922);
nor UO_972 (O_972,N_8542,N_8538);
and UO_973 (O_973,N_9092,N_8447);
and UO_974 (O_974,N_8267,N_9233);
and UO_975 (O_975,N_7962,N_9859);
and UO_976 (O_976,N_8728,N_9718);
and UO_977 (O_977,N_8864,N_7929);
xor UO_978 (O_978,N_9411,N_9878);
and UO_979 (O_979,N_7670,N_9195);
xnor UO_980 (O_980,N_8134,N_8940);
and UO_981 (O_981,N_9337,N_9390);
nor UO_982 (O_982,N_9896,N_8067);
or UO_983 (O_983,N_9640,N_9836);
or UO_984 (O_984,N_9630,N_9459);
nor UO_985 (O_985,N_8587,N_7858);
or UO_986 (O_986,N_8052,N_9653);
nand UO_987 (O_987,N_9665,N_9716);
nand UO_988 (O_988,N_9145,N_8635);
and UO_989 (O_989,N_9165,N_8936);
and UO_990 (O_990,N_9689,N_9876);
and UO_991 (O_991,N_8722,N_9946);
nand UO_992 (O_992,N_8666,N_8881);
nor UO_993 (O_993,N_9097,N_9817);
and UO_994 (O_994,N_9033,N_8259);
nand UO_995 (O_995,N_7823,N_7987);
nor UO_996 (O_996,N_7617,N_9059);
or UO_997 (O_997,N_8028,N_8709);
and UO_998 (O_998,N_8060,N_8719);
or UO_999 (O_999,N_8723,N_9690);
and UO_1000 (O_1000,N_9333,N_9697);
or UO_1001 (O_1001,N_8788,N_8265);
nor UO_1002 (O_1002,N_9124,N_7586);
nor UO_1003 (O_1003,N_9617,N_8906);
xor UO_1004 (O_1004,N_8326,N_9116);
nor UO_1005 (O_1005,N_9104,N_8422);
and UO_1006 (O_1006,N_8882,N_8163);
nand UO_1007 (O_1007,N_9388,N_7512);
and UO_1008 (O_1008,N_9132,N_8866);
nand UO_1009 (O_1009,N_9654,N_8814);
and UO_1010 (O_1010,N_9178,N_9687);
or UO_1011 (O_1011,N_9257,N_8193);
nand UO_1012 (O_1012,N_8733,N_9009);
or UO_1013 (O_1013,N_8461,N_9090);
or UO_1014 (O_1014,N_9078,N_7842);
nor UO_1015 (O_1015,N_9473,N_7820);
xor UO_1016 (O_1016,N_9435,N_8317);
and UO_1017 (O_1017,N_8017,N_8263);
and UO_1018 (O_1018,N_9286,N_8255);
nand UO_1019 (O_1019,N_9402,N_9468);
nand UO_1020 (O_1020,N_8324,N_7563);
nor UO_1021 (O_1021,N_8820,N_8180);
nor UO_1022 (O_1022,N_8385,N_9907);
nand UO_1023 (O_1023,N_8870,N_7806);
or UO_1024 (O_1024,N_8551,N_9049);
or UO_1025 (O_1025,N_9425,N_7702);
nand UO_1026 (O_1026,N_8909,N_9674);
nand UO_1027 (O_1027,N_9004,N_8352);
or UO_1028 (O_1028,N_9967,N_9563);
and UO_1029 (O_1029,N_9177,N_8295);
nand UO_1030 (O_1030,N_7618,N_8243);
nand UO_1031 (O_1031,N_9019,N_9739);
or UO_1032 (O_1032,N_9216,N_7927);
nand UO_1033 (O_1033,N_9587,N_7766);
nor UO_1034 (O_1034,N_8444,N_8935);
nand UO_1035 (O_1035,N_9113,N_8917);
and UO_1036 (O_1036,N_9115,N_8828);
and UO_1037 (O_1037,N_9679,N_7587);
or UO_1038 (O_1038,N_8403,N_8057);
nor UO_1039 (O_1039,N_7828,N_8844);
and UO_1040 (O_1040,N_8573,N_8298);
nand UO_1041 (O_1041,N_9006,N_8982);
nand UO_1042 (O_1042,N_8189,N_8596);
nand UO_1043 (O_1043,N_9308,N_8883);
and UO_1044 (O_1044,N_8978,N_8756);
or UO_1045 (O_1045,N_9123,N_9709);
nor UO_1046 (O_1046,N_8802,N_8142);
nor UO_1047 (O_1047,N_8077,N_7653);
xnor UO_1048 (O_1048,N_7932,N_9589);
and UO_1049 (O_1049,N_9240,N_7878);
or UO_1050 (O_1050,N_7668,N_9428);
and UO_1051 (O_1051,N_8729,N_7918);
nand UO_1052 (O_1052,N_7648,N_8048);
and UO_1053 (O_1053,N_7621,N_9806);
nand UO_1054 (O_1054,N_8806,N_8879);
and UO_1055 (O_1055,N_9875,N_7684);
or UO_1056 (O_1056,N_9327,N_8888);
and UO_1057 (O_1057,N_7944,N_8637);
nor UO_1058 (O_1058,N_9977,N_9433);
or UO_1059 (O_1059,N_8200,N_9763);
or UO_1060 (O_1060,N_9481,N_9556);
and UO_1061 (O_1061,N_9380,N_7559);
and UO_1062 (O_1062,N_8919,N_9942);
or UO_1063 (O_1063,N_7719,N_7726);
nand UO_1064 (O_1064,N_9933,N_9448);
nor UO_1065 (O_1065,N_9483,N_9725);
nand UO_1066 (O_1066,N_7674,N_9066);
and UO_1067 (O_1067,N_9796,N_8872);
nand UO_1068 (O_1068,N_8995,N_9720);
xor UO_1069 (O_1069,N_9409,N_9401);
nor UO_1070 (O_1070,N_9183,N_7862);
nand UO_1071 (O_1071,N_7501,N_9602);
and UO_1072 (O_1072,N_8395,N_9624);
nor UO_1073 (O_1073,N_8242,N_9452);
nand UO_1074 (O_1074,N_8845,N_9021);
or UO_1075 (O_1075,N_7509,N_8271);
or UO_1076 (O_1076,N_9509,N_7796);
and UO_1077 (O_1077,N_8486,N_7837);
and UO_1078 (O_1078,N_9243,N_8875);
or UO_1079 (O_1079,N_8115,N_9083);
nor UO_1080 (O_1080,N_8202,N_9773);
nor UO_1081 (O_1081,N_8769,N_7947);
and UO_1082 (O_1082,N_8548,N_8018);
and UO_1083 (O_1083,N_8405,N_8043);
and UO_1084 (O_1084,N_8230,N_7688);
nand UO_1085 (O_1085,N_8550,N_9284);
nor UO_1086 (O_1086,N_8578,N_9811);
nand UO_1087 (O_1087,N_8244,N_8487);
nor UO_1088 (O_1088,N_8497,N_8884);
and UO_1089 (O_1089,N_9110,N_9691);
and UO_1090 (O_1090,N_9839,N_8743);
nor UO_1091 (O_1091,N_9619,N_7754);
nand UO_1092 (O_1092,N_7835,N_9642);
or UO_1093 (O_1093,N_8944,N_7905);
or UO_1094 (O_1094,N_9419,N_9614);
and UO_1095 (O_1095,N_8196,N_8628);
and UO_1096 (O_1096,N_9063,N_7528);
nand UO_1097 (O_1097,N_8511,N_7965);
nand UO_1098 (O_1098,N_8449,N_8384);
or UO_1099 (O_1099,N_8315,N_7697);
and UO_1100 (O_1100,N_9453,N_9740);
nand UO_1101 (O_1101,N_7523,N_8685);
nand UO_1102 (O_1102,N_9793,N_9122);
or UO_1103 (O_1103,N_7930,N_9995);
nand UO_1104 (O_1104,N_7995,N_7780);
and UO_1105 (O_1105,N_8730,N_8602);
or UO_1106 (O_1106,N_8726,N_9202);
or UO_1107 (O_1107,N_9949,N_9443);
nor UO_1108 (O_1108,N_9650,N_9547);
or UO_1109 (O_1109,N_8000,N_8059);
or UO_1110 (O_1110,N_9251,N_9002);
nand UO_1111 (O_1111,N_7785,N_8011);
nor UO_1112 (O_1112,N_9223,N_7744);
nand UO_1113 (O_1113,N_9134,N_7681);
nand UO_1114 (O_1114,N_8988,N_9825);
nor UO_1115 (O_1115,N_8901,N_9117);
or UO_1116 (O_1116,N_9685,N_8140);
nor UO_1117 (O_1117,N_7710,N_8963);
nor UO_1118 (O_1118,N_7667,N_8691);
and UO_1119 (O_1119,N_8953,N_7596);
xor UO_1120 (O_1120,N_9418,N_9884);
nand UO_1121 (O_1121,N_9787,N_8055);
and UO_1122 (O_1122,N_8380,N_8062);
or UO_1123 (O_1123,N_9209,N_7949);
nor UO_1124 (O_1124,N_7892,N_8463);
and UO_1125 (O_1125,N_9405,N_9762);
nor UO_1126 (O_1126,N_8291,N_7524);
xnor UO_1127 (O_1127,N_9192,N_7797);
xnor UO_1128 (O_1128,N_7606,N_9867);
nand UO_1129 (O_1129,N_8095,N_9157);
or UO_1130 (O_1130,N_8023,N_8699);
or UO_1131 (O_1131,N_9931,N_8731);
xor UO_1132 (O_1132,N_9757,N_9727);
nor UO_1133 (O_1133,N_9276,N_9633);
and UO_1134 (O_1134,N_7849,N_9574);
nor UO_1135 (O_1135,N_7669,N_8702);
nand UO_1136 (O_1136,N_7777,N_9096);
nor UO_1137 (O_1137,N_8501,N_8529);
or UO_1138 (O_1138,N_9310,N_8113);
nand UO_1139 (O_1139,N_9997,N_7562);
nor UO_1140 (O_1140,N_8481,N_9328);
nand UO_1141 (O_1141,N_9444,N_8572);
nor UO_1142 (O_1142,N_9937,N_7713);
nand UO_1143 (O_1143,N_8452,N_8417);
nor UO_1144 (O_1144,N_7948,N_9715);
or UO_1145 (O_1145,N_8484,N_7652);
or UO_1146 (O_1146,N_9457,N_9513);
or UO_1147 (O_1147,N_7755,N_8856);
or UO_1148 (O_1148,N_8046,N_8639);
or UO_1149 (O_1149,N_7800,N_7554);
and UO_1150 (O_1150,N_7966,N_8251);
nor UO_1151 (O_1151,N_8932,N_9657);
nor UO_1152 (O_1152,N_8392,N_8605);
nand UO_1153 (O_1153,N_9467,N_8049);
nor UO_1154 (O_1154,N_9320,N_9325);
nor UO_1155 (O_1155,N_8143,N_8340);
nand UO_1156 (O_1156,N_9039,N_9823);
and UO_1157 (O_1157,N_7698,N_7551);
and UO_1158 (O_1158,N_9075,N_9872);
or UO_1159 (O_1159,N_7700,N_9915);
and UO_1160 (O_1160,N_8120,N_8968);
nand UO_1161 (O_1161,N_8608,N_9357);
nor UO_1162 (O_1162,N_8588,N_8414);
nand UO_1163 (O_1163,N_8091,N_8170);
or UO_1164 (O_1164,N_8861,N_9103);
nand UO_1165 (O_1165,N_7802,N_8574);
nor UO_1166 (O_1166,N_8761,N_9906);
nand UO_1167 (O_1167,N_9729,N_9041);
or UO_1168 (O_1168,N_7832,N_7887);
nor UO_1169 (O_1169,N_9180,N_8238);
nor UO_1170 (O_1170,N_9525,N_7679);
nor UO_1171 (O_1171,N_9889,N_9446);
nor UO_1172 (O_1172,N_9662,N_8964);
or UO_1173 (O_1173,N_8570,N_7801);
or UO_1174 (O_1174,N_9940,N_9363);
and UO_1175 (O_1175,N_8350,N_8256);
or UO_1176 (O_1176,N_8670,N_7661);
xor UO_1177 (O_1177,N_8286,N_7629);
and UO_1178 (O_1178,N_9705,N_7884);
or UO_1179 (O_1179,N_7565,N_9973);
or UO_1180 (O_1180,N_8784,N_9138);
and UO_1181 (O_1181,N_8003,N_8658);
nand UO_1182 (O_1182,N_9586,N_8660);
or UO_1183 (O_1183,N_9163,N_8367);
or UO_1184 (O_1184,N_9644,N_8716);
or UO_1185 (O_1185,N_9711,N_7759);
or UO_1186 (O_1186,N_7638,N_7787);
and UO_1187 (O_1187,N_8083,N_8031);
nand UO_1188 (O_1188,N_9480,N_8986);
and UO_1189 (O_1189,N_8895,N_8135);
or UO_1190 (O_1190,N_9571,N_8436);
or UO_1191 (O_1191,N_8934,N_8880);
or UO_1192 (O_1192,N_7928,N_8869);
nand UO_1193 (O_1193,N_8946,N_9008);
and UO_1194 (O_1194,N_7716,N_8854);
xor UO_1195 (O_1195,N_9133,N_9543);
nor UO_1196 (O_1196,N_9470,N_8683);
and UO_1197 (O_1197,N_9016,N_8819);
or UO_1198 (O_1198,N_9154,N_7752);
or UO_1199 (O_1199,N_8136,N_8400);
nand UO_1200 (O_1200,N_9449,N_8345);
nor UO_1201 (O_1201,N_7520,N_8362);
or UO_1202 (O_1202,N_8192,N_9227);
nor UO_1203 (O_1203,N_9590,N_9309);
nand UO_1204 (O_1204,N_8333,N_9348);
or UO_1205 (O_1205,N_9184,N_7967);
nand UO_1206 (O_1206,N_9355,N_9052);
and UO_1207 (O_1207,N_8793,N_9230);
or UO_1208 (O_1208,N_8065,N_9249);
or UO_1209 (O_1209,N_9786,N_9005);
or UO_1210 (O_1210,N_7753,N_9232);
or UO_1211 (O_1211,N_8480,N_8838);
nor UO_1212 (O_1212,N_9265,N_8312);
nand UO_1213 (O_1213,N_8569,N_8079);
or UO_1214 (O_1214,N_8778,N_7539);
or UO_1215 (O_1215,N_8110,N_8132);
and UO_1216 (O_1216,N_7870,N_9319);
or UO_1217 (O_1217,N_8126,N_7830);
and UO_1218 (O_1218,N_8394,N_9917);
nand UO_1219 (O_1219,N_9014,N_7643);
and UO_1220 (O_1220,N_7954,N_9770);
or UO_1221 (O_1221,N_8738,N_9300);
and UO_1222 (O_1222,N_8695,N_7640);
nand UO_1223 (O_1223,N_9386,N_8663);
nor UO_1224 (O_1224,N_8279,N_7853);
and UO_1225 (O_1225,N_9187,N_9520);
xnor UO_1226 (O_1226,N_7851,N_8093);
and UO_1227 (O_1227,N_7662,N_9935);
nand UO_1228 (O_1228,N_8358,N_9958);
or UO_1229 (O_1229,N_9717,N_9686);
nand UO_1230 (O_1230,N_8720,N_7663);
xor UO_1231 (O_1231,N_8531,N_7772);
or UO_1232 (O_1232,N_9023,N_7825);
nor UO_1233 (O_1233,N_8780,N_9597);
and UO_1234 (O_1234,N_7537,N_7871);
or UO_1235 (O_1235,N_9759,N_8792);
and UO_1236 (O_1236,N_9821,N_8682);
nand UO_1237 (O_1237,N_7646,N_7644);
nand UO_1238 (O_1238,N_7989,N_9466);
nand UO_1239 (O_1239,N_9539,N_8977);
and UO_1240 (O_1240,N_9922,N_8280);
nor UO_1241 (O_1241,N_8672,N_8725);
and UO_1242 (O_1242,N_7602,N_8773);
and UO_1243 (O_1243,N_7548,N_7896);
nand UO_1244 (O_1244,N_8627,N_9514);
nand UO_1245 (O_1245,N_9502,N_8008);
xnor UO_1246 (O_1246,N_7809,N_8476);
nand UO_1247 (O_1247,N_9164,N_8081);
and UO_1248 (O_1248,N_9001,N_7882);
nand UO_1249 (O_1249,N_8327,N_7535);
or UO_1250 (O_1250,N_8473,N_9540);
or UO_1251 (O_1251,N_8569,N_9513);
and UO_1252 (O_1252,N_8877,N_7875);
or UO_1253 (O_1253,N_9674,N_8848);
nand UO_1254 (O_1254,N_9480,N_8167);
xnor UO_1255 (O_1255,N_9169,N_9754);
and UO_1256 (O_1256,N_7605,N_8642);
nor UO_1257 (O_1257,N_8953,N_9512);
nor UO_1258 (O_1258,N_8596,N_9641);
nor UO_1259 (O_1259,N_7663,N_7682);
or UO_1260 (O_1260,N_9501,N_9724);
nor UO_1261 (O_1261,N_8954,N_9345);
nand UO_1262 (O_1262,N_7881,N_8198);
and UO_1263 (O_1263,N_9865,N_8015);
and UO_1264 (O_1264,N_7743,N_8890);
or UO_1265 (O_1265,N_9662,N_7551);
nor UO_1266 (O_1266,N_9845,N_7727);
xnor UO_1267 (O_1267,N_8820,N_7800);
nand UO_1268 (O_1268,N_9701,N_9402);
and UO_1269 (O_1269,N_7942,N_9406);
and UO_1270 (O_1270,N_8707,N_9498);
and UO_1271 (O_1271,N_9432,N_8343);
nor UO_1272 (O_1272,N_9980,N_9628);
nand UO_1273 (O_1273,N_9700,N_9612);
or UO_1274 (O_1274,N_8460,N_8668);
nor UO_1275 (O_1275,N_7813,N_9277);
nand UO_1276 (O_1276,N_7622,N_8706);
and UO_1277 (O_1277,N_8908,N_9032);
and UO_1278 (O_1278,N_8695,N_8181);
and UO_1279 (O_1279,N_7688,N_8769);
and UO_1280 (O_1280,N_8923,N_9781);
nor UO_1281 (O_1281,N_9829,N_8515);
and UO_1282 (O_1282,N_9105,N_8998);
or UO_1283 (O_1283,N_9148,N_8844);
and UO_1284 (O_1284,N_8978,N_9447);
and UO_1285 (O_1285,N_9621,N_8330);
or UO_1286 (O_1286,N_9760,N_9599);
or UO_1287 (O_1287,N_7945,N_7627);
and UO_1288 (O_1288,N_7748,N_7722);
and UO_1289 (O_1289,N_8219,N_8759);
nor UO_1290 (O_1290,N_9347,N_8833);
nand UO_1291 (O_1291,N_9011,N_8724);
nand UO_1292 (O_1292,N_7554,N_8900);
or UO_1293 (O_1293,N_9923,N_8430);
nor UO_1294 (O_1294,N_8533,N_9780);
and UO_1295 (O_1295,N_8637,N_7517);
nor UO_1296 (O_1296,N_8886,N_9006);
nand UO_1297 (O_1297,N_8296,N_8310);
nand UO_1298 (O_1298,N_8896,N_8665);
nor UO_1299 (O_1299,N_7861,N_8831);
nor UO_1300 (O_1300,N_9691,N_9163);
nand UO_1301 (O_1301,N_8455,N_9916);
and UO_1302 (O_1302,N_8200,N_9749);
nor UO_1303 (O_1303,N_8980,N_9019);
and UO_1304 (O_1304,N_8982,N_8564);
nor UO_1305 (O_1305,N_9610,N_8723);
or UO_1306 (O_1306,N_7995,N_7625);
nor UO_1307 (O_1307,N_7551,N_8705);
nor UO_1308 (O_1308,N_9578,N_8411);
nand UO_1309 (O_1309,N_9194,N_8369);
and UO_1310 (O_1310,N_9072,N_9165);
nor UO_1311 (O_1311,N_8820,N_8122);
nand UO_1312 (O_1312,N_9811,N_8566);
nand UO_1313 (O_1313,N_9916,N_8435);
and UO_1314 (O_1314,N_9853,N_9178);
nand UO_1315 (O_1315,N_8076,N_9405);
and UO_1316 (O_1316,N_9007,N_9189);
nand UO_1317 (O_1317,N_7923,N_8444);
nor UO_1318 (O_1318,N_9438,N_9771);
nor UO_1319 (O_1319,N_8382,N_9012);
nand UO_1320 (O_1320,N_8321,N_8314);
nor UO_1321 (O_1321,N_8280,N_7817);
and UO_1322 (O_1322,N_7976,N_8255);
nand UO_1323 (O_1323,N_7550,N_8899);
nand UO_1324 (O_1324,N_8094,N_8339);
and UO_1325 (O_1325,N_8721,N_8984);
or UO_1326 (O_1326,N_8877,N_9684);
nor UO_1327 (O_1327,N_8265,N_9812);
nand UO_1328 (O_1328,N_8355,N_9287);
nor UO_1329 (O_1329,N_9533,N_9681);
or UO_1330 (O_1330,N_7502,N_9033);
nand UO_1331 (O_1331,N_8335,N_9282);
or UO_1332 (O_1332,N_9124,N_9754);
xor UO_1333 (O_1333,N_7926,N_9420);
nand UO_1334 (O_1334,N_7560,N_8377);
nor UO_1335 (O_1335,N_7741,N_8940);
and UO_1336 (O_1336,N_7727,N_8828);
and UO_1337 (O_1337,N_9024,N_8683);
nand UO_1338 (O_1338,N_7974,N_7992);
and UO_1339 (O_1339,N_9454,N_9441);
or UO_1340 (O_1340,N_7568,N_9485);
and UO_1341 (O_1341,N_9681,N_8932);
or UO_1342 (O_1342,N_8964,N_9741);
and UO_1343 (O_1343,N_8763,N_7967);
nand UO_1344 (O_1344,N_8259,N_8486);
and UO_1345 (O_1345,N_8464,N_9707);
nand UO_1346 (O_1346,N_9105,N_8146);
xor UO_1347 (O_1347,N_8538,N_7968);
and UO_1348 (O_1348,N_9929,N_8440);
or UO_1349 (O_1349,N_8785,N_9602);
or UO_1350 (O_1350,N_8807,N_7676);
nand UO_1351 (O_1351,N_9170,N_9788);
nand UO_1352 (O_1352,N_8254,N_9367);
nand UO_1353 (O_1353,N_7635,N_9635);
xor UO_1354 (O_1354,N_8168,N_9280);
or UO_1355 (O_1355,N_8854,N_9081);
nor UO_1356 (O_1356,N_9945,N_9297);
nand UO_1357 (O_1357,N_8691,N_9127);
nand UO_1358 (O_1358,N_9102,N_8337);
nor UO_1359 (O_1359,N_9762,N_9136);
or UO_1360 (O_1360,N_9697,N_9822);
nor UO_1361 (O_1361,N_8824,N_8844);
or UO_1362 (O_1362,N_9422,N_8455);
or UO_1363 (O_1363,N_9383,N_9075);
or UO_1364 (O_1364,N_9044,N_8767);
nor UO_1365 (O_1365,N_7680,N_7555);
nand UO_1366 (O_1366,N_8278,N_7966);
xnor UO_1367 (O_1367,N_9646,N_7907);
and UO_1368 (O_1368,N_7503,N_7588);
or UO_1369 (O_1369,N_8541,N_7864);
or UO_1370 (O_1370,N_8383,N_7793);
and UO_1371 (O_1371,N_9383,N_9066);
nor UO_1372 (O_1372,N_7799,N_8421);
and UO_1373 (O_1373,N_8203,N_8427);
or UO_1374 (O_1374,N_9427,N_8736);
or UO_1375 (O_1375,N_7709,N_8677);
and UO_1376 (O_1376,N_8481,N_8864);
nor UO_1377 (O_1377,N_9812,N_9373);
and UO_1378 (O_1378,N_9413,N_8834);
nand UO_1379 (O_1379,N_9479,N_9789);
or UO_1380 (O_1380,N_8281,N_8205);
and UO_1381 (O_1381,N_8892,N_8956);
nand UO_1382 (O_1382,N_9479,N_8362);
nor UO_1383 (O_1383,N_9087,N_8065);
nor UO_1384 (O_1384,N_8519,N_9578);
and UO_1385 (O_1385,N_8660,N_9489);
nor UO_1386 (O_1386,N_8330,N_9599);
and UO_1387 (O_1387,N_7864,N_9227);
nor UO_1388 (O_1388,N_9768,N_9293);
and UO_1389 (O_1389,N_7898,N_9261);
and UO_1390 (O_1390,N_7668,N_7902);
nand UO_1391 (O_1391,N_9207,N_8716);
nor UO_1392 (O_1392,N_7561,N_8124);
and UO_1393 (O_1393,N_8668,N_8017);
nand UO_1394 (O_1394,N_8491,N_9559);
and UO_1395 (O_1395,N_8326,N_8092);
nand UO_1396 (O_1396,N_7644,N_7709);
nor UO_1397 (O_1397,N_8932,N_9723);
nor UO_1398 (O_1398,N_8462,N_7894);
and UO_1399 (O_1399,N_8004,N_9294);
nand UO_1400 (O_1400,N_8886,N_9290);
or UO_1401 (O_1401,N_8713,N_7630);
nand UO_1402 (O_1402,N_8055,N_8332);
or UO_1403 (O_1403,N_8064,N_8137);
or UO_1404 (O_1404,N_7560,N_8509);
and UO_1405 (O_1405,N_9348,N_9832);
nor UO_1406 (O_1406,N_9681,N_9933);
nand UO_1407 (O_1407,N_7902,N_9343);
nand UO_1408 (O_1408,N_8680,N_9151);
or UO_1409 (O_1409,N_8625,N_8547);
nor UO_1410 (O_1410,N_7601,N_9550);
and UO_1411 (O_1411,N_9551,N_9439);
nor UO_1412 (O_1412,N_7635,N_9130);
nor UO_1413 (O_1413,N_8850,N_9580);
and UO_1414 (O_1414,N_8689,N_9272);
and UO_1415 (O_1415,N_9439,N_8038);
nor UO_1416 (O_1416,N_9185,N_9829);
or UO_1417 (O_1417,N_8841,N_7970);
or UO_1418 (O_1418,N_9498,N_8290);
and UO_1419 (O_1419,N_7984,N_8600);
nand UO_1420 (O_1420,N_7546,N_8510);
nand UO_1421 (O_1421,N_7705,N_8203);
nand UO_1422 (O_1422,N_7964,N_8971);
or UO_1423 (O_1423,N_8742,N_9584);
nor UO_1424 (O_1424,N_9662,N_9140);
or UO_1425 (O_1425,N_9155,N_8347);
and UO_1426 (O_1426,N_8969,N_8819);
nand UO_1427 (O_1427,N_7960,N_8213);
nor UO_1428 (O_1428,N_9563,N_8201);
nand UO_1429 (O_1429,N_8173,N_7969);
or UO_1430 (O_1430,N_7934,N_9375);
nor UO_1431 (O_1431,N_8443,N_8295);
or UO_1432 (O_1432,N_9269,N_8799);
nor UO_1433 (O_1433,N_9020,N_9072);
and UO_1434 (O_1434,N_9878,N_8297);
nand UO_1435 (O_1435,N_9074,N_9752);
nand UO_1436 (O_1436,N_8073,N_9925);
nand UO_1437 (O_1437,N_8243,N_7970);
nor UO_1438 (O_1438,N_9825,N_8022);
or UO_1439 (O_1439,N_9312,N_9877);
nor UO_1440 (O_1440,N_7938,N_9051);
or UO_1441 (O_1441,N_9553,N_9763);
nand UO_1442 (O_1442,N_9840,N_8494);
or UO_1443 (O_1443,N_8360,N_7805);
or UO_1444 (O_1444,N_8044,N_8073);
nand UO_1445 (O_1445,N_9208,N_8725);
nor UO_1446 (O_1446,N_7941,N_9148);
or UO_1447 (O_1447,N_7637,N_7917);
and UO_1448 (O_1448,N_8623,N_8045);
nand UO_1449 (O_1449,N_8403,N_8952);
and UO_1450 (O_1450,N_9050,N_8516);
nand UO_1451 (O_1451,N_9553,N_7678);
nand UO_1452 (O_1452,N_9088,N_8095);
nand UO_1453 (O_1453,N_8111,N_9823);
nand UO_1454 (O_1454,N_9361,N_7645);
or UO_1455 (O_1455,N_8728,N_8005);
or UO_1456 (O_1456,N_9624,N_7717);
nor UO_1457 (O_1457,N_8504,N_9039);
and UO_1458 (O_1458,N_9606,N_9439);
nor UO_1459 (O_1459,N_8202,N_9491);
and UO_1460 (O_1460,N_9246,N_7591);
or UO_1461 (O_1461,N_8472,N_8003);
nand UO_1462 (O_1462,N_8772,N_8745);
or UO_1463 (O_1463,N_7828,N_8431);
and UO_1464 (O_1464,N_8375,N_8237);
nor UO_1465 (O_1465,N_9923,N_7523);
nor UO_1466 (O_1466,N_9606,N_8662);
and UO_1467 (O_1467,N_8008,N_9858);
nand UO_1468 (O_1468,N_7651,N_9124);
nand UO_1469 (O_1469,N_9991,N_9131);
nand UO_1470 (O_1470,N_8407,N_8740);
nand UO_1471 (O_1471,N_8588,N_9395);
and UO_1472 (O_1472,N_8239,N_9027);
nor UO_1473 (O_1473,N_8985,N_9238);
and UO_1474 (O_1474,N_9234,N_8460);
or UO_1475 (O_1475,N_7741,N_7768);
nor UO_1476 (O_1476,N_9434,N_7782);
nand UO_1477 (O_1477,N_8735,N_9164);
nor UO_1478 (O_1478,N_9565,N_9728);
or UO_1479 (O_1479,N_8498,N_7974);
and UO_1480 (O_1480,N_7685,N_7698);
nand UO_1481 (O_1481,N_9264,N_8493);
and UO_1482 (O_1482,N_9933,N_9969);
nor UO_1483 (O_1483,N_9489,N_9291);
nor UO_1484 (O_1484,N_9091,N_8339);
and UO_1485 (O_1485,N_8230,N_9333);
or UO_1486 (O_1486,N_9305,N_7986);
and UO_1487 (O_1487,N_7953,N_9668);
nor UO_1488 (O_1488,N_7697,N_9507);
or UO_1489 (O_1489,N_8860,N_9618);
and UO_1490 (O_1490,N_9796,N_9631);
nor UO_1491 (O_1491,N_7644,N_9482);
nor UO_1492 (O_1492,N_7973,N_7760);
or UO_1493 (O_1493,N_9161,N_9324);
and UO_1494 (O_1494,N_8568,N_9204);
nor UO_1495 (O_1495,N_9039,N_9231);
nor UO_1496 (O_1496,N_9852,N_8684);
or UO_1497 (O_1497,N_8287,N_8116);
nor UO_1498 (O_1498,N_9901,N_8579);
and UO_1499 (O_1499,N_9315,N_9022);
endmodule