module basic_1000_10000_1500_20_levels_5xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nand U0 (N_0,In_868,In_172);
nor U1 (N_1,In_80,In_971);
nor U2 (N_2,In_321,In_715);
nor U3 (N_3,In_532,In_422);
nand U4 (N_4,In_564,In_293);
nand U5 (N_5,In_645,In_741);
nand U6 (N_6,In_704,In_800);
or U7 (N_7,In_947,In_765);
nor U8 (N_8,In_539,In_614);
and U9 (N_9,In_142,In_571);
nand U10 (N_10,In_607,In_748);
nand U11 (N_11,In_727,In_18);
nand U12 (N_12,In_239,In_481);
nand U13 (N_13,In_753,In_884);
and U14 (N_14,In_109,In_275);
or U15 (N_15,In_984,In_940);
or U16 (N_16,In_896,In_937);
nor U17 (N_17,In_465,In_955);
nand U18 (N_18,In_7,In_804);
nor U19 (N_19,In_905,In_276);
or U20 (N_20,In_232,In_813);
nand U21 (N_21,In_624,In_912);
and U22 (N_22,In_808,In_633);
xnor U23 (N_23,In_987,In_62);
nor U24 (N_24,In_916,In_157);
nand U25 (N_25,In_6,In_897);
xor U26 (N_26,In_272,In_784);
nand U27 (N_27,In_587,In_924);
nand U28 (N_28,In_467,In_212);
nor U29 (N_29,In_156,In_977);
or U30 (N_30,In_166,In_304);
or U31 (N_31,In_821,In_299);
nor U32 (N_32,In_552,In_946);
nand U33 (N_33,In_345,In_12);
and U34 (N_34,In_577,In_181);
nand U35 (N_35,In_42,In_547);
and U36 (N_36,In_835,In_891);
nor U37 (N_37,In_187,In_469);
nor U38 (N_38,In_883,In_847);
or U39 (N_39,In_416,In_589);
or U40 (N_40,In_854,In_330);
nor U41 (N_41,In_147,In_529);
nand U42 (N_42,In_122,In_637);
and U43 (N_43,In_355,In_494);
nand U44 (N_44,In_747,In_409);
xnor U45 (N_45,In_68,In_178);
and U46 (N_46,In_591,In_592);
nor U47 (N_47,In_100,In_491);
nor U48 (N_48,In_931,In_849);
xnor U49 (N_49,In_632,In_191);
or U50 (N_50,In_28,In_322);
or U51 (N_51,In_240,In_521);
or U52 (N_52,In_381,In_489);
and U53 (N_53,In_86,In_132);
and U54 (N_54,In_600,In_795);
xor U55 (N_55,In_210,In_586);
and U56 (N_56,In_155,In_549);
and U57 (N_57,In_890,In_346);
nor U58 (N_58,In_113,In_387);
nand U59 (N_59,In_140,In_995);
nand U60 (N_60,In_966,In_92);
or U61 (N_61,In_329,In_828);
nand U62 (N_62,In_368,In_930);
or U63 (N_63,In_201,In_697);
xor U64 (N_64,In_510,In_246);
or U65 (N_65,In_986,In_651);
nor U66 (N_66,In_812,In_582);
nor U67 (N_67,In_110,In_38);
or U68 (N_68,In_681,In_593);
xnor U69 (N_69,In_174,In_935);
nor U70 (N_70,In_39,In_457);
and U71 (N_71,In_815,In_135);
and U72 (N_72,In_5,In_447);
and U73 (N_73,In_833,In_320);
nand U74 (N_74,In_117,In_779);
nand U75 (N_75,In_856,In_985);
and U76 (N_76,In_388,In_885);
nor U77 (N_77,In_126,In_256);
or U78 (N_78,In_899,In_273);
nand U79 (N_79,In_504,In_151);
or U80 (N_80,In_588,In_572);
and U81 (N_81,In_575,In_215);
nor U82 (N_82,In_9,In_291);
nand U83 (N_83,In_186,In_628);
and U84 (N_84,In_541,In_846);
or U85 (N_85,In_162,In_486);
nand U86 (N_86,In_520,In_604);
or U87 (N_87,In_200,In_373);
or U88 (N_88,In_456,In_376);
or U89 (N_89,In_347,In_20);
or U90 (N_90,In_507,In_745);
or U91 (N_91,In_743,In_356);
nand U92 (N_92,In_620,In_769);
or U93 (N_93,In_53,In_669);
or U94 (N_94,In_115,In_725);
nand U95 (N_95,In_663,In_889);
and U96 (N_96,In_440,In_943);
and U97 (N_97,In_973,In_951);
nand U98 (N_98,In_948,In_735);
nand U99 (N_99,In_662,In_701);
nor U100 (N_100,In_83,In_423);
and U101 (N_101,In_114,In_400);
or U102 (N_102,In_960,In_404);
nand U103 (N_103,In_517,In_907);
nand U104 (N_104,In_466,In_194);
and U105 (N_105,In_768,In_406);
or U106 (N_106,In_622,In_313);
nand U107 (N_107,In_359,In_585);
nand U108 (N_108,In_554,In_534);
or U109 (N_109,In_934,In_683);
nand U110 (N_110,In_206,In_432);
and U111 (N_111,In_125,In_842);
nand U112 (N_112,In_926,In_249);
or U113 (N_113,In_69,In_384);
nand U114 (N_114,In_789,In_402);
nand U115 (N_115,In_556,In_665);
nand U116 (N_116,In_158,In_791);
or U117 (N_117,In_403,In_807);
nand U118 (N_118,In_454,In_234);
nand U119 (N_119,In_785,In_288);
or U120 (N_120,In_268,In_188);
or U121 (N_121,In_182,In_859);
xnor U122 (N_122,In_225,In_143);
nor U123 (N_123,In_555,In_991);
nor U124 (N_124,In_533,In_13);
nand U125 (N_125,In_325,In_141);
xnor U126 (N_126,In_711,In_380);
nor U127 (N_127,In_668,In_640);
nand U128 (N_128,In_138,In_619);
nor U129 (N_129,In_327,In_929);
nand U130 (N_130,In_505,In_183);
or U131 (N_131,In_963,In_328);
nor U132 (N_132,In_999,In_26);
nor U133 (N_133,In_817,In_365);
nand U134 (N_134,In_244,In_612);
nor U135 (N_135,In_371,In_750);
xor U136 (N_136,In_30,In_261);
or U137 (N_137,In_524,In_468);
and U138 (N_138,In_776,In_379);
and U139 (N_139,In_732,In_220);
and U140 (N_140,In_148,In_687);
or U141 (N_141,In_602,In_267);
or U142 (N_142,In_566,In_513);
nand U143 (N_143,In_265,In_294);
and U144 (N_144,In_251,In_694);
or U145 (N_145,In_527,In_230);
xor U146 (N_146,In_95,In_199);
nor U147 (N_147,In_672,In_799);
nand U148 (N_148,In_969,In_198);
or U149 (N_149,In_439,In_255);
nand U150 (N_150,In_87,In_67);
nand U151 (N_151,In_480,In_642);
nand U152 (N_152,In_271,In_302);
and U153 (N_153,In_975,In_19);
or U154 (N_154,In_522,In_146);
and U155 (N_155,In_295,In_836);
nor U156 (N_156,In_892,In_248);
nand U157 (N_157,In_362,In_245);
nand U158 (N_158,In_431,In_264);
and U159 (N_159,In_543,In_340);
nand U160 (N_160,In_15,In_184);
or U161 (N_161,In_305,In_176);
and U162 (N_162,In_703,In_2);
and U163 (N_163,In_563,In_528);
nand U164 (N_164,In_129,In_959);
and U165 (N_165,In_565,In_675);
or U166 (N_166,In_464,In_414);
and U167 (N_167,In_170,In_385);
nand U168 (N_168,In_133,In_914);
or U169 (N_169,In_211,In_636);
xor U170 (N_170,In_280,In_797);
nor U171 (N_171,In_853,In_289);
and U172 (N_172,In_569,In_269);
nor U173 (N_173,In_686,In_11);
nand U174 (N_174,In_980,In_196);
nand U175 (N_175,In_60,In_8);
or U176 (N_176,In_942,In_514);
xnor U177 (N_177,In_945,In_992);
and U178 (N_178,In_661,In_644);
or U179 (N_179,In_226,In_185);
or U180 (N_180,In_578,In_886);
nor U181 (N_181,In_242,In_277);
or U182 (N_182,In_775,In_746);
xnor U183 (N_183,In_428,In_670);
or U184 (N_184,In_145,In_780);
or U185 (N_185,In_258,In_895);
and U186 (N_186,In_219,In_879);
and U187 (N_187,In_699,In_643);
or U188 (N_188,In_377,In_845);
nand U189 (N_189,In_771,In_820);
xor U190 (N_190,In_103,In_284);
nand U191 (N_191,In_153,In_994);
or U192 (N_192,In_502,In_337);
xor U193 (N_193,In_306,In_736);
and U194 (N_194,In_819,In_606);
nor U195 (N_195,In_236,In_579);
xnor U196 (N_196,In_237,In_667);
nand U197 (N_197,In_460,In_352);
nor U198 (N_198,In_674,In_487);
nand U199 (N_199,In_283,In_950);
and U200 (N_200,In_250,In_372);
nand U201 (N_201,In_827,In_72);
nor U202 (N_202,In_584,In_621);
nand U203 (N_203,In_99,In_709);
nor U204 (N_204,In_550,In_843);
nor U205 (N_205,In_506,In_231);
and U206 (N_206,In_4,In_292);
nor U207 (N_207,In_673,In_485);
and U208 (N_208,In_296,In_35);
and U209 (N_209,In_475,In_855);
or U210 (N_210,In_898,In_708);
and U211 (N_211,In_266,In_446);
nor U212 (N_212,In_48,In_253);
nor U213 (N_213,In_36,In_370);
or U214 (N_214,In_676,In_417);
nand U215 (N_215,In_364,In_197);
or U216 (N_216,In_548,In_262);
or U217 (N_217,In_297,In_334);
or U218 (N_218,In_77,In_783);
and U219 (N_219,In_171,In_756);
or U220 (N_220,In_10,In_832);
nor U221 (N_221,In_259,In_315);
nor U222 (N_222,In_802,In_906);
nand U223 (N_223,In_221,In_411);
nand U224 (N_224,In_875,In_106);
or U225 (N_225,In_169,In_45);
xor U226 (N_226,In_508,In_326);
nor U227 (N_227,In_649,In_625);
nor U228 (N_228,In_722,In_23);
or U229 (N_229,In_168,In_43);
and U230 (N_230,In_415,In_434);
nand U231 (N_231,In_85,In_323);
nor U232 (N_232,In_243,In_961);
xor U233 (N_233,In_119,In_438);
nor U234 (N_234,In_707,In_887);
xor U235 (N_235,In_751,In_163);
nand U236 (N_236,In_344,In_495);
and U237 (N_237,In_925,In_204);
or U238 (N_238,In_123,In_613);
nor U239 (N_239,In_413,In_816);
nor U240 (N_240,In_826,In_656);
and U241 (N_241,In_616,In_610);
nand U242 (N_242,In_37,In_848);
and U243 (N_243,In_623,In_611);
and U244 (N_244,In_331,In_837);
nor U245 (N_245,In_974,In_300);
or U246 (N_246,In_471,In_858);
or U247 (N_247,In_40,In_378);
nand U248 (N_248,In_778,In_764);
nor U249 (N_249,In_958,In_173);
nor U250 (N_250,In_801,In_354);
nor U251 (N_251,In_358,In_719);
or U252 (N_252,In_928,In_97);
nor U253 (N_253,In_570,In_536);
xor U254 (N_254,In_693,In_923);
and U255 (N_255,In_429,In_224);
and U256 (N_256,In_882,In_71);
or U257 (N_257,In_617,In_44);
nor U258 (N_258,In_64,In_618);
nor U259 (N_259,In_518,In_583);
nor U260 (N_260,In_702,In_574);
nand U261 (N_261,In_729,In_758);
and U262 (N_262,In_763,In_105);
nand U263 (N_263,In_629,In_918);
nor U264 (N_264,In_314,In_81);
xor U265 (N_265,In_630,In_312);
and U266 (N_266,In_876,In_130);
xnor U267 (N_267,In_452,In_58);
nand U268 (N_268,In_634,In_410);
and U269 (N_269,In_692,In_399);
and U270 (N_270,In_360,In_93);
or U271 (N_271,In_691,In_685);
nor U272 (N_272,In_705,In_782);
or U273 (N_273,In_316,In_332);
or U274 (N_274,In_559,In_567);
nor U275 (N_275,In_988,In_476);
or U276 (N_276,In_956,In_531);
or U277 (N_277,In_757,In_363);
and U278 (N_278,In_671,In_73);
and U279 (N_279,In_852,In_754);
or U280 (N_280,In_728,In_154);
and U281 (N_281,In_558,In_927);
or U282 (N_282,In_420,In_866);
and U283 (N_283,In_762,In_461);
xnor U284 (N_284,In_235,In_160);
nand U285 (N_285,In_398,In_850);
nand U286 (N_286,In_121,In_396);
and U287 (N_287,In_957,In_752);
and U288 (N_288,In_418,In_760);
and U289 (N_289,In_336,In_482);
nand U290 (N_290,In_823,In_677);
xor U291 (N_291,In_989,In_63);
nand U292 (N_292,In_473,In_915);
and U293 (N_293,In_490,In_165);
and U294 (N_294,In_968,In_825);
nor U295 (N_295,In_700,In_793);
nor U296 (N_296,In_523,In_311);
nand U297 (N_297,In_860,In_167);
or U298 (N_298,In_734,In_537);
nor U299 (N_299,In_773,In_605);
nand U300 (N_300,In_310,In_118);
or U301 (N_301,In_497,In_803);
nand U302 (N_302,In_688,In_839);
nor U303 (N_303,In_1,In_79);
nor U304 (N_304,In_357,In_120);
and U305 (N_305,In_208,In_116);
or U306 (N_306,In_361,In_350);
nor U307 (N_307,In_449,In_862);
nand U308 (N_308,In_213,In_82);
nor U309 (N_309,In_192,In_479);
nand U310 (N_310,In_412,In_718);
nor U311 (N_311,In_52,In_695);
or U312 (N_312,In_144,In_519);
and U313 (N_313,In_888,In_721);
nand U314 (N_314,In_444,In_54);
nand U315 (N_315,In_421,In_603);
nand U316 (N_316,In_822,In_104);
and U317 (N_317,In_70,In_279);
and U318 (N_318,In_902,In_720);
nor U319 (N_319,In_561,In_838);
and U320 (N_320,In_921,In_581);
and U321 (N_321,In_349,In_731);
nand U322 (N_322,In_809,In_425);
nor U323 (N_323,In_458,In_137);
nor U324 (N_324,In_638,In_499);
and U325 (N_325,In_75,In_910);
xor U326 (N_326,In_366,In_98);
nor U327 (N_327,In_515,In_228);
and U328 (N_328,In_874,In_512);
nor U329 (N_329,In_919,In_430);
or U330 (N_330,In_737,In_865);
nand U331 (N_331,In_500,In_319);
or U332 (N_332,In_938,In_911);
nand U333 (N_333,In_426,In_223);
and U334 (N_334,In_792,In_904);
nor U335 (N_335,In_287,In_786);
xnor U336 (N_336,In_599,In_341);
nor U337 (N_337,In_682,In_798);
nand U338 (N_338,In_608,In_351);
nor U339 (N_339,In_450,In_657);
and U340 (N_340,In_180,In_716);
nand U341 (N_341,In_857,In_998);
xnor U342 (N_342,In_690,In_134);
nor U343 (N_343,In_94,In_979);
nand U344 (N_344,In_596,In_867);
and U345 (N_345,In_818,In_900);
or U346 (N_346,In_560,In_774);
or U347 (N_347,In_260,In_553);
or U348 (N_348,In_841,In_679);
or U349 (N_349,In_913,In_546);
and U350 (N_350,In_724,In_335);
nand U351 (N_351,In_342,In_189);
and U352 (N_352,In_107,In_427);
nor U353 (N_353,In_573,In_65);
nor U354 (N_354,In_698,In_57);
xnor U355 (N_355,In_477,In_562);
nand U356 (N_356,In_241,In_492);
and U357 (N_357,In_723,In_650);
or U358 (N_358,In_324,In_829);
or U359 (N_359,In_161,In_834);
or U360 (N_360,In_863,In_538);
and U361 (N_361,In_395,In_767);
nor U362 (N_362,In_917,In_31);
and U363 (N_363,In_353,In_759);
nand U364 (N_364,In_831,In_944);
or U365 (N_365,In_257,In_595);
and U366 (N_366,In_932,In_348);
or U367 (N_367,In_684,In_824);
nand U368 (N_368,In_503,In_463);
or U369 (N_369,In_659,In_392);
or U370 (N_370,In_953,In_405);
nor U371 (N_371,In_34,In_811);
nor U372 (N_372,In_127,In_175);
xnor U373 (N_373,In_96,In_794);
and U374 (N_374,In_216,In_136);
xor U375 (N_375,In_761,In_787);
nand U376 (N_376,In_796,In_997);
or U377 (N_377,In_949,In_526);
nor U378 (N_378,In_66,In_710);
or U379 (N_379,In_954,In_22);
nor U380 (N_380,In_89,In_788);
or U381 (N_381,In_478,In_501);
nor U382 (N_382,In_733,In_941);
nand U383 (N_383,In_726,In_993);
nand U384 (N_384,In_666,In_646);
and U385 (N_385,In_445,In_655);
nor U386 (N_386,In_777,In_551);
or U387 (N_387,In_386,In_483);
and U388 (N_388,In_47,In_576);
nor U389 (N_389,In_227,In_990);
nand U390 (N_390,In_338,In_511);
nand U391 (N_391,In_738,In_76);
nor U392 (N_392,In_55,In_755);
and U393 (N_393,In_195,In_936);
and U394 (N_394,In_689,In_790);
nor U395 (N_395,In_772,In_74);
nand U396 (N_396,In_920,In_88);
and U397 (N_397,In_844,In_205);
or U398 (N_398,In_877,In_781);
nor U399 (N_399,In_870,In_880);
or U400 (N_400,In_909,In_263);
nand U401 (N_401,In_301,In_601);
nor U402 (N_402,In_568,In_627);
xnor U403 (N_403,In_744,In_393);
nand U404 (N_404,In_470,In_871);
nand U405 (N_405,In_922,In_17);
and U406 (N_406,In_878,In_982);
and U407 (N_407,In_648,In_408);
nor U408 (N_408,In_742,In_29);
nor U409 (N_409,In_952,In_660);
and U410 (N_410,In_965,In_308);
or U411 (N_411,In_49,In_32);
or U412 (N_412,In_540,In_442);
nand U413 (N_413,In_493,In_474);
xor U414 (N_414,In_25,In_881);
and U415 (N_415,In_298,In_309);
and U416 (N_416,In_278,In_436);
nor U417 (N_417,In_401,In_840);
nor U418 (N_418,In_978,In_459);
and U419 (N_419,In_626,In_545);
or U420 (N_420,In_641,In_962);
nor U421 (N_421,In_90,In_150);
or U422 (N_422,In_441,In_706);
nor U423 (N_423,In_318,In_714);
or U424 (N_424,In_903,In_805);
nand U425 (N_425,In_873,In_27);
nor U426 (N_426,In_317,In_339);
nand U427 (N_427,In_3,In_967);
nor U428 (N_428,In_383,In_713);
and U429 (N_429,In_557,In_407);
or U430 (N_430,In_981,In_207);
nor U431 (N_431,In_307,In_484);
and U432 (N_432,In_597,In_149);
or U433 (N_433,In_433,In_810);
or U434 (N_434,In_391,In_766);
or U435 (N_435,In_290,In_56);
or U436 (N_436,In_647,In_50);
nor U437 (N_437,In_159,In_394);
or U438 (N_438,In_124,In_964);
nor U439 (N_439,In_509,In_41);
nor U440 (N_440,In_303,In_631);
xnor U441 (N_441,In_525,In_369);
nor U442 (N_442,In_437,In_84);
nor U443 (N_443,In_102,In_488);
nand U444 (N_444,In_594,In_609);
and U445 (N_445,In_893,In_740);
or U446 (N_446,In_749,In_131);
and U447 (N_447,In_639,In_535);
nand U448 (N_448,In_374,In_128);
or U449 (N_449,In_544,In_635);
and U450 (N_450,In_229,In_238);
and U451 (N_451,In_164,In_983);
nand U452 (N_452,In_462,In_190);
nand U453 (N_453,In_901,In_654);
or U454 (N_454,In_770,In_0);
nor U455 (N_455,In_996,In_448);
nor U456 (N_456,In_869,In_658);
nor U457 (N_457,In_247,In_976);
or U458 (N_458,In_21,In_179);
and U459 (N_459,In_443,In_453);
nand U460 (N_460,In_598,In_222);
xor U461 (N_461,In_516,In_375);
xor U462 (N_462,In_894,In_972);
or U463 (N_463,In_343,In_14);
nand U464 (N_464,In_152,In_664);
nor U465 (N_465,In_217,In_270);
and U466 (N_466,In_970,In_419);
and U467 (N_467,In_46,In_939);
and U468 (N_468,In_218,In_542);
and U469 (N_469,In_451,In_615);
and U470 (N_470,In_193,In_590);
nor U471 (N_471,In_908,In_139);
or U472 (N_472,In_814,In_252);
or U473 (N_473,In_397,In_696);
or U474 (N_474,In_16,In_496);
nand U475 (N_475,In_367,In_861);
nor U476 (N_476,In_712,In_233);
nand U477 (N_477,In_51,In_389);
nor U478 (N_478,In_112,In_203);
and U479 (N_479,In_455,In_717);
nand U480 (N_480,In_111,In_806);
nand U481 (N_481,In_498,In_254);
or U482 (N_482,In_864,In_739);
xor U483 (N_483,In_333,In_24);
or U484 (N_484,In_851,In_274);
nand U485 (N_485,In_91,In_872);
nand U486 (N_486,In_101,In_59);
nand U487 (N_487,In_108,In_214);
nor U488 (N_488,In_678,In_33);
and U489 (N_489,In_382,In_285);
and U490 (N_490,In_281,In_730);
or U491 (N_491,In_530,In_652);
xnor U492 (N_492,In_435,In_78);
and U493 (N_493,In_830,In_282);
or U494 (N_494,In_680,In_424);
or U495 (N_495,In_472,In_933);
nand U496 (N_496,In_202,In_177);
nand U497 (N_497,In_209,In_390);
nor U498 (N_498,In_61,In_286);
or U499 (N_499,In_580,In_653);
xor U500 (N_500,N_417,N_487);
xor U501 (N_501,N_243,N_126);
nand U502 (N_502,N_16,N_175);
xnor U503 (N_503,N_477,N_202);
and U504 (N_504,N_332,N_107);
nor U505 (N_505,N_427,N_342);
and U506 (N_506,N_220,N_372);
nand U507 (N_507,N_6,N_266);
xor U508 (N_508,N_436,N_5);
and U509 (N_509,N_203,N_413);
and U510 (N_510,N_249,N_9);
and U511 (N_511,N_331,N_358);
or U512 (N_512,N_221,N_247);
and U513 (N_513,N_218,N_44);
nor U514 (N_514,N_227,N_2);
or U515 (N_515,N_379,N_228);
nand U516 (N_516,N_256,N_190);
xnor U517 (N_517,N_398,N_22);
or U518 (N_518,N_482,N_262);
and U519 (N_519,N_181,N_403);
or U520 (N_520,N_86,N_248);
and U521 (N_521,N_21,N_172);
nor U522 (N_522,N_324,N_38);
nor U523 (N_523,N_122,N_49);
nand U524 (N_524,N_235,N_307);
and U525 (N_525,N_41,N_498);
nand U526 (N_526,N_215,N_466);
or U527 (N_527,N_278,N_164);
xor U528 (N_528,N_40,N_318);
nor U529 (N_529,N_406,N_230);
nand U530 (N_530,N_418,N_73);
nor U531 (N_531,N_29,N_98);
nand U532 (N_532,N_66,N_407);
or U533 (N_533,N_17,N_113);
or U534 (N_534,N_183,N_286);
nand U535 (N_535,N_327,N_36);
or U536 (N_536,N_238,N_82);
nor U537 (N_537,N_223,N_316);
or U538 (N_538,N_188,N_132);
and U539 (N_539,N_51,N_14);
or U540 (N_540,N_37,N_153);
or U541 (N_541,N_437,N_289);
or U542 (N_542,N_157,N_411);
and U543 (N_543,N_27,N_155);
nor U544 (N_544,N_401,N_18);
nand U545 (N_545,N_280,N_294);
xor U546 (N_546,N_260,N_75);
and U547 (N_547,N_370,N_217);
nor U548 (N_548,N_396,N_297);
and U549 (N_549,N_321,N_384);
nand U550 (N_550,N_283,N_269);
nor U551 (N_551,N_369,N_293);
xnor U552 (N_552,N_15,N_141);
and U553 (N_553,N_474,N_208);
and U554 (N_554,N_140,N_363);
or U555 (N_555,N_494,N_77);
nand U556 (N_556,N_79,N_391);
nand U557 (N_557,N_313,N_479);
and U558 (N_558,N_186,N_351);
nor U559 (N_559,N_152,N_224);
nand U560 (N_560,N_233,N_60);
nor U561 (N_561,N_315,N_275);
or U562 (N_562,N_345,N_88);
or U563 (N_563,N_287,N_229);
nand U564 (N_564,N_291,N_168);
nor U565 (N_565,N_251,N_435);
or U566 (N_566,N_469,N_421);
nand U567 (N_567,N_232,N_400);
nor U568 (N_568,N_288,N_47);
and U569 (N_569,N_408,N_226);
nor U570 (N_570,N_94,N_463);
or U571 (N_571,N_246,N_454);
nor U572 (N_572,N_445,N_133);
nand U573 (N_573,N_32,N_399);
nand U574 (N_574,N_440,N_13);
xor U575 (N_575,N_144,N_154);
and U576 (N_576,N_424,N_7);
nand U577 (N_577,N_458,N_446);
and U578 (N_578,N_137,N_365);
and U579 (N_579,N_110,N_268);
or U580 (N_580,N_91,N_285);
nor U581 (N_581,N_150,N_491);
or U582 (N_582,N_284,N_339);
and U583 (N_583,N_359,N_102);
nand U584 (N_584,N_78,N_195);
nor U585 (N_585,N_120,N_74);
nand U586 (N_586,N_39,N_376);
or U587 (N_587,N_241,N_131);
nand U588 (N_588,N_302,N_33);
or U589 (N_589,N_308,N_130);
nor U590 (N_590,N_146,N_24);
nor U591 (N_591,N_386,N_389);
nand U592 (N_592,N_201,N_67);
or U593 (N_593,N_192,N_70);
nor U594 (N_594,N_84,N_111);
and U595 (N_595,N_444,N_206);
or U596 (N_596,N_304,N_20);
xnor U597 (N_597,N_387,N_449);
xor U598 (N_598,N_199,N_329);
nand U599 (N_599,N_101,N_300);
and U600 (N_600,N_340,N_197);
nand U601 (N_601,N_92,N_456);
nor U602 (N_602,N_58,N_416);
or U603 (N_603,N_65,N_166);
nand U604 (N_604,N_129,N_207);
nand U605 (N_605,N_158,N_263);
nand U606 (N_606,N_265,N_356);
and U607 (N_607,N_50,N_156);
xnor U608 (N_608,N_204,N_214);
xnor U609 (N_609,N_1,N_336);
nand U610 (N_610,N_355,N_198);
or U611 (N_611,N_72,N_279);
nand U612 (N_612,N_179,N_362);
nand U613 (N_613,N_34,N_160);
or U614 (N_614,N_116,N_305);
or U615 (N_615,N_222,N_167);
nor U616 (N_616,N_142,N_303);
nor U617 (N_617,N_295,N_97);
or U618 (N_618,N_447,N_12);
nand U619 (N_619,N_346,N_185);
nor U620 (N_620,N_320,N_377);
xor U621 (N_621,N_105,N_83);
or U622 (N_622,N_371,N_419);
xnor U623 (N_623,N_353,N_257);
and U624 (N_624,N_148,N_290);
nand U625 (N_625,N_219,N_465);
or U626 (N_626,N_169,N_53);
nor U627 (N_627,N_149,N_486);
nor U628 (N_628,N_68,N_488);
and U629 (N_629,N_405,N_46);
or U630 (N_630,N_347,N_471);
or U631 (N_631,N_461,N_373);
nor U632 (N_632,N_213,N_250);
and U633 (N_633,N_258,N_434);
nand U634 (N_634,N_138,N_431);
nor U635 (N_635,N_147,N_25);
and U636 (N_636,N_468,N_87);
nor U637 (N_637,N_100,N_253);
nand U638 (N_638,N_484,N_442);
nand U639 (N_639,N_483,N_19);
nand U640 (N_640,N_412,N_124);
or U641 (N_641,N_364,N_182);
nand U642 (N_642,N_441,N_443);
nor U643 (N_643,N_187,N_385);
or U644 (N_644,N_333,N_309);
and U645 (N_645,N_52,N_292);
and U646 (N_646,N_30,N_281);
or U647 (N_647,N_352,N_143);
nor U648 (N_648,N_242,N_109);
nor U649 (N_649,N_395,N_261);
nor U650 (N_650,N_127,N_145);
xor U651 (N_651,N_277,N_448);
nor U652 (N_652,N_205,N_452);
nor U653 (N_653,N_62,N_139);
and U654 (N_654,N_23,N_189);
or U655 (N_655,N_432,N_335);
xor U656 (N_656,N_374,N_259);
and U657 (N_657,N_173,N_267);
nor U658 (N_658,N_121,N_42);
nor U659 (N_659,N_254,N_3);
nor U660 (N_660,N_328,N_306);
nor U661 (N_661,N_455,N_0);
nor U662 (N_662,N_392,N_55);
or U663 (N_663,N_338,N_134);
nand U664 (N_664,N_489,N_252);
nor U665 (N_665,N_462,N_433);
or U666 (N_666,N_106,N_245);
nor U667 (N_667,N_480,N_270);
nor U668 (N_668,N_136,N_390);
xnor U669 (N_669,N_69,N_380);
and U670 (N_670,N_414,N_171);
or U671 (N_671,N_459,N_366);
or U672 (N_672,N_196,N_420);
nand U673 (N_673,N_117,N_56);
nor U674 (N_674,N_180,N_354);
nand U675 (N_675,N_425,N_191);
or U676 (N_676,N_90,N_439);
or U677 (N_677,N_282,N_337);
and U678 (N_678,N_240,N_475);
xnor U679 (N_679,N_312,N_236);
nor U680 (N_680,N_61,N_225);
nor U681 (N_681,N_368,N_170);
nor U682 (N_682,N_28,N_499);
nand U683 (N_683,N_244,N_193);
nand U684 (N_684,N_375,N_457);
or U685 (N_685,N_184,N_311);
nand U686 (N_686,N_357,N_476);
nand U687 (N_687,N_35,N_11);
nor U688 (N_688,N_108,N_161);
nand U689 (N_689,N_93,N_367);
nor U690 (N_690,N_274,N_118);
nor U691 (N_691,N_31,N_112);
and U692 (N_692,N_231,N_326);
or U693 (N_693,N_271,N_467);
or U694 (N_694,N_85,N_453);
nand U695 (N_695,N_209,N_264);
or U696 (N_696,N_114,N_478);
and U697 (N_697,N_349,N_410);
or U698 (N_698,N_430,N_317);
nor U699 (N_699,N_211,N_323);
nand U700 (N_700,N_125,N_299);
nor U701 (N_701,N_438,N_378);
nor U702 (N_702,N_162,N_212);
and U703 (N_703,N_104,N_176);
nor U704 (N_704,N_422,N_409);
xnor U705 (N_705,N_76,N_273);
or U706 (N_706,N_361,N_54);
nand U707 (N_707,N_71,N_89);
and U708 (N_708,N_341,N_481);
and U709 (N_709,N_415,N_10);
nor U710 (N_710,N_428,N_360);
nand U711 (N_711,N_8,N_234);
nor U712 (N_712,N_165,N_57);
nand U713 (N_713,N_99,N_383);
nand U714 (N_714,N_63,N_493);
or U715 (N_715,N_210,N_194);
nand U716 (N_716,N_485,N_382);
and U717 (N_717,N_426,N_64);
and U718 (N_718,N_490,N_177);
and U719 (N_719,N_45,N_397);
and U720 (N_720,N_81,N_393);
nand U721 (N_721,N_200,N_115);
nand U722 (N_722,N_163,N_496);
nor U723 (N_723,N_159,N_495);
or U724 (N_724,N_473,N_80);
and U725 (N_725,N_96,N_239);
and U726 (N_726,N_298,N_460);
nand U727 (N_727,N_322,N_26);
or U728 (N_728,N_470,N_464);
or U729 (N_729,N_381,N_423);
nand U730 (N_730,N_296,N_450);
and U731 (N_731,N_429,N_492);
nand U732 (N_732,N_151,N_237);
nor U733 (N_733,N_343,N_497);
and U734 (N_734,N_394,N_314);
nor U735 (N_735,N_59,N_330);
or U736 (N_736,N_325,N_334);
nor U737 (N_737,N_216,N_119);
and U738 (N_738,N_95,N_43);
and U739 (N_739,N_272,N_178);
xnor U740 (N_740,N_319,N_276);
nand U741 (N_741,N_123,N_472);
nand U742 (N_742,N_344,N_301);
nor U743 (N_743,N_135,N_350);
or U744 (N_744,N_451,N_402);
or U745 (N_745,N_404,N_103);
nand U746 (N_746,N_388,N_128);
nor U747 (N_747,N_310,N_4);
and U748 (N_748,N_348,N_174);
xnor U749 (N_749,N_48,N_255);
nor U750 (N_750,N_359,N_176);
or U751 (N_751,N_249,N_79);
or U752 (N_752,N_281,N_292);
nor U753 (N_753,N_392,N_336);
or U754 (N_754,N_440,N_344);
nor U755 (N_755,N_155,N_183);
nand U756 (N_756,N_122,N_265);
xnor U757 (N_757,N_497,N_439);
and U758 (N_758,N_141,N_209);
and U759 (N_759,N_221,N_408);
nand U760 (N_760,N_238,N_253);
and U761 (N_761,N_345,N_258);
and U762 (N_762,N_391,N_370);
or U763 (N_763,N_195,N_34);
nand U764 (N_764,N_188,N_257);
nand U765 (N_765,N_397,N_311);
and U766 (N_766,N_14,N_135);
nand U767 (N_767,N_110,N_116);
and U768 (N_768,N_274,N_147);
nor U769 (N_769,N_133,N_93);
or U770 (N_770,N_323,N_339);
nor U771 (N_771,N_464,N_174);
or U772 (N_772,N_122,N_135);
and U773 (N_773,N_257,N_179);
and U774 (N_774,N_34,N_1);
nor U775 (N_775,N_324,N_188);
or U776 (N_776,N_100,N_51);
nor U777 (N_777,N_172,N_400);
nand U778 (N_778,N_281,N_465);
nor U779 (N_779,N_54,N_84);
or U780 (N_780,N_138,N_4);
nor U781 (N_781,N_99,N_418);
or U782 (N_782,N_363,N_345);
or U783 (N_783,N_475,N_51);
nor U784 (N_784,N_320,N_288);
nor U785 (N_785,N_422,N_231);
nand U786 (N_786,N_23,N_413);
xnor U787 (N_787,N_350,N_149);
nor U788 (N_788,N_50,N_313);
and U789 (N_789,N_380,N_95);
or U790 (N_790,N_342,N_472);
or U791 (N_791,N_140,N_1);
nand U792 (N_792,N_258,N_290);
nor U793 (N_793,N_20,N_466);
nor U794 (N_794,N_371,N_328);
nor U795 (N_795,N_333,N_319);
nor U796 (N_796,N_492,N_463);
and U797 (N_797,N_490,N_238);
and U798 (N_798,N_177,N_239);
nor U799 (N_799,N_3,N_468);
nand U800 (N_800,N_487,N_235);
and U801 (N_801,N_411,N_167);
and U802 (N_802,N_332,N_164);
or U803 (N_803,N_455,N_374);
nand U804 (N_804,N_103,N_452);
nor U805 (N_805,N_167,N_497);
and U806 (N_806,N_211,N_443);
and U807 (N_807,N_307,N_169);
nor U808 (N_808,N_197,N_433);
or U809 (N_809,N_197,N_458);
xor U810 (N_810,N_130,N_205);
nand U811 (N_811,N_100,N_26);
nor U812 (N_812,N_162,N_301);
or U813 (N_813,N_119,N_39);
and U814 (N_814,N_39,N_456);
nand U815 (N_815,N_156,N_81);
nand U816 (N_816,N_70,N_446);
nor U817 (N_817,N_80,N_282);
xnor U818 (N_818,N_318,N_369);
or U819 (N_819,N_491,N_89);
or U820 (N_820,N_134,N_404);
or U821 (N_821,N_448,N_258);
and U822 (N_822,N_360,N_389);
and U823 (N_823,N_474,N_487);
and U824 (N_824,N_105,N_407);
nor U825 (N_825,N_285,N_151);
or U826 (N_826,N_44,N_437);
nor U827 (N_827,N_185,N_400);
xnor U828 (N_828,N_404,N_355);
or U829 (N_829,N_303,N_317);
nand U830 (N_830,N_354,N_358);
or U831 (N_831,N_368,N_258);
or U832 (N_832,N_398,N_101);
nor U833 (N_833,N_369,N_270);
nor U834 (N_834,N_411,N_206);
nand U835 (N_835,N_488,N_169);
and U836 (N_836,N_78,N_486);
nor U837 (N_837,N_345,N_332);
xor U838 (N_838,N_334,N_363);
and U839 (N_839,N_92,N_285);
and U840 (N_840,N_199,N_225);
xnor U841 (N_841,N_61,N_201);
nand U842 (N_842,N_466,N_145);
or U843 (N_843,N_490,N_170);
xnor U844 (N_844,N_233,N_231);
nand U845 (N_845,N_350,N_37);
nand U846 (N_846,N_171,N_415);
and U847 (N_847,N_445,N_373);
and U848 (N_848,N_196,N_344);
nor U849 (N_849,N_212,N_33);
nor U850 (N_850,N_431,N_242);
or U851 (N_851,N_67,N_300);
or U852 (N_852,N_454,N_457);
nand U853 (N_853,N_375,N_27);
and U854 (N_854,N_88,N_314);
and U855 (N_855,N_112,N_274);
nor U856 (N_856,N_59,N_76);
and U857 (N_857,N_250,N_348);
or U858 (N_858,N_347,N_294);
nor U859 (N_859,N_204,N_268);
nor U860 (N_860,N_294,N_239);
xnor U861 (N_861,N_493,N_426);
nand U862 (N_862,N_279,N_447);
nand U863 (N_863,N_162,N_195);
or U864 (N_864,N_481,N_350);
or U865 (N_865,N_197,N_324);
or U866 (N_866,N_267,N_303);
nor U867 (N_867,N_132,N_323);
or U868 (N_868,N_323,N_477);
nand U869 (N_869,N_175,N_1);
nand U870 (N_870,N_369,N_64);
nand U871 (N_871,N_497,N_58);
or U872 (N_872,N_380,N_345);
and U873 (N_873,N_207,N_488);
xor U874 (N_874,N_442,N_20);
nand U875 (N_875,N_115,N_114);
nor U876 (N_876,N_201,N_397);
nand U877 (N_877,N_27,N_410);
and U878 (N_878,N_311,N_250);
nor U879 (N_879,N_150,N_337);
xor U880 (N_880,N_345,N_181);
or U881 (N_881,N_397,N_82);
xor U882 (N_882,N_107,N_460);
and U883 (N_883,N_301,N_321);
xnor U884 (N_884,N_375,N_346);
nor U885 (N_885,N_334,N_215);
nor U886 (N_886,N_140,N_308);
or U887 (N_887,N_2,N_144);
nand U888 (N_888,N_328,N_247);
nand U889 (N_889,N_55,N_1);
nor U890 (N_890,N_475,N_337);
xnor U891 (N_891,N_308,N_121);
or U892 (N_892,N_0,N_423);
nor U893 (N_893,N_145,N_268);
or U894 (N_894,N_155,N_293);
and U895 (N_895,N_321,N_164);
or U896 (N_896,N_172,N_91);
nand U897 (N_897,N_165,N_275);
or U898 (N_898,N_50,N_405);
nor U899 (N_899,N_308,N_459);
nand U900 (N_900,N_344,N_336);
and U901 (N_901,N_292,N_458);
or U902 (N_902,N_94,N_310);
xor U903 (N_903,N_130,N_328);
nor U904 (N_904,N_136,N_244);
and U905 (N_905,N_332,N_241);
nand U906 (N_906,N_453,N_10);
or U907 (N_907,N_107,N_377);
or U908 (N_908,N_156,N_219);
or U909 (N_909,N_406,N_318);
nand U910 (N_910,N_298,N_34);
and U911 (N_911,N_26,N_72);
nor U912 (N_912,N_79,N_11);
and U913 (N_913,N_51,N_230);
or U914 (N_914,N_215,N_357);
and U915 (N_915,N_186,N_274);
nand U916 (N_916,N_405,N_378);
nor U917 (N_917,N_227,N_91);
nor U918 (N_918,N_45,N_372);
xor U919 (N_919,N_214,N_484);
nand U920 (N_920,N_306,N_240);
and U921 (N_921,N_17,N_162);
nand U922 (N_922,N_122,N_226);
nor U923 (N_923,N_261,N_403);
and U924 (N_924,N_319,N_387);
or U925 (N_925,N_427,N_491);
nor U926 (N_926,N_17,N_163);
nor U927 (N_927,N_397,N_12);
or U928 (N_928,N_483,N_394);
or U929 (N_929,N_414,N_193);
and U930 (N_930,N_310,N_261);
and U931 (N_931,N_496,N_433);
nor U932 (N_932,N_221,N_56);
and U933 (N_933,N_451,N_346);
and U934 (N_934,N_329,N_30);
or U935 (N_935,N_291,N_462);
xnor U936 (N_936,N_405,N_457);
and U937 (N_937,N_182,N_499);
or U938 (N_938,N_475,N_217);
nand U939 (N_939,N_35,N_129);
nand U940 (N_940,N_191,N_442);
nand U941 (N_941,N_493,N_119);
nand U942 (N_942,N_488,N_264);
and U943 (N_943,N_367,N_178);
and U944 (N_944,N_1,N_487);
or U945 (N_945,N_384,N_412);
nand U946 (N_946,N_467,N_281);
nor U947 (N_947,N_153,N_177);
xor U948 (N_948,N_294,N_188);
nand U949 (N_949,N_484,N_267);
and U950 (N_950,N_135,N_239);
or U951 (N_951,N_68,N_10);
xnor U952 (N_952,N_375,N_386);
nand U953 (N_953,N_407,N_70);
xor U954 (N_954,N_190,N_40);
or U955 (N_955,N_492,N_140);
nand U956 (N_956,N_246,N_13);
and U957 (N_957,N_187,N_435);
or U958 (N_958,N_366,N_31);
xor U959 (N_959,N_11,N_78);
or U960 (N_960,N_52,N_374);
nor U961 (N_961,N_79,N_42);
xor U962 (N_962,N_275,N_333);
and U963 (N_963,N_170,N_203);
xnor U964 (N_964,N_151,N_174);
or U965 (N_965,N_32,N_433);
or U966 (N_966,N_143,N_51);
nand U967 (N_967,N_113,N_200);
and U968 (N_968,N_397,N_63);
or U969 (N_969,N_66,N_150);
nor U970 (N_970,N_231,N_341);
and U971 (N_971,N_466,N_267);
nor U972 (N_972,N_146,N_145);
or U973 (N_973,N_420,N_3);
nor U974 (N_974,N_56,N_174);
nor U975 (N_975,N_437,N_264);
nand U976 (N_976,N_278,N_367);
nor U977 (N_977,N_100,N_28);
or U978 (N_978,N_480,N_106);
and U979 (N_979,N_328,N_56);
or U980 (N_980,N_403,N_127);
and U981 (N_981,N_199,N_298);
nor U982 (N_982,N_232,N_260);
or U983 (N_983,N_291,N_398);
or U984 (N_984,N_312,N_85);
or U985 (N_985,N_394,N_92);
nand U986 (N_986,N_417,N_341);
nor U987 (N_987,N_167,N_195);
or U988 (N_988,N_103,N_66);
and U989 (N_989,N_317,N_320);
nand U990 (N_990,N_111,N_460);
nor U991 (N_991,N_142,N_57);
nor U992 (N_992,N_276,N_376);
xor U993 (N_993,N_348,N_1);
xor U994 (N_994,N_491,N_141);
or U995 (N_995,N_280,N_235);
and U996 (N_996,N_62,N_484);
xor U997 (N_997,N_6,N_137);
nor U998 (N_998,N_320,N_249);
nor U999 (N_999,N_453,N_302);
and U1000 (N_1000,N_550,N_990);
or U1001 (N_1001,N_635,N_825);
or U1002 (N_1002,N_549,N_960);
or U1003 (N_1003,N_605,N_511);
nor U1004 (N_1004,N_848,N_526);
nor U1005 (N_1005,N_741,N_884);
or U1006 (N_1006,N_671,N_765);
nor U1007 (N_1007,N_650,N_963);
or U1008 (N_1008,N_573,N_629);
nand U1009 (N_1009,N_852,N_543);
and U1010 (N_1010,N_944,N_937);
or U1011 (N_1011,N_762,N_930);
nor U1012 (N_1012,N_870,N_844);
or U1013 (N_1013,N_767,N_538);
or U1014 (N_1014,N_782,N_875);
or U1015 (N_1015,N_789,N_598);
or U1016 (N_1016,N_522,N_745);
nand U1017 (N_1017,N_562,N_818);
nand U1018 (N_1018,N_524,N_828);
nor U1019 (N_1019,N_871,N_591);
or U1020 (N_1020,N_939,N_673);
or U1021 (N_1021,N_863,N_530);
and U1022 (N_1022,N_729,N_865);
and U1023 (N_1023,N_571,N_817);
nor U1024 (N_1024,N_560,N_839);
nand U1025 (N_1025,N_798,N_921);
or U1026 (N_1026,N_666,N_809);
xor U1027 (N_1027,N_730,N_862);
nor U1028 (N_1028,N_567,N_685);
or U1029 (N_1029,N_954,N_933);
nor U1030 (N_1030,N_754,N_904);
or U1031 (N_1031,N_647,N_945);
nand U1032 (N_1032,N_893,N_755);
nand U1033 (N_1033,N_634,N_531);
nand U1034 (N_1034,N_972,N_544);
or U1035 (N_1035,N_734,N_581);
nor U1036 (N_1036,N_689,N_829);
and U1037 (N_1037,N_508,N_514);
nand U1038 (N_1038,N_711,N_858);
or U1039 (N_1039,N_720,N_636);
xnor U1040 (N_1040,N_905,N_777);
or U1041 (N_1041,N_861,N_927);
or U1042 (N_1042,N_879,N_648);
nor U1043 (N_1043,N_616,N_715);
xnor U1044 (N_1044,N_780,N_796);
and U1045 (N_1045,N_620,N_743);
nand U1046 (N_1046,N_747,N_831);
xor U1047 (N_1047,N_646,N_947);
or U1048 (N_1048,N_942,N_710);
xnor U1049 (N_1049,N_984,N_955);
and U1050 (N_1050,N_696,N_682);
or U1051 (N_1051,N_702,N_769);
nor U1052 (N_1052,N_694,N_717);
and U1053 (N_1053,N_814,N_832);
or U1054 (N_1054,N_719,N_851);
and U1055 (N_1055,N_982,N_837);
or U1056 (N_1056,N_695,N_570);
and U1057 (N_1057,N_776,N_792);
and U1058 (N_1058,N_830,N_897);
nand U1059 (N_1059,N_811,N_768);
nand U1060 (N_1060,N_513,N_980);
nor U1061 (N_1061,N_838,N_759);
nand U1062 (N_1062,N_582,N_618);
or U1063 (N_1063,N_527,N_708);
and U1064 (N_1064,N_726,N_888);
nor U1065 (N_1065,N_516,N_592);
or U1066 (N_1066,N_662,N_894);
nand U1067 (N_1067,N_542,N_752);
or U1068 (N_1068,N_692,N_899);
nand U1069 (N_1069,N_709,N_775);
nand U1070 (N_1070,N_840,N_766);
or U1071 (N_1071,N_974,N_749);
or U1072 (N_1072,N_630,N_866);
nand U1073 (N_1073,N_928,N_608);
nor U1074 (N_1074,N_951,N_773);
nor U1075 (N_1075,N_908,N_533);
nand U1076 (N_1076,N_868,N_819);
or U1077 (N_1077,N_701,N_987);
and U1078 (N_1078,N_740,N_532);
nand U1079 (N_1079,N_900,N_691);
or U1080 (N_1080,N_800,N_949);
nand U1081 (N_1081,N_744,N_553);
nor U1082 (N_1082,N_523,N_845);
xor U1083 (N_1083,N_529,N_521);
nand U1084 (N_1084,N_609,N_574);
or U1085 (N_1085,N_751,N_907);
nand U1086 (N_1086,N_746,N_596);
and U1087 (N_1087,N_836,N_975);
nand U1088 (N_1088,N_654,N_753);
and U1089 (N_1089,N_995,N_727);
nand U1090 (N_1090,N_724,N_965);
and U1091 (N_1091,N_735,N_528);
nor U1092 (N_1092,N_756,N_916);
and U1093 (N_1093,N_507,N_610);
nor U1094 (N_1094,N_878,N_690);
or U1095 (N_1095,N_614,N_781);
nor U1096 (N_1096,N_989,N_812);
or U1097 (N_1097,N_834,N_577);
nand U1098 (N_1098,N_988,N_786);
nor U1099 (N_1099,N_737,N_505);
nor U1100 (N_1100,N_742,N_909);
nand U1101 (N_1101,N_968,N_827);
nand U1102 (N_1102,N_540,N_502);
nand U1103 (N_1103,N_892,N_669);
nand U1104 (N_1104,N_958,N_536);
and U1105 (N_1105,N_978,N_859);
and U1106 (N_1106,N_822,N_788);
and U1107 (N_1107,N_842,N_967);
nor U1108 (N_1108,N_889,N_625);
or U1109 (N_1109,N_597,N_804);
nand U1110 (N_1110,N_575,N_874);
and U1111 (N_1111,N_977,N_999);
nor U1112 (N_1112,N_552,N_733);
and U1113 (N_1113,N_760,N_813);
xor U1114 (N_1114,N_764,N_686);
and U1115 (N_1115,N_854,N_518);
and U1116 (N_1116,N_805,N_956);
nor U1117 (N_1117,N_551,N_566);
nand U1118 (N_1118,N_902,N_993);
or U1119 (N_1119,N_564,N_994);
or U1120 (N_1120,N_996,N_699);
and U1121 (N_1121,N_739,N_799);
or U1122 (N_1122,N_802,N_652);
nand U1123 (N_1123,N_664,N_821);
and U1124 (N_1124,N_801,N_912);
nor U1125 (N_1125,N_604,N_722);
nor U1126 (N_1126,N_590,N_816);
nor U1127 (N_1127,N_957,N_679);
and U1128 (N_1128,N_815,N_644);
and U1129 (N_1129,N_943,N_846);
nand U1130 (N_1130,N_932,N_563);
nor U1131 (N_1131,N_557,N_992);
and U1132 (N_1132,N_602,N_678);
or U1133 (N_1133,N_983,N_959);
nor U1134 (N_1134,N_847,N_661);
nand U1135 (N_1135,N_873,N_638);
nand U1136 (N_1136,N_774,N_898);
nand U1137 (N_1137,N_594,N_698);
nor U1138 (N_1138,N_856,N_503);
and U1139 (N_1139,N_855,N_642);
or U1140 (N_1140,N_643,N_510);
nor U1141 (N_1141,N_587,N_593);
nor U1142 (N_1142,N_535,N_895);
nor U1143 (N_1143,N_509,N_684);
nor U1144 (N_1144,N_504,N_672);
or U1145 (N_1145,N_639,N_785);
nor U1146 (N_1146,N_586,N_565);
or U1147 (N_1147,N_599,N_867);
or U1148 (N_1148,N_911,N_929);
and U1149 (N_1149,N_883,N_576);
nand U1150 (N_1150,N_890,N_946);
nor U1151 (N_1151,N_637,N_569);
xnor U1152 (N_1152,N_797,N_706);
or U1153 (N_1153,N_603,N_624);
or U1154 (N_1154,N_725,N_877);
or U1155 (N_1155,N_600,N_548);
and U1156 (N_1156,N_910,N_770);
xor U1157 (N_1157,N_833,N_934);
xor U1158 (N_1158,N_721,N_649);
and U1159 (N_1159,N_626,N_979);
or U1160 (N_1160,N_824,N_541);
or U1161 (N_1161,N_935,N_807);
nand U1162 (N_1162,N_501,N_918);
or U1163 (N_1163,N_948,N_880);
nand U1164 (N_1164,N_761,N_885);
nand U1165 (N_1165,N_619,N_941);
or U1166 (N_1166,N_559,N_525);
and U1167 (N_1167,N_876,N_869);
or U1168 (N_1168,N_860,N_731);
xnor U1169 (N_1169,N_962,N_519);
and U1170 (N_1170,N_580,N_903);
nor U1171 (N_1171,N_687,N_841);
nor U1172 (N_1172,N_683,N_655);
xnor U1173 (N_1173,N_633,N_906);
nand U1174 (N_1174,N_556,N_917);
xnor U1175 (N_1175,N_613,N_779);
and U1176 (N_1176,N_950,N_680);
or U1177 (N_1177,N_940,N_641);
nand U1178 (N_1178,N_640,N_793);
nor U1179 (N_1179,N_966,N_826);
nor U1180 (N_1180,N_808,N_969);
and U1181 (N_1181,N_707,N_668);
xor U1182 (N_1182,N_718,N_991);
or U1183 (N_1183,N_612,N_693);
and U1184 (N_1184,N_891,N_623);
and U1185 (N_1185,N_872,N_589);
nor U1186 (N_1186,N_645,N_539);
and U1187 (N_1187,N_938,N_506);
and U1188 (N_1188,N_843,N_772);
nor U1189 (N_1189,N_976,N_584);
nor U1190 (N_1190,N_611,N_723);
or U1191 (N_1191,N_728,N_627);
nor U1192 (N_1192,N_810,N_750);
or U1193 (N_1193,N_676,N_936);
or U1194 (N_1194,N_732,N_716);
nor U1195 (N_1195,N_546,N_500);
xor U1196 (N_1196,N_656,N_705);
xnor U1197 (N_1197,N_914,N_714);
xor U1198 (N_1198,N_926,N_585);
or U1199 (N_1199,N_607,N_632);
and U1200 (N_1200,N_628,N_881);
or U1201 (N_1201,N_738,N_558);
nor U1202 (N_1202,N_835,N_887);
nand U1203 (N_1203,N_981,N_771);
nor U1204 (N_1204,N_621,N_583);
or U1205 (N_1205,N_920,N_997);
or U1206 (N_1206,N_554,N_795);
nand U1207 (N_1207,N_665,N_806);
nor U1208 (N_1208,N_700,N_922);
xor U1209 (N_1209,N_675,N_515);
or U1210 (N_1210,N_667,N_663);
nand U1211 (N_1211,N_704,N_588);
and U1212 (N_1212,N_537,N_622);
or U1213 (N_1213,N_601,N_688);
and U1214 (N_1214,N_748,N_697);
nand U1215 (N_1215,N_657,N_713);
nand U1216 (N_1216,N_763,N_971);
and U1217 (N_1217,N_791,N_896);
and U1218 (N_1218,N_578,N_924);
or U1219 (N_1219,N_615,N_973);
nor U1220 (N_1220,N_986,N_998);
or U1221 (N_1221,N_555,N_849);
nand U1222 (N_1222,N_677,N_520);
nor U1223 (N_1223,N_545,N_595);
nor U1224 (N_1224,N_651,N_736);
nor U1225 (N_1225,N_961,N_964);
or U1226 (N_1226,N_790,N_953);
nor U1227 (N_1227,N_703,N_923);
nand U1228 (N_1228,N_561,N_617);
xor U1229 (N_1229,N_568,N_517);
nor U1230 (N_1230,N_534,N_512);
or U1231 (N_1231,N_915,N_659);
and U1232 (N_1232,N_547,N_925);
and U1233 (N_1233,N_787,N_712);
and U1234 (N_1234,N_572,N_784);
nand U1235 (N_1235,N_853,N_778);
or U1236 (N_1236,N_631,N_794);
nand U1237 (N_1237,N_886,N_820);
nand U1238 (N_1238,N_758,N_919);
nand U1239 (N_1239,N_913,N_783);
nor U1240 (N_1240,N_970,N_882);
and U1241 (N_1241,N_660,N_803);
nand U1242 (N_1242,N_658,N_681);
or U1243 (N_1243,N_952,N_864);
nand U1244 (N_1244,N_850,N_653);
nor U1245 (N_1245,N_931,N_757);
and U1246 (N_1246,N_823,N_579);
nor U1247 (N_1247,N_670,N_606);
and U1248 (N_1248,N_985,N_901);
nor U1249 (N_1249,N_857,N_674);
nor U1250 (N_1250,N_541,N_966);
or U1251 (N_1251,N_954,N_546);
or U1252 (N_1252,N_699,N_547);
nor U1253 (N_1253,N_578,N_660);
nor U1254 (N_1254,N_525,N_852);
or U1255 (N_1255,N_942,N_616);
or U1256 (N_1256,N_626,N_783);
nand U1257 (N_1257,N_756,N_558);
and U1258 (N_1258,N_723,N_911);
or U1259 (N_1259,N_502,N_831);
and U1260 (N_1260,N_994,N_512);
or U1261 (N_1261,N_870,N_699);
nand U1262 (N_1262,N_557,N_701);
nand U1263 (N_1263,N_946,N_721);
or U1264 (N_1264,N_547,N_926);
nor U1265 (N_1265,N_662,N_657);
and U1266 (N_1266,N_586,N_594);
and U1267 (N_1267,N_819,N_845);
nand U1268 (N_1268,N_879,N_502);
and U1269 (N_1269,N_904,N_854);
and U1270 (N_1270,N_692,N_562);
nor U1271 (N_1271,N_911,N_973);
or U1272 (N_1272,N_848,N_814);
nand U1273 (N_1273,N_750,N_984);
nand U1274 (N_1274,N_832,N_544);
and U1275 (N_1275,N_500,N_598);
or U1276 (N_1276,N_687,N_811);
or U1277 (N_1277,N_724,N_575);
nand U1278 (N_1278,N_647,N_574);
and U1279 (N_1279,N_787,N_655);
or U1280 (N_1280,N_784,N_833);
or U1281 (N_1281,N_625,N_822);
or U1282 (N_1282,N_851,N_581);
and U1283 (N_1283,N_800,N_592);
and U1284 (N_1284,N_618,N_810);
and U1285 (N_1285,N_830,N_516);
nand U1286 (N_1286,N_600,N_604);
and U1287 (N_1287,N_973,N_502);
nand U1288 (N_1288,N_915,N_541);
nor U1289 (N_1289,N_773,N_898);
or U1290 (N_1290,N_703,N_506);
nor U1291 (N_1291,N_820,N_798);
or U1292 (N_1292,N_659,N_874);
xor U1293 (N_1293,N_547,N_863);
xor U1294 (N_1294,N_730,N_838);
nand U1295 (N_1295,N_528,N_810);
xnor U1296 (N_1296,N_828,N_814);
and U1297 (N_1297,N_685,N_643);
xnor U1298 (N_1298,N_506,N_658);
or U1299 (N_1299,N_772,N_560);
nand U1300 (N_1300,N_916,N_788);
nor U1301 (N_1301,N_863,N_612);
nor U1302 (N_1302,N_537,N_739);
nor U1303 (N_1303,N_776,N_570);
nor U1304 (N_1304,N_803,N_829);
nor U1305 (N_1305,N_594,N_992);
and U1306 (N_1306,N_916,N_691);
nand U1307 (N_1307,N_813,N_928);
or U1308 (N_1308,N_809,N_827);
or U1309 (N_1309,N_563,N_994);
xor U1310 (N_1310,N_861,N_937);
and U1311 (N_1311,N_646,N_568);
and U1312 (N_1312,N_699,N_924);
nand U1313 (N_1313,N_606,N_581);
or U1314 (N_1314,N_788,N_852);
nor U1315 (N_1315,N_915,N_534);
nand U1316 (N_1316,N_885,N_844);
nor U1317 (N_1317,N_995,N_554);
nor U1318 (N_1318,N_517,N_673);
nand U1319 (N_1319,N_763,N_585);
nand U1320 (N_1320,N_913,N_555);
and U1321 (N_1321,N_759,N_886);
nand U1322 (N_1322,N_671,N_998);
or U1323 (N_1323,N_976,N_725);
nand U1324 (N_1324,N_812,N_665);
or U1325 (N_1325,N_635,N_555);
nand U1326 (N_1326,N_597,N_518);
and U1327 (N_1327,N_594,N_890);
nand U1328 (N_1328,N_630,N_706);
or U1329 (N_1329,N_990,N_630);
or U1330 (N_1330,N_501,N_948);
nor U1331 (N_1331,N_964,N_850);
and U1332 (N_1332,N_508,N_794);
nor U1333 (N_1333,N_949,N_802);
or U1334 (N_1334,N_691,N_919);
nor U1335 (N_1335,N_716,N_674);
or U1336 (N_1336,N_741,N_645);
or U1337 (N_1337,N_905,N_579);
xnor U1338 (N_1338,N_672,N_767);
xnor U1339 (N_1339,N_921,N_945);
or U1340 (N_1340,N_622,N_617);
nand U1341 (N_1341,N_944,N_856);
and U1342 (N_1342,N_805,N_577);
or U1343 (N_1343,N_588,N_974);
nor U1344 (N_1344,N_602,N_740);
nand U1345 (N_1345,N_721,N_821);
or U1346 (N_1346,N_838,N_608);
and U1347 (N_1347,N_975,N_605);
nor U1348 (N_1348,N_961,N_877);
nor U1349 (N_1349,N_620,N_966);
nand U1350 (N_1350,N_857,N_791);
nand U1351 (N_1351,N_735,N_581);
xor U1352 (N_1352,N_953,N_523);
xor U1353 (N_1353,N_629,N_772);
nand U1354 (N_1354,N_687,N_897);
nor U1355 (N_1355,N_760,N_872);
or U1356 (N_1356,N_888,N_724);
nand U1357 (N_1357,N_663,N_556);
and U1358 (N_1358,N_513,N_604);
and U1359 (N_1359,N_749,N_946);
or U1360 (N_1360,N_573,N_634);
nand U1361 (N_1361,N_733,N_806);
and U1362 (N_1362,N_777,N_731);
nand U1363 (N_1363,N_850,N_766);
nand U1364 (N_1364,N_849,N_641);
and U1365 (N_1365,N_759,N_870);
nand U1366 (N_1366,N_744,N_770);
and U1367 (N_1367,N_517,N_860);
or U1368 (N_1368,N_814,N_757);
nor U1369 (N_1369,N_583,N_624);
nor U1370 (N_1370,N_892,N_825);
nand U1371 (N_1371,N_614,N_624);
nand U1372 (N_1372,N_530,N_775);
xor U1373 (N_1373,N_527,N_552);
and U1374 (N_1374,N_600,N_738);
nor U1375 (N_1375,N_529,N_572);
nor U1376 (N_1376,N_883,N_591);
and U1377 (N_1377,N_972,N_859);
nor U1378 (N_1378,N_827,N_609);
and U1379 (N_1379,N_894,N_691);
nor U1380 (N_1380,N_825,N_649);
or U1381 (N_1381,N_908,N_701);
nand U1382 (N_1382,N_787,N_819);
nand U1383 (N_1383,N_600,N_871);
nor U1384 (N_1384,N_552,N_730);
nand U1385 (N_1385,N_813,N_575);
and U1386 (N_1386,N_715,N_997);
nand U1387 (N_1387,N_875,N_565);
xnor U1388 (N_1388,N_581,N_509);
nand U1389 (N_1389,N_770,N_811);
nand U1390 (N_1390,N_798,N_598);
xnor U1391 (N_1391,N_818,N_994);
and U1392 (N_1392,N_769,N_571);
and U1393 (N_1393,N_828,N_742);
xnor U1394 (N_1394,N_629,N_807);
nor U1395 (N_1395,N_646,N_642);
nand U1396 (N_1396,N_816,N_713);
or U1397 (N_1397,N_711,N_714);
nand U1398 (N_1398,N_618,N_654);
xnor U1399 (N_1399,N_593,N_531);
nand U1400 (N_1400,N_575,N_797);
nand U1401 (N_1401,N_606,N_911);
and U1402 (N_1402,N_825,N_773);
nor U1403 (N_1403,N_521,N_852);
xor U1404 (N_1404,N_551,N_735);
xor U1405 (N_1405,N_915,N_765);
nand U1406 (N_1406,N_603,N_600);
or U1407 (N_1407,N_518,N_558);
and U1408 (N_1408,N_612,N_653);
or U1409 (N_1409,N_790,N_973);
nor U1410 (N_1410,N_597,N_800);
xor U1411 (N_1411,N_936,N_500);
nand U1412 (N_1412,N_992,N_928);
nand U1413 (N_1413,N_705,N_842);
or U1414 (N_1414,N_546,N_801);
nand U1415 (N_1415,N_910,N_585);
or U1416 (N_1416,N_737,N_722);
and U1417 (N_1417,N_676,N_723);
or U1418 (N_1418,N_602,N_832);
nor U1419 (N_1419,N_756,N_507);
nand U1420 (N_1420,N_747,N_984);
and U1421 (N_1421,N_926,N_548);
nor U1422 (N_1422,N_981,N_744);
or U1423 (N_1423,N_561,N_669);
or U1424 (N_1424,N_519,N_622);
nand U1425 (N_1425,N_731,N_896);
nand U1426 (N_1426,N_808,N_662);
xor U1427 (N_1427,N_855,N_702);
nand U1428 (N_1428,N_675,N_501);
nor U1429 (N_1429,N_878,N_665);
nand U1430 (N_1430,N_863,N_875);
nor U1431 (N_1431,N_636,N_740);
or U1432 (N_1432,N_681,N_981);
or U1433 (N_1433,N_606,N_985);
nand U1434 (N_1434,N_898,N_918);
or U1435 (N_1435,N_553,N_873);
nand U1436 (N_1436,N_796,N_630);
and U1437 (N_1437,N_711,N_981);
xnor U1438 (N_1438,N_994,N_524);
or U1439 (N_1439,N_891,N_930);
or U1440 (N_1440,N_760,N_730);
nor U1441 (N_1441,N_793,N_977);
and U1442 (N_1442,N_952,N_873);
and U1443 (N_1443,N_963,N_574);
or U1444 (N_1444,N_820,N_702);
nor U1445 (N_1445,N_816,N_605);
nor U1446 (N_1446,N_985,N_910);
and U1447 (N_1447,N_758,N_910);
nand U1448 (N_1448,N_505,N_864);
and U1449 (N_1449,N_677,N_527);
nor U1450 (N_1450,N_805,N_638);
or U1451 (N_1451,N_657,N_721);
nor U1452 (N_1452,N_527,N_931);
or U1453 (N_1453,N_977,N_501);
or U1454 (N_1454,N_506,N_604);
nor U1455 (N_1455,N_558,N_616);
xnor U1456 (N_1456,N_698,N_976);
nand U1457 (N_1457,N_863,N_722);
and U1458 (N_1458,N_506,N_983);
nand U1459 (N_1459,N_993,N_842);
or U1460 (N_1460,N_734,N_941);
or U1461 (N_1461,N_959,N_964);
nand U1462 (N_1462,N_809,N_677);
and U1463 (N_1463,N_926,N_601);
xor U1464 (N_1464,N_683,N_951);
xnor U1465 (N_1465,N_871,N_522);
nand U1466 (N_1466,N_838,N_892);
and U1467 (N_1467,N_878,N_833);
nand U1468 (N_1468,N_971,N_656);
or U1469 (N_1469,N_619,N_704);
or U1470 (N_1470,N_717,N_984);
nand U1471 (N_1471,N_977,N_693);
nand U1472 (N_1472,N_867,N_633);
or U1473 (N_1473,N_793,N_934);
or U1474 (N_1474,N_872,N_633);
and U1475 (N_1475,N_757,N_628);
or U1476 (N_1476,N_790,N_626);
and U1477 (N_1477,N_828,N_634);
nor U1478 (N_1478,N_588,N_862);
nor U1479 (N_1479,N_628,N_736);
nand U1480 (N_1480,N_920,N_642);
nand U1481 (N_1481,N_840,N_939);
or U1482 (N_1482,N_746,N_553);
or U1483 (N_1483,N_823,N_641);
nor U1484 (N_1484,N_995,N_736);
or U1485 (N_1485,N_801,N_971);
nor U1486 (N_1486,N_727,N_524);
nor U1487 (N_1487,N_663,N_501);
nand U1488 (N_1488,N_724,N_763);
nor U1489 (N_1489,N_508,N_580);
or U1490 (N_1490,N_635,N_904);
nor U1491 (N_1491,N_756,N_929);
nand U1492 (N_1492,N_868,N_762);
or U1493 (N_1493,N_799,N_883);
or U1494 (N_1494,N_804,N_671);
or U1495 (N_1495,N_636,N_736);
nor U1496 (N_1496,N_654,N_504);
nand U1497 (N_1497,N_824,N_749);
and U1498 (N_1498,N_826,N_748);
nand U1499 (N_1499,N_915,N_503);
or U1500 (N_1500,N_1247,N_1334);
or U1501 (N_1501,N_1387,N_1228);
or U1502 (N_1502,N_1490,N_1158);
nand U1503 (N_1503,N_1224,N_1100);
and U1504 (N_1504,N_1260,N_1036);
nand U1505 (N_1505,N_1434,N_1453);
and U1506 (N_1506,N_1337,N_1383);
or U1507 (N_1507,N_1327,N_1249);
or U1508 (N_1508,N_1390,N_1190);
or U1509 (N_1509,N_1465,N_1317);
nor U1510 (N_1510,N_1478,N_1369);
and U1511 (N_1511,N_1172,N_1042);
and U1512 (N_1512,N_1410,N_1267);
nor U1513 (N_1513,N_1041,N_1002);
nor U1514 (N_1514,N_1236,N_1424);
or U1515 (N_1515,N_1215,N_1365);
or U1516 (N_1516,N_1229,N_1213);
and U1517 (N_1517,N_1026,N_1308);
and U1518 (N_1518,N_1310,N_1051);
nand U1519 (N_1519,N_1094,N_1354);
nand U1520 (N_1520,N_1340,N_1281);
and U1521 (N_1521,N_1148,N_1070);
and U1522 (N_1522,N_1117,N_1014);
and U1523 (N_1523,N_1018,N_1336);
and U1524 (N_1524,N_1198,N_1149);
nor U1525 (N_1525,N_1031,N_1353);
or U1526 (N_1526,N_1009,N_1399);
nor U1527 (N_1527,N_1345,N_1450);
or U1528 (N_1528,N_1167,N_1015);
and U1529 (N_1529,N_1174,N_1253);
or U1530 (N_1530,N_1451,N_1201);
nor U1531 (N_1531,N_1222,N_1409);
nand U1532 (N_1532,N_1344,N_1211);
nor U1533 (N_1533,N_1244,N_1072);
or U1534 (N_1534,N_1087,N_1164);
and U1535 (N_1535,N_1494,N_1357);
or U1536 (N_1536,N_1062,N_1420);
or U1537 (N_1537,N_1426,N_1169);
and U1538 (N_1538,N_1126,N_1292);
xor U1539 (N_1539,N_1343,N_1056);
nand U1540 (N_1540,N_1135,N_1032);
nand U1541 (N_1541,N_1103,N_1485);
and U1542 (N_1542,N_1279,N_1077);
nand U1543 (N_1543,N_1256,N_1379);
nand U1544 (N_1544,N_1181,N_1455);
nand U1545 (N_1545,N_1199,N_1367);
nand U1546 (N_1546,N_1024,N_1444);
and U1547 (N_1547,N_1276,N_1205);
or U1548 (N_1548,N_1239,N_1075);
or U1549 (N_1549,N_1161,N_1411);
and U1550 (N_1550,N_1227,N_1449);
xor U1551 (N_1551,N_1145,N_1347);
or U1552 (N_1552,N_1315,N_1218);
and U1553 (N_1553,N_1309,N_1432);
nor U1554 (N_1554,N_1303,N_1293);
and U1555 (N_1555,N_1074,N_1484);
nand U1556 (N_1556,N_1392,N_1150);
nor U1557 (N_1557,N_1132,N_1003);
or U1558 (N_1558,N_1417,N_1352);
and U1559 (N_1559,N_1361,N_1155);
and U1560 (N_1560,N_1333,N_1127);
or U1561 (N_1561,N_1427,N_1243);
and U1562 (N_1562,N_1023,N_1391);
nor U1563 (N_1563,N_1439,N_1382);
nand U1564 (N_1564,N_1288,N_1186);
nor U1565 (N_1565,N_1405,N_1498);
nand U1566 (N_1566,N_1324,N_1095);
nand U1567 (N_1567,N_1375,N_1445);
nor U1568 (N_1568,N_1396,N_1129);
and U1569 (N_1569,N_1082,N_1266);
nand U1570 (N_1570,N_1318,N_1313);
or U1571 (N_1571,N_1143,N_1097);
nor U1572 (N_1572,N_1008,N_1322);
nand U1573 (N_1573,N_1049,N_1269);
nand U1574 (N_1574,N_1136,N_1170);
nand U1575 (N_1575,N_1338,N_1294);
or U1576 (N_1576,N_1221,N_1487);
xnor U1577 (N_1577,N_1177,N_1217);
and U1578 (N_1578,N_1251,N_1299);
nor U1579 (N_1579,N_1089,N_1054);
or U1580 (N_1580,N_1027,N_1080);
nor U1581 (N_1581,N_1055,N_1330);
nand U1582 (N_1582,N_1246,N_1374);
or U1583 (N_1583,N_1028,N_1109);
nor U1584 (N_1584,N_1316,N_1389);
nor U1585 (N_1585,N_1098,N_1402);
nand U1586 (N_1586,N_1335,N_1168);
nor U1587 (N_1587,N_1182,N_1438);
nor U1588 (N_1588,N_1372,N_1339);
nand U1589 (N_1589,N_1386,N_1033);
nor U1590 (N_1590,N_1096,N_1187);
nand U1591 (N_1591,N_1297,N_1452);
nor U1592 (N_1592,N_1433,N_1195);
or U1593 (N_1593,N_1472,N_1464);
nand U1594 (N_1594,N_1423,N_1066);
and U1595 (N_1595,N_1004,N_1306);
nand U1596 (N_1596,N_1131,N_1348);
and U1597 (N_1597,N_1346,N_1084);
nand U1598 (N_1598,N_1151,N_1202);
and U1599 (N_1599,N_1377,N_1425);
nand U1600 (N_1600,N_1064,N_1270);
and U1601 (N_1601,N_1265,N_1192);
or U1602 (N_1602,N_1111,N_1466);
nand U1603 (N_1603,N_1471,N_1441);
and U1604 (N_1604,N_1406,N_1285);
and U1605 (N_1605,N_1404,N_1370);
or U1606 (N_1606,N_1255,N_1144);
nor U1607 (N_1607,N_1025,N_1063);
nor U1608 (N_1608,N_1130,N_1488);
nor U1609 (N_1609,N_1262,N_1289);
or U1610 (N_1610,N_1314,N_1457);
xor U1611 (N_1611,N_1291,N_1312);
or U1612 (N_1612,N_1469,N_1007);
nand U1613 (N_1613,N_1416,N_1044);
nand U1614 (N_1614,N_1180,N_1016);
nand U1615 (N_1615,N_1319,N_1108);
and U1616 (N_1616,N_1173,N_1152);
nor U1617 (N_1617,N_1238,N_1088);
or U1618 (N_1618,N_1364,N_1491);
nand U1619 (N_1619,N_1142,N_1477);
or U1620 (N_1620,N_1107,N_1325);
or U1621 (N_1621,N_1006,N_1017);
and U1622 (N_1622,N_1429,N_1278);
nand U1623 (N_1623,N_1263,N_1418);
nand U1624 (N_1624,N_1153,N_1081);
nor U1625 (N_1625,N_1329,N_1000);
nand U1626 (N_1626,N_1124,N_1384);
nor U1627 (N_1627,N_1073,N_1493);
xnor U1628 (N_1628,N_1298,N_1323);
nor U1629 (N_1629,N_1388,N_1101);
and U1630 (N_1630,N_1092,N_1400);
nor U1631 (N_1631,N_1385,N_1250);
nor U1632 (N_1632,N_1414,N_1118);
nor U1633 (N_1633,N_1476,N_1280);
nand U1634 (N_1634,N_1133,N_1245);
nand U1635 (N_1635,N_1012,N_1110);
or U1636 (N_1636,N_1286,N_1138);
and U1637 (N_1637,N_1059,N_1301);
xnor U1638 (N_1638,N_1436,N_1373);
nand U1639 (N_1639,N_1496,N_1480);
nor U1640 (N_1640,N_1380,N_1102);
and U1641 (N_1641,N_1394,N_1328);
or U1642 (N_1642,N_1296,N_1210);
or U1643 (N_1643,N_1483,N_1001);
and U1644 (N_1644,N_1401,N_1235);
nor U1645 (N_1645,N_1034,N_1204);
xor U1646 (N_1646,N_1035,N_1159);
and U1647 (N_1647,N_1460,N_1165);
or U1648 (N_1648,N_1259,N_1492);
xor U1649 (N_1649,N_1290,N_1068);
and U1650 (N_1650,N_1234,N_1381);
or U1651 (N_1651,N_1456,N_1219);
or U1652 (N_1652,N_1171,N_1470);
nand U1653 (N_1653,N_1178,N_1112);
nand U1654 (N_1654,N_1359,N_1311);
nand U1655 (N_1655,N_1185,N_1341);
xor U1656 (N_1656,N_1079,N_1175);
nand U1657 (N_1657,N_1368,N_1115);
and U1658 (N_1658,N_1057,N_1331);
nand U1659 (N_1659,N_1355,N_1120);
nand U1660 (N_1660,N_1093,N_1099);
nand U1661 (N_1661,N_1113,N_1189);
or U1662 (N_1662,N_1021,N_1209);
nand U1663 (N_1663,N_1304,N_1162);
and U1664 (N_1664,N_1226,N_1086);
nor U1665 (N_1665,N_1040,N_1156);
or U1666 (N_1666,N_1157,N_1408);
xnor U1667 (N_1667,N_1214,N_1067);
nor U1668 (N_1668,N_1200,N_1240);
nand U1669 (N_1669,N_1078,N_1196);
or U1670 (N_1670,N_1065,N_1443);
and U1671 (N_1671,N_1123,N_1085);
nand U1672 (N_1672,N_1011,N_1119);
or U1673 (N_1673,N_1043,N_1128);
nand U1674 (N_1674,N_1479,N_1154);
or U1675 (N_1675,N_1020,N_1038);
nor U1676 (N_1676,N_1287,N_1447);
nand U1677 (N_1677,N_1203,N_1258);
or U1678 (N_1678,N_1497,N_1378);
or U1679 (N_1679,N_1275,N_1448);
and U1680 (N_1680,N_1431,N_1242);
or U1681 (N_1681,N_1030,N_1212);
or U1682 (N_1682,N_1489,N_1282);
nand U1683 (N_1683,N_1468,N_1366);
nand U1684 (N_1684,N_1274,N_1223);
and U1685 (N_1685,N_1332,N_1273);
xnor U1686 (N_1686,N_1179,N_1069);
nor U1687 (N_1687,N_1362,N_1305);
xor U1688 (N_1688,N_1398,N_1295);
nand U1689 (N_1689,N_1300,N_1252);
nand U1690 (N_1690,N_1013,N_1428);
and U1691 (N_1691,N_1039,N_1125);
nand U1692 (N_1692,N_1183,N_1166);
and U1693 (N_1693,N_1397,N_1220);
nor U1694 (N_1694,N_1422,N_1045);
xnor U1695 (N_1695,N_1261,N_1019);
xnor U1696 (N_1696,N_1415,N_1283);
or U1697 (N_1697,N_1349,N_1358);
and U1698 (N_1698,N_1454,N_1277);
nand U1699 (N_1699,N_1499,N_1421);
nand U1700 (N_1700,N_1351,N_1005);
nor U1701 (N_1701,N_1114,N_1430);
or U1702 (N_1702,N_1463,N_1393);
nor U1703 (N_1703,N_1412,N_1495);
nand U1704 (N_1704,N_1116,N_1264);
and U1705 (N_1705,N_1474,N_1473);
nor U1706 (N_1706,N_1241,N_1232);
xnor U1707 (N_1707,N_1284,N_1083);
or U1708 (N_1708,N_1435,N_1121);
nor U1709 (N_1709,N_1350,N_1395);
nand U1710 (N_1710,N_1053,N_1207);
or U1711 (N_1711,N_1486,N_1176);
nor U1712 (N_1712,N_1147,N_1482);
nand U1713 (N_1713,N_1104,N_1307);
or U1714 (N_1714,N_1225,N_1140);
and U1715 (N_1715,N_1022,N_1440);
nor U1716 (N_1716,N_1419,N_1231);
nor U1717 (N_1717,N_1481,N_1091);
and U1718 (N_1718,N_1271,N_1403);
xor U1719 (N_1719,N_1320,N_1050);
or U1720 (N_1720,N_1141,N_1254);
nor U1721 (N_1721,N_1060,N_1467);
and U1722 (N_1722,N_1446,N_1326);
nand U1723 (N_1723,N_1052,N_1188);
and U1724 (N_1724,N_1193,N_1010);
or U1725 (N_1725,N_1090,N_1237);
and U1726 (N_1726,N_1413,N_1137);
xnor U1727 (N_1727,N_1106,N_1139);
and U1728 (N_1728,N_1363,N_1191);
and U1729 (N_1729,N_1230,N_1134);
and U1730 (N_1730,N_1376,N_1216);
nand U1731 (N_1731,N_1047,N_1029);
or U1732 (N_1732,N_1321,N_1046);
or U1733 (N_1733,N_1268,N_1461);
or U1734 (N_1734,N_1233,N_1356);
or U1735 (N_1735,N_1037,N_1071);
nand U1736 (N_1736,N_1462,N_1197);
nor U1737 (N_1737,N_1371,N_1194);
nand U1738 (N_1738,N_1122,N_1342);
nor U1739 (N_1739,N_1302,N_1061);
nor U1740 (N_1740,N_1248,N_1206);
or U1741 (N_1741,N_1360,N_1272);
nand U1742 (N_1742,N_1163,N_1076);
nor U1743 (N_1743,N_1160,N_1458);
and U1744 (N_1744,N_1257,N_1184);
nand U1745 (N_1745,N_1437,N_1442);
or U1746 (N_1746,N_1459,N_1208);
or U1747 (N_1747,N_1058,N_1407);
nand U1748 (N_1748,N_1475,N_1146);
or U1749 (N_1749,N_1105,N_1048);
or U1750 (N_1750,N_1302,N_1176);
or U1751 (N_1751,N_1062,N_1303);
and U1752 (N_1752,N_1451,N_1047);
nor U1753 (N_1753,N_1462,N_1332);
nor U1754 (N_1754,N_1012,N_1262);
nor U1755 (N_1755,N_1032,N_1241);
and U1756 (N_1756,N_1380,N_1103);
nor U1757 (N_1757,N_1499,N_1049);
nand U1758 (N_1758,N_1344,N_1135);
and U1759 (N_1759,N_1406,N_1328);
nor U1760 (N_1760,N_1396,N_1190);
nand U1761 (N_1761,N_1276,N_1458);
nand U1762 (N_1762,N_1208,N_1138);
or U1763 (N_1763,N_1151,N_1416);
nand U1764 (N_1764,N_1416,N_1144);
nor U1765 (N_1765,N_1252,N_1402);
nor U1766 (N_1766,N_1413,N_1187);
nor U1767 (N_1767,N_1098,N_1168);
nand U1768 (N_1768,N_1059,N_1164);
or U1769 (N_1769,N_1166,N_1011);
nand U1770 (N_1770,N_1341,N_1299);
or U1771 (N_1771,N_1497,N_1253);
and U1772 (N_1772,N_1211,N_1339);
and U1773 (N_1773,N_1348,N_1005);
or U1774 (N_1774,N_1300,N_1316);
nand U1775 (N_1775,N_1185,N_1118);
xor U1776 (N_1776,N_1309,N_1279);
xnor U1777 (N_1777,N_1458,N_1400);
and U1778 (N_1778,N_1083,N_1293);
nor U1779 (N_1779,N_1472,N_1450);
and U1780 (N_1780,N_1244,N_1031);
and U1781 (N_1781,N_1496,N_1080);
or U1782 (N_1782,N_1275,N_1268);
or U1783 (N_1783,N_1200,N_1414);
or U1784 (N_1784,N_1019,N_1396);
nor U1785 (N_1785,N_1354,N_1451);
nand U1786 (N_1786,N_1428,N_1219);
and U1787 (N_1787,N_1275,N_1182);
nand U1788 (N_1788,N_1254,N_1271);
and U1789 (N_1789,N_1087,N_1021);
nand U1790 (N_1790,N_1255,N_1182);
nand U1791 (N_1791,N_1127,N_1354);
and U1792 (N_1792,N_1321,N_1409);
or U1793 (N_1793,N_1273,N_1090);
nor U1794 (N_1794,N_1246,N_1191);
nand U1795 (N_1795,N_1461,N_1171);
nor U1796 (N_1796,N_1335,N_1175);
xnor U1797 (N_1797,N_1211,N_1296);
or U1798 (N_1798,N_1288,N_1462);
and U1799 (N_1799,N_1051,N_1249);
and U1800 (N_1800,N_1290,N_1255);
nor U1801 (N_1801,N_1140,N_1158);
or U1802 (N_1802,N_1088,N_1347);
nand U1803 (N_1803,N_1272,N_1133);
xnor U1804 (N_1804,N_1475,N_1190);
or U1805 (N_1805,N_1182,N_1337);
and U1806 (N_1806,N_1182,N_1450);
or U1807 (N_1807,N_1447,N_1040);
and U1808 (N_1808,N_1253,N_1388);
or U1809 (N_1809,N_1058,N_1254);
and U1810 (N_1810,N_1118,N_1423);
and U1811 (N_1811,N_1306,N_1033);
nand U1812 (N_1812,N_1369,N_1197);
and U1813 (N_1813,N_1315,N_1338);
or U1814 (N_1814,N_1275,N_1342);
nor U1815 (N_1815,N_1461,N_1066);
nor U1816 (N_1816,N_1260,N_1499);
xnor U1817 (N_1817,N_1160,N_1092);
nor U1818 (N_1818,N_1459,N_1284);
nand U1819 (N_1819,N_1229,N_1367);
nand U1820 (N_1820,N_1164,N_1260);
nand U1821 (N_1821,N_1380,N_1224);
nor U1822 (N_1822,N_1428,N_1327);
and U1823 (N_1823,N_1386,N_1129);
xor U1824 (N_1824,N_1061,N_1173);
or U1825 (N_1825,N_1449,N_1319);
nor U1826 (N_1826,N_1465,N_1276);
xor U1827 (N_1827,N_1092,N_1246);
nor U1828 (N_1828,N_1025,N_1415);
nor U1829 (N_1829,N_1398,N_1148);
or U1830 (N_1830,N_1307,N_1435);
and U1831 (N_1831,N_1373,N_1163);
or U1832 (N_1832,N_1452,N_1227);
and U1833 (N_1833,N_1117,N_1185);
xor U1834 (N_1834,N_1488,N_1460);
xor U1835 (N_1835,N_1396,N_1380);
and U1836 (N_1836,N_1485,N_1080);
or U1837 (N_1837,N_1141,N_1268);
nand U1838 (N_1838,N_1338,N_1326);
nand U1839 (N_1839,N_1078,N_1333);
and U1840 (N_1840,N_1118,N_1074);
nand U1841 (N_1841,N_1234,N_1207);
and U1842 (N_1842,N_1493,N_1174);
nor U1843 (N_1843,N_1396,N_1164);
and U1844 (N_1844,N_1313,N_1215);
xor U1845 (N_1845,N_1096,N_1125);
nand U1846 (N_1846,N_1122,N_1030);
or U1847 (N_1847,N_1151,N_1362);
nand U1848 (N_1848,N_1335,N_1045);
and U1849 (N_1849,N_1038,N_1004);
and U1850 (N_1850,N_1178,N_1002);
nor U1851 (N_1851,N_1258,N_1015);
or U1852 (N_1852,N_1321,N_1431);
and U1853 (N_1853,N_1355,N_1301);
xor U1854 (N_1854,N_1210,N_1274);
nor U1855 (N_1855,N_1238,N_1001);
nor U1856 (N_1856,N_1056,N_1374);
nor U1857 (N_1857,N_1404,N_1264);
xnor U1858 (N_1858,N_1354,N_1138);
or U1859 (N_1859,N_1012,N_1293);
xor U1860 (N_1860,N_1445,N_1457);
or U1861 (N_1861,N_1184,N_1338);
nand U1862 (N_1862,N_1306,N_1133);
nor U1863 (N_1863,N_1140,N_1289);
nand U1864 (N_1864,N_1041,N_1390);
nor U1865 (N_1865,N_1468,N_1297);
nand U1866 (N_1866,N_1182,N_1204);
and U1867 (N_1867,N_1442,N_1475);
nor U1868 (N_1868,N_1151,N_1192);
nand U1869 (N_1869,N_1390,N_1155);
nand U1870 (N_1870,N_1336,N_1061);
nand U1871 (N_1871,N_1048,N_1431);
or U1872 (N_1872,N_1105,N_1015);
nor U1873 (N_1873,N_1199,N_1455);
and U1874 (N_1874,N_1421,N_1331);
and U1875 (N_1875,N_1351,N_1107);
or U1876 (N_1876,N_1174,N_1341);
or U1877 (N_1877,N_1064,N_1268);
nor U1878 (N_1878,N_1445,N_1024);
or U1879 (N_1879,N_1207,N_1285);
xnor U1880 (N_1880,N_1323,N_1082);
or U1881 (N_1881,N_1076,N_1094);
nand U1882 (N_1882,N_1333,N_1198);
nor U1883 (N_1883,N_1261,N_1458);
nor U1884 (N_1884,N_1467,N_1045);
or U1885 (N_1885,N_1074,N_1425);
or U1886 (N_1886,N_1278,N_1271);
nand U1887 (N_1887,N_1053,N_1196);
nand U1888 (N_1888,N_1045,N_1229);
and U1889 (N_1889,N_1225,N_1166);
nand U1890 (N_1890,N_1034,N_1298);
and U1891 (N_1891,N_1471,N_1336);
and U1892 (N_1892,N_1449,N_1099);
nor U1893 (N_1893,N_1281,N_1225);
nand U1894 (N_1894,N_1050,N_1202);
nor U1895 (N_1895,N_1110,N_1146);
or U1896 (N_1896,N_1071,N_1195);
nand U1897 (N_1897,N_1219,N_1442);
nor U1898 (N_1898,N_1267,N_1168);
or U1899 (N_1899,N_1365,N_1419);
nor U1900 (N_1900,N_1102,N_1068);
and U1901 (N_1901,N_1307,N_1450);
nand U1902 (N_1902,N_1104,N_1003);
nor U1903 (N_1903,N_1109,N_1093);
xor U1904 (N_1904,N_1286,N_1351);
nand U1905 (N_1905,N_1305,N_1455);
or U1906 (N_1906,N_1008,N_1206);
or U1907 (N_1907,N_1036,N_1262);
and U1908 (N_1908,N_1384,N_1353);
or U1909 (N_1909,N_1332,N_1127);
and U1910 (N_1910,N_1133,N_1332);
nor U1911 (N_1911,N_1033,N_1270);
and U1912 (N_1912,N_1011,N_1388);
nand U1913 (N_1913,N_1162,N_1369);
xor U1914 (N_1914,N_1406,N_1391);
and U1915 (N_1915,N_1431,N_1384);
xnor U1916 (N_1916,N_1469,N_1459);
and U1917 (N_1917,N_1241,N_1381);
nor U1918 (N_1918,N_1225,N_1431);
or U1919 (N_1919,N_1384,N_1295);
nor U1920 (N_1920,N_1138,N_1431);
nor U1921 (N_1921,N_1179,N_1448);
and U1922 (N_1922,N_1358,N_1490);
nor U1923 (N_1923,N_1332,N_1216);
and U1924 (N_1924,N_1103,N_1081);
and U1925 (N_1925,N_1479,N_1207);
nor U1926 (N_1926,N_1133,N_1118);
nor U1927 (N_1927,N_1041,N_1425);
xor U1928 (N_1928,N_1157,N_1294);
nand U1929 (N_1929,N_1125,N_1091);
nand U1930 (N_1930,N_1496,N_1069);
nand U1931 (N_1931,N_1473,N_1190);
nand U1932 (N_1932,N_1303,N_1464);
nand U1933 (N_1933,N_1396,N_1086);
nor U1934 (N_1934,N_1089,N_1182);
nand U1935 (N_1935,N_1489,N_1164);
and U1936 (N_1936,N_1493,N_1185);
and U1937 (N_1937,N_1287,N_1253);
nor U1938 (N_1938,N_1070,N_1258);
or U1939 (N_1939,N_1142,N_1027);
nor U1940 (N_1940,N_1079,N_1238);
or U1941 (N_1941,N_1056,N_1117);
and U1942 (N_1942,N_1339,N_1480);
nand U1943 (N_1943,N_1475,N_1219);
xnor U1944 (N_1944,N_1056,N_1012);
nand U1945 (N_1945,N_1275,N_1247);
or U1946 (N_1946,N_1432,N_1412);
nand U1947 (N_1947,N_1163,N_1351);
nor U1948 (N_1948,N_1008,N_1048);
or U1949 (N_1949,N_1044,N_1372);
nand U1950 (N_1950,N_1298,N_1450);
or U1951 (N_1951,N_1454,N_1494);
nor U1952 (N_1952,N_1008,N_1238);
nor U1953 (N_1953,N_1261,N_1088);
or U1954 (N_1954,N_1043,N_1021);
nand U1955 (N_1955,N_1084,N_1078);
and U1956 (N_1956,N_1489,N_1306);
and U1957 (N_1957,N_1115,N_1378);
nand U1958 (N_1958,N_1049,N_1332);
or U1959 (N_1959,N_1361,N_1223);
or U1960 (N_1960,N_1460,N_1385);
and U1961 (N_1961,N_1099,N_1173);
or U1962 (N_1962,N_1185,N_1298);
nor U1963 (N_1963,N_1195,N_1302);
or U1964 (N_1964,N_1493,N_1305);
or U1965 (N_1965,N_1445,N_1314);
nand U1966 (N_1966,N_1264,N_1359);
or U1967 (N_1967,N_1182,N_1149);
or U1968 (N_1968,N_1496,N_1351);
or U1969 (N_1969,N_1259,N_1249);
nor U1970 (N_1970,N_1351,N_1078);
nand U1971 (N_1971,N_1300,N_1020);
xnor U1972 (N_1972,N_1191,N_1379);
and U1973 (N_1973,N_1114,N_1148);
nand U1974 (N_1974,N_1434,N_1416);
nor U1975 (N_1975,N_1225,N_1487);
nand U1976 (N_1976,N_1362,N_1495);
nand U1977 (N_1977,N_1116,N_1115);
and U1978 (N_1978,N_1489,N_1349);
nor U1979 (N_1979,N_1180,N_1243);
nor U1980 (N_1980,N_1167,N_1206);
nor U1981 (N_1981,N_1153,N_1301);
and U1982 (N_1982,N_1075,N_1202);
nand U1983 (N_1983,N_1304,N_1320);
nor U1984 (N_1984,N_1149,N_1044);
and U1985 (N_1985,N_1028,N_1458);
or U1986 (N_1986,N_1413,N_1017);
nor U1987 (N_1987,N_1011,N_1462);
nor U1988 (N_1988,N_1335,N_1255);
nand U1989 (N_1989,N_1111,N_1104);
nand U1990 (N_1990,N_1007,N_1073);
nor U1991 (N_1991,N_1301,N_1162);
or U1992 (N_1992,N_1272,N_1018);
nor U1993 (N_1993,N_1314,N_1019);
and U1994 (N_1994,N_1388,N_1160);
and U1995 (N_1995,N_1246,N_1239);
xor U1996 (N_1996,N_1074,N_1410);
and U1997 (N_1997,N_1149,N_1320);
or U1998 (N_1998,N_1483,N_1195);
or U1999 (N_1999,N_1326,N_1084);
nor U2000 (N_2000,N_1763,N_1900);
or U2001 (N_2001,N_1707,N_1932);
and U2002 (N_2002,N_1630,N_1990);
and U2003 (N_2003,N_1804,N_1818);
or U2004 (N_2004,N_1935,N_1758);
xor U2005 (N_2005,N_1983,N_1757);
and U2006 (N_2006,N_1565,N_1819);
or U2007 (N_2007,N_1860,N_1993);
xor U2008 (N_2008,N_1610,N_1748);
nand U2009 (N_2009,N_1674,N_1696);
or U2010 (N_2010,N_1655,N_1967);
nand U2011 (N_2011,N_1977,N_1936);
nor U2012 (N_2012,N_1994,N_1880);
and U2013 (N_2013,N_1780,N_1568);
and U2014 (N_2014,N_1843,N_1584);
and U2015 (N_2015,N_1523,N_1593);
nand U2016 (N_2016,N_1502,N_1745);
or U2017 (N_2017,N_1531,N_1778);
xnor U2018 (N_2018,N_1850,N_1576);
nor U2019 (N_2019,N_1641,N_1891);
nor U2020 (N_2020,N_1762,N_1901);
and U2021 (N_2021,N_1734,N_1546);
nand U2022 (N_2022,N_1680,N_1938);
nand U2023 (N_2023,N_1837,N_1585);
nor U2024 (N_2024,N_1689,N_1879);
and U2025 (N_2025,N_1806,N_1526);
and U2026 (N_2026,N_1826,N_1720);
nand U2027 (N_2027,N_1809,N_1892);
nor U2028 (N_2028,N_1515,N_1697);
and U2029 (N_2029,N_1844,N_1686);
nand U2030 (N_2030,N_1840,N_1521);
nand U2031 (N_2031,N_1652,N_1767);
or U2032 (N_2032,N_1574,N_1627);
or U2033 (N_2033,N_1611,N_1975);
or U2034 (N_2034,N_1862,N_1501);
or U2035 (N_2035,N_1668,N_1999);
or U2036 (N_2036,N_1561,N_1594);
nor U2037 (N_2037,N_1859,N_1898);
and U2038 (N_2038,N_1598,N_1532);
xor U2039 (N_2039,N_1823,N_1604);
and U2040 (N_2040,N_1789,N_1884);
xor U2041 (N_2041,N_1587,N_1529);
and U2042 (N_2042,N_1519,N_1772);
nor U2043 (N_2043,N_1817,N_1712);
or U2044 (N_2044,N_1897,N_1960);
nand U2045 (N_2045,N_1916,N_1640);
xor U2046 (N_2046,N_1729,N_1846);
or U2047 (N_2047,N_1797,N_1746);
or U2048 (N_2048,N_1908,N_1943);
nand U2049 (N_2049,N_1638,N_1777);
nor U2050 (N_2050,N_1774,N_1595);
nor U2051 (N_2051,N_1941,N_1863);
or U2052 (N_2052,N_1728,N_1933);
nor U2053 (N_2053,N_1613,N_1549);
or U2054 (N_2054,N_1962,N_1682);
or U2055 (N_2055,N_1937,N_1873);
nand U2056 (N_2056,N_1779,N_1539);
or U2057 (N_2057,N_1925,N_1876);
and U2058 (N_2058,N_1713,N_1725);
xnor U2059 (N_2059,N_1737,N_1679);
or U2060 (N_2060,N_1827,N_1555);
nor U2061 (N_2061,N_1554,N_1537);
nor U2062 (N_2062,N_1899,N_1822);
nand U2063 (N_2063,N_1566,N_1601);
and U2064 (N_2064,N_1885,N_1909);
and U2065 (N_2065,N_1735,N_1731);
and U2066 (N_2066,N_1978,N_1761);
nand U2067 (N_2067,N_1877,N_1509);
nand U2068 (N_2068,N_1872,N_1619);
nor U2069 (N_2069,N_1802,N_1784);
nand U2070 (N_2070,N_1514,N_1996);
xor U2071 (N_2071,N_1952,N_1698);
nand U2072 (N_2072,N_1550,N_1547);
and U2073 (N_2073,N_1847,N_1985);
nor U2074 (N_2074,N_1869,N_1914);
nand U2075 (N_2075,N_1959,N_1646);
nand U2076 (N_2076,N_1542,N_1934);
nand U2077 (N_2077,N_1830,N_1670);
and U2078 (N_2078,N_1856,N_1692);
or U2079 (N_2079,N_1991,N_1560);
nand U2080 (N_2080,N_1849,N_1683);
and U2081 (N_2081,N_1868,N_1551);
xnor U2082 (N_2082,N_1717,N_1792);
and U2083 (N_2083,N_1583,N_1518);
and U2084 (N_2084,N_1520,N_1663);
and U2085 (N_2085,N_1552,N_1870);
nand U2086 (N_2086,N_1808,N_1988);
or U2087 (N_2087,N_1597,N_1970);
or U2088 (N_2088,N_1716,N_1824);
and U2089 (N_2089,N_1634,N_1562);
or U2090 (N_2090,N_1851,N_1785);
nor U2091 (N_2091,N_1966,N_1752);
and U2092 (N_2092,N_1558,N_1599);
or U2093 (N_2093,N_1760,N_1660);
nand U2094 (N_2094,N_1825,N_1838);
and U2095 (N_2095,N_1968,N_1906);
nor U2096 (N_2096,N_1563,N_1794);
nor U2097 (N_2097,N_1878,N_1861);
and U2098 (N_2098,N_1733,N_1724);
nand U2099 (N_2099,N_1675,N_1889);
xor U2100 (N_2100,N_1928,N_1704);
nor U2101 (N_2101,N_1754,N_1582);
and U2102 (N_2102,N_1807,N_1931);
or U2103 (N_2103,N_1755,N_1955);
nand U2104 (N_2104,N_1556,N_1687);
nor U2105 (N_2105,N_1572,N_1649);
and U2106 (N_2106,N_1617,N_1522);
or U2107 (N_2107,N_1917,N_1592);
nor U2108 (N_2108,N_1886,N_1756);
or U2109 (N_2109,N_1940,N_1678);
or U2110 (N_2110,N_1658,N_1616);
nand U2111 (N_2111,N_1622,N_1694);
nand U2112 (N_2112,N_1912,N_1915);
nor U2113 (N_2113,N_1691,N_1987);
nor U2114 (N_2114,N_1533,N_1570);
or U2115 (N_2115,N_1929,N_1633);
xor U2116 (N_2116,N_1647,N_1816);
and U2117 (N_2117,N_1528,N_1544);
nand U2118 (N_2118,N_1581,N_1930);
nand U2119 (N_2119,N_1773,N_1685);
nor U2120 (N_2120,N_1578,N_1510);
and U2121 (N_2121,N_1895,N_1858);
nand U2122 (N_2122,N_1922,N_1703);
nand U2123 (N_2123,N_1971,N_1636);
nand U2124 (N_2124,N_1618,N_1961);
nand U2125 (N_2125,N_1946,N_1771);
or U2126 (N_2126,N_1710,N_1524);
nand U2127 (N_2127,N_1783,N_1839);
and U2128 (N_2128,N_1577,N_1702);
nand U2129 (N_2129,N_1676,N_1919);
and U2130 (N_2130,N_1596,N_1871);
or U2131 (N_2131,N_1648,N_1708);
nor U2132 (N_2132,N_1516,N_1650);
nor U2133 (N_2133,N_1654,N_1671);
xor U2134 (N_2134,N_1743,N_1688);
nand U2135 (N_2135,N_1637,N_1815);
and U2136 (N_2136,N_1951,N_1764);
nor U2137 (N_2137,N_1672,N_1681);
nand U2138 (N_2138,N_1645,N_1997);
and U2139 (N_2139,N_1927,N_1662);
and U2140 (N_2140,N_1606,N_1864);
nor U2141 (N_2141,N_1958,N_1677);
nor U2142 (N_2142,N_1793,N_1569);
or U2143 (N_2143,N_1984,N_1913);
nand U2144 (N_2144,N_1625,N_1736);
nand U2145 (N_2145,N_1727,N_1765);
nor U2146 (N_2146,N_1890,N_1669);
nor U2147 (N_2147,N_1742,N_1998);
nand U2148 (N_2148,N_1911,N_1656);
and U2149 (N_2149,N_1706,N_1799);
nand U2150 (N_2150,N_1882,N_1881);
and U2151 (N_2151,N_1836,N_1541);
nor U2152 (N_2152,N_1699,N_1974);
xor U2153 (N_2153,N_1982,N_1992);
xor U2154 (N_2154,N_1530,N_1540);
nor U2155 (N_2155,N_1673,N_1575);
or U2156 (N_2156,N_1798,N_1953);
nand U2157 (N_2157,N_1776,N_1795);
or U2158 (N_2158,N_1621,N_1722);
nor U2159 (N_2159,N_1666,N_1718);
nor U2160 (N_2160,N_1829,N_1883);
or U2161 (N_2161,N_1588,N_1723);
nand U2162 (N_2162,N_1709,N_1508);
nor U2163 (N_2163,N_1715,N_1989);
and U2164 (N_2164,N_1517,N_1602);
and U2165 (N_2165,N_1741,N_1923);
and U2166 (N_2166,N_1853,N_1609);
or U2167 (N_2167,N_1865,N_1976);
xor U2168 (N_2168,N_1845,N_1738);
xor U2169 (N_2169,N_1639,N_1848);
and U2170 (N_2170,N_1769,N_1814);
nand U2171 (N_2171,N_1553,N_1732);
nor U2172 (N_2172,N_1980,N_1600);
and U2173 (N_2173,N_1750,N_1714);
nand U2174 (N_2174,N_1907,N_1632);
nand U2175 (N_2175,N_1896,N_1721);
and U2176 (N_2176,N_1507,N_1605);
or U2177 (N_2177,N_1614,N_1973);
nor U2178 (N_2178,N_1512,N_1903);
or U2179 (N_2179,N_1854,N_1749);
and U2180 (N_2180,N_1875,N_1950);
nand U2181 (N_2181,N_1500,N_1665);
and U2182 (N_2182,N_1753,N_1653);
nand U2183 (N_2183,N_1589,N_1527);
or U2184 (N_2184,N_1801,N_1800);
nor U2185 (N_2185,N_1945,N_1924);
nand U2186 (N_2186,N_1820,N_1964);
nand U2187 (N_2187,N_1894,N_1511);
and U2188 (N_2188,N_1813,N_1770);
nand U2189 (N_2189,N_1834,N_1835);
xor U2190 (N_2190,N_1571,N_1701);
and U2191 (N_2191,N_1579,N_1874);
and U2192 (N_2192,N_1586,N_1751);
or U2193 (N_2193,N_1690,N_1759);
nor U2194 (N_2194,N_1643,N_1888);
or U2195 (N_2195,N_1969,N_1624);
nand U2196 (N_2196,N_1791,N_1657);
nand U2197 (N_2197,N_1812,N_1534);
xnor U2198 (N_2198,N_1504,N_1719);
nor U2199 (N_2199,N_1766,N_1543);
nor U2200 (N_2200,N_1661,N_1920);
nand U2201 (N_2201,N_1893,N_1603);
or U2202 (N_2202,N_1867,N_1536);
or U2203 (N_2203,N_1944,N_1538);
nand U2204 (N_2204,N_1525,N_1902);
and U2205 (N_2205,N_1573,N_1942);
nor U2206 (N_2206,N_1535,N_1623);
and U2207 (N_2207,N_1744,N_1629);
nor U2208 (N_2208,N_1833,N_1910);
nand U2209 (N_2209,N_1904,N_1866);
nor U2210 (N_2210,N_1805,N_1796);
nand U2211 (N_2211,N_1986,N_1981);
and U2212 (N_2212,N_1659,N_1995);
nand U2213 (N_2213,N_1612,N_1857);
nor U2214 (N_2214,N_1972,N_1887);
nand U2215 (N_2215,N_1954,N_1747);
xor U2216 (N_2216,N_1548,N_1726);
nor U2217 (N_2217,N_1580,N_1787);
xnor U2218 (N_2218,N_1842,N_1810);
nor U2219 (N_2219,N_1768,N_1608);
or U2220 (N_2220,N_1664,N_1979);
nor U2221 (N_2221,N_1607,N_1841);
nor U2222 (N_2222,N_1947,N_1926);
and U2223 (N_2223,N_1545,N_1786);
nand U2224 (N_2224,N_1918,N_1831);
and U2225 (N_2225,N_1739,N_1921);
nand U2226 (N_2226,N_1642,N_1700);
and U2227 (N_2227,N_1939,N_1855);
nor U2228 (N_2228,N_1503,N_1505);
or U2229 (N_2229,N_1905,N_1711);
or U2230 (N_2230,N_1788,N_1828);
nor U2231 (N_2231,N_1591,N_1811);
xnor U2232 (N_2232,N_1730,N_1693);
xor U2233 (N_2233,N_1626,N_1631);
nand U2234 (N_2234,N_1635,N_1782);
nand U2235 (N_2235,N_1775,N_1852);
or U2236 (N_2236,N_1644,N_1790);
or U2237 (N_2237,N_1513,N_1957);
nor U2238 (N_2238,N_1590,N_1620);
nor U2239 (N_2239,N_1963,N_1651);
xnor U2240 (N_2240,N_1567,N_1667);
nor U2241 (N_2241,N_1949,N_1506);
or U2242 (N_2242,N_1821,N_1705);
nor U2243 (N_2243,N_1564,N_1956);
or U2244 (N_2244,N_1559,N_1628);
or U2245 (N_2245,N_1803,N_1781);
xnor U2246 (N_2246,N_1965,N_1948);
and U2247 (N_2247,N_1695,N_1740);
xor U2248 (N_2248,N_1832,N_1615);
or U2249 (N_2249,N_1557,N_1684);
nand U2250 (N_2250,N_1833,N_1594);
and U2251 (N_2251,N_1754,N_1748);
nand U2252 (N_2252,N_1853,N_1665);
or U2253 (N_2253,N_1920,N_1590);
nor U2254 (N_2254,N_1632,N_1816);
or U2255 (N_2255,N_1956,N_1835);
and U2256 (N_2256,N_1572,N_1685);
or U2257 (N_2257,N_1913,N_1602);
nor U2258 (N_2258,N_1694,N_1563);
nor U2259 (N_2259,N_1575,N_1595);
nand U2260 (N_2260,N_1540,N_1997);
and U2261 (N_2261,N_1988,N_1897);
or U2262 (N_2262,N_1885,N_1671);
nor U2263 (N_2263,N_1692,N_1847);
or U2264 (N_2264,N_1892,N_1945);
nand U2265 (N_2265,N_1997,N_1587);
nand U2266 (N_2266,N_1858,N_1536);
nand U2267 (N_2267,N_1758,N_1607);
xnor U2268 (N_2268,N_1890,N_1816);
or U2269 (N_2269,N_1543,N_1679);
nand U2270 (N_2270,N_1960,N_1601);
nor U2271 (N_2271,N_1781,N_1860);
nand U2272 (N_2272,N_1591,N_1602);
or U2273 (N_2273,N_1574,N_1599);
xor U2274 (N_2274,N_1979,N_1591);
nand U2275 (N_2275,N_1766,N_1678);
nor U2276 (N_2276,N_1732,N_1974);
or U2277 (N_2277,N_1983,N_1575);
and U2278 (N_2278,N_1799,N_1857);
nor U2279 (N_2279,N_1525,N_1667);
nor U2280 (N_2280,N_1783,N_1706);
nor U2281 (N_2281,N_1721,N_1801);
or U2282 (N_2282,N_1695,N_1569);
and U2283 (N_2283,N_1769,N_1574);
nor U2284 (N_2284,N_1951,N_1788);
or U2285 (N_2285,N_1724,N_1647);
or U2286 (N_2286,N_1979,N_1594);
or U2287 (N_2287,N_1968,N_1865);
or U2288 (N_2288,N_1709,N_1532);
nand U2289 (N_2289,N_1769,N_1880);
xnor U2290 (N_2290,N_1907,N_1890);
nand U2291 (N_2291,N_1628,N_1668);
nor U2292 (N_2292,N_1914,N_1874);
or U2293 (N_2293,N_1988,N_1916);
or U2294 (N_2294,N_1547,N_1886);
and U2295 (N_2295,N_1699,N_1940);
or U2296 (N_2296,N_1973,N_1805);
nor U2297 (N_2297,N_1668,N_1620);
nand U2298 (N_2298,N_1930,N_1924);
nor U2299 (N_2299,N_1786,N_1713);
nand U2300 (N_2300,N_1734,N_1898);
and U2301 (N_2301,N_1741,N_1564);
nor U2302 (N_2302,N_1969,N_1825);
nor U2303 (N_2303,N_1998,N_1959);
nor U2304 (N_2304,N_1775,N_1987);
or U2305 (N_2305,N_1846,N_1644);
nand U2306 (N_2306,N_1669,N_1895);
nand U2307 (N_2307,N_1860,N_1784);
or U2308 (N_2308,N_1886,N_1968);
xor U2309 (N_2309,N_1578,N_1520);
nor U2310 (N_2310,N_1942,N_1506);
nand U2311 (N_2311,N_1965,N_1667);
and U2312 (N_2312,N_1535,N_1516);
xor U2313 (N_2313,N_1947,N_1622);
xnor U2314 (N_2314,N_1706,N_1595);
nand U2315 (N_2315,N_1705,N_1743);
and U2316 (N_2316,N_1835,N_1912);
xnor U2317 (N_2317,N_1938,N_1925);
or U2318 (N_2318,N_1550,N_1573);
nor U2319 (N_2319,N_1994,N_1774);
or U2320 (N_2320,N_1725,N_1507);
and U2321 (N_2321,N_1986,N_1615);
nor U2322 (N_2322,N_1762,N_1940);
or U2323 (N_2323,N_1943,N_1719);
nor U2324 (N_2324,N_1642,N_1726);
nand U2325 (N_2325,N_1530,N_1746);
nor U2326 (N_2326,N_1684,N_1965);
or U2327 (N_2327,N_1646,N_1853);
or U2328 (N_2328,N_1988,N_1830);
and U2329 (N_2329,N_1595,N_1839);
and U2330 (N_2330,N_1592,N_1955);
or U2331 (N_2331,N_1657,N_1937);
nor U2332 (N_2332,N_1899,N_1845);
nor U2333 (N_2333,N_1774,N_1917);
nor U2334 (N_2334,N_1900,N_1891);
or U2335 (N_2335,N_1678,N_1597);
or U2336 (N_2336,N_1605,N_1909);
or U2337 (N_2337,N_1939,N_1761);
and U2338 (N_2338,N_1874,N_1973);
or U2339 (N_2339,N_1505,N_1846);
xor U2340 (N_2340,N_1761,N_1676);
nor U2341 (N_2341,N_1547,N_1564);
or U2342 (N_2342,N_1659,N_1710);
or U2343 (N_2343,N_1934,N_1681);
or U2344 (N_2344,N_1599,N_1729);
nand U2345 (N_2345,N_1671,N_1893);
or U2346 (N_2346,N_1776,N_1972);
and U2347 (N_2347,N_1584,N_1748);
xor U2348 (N_2348,N_1897,N_1905);
and U2349 (N_2349,N_1992,N_1886);
xor U2350 (N_2350,N_1768,N_1641);
or U2351 (N_2351,N_1803,N_1948);
nand U2352 (N_2352,N_1591,N_1905);
and U2353 (N_2353,N_1551,N_1580);
nand U2354 (N_2354,N_1677,N_1581);
and U2355 (N_2355,N_1703,N_1926);
nor U2356 (N_2356,N_1708,N_1596);
nand U2357 (N_2357,N_1600,N_1537);
nand U2358 (N_2358,N_1579,N_1573);
and U2359 (N_2359,N_1738,N_1826);
and U2360 (N_2360,N_1652,N_1900);
nand U2361 (N_2361,N_1960,N_1659);
or U2362 (N_2362,N_1598,N_1629);
or U2363 (N_2363,N_1711,N_1741);
and U2364 (N_2364,N_1857,N_1600);
xnor U2365 (N_2365,N_1519,N_1645);
or U2366 (N_2366,N_1804,N_1581);
nand U2367 (N_2367,N_1924,N_1568);
or U2368 (N_2368,N_1664,N_1999);
nor U2369 (N_2369,N_1879,N_1960);
xnor U2370 (N_2370,N_1932,N_1626);
or U2371 (N_2371,N_1721,N_1524);
or U2372 (N_2372,N_1525,N_1612);
nand U2373 (N_2373,N_1962,N_1949);
xnor U2374 (N_2374,N_1861,N_1530);
and U2375 (N_2375,N_1802,N_1696);
or U2376 (N_2376,N_1734,N_1739);
nor U2377 (N_2377,N_1972,N_1628);
or U2378 (N_2378,N_1697,N_1746);
and U2379 (N_2379,N_1672,N_1790);
nor U2380 (N_2380,N_1544,N_1510);
nand U2381 (N_2381,N_1881,N_1974);
nand U2382 (N_2382,N_1606,N_1884);
nand U2383 (N_2383,N_1967,N_1725);
and U2384 (N_2384,N_1974,N_1515);
or U2385 (N_2385,N_1904,N_1952);
and U2386 (N_2386,N_1901,N_1892);
and U2387 (N_2387,N_1726,N_1969);
nor U2388 (N_2388,N_1680,N_1943);
and U2389 (N_2389,N_1732,N_1900);
xnor U2390 (N_2390,N_1859,N_1648);
or U2391 (N_2391,N_1601,N_1727);
xor U2392 (N_2392,N_1978,N_1941);
or U2393 (N_2393,N_1891,N_1763);
or U2394 (N_2394,N_1909,N_1945);
nand U2395 (N_2395,N_1682,N_1519);
nand U2396 (N_2396,N_1678,N_1677);
nor U2397 (N_2397,N_1927,N_1762);
nor U2398 (N_2398,N_1731,N_1524);
xnor U2399 (N_2399,N_1742,N_1983);
and U2400 (N_2400,N_1925,N_1546);
or U2401 (N_2401,N_1813,N_1555);
and U2402 (N_2402,N_1963,N_1530);
nand U2403 (N_2403,N_1953,N_1974);
nor U2404 (N_2404,N_1562,N_1809);
xor U2405 (N_2405,N_1618,N_1541);
nor U2406 (N_2406,N_1647,N_1859);
xnor U2407 (N_2407,N_1704,N_1656);
nand U2408 (N_2408,N_1538,N_1856);
and U2409 (N_2409,N_1610,N_1811);
and U2410 (N_2410,N_1683,N_1816);
nor U2411 (N_2411,N_1615,N_1710);
nor U2412 (N_2412,N_1690,N_1869);
and U2413 (N_2413,N_1557,N_1564);
and U2414 (N_2414,N_1942,N_1599);
nand U2415 (N_2415,N_1873,N_1691);
nor U2416 (N_2416,N_1812,N_1961);
or U2417 (N_2417,N_1799,N_1568);
nand U2418 (N_2418,N_1800,N_1694);
nand U2419 (N_2419,N_1773,N_1853);
nand U2420 (N_2420,N_1999,N_1975);
nor U2421 (N_2421,N_1998,N_1549);
nor U2422 (N_2422,N_1842,N_1676);
or U2423 (N_2423,N_1746,N_1931);
or U2424 (N_2424,N_1564,N_1959);
xnor U2425 (N_2425,N_1839,N_1735);
or U2426 (N_2426,N_1997,N_1960);
or U2427 (N_2427,N_1970,N_1929);
nand U2428 (N_2428,N_1717,N_1640);
and U2429 (N_2429,N_1639,N_1770);
and U2430 (N_2430,N_1627,N_1975);
or U2431 (N_2431,N_1954,N_1586);
nand U2432 (N_2432,N_1990,N_1512);
nor U2433 (N_2433,N_1692,N_1537);
nor U2434 (N_2434,N_1908,N_1851);
nor U2435 (N_2435,N_1527,N_1927);
nor U2436 (N_2436,N_1700,N_1997);
nor U2437 (N_2437,N_1541,N_1907);
or U2438 (N_2438,N_1865,N_1790);
nand U2439 (N_2439,N_1643,N_1779);
or U2440 (N_2440,N_1791,N_1546);
nand U2441 (N_2441,N_1862,N_1536);
or U2442 (N_2442,N_1962,N_1622);
or U2443 (N_2443,N_1775,N_1930);
or U2444 (N_2444,N_1677,N_1616);
nand U2445 (N_2445,N_1961,N_1566);
or U2446 (N_2446,N_1620,N_1585);
or U2447 (N_2447,N_1622,N_1887);
nand U2448 (N_2448,N_1942,N_1687);
and U2449 (N_2449,N_1557,N_1783);
nor U2450 (N_2450,N_1785,N_1730);
nand U2451 (N_2451,N_1916,N_1516);
nor U2452 (N_2452,N_1980,N_1787);
xor U2453 (N_2453,N_1728,N_1928);
or U2454 (N_2454,N_1807,N_1886);
xnor U2455 (N_2455,N_1921,N_1909);
or U2456 (N_2456,N_1901,N_1671);
or U2457 (N_2457,N_1703,N_1745);
nand U2458 (N_2458,N_1951,N_1629);
or U2459 (N_2459,N_1698,N_1579);
nor U2460 (N_2460,N_1589,N_1897);
nor U2461 (N_2461,N_1729,N_1738);
or U2462 (N_2462,N_1780,N_1565);
or U2463 (N_2463,N_1945,N_1548);
nand U2464 (N_2464,N_1749,N_1799);
or U2465 (N_2465,N_1941,N_1548);
nor U2466 (N_2466,N_1682,N_1869);
and U2467 (N_2467,N_1627,N_1626);
and U2468 (N_2468,N_1607,N_1556);
nor U2469 (N_2469,N_1797,N_1510);
and U2470 (N_2470,N_1793,N_1602);
nand U2471 (N_2471,N_1854,N_1774);
nor U2472 (N_2472,N_1517,N_1896);
or U2473 (N_2473,N_1521,N_1901);
or U2474 (N_2474,N_1605,N_1876);
nand U2475 (N_2475,N_1971,N_1673);
xnor U2476 (N_2476,N_1990,N_1766);
nor U2477 (N_2477,N_1834,N_1913);
nor U2478 (N_2478,N_1668,N_1923);
xor U2479 (N_2479,N_1756,N_1929);
and U2480 (N_2480,N_1817,N_1704);
nand U2481 (N_2481,N_1719,N_1770);
nand U2482 (N_2482,N_1979,N_1682);
or U2483 (N_2483,N_1605,N_1738);
nand U2484 (N_2484,N_1502,N_1680);
nand U2485 (N_2485,N_1596,N_1515);
nand U2486 (N_2486,N_1968,N_1885);
nor U2487 (N_2487,N_1649,N_1872);
and U2488 (N_2488,N_1799,N_1698);
or U2489 (N_2489,N_1649,N_1875);
or U2490 (N_2490,N_1643,N_1588);
nor U2491 (N_2491,N_1956,N_1586);
or U2492 (N_2492,N_1900,N_1667);
nor U2493 (N_2493,N_1910,N_1538);
or U2494 (N_2494,N_1836,N_1720);
nand U2495 (N_2495,N_1858,N_1780);
or U2496 (N_2496,N_1761,N_1678);
nor U2497 (N_2497,N_1830,N_1995);
and U2498 (N_2498,N_1541,N_1982);
nand U2499 (N_2499,N_1757,N_1803);
or U2500 (N_2500,N_2291,N_2169);
nor U2501 (N_2501,N_2316,N_2397);
and U2502 (N_2502,N_2073,N_2077);
nor U2503 (N_2503,N_2005,N_2284);
or U2504 (N_2504,N_2434,N_2238);
nand U2505 (N_2505,N_2301,N_2456);
and U2506 (N_2506,N_2300,N_2455);
or U2507 (N_2507,N_2369,N_2231);
nor U2508 (N_2508,N_2287,N_2004);
or U2509 (N_2509,N_2362,N_2071);
nand U2510 (N_2510,N_2090,N_2143);
nand U2511 (N_2511,N_2003,N_2123);
and U2512 (N_2512,N_2440,N_2364);
and U2513 (N_2513,N_2172,N_2002);
nor U2514 (N_2514,N_2407,N_2086);
and U2515 (N_2515,N_2280,N_2279);
and U2516 (N_2516,N_2351,N_2135);
xor U2517 (N_2517,N_2368,N_2055);
and U2518 (N_2518,N_2386,N_2251);
and U2519 (N_2519,N_2059,N_2042);
nand U2520 (N_2520,N_2022,N_2179);
xnor U2521 (N_2521,N_2008,N_2140);
or U2522 (N_2522,N_2085,N_2379);
nor U2523 (N_2523,N_2234,N_2147);
or U2524 (N_2524,N_2239,N_2396);
nor U2525 (N_2525,N_2117,N_2484);
or U2526 (N_2526,N_2425,N_2120);
and U2527 (N_2527,N_2095,N_2034);
nand U2528 (N_2528,N_2339,N_2448);
nor U2529 (N_2529,N_2205,N_2395);
nor U2530 (N_2530,N_2132,N_2373);
and U2531 (N_2531,N_2359,N_2378);
or U2532 (N_2532,N_2346,N_2099);
or U2533 (N_2533,N_2427,N_2430);
and U2534 (N_2534,N_2019,N_2009);
or U2535 (N_2535,N_2489,N_2052);
xor U2536 (N_2536,N_2341,N_2311);
nor U2537 (N_2537,N_2358,N_2289);
nand U2538 (N_2538,N_2146,N_2124);
nor U2539 (N_2539,N_2370,N_2098);
nor U2540 (N_2540,N_2389,N_2190);
nor U2541 (N_2541,N_2277,N_2497);
nor U2542 (N_2542,N_2492,N_2111);
nor U2543 (N_2543,N_2292,N_2193);
nand U2544 (N_2544,N_2417,N_2018);
xor U2545 (N_2545,N_2138,N_2480);
xnor U2546 (N_2546,N_2007,N_2282);
or U2547 (N_2547,N_2000,N_2337);
nor U2548 (N_2548,N_2254,N_2475);
nand U2549 (N_2549,N_2050,N_2366);
nand U2550 (N_2550,N_2357,N_2258);
xnor U2551 (N_2551,N_2079,N_2353);
nor U2552 (N_2552,N_2318,N_2377);
xor U2553 (N_2553,N_2394,N_2092);
nor U2554 (N_2554,N_2107,N_2257);
and U2555 (N_2555,N_2130,N_2259);
and U2556 (N_2556,N_2221,N_2200);
nor U2557 (N_2557,N_2473,N_2442);
xor U2558 (N_2558,N_2435,N_2367);
nand U2559 (N_2559,N_2348,N_2177);
and U2560 (N_2560,N_2250,N_2420);
nand U2561 (N_2561,N_2013,N_2211);
nand U2562 (N_2562,N_2412,N_2436);
nor U2563 (N_2563,N_2468,N_2392);
and U2564 (N_2564,N_2227,N_2184);
or U2565 (N_2565,N_2422,N_2269);
or U2566 (N_2566,N_2155,N_2060);
and U2567 (N_2567,N_2160,N_2192);
nand U2568 (N_2568,N_2262,N_2383);
and U2569 (N_2569,N_2495,N_2167);
nand U2570 (N_2570,N_2183,N_2186);
and U2571 (N_2571,N_2129,N_2108);
nand U2572 (N_2572,N_2446,N_2087);
or U2573 (N_2573,N_2125,N_2290);
nor U2574 (N_2574,N_2161,N_2461);
or U2575 (N_2575,N_2173,N_2295);
and U2576 (N_2576,N_2240,N_2175);
or U2577 (N_2577,N_2064,N_2083);
nor U2578 (N_2578,N_2381,N_2118);
nor U2579 (N_2579,N_2401,N_2325);
or U2580 (N_2580,N_2498,N_2178);
and U2581 (N_2581,N_2260,N_2452);
nand U2582 (N_2582,N_2197,N_2074);
and U2583 (N_2583,N_2017,N_2350);
and U2584 (N_2584,N_2486,N_2168);
nor U2585 (N_2585,N_2032,N_2023);
or U2586 (N_2586,N_2462,N_2218);
or U2587 (N_2587,N_2274,N_2199);
and U2588 (N_2588,N_2443,N_2049);
nor U2589 (N_2589,N_2418,N_2365);
nand U2590 (N_2590,N_2115,N_2445);
and U2591 (N_2591,N_2037,N_2208);
xor U2592 (N_2592,N_2011,N_2390);
nor U2593 (N_2593,N_2058,N_2447);
xor U2594 (N_2594,N_2431,N_2453);
nand U2595 (N_2595,N_2276,N_2194);
nand U2596 (N_2596,N_2171,N_2457);
nor U2597 (N_2597,N_2051,N_2158);
or U2598 (N_2598,N_2066,N_2236);
and U2599 (N_2599,N_2206,N_2075);
nor U2600 (N_2600,N_2048,N_2329);
and U2601 (N_2601,N_2162,N_2265);
xnor U2602 (N_2602,N_2256,N_2310);
nand U2603 (N_2603,N_2356,N_2454);
xor U2604 (N_2604,N_2212,N_2253);
and U2605 (N_2605,N_2345,N_2398);
and U2606 (N_2606,N_2424,N_2245);
or U2607 (N_2607,N_2261,N_2235);
nor U2608 (N_2608,N_2444,N_2209);
or U2609 (N_2609,N_2148,N_2312);
or U2610 (N_2610,N_2187,N_2413);
nor U2611 (N_2611,N_2467,N_2065);
or U2612 (N_2612,N_2237,N_2415);
nor U2613 (N_2613,N_2450,N_2298);
xnor U2614 (N_2614,N_2408,N_2196);
or U2615 (N_2615,N_2402,N_2294);
or U2616 (N_2616,N_2174,N_2268);
xnor U2617 (N_2617,N_2433,N_2399);
or U2618 (N_2618,N_2244,N_2204);
nor U2619 (N_2619,N_2163,N_2061);
or U2620 (N_2620,N_2286,N_2296);
nor U2621 (N_2621,N_2423,N_2152);
nor U2622 (N_2622,N_2222,N_2264);
and U2623 (N_2623,N_2376,N_2278);
nand U2624 (N_2624,N_2069,N_2101);
nor U2625 (N_2625,N_2217,N_2414);
and U2626 (N_2626,N_2159,N_2141);
xor U2627 (N_2627,N_2273,N_2045);
and U2628 (N_2628,N_2046,N_2460);
nand U2629 (N_2629,N_2067,N_2463);
nor U2630 (N_2630,N_2047,N_2384);
or U2631 (N_2631,N_2488,N_2416);
xor U2632 (N_2632,N_2479,N_2170);
or U2633 (N_2633,N_2012,N_2331);
xnor U2634 (N_2634,N_2410,N_2084);
or U2635 (N_2635,N_2082,N_2441);
nor U2636 (N_2636,N_2121,N_2080);
nor U2637 (N_2637,N_2029,N_2180);
and U2638 (N_2638,N_2097,N_2491);
nand U2639 (N_2639,N_2149,N_2031);
nor U2640 (N_2640,N_2142,N_2426);
and U2641 (N_2641,N_2131,N_2033);
nor U2642 (N_2642,N_2156,N_2288);
or U2643 (N_2643,N_2382,N_2409);
nor U2644 (N_2644,N_2363,N_2122);
and U2645 (N_2645,N_2249,N_2299);
and U2646 (N_2646,N_2466,N_2308);
nor U2647 (N_2647,N_2478,N_2188);
or U2648 (N_2648,N_2181,N_2411);
nor U2649 (N_2649,N_2499,N_2465);
or U2650 (N_2650,N_2347,N_2469);
nand U2651 (N_2651,N_2203,N_2342);
or U2652 (N_2652,N_2232,N_2028);
or U2653 (N_2653,N_2438,N_2474);
or U2654 (N_2654,N_2354,N_2116);
nor U2655 (N_2655,N_2493,N_2242);
xnor U2656 (N_2656,N_2210,N_2136);
nor U2657 (N_2657,N_2025,N_2151);
nand U2658 (N_2658,N_2113,N_2272);
nor U2659 (N_2659,N_2038,N_2229);
and U2660 (N_2660,N_2063,N_2223);
or U2661 (N_2661,N_2057,N_2195);
or U2662 (N_2662,N_2380,N_2314);
nand U2663 (N_2663,N_2419,N_2248);
nand U2664 (N_2664,N_2010,N_2246);
or U2665 (N_2665,N_2053,N_2020);
and U2666 (N_2666,N_2360,N_2014);
and U2667 (N_2667,N_2094,N_2428);
and U2668 (N_2668,N_2088,N_2207);
xor U2669 (N_2669,N_2070,N_2214);
nand U2670 (N_2670,N_2213,N_2027);
nor U2671 (N_2671,N_2315,N_2112);
nand U2672 (N_2672,N_2145,N_2432);
or U2673 (N_2673,N_2470,N_2429);
or U2674 (N_2674,N_2344,N_2165);
xor U2675 (N_2675,N_2330,N_2166);
nand U2676 (N_2676,N_2001,N_2157);
or U2677 (N_2677,N_2198,N_2103);
nand U2678 (N_2678,N_2355,N_2281);
nor U2679 (N_2679,N_2109,N_2243);
nand U2680 (N_2680,N_2391,N_2285);
and U2681 (N_2681,N_2283,N_2039);
nand U2682 (N_2682,N_2106,N_2437);
and U2683 (N_2683,N_2313,N_2458);
and U2684 (N_2684,N_2078,N_2326);
nand U2685 (N_2685,N_2263,N_2275);
or U2686 (N_2686,N_2150,N_2482);
nand U2687 (N_2687,N_2476,N_2388);
or U2688 (N_2688,N_2089,N_2056);
or U2689 (N_2689,N_2338,N_2040);
nor U2690 (N_2690,N_2024,N_2182);
and U2691 (N_2691,N_2006,N_2439);
and U2692 (N_2692,N_2374,N_2026);
or U2693 (N_2693,N_2119,N_2228);
or U2694 (N_2694,N_2164,N_2105);
and U2695 (N_2695,N_2247,N_2270);
and U2696 (N_2696,N_2036,N_2335);
nand U2697 (N_2697,N_2322,N_2321);
xnor U2698 (N_2698,N_2307,N_2340);
and U2699 (N_2699,N_2093,N_2303);
nor U2700 (N_2700,N_2449,N_2076);
or U2701 (N_2701,N_2334,N_2371);
or U2702 (N_2702,N_2323,N_2464);
nand U2703 (N_2703,N_2459,N_2387);
or U2704 (N_2704,N_2021,N_2267);
and U2705 (N_2705,N_2044,N_2134);
or U2706 (N_2706,N_2403,N_2271);
and U2707 (N_2707,N_2483,N_2343);
or U2708 (N_2708,N_2471,N_2041);
or U2709 (N_2709,N_2302,N_2100);
xnor U2710 (N_2710,N_2255,N_2015);
xor U2711 (N_2711,N_2081,N_2324);
or U2712 (N_2712,N_2230,N_2224);
nor U2713 (N_2713,N_2490,N_2241);
nand U2714 (N_2714,N_2225,N_2215);
and U2715 (N_2715,N_2266,N_2317);
nand U2716 (N_2716,N_2297,N_2494);
xnor U2717 (N_2717,N_2406,N_2472);
and U2718 (N_2718,N_2304,N_2349);
and U2719 (N_2719,N_2400,N_2352);
nor U2720 (N_2720,N_2404,N_2309);
nor U2721 (N_2721,N_2385,N_2293);
or U2722 (N_2722,N_2104,N_2185);
nor U2723 (N_2723,N_2333,N_2072);
nand U2724 (N_2724,N_2062,N_2477);
nand U2725 (N_2725,N_2216,N_2252);
nand U2726 (N_2726,N_2421,N_2332);
xnor U2727 (N_2727,N_2191,N_2153);
and U2728 (N_2728,N_2393,N_2016);
nor U2729 (N_2729,N_2372,N_2405);
and U2730 (N_2730,N_2496,N_2220);
and U2731 (N_2731,N_2202,N_2091);
nor U2732 (N_2732,N_2361,N_2201);
nor U2733 (N_2733,N_2306,N_2128);
nand U2734 (N_2734,N_2114,N_2043);
and U2735 (N_2735,N_2176,N_2319);
or U2736 (N_2736,N_2127,N_2068);
nand U2737 (N_2737,N_2487,N_2126);
nor U2738 (N_2738,N_2030,N_2139);
nand U2739 (N_2739,N_2375,N_2144);
nor U2740 (N_2740,N_2054,N_2485);
nand U2741 (N_2741,N_2305,N_2189);
and U2742 (N_2742,N_2328,N_2096);
nand U2743 (N_2743,N_2133,N_2219);
and U2744 (N_2744,N_2137,N_2226);
xor U2745 (N_2745,N_2320,N_2481);
or U2746 (N_2746,N_2336,N_2327);
xnor U2747 (N_2747,N_2035,N_2451);
and U2748 (N_2748,N_2110,N_2154);
nor U2749 (N_2749,N_2102,N_2233);
nand U2750 (N_2750,N_2480,N_2430);
nand U2751 (N_2751,N_2468,N_2136);
nor U2752 (N_2752,N_2253,N_2449);
nor U2753 (N_2753,N_2286,N_2037);
or U2754 (N_2754,N_2071,N_2486);
and U2755 (N_2755,N_2071,N_2370);
xor U2756 (N_2756,N_2089,N_2241);
and U2757 (N_2757,N_2047,N_2120);
xor U2758 (N_2758,N_2465,N_2105);
or U2759 (N_2759,N_2341,N_2094);
nor U2760 (N_2760,N_2268,N_2343);
nand U2761 (N_2761,N_2486,N_2008);
nand U2762 (N_2762,N_2209,N_2134);
or U2763 (N_2763,N_2360,N_2363);
nor U2764 (N_2764,N_2430,N_2417);
nand U2765 (N_2765,N_2206,N_2142);
nor U2766 (N_2766,N_2431,N_2123);
and U2767 (N_2767,N_2472,N_2087);
nand U2768 (N_2768,N_2101,N_2100);
and U2769 (N_2769,N_2054,N_2454);
nand U2770 (N_2770,N_2460,N_2082);
nand U2771 (N_2771,N_2172,N_2226);
or U2772 (N_2772,N_2303,N_2062);
and U2773 (N_2773,N_2420,N_2036);
or U2774 (N_2774,N_2267,N_2007);
nand U2775 (N_2775,N_2182,N_2497);
and U2776 (N_2776,N_2160,N_2138);
xor U2777 (N_2777,N_2041,N_2306);
or U2778 (N_2778,N_2346,N_2277);
or U2779 (N_2779,N_2363,N_2167);
nand U2780 (N_2780,N_2306,N_2002);
and U2781 (N_2781,N_2059,N_2309);
nor U2782 (N_2782,N_2075,N_2449);
or U2783 (N_2783,N_2269,N_2383);
and U2784 (N_2784,N_2370,N_2142);
xor U2785 (N_2785,N_2157,N_2388);
nand U2786 (N_2786,N_2188,N_2028);
and U2787 (N_2787,N_2013,N_2340);
nor U2788 (N_2788,N_2344,N_2198);
nand U2789 (N_2789,N_2379,N_2029);
and U2790 (N_2790,N_2389,N_2164);
and U2791 (N_2791,N_2260,N_2227);
nand U2792 (N_2792,N_2074,N_2313);
and U2793 (N_2793,N_2228,N_2336);
nand U2794 (N_2794,N_2119,N_2369);
xor U2795 (N_2795,N_2275,N_2132);
nand U2796 (N_2796,N_2452,N_2412);
xnor U2797 (N_2797,N_2458,N_2058);
xor U2798 (N_2798,N_2374,N_2456);
and U2799 (N_2799,N_2387,N_2313);
and U2800 (N_2800,N_2302,N_2346);
xor U2801 (N_2801,N_2291,N_2272);
nor U2802 (N_2802,N_2114,N_2072);
nor U2803 (N_2803,N_2342,N_2386);
nand U2804 (N_2804,N_2352,N_2123);
nor U2805 (N_2805,N_2269,N_2340);
or U2806 (N_2806,N_2172,N_2273);
nand U2807 (N_2807,N_2486,N_2437);
or U2808 (N_2808,N_2010,N_2358);
nor U2809 (N_2809,N_2320,N_2428);
and U2810 (N_2810,N_2116,N_2284);
nand U2811 (N_2811,N_2114,N_2442);
or U2812 (N_2812,N_2405,N_2354);
or U2813 (N_2813,N_2035,N_2181);
nor U2814 (N_2814,N_2091,N_2430);
nor U2815 (N_2815,N_2291,N_2082);
or U2816 (N_2816,N_2241,N_2013);
nor U2817 (N_2817,N_2101,N_2429);
or U2818 (N_2818,N_2370,N_2091);
or U2819 (N_2819,N_2119,N_2330);
nor U2820 (N_2820,N_2367,N_2206);
and U2821 (N_2821,N_2205,N_2476);
nor U2822 (N_2822,N_2240,N_2361);
or U2823 (N_2823,N_2131,N_2300);
nand U2824 (N_2824,N_2044,N_2377);
and U2825 (N_2825,N_2279,N_2226);
nor U2826 (N_2826,N_2271,N_2120);
or U2827 (N_2827,N_2253,N_2071);
and U2828 (N_2828,N_2323,N_2074);
and U2829 (N_2829,N_2059,N_2394);
nor U2830 (N_2830,N_2172,N_2496);
nor U2831 (N_2831,N_2016,N_2461);
and U2832 (N_2832,N_2097,N_2071);
nand U2833 (N_2833,N_2437,N_2028);
nor U2834 (N_2834,N_2080,N_2013);
and U2835 (N_2835,N_2256,N_2214);
nor U2836 (N_2836,N_2240,N_2348);
nand U2837 (N_2837,N_2424,N_2185);
nor U2838 (N_2838,N_2227,N_2225);
and U2839 (N_2839,N_2022,N_2065);
xor U2840 (N_2840,N_2464,N_2280);
nor U2841 (N_2841,N_2038,N_2415);
nor U2842 (N_2842,N_2366,N_2174);
nand U2843 (N_2843,N_2074,N_2163);
nor U2844 (N_2844,N_2363,N_2339);
nor U2845 (N_2845,N_2303,N_2006);
and U2846 (N_2846,N_2446,N_2307);
nor U2847 (N_2847,N_2062,N_2230);
and U2848 (N_2848,N_2278,N_2044);
and U2849 (N_2849,N_2189,N_2467);
nand U2850 (N_2850,N_2018,N_2060);
nor U2851 (N_2851,N_2371,N_2443);
and U2852 (N_2852,N_2223,N_2087);
nand U2853 (N_2853,N_2031,N_2430);
nor U2854 (N_2854,N_2131,N_2410);
nor U2855 (N_2855,N_2347,N_2158);
nand U2856 (N_2856,N_2307,N_2253);
nand U2857 (N_2857,N_2132,N_2061);
xnor U2858 (N_2858,N_2047,N_2209);
or U2859 (N_2859,N_2380,N_2004);
nand U2860 (N_2860,N_2320,N_2069);
nor U2861 (N_2861,N_2447,N_2468);
and U2862 (N_2862,N_2146,N_2177);
or U2863 (N_2863,N_2284,N_2431);
and U2864 (N_2864,N_2269,N_2230);
xnor U2865 (N_2865,N_2497,N_2414);
nor U2866 (N_2866,N_2336,N_2292);
xor U2867 (N_2867,N_2472,N_2225);
and U2868 (N_2868,N_2301,N_2452);
xor U2869 (N_2869,N_2129,N_2291);
nand U2870 (N_2870,N_2030,N_2301);
nor U2871 (N_2871,N_2326,N_2134);
or U2872 (N_2872,N_2251,N_2266);
nor U2873 (N_2873,N_2126,N_2113);
nor U2874 (N_2874,N_2168,N_2045);
or U2875 (N_2875,N_2235,N_2297);
nor U2876 (N_2876,N_2266,N_2283);
or U2877 (N_2877,N_2497,N_2031);
nor U2878 (N_2878,N_2195,N_2212);
or U2879 (N_2879,N_2166,N_2103);
nor U2880 (N_2880,N_2025,N_2340);
or U2881 (N_2881,N_2305,N_2471);
and U2882 (N_2882,N_2148,N_2057);
nor U2883 (N_2883,N_2226,N_2155);
and U2884 (N_2884,N_2187,N_2407);
or U2885 (N_2885,N_2195,N_2099);
xnor U2886 (N_2886,N_2305,N_2350);
nor U2887 (N_2887,N_2132,N_2092);
nand U2888 (N_2888,N_2303,N_2330);
or U2889 (N_2889,N_2164,N_2140);
nor U2890 (N_2890,N_2015,N_2135);
nor U2891 (N_2891,N_2310,N_2283);
and U2892 (N_2892,N_2458,N_2415);
nor U2893 (N_2893,N_2303,N_2116);
nand U2894 (N_2894,N_2179,N_2162);
nor U2895 (N_2895,N_2290,N_2145);
and U2896 (N_2896,N_2243,N_2089);
and U2897 (N_2897,N_2332,N_2051);
and U2898 (N_2898,N_2255,N_2331);
nand U2899 (N_2899,N_2463,N_2293);
and U2900 (N_2900,N_2050,N_2418);
nand U2901 (N_2901,N_2072,N_2087);
nand U2902 (N_2902,N_2459,N_2406);
and U2903 (N_2903,N_2135,N_2438);
nor U2904 (N_2904,N_2100,N_2127);
nand U2905 (N_2905,N_2472,N_2497);
nand U2906 (N_2906,N_2052,N_2497);
or U2907 (N_2907,N_2059,N_2305);
or U2908 (N_2908,N_2387,N_2411);
nor U2909 (N_2909,N_2159,N_2042);
nand U2910 (N_2910,N_2102,N_2196);
or U2911 (N_2911,N_2113,N_2191);
nor U2912 (N_2912,N_2468,N_2257);
or U2913 (N_2913,N_2103,N_2291);
and U2914 (N_2914,N_2415,N_2334);
or U2915 (N_2915,N_2377,N_2190);
nand U2916 (N_2916,N_2397,N_2137);
or U2917 (N_2917,N_2397,N_2259);
nor U2918 (N_2918,N_2111,N_2304);
or U2919 (N_2919,N_2268,N_2189);
nor U2920 (N_2920,N_2009,N_2017);
or U2921 (N_2921,N_2096,N_2396);
nor U2922 (N_2922,N_2449,N_2034);
nand U2923 (N_2923,N_2051,N_2392);
xnor U2924 (N_2924,N_2335,N_2220);
nand U2925 (N_2925,N_2490,N_2336);
nand U2926 (N_2926,N_2214,N_2378);
or U2927 (N_2927,N_2460,N_2377);
or U2928 (N_2928,N_2381,N_2104);
and U2929 (N_2929,N_2408,N_2448);
or U2930 (N_2930,N_2479,N_2181);
or U2931 (N_2931,N_2448,N_2287);
nor U2932 (N_2932,N_2290,N_2130);
and U2933 (N_2933,N_2195,N_2138);
nand U2934 (N_2934,N_2237,N_2258);
xnor U2935 (N_2935,N_2063,N_2266);
or U2936 (N_2936,N_2232,N_2115);
xnor U2937 (N_2937,N_2418,N_2002);
and U2938 (N_2938,N_2359,N_2345);
and U2939 (N_2939,N_2253,N_2146);
nor U2940 (N_2940,N_2181,N_2130);
or U2941 (N_2941,N_2214,N_2382);
and U2942 (N_2942,N_2456,N_2465);
xor U2943 (N_2943,N_2495,N_2235);
nor U2944 (N_2944,N_2311,N_2114);
xnor U2945 (N_2945,N_2111,N_2038);
or U2946 (N_2946,N_2060,N_2059);
nand U2947 (N_2947,N_2146,N_2474);
nor U2948 (N_2948,N_2445,N_2239);
or U2949 (N_2949,N_2490,N_2386);
or U2950 (N_2950,N_2118,N_2223);
and U2951 (N_2951,N_2182,N_2071);
nand U2952 (N_2952,N_2413,N_2377);
or U2953 (N_2953,N_2269,N_2486);
and U2954 (N_2954,N_2354,N_2073);
nor U2955 (N_2955,N_2268,N_2323);
and U2956 (N_2956,N_2368,N_2098);
nand U2957 (N_2957,N_2068,N_2271);
xor U2958 (N_2958,N_2491,N_2472);
and U2959 (N_2959,N_2382,N_2204);
nor U2960 (N_2960,N_2380,N_2233);
and U2961 (N_2961,N_2481,N_2382);
nor U2962 (N_2962,N_2413,N_2113);
nor U2963 (N_2963,N_2283,N_2293);
nor U2964 (N_2964,N_2287,N_2389);
xnor U2965 (N_2965,N_2485,N_2496);
and U2966 (N_2966,N_2219,N_2298);
nand U2967 (N_2967,N_2034,N_2114);
and U2968 (N_2968,N_2397,N_2191);
and U2969 (N_2969,N_2186,N_2475);
and U2970 (N_2970,N_2223,N_2314);
nand U2971 (N_2971,N_2375,N_2485);
and U2972 (N_2972,N_2186,N_2122);
nor U2973 (N_2973,N_2072,N_2263);
nand U2974 (N_2974,N_2321,N_2367);
nor U2975 (N_2975,N_2291,N_2215);
or U2976 (N_2976,N_2406,N_2442);
and U2977 (N_2977,N_2258,N_2333);
xor U2978 (N_2978,N_2233,N_2479);
nor U2979 (N_2979,N_2363,N_2182);
nor U2980 (N_2980,N_2327,N_2243);
nor U2981 (N_2981,N_2489,N_2370);
nor U2982 (N_2982,N_2250,N_2236);
and U2983 (N_2983,N_2345,N_2115);
and U2984 (N_2984,N_2086,N_2136);
nor U2985 (N_2985,N_2440,N_2180);
nand U2986 (N_2986,N_2272,N_2178);
nor U2987 (N_2987,N_2339,N_2345);
nand U2988 (N_2988,N_2232,N_2368);
or U2989 (N_2989,N_2458,N_2190);
and U2990 (N_2990,N_2451,N_2472);
and U2991 (N_2991,N_2072,N_2399);
xnor U2992 (N_2992,N_2349,N_2313);
nor U2993 (N_2993,N_2461,N_2261);
or U2994 (N_2994,N_2095,N_2173);
and U2995 (N_2995,N_2224,N_2265);
xnor U2996 (N_2996,N_2421,N_2167);
or U2997 (N_2997,N_2406,N_2078);
and U2998 (N_2998,N_2315,N_2038);
nor U2999 (N_2999,N_2442,N_2244);
and U3000 (N_3000,N_2853,N_2778);
nor U3001 (N_3001,N_2733,N_2550);
nand U3002 (N_3002,N_2839,N_2798);
nand U3003 (N_3003,N_2593,N_2732);
xnor U3004 (N_3004,N_2789,N_2634);
and U3005 (N_3005,N_2785,N_2511);
nor U3006 (N_3006,N_2840,N_2714);
or U3007 (N_3007,N_2543,N_2862);
or U3008 (N_3008,N_2501,N_2705);
and U3009 (N_3009,N_2812,N_2804);
nor U3010 (N_3010,N_2808,N_2528);
nand U3011 (N_3011,N_2612,N_2775);
nor U3012 (N_3012,N_2925,N_2906);
nand U3013 (N_3013,N_2769,N_2773);
nand U3014 (N_3014,N_2751,N_2841);
and U3015 (N_3015,N_2629,N_2558);
xnor U3016 (N_3016,N_2847,N_2968);
and U3017 (N_3017,N_2996,N_2577);
or U3018 (N_3018,N_2943,N_2991);
and U3019 (N_3019,N_2663,N_2805);
xor U3020 (N_3020,N_2843,N_2615);
nand U3021 (N_3021,N_2519,N_2890);
or U3022 (N_3022,N_2931,N_2692);
nor U3023 (N_3023,N_2978,N_2573);
or U3024 (N_3024,N_2831,N_2693);
nor U3025 (N_3025,N_2706,N_2971);
nand U3026 (N_3026,N_2886,N_2622);
or U3027 (N_3027,N_2707,N_2761);
nor U3028 (N_3028,N_2608,N_2735);
nor U3029 (N_3029,N_2837,N_2635);
nor U3030 (N_3030,N_2688,N_2517);
or U3031 (N_3031,N_2649,N_2810);
nor U3032 (N_3032,N_2913,N_2620);
nand U3033 (N_3033,N_2796,N_2950);
nand U3034 (N_3034,N_2855,N_2587);
nand U3035 (N_3035,N_2594,N_2532);
nor U3036 (N_3036,N_2763,N_2907);
nand U3037 (N_3037,N_2894,N_2514);
nor U3038 (N_3038,N_2788,N_2530);
or U3039 (N_3039,N_2526,N_2901);
or U3040 (N_3040,N_2835,N_2570);
and U3041 (N_3041,N_2624,N_2562);
and U3042 (N_3042,N_2586,N_2874);
and U3043 (N_3043,N_2680,N_2818);
nand U3044 (N_3044,N_2630,N_2986);
nor U3045 (N_3045,N_2613,N_2740);
and U3046 (N_3046,N_2914,N_2569);
and U3047 (N_3047,N_2975,N_2916);
nor U3048 (N_3048,N_2784,N_2933);
nand U3049 (N_3049,N_2972,N_2786);
and U3050 (N_3050,N_2934,N_2701);
and U3051 (N_3051,N_2891,N_2552);
and U3052 (N_3052,N_2523,N_2736);
or U3053 (N_3053,N_2849,N_2961);
or U3054 (N_3054,N_2538,N_2540);
nand U3055 (N_3055,N_2715,N_2670);
or U3056 (N_3056,N_2844,N_2506);
nand U3057 (N_3057,N_2604,N_2529);
nand U3058 (N_3058,N_2960,N_2883);
nor U3059 (N_3059,N_2505,N_2524);
nor U3060 (N_3060,N_2800,N_2994);
or U3061 (N_3061,N_2926,N_2783);
or U3062 (N_3062,N_2721,N_2713);
and U3063 (N_3063,N_2534,N_2575);
nor U3064 (N_3064,N_2762,N_2557);
xor U3065 (N_3065,N_2776,N_2957);
and U3066 (N_3066,N_2730,N_2589);
or U3067 (N_3067,N_2754,N_2878);
xor U3068 (N_3068,N_2921,N_2584);
and U3069 (N_3069,N_2610,N_2764);
and U3070 (N_3070,N_2691,N_2774);
nand U3071 (N_3071,N_2621,N_2669);
or U3072 (N_3072,N_2535,N_2806);
xnor U3073 (N_3073,N_2899,N_2625);
and U3074 (N_3074,N_2865,N_2728);
or U3075 (N_3075,N_2606,N_2507);
nand U3076 (N_3076,N_2823,N_2866);
nand U3077 (N_3077,N_2725,N_2709);
nand U3078 (N_3078,N_2717,N_2545);
or U3079 (N_3079,N_2537,N_2675);
nand U3080 (N_3080,N_2869,N_2859);
or U3081 (N_3081,N_2718,N_2565);
or U3082 (N_3082,N_2903,N_2690);
nand U3083 (N_3083,N_2563,N_2574);
nor U3084 (N_3084,N_2851,N_2820);
or U3085 (N_3085,N_2790,N_2739);
or U3086 (N_3086,N_2516,N_2898);
or U3087 (N_3087,N_2908,N_2932);
or U3088 (N_3088,N_2568,N_2902);
and U3089 (N_3089,N_2638,N_2581);
or U3090 (N_3090,N_2640,N_2989);
nand U3091 (N_3091,N_2602,N_2973);
nand U3092 (N_3092,N_2611,N_2567);
nand U3093 (N_3093,N_2648,N_2928);
nand U3094 (N_3094,N_2845,N_2734);
nand U3095 (N_3095,N_2647,N_2860);
or U3096 (N_3096,N_2527,N_2665);
and U3097 (N_3097,N_2920,N_2927);
nor U3098 (N_3098,N_2503,N_2544);
and U3099 (N_3099,N_2904,N_2814);
xor U3100 (N_3100,N_2546,N_2885);
xor U3101 (N_3101,N_2689,N_2872);
or U3102 (N_3102,N_2864,N_2828);
nand U3103 (N_3103,N_2681,N_2678);
nand U3104 (N_3104,N_2875,N_2645);
nor U3105 (N_3105,N_2836,N_2623);
and U3106 (N_3106,N_2937,N_2838);
nor U3107 (N_3107,N_2876,N_2958);
or U3108 (N_3108,N_2772,N_2609);
or U3109 (N_3109,N_2664,N_2848);
and U3110 (N_3110,N_2826,N_2755);
or U3111 (N_3111,N_2905,N_2659);
nor U3112 (N_3112,N_2564,N_2591);
nor U3113 (N_3113,N_2795,N_2935);
and U3114 (N_3114,N_2737,N_2652);
and U3115 (N_3115,N_2852,N_2504);
and U3116 (N_3116,N_2533,N_2520);
or U3117 (N_3117,N_2671,N_2854);
nand U3118 (N_3118,N_2997,N_2555);
nor U3119 (N_3119,N_2953,N_2909);
nor U3120 (N_3120,N_2787,N_2742);
nand U3121 (N_3121,N_2596,N_2666);
nand U3122 (N_3122,N_2607,N_2792);
nor U3123 (N_3123,N_2977,N_2939);
nor U3124 (N_3124,N_2729,N_2551);
nor U3125 (N_3125,N_2633,N_2676);
nor U3126 (N_3126,N_2745,N_2618);
xor U3127 (N_3127,N_2830,N_2576);
or U3128 (N_3128,N_2767,N_2873);
xor U3129 (N_3129,N_2685,N_2871);
or U3130 (N_3130,N_2896,N_2897);
nor U3131 (N_3131,N_2829,N_2768);
nand U3132 (N_3132,N_2992,N_2547);
and U3133 (N_3133,N_2657,N_2821);
nor U3134 (N_3134,N_2879,N_2702);
and U3135 (N_3135,N_2695,N_2601);
xnor U3136 (N_3136,N_2964,N_2794);
nand U3137 (N_3137,N_2779,N_2956);
nor U3138 (N_3138,N_2893,N_2756);
or U3139 (N_3139,N_2797,N_2915);
or U3140 (N_3140,N_2556,N_2868);
and U3141 (N_3141,N_2616,N_2674);
and U3142 (N_3142,N_2811,N_2753);
nand U3143 (N_3143,N_2655,N_2880);
nand U3144 (N_3144,N_2936,N_2982);
nand U3145 (N_3145,N_2832,N_2700);
and U3146 (N_3146,N_2605,N_2765);
or U3147 (N_3147,N_2566,N_2910);
xnor U3148 (N_3148,N_2703,N_2815);
nand U3149 (N_3149,N_2819,N_2770);
nand U3150 (N_3150,N_2636,N_2749);
or U3151 (N_3151,N_2791,N_2870);
xor U3152 (N_3152,N_2747,N_2541);
nor U3153 (N_3153,N_2863,N_2580);
xnor U3154 (N_3154,N_2882,N_2627);
and U3155 (N_3155,N_2578,N_2807);
and U3156 (N_3156,N_2799,N_2599);
nand U3157 (N_3157,N_2661,N_2881);
nor U3158 (N_3158,N_2827,N_2962);
and U3159 (N_3159,N_2628,N_2919);
and U3160 (N_3160,N_2559,N_2757);
nor U3161 (N_3161,N_2743,N_2603);
nor U3162 (N_3162,N_2549,N_2704);
nor U3163 (N_3163,N_2637,N_2597);
xnor U3164 (N_3164,N_2766,N_2752);
nor U3165 (N_3165,N_2720,N_2656);
and U3166 (N_3166,N_2738,N_2900);
or U3167 (N_3167,N_2641,N_2833);
or U3168 (N_3168,N_2710,N_2824);
nor U3169 (N_3169,N_2646,N_2942);
or U3170 (N_3170,N_2698,N_2583);
nand U3171 (N_3171,N_2711,N_2946);
nand U3172 (N_3172,N_2887,N_2758);
xor U3173 (N_3173,N_2748,N_2508);
nand U3174 (N_3174,N_2662,N_2554);
xor U3175 (N_3175,N_2782,N_2995);
nor U3176 (N_3176,N_2781,N_2502);
or U3177 (N_3177,N_2561,N_2944);
and U3178 (N_3178,N_2974,N_2917);
xor U3179 (N_3179,N_2941,N_2817);
nor U3180 (N_3180,N_2912,N_2858);
or U3181 (N_3181,N_2726,N_2697);
or U3182 (N_3182,N_2500,N_2512);
or U3183 (N_3183,N_2809,N_2983);
and U3184 (N_3184,N_2684,N_2619);
xor U3185 (N_3185,N_2677,N_2553);
and U3186 (N_3186,N_2572,N_2571);
or U3187 (N_3187,N_2813,N_2780);
xnor U3188 (N_3188,N_2643,N_2988);
and U3189 (N_3189,N_2667,N_2803);
nor U3190 (N_3190,N_2970,N_2585);
and U3191 (N_3191,N_2683,N_2948);
nor U3192 (N_3192,N_2531,N_2724);
or U3193 (N_3193,N_2746,N_2539);
nand U3194 (N_3194,N_2642,N_2548);
xnor U3195 (N_3195,N_2639,N_2509);
or U3196 (N_3196,N_2966,N_2842);
or U3197 (N_3197,N_2708,N_2595);
nor U3198 (N_3198,N_2825,N_2522);
and U3199 (N_3199,N_2600,N_2632);
and U3200 (N_3200,N_2727,N_2687);
nand U3201 (N_3201,N_2981,N_2861);
nor U3202 (N_3202,N_2521,N_2918);
nand U3203 (N_3203,N_2967,N_2955);
xor U3204 (N_3204,N_2617,N_2985);
nand U3205 (N_3205,N_2686,N_2949);
xor U3206 (N_3206,N_2771,N_2923);
and U3207 (N_3207,N_2987,N_2679);
nand U3208 (N_3208,N_2682,N_2895);
nand U3209 (N_3209,N_2938,N_2924);
and U3210 (N_3210,N_2802,N_2979);
or U3211 (N_3211,N_2990,N_2660);
nand U3212 (N_3212,N_2930,N_2536);
xor U3213 (N_3213,N_2614,N_2889);
xnor U3214 (N_3214,N_2696,N_2582);
nor U3215 (N_3215,N_2750,N_2963);
or U3216 (N_3216,N_2984,N_2947);
and U3217 (N_3217,N_2888,N_2525);
and U3218 (N_3218,N_2976,N_2510);
or U3219 (N_3219,N_2651,N_2712);
nor U3220 (N_3220,N_2644,N_2654);
or U3221 (N_3221,N_2945,N_2694);
and U3222 (N_3222,N_2969,N_2884);
and U3223 (N_3223,N_2598,N_2759);
nand U3224 (N_3224,N_2653,N_2513);
nand U3225 (N_3225,N_2965,N_2560);
and U3226 (N_3226,N_2959,N_2744);
and U3227 (N_3227,N_2999,N_2542);
and U3228 (N_3228,N_2857,N_2892);
or U3229 (N_3229,N_2911,N_2816);
nor U3230 (N_3230,N_2951,N_2631);
nor U3231 (N_3231,N_2777,N_2626);
and U3232 (N_3232,N_2673,N_2723);
nand U3233 (N_3233,N_2722,N_2515);
and U3234 (N_3234,N_2856,N_2793);
or U3235 (N_3235,N_2760,N_2834);
nor U3236 (N_3236,N_2867,N_2929);
xnor U3237 (N_3237,N_2952,N_2822);
nand U3238 (N_3238,N_2846,N_2998);
nand U3239 (N_3239,N_2650,N_2741);
or U3240 (N_3240,N_2922,N_2801);
nand U3241 (N_3241,N_2850,N_2940);
nand U3242 (N_3242,N_2877,N_2590);
nor U3243 (N_3243,N_2579,N_2518);
nor U3244 (N_3244,N_2980,N_2719);
nand U3245 (N_3245,N_2658,N_2993);
xnor U3246 (N_3246,N_2731,N_2716);
nor U3247 (N_3247,N_2588,N_2699);
nand U3248 (N_3248,N_2592,N_2954);
nand U3249 (N_3249,N_2668,N_2672);
and U3250 (N_3250,N_2824,N_2995);
or U3251 (N_3251,N_2754,N_2852);
nor U3252 (N_3252,N_2725,N_2930);
and U3253 (N_3253,N_2544,N_2687);
nor U3254 (N_3254,N_2672,N_2917);
or U3255 (N_3255,N_2514,N_2619);
nor U3256 (N_3256,N_2750,N_2578);
and U3257 (N_3257,N_2581,N_2869);
nand U3258 (N_3258,N_2687,N_2838);
nor U3259 (N_3259,N_2759,N_2568);
nand U3260 (N_3260,N_2645,N_2989);
nand U3261 (N_3261,N_2858,N_2789);
or U3262 (N_3262,N_2635,N_2826);
nor U3263 (N_3263,N_2612,N_2815);
and U3264 (N_3264,N_2696,N_2546);
nor U3265 (N_3265,N_2610,N_2883);
nor U3266 (N_3266,N_2985,N_2508);
nor U3267 (N_3267,N_2970,N_2835);
and U3268 (N_3268,N_2559,N_2523);
nand U3269 (N_3269,N_2747,N_2740);
xnor U3270 (N_3270,N_2690,N_2808);
and U3271 (N_3271,N_2634,N_2915);
nor U3272 (N_3272,N_2742,N_2898);
nand U3273 (N_3273,N_2523,N_2934);
and U3274 (N_3274,N_2905,N_2701);
and U3275 (N_3275,N_2629,N_2572);
nor U3276 (N_3276,N_2599,N_2825);
nand U3277 (N_3277,N_2605,N_2735);
and U3278 (N_3278,N_2979,N_2801);
nand U3279 (N_3279,N_2807,N_2592);
or U3280 (N_3280,N_2546,N_2759);
and U3281 (N_3281,N_2768,N_2507);
nand U3282 (N_3282,N_2681,N_2724);
nor U3283 (N_3283,N_2845,N_2868);
nand U3284 (N_3284,N_2870,N_2612);
nor U3285 (N_3285,N_2756,N_2818);
or U3286 (N_3286,N_2589,N_2664);
or U3287 (N_3287,N_2623,N_2718);
or U3288 (N_3288,N_2965,N_2983);
nand U3289 (N_3289,N_2587,N_2558);
nor U3290 (N_3290,N_2788,N_2898);
or U3291 (N_3291,N_2523,N_2774);
nor U3292 (N_3292,N_2797,N_2830);
xnor U3293 (N_3293,N_2811,N_2981);
nand U3294 (N_3294,N_2700,N_2613);
nand U3295 (N_3295,N_2504,N_2748);
xor U3296 (N_3296,N_2774,N_2712);
nor U3297 (N_3297,N_2801,N_2729);
nand U3298 (N_3298,N_2957,N_2975);
or U3299 (N_3299,N_2701,N_2762);
nor U3300 (N_3300,N_2998,N_2990);
and U3301 (N_3301,N_2568,N_2637);
and U3302 (N_3302,N_2659,N_2676);
and U3303 (N_3303,N_2707,N_2811);
or U3304 (N_3304,N_2722,N_2551);
and U3305 (N_3305,N_2803,N_2940);
and U3306 (N_3306,N_2853,N_2675);
nand U3307 (N_3307,N_2745,N_2967);
or U3308 (N_3308,N_2692,N_2544);
nand U3309 (N_3309,N_2896,N_2660);
nor U3310 (N_3310,N_2523,N_2782);
nand U3311 (N_3311,N_2929,N_2568);
xnor U3312 (N_3312,N_2841,N_2863);
and U3313 (N_3313,N_2776,N_2711);
and U3314 (N_3314,N_2558,N_2638);
nand U3315 (N_3315,N_2779,N_2995);
nor U3316 (N_3316,N_2744,N_2606);
nand U3317 (N_3317,N_2853,N_2547);
or U3318 (N_3318,N_2860,N_2720);
and U3319 (N_3319,N_2812,N_2519);
and U3320 (N_3320,N_2716,N_2588);
or U3321 (N_3321,N_2818,N_2585);
nand U3322 (N_3322,N_2948,N_2913);
nand U3323 (N_3323,N_2968,N_2988);
nand U3324 (N_3324,N_2865,N_2647);
or U3325 (N_3325,N_2851,N_2996);
nand U3326 (N_3326,N_2887,N_2982);
and U3327 (N_3327,N_2639,N_2520);
nand U3328 (N_3328,N_2862,N_2975);
and U3329 (N_3329,N_2632,N_2584);
xor U3330 (N_3330,N_2750,N_2898);
nand U3331 (N_3331,N_2615,N_2946);
and U3332 (N_3332,N_2855,N_2718);
and U3333 (N_3333,N_2990,N_2845);
and U3334 (N_3334,N_2991,N_2969);
and U3335 (N_3335,N_2762,N_2829);
nor U3336 (N_3336,N_2896,N_2669);
or U3337 (N_3337,N_2552,N_2774);
nand U3338 (N_3338,N_2927,N_2703);
or U3339 (N_3339,N_2791,N_2933);
nand U3340 (N_3340,N_2687,N_2705);
xor U3341 (N_3341,N_2722,N_2804);
xnor U3342 (N_3342,N_2616,N_2833);
nand U3343 (N_3343,N_2710,N_2807);
nand U3344 (N_3344,N_2775,N_2709);
nor U3345 (N_3345,N_2966,N_2721);
xor U3346 (N_3346,N_2594,N_2848);
or U3347 (N_3347,N_2536,N_2677);
and U3348 (N_3348,N_2967,N_2637);
and U3349 (N_3349,N_2628,N_2788);
or U3350 (N_3350,N_2501,N_2531);
or U3351 (N_3351,N_2751,N_2538);
and U3352 (N_3352,N_2807,N_2771);
nor U3353 (N_3353,N_2574,N_2912);
and U3354 (N_3354,N_2690,N_2528);
nor U3355 (N_3355,N_2771,N_2635);
nand U3356 (N_3356,N_2994,N_2720);
and U3357 (N_3357,N_2901,N_2620);
nand U3358 (N_3358,N_2514,N_2637);
xnor U3359 (N_3359,N_2690,N_2961);
xor U3360 (N_3360,N_2607,N_2723);
and U3361 (N_3361,N_2623,N_2862);
or U3362 (N_3362,N_2606,N_2826);
and U3363 (N_3363,N_2939,N_2918);
and U3364 (N_3364,N_2653,N_2918);
nor U3365 (N_3365,N_2532,N_2694);
xnor U3366 (N_3366,N_2524,N_2964);
or U3367 (N_3367,N_2754,N_2811);
nor U3368 (N_3368,N_2646,N_2795);
xor U3369 (N_3369,N_2796,N_2907);
nand U3370 (N_3370,N_2878,N_2795);
nand U3371 (N_3371,N_2988,N_2950);
nand U3372 (N_3372,N_2972,N_2804);
xor U3373 (N_3373,N_2568,N_2895);
nor U3374 (N_3374,N_2954,N_2568);
or U3375 (N_3375,N_2854,N_2826);
nand U3376 (N_3376,N_2502,N_2734);
xor U3377 (N_3377,N_2956,N_2981);
nand U3378 (N_3378,N_2863,N_2874);
nor U3379 (N_3379,N_2516,N_2963);
nor U3380 (N_3380,N_2500,N_2994);
or U3381 (N_3381,N_2670,N_2687);
nor U3382 (N_3382,N_2936,N_2586);
or U3383 (N_3383,N_2531,N_2551);
nor U3384 (N_3384,N_2763,N_2661);
nor U3385 (N_3385,N_2876,N_2949);
and U3386 (N_3386,N_2605,N_2843);
nand U3387 (N_3387,N_2994,N_2504);
xor U3388 (N_3388,N_2772,N_2537);
or U3389 (N_3389,N_2948,N_2704);
nand U3390 (N_3390,N_2744,N_2937);
nand U3391 (N_3391,N_2555,N_2549);
nor U3392 (N_3392,N_2771,N_2688);
nor U3393 (N_3393,N_2710,N_2652);
xor U3394 (N_3394,N_2644,N_2578);
or U3395 (N_3395,N_2776,N_2741);
xor U3396 (N_3396,N_2954,N_2716);
nor U3397 (N_3397,N_2853,N_2558);
nand U3398 (N_3398,N_2845,N_2944);
nor U3399 (N_3399,N_2918,N_2503);
xnor U3400 (N_3400,N_2563,N_2681);
nand U3401 (N_3401,N_2977,N_2955);
nor U3402 (N_3402,N_2666,N_2509);
nand U3403 (N_3403,N_2881,N_2771);
or U3404 (N_3404,N_2882,N_2895);
xnor U3405 (N_3405,N_2919,N_2697);
xnor U3406 (N_3406,N_2577,N_2989);
nor U3407 (N_3407,N_2950,N_2846);
nor U3408 (N_3408,N_2977,N_2518);
or U3409 (N_3409,N_2700,N_2583);
nor U3410 (N_3410,N_2707,N_2976);
nor U3411 (N_3411,N_2631,N_2830);
and U3412 (N_3412,N_2729,N_2560);
nand U3413 (N_3413,N_2543,N_2610);
nand U3414 (N_3414,N_2718,N_2899);
and U3415 (N_3415,N_2826,N_2915);
nand U3416 (N_3416,N_2927,N_2903);
nor U3417 (N_3417,N_2882,N_2808);
nand U3418 (N_3418,N_2558,N_2593);
xnor U3419 (N_3419,N_2594,N_2723);
xnor U3420 (N_3420,N_2505,N_2815);
nor U3421 (N_3421,N_2879,N_2783);
nand U3422 (N_3422,N_2833,N_2705);
nor U3423 (N_3423,N_2842,N_2604);
nor U3424 (N_3424,N_2779,N_2545);
and U3425 (N_3425,N_2897,N_2858);
nor U3426 (N_3426,N_2639,N_2710);
or U3427 (N_3427,N_2648,N_2539);
or U3428 (N_3428,N_2647,N_2594);
nor U3429 (N_3429,N_2560,N_2656);
nor U3430 (N_3430,N_2826,N_2597);
nor U3431 (N_3431,N_2555,N_2702);
xor U3432 (N_3432,N_2519,N_2669);
nor U3433 (N_3433,N_2565,N_2741);
or U3434 (N_3434,N_2727,N_2712);
and U3435 (N_3435,N_2775,N_2946);
or U3436 (N_3436,N_2903,N_2854);
nand U3437 (N_3437,N_2723,N_2638);
xor U3438 (N_3438,N_2526,N_2931);
or U3439 (N_3439,N_2509,N_2570);
and U3440 (N_3440,N_2884,N_2757);
and U3441 (N_3441,N_2777,N_2837);
nor U3442 (N_3442,N_2639,N_2516);
or U3443 (N_3443,N_2982,N_2987);
nor U3444 (N_3444,N_2929,N_2596);
nor U3445 (N_3445,N_2877,N_2632);
and U3446 (N_3446,N_2828,N_2935);
nor U3447 (N_3447,N_2934,N_2969);
nor U3448 (N_3448,N_2965,N_2648);
and U3449 (N_3449,N_2573,N_2768);
nand U3450 (N_3450,N_2898,N_2888);
and U3451 (N_3451,N_2775,N_2975);
nand U3452 (N_3452,N_2891,N_2651);
nor U3453 (N_3453,N_2630,N_2887);
nor U3454 (N_3454,N_2866,N_2646);
nand U3455 (N_3455,N_2803,N_2653);
xnor U3456 (N_3456,N_2508,N_2909);
and U3457 (N_3457,N_2728,N_2700);
xnor U3458 (N_3458,N_2915,N_2588);
nand U3459 (N_3459,N_2627,N_2892);
or U3460 (N_3460,N_2671,N_2866);
or U3461 (N_3461,N_2876,N_2991);
nor U3462 (N_3462,N_2683,N_2600);
nor U3463 (N_3463,N_2709,N_2729);
nand U3464 (N_3464,N_2885,N_2815);
nor U3465 (N_3465,N_2897,N_2578);
or U3466 (N_3466,N_2890,N_2920);
or U3467 (N_3467,N_2703,N_2952);
nand U3468 (N_3468,N_2858,N_2948);
nand U3469 (N_3469,N_2670,N_2523);
nor U3470 (N_3470,N_2712,N_2697);
xor U3471 (N_3471,N_2696,N_2715);
and U3472 (N_3472,N_2647,N_2511);
nand U3473 (N_3473,N_2708,N_2787);
and U3474 (N_3474,N_2901,N_2612);
and U3475 (N_3475,N_2817,N_2660);
xor U3476 (N_3476,N_2535,N_2872);
nand U3477 (N_3477,N_2772,N_2581);
nand U3478 (N_3478,N_2840,N_2730);
nor U3479 (N_3479,N_2869,N_2750);
nor U3480 (N_3480,N_2991,N_2691);
nand U3481 (N_3481,N_2608,N_2802);
or U3482 (N_3482,N_2858,N_2859);
nor U3483 (N_3483,N_2677,N_2818);
nand U3484 (N_3484,N_2680,N_2611);
or U3485 (N_3485,N_2684,N_2972);
nor U3486 (N_3486,N_2543,N_2545);
and U3487 (N_3487,N_2872,N_2824);
and U3488 (N_3488,N_2993,N_2973);
and U3489 (N_3489,N_2970,N_2997);
nor U3490 (N_3490,N_2849,N_2693);
or U3491 (N_3491,N_2900,N_2961);
or U3492 (N_3492,N_2769,N_2629);
nor U3493 (N_3493,N_2703,N_2749);
and U3494 (N_3494,N_2752,N_2744);
nand U3495 (N_3495,N_2621,N_2715);
and U3496 (N_3496,N_2927,N_2504);
nand U3497 (N_3497,N_2503,N_2638);
nor U3498 (N_3498,N_2730,N_2911);
xor U3499 (N_3499,N_2670,N_2877);
nor U3500 (N_3500,N_3267,N_3184);
nor U3501 (N_3501,N_3341,N_3284);
nor U3502 (N_3502,N_3066,N_3421);
or U3503 (N_3503,N_3114,N_3166);
nor U3504 (N_3504,N_3440,N_3151);
or U3505 (N_3505,N_3357,N_3343);
or U3506 (N_3506,N_3461,N_3288);
or U3507 (N_3507,N_3479,N_3367);
and U3508 (N_3508,N_3067,N_3350);
nor U3509 (N_3509,N_3282,N_3306);
or U3510 (N_3510,N_3108,N_3331);
nor U3511 (N_3511,N_3059,N_3415);
xor U3512 (N_3512,N_3434,N_3293);
nor U3513 (N_3513,N_3241,N_3125);
xor U3514 (N_3514,N_3443,N_3477);
and U3515 (N_3515,N_3314,N_3140);
nor U3516 (N_3516,N_3061,N_3130);
nor U3517 (N_3517,N_3433,N_3080);
nand U3518 (N_3518,N_3002,N_3397);
and U3519 (N_3519,N_3276,N_3418);
nand U3520 (N_3520,N_3329,N_3243);
xor U3521 (N_3521,N_3024,N_3322);
nor U3522 (N_3522,N_3225,N_3386);
or U3523 (N_3523,N_3469,N_3256);
or U3524 (N_3524,N_3044,N_3152);
nor U3525 (N_3525,N_3129,N_3368);
nand U3526 (N_3526,N_3218,N_3029);
nand U3527 (N_3527,N_3013,N_3320);
nand U3528 (N_3528,N_3192,N_3003);
nor U3529 (N_3529,N_3348,N_3191);
nand U3530 (N_3530,N_3064,N_3233);
nor U3531 (N_3531,N_3285,N_3011);
and U3532 (N_3532,N_3212,N_3197);
nor U3533 (N_3533,N_3303,N_3045);
or U3534 (N_3534,N_3253,N_3091);
or U3535 (N_3535,N_3093,N_3336);
xor U3536 (N_3536,N_3100,N_3422);
or U3537 (N_3537,N_3221,N_3112);
nor U3538 (N_3538,N_3297,N_3056);
or U3539 (N_3539,N_3416,N_3424);
and U3540 (N_3540,N_3473,N_3089);
or U3541 (N_3541,N_3312,N_3131);
nor U3542 (N_3542,N_3485,N_3326);
nor U3543 (N_3543,N_3070,N_3370);
nand U3544 (N_3544,N_3387,N_3224);
nor U3545 (N_3545,N_3120,N_3196);
or U3546 (N_3546,N_3028,N_3385);
or U3547 (N_3547,N_3475,N_3085);
and U3548 (N_3548,N_3279,N_3301);
xnor U3549 (N_3549,N_3337,N_3481);
or U3550 (N_3550,N_3082,N_3441);
nor U3551 (N_3551,N_3174,N_3142);
and U3552 (N_3552,N_3173,N_3194);
nand U3553 (N_3553,N_3018,N_3496);
and U3554 (N_3554,N_3217,N_3380);
or U3555 (N_3555,N_3494,N_3497);
or U3556 (N_3556,N_3261,N_3262);
nand U3557 (N_3557,N_3170,N_3404);
and U3558 (N_3558,N_3292,N_3396);
nor U3559 (N_3559,N_3086,N_3209);
nand U3560 (N_3560,N_3203,N_3403);
nor U3561 (N_3561,N_3081,N_3451);
and U3562 (N_3562,N_3156,N_3169);
and U3563 (N_3563,N_3417,N_3258);
nand U3564 (N_3564,N_3486,N_3283);
and U3565 (N_3565,N_3406,N_3153);
and U3566 (N_3566,N_3049,N_3340);
or U3567 (N_3567,N_3269,N_3090);
nand U3568 (N_3568,N_3408,N_3210);
and U3569 (N_3569,N_3448,N_3105);
and U3570 (N_3570,N_3239,N_3004);
nand U3571 (N_3571,N_3150,N_3463);
nand U3572 (N_3572,N_3182,N_3458);
and U3573 (N_3573,N_3495,N_3400);
or U3574 (N_3574,N_3157,N_3489);
xnor U3575 (N_3575,N_3007,N_3374);
nand U3576 (N_3576,N_3155,N_3286);
and U3577 (N_3577,N_3316,N_3015);
or U3578 (N_3578,N_3391,N_3001);
and U3579 (N_3579,N_3035,N_3206);
or U3580 (N_3580,N_3117,N_3077);
or U3581 (N_3581,N_3470,N_3447);
or U3582 (N_3582,N_3345,N_3071);
and U3583 (N_3583,N_3296,N_3446);
nand U3584 (N_3584,N_3321,N_3493);
xor U3585 (N_3585,N_3144,N_3094);
or U3586 (N_3586,N_3058,N_3092);
and U3587 (N_3587,N_3228,N_3299);
and U3588 (N_3588,N_3216,N_3298);
or U3589 (N_3589,N_3278,N_3222);
and U3590 (N_3590,N_3020,N_3188);
and U3591 (N_3591,N_3444,N_3232);
and U3592 (N_3592,N_3214,N_3275);
nor U3593 (N_3593,N_3402,N_3236);
and U3594 (N_3594,N_3038,N_3344);
and U3595 (N_3595,N_3375,N_3005);
and U3596 (N_3596,N_3354,N_3043);
and U3597 (N_3597,N_3355,N_3146);
and U3598 (N_3598,N_3454,N_3022);
or U3599 (N_3599,N_3250,N_3290);
or U3600 (N_3600,N_3132,N_3145);
nor U3601 (N_3601,N_3468,N_3484);
or U3602 (N_3602,N_3136,N_3181);
xor U3603 (N_3603,N_3229,N_3358);
nor U3604 (N_3604,N_3010,N_3478);
nand U3605 (N_3605,N_3462,N_3054);
or U3606 (N_3606,N_3069,N_3376);
or U3607 (N_3607,N_3378,N_3442);
nor U3608 (N_3608,N_3012,N_3420);
nand U3609 (N_3609,N_3323,N_3041);
nor U3610 (N_3610,N_3488,N_3052);
nand U3611 (N_3611,N_3180,N_3167);
or U3612 (N_3612,N_3172,N_3338);
xnor U3613 (N_3613,N_3472,N_3234);
or U3614 (N_3614,N_3356,N_3393);
nor U3615 (N_3615,N_3128,N_3096);
nand U3616 (N_3616,N_3245,N_3074);
xor U3617 (N_3617,N_3088,N_3017);
xor U3618 (N_3618,N_3110,N_3466);
or U3619 (N_3619,N_3425,N_3289);
nand U3620 (N_3620,N_3242,N_3366);
nand U3621 (N_3621,N_3102,N_3154);
and U3622 (N_3622,N_3474,N_3023);
or U3623 (N_3623,N_3265,N_3411);
nor U3624 (N_3624,N_3464,N_3349);
xnor U3625 (N_3625,N_3310,N_3491);
nand U3626 (N_3626,N_3032,N_3377);
or U3627 (N_3627,N_3240,N_3309);
and U3628 (N_3628,N_3042,N_3359);
nor U3629 (N_3629,N_3270,N_3414);
nor U3630 (N_3630,N_3457,N_3099);
xor U3631 (N_3631,N_3383,N_3268);
and U3632 (N_3632,N_3437,N_3025);
or U3633 (N_3633,N_3249,N_3302);
and U3634 (N_3634,N_3459,N_3410);
xnor U3635 (N_3635,N_3360,N_3238);
or U3636 (N_3636,N_3073,N_3040);
nand U3637 (N_3637,N_3116,N_3213);
nand U3638 (N_3638,N_3260,N_3304);
and U3639 (N_3639,N_3492,N_3412);
or U3640 (N_3640,N_3202,N_3113);
nand U3641 (N_3641,N_3429,N_3207);
nor U3642 (N_3642,N_3389,N_3127);
nor U3643 (N_3643,N_3295,N_3291);
and U3644 (N_3644,N_3257,N_3307);
nand U3645 (N_3645,N_3193,N_3055);
nand U3646 (N_3646,N_3438,N_3333);
or U3647 (N_3647,N_3183,N_3395);
nand U3648 (N_3648,N_3060,N_3141);
nand U3649 (N_3649,N_3171,N_3328);
and U3650 (N_3650,N_3065,N_3204);
nor U3651 (N_3651,N_3430,N_3254);
nor U3652 (N_3652,N_3379,N_3401);
nor U3653 (N_3653,N_3095,N_3124);
nand U3654 (N_3654,N_3220,N_3000);
or U3655 (N_3655,N_3432,N_3247);
nand U3656 (N_3656,N_3158,N_3162);
or U3657 (N_3657,N_3137,N_3159);
xnor U3658 (N_3658,N_3445,N_3205);
nand U3659 (N_3659,N_3050,N_3390);
xnor U3660 (N_3660,N_3198,N_3319);
nor U3661 (N_3661,N_3147,N_3009);
nor U3662 (N_3662,N_3101,N_3436);
nand U3663 (N_3663,N_3201,N_3072);
nand U3664 (N_3664,N_3460,N_3334);
nor U3665 (N_3665,N_3115,N_3034);
nor U3666 (N_3666,N_3263,N_3143);
or U3667 (N_3667,N_3030,N_3453);
or U3668 (N_3668,N_3031,N_3109);
nand U3669 (N_3669,N_3272,N_3398);
or U3670 (N_3670,N_3450,N_3037);
and U3671 (N_3671,N_3103,N_3185);
nor U3672 (N_3672,N_3409,N_3369);
and U3673 (N_3673,N_3394,N_3189);
or U3674 (N_3674,N_3428,N_3122);
or U3675 (N_3675,N_3123,N_3255);
and U3676 (N_3676,N_3008,N_3176);
nor U3677 (N_3677,N_3244,N_3305);
and U3678 (N_3678,N_3364,N_3271);
nor U3679 (N_3679,N_3465,N_3476);
nor U3680 (N_3680,N_3036,N_3178);
xor U3681 (N_3681,N_3019,N_3039);
or U3682 (N_3682,N_3317,N_3281);
nand U3683 (N_3683,N_3021,N_3148);
nand U3684 (N_3684,N_3413,N_3160);
or U3685 (N_3685,N_3164,N_3273);
nor U3686 (N_3686,N_3133,N_3161);
nand U3687 (N_3687,N_3427,N_3175);
nand U3688 (N_3688,N_3200,N_3219);
nand U3689 (N_3689,N_3208,N_3063);
xnor U3690 (N_3690,N_3480,N_3456);
nand U3691 (N_3691,N_3006,N_3365);
and U3692 (N_3692,N_3499,N_3455);
or U3693 (N_3693,N_3259,N_3382);
nor U3694 (N_3694,N_3313,N_3235);
or U3695 (N_3695,N_3311,N_3287);
and U3696 (N_3696,N_3361,N_3252);
and U3697 (N_3697,N_3426,N_3373);
nor U3698 (N_3698,N_3315,N_3352);
or U3699 (N_3699,N_3149,N_3467);
nand U3700 (N_3700,N_3423,N_3014);
nand U3701 (N_3701,N_3068,N_3237);
or U3702 (N_3702,N_3199,N_3076);
nand U3703 (N_3703,N_3078,N_3318);
and U3704 (N_3704,N_3483,N_3084);
nand U3705 (N_3705,N_3435,N_3330);
nor U3706 (N_3706,N_3016,N_3223);
and U3707 (N_3707,N_3165,N_3168);
or U3708 (N_3708,N_3177,N_3126);
xor U3709 (N_3709,N_3274,N_3388);
or U3710 (N_3710,N_3405,N_3308);
nor U3711 (N_3711,N_3231,N_3087);
or U3712 (N_3712,N_3057,N_3118);
or U3713 (N_3713,N_3399,N_3339);
nor U3714 (N_3714,N_3294,N_3346);
nand U3715 (N_3715,N_3121,N_3487);
and U3716 (N_3716,N_3439,N_3195);
nor U3717 (N_3717,N_3179,N_3226);
and U3718 (N_3718,N_3138,N_3135);
xnor U3719 (N_3719,N_3187,N_3246);
or U3720 (N_3720,N_3163,N_3363);
and U3721 (N_3721,N_3392,N_3407);
xor U3722 (N_3722,N_3098,N_3053);
xor U3723 (N_3723,N_3482,N_3139);
nand U3724 (N_3724,N_3300,N_3111);
nand U3725 (N_3725,N_3062,N_3362);
and U3726 (N_3726,N_3047,N_3083);
and U3727 (N_3727,N_3106,N_3264);
and U3728 (N_3728,N_3371,N_3266);
nor U3729 (N_3729,N_3046,N_3351);
nand U3730 (N_3730,N_3190,N_3051);
nand U3731 (N_3731,N_3332,N_3419);
xor U3732 (N_3732,N_3227,N_3471);
nand U3733 (N_3733,N_3107,N_3342);
nor U3734 (N_3734,N_3211,N_3372);
nor U3735 (N_3735,N_3490,N_3033);
nand U3736 (N_3736,N_3449,N_3075);
xor U3737 (N_3737,N_3134,N_3325);
nand U3738 (N_3738,N_3104,N_3327);
nand U3739 (N_3739,N_3431,N_3347);
and U3740 (N_3740,N_3248,N_3384);
or U3741 (N_3741,N_3335,N_3079);
xor U3742 (N_3742,N_3280,N_3498);
nor U3743 (N_3743,N_3381,N_3119);
and U3744 (N_3744,N_3215,N_3048);
xor U3745 (N_3745,N_3353,N_3452);
nor U3746 (N_3746,N_3027,N_3230);
or U3747 (N_3747,N_3186,N_3251);
xor U3748 (N_3748,N_3097,N_3026);
xnor U3749 (N_3749,N_3277,N_3324);
nand U3750 (N_3750,N_3244,N_3302);
and U3751 (N_3751,N_3164,N_3320);
nor U3752 (N_3752,N_3340,N_3174);
nor U3753 (N_3753,N_3063,N_3433);
or U3754 (N_3754,N_3284,N_3298);
or U3755 (N_3755,N_3125,N_3483);
or U3756 (N_3756,N_3052,N_3196);
xnor U3757 (N_3757,N_3183,N_3196);
or U3758 (N_3758,N_3408,N_3185);
and U3759 (N_3759,N_3287,N_3169);
or U3760 (N_3760,N_3128,N_3452);
nand U3761 (N_3761,N_3206,N_3061);
nor U3762 (N_3762,N_3359,N_3438);
nand U3763 (N_3763,N_3131,N_3372);
and U3764 (N_3764,N_3270,N_3214);
or U3765 (N_3765,N_3277,N_3181);
nand U3766 (N_3766,N_3056,N_3095);
and U3767 (N_3767,N_3056,N_3263);
or U3768 (N_3768,N_3363,N_3130);
or U3769 (N_3769,N_3283,N_3388);
nand U3770 (N_3770,N_3097,N_3041);
nand U3771 (N_3771,N_3156,N_3172);
nand U3772 (N_3772,N_3247,N_3235);
nand U3773 (N_3773,N_3248,N_3196);
or U3774 (N_3774,N_3314,N_3070);
nor U3775 (N_3775,N_3470,N_3278);
or U3776 (N_3776,N_3158,N_3252);
and U3777 (N_3777,N_3388,N_3064);
nand U3778 (N_3778,N_3468,N_3459);
nor U3779 (N_3779,N_3469,N_3410);
nand U3780 (N_3780,N_3228,N_3260);
and U3781 (N_3781,N_3087,N_3436);
or U3782 (N_3782,N_3320,N_3409);
and U3783 (N_3783,N_3463,N_3005);
nor U3784 (N_3784,N_3440,N_3387);
or U3785 (N_3785,N_3361,N_3148);
xor U3786 (N_3786,N_3334,N_3483);
or U3787 (N_3787,N_3076,N_3380);
and U3788 (N_3788,N_3420,N_3132);
nand U3789 (N_3789,N_3031,N_3318);
or U3790 (N_3790,N_3067,N_3134);
nor U3791 (N_3791,N_3430,N_3001);
nand U3792 (N_3792,N_3468,N_3402);
and U3793 (N_3793,N_3288,N_3380);
nand U3794 (N_3794,N_3066,N_3217);
and U3795 (N_3795,N_3476,N_3070);
and U3796 (N_3796,N_3171,N_3460);
or U3797 (N_3797,N_3254,N_3120);
and U3798 (N_3798,N_3261,N_3293);
nor U3799 (N_3799,N_3216,N_3159);
nand U3800 (N_3800,N_3263,N_3309);
nand U3801 (N_3801,N_3425,N_3032);
and U3802 (N_3802,N_3281,N_3166);
and U3803 (N_3803,N_3277,N_3176);
xor U3804 (N_3804,N_3456,N_3258);
and U3805 (N_3805,N_3412,N_3174);
and U3806 (N_3806,N_3431,N_3099);
and U3807 (N_3807,N_3217,N_3198);
or U3808 (N_3808,N_3101,N_3097);
xnor U3809 (N_3809,N_3395,N_3342);
nor U3810 (N_3810,N_3461,N_3205);
nor U3811 (N_3811,N_3265,N_3463);
xnor U3812 (N_3812,N_3008,N_3244);
and U3813 (N_3813,N_3264,N_3144);
xnor U3814 (N_3814,N_3306,N_3039);
or U3815 (N_3815,N_3498,N_3394);
nand U3816 (N_3816,N_3138,N_3037);
and U3817 (N_3817,N_3397,N_3245);
or U3818 (N_3818,N_3031,N_3377);
nand U3819 (N_3819,N_3329,N_3003);
nand U3820 (N_3820,N_3076,N_3373);
nor U3821 (N_3821,N_3261,N_3347);
or U3822 (N_3822,N_3422,N_3227);
and U3823 (N_3823,N_3018,N_3413);
nand U3824 (N_3824,N_3271,N_3201);
or U3825 (N_3825,N_3485,N_3009);
or U3826 (N_3826,N_3190,N_3435);
nand U3827 (N_3827,N_3470,N_3279);
nand U3828 (N_3828,N_3033,N_3416);
xor U3829 (N_3829,N_3435,N_3201);
and U3830 (N_3830,N_3269,N_3479);
nand U3831 (N_3831,N_3346,N_3398);
xnor U3832 (N_3832,N_3138,N_3076);
xor U3833 (N_3833,N_3211,N_3099);
nand U3834 (N_3834,N_3128,N_3226);
or U3835 (N_3835,N_3290,N_3082);
and U3836 (N_3836,N_3248,N_3128);
nand U3837 (N_3837,N_3368,N_3355);
nand U3838 (N_3838,N_3423,N_3387);
xnor U3839 (N_3839,N_3201,N_3122);
nor U3840 (N_3840,N_3394,N_3107);
nand U3841 (N_3841,N_3134,N_3104);
and U3842 (N_3842,N_3454,N_3340);
xor U3843 (N_3843,N_3416,N_3369);
nor U3844 (N_3844,N_3375,N_3158);
nor U3845 (N_3845,N_3225,N_3022);
nor U3846 (N_3846,N_3269,N_3263);
or U3847 (N_3847,N_3302,N_3304);
nand U3848 (N_3848,N_3320,N_3338);
nand U3849 (N_3849,N_3129,N_3480);
or U3850 (N_3850,N_3276,N_3026);
and U3851 (N_3851,N_3414,N_3252);
and U3852 (N_3852,N_3488,N_3303);
and U3853 (N_3853,N_3191,N_3110);
nor U3854 (N_3854,N_3228,N_3249);
nor U3855 (N_3855,N_3476,N_3244);
nor U3856 (N_3856,N_3214,N_3450);
or U3857 (N_3857,N_3398,N_3145);
nand U3858 (N_3858,N_3085,N_3357);
or U3859 (N_3859,N_3192,N_3398);
or U3860 (N_3860,N_3323,N_3436);
nand U3861 (N_3861,N_3035,N_3225);
nor U3862 (N_3862,N_3318,N_3391);
and U3863 (N_3863,N_3089,N_3494);
nor U3864 (N_3864,N_3279,N_3061);
and U3865 (N_3865,N_3263,N_3253);
nand U3866 (N_3866,N_3435,N_3272);
nor U3867 (N_3867,N_3052,N_3257);
xnor U3868 (N_3868,N_3382,N_3291);
or U3869 (N_3869,N_3474,N_3099);
and U3870 (N_3870,N_3313,N_3426);
nor U3871 (N_3871,N_3071,N_3013);
nand U3872 (N_3872,N_3404,N_3214);
nand U3873 (N_3873,N_3095,N_3182);
and U3874 (N_3874,N_3191,N_3362);
xor U3875 (N_3875,N_3499,N_3467);
or U3876 (N_3876,N_3150,N_3292);
nand U3877 (N_3877,N_3428,N_3228);
nand U3878 (N_3878,N_3305,N_3151);
and U3879 (N_3879,N_3390,N_3090);
or U3880 (N_3880,N_3379,N_3454);
xor U3881 (N_3881,N_3436,N_3153);
or U3882 (N_3882,N_3108,N_3438);
nor U3883 (N_3883,N_3196,N_3108);
and U3884 (N_3884,N_3210,N_3389);
or U3885 (N_3885,N_3499,N_3223);
and U3886 (N_3886,N_3324,N_3321);
and U3887 (N_3887,N_3017,N_3416);
nand U3888 (N_3888,N_3412,N_3384);
and U3889 (N_3889,N_3026,N_3169);
or U3890 (N_3890,N_3205,N_3000);
nor U3891 (N_3891,N_3444,N_3090);
nand U3892 (N_3892,N_3464,N_3179);
xnor U3893 (N_3893,N_3425,N_3048);
or U3894 (N_3894,N_3006,N_3044);
nand U3895 (N_3895,N_3101,N_3455);
nand U3896 (N_3896,N_3099,N_3224);
nor U3897 (N_3897,N_3110,N_3315);
or U3898 (N_3898,N_3208,N_3007);
nand U3899 (N_3899,N_3006,N_3294);
and U3900 (N_3900,N_3474,N_3294);
xor U3901 (N_3901,N_3359,N_3180);
nor U3902 (N_3902,N_3368,N_3434);
xor U3903 (N_3903,N_3196,N_3227);
and U3904 (N_3904,N_3444,N_3227);
xor U3905 (N_3905,N_3490,N_3424);
nor U3906 (N_3906,N_3337,N_3472);
or U3907 (N_3907,N_3162,N_3088);
and U3908 (N_3908,N_3266,N_3468);
xor U3909 (N_3909,N_3129,N_3067);
nor U3910 (N_3910,N_3418,N_3132);
nor U3911 (N_3911,N_3137,N_3383);
nor U3912 (N_3912,N_3041,N_3248);
and U3913 (N_3913,N_3025,N_3299);
or U3914 (N_3914,N_3238,N_3044);
or U3915 (N_3915,N_3213,N_3030);
nor U3916 (N_3916,N_3258,N_3485);
nor U3917 (N_3917,N_3059,N_3306);
nand U3918 (N_3918,N_3453,N_3425);
nor U3919 (N_3919,N_3150,N_3289);
nor U3920 (N_3920,N_3114,N_3136);
nor U3921 (N_3921,N_3140,N_3448);
or U3922 (N_3922,N_3046,N_3350);
and U3923 (N_3923,N_3279,N_3476);
or U3924 (N_3924,N_3220,N_3378);
and U3925 (N_3925,N_3061,N_3264);
and U3926 (N_3926,N_3107,N_3194);
or U3927 (N_3927,N_3437,N_3014);
nand U3928 (N_3928,N_3274,N_3072);
xnor U3929 (N_3929,N_3073,N_3463);
nand U3930 (N_3930,N_3219,N_3110);
nand U3931 (N_3931,N_3061,N_3157);
or U3932 (N_3932,N_3351,N_3405);
nor U3933 (N_3933,N_3158,N_3408);
and U3934 (N_3934,N_3151,N_3334);
nor U3935 (N_3935,N_3040,N_3096);
or U3936 (N_3936,N_3340,N_3279);
nor U3937 (N_3937,N_3092,N_3195);
nor U3938 (N_3938,N_3403,N_3011);
nand U3939 (N_3939,N_3454,N_3347);
nor U3940 (N_3940,N_3364,N_3423);
nand U3941 (N_3941,N_3108,N_3375);
nor U3942 (N_3942,N_3489,N_3452);
or U3943 (N_3943,N_3483,N_3385);
nor U3944 (N_3944,N_3441,N_3342);
and U3945 (N_3945,N_3226,N_3260);
or U3946 (N_3946,N_3296,N_3185);
and U3947 (N_3947,N_3001,N_3225);
nor U3948 (N_3948,N_3323,N_3154);
nor U3949 (N_3949,N_3438,N_3320);
and U3950 (N_3950,N_3349,N_3359);
and U3951 (N_3951,N_3257,N_3402);
nor U3952 (N_3952,N_3389,N_3068);
and U3953 (N_3953,N_3302,N_3342);
nor U3954 (N_3954,N_3107,N_3106);
and U3955 (N_3955,N_3123,N_3118);
nor U3956 (N_3956,N_3313,N_3043);
nand U3957 (N_3957,N_3193,N_3115);
and U3958 (N_3958,N_3441,N_3181);
or U3959 (N_3959,N_3476,N_3354);
xor U3960 (N_3960,N_3194,N_3144);
nand U3961 (N_3961,N_3471,N_3075);
or U3962 (N_3962,N_3199,N_3145);
or U3963 (N_3963,N_3141,N_3398);
xor U3964 (N_3964,N_3389,N_3106);
nand U3965 (N_3965,N_3333,N_3008);
nor U3966 (N_3966,N_3278,N_3035);
nand U3967 (N_3967,N_3341,N_3285);
and U3968 (N_3968,N_3066,N_3268);
nand U3969 (N_3969,N_3130,N_3365);
and U3970 (N_3970,N_3008,N_3374);
or U3971 (N_3971,N_3268,N_3241);
nor U3972 (N_3972,N_3342,N_3414);
nand U3973 (N_3973,N_3248,N_3336);
nor U3974 (N_3974,N_3480,N_3205);
nor U3975 (N_3975,N_3479,N_3218);
and U3976 (N_3976,N_3069,N_3020);
or U3977 (N_3977,N_3447,N_3426);
and U3978 (N_3978,N_3360,N_3252);
and U3979 (N_3979,N_3188,N_3283);
or U3980 (N_3980,N_3261,N_3321);
nand U3981 (N_3981,N_3187,N_3126);
nor U3982 (N_3982,N_3416,N_3367);
nor U3983 (N_3983,N_3467,N_3351);
nand U3984 (N_3984,N_3162,N_3023);
nand U3985 (N_3985,N_3288,N_3407);
nor U3986 (N_3986,N_3341,N_3247);
and U3987 (N_3987,N_3022,N_3270);
and U3988 (N_3988,N_3312,N_3326);
nand U3989 (N_3989,N_3398,N_3222);
xor U3990 (N_3990,N_3012,N_3297);
and U3991 (N_3991,N_3489,N_3299);
nand U3992 (N_3992,N_3289,N_3420);
or U3993 (N_3993,N_3345,N_3281);
nor U3994 (N_3994,N_3388,N_3403);
nor U3995 (N_3995,N_3010,N_3401);
nor U3996 (N_3996,N_3473,N_3437);
xor U3997 (N_3997,N_3026,N_3168);
nor U3998 (N_3998,N_3340,N_3096);
and U3999 (N_3999,N_3421,N_3039);
xor U4000 (N_4000,N_3523,N_3644);
xor U4001 (N_4001,N_3935,N_3954);
or U4002 (N_4002,N_3869,N_3512);
and U4003 (N_4003,N_3896,N_3544);
xor U4004 (N_4004,N_3876,N_3841);
and U4005 (N_4005,N_3934,N_3984);
nor U4006 (N_4006,N_3820,N_3967);
and U4007 (N_4007,N_3905,N_3835);
xnor U4008 (N_4008,N_3939,N_3847);
and U4009 (N_4009,N_3626,N_3949);
nor U4010 (N_4010,N_3510,N_3638);
nand U4011 (N_4011,N_3814,N_3628);
nand U4012 (N_4012,N_3543,N_3972);
nor U4013 (N_4013,N_3586,N_3658);
nand U4014 (N_4014,N_3988,N_3800);
or U4015 (N_4015,N_3824,N_3948);
or U4016 (N_4016,N_3643,N_3887);
and U4017 (N_4017,N_3808,N_3529);
or U4018 (N_4018,N_3855,N_3928);
nand U4019 (N_4019,N_3581,N_3969);
xor U4020 (N_4020,N_3840,N_3873);
and U4021 (N_4021,N_3675,N_3990);
or U4022 (N_4022,N_3993,N_3868);
and U4023 (N_4023,N_3827,N_3974);
nor U4024 (N_4024,N_3627,N_3513);
and U4025 (N_4025,N_3966,N_3561);
or U4026 (N_4026,N_3670,N_3812);
xnor U4027 (N_4027,N_3556,N_3728);
nor U4028 (N_4028,N_3721,N_3906);
or U4029 (N_4029,N_3530,N_3573);
nand U4030 (N_4030,N_3958,N_3851);
and U4031 (N_4031,N_3802,N_3551);
xnor U4032 (N_4032,N_3878,N_3514);
nor U4033 (N_4033,N_3631,N_3539);
and U4034 (N_4034,N_3674,N_3596);
or U4035 (N_4035,N_3546,N_3953);
and U4036 (N_4036,N_3532,N_3985);
nand U4037 (N_4037,N_3863,N_3616);
xor U4038 (N_4038,N_3772,N_3785);
nor U4039 (N_4039,N_3766,N_3642);
and U4040 (N_4040,N_3667,N_3611);
nand U4041 (N_4041,N_3600,N_3940);
nor U4042 (N_4042,N_3655,N_3646);
nor U4043 (N_4043,N_3649,N_3701);
or U4044 (N_4044,N_3923,N_3787);
nand U4045 (N_4045,N_3957,N_3996);
and U4046 (N_4046,N_3740,N_3941);
or U4047 (N_4047,N_3621,N_3994);
nor U4048 (N_4048,N_3811,N_3942);
or U4049 (N_4049,N_3592,N_3682);
or U4050 (N_4050,N_3566,N_3977);
nor U4051 (N_4051,N_3915,N_3843);
or U4052 (N_4052,N_3760,N_3577);
nor U4053 (N_4053,N_3755,N_3515);
and U4054 (N_4054,N_3562,N_3689);
xnor U4055 (N_4055,N_3589,N_3833);
nand U4056 (N_4056,N_3860,N_3872);
and U4057 (N_4057,N_3837,N_3792);
xnor U4058 (N_4058,N_3893,N_3735);
xor U4059 (N_4059,N_3538,N_3799);
or U4060 (N_4060,N_3697,N_3859);
nor U4061 (N_4061,N_3681,N_3956);
nor U4062 (N_4062,N_3997,N_3550);
or U4063 (N_4063,N_3509,N_3503);
nor U4064 (N_4064,N_3895,N_3920);
nor U4065 (N_4065,N_3610,N_3575);
and U4066 (N_4066,N_3962,N_3633);
and U4067 (N_4067,N_3933,N_3846);
or U4068 (N_4068,N_3622,N_3796);
nand U4069 (N_4069,N_3866,N_3756);
nor U4070 (N_4070,N_3517,N_3725);
nor U4071 (N_4071,N_3639,N_3629);
and U4072 (N_4072,N_3914,N_3640);
and U4073 (N_4073,N_3845,N_3788);
or U4074 (N_4074,N_3867,N_3922);
or U4075 (N_4075,N_3804,N_3572);
and U4076 (N_4076,N_3998,N_3630);
and U4077 (N_4077,N_3729,N_3927);
and U4078 (N_4078,N_3542,N_3854);
and U4079 (N_4079,N_3753,N_3778);
and U4080 (N_4080,N_3931,N_3618);
or U4081 (N_4081,N_3983,N_3715);
nor U4082 (N_4082,N_3909,N_3856);
nor U4083 (N_4083,N_3656,N_3738);
and U4084 (N_4084,N_3825,N_3897);
nor U4085 (N_4085,N_3890,N_3797);
nor U4086 (N_4086,N_3961,N_3813);
xor U4087 (N_4087,N_3696,N_3694);
or U4088 (N_4088,N_3617,N_3992);
or U4089 (N_4089,N_3698,N_3625);
xor U4090 (N_4090,N_3786,N_3613);
or U4091 (N_4091,N_3522,N_3917);
and U4092 (N_4092,N_3870,N_3724);
nor U4093 (N_4093,N_3536,N_3659);
or U4094 (N_4094,N_3826,N_3925);
or U4095 (N_4095,N_3816,N_3502);
or U4096 (N_4096,N_3557,N_3937);
nand U4097 (N_4097,N_3565,N_3938);
xor U4098 (N_4098,N_3865,N_3676);
nor U4099 (N_4099,N_3615,N_3518);
and U4100 (N_4100,N_3757,N_3593);
and U4101 (N_4101,N_3970,N_3834);
and U4102 (N_4102,N_3641,N_3590);
or U4103 (N_4103,N_3947,N_3660);
nand U4104 (N_4104,N_3844,N_3853);
or U4105 (N_4105,N_3582,N_3603);
or U4106 (N_4106,N_3708,N_3780);
and U4107 (N_4107,N_3535,N_3741);
and U4108 (N_4108,N_3946,N_3723);
nand U4109 (N_4109,N_3665,N_3894);
nor U4110 (N_4110,N_3885,N_3680);
or U4111 (N_4111,N_3547,N_3730);
and U4112 (N_4112,N_3995,N_3910);
xnor U4113 (N_4113,N_3533,N_3761);
and U4114 (N_4114,N_3850,N_3700);
or U4115 (N_4115,N_3763,N_3736);
nand U4116 (N_4116,N_3886,N_3806);
or U4117 (N_4117,N_3637,N_3776);
or U4118 (N_4118,N_3548,N_3880);
or U4119 (N_4119,N_3884,N_3688);
nor U4120 (N_4120,N_3570,N_3768);
and U4121 (N_4121,N_3727,N_3559);
nor U4122 (N_4122,N_3511,N_3580);
nand U4123 (N_4123,N_3764,N_3705);
nand U4124 (N_4124,N_3653,N_3801);
nand U4125 (N_4125,N_3554,N_3798);
or U4126 (N_4126,N_3569,N_3810);
or U4127 (N_4127,N_3578,N_3881);
or U4128 (N_4128,N_3982,N_3500);
or U4129 (N_4129,N_3683,N_3750);
nand U4130 (N_4130,N_3703,N_3684);
nor U4131 (N_4131,N_3709,N_3823);
or U4132 (N_4132,N_3747,N_3545);
nor U4133 (N_4133,N_3980,N_3504);
xor U4134 (N_4134,N_3775,N_3534);
nand U4135 (N_4135,N_3508,N_3516);
and U4136 (N_4136,N_3902,N_3930);
or U4137 (N_4137,N_3889,N_3558);
nor U4138 (N_4138,N_3832,N_3913);
nand U4139 (N_4139,N_3563,N_3612);
and U4140 (N_4140,N_3849,N_3744);
nand U4141 (N_4141,N_3652,N_3521);
xnor U4142 (N_4142,N_3525,N_3691);
xnor U4143 (N_4143,N_3790,N_3916);
nand U4144 (N_4144,N_3695,N_3891);
or U4145 (N_4145,N_3829,N_3791);
nor U4146 (N_4146,N_3609,N_3842);
nor U4147 (N_4147,N_3921,N_3720);
and U4148 (N_4148,N_3541,N_3782);
nand U4149 (N_4149,N_3686,N_3944);
nand U4150 (N_4150,N_3879,N_3672);
nor U4151 (N_4151,N_3943,N_3882);
and U4152 (N_4152,N_3751,N_3762);
or U4153 (N_4153,N_3874,N_3583);
nand U4154 (N_4154,N_3506,N_3978);
or U4155 (N_4155,N_3588,N_3901);
nand U4156 (N_4156,N_3828,N_3531);
or U4157 (N_4157,N_3819,N_3809);
nor U4158 (N_4158,N_3770,N_3524);
xnor U4159 (N_4159,N_3731,N_3699);
xnor U4160 (N_4160,N_3662,N_3945);
and U4161 (N_4161,N_3929,N_3779);
nor U4162 (N_4162,N_3784,N_3737);
nor U4163 (N_4163,N_3754,N_3888);
nand U4164 (N_4164,N_3900,N_3955);
nand U4165 (N_4165,N_3991,N_3601);
xor U4166 (N_4166,N_3803,N_3607);
or U4167 (N_4167,N_3950,N_3677);
nor U4168 (N_4168,N_3794,N_3789);
nor U4169 (N_4169,N_3857,N_3599);
and U4170 (N_4170,N_3769,N_3707);
or U4171 (N_4171,N_3719,N_3574);
nand U4172 (N_4172,N_3952,N_3702);
xor U4173 (N_4173,N_3687,N_3604);
or U4174 (N_4174,N_3734,N_3919);
nor U4175 (N_4175,N_3759,N_3752);
nand U4176 (N_4176,N_3654,N_3528);
nor U4177 (N_4177,N_3777,N_3714);
nand U4178 (N_4178,N_3908,N_3598);
or U4179 (N_4179,N_3911,N_3624);
or U4180 (N_4180,N_3567,N_3620);
xnor U4181 (N_4181,N_3903,N_3979);
xor U4182 (N_4182,N_3527,N_3713);
xor U4183 (N_4183,N_3669,N_3739);
nand U4184 (N_4184,N_3822,N_3717);
and U4185 (N_4185,N_3960,N_3963);
or U4186 (N_4186,N_3671,N_3585);
nor U4187 (N_4187,N_3838,N_3711);
or U4188 (N_4188,N_3564,N_3732);
or U4189 (N_4189,N_3975,N_3795);
nor U4190 (N_4190,N_3807,N_3999);
nand U4191 (N_4191,N_3666,N_3733);
xor U4192 (N_4192,N_3924,N_3726);
or U4193 (N_4193,N_3595,N_3718);
xor U4194 (N_4194,N_3877,N_3986);
and U4195 (N_4195,N_3875,N_3597);
and U4196 (N_4196,N_3571,N_3679);
and U4197 (N_4197,N_3553,N_3634);
nand U4198 (N_4198,N_3805,N_3836);
and U4199 (N_4199,N_3605,N_3712);
and U4200 (N_4200,N_3647,N_3650);
nor U4201 (N_4201,N_3651,N_3526);
and U4202 (N_4202,N_3552,N_3918);
nand U4203 (N_4203,N_3758,N_3663);
xnor U4204 (N_4204,N_3668,N_3987);
nor U4205 (N_4205,N_3959,N_3507);
nor U4206 (N_4206,N_3830,N_3587);
nand U4207 (N_4207,N_3576,N_3594);
or U4208 (N_4208,N_3746,N_3549);
and U4209 (N_4209,N_3965,N_3560);
nand U4210 (N_4210,N_3716,N_3602);
xnor U4211 (N_4211,N_3648,N_3861);
nor U4212 (N_4212,N_3774,N_3971);
nor U4213 (N_4213,N_3608,N_3821);
or U4214 (N_4214,N_3765,N_3661);
nor U4215 (N_4215,N_3781,N_3520);
or U4216 (N_4216,N_3907,N_3704);
or U4217 (N_4217,N_3818,N_3926);
or U4218 (N_4218,N_3817,N_3748);
and U4219 (N_4219,N_3951,N_3614);
or U4220 (N_4220,N_3690,N_3981);
nand U4221 (N_4221,N_3831,N_3606);
nor U4222 (N_4222,N_3793,N_3767);
nor U4223 (N_4223,N_3505,N_3657);
nor U4224 (N_4224,N_3976,N_3636);
nor U4225 (N_4225,N_3501,N_3664);
or U4226 (N_4226,N_3745,N_3852);
and U4227 (N_4227,N_3749,N_3871);
or U4228 (N_4228,N_3742,N_3904);
or U4229 (N_4229,N_3864,N_3519);
nor U4230 (N_4230,N_3862,N_3623);
nor U4231 (N_4231,N_3912,N_3899);
nand U4232 (N_4232,N_3898,N_3773);
nand U4233 (N_4233,N_3685,N_3692);
xor U4234 (N_4234,N_3678,N_3632);
and U4235 (N_4235,N_3568,N_3848);
or U4236 (N_4236,N_3839,N_3537);
xor U4237 (N_4237,N_3635,N_3883);
xnor U4238 (N_4238,N_3710,N_3673);
and U4239 (N_4239,N_3968,N_3743);
and U4240 (N_4240,N_3858,N_3932);
nor U4241 (N_4241,N_3619,N_3973);
nor U4242 (N_4242,N_3579,N_3693);
nor U4243 (N_4243,N_3892,N_3783);
nand U4244 (N_4244,N_3645,N_3964);
nor U4245 (N_4245,N_3936,N_3540);
or U4246 (N_4246,N_3584,N_3706);
nand U4247 (N_4247,N_3989,N_3771);
nor U4248 (N_4248,N_3722,N_3815);
and U4249 (N_4249,N_3591,N_3555);
nor U4250 (N_4250,N_3769,N_3886);
nand U4251 (N_4251,N_3649,N_3994);
nand U4252 (N_4252,N_3897,N_3770);
nand U4253 (N_4253,N_3587,N_3688);
nor U4254 (N_4254,N_3687,N_3933);
and U4255 (N_4255,N_3608,N_3575);
or U4256 (N_4256,N_3562,N_3505);
nor U4257 (N_4257,N_3618,N_3844);
or U4258 (N_4258,N_3926,N_3542);
and U4259 (N_4259,N_3533,N_3675);
nand U4260 (N_4260,N_3558,N_3685);
xor U4261 (N_4261,N_3642,N_3783);
nor U4262 (N_4262,N_3741,N_3711);
and U4263 (N_4263,N_3710,N_3590);
and U4264 (N_4264,N_3725,N_3562);
or U4265 (N_4265,N_3891,N_3688);
nor U4266 (N_4266,N_3628,N_3663);
or U4267 (N_4267,N_3686,N_3704);
nor U4268 (N_4268,N_3524,N_3638);
nand U4269 (N_4269,N_3885,N_3922);
xnor U4270 (N_4270,N_3661,N_3693);
and U4271 (N_4271,N_3962,N_3814);
or U4272 (N_4272,N_3838,N_3808);
or U4273 (N_4273,N_3657,N_3739);
nand U4274 (N_4274,N_3587,N_3753);
or U4275 (N_4275,N_3792,N_3588);
or U4276 (N_4276,N_3616,N_3875);
or U4277 (N_4277,N_3902,N_3671);
nor U4278 (N_4278,N_3952,N_3877);
nand U4279 (N_4279,N_3656,N_3975);
nand U4280 (N_4280,N_3946,N_3638);
or U4281 (N_4281,N_3808,N_3687);
or U4282 (N_4282,N_3764,N_3796);
or U4283 (N_4283,N_3723,N_3820);
and U4284 (N_4284,N_3878,N_3744);
and U4285 (N_4285,N_3524,N_3602);
or U4286 (N_4286,N_3878,N_3812);
xnor U4287 (N_4287,N_3678,N_3574);
nor U4288 (N_4288,N_3773,N_3737);
or U4289 (N_4289,N_3625,N_3772);
nand U4290 (N_4290,N_3918,N_3791);
nand U4291 (N_4291,N_3559,N_3924);
and U4292 (N_4292,N_3799,N_3775);
nor U4293 (N_4293,N_3806,N_3881);
or U4294 (N_4294,N_3698,N_3578);
or U4295 (N_4295,N_3676,N_3962);
nand U4296 (N_4296,N_3959,N_3699);
or U4297 (N_4297,N_3720,N_3662);
or U4298 (N_4298,N_3749,N_3989);
nand U4299 (N_4299,N_3720,N_3693);
nor U4300 (N_4300,N_3577,N_3940);
or U4301 (N_4301,N_3973,N_3637);
or U4302 (N_4302,N_3582,N_3899);
nand U4303 (N_4303,N_3629,N_3884);
nor U4304 (N_4304,N_3765,N_3815);
xor U4305 (N_4305,N_3570,N_3644);
or U4306 (N_4306,N_3765,N_3628);
and U4307 (N_4307,N_3745,N_3697);
xnor U4308 (N_4308,N_3792,N_3629);
or U4309 (N_4309,N_3629,N_3645);
nor U4310 (N_4310,N_3663,N_3762);
xor U4311 (N_4311,N_3834,N_3756);
and U4312 (N_4312,N_3984,N_3734);
xnor U4313 (N_4313,N_3714,N_3643);
or U4314 (N_4314,N_3544,N_3713);
nor U4315 (N_4315,N_3604,N_3764);
or U4316 (N_4316,N_3885,N_3517);
nor U4317 (N_4317,N_3786,N_3690);
or U4318 (N_4318,N_3960,N_3771);
nand U4319 (N_4319,N_3612,N_3764);
or U4320 (N_4320,N_3843,N_3571);
and U4321 (N_4321,N_3935,N_3593);
and U4322 (N_4322,N_3891,N_3843);
or U4323 (N_4323,N_3827,N_3676);
and U4324 (N_4324,N_3716,N_3916);
nor U4325 (N_4325,N_3740,N_3990);
nand U4326 (N_4326,N_3810,N_3842);
or U4327 (N_4327,N_3873,N_3948);
nand U4328 (N_4328,N_3787,N_3559);
nor U4329 (N_4329,N_3966,N_3902);
and U4330 (N_4330,N_3978,N_3755);
or U4331 (N_4331,N_3899,N_3539);
or U4332 (N_4332,N_3948,N_3649);
and U4333 (N_4333,N_3843,N_3663);
nand U4334 (N_4334,N_3767,N_3867);
or U4335 (N_4335,N_3692,N_3812);
nor U4336 (N_4336,N_3848,N_3684);
nor U4337 (N_4337,N_3653,N_3513);
and U4338 (N_4338,N_3719,N_3910);
or U4339 (N_4339,N_3653,N_3892);
or U4340 (N_4340,N_3935,N_3878);
and U4341 (N_4341,N_3515,N_3639);
or U4342 (N_4342,N_3623,N_3827);
nor U4343 (N_4343,N_3709,N_3597);
and U4344 (N_4344,N_3615,N_3735);
or U4345 (N_4345,N_3824,N_3651);
and U4346 (N_4346,N_3639,N_3844);
nand U4347 (N_4347,N_3797,N_3893);
and U4348 (N_4348,N_3714,N_3901);
nor U4349 (N_4349,N_3995,N_3979);
nor U4350 (N_4350,N_3614,N_3917);
or U4351 (N_4351,N_3616,N_3695);
nor U4352 (N_4352,N_3611,N_3985);
nand U4353 (N_4353,N_3559,N_3780);
nand U4354 (N_4354,N_3808,N_3724);
and U4355 (N_4355,N_3962,N_3598);
nand U4356 (N_4356,N_3922,N_3587);
and U4357 (N_4357,N_3837,N_3684);
nor U4358 (N_4358,N_3799,N_3578);
nor U4359 (N_4359,N_3903,N_3780);
nor U4360 (N_4360,N_3816,N_3641);
or U4361 (N_4361,N_3611,N_3626);
xor U4362 (N_4362,N_3617,N_3941);
nand U4363 (N_4363,N_3834,N_3767);
nor U4364 (N_4364,N_3537,N_3652);
or U4365 (N_4365,N_3786,N_3919);
and U4366 (N_4366,N_3870,N_3951);
or U4367 (N_4367,N_3790,N_3651);
nor U4368 (N_4368,N_3988,N_3612);
and U4369 (N_4369,N_3571,N_3855);
nand U4370 (N_4370,N_3909,N_3810);
nor U4371 (N_4371,N_3527,N_3814);
and U4372 (N_4372,N_3730,N_3508);
nand U4373 (N_4373,N_3602,N_3571);
nor U4374 (N_4374,N_3881,N_3956);
nor U4375 (N_4375,N_3824,N_3806);
and U4376 (N_4376,N_3614,N_3797);
xnor U4377 (N_4377,N_3837,N_3804);
and U4378 (N_4378,N_3507,N_3680);
and U4379 (N_4379,N_3541,N_3616);
nor U4380 (N_4380,N_3818,N_3650);
or U4381 (N_4381,N_3824,N_3905);
and U4382 (N_4382,N_3567,N_3922);
and U4383 (N_4383,N_3671,N_3600);
nor U4384 (N_4384,N_3779,N_3978);
nand U4385 (N_4385,N_3850,N_3797);
and U4386 (N_4386,N_3748,N_3979);
nor U4387 (N_4387,N_3691,N_3915);
nand U4388 (N_4388,N_3526,N_3686);
and U4389 (N_4389,N_3964,N_3717);
and U4390 (N_4390,N_3542,N_3541);
xnor U4391 (N_4391,N_3564,N_3627);
or U4392 (N_4392,N_3685,N_3704);
nor U4393 (N_4393,N_3778,N_3997);
nand U4394 (N_4394,N_3658,N_3508);
and U4395 (N_4395,N_3814,N_3815);
and U4396 (N_4396,N_3679,N_3557);
nand U4397 (N_4397,N_3580,N_3932);
and U4398 (N_4398,N_3546,N_3628);
nor U4399 (N_4399,N_3859,N_3753);
and U4400 (N_4400,N_3501,N_3899);
nor U4401 (N_4401,N_3922,N_3651);
or U4402 (N_4402,N_3919,N_3907);
or U4403 (N_4403,N_3538,N_3573);
nand U4404 (N_4404,N_3926,N_3563);
nand U4405 (N_4405,N_3701,N_3922);
nand U4406 (N_4406,N_3581,N_3832);
or U4407 (N_4407,N_3697,N_3989);
nand U4408 (N_4408,N_3620,N_3876);
nor U4409 (N_4409,N_3911,N_3719);
or U4410 (N_4410,N_3532,N_3838);
nand U4411 (N_4411,N_3803,N_3954);
or U4412 (N_4412,N_3823,N_3960);
nor U4413 (N_4413,N_3669,N_3579);
nor U4414 (N_4414,N_3833,N_3585);
nand U4415 (N_4415,N_3730,N_3620);
nor U4416 (N_4416,N_3724,N_3922);
nor U4417 (N_4417,N_3533,N_3907);
nand U4418 (N_4418,N_3983,N_3718);
or U4419 (N_4419,N_3937,N_3901);
or U4420 (N_4420,N_3951,N_3603);
or U4421 (N_4421,N_3510,N_3901);
nand U4422 (N_4422,N_3575,N_3727);
and U4423 (N_4423,N_3560,N_3659);
xor U4424 (N_4424,N_3625,N_3786);
nor U4425 (N_4425,N_3978,N_3600);
nand U4426 (N_4426,N_3617,N_3838);
nand U4427 (N_4427,N_3703,N_3664);
and U4428 (N_4428,N_3797,N_3927);
and U4429 (N_4429,N_3993,N_3856);
and U4430 (N_4430,N_3558,N_3887);
and U4431 (N_4431,N_3502,N_3937);
xnor U4432 (N_4432,N_3752,N_3900);
nor U4433 (N_4433,N_3762,N_3562);
or U4434 (N_4434,N_3708,N_3949);
nand U4435 (N_4435,N_3811,N_3798);
or U4436 (N_4436,N_3732,N_3913);
xnor U4437 (N_4437,N_3681,N_3657);
or U4438 (N_4438,N_3698,N_3580);
nor U4439 (N_4439,N_3596,N_3743);
and U4440 (N_4440,N_3513,N_3943);
nor U4441 (N_4441,N_3589,N_3723);
nand U4442 (N_4442,N_3566,N_3507);
or U4443 (N_4443,N_3775,N_3725);
xor U4444 (N_4444,N_3831,N_3820);
nor U4445 (N_4445,N_3678,N_3989);
or U4446 (N_4446,N_3550,N_3946);
nand U4447 (N_4447,N_3517,N_3970);
nor U4448 (N_4448,N_3925,N_3969);
and U4449 (N_4449,N_3624,N_3811);
nand U4450 (N_4450,N_3631,N_3787);
and U4451 (N_4451,N_3596,N_3943);
or U4452 (N_4452,N_3764,N_3728);
nor U4453 (N_4453,N_3897,N_3647);
nand U4454 (N_4454,N_3581,N_3799);
nand U4455 (N_4455,N_3955,N_3841);
or U4456 (N_4456,N_3954,N_3952);
nor U4457 (N_4457,N_3615,N_3982);
and U4458 (N_4458,N_3837,N_3784);
nor U4459 (N_4459,N_3762,N_3799);
nor U4460 (N_4460,N_3913,N_3882);
nor U4461 (N_4461,N_3715,N_3779);
and U4462 (N_4462,N_3877,N_3585);
or U4463 (N_4463,N_3774,N_3667);
nand U4464 (N_4464,N_3556,N_3834);
nand U4465 (N_4465,N_3848,N_3596);
xor U4466 (N_4466,N_3873,N_3926);
nor U4467 (N_4467,N_3930,N_3608);
or U4468 (N_4468,N_3606,N_3894);
nor U4469 (N_4469,N_3754,N_3835);
nor U4470 (N_4470,N_3955,N_3611);
xnor U4471 (N_4471,N_3844,N_3536);
nand U4472 (N_4472,N_3893,N_3647);
and U4473 (N_4473,N_3940,N_3588);
nand U4474 (N_4474,N_3633,N_3830);
nand U4475 (N_4475,N_3831,N_3674);
and U4476 (N_4476,N_3803,N_3983);
and U4477 (N_4477,N_3973,N_3542);
or U4478 (N_4478,N_3833,N_3651);
nor U4479 (N_4479,N_3788,N_3575);
or U4480 (N_4480,N_3894,N_3924);
and U4481 (N_4481,N_3543,N_3634);
and U4482 (N_4482,N_3912,N_3578);
and U4483 (N_4483,N_3859,N_3763);
or U4484 (N_4484,N_3932,N_3965);
xor U4485 (N_4485,N_3744,N_3644);
or U4486 (N_4486,N_3976,N_3926);
and U4487 (N_4487,N_3500,N_3881);
nor U4488 (N_4488,N_3867,N_3693);
xnor U4489 (N_4489,N_3625,N_3791);
or U4490 (N_4490,N_3746,N_3608);
and U4491 (N_4491,N_3758,N_3500);
nor U4492 (N_4492,N_3678,N_3817);
nand U4493 (N_4493,N_3905,N_3787);
and U4494 (N_4494,N_3521,N_3769);
nand U4495 (N_4495,N_3637,N_3981);
or U4496 (N_4496,N_3728,N_3703);
or U4497 (N_4497,N_3832,N_3988);
and U4498 (N_4498,N_3937,N_3737);
nor U4499 (N_4499,N_3620,N_3776);
nor U4500 (N_4500,N_4418,N_4312);
xor U4501 (N_4501,N_4081,N_4212);
or U4502 (N_4502,N_4356,N_4468);
and U4503 (N_4503,N_4173,N_4238);
nand U4504 (N_4504,N_4384,N_4264);
nand U4505 (N_4505,N_4337,N_4358);
or U4506 (N_4506,N_4300,N_4276);
nor U4507 (N_4507,N_4410,N_4028);
and U4508 (N_4508,N_4096,N_4421);
or U4509 (N_4509,N_4495,N_4326);
or U4510 (N_4510,N_4402,N_4139);
and U4511 (N_4511,N_4279,N_4443);
or U4512 (N_4512,N_4253,N_4455);
nor U4513 (N_4513,N_4259,N_4146);
nand U4514 (N_4514,N_4088,N_4460);
or U4515 (N_4515,N_4446,N_4226);
nand U4516 (N_4516,N_4031,N_4019);
xnor U4517 (N_4517,N_4108,N_4383);
nor U4518 (N_4518,N_4044,N_4271);
or U4519 (N_4519,N_4313,N_4491);
nand U4520 (N_4520,N_4397,N_4024);
xnor U4521 (N_4521,N_4317,N_4377);
and U4522 (N_4522,N_4154,N_4355);
nor U4523 (N_4523,N_4296,N_4207);
nand U4524 (N_4524,N_4021,N_4042);
nor U4525 (N_4525,N_4182,N_4122);
and U4526 (N_4526,N_4060,N_4396);
or U4527 (N_4527,N_4181,N_4140);
nand U4528 (N_4528,N_4408,N_4353);
and U4529 (N_4529,N_4391,N_4417);
or U4530 (N_4530,N_4399,N_4006);
or U4531 (N_4531,N_4252,N_4255);
nor U4532 (N_4532,N_4117,N_4000);
nand U4533 (N_4533,N_4304,N_4363);
nand U4534 (N_4534,N_4265,N_4289);
and U4535 (N_4535,N_4111,N_4013);
nand U4536 (N_4536,N_4215,N_4053);
and U4537 (N_4537,N_4071,N_4423);
and U4538 (N_4538,N_4229,N_4109);
nor U4539 (N_4539,N_4392,N_4321);
nor U4540 (N_4540,N_4038,N_4022);
and U4541 (N_4541,N_4406,N_4453);
nand U4542 (N_4542,N_4436,N_4197);
nor U4543 (N_4543,N_4156,N_4112);
nand U4544 (N_4544,N_4341,N_4496);
nor U4545 (N_4545,N_4454,N_4280);
nand U4546 (N_4546,N_4307,N_4340);
and U4547 (N_4547,N_4159,N_4049);
nor U4548 (N_4548,N_4316,N_4338);
and U4549 (N_4549,N_4190,N_4262);
nor U4550 (N_4550,N_4447,N_4388);
and U4551 (N_4551,N_4348,N_4195);
nor U4552 (N_4552,N_4375,N_4005);
and U4553 (N_4553,N_4135,N_4148);
or U4554 (N_4554,N_4281,N_4075);
nand U4555 (N_4555,N_4339,N_4235);
nor U4556 (N_4556,N_4089,N_4043);
nand U4557 (N_4557,N_4439,N_4016);
nand U4558 (N_4558,N_4441,N_4234);
xor U4559 (N_4559,N_4116,N_4133);
nand U4560 (N_4560,N_4036,N_4301);
nand U4561 (N_4561,N_4103,N_4023);
and U4562 (N_4562,N_4012,N_4477);
nor U4563 (N_4563,N_4039,N_4303);
nand U4564 (N_4564,N_4311,N_4427);
and U4565 (N_4565,N_4284,N_4216);
and U4566 (N_4566,N_4149,N_4020);
nor U4567 (N_4567,N_4115,N_4369);
xor U4568 (N_4568,N_4170,N_4177);
nand U4569 (N_4569,N_4451,N_4457);
nand U4570 (N_4570,N_4153,N_4275);
or U4571 (N_4571,N_4346,N_4249);
nand U4572 (N_4572,N_4017,N_4186);
or U4573 (N_4573,N_4260,N_4445);
and U4574 (N_4574,N_4068,N_4113);
nor U4575 (N_4575,N_4498,N_4136);
nand U4576 (N_4576,N_4327,N_4150);
and U4577 (N_4577,N_4352,N_4329);
xnor U4578 (N_4578,N_4448,N_4094);
and U4579 (N_4579,N_4489,N_4175);
nand U4580 (N_4580,N_4095,N_4084);
nand U4581 (N_4581,N_4400,N_4343);
and U4582 (N_4582,N_4488,N_4227);
nand U4583 (N_4583,N_4290,N_4099);
or U4584 (N_4584,N_4211,N_4332);
or U4585 (N_4585,N_4359,N_4458);
nand U4586 (N_4586,N_4003,N_4376);
and U4587 (N_4587,N_4493,N_4134);
nand U4588 (N_4588,N_4032,N_4404);
nor U4589 (N_4589,N_4002,N_4041);
xnor U4590 (N_4590,N_4231,N_4459);
nor U4591 (N_4591,N_4239,N_4333);
xnor U4592 (N_4592,N_4106,N_4387);
xnor U4593 (N_4593,N_4054,N_4419);
nor U4594 (N_4594,N_4413,N_4490);
nor U4595 (N_4595,N_4344,N_4442);
xor U4596 (N_4596,N_4070,N_4082);
nor U4597 (N_4597,N_4449,N_4014);
nor U4598 (N_4598,N_4285,N_4478);
nand U4599 (N_4599,N_4138,N_4288);
and U4600 (N_4600,N_4090,N_4072);
xnor U4601 (N_4601,N_4011,N_4100);
and U4602 (N_4602,N_4223,N_4292);
nor U4603 (N_4603,N_4293,N_4401);
xnor U4604 (N_4604,N_4168,N_4322);
nand U4605 (N_4605,N_4001,N_4204);
or U4606 (N_4606,N_4143,N_4233);
nor U4607 (N_4607,N_4432,N_4015);
nor U4608 (N_4608,N_4169,N_4192);
and U4609 (N_4609,N_4347,N_4373);
nor U4610 (N_4610,N_4467,N_4077);
nand U4611 (N_4611,N_4374,N_4205);
nand U4612 (N_4612,N_4045,N_4472);
nand U4613 (N_4613,N_4354,N_4294);
nand U4614 (N_4614,N_4208,N_4364);
xor U4615 (N_4615,N_4127,N_4161);
and U4616 (N_4616,N_4405,N_4416);
nand U4617 (N_4617,N_4297,N_4128);
and U4618 (N_4618,N_4033,N_4415);
or U4619 (N_4619,N_4365,N_4147);
nand U4620 (N_4620,N_4282,N_4270);
xnor U4621 (N_4621,N_4050,N_4087);
and U4622 (N_4622,N_4200,N_4395);
xor U4623 (N_4623,N_4209,N_4393);
and U4624 (N_4624,N_4360,N_4267);
nand U4625 (N_4625,N_4184,N_4480);
and U4626 (N_4626,N_4172,N_4120);
and U4627 (N_4627,N_4121,N_4218);
nor U4628 (N_4628,N_4057,N_4487);
nand U4629 (N_4629,N_4118,N_4382);
nand U4630 (N_4630,N_4222,N_4034);
nand U4631 (N_4631,N_4114,N_4225);
nor U4632 (N_4632,N_4398,N_4484);
nor U4633 (N_4633,N_4193,N_4386);
and U4634 (N_4634,N_4247,N_4283);
and U4635 (N_4635,N_4244,N_4243);
nand U4636 (N_4636,N_4318,N_4403);
or U4637 (N_4637,N_4126,N_4046);
or U4638 (N_4638,N_4309,N_4425);
nor U4639 (N_4639,N_4492,N_4479);
nor U4640 (N_4640,N_4461,N_4105);
and U4641 (N_4641,N_4018,N_4381);
nor U4642 (N_4642,N_4232,N_4132);
nand U4643 (N_4643,N_4051,N_4379);
or U4644 (N_4644,N_4066,N_4269);
nand U4645 (N_4645,N_4083,N_4250);
nand U4646 (N_4646,N_4119,N_4217);
or U4647 (N_4647,N_4263,N_4058);
nand U4648 (N_4648,N_4334,N_4009);
and U4649 (N_4649,N_4361,N_4142);
nand U4650 (N_4650,N_4366,N_4007);
nor U4651 (N_4651,N_4214,N_4074);
or U4652 (N_4652,N_4470,N_4213);
or U4653 (N_4653,N_4463,N_4131);
nor U4654 (N_4654,N_4412,N_4409);
nand U4655 (N_4655,N_4076,N_4420);
nor U4656 (N_4656,N_4278,N_4310);
xor U4657 (N_4657,N_4314,N_4004);
and U4658 (N_4658,N_4224,N_4299);
nor U4659 (N_4659,N_4273,N_4221);
xor U4660 (N_4660,N_4437,N_4483);
and U4661 (N_4661,N_4151,N_4362);
or U4662 (N_4662,N_4305,N_4345);
and U4663 (N_4663,N_4433,N_4174);
nor U4664 (N_4664,N_4245,N_4380);
nand U4665 (N_4665,N_4080,N_4471);
and U4666 (N_4666,N_4164,N_4335);
nand U4667 (N_4667,N_4085,N_4378);
nand U4668 (N_4668,N_4368,N_4469);
or U4669 (N_4669,N_4258,N_4160);
nor U4670 (N_4670,N_4424,N_4274);
nand U4671 (N_4671,N_4165,N_4367);
nor U4672 (N_4672,N_4130,N_4256);
nand U4673 (N_4673,N_4444,N_4254);
nor U4674 (N_4674,N_4196,N_4440);
or U4675 (N_4675,N_4097,N_4320);
nand U4676 (N_4676,N_4246,N_4157);
and U4677 (N_4677,N_4187,N_4063);
and U4678 (N_4678,N_4123,N_4237);
xor U4679 (N_4679,N_4155,N_4037);
and U4680 (N_4680,N_4315,N_4462);
nor U4681 (N_4681,N_4065,N_4210);
nand U4682 (N_4682,N_4466,N_4240);
nand U4683 (N_4683,N_4272,N_4473);
and U4684 (N_4684,N_4104,N_4474);
nor U4685 (N_4685,N_4266,N_4203);
nor U4686 (N_4686,N_4298,N_4093);
nor U4687 (N_4687,N_4129,N_4008);
nor U4688 (N_4688,N_4286,N_4319);
or U4689 (N_4689,N_4047,N_4438);
and U4690 (N_4690,N_4055,N_4062);
nor U4691 (N_4691,N_4497,N_4158);
nor U4692 (N_4692,N_4167,N_4428);
and U4693 (N_4693,N_4180,N_4342);
nor U4694 (N_4694,N_4079,N_4086);
and U4695 (N_4695,N_4191,N_4189);
nor U4696 (N_4696,N_4199,N_4435);
or U4697 (N_4697,N_4026,N_4251);
or U4698 (N_4698,N_4152,N_4052);
xnor U4699 (N_4699,N_4107,N_4414);
or U4700 (N_4700,N_4178,N_4464);
nor U4701 (N_4701,N_4350,N_4179);
or U4702 (N_4702,N_4176,N_4185);
nand U4703 (N_4703,N_4124,N_4434);
or U4704 (N_4704,N_4475,N_4069);
or U4705 (N_4705,N_4188,N_4029);
nor U4706 (N_4706,N_4040,N_4308);
nor U4707 (N_4707,N_4220,N_4248);
and U4708 (N_4708,N_4485,N_4257);
nor U4709 (N_4709,N_4183,N_4141);
and U4710 (N_4710,N_4394,N_4241);
nor U4711 (N_4711,N_4494,N_4166);
xnor U4712 (N_4712,N_4349,N_4325);
nand U4713 (N_4713,N_4056,N_4302);
nand U4714 (N_4714,N_4162,N_4064);
xor U4715 (N_4715,N_4230,N_4236);
or U4716 (N_4716,N_4411,N_4035);
nor U4717 (N_4717,N_4291,N_4486);
or U4718 (N_4718,N_4098,N_4202);
nand U4719 (N_4719,N_4407,N_4092);
and U4720 (N_4720,N_4030,N_4429);
or U4721 (N_4721,N_4073,N_4430);
nor U4722 (N_4722,N_4306,N_4201);
and U4723 (N_4723,N_4371,N_4102);
nor U4724 (N_4724,N_4194,N_4357);
nand U4725 (N_4725,N_4431,N_4370);
nand U4726 (N_4726,N_4330,N_4324);
nor U4727 (N_4727,N_4061,N_4372);
and U4728 (N_4728,N_4091,N_4125);
nand U4729 (N_4729,N_4219,N_4010);
and U4730 (N_4730,N_4242,N_4110);
nand U4731 (N_4731,N_4328,N_4426);
or U4732 (N_4732,N_4476,N_4025);
and U4733 (N_4733,N_4059,N_4228);
nor U4734 (N_4734,N_4336,N_4145);
or U4735 (N_4735,N_4101,N_4027);
and U4736 (N_4736,N_4465,N_4385);
nor U4737 (N_4737,N_4067,N_4048);
nand U4738 (N_4738,N_4351,N_4450);
nor U4739 (N_4739,N_4261,N_4456);
nor U4740 (N_4740,N_4422,N_4390);
or U4741 (N_4741,N_4144,N_4452);
nand U4742 (N_4742,N_4481,N_4287);
and U4743 (N_4743,N_4499,N_4323);
nand U4744 (N_4744,N_4137,N_4268);
nor U4745 (N_4745,N_4331,N_4277);
or U4746 (N_4746,N_4171,N_4163);
nand U4747 (N_4747,N_4078,N_4295);
and U4748 (N_4748,N_4389,N_4198);
nor U4749 (N_4749,N_4206,N_4482);
or U4750 (N_4750,N_4498,N_4304);
and U4751 (N_4751,N_4201,N_4072);
and U4752 (N_4752,N_4000,N_4178);
nor U4753 (N_4753,N_4155,N_4101);
and U4754 (N_4754,N_4185,N_4199);
and U4755 (N_4755,N_4267,N_4224);
or U4756 (N_4756,N_4321,N_4252);
xor U4757 (N_4757,N_4340,N_4105);
nor U4758 (N_4758,N_4330,N_4190);
or U4759 (N_4759,N_4328,N_4252);
nand U4760 (N_4760,N_4139,N_4269);
or U4761 (N_4761,N_4490,N_4374);
nand U4762 (N_4762,N_4437,N_4024);
or U4763 (N_4763,N_4319,N_4484);
nand U4764 (N_4764,N_4336,N_4459);
or U4765 (N_4765,N_4095,N_4390);
nor U4766 (N_4766,N_4343,N_4272);
nor U4767 (N_4767,N_4200,N_4139);
and U4768 (N_4768,N_4014,N_4264);
nor U4769 (N_4769,N_4134,N_4192);
nor U4770 (N_4770,N_4356,N_4040);
and U4771 (N_4771,N_4495,N_4091);
nor U4772 (N_4772,N_4231,N_4042);
nor U4773 (N_4773,N_4388,N_4333);
or U4774 (N_4774,N_4499,N_4362);
and U4775 (N_4775,N_4063,N_4323);
xor U4776 (N_4776,N_4400,N_4078);
nand U4777 (N_4777,N_4126,N_4035);
or U4778 (N_4778,N_4468,N_4311);
or U4779 (N_4779,N_4254,N_4427);
nor U4780 (N_4780,N_4247,N_4225);
nand U4781 (N_4781,N_4273,N_4113);
xor U4782 (N_4782,N_4311,N_4001);
nor U4783 (N_4783,N_4412,N_4439);
or U4784 (N_4784,N_4318,N_4253);
nor U4785 (N_4785,N_4091,N_4130);
and U4786 (N_4786,N_4491,N_4035);
or U4787 (N_4787,N_4192,N_4184);
and U4788 (N_4788,N_4482,N_4440);
nor U4789 (N_4789,N_4331,N_4351);
or U4790 (N_4790,N_4480,N_4331);
or U4791 (N_4791,N_4381,N_4328);
nand U4792 (N_4792,N_4446,N_4341);
nor U4793 (N_4793,N_4094,N_4490);
nor U4794 (N_4794,N_4109,N_4227);
nand U4795 (N_4795,N_4453,N_4199);
nor U4796 (N_4796,N_4116,N_4265);
and U4797 (N_4797,N_4189,N_4211);
and U4798 (N_4798,N_4231,N_4088);
nor U4799 (N_4799,N_4454,N_4260);
and U4800 (N_4800,N_4211,N_4255);
nand U4801 (N_4801,N_4127,N_4220);
nor U4802 (N_4802,N_4053,N_4391);
nand U4803 (N_4803,N_4060,N_4076);
and U4804 (N_4804,N_4394,N_4328);
and U4805 (N_4805,N_4209,N_4237);
and U4806 (N_4806,N_4231,N_4154);
nand U4807 (N_4807,N_4256,N_4461);
xnor U4808 (N_4808,N_4471,N_4158);
xnor U4809 (N_4809,N_4298,N_4444);
and U4810 (N_4810,N_4312,N_4280);
nand U4811 (N_4811,N_4180,N_4474);
nand U4812 (N_4812,N_4162,N_4286);
nor U4813 (N_4813,N_4113,N_4301);
nand U4814 (N_4814,N_4105,N_4495);
and U4815 (N_4815,N_4131,N_4177);
and U4816 (N_4816,N_4077,N_4069);
or U4817 (N_4817,N_4093,N_4246);
and U4818 (N_4818,N_4386,N_4151);
or U4819 (N_4819,N_4022,N_4458);
or U4820 (N_4820,N_4474,N_4324);
nor U4821 (N_4821,N_4386,N_4084);
nor U4822 (N_4822,N_4230,N_4176);
nand U4823 (N_4823,N_4062,N_4085);
nand U4824 (N_4824,N_4458,N_4345);
nand U4825 (N_4825,N_4444,N_4469);
nor U4826 (N_4826,N_4162,N_4151);
and U4827 (N_4827,N_4494,N_4372);
nor U4828 (N_4828,N_4123,N_4428);
xnor U4829 (N_4829,N_4061,N_4356);
and U4830 (N_4830,N_4061,N_4229);
and U4831 (N_4831,N_4164,N_4299);
or U4832 (N_4832,N_4183,N_4469);
and U4833 (N_4833,N_4306,N_4104);
and U4834 (N_4834,N_4271,N_4007);
and U4835 (N_4835,N_4268,N_4307);
nand U4836 (N_4836,N_4064,N_4366);
and U4837 (N_4837,N_4229,N_4292);
nor U4838 (N_4838,N_4135,N_4198);
and U4839 (N_4839,N_4111,N_4271);
nand U4840 (N_4840,N_4214,N_4381);
nand U4841 (N_4841,N_4400,N_4494);
or U4842 (N_4842,N_4379,N_4133);
and U4843 (N_4843,N_4127,N_4086);
xor U4844 (N_4844,N_4486,N_4490);
or U4845 (N_4845,N_4122,N_4448);
or U4846 (N_4846,N_4463,N_4467);
nor U4847 (N_4847,N_4134,N_4317);
or U4848 (N_4848,N_4159,N_4280);
or U4849 (N_4849,N_4352,N_4097);
nand U4850 (N_4850,N_4163,N_4179);
or U4851 (N_4851,N_4046,N_4409);
nor U4852 (N_4852,N_4099,N_4097);
nand U4853 (N_4853,N_4166,N_4338);
or U4854 (N_4854,N_4387,N_4161);
nor U4855 (N_4855,N_4454,N_4104);
xnor U4856 (N_4856,N_4261,N_4471);
or U4857 (N_4857,N_4055,N_4219);
or U4858 (N_4858,N_4247,N_4432);
nand U4859 (N_4859,N_4421,N_4356);
xor U4860 (N_4860,N_4432,N_4087);
and U4861 (N_4861,N_4351,N_4384);
or U4862 (N_4862,N_4392,N_4273);
nand U4863 (N_4863,N_4235,N_4142);
nand U4864 (N_4864,N_4272,N_4119);
or U4865 (N_4865,N_4167,N_4397);
nor U4866 (N_4866,N_4415,N_4407);
nor U4867 (N_4867,N_4055,N_4113);
nand U4868 (N_4868,N_4262,N_4189);
nand U4869 (N_4869,N_4010,N_4009);
xnor U4870 (N_4870,N_4080,N_4085);
and U4871 (N_4871,N_4226,N_4132);
nand U4872 (N_4872,N_4063,N_4201);
and U4873 (N_4873,N_4269,N_4349);
xnor U4874 (N_4874,N_4401,N_4021);
nand U4875 (N_4875,N_4118,N_4241);
nand U4876 (N_4876,N_4145,N_4458);
nor U4877 (N_4877,N_4297,N_4039);
and U4878 (N_4878,N_4094,N_4220);
xor U4879 (N_4879,N_4352,N_4445);
nand U4880 (N_4880,N_4452,N_4374);
nand U4881 (N_4881,N_4076,N_4438);
or U4882 (N_4882,N_4125,N_4359);
and U4883 (N_4883,N_4257,N_4499);
and U4884 (N_4884,N_4235,N_4483);
or U4885 (N_4885,N_4451,N_4141);
nand U4886 (N_4886,N_4379,N_4328);
and U4887 (N_4887,N_4036,N_4325);
and U4888 (N_4888,N_4436,N_4136);
nor U4889 (N_4889,N_4219,N_4146);
nor U4890 (N_4890,N_4411,N_4308);
and U4891 (N_4891,N_4294,N_4379);
nor U4892 (N_4892,N_4365,N_4097);
nor U4893 (N_4893,N_4010,N_4384);
nor U4894 (N_4894,N_4468,N_4234);
nand U4895 (N_4895,N_4026,N_4292);
or U4896 (N_4896,N_4187,N_4127);
nand U4897 (N_4897,N_4284,N_4351);
nor U4898 (N_4898,N_4439,N_4401);
and U4899 (N_4899,N_4137,N_4163);
or U4900 (N_4900,N_4482,N_4252);
or U4901 (N_4901,N_4484,N_4428);
xor U4902 (N_4902,N_4277,N_4107);
nand U4903 (N_4903,N_4414,N_4293);
nand U4904 (N_4904,N_4018,N_4248);
nor U4905 (N_4905,N_4102,N_4277);
xnor U4906 (N_4906,N_4381,N_4273);
or U4907 (N_4907,N_4315,N_4421);
and U4908 (N_4908,N_4079,N_4336);
and U4909 (N_4909,N_4012,N_4234);
nor U4910 (N_4910,N_4189,N_4402);
or U4911 (N_4911,N_4323,N_4262);
xor U4912 (N_4912,N_4474,N_4486);
and U4913 (N_4913,N_4452,N_4018);
and U4914 (N_4914,N_4222,N_4497);
xnor U4915 (N_4915,N_4484,N_4269);
or U4916 (N_4916,N_4482,N_4415);
nor U4917 (N_4917,N_4132,N_4304);
nand U4918 (N_4918,N_4274,N_4435);
and U4919 (N_4919,N_4479,N_4365);
nor U4920 (N_4920,N_4092,N_4098);
or U4921 (N_4921,N_4488,N_4005);
nand U4922 (N_4922,N_4108,N_4439);
nor U4923 (N_4923,N_4314,N_4036);
or U4924 (N_4924,N_4189,N_4323);
nor U4925 (N_4925,N_4181,N_4366);
nand U4926 (N_4926,N_4162,N_4154);
and U4927 (N_4927,N_4430,N_4317);
xor U4928 (N_4928,N_4267,N_4455);
and U4929 (N_4929,N_4392,N_4438);
and U4930 (N_4930,N_4049,N_4316);
and U4931 (N_4931,N_4069,N_4067);
and U4932 (N_4932,N_4401,N_4037);
or U4933 (N_4933,N_4059,N_4349);
nor U4934 (N_4934,N_4037,N_4417);
nand U4935 (N_4935,N_4196,N_4458);
nor U4936 (N_4936,N_4180,N_4359);
and U4937 (N_4937,N_4367,N_4256);
nand U4938 (N_4938,N_4173,N_4149);
nand U4939 (N_4939,N_4398,N_4041);
nand U4940 (N_4940,N_4288,N_4206);
nor U4941 (N_4941,N_4467,N_4365);
and U4942 (N_4942,N_4340,N_4082);
or U4943 (N_4943,N_4426,N_4326);
nand U4944 (N_4944,N_4087,N_4204);
nor U4945 (N_4945,N_4212,N_4056);
or U4946 (N_4946,N_4138,N_4470);
and U4947 (N_4947,N_4315,N_4181);
nor U4948 (N_4948,N_4492,N_4396);
nand U4949 (N_4949,N_4138,N_4394);
xnor U4950 (N_4950,N_4063,N_4079);
or U4951 (N_4951,N_4373,N_4166);
or U4952 (N_4952,N_4240,N_4369);
and U4953 (N_4953,N_4423,N_4043);
nand U4954 (N_4954,N_4359,N_4374);
or U4955 (N_4955,N_4016,N_4230);
and U4956 (N_4956,N_4407,N_4116);
or U4957 (N_4957,N_4001,N_4127);
or U4958 (N_4958,N_4105,N_4099);
nor U4959 (N_4959,N_4397,N_4191);
and U4960 (N_4960,N_4036,N_4006);
xor U4961 (N_4961,N_4347,N_4004);
nor U4962 (N_4962,N_4238,N_4292);
nor U4963 (N_4963,N_4232,N_4481);
nor U4964 (N_4964,N_4289,N_4128);
or U4965 (N_4965,N_4100,N_4075);
and U4966 (N_4966,N_4027,N_4000);
nand U4967 (N_4967,N_4380,N_4172);
and U4968 (N_4968,N_4362,N_4126);
xnor U4969 (N_4969,N_4259,N_4391);
nand U4970 (N_4970,N_4352,N_4176);
and U4971 (N_4971,N_4038,N_4241);
nor U4972 (N_4972,N_4156,N_4064);
nand U4973 (N_4973,N_4483,N_4306);
and U4974 (N_4974,N_4460,N_4191);
and U4975 (N_4975,N_4166,N_4384);
nor U4976 (N_4976,N_4333,N_4322);
nor U4977 (N_4977,N_4289,N_4166);
nand U4978 (N_4978,N_4016,N_4266);
or U4979 (N_4979,N_4040,N_4438);
or U4980 (N_4980,N_4128,N_4474);
nand U4981 (N_4981,N_4315,N_4425);
or U4982 (N_4982,N_4262,N_4098);
or U4983 (N_4983,N_4278,N_4239);
and U4984 (N_4984,N_4346,N_4425);
nor U4985 (N_4985,N_4453,N_4175);
and U4986 (N_4986,N_4025,N_4387);
nor U4987 (N_4987,N_4302,N_4028);
nor U4988 (N_4988,N_4316,N_4451);
or U4989 (N_4989,N_4443,N_4201);
nor U4990 (N_4990,N_4201,N_4315);
nand U4991 (N_4991,N_4154,N_4487);
nand U4992 (N_4992,N_4221,N_4322);
and U4993 (N_4993,N_4491,N_4317);
nand U4994 (N_4994,N_4176,N_4226);
nand U4995 (N_4995,N_4175,N_4279);
and U4996 (N_4996,N_4464,N_4298);
nand U4997 (N_4997,N_4042,N_4314);
xor U4998 (N_4998,N_4353,N_4387);
xnor U4999 (N_4999,N_4172,N_4176);
nor U5000 (N_5000,N_4678,N_4915);
and U5001 (N_5001,N_4842,N_4716);
or U5002 (N_5002,N_4742,N_4932);
nor U5003 (N_5003,N_4775,N_4816);
and U5004 (N_5004,N_4641,N_4905);
nand U5005 (N_5005,N_4501,N_4783);
and U5006 (N_5006,N_4881,N_4587);
nor U5007 (N_5007,N_4500,N_4575);
nand U5008 (N_5008,N_4569,N_4822);
nand U5009 (N_5009,N_4829,N_4523);
nor U5010 (N_5010,N_4752,N_4647);
or U5011 (N_5011,N_4764,N_4962);
and U5012 (N_5012,N_4815,N_4632);
xnor U5013 (N_5013,N_4563,N_4703);
nor U5014 (N_5014,N_4668,N_4934);
or U5015 (N_5015,N_4991,N_4894);
xnor U5016 (N_5016,N_4929,N_4795);
nand U5017 (N_5017,N_4824,N_4719);
and U5018 (N_5018,N_4707,N_4662);
and U5019 (N_5019,N_4768,N_4924);
or U5020 (N_5020,N_4959,N_4511);
or U5021 (N_5021,N_4540,N_4698);
or U5022 (N_5022,N_4600,N_4780);
and U5023 (N_5023,N_4903,N_4895);
nor U5024 (N_5024,N_4510,N_4708);
nand U5025 (N_5025,N_4793,N_4610);
nor U5026 (N_5026,N_4787,N_4611);
xnor U5027 (N_5027,N_4670,N_4725);
or U5028 (N_5028,N_4505,N_4831);
and U5029 (N_5029,N_4536,N_4811);
nor U5030 (N_5030,N_4933,N_4539);
or U5031 (N_5031,N_4701,N_4590);
nor U5032 (N_5032,N_4858,N_4608);
or U5033 (N_5033,N_4530,N_4772);
nand U5034 (N_5034,N_4603,N_4799);
nand U5035 (N_5035,N_4748,N_4879);
nand U5036 (N_5036,N_4872,N_4550);
nor U5037 (N_5037,N_4908,N_4502);
or U5038 (N_5038,N_4524,N_4847);
and U5039 (N_5039,N_4759,N_4766);
nand U5040 (N_5040,N_4921,N_4615);
or U5041 (N_5041,N_4627,N_4869);
nand U5042 (N_5042,N_4970,N_4784);
nor U5043 (N_5043,N_4988,N_4901);
nand U5044 (N_5044,N_4947,N_4837);
nor U5045 (N_5045,N_4572,N_4955);
nand U5046 (N_5046,N_4973,N_4843);
or U5047 (N_5047,N_4601,N_4612);
nand U5048 (N_5048,N_4969,N_4711);
or U5049 (N_5049,N_4674,N_4567);
nor U5050 (N_5050,N_4856,N_4570);
and U5051 (N_5051,N_4941,N_4622);
and U5052 (N_5052,N_4981,N_4907);
and U5053 (N_5053,N_4912,N_4534);
and U5054 (N_5054,N_4938,N_4994);
or U5055 (N_5055,N_4697,N_4814);
and U5056 (N_5056,N_4520,N_4864);
and U5057 (N_5057,N_4918,N_4914);
or U5058 (N_5058,N_4650,N_4866);
xor U5059 (N_5059,N_4800,N_4586);
nor U5060 (N_5060,N_4626,N_4585);
or U5061 (N_5061,N_4840,N_4664);
nand U5062 (N_5062,N_4635,N_4685);
nand U5063 (N_5063,N_4559,N_4598);
and U5064 (N_5064,N_4715,N_4712);
and U5065 (N_5065,N_4553,N_4614);
nand U5066 (N_5066,N_4665,N_4873);
nand U5067 (N_5067,N_4757,N_4740);
nand U5068 (N_5068,N_4850,N_4582);
nand U5069 (N_5069,N_4583,N_4737);
nor U5070 (N_5070,N_4648,N_4566);
nor U5071 (N_5071,N_4589,N_4761);
nand U5072 (N_5072,N_4944,N_4892);
nand U5073 (N_5073,N_4628,N_4774);
and U5074 (N_5074,N_4871,N_4957);
and U5075 (N_5075,N_4637,N_4532);
nand U5076 (N_5076,N_4667,N_4960);
xnor U5077 (N_5077,N_4926,N_4722);
nand U5078 (N_5078,N_4909,N_4721);
or U5079 (N_5079,N_4578,N_4998);
or U5080 (N_5080,N_4581,N_4560);
and U5081 (N_5081,N_4913,N_4541);
xor U5082 (N_5082,N_4551,N_4887);
and U5083 (N_5083,N_4577,N_4718);
and U5084 (N_5084,N_4651,N_4948);
or U5085 (N_5085,N_4939,N_4522);
nor U5086 (N_5086,N_4896,N_4971);
nor U5087 (N_5087,N_4936,N_4773);
nor U5088 (N_5088,N_4823,N_4609);
nor U5089 (N_5089,N_4630,N_4855);
or U5090 (N_5090,N_4834,N_4576);
xor U5091 (N_5091,N_4767,N_4555);
or U5092 (N_5092,N_4841,N_4789);
nor U5093 (N_5093,N_4958,N_4681);
nor U5094 (N_5094,N_4504,N_4616);
xnor U5095 (N_5095,N_4977,N_4805);
xor U5096 (N_5096,N_4758,N_4756);
nand U5097 (N_5097,N_4556,N_4839);
or U5098 (N_5098,N_4952,N_4561);
nand U5099 (N_5099,N_4531,N_4770);
nand U5100 (N_5100,N_4683,N_4862);
or U5101 (N_5101,N_4516,N_4597);
or U5102 (N_5102,N_4514,N_4705);
and U5103 (N_5103,N_4694,N_4785);
and U5104 (N_5104,N_4911,N_4621);
or U5105 (N_5105,N_4517,N_4638);
and U5106 (N_5106,N_4591,N_4853);
xnor U5107 (N_5107,N_4821,N_4830);
nand U5108 (N_5108,N_4910,N_4927);
nor U5109 (N_5109,N_4673,N_4968);
xor U5110 (N_5110,N_4620,N_4663);
xnor U5111 (N_5111,N_4644,N_4642);
nor U5112 (N_5112,N_4671,N_4844);
nor U5113 (N_5113,N_4564,N_4845);
and U5114 (N_5114,N_4739,N_4625);
nor U5115 (N_5115,N_4992,N_4966);
nand U5116 (N_5116,N_4538,N_4906);
nor U5117 (N_5117,N_4643,N_4868);
nor U5118 (N_5118,N_4863,N_4798);
nand U5119 (N_5119,N_4930,N_4696);
nand U5120 (N_5120,N_4940,N_4754);
nand U5121 (N_5121,N_4883,N_4857);
nor U5122 (N_5122,N_4702,N_4714);
xnor U5123 (N_5123,N_4506,N_4931);
xnor U5124 (N_5124,N_4976,N_4942);
nand U5125 (N_5125,N_4736,N_4848);
or U5126 (N_5126,N_4937,N_4781);
nor U5127 (N_5127,N_4552,N_4579);
and U5128 (N_5128,N_4755,N_4897);
nand U5129 (N_5129,N_4746,N_4717);
nand U5130 (N_5130,N_4794,N_4870);
or U5131 (N_5131,N_4972,N_4571);
or U5132 (N_5132,N_4568,N_4880);
or U5133 (N_5133,N_4710,N_4509);
or U5134 (N_5134,N_4623,N_4996);
nor U5135 (N_5135,N_4886,N_4920);
and U5136 (N_5136,N_4828,N_4750);
nand U5137 (N_5137,N_4777,N_4956);
nor U5138 (N_5138,N_4876,N_4513);
nor U5139 (N_5139,N_4925,N_4846);
or U5140 (N_5140,N_4558,N_4923);
nand U5141 (N_5141,N_4993,N_4796);
nand U5142 (N_5142,N_4877,N_4535);
and U5143 (N_5143,N_4657,N_4729);
and U5144 (N_5144,N_4954,N_4951);
nor U5145 (N_5145,N_4744,N_4860);
and U5146 (N_5146,N_4997,N_4990);
nor U5147 (N_5147,N_4688,N_4604);
or U5148 (N_5148,N_4779,N_4606);
nor U5149 (N_5149,N_4659,N_4987);
or U5150 (N_5150,N_4809,N_4691);
or U5151 (N_5151,N_4543,N_4588);
or U5152 (N_5152,N_4782,N_4889);
and U5153 (N_5153,N_4602,N_4618);
nor U5154 (N_5154,N_4521,N_4653);
nor U5155 (N_5155,N_4825,N_4900);
nand U5156 (N_5156,N_4527,N_4593);
or U5157 (N_5157,N_4528,N_4695);
and U5158 (N_5158,N_4935,N_4649);
nor U5159 (N_5159,N_4919,N_4646);
and U5160 (N_5160,N_4542,N_4961);
xor U5161 (N_5161,N_4833,N_4865);
and U5162 (N_5162,N_4666,N_4804);
nor U5163 (N_5163,N_4978,N_4675);
nand U5164 (N_5164,N_4726,N_4706);
or U5165 (N_5165,N_4854,N_4749);
nand U5166 (N_5166,N_4633,N_4786);
nand U5167 (N_5167,N_4547,N_4916);
or U5168 (N_5168,N_4946,N_4745);
nand U5169 (N_5169,N_4503,N_4967);
or U5170 (N_5170,N_4806,N_4557);
nand U5171 (N_5171,N_4669,N_4732);
nor U5172 (N_5172,N_4629,N_4899);
or U5173 (N_5173,N_4655,N_4974);
nor U5174 (N_5174,N_4596,N_4682);
nor U5175 (N_5175,N_4819,N_4891);
or U5176 (N_5176,N_4676,N_4943);
nor U5177 (N_5177,N_4645,N_4904);
and U5178 (N_5178,N_4617,N_4874);
nand U5179 (N_5179,N_4654,N_4738);
nand U5180 (N_5180,N_4922,N_4700);
or U5181 (N_5181,N_4763,N_4660);
xnor U5182 (N_5182,N_4677,N_4776);
nor U5183 (N_5183,N_4580,N_4661);
nand U5184 (N_5184,N_4544,N_4562);
nor U5185 (N_5185,N_4803,N_4975);
xor U5186 (N_5186,N_4747,N_4945);
or U5187 (N_5187,N_4686,N_4788);
nand U5188 (N_5188,N_4753,N_4512);
or U5189 (N_5189,N_4878,N_4999);
nor U5190 (N_5190,N_4672,N_4679);
nor U5191 (N_5191,N_4802,N_4594);
nor U5192 (N_5192,N_4709,N_4765);
xnor U5193 (N_5193,N_4545,N_4734);
nor U5194 (N_5194,N_4985,N_4508);
nand U5195 (N_5195,N_4861,N_4989);
nand U5196 (N_5196,N_4515,N_4980);
or U5197 (N_5197,N_4890,N_4902);
nand U5198 (N_5198,N_4982,N_4859);
xnor U5199 (N_5199,N_4525,N_4573);
nor U5200 (N_5200,N_4790,N_4713);
or U5201 (N_5201,N_4727,N_4760);
and U5202 (N_5202,N_4885,N_4546);
nor U5203 (N_5203,N_4995,N_4875);
and U5204 (N_5204,N_4537,N_4983);
xor U5205 (N_5205,N_4963,N_4986);
nor U5206 (N_5206,N_4704,N_4827);
nor U5207 (N_5207,N_4836,N_4979);
nand U5208 (N_5208,N_4605,N_4826);
and U5209 (N_5209,N_4634,N_4818);
or U5210 (N_5210,N_4730,N_4928);
or U5211 (N_5211,N_4797,N_4518);
and U5212 (N_5212,N_4820,N_4882);
nand U5213 (N_5213,N_4852,N_4807);
nand U5214 (N_5214,N_4964,N_4689);
nor U5215 (N_5215,N_4751,N_4771);
and U5216 (N_5216,N_4731,N_4724);
and U5217 (N_5217,N_4808,N_4723);
and U5218 (N_5218,N_4624,N_4743);
nand U5219 (N_5219,N_4599,N_4680);
and U5220 (N_5220,N_4526,N_4607);
nor U5221 (N_5221,N_4838,N_4817);
nor U5222 (N_5222,N_4762,N_4699);
nand U5223 (N_5223,N_4953,N_4574);
and U5224 (N_5224,N_4984,N_4720);
nand U5225 (N_5225,N_4884,N_4554);
nor U5226 (N_5226,N_4832,N_4965);
nand U5227 (N_5227,N_4584,N_4619);
or U5228 (N_5228,N_4733,N_4684);
and U5229 (N_5229,N_4813,N_4636);
and U5230 (N_5230,N_4549,N_4507);
nand U5231 (N_5231,N_4791,N_4640);
nor U5232 (N_5232,N_4656,N_4565);
and U5233 (N_5233,N_4810,N_4851);
nand U5234 (N_5234,N_4867,N_4592);
or U5235 (N_5235,N_4769,N_4658);
or U5236 (N_5236,N_4898,N_4693);
nor U5237 (N_5237,N_4835,N_4690);
or U5238 (N_5238,N_4893,N_4917);
and U5239 (N_5239,N_4639,N_4950);
or U5240 (N_5240,N_4548,N_4687);
or U5241 (N_5241,N_4741,N_4888);
nor U5242 (N_5242,N_4533,N_4519);
and U5243 (N_5243,N_4778,N_4595);
or U5244 (N_5244,N_4631,N_4812);
or U5245 (N_5245,N_4801,N_4735);
or U5246 (N_5246,N_4792,N_4613);
nand U5247 (N_5247,N_4692,N_4849);
nor U5248 (N_5248,N_4949,N_4728);
or U5249 (N_5249,N_4529,N_4652);
or U5250 (N_5250,N_4509,N_4954);
nor U5251 (N_5251,N_4876,N_4917);
nand U5252 (N_5252,N_4592,N_4939);
or U5253 (N_5253,N_4633,N_4534);
or U5254 (N_5254,N_4558,N_4851);
xnor U5255 (N_5255,N_4937,N_4577);
or U5256 (N_5256,N_4906,N_4715);
nor U5257 (N_5257,N_4567,N_4635);
and U5258 (N_5258,N_4561,N_4709);
nor U5259 (N_5259,N_4876,N_4720);
nand U5260 (N_5260,N_4806,N_4779);
and U5261 (N_5261,N_4610,N_4963);
or U5262 (N_5262,N_4927,N_4647);
nand U5263 (N_5263,N_4692,N_4770);
xor U5264 (N_5264,N_4615,N_4821);
or U5265 (N_5265,N_4730,N_4520);
nand U5266 (N_5266,N_4725,N_4558);
xnor U5267 (N_5267,N_4757,N_4858);
nand U5268 (N_5268,N_4803,N_4831);
or U5269 (N_5269,N_4868,N_4754);
nand U5270 (N_5270,N_4711,N_4867);
and U5271 (N_5271,N_4774,N_4962);
and U5272 (N_5272,N_4915,N_4640);
xor U5273 (N_5273,N_4734,N_4618);
and U5274 (N_5274,N_4630,N_4794);
xor U5275 (N_5275,N_4972,N_4927);
and U5276 (N_5276,N_4741,N_4870);
or U5277 (N_5277,N_4821,N_4543);
xor U5278 (N_5278,N_4555,N_4709);
nor U5279 (N_5279,N_4555,N_4507);
and U5280 (N_5280,N_4973,N_4965);
or U5281 (N_5281,N_4603,N_4635);
or U5282 (N_5282,N_4706,N_4985);
nand U5283 (N_5283,N_4680,N_4986);
or U5284 (N_5284,N_4966,N_4834);
nand U5285 (N_5285,N_4860,N_4612);
xor U5286 (N_5286,N_4955,N_4901);
or U5287 (N_5287,N_4623,N_4982);
nor U5288 (N_5288,N_4910,N_4906);
or U5289 (N_5289,N_4987,N_4502);
xor U5290 (N_5290,N_4661,N_4850);
nand U5291 (N_5291,N_4679,N_4697);
nand U5292 (N_5292,N_4857,N_4783);
or U5293 (N_5293,N_4970,N_4662);
nor U5294 (N_5294,N_4507,N_4900);
or U5295 (N_5295,N_4706,N_4652);
xnor U5296 (N_5296,N_4998,N_4593);
nor U5297 (N_5297,N_4824,N_4764);
nand U5298 (N_5298,N_4816,N_4785);
and U5299 (N_5299,N_4966,N_4752);
and U5300 (N_5300,N_4882,N_4939);
and U5301 (N_5301,N_4865,N_4824);
nand U5302 (N_5302,N_4736,N_4953);
nor U5303 (N_5303,N_4814,N_4924);
and U5304 (N_5304,N_4958,N_4515);
or U5305 (N_5305,N_4799,N_4804);
nor U5306 (N_5306,N_4644,N_4505);
and U5307 (N_5307,N_4541,N_4600);
nor U5308 (N_5308,N_4509,N_4564);
nand U5309 (N_5309,N_4665,N_4744);
xor U5310 (N_5310,N_4670,N_4916);
or U5311 (N_5311,N_4662,N_4895);
nand U5312 (N_5312,N_4720,N_4520);
or U5313 (N_5313,N_4792,N_4666);
and U5314 (N_5314,N_4922,N_4829);
or U5315 (N_5315,N_4613,N_4848);
and U5316 (N_5316,N_4628,N_4678);
and U5317 (N_5317,N_4706,N_4621);
nor U5318 (N_5318,N_4640,N_4944);
and U5319 (N_5319,N_4649,N_4780);
and U5320 (N_5320,N_4711,N_4933);
nand U5321 (N_5321,N_4873,N_4868);
nor U5322 (N_5322,N_4939,N_4684);
and U5323 (N_5323,N_4794,N_4791);
nor U5324 (N_5324,N_4976,N_4627);
or U5325 (N_5325,N_4819,N_4514);
nor U5326 (N_5326,N_4746,N_4572);
nand U5327 (N_5327,N_4904,N_4924);
xnor U5328 (N_5328,N_4843,N_4965);
or U5329 (N_5329,N_4863,N_4711);
or U5330 (N_5330,N_4550,N_4570);
and U5331 (N_5331,N_4719,N_4651);
or U5332 (N_5332,N_4697,N_4563);
nand U5333 (N_5333,N_4575,N_4508);
and U5334 (N_5334,N_4838,N_4502);
nand U5335 (N_5335,N_4600,N_4863);
nor U5336 (N_5336,N_4778,N_4922);
or U5337 (N_5337,N_4958,N_4585);
nand U5338 (N_5338,N_4816,N_4923);
nor U5339 (N_5339,N_4559,N_4719);
or U5340 (N_5340,N_4923,N_4686);
nand U5341 (N_5341,N_4643,N_4874);
nor U5342 (N_5342,N_4996,N_4867);
nor U5343 (N_5343,N_4830,N_4799);
or U5344 (N_5344,N_4831,N_4845);
nand U5345 (N_5345,N_4711,N_4773);
nor U5346 (N_5346,N_4697,N_4925);
and U5347 (N_5347,N_4738,N_4616);
nor U5348 (N_5348,N_4676,N_4784);
xnor U5349 (N_5349,N_4669,N_4639);
and U5350 (N_5350,N_4654,N_4546);
nor U5351 (N_5351,N_4945,N_4719);
nand U5352 (N_5352,N_4751,N_4997);
xor U5353 (N_5353,N_4647,N_4877);
xnor U5354 (N_5354,N_4908,N_4941);
or U5355 (N_5355,N_4994,N_4808);
and U5356 (N_5356,N_4735,N_4506);
and U5357 (N_5357,N_4912,N_4872);
nor U5358 (N_5358,N_4776,N_4847);
nand U5359 (N_5359,N_4637,N_4821);
nand U5360 (N_5360,N_4734,N_4680);
nand U5361 (N_5361,N_4509,N_4732);
nor U5362 (N_5362,N_4613,N_4892);
nand U5363 (N_5363,N_4864,N_4890);
and U5364 (N_5364,N_4777,N_4703);
and U5365 (N_5365,N_4982,N_4864);
or U5366 (N_5366,N_4513,N_4694);
xnor U5367 (N_5367,N_4983,N_4648);
and U5368 (N_5368,N_4994,N_4715);
nand U5369 (N_5369,N_4852,N_4530);
or U5370 (N_5370,N_4506,N_4997);
and U5371 (N_5371,N_4576,N_4949);
nor U5372 (N_5372,N_4819,N_4848);
nand U5373 (N_5373,N_4955,N_4927);
and U5374 (N_5374,N_4928,N_4503);
nor U5375 (N_5375,N_4773,N_4971);
nand U5376 (N_5376,N_4630,N_4567);
nand U5377 (N_5377,N_4846,N_4937);
or U5378 (N_5378,N_4899,N_4757);
nand U5379 (N_5379,N_4883,N_4582);
or U5380 (N_5380,N_4932,N_4901);
nand U5381 (N_5381,N_4807,N_4979);
and U5382 (N_5382,N_4538,N_4844);
and U5383 (N_5383,N_4774,N_4688);
or U5384 (N_5384,N_4573,N_4700);
or U5385 (N_5385,N_4749,N_4650);
and U5386 (N_5386,N_4901,N_4761);
and U5387 (N_5387,N_4965,N_4852);
or U5388 (N_5388,N_4889,N_4883);
or U5389 (N_5389,N_4887,N_4866);
nand U5390 (N_5390,N_4502,N_4955);
or U5391 (N_5391,N_4659,N_4705);
or U5392 (N_5392,N_4504,N_4505);
and U5393 (N_5393,N_4542,N_4932);
or U5394 (N_5394,N_4856,N_4780);
or U5395 (N_5395,N_4665,N_4620);
nor U5396 (N_5396,N_4825,N_4528);
and U5397 (N_5397,N_4890,N_4827);
nand U5398 (N_5398,N_4535,N_4558);
nand U5399 (N_5399,N_4805,N_4994);
and U5400 (N_5400,N_4766,N_4850);
or U5401 (N_5401,N_4903,N_4955);
xnor U5402 (N_5402,N_4673,N_4680);
nand U5403 (N_5403,N_4864,N_4730);
nor U5404 (N_5404,N_4718,N_4867);
and U5405 (N_5405,N_4607,N_4844);
or U5406 (N_5406,N_4589,N_4814);
nand U5407 (N_5407,N_4746,N_4820);
or U5408 (N_5408,N_4969,N_4999);
and U5409 (N_5409,N_4833,N_4705);
nor U5410 (N_5410,N_4604,N_4961);
nand U5411 (N_5411,N_4614,N_4522);
and U5412 (N_5412,N_4615,N_4583);
or U5413 (N_5413,N_4706,N_4728);
or U5414 (N_5414,N_4939,N_4969);
nand U5415 (N_5415,N_4612,N_4917);
nor U5416 (N_5416,N_4931,N_4787);
or U5417 (N_5417,N_4869,N_4825);
nor U5418 (N_5418,N_4946,N_4630);
nor U5419 (N_5419,N_4592,N_4824);
xnor U5420 (N_5420,N_4983,N_4729);
or U5421 (N_5421,N_4856,N_4764);
xor U5422 (N_5422,N_4717,N_4603);
or U5423 (N_5423,N_4609,N_4535);
nor U5424 (N_5424,N_4697,N_4712);
nand U5425 (N_5425,N_4770,N_4968);
nand U5426 (N_5426,N_4632,N_4980);
and U5427 (N_5427,N_4984,N_4777);
and U5428 (N_5428,N_4800,N_4683);
nor U5429 (N_5429,N_4518,N_4593);
or U5430 (N_5430,N_4537,N_4973);
and U5431 (N_5431,N_4597,N_4909);
nor U5432 (N_5432,N_4653,N_4627);
or U5433 (N_5433,N_4742,N_4773);
nor U5434 (N_5434,N_4766,N_4546);
nor U5435 (N_5435,N_4874,N_4554);
or U5436 (N_5436,N_4822,N_4760);
or U5437 (N_5437,N_4778,N_4868);
nand U5438 (N_5438,N_4681,N_4857);
and U5439 (N_5439,N_4711,N_4600);
nand U5440 (N_5440,N_4815,N_4505);
nor U5441 (N_5441,N_4566,N_4773);
nor U5442 (N_5442,N_4605,N_4618);
nor U5443 (N_5443,N_4707,N_4716);
nand U5444 (N_5444,N_4568,N_4967);
or U5445 (N_5445,N_4967,N_4666);
or U5446 (N_5446,N_4585,N_4993);
nand U5447 (N_5447,N_4567,N_4818);
nor U5448 (N_5448,N_4937,N_4581);
or U5449 (N_5449,N_4592,N_4953);
or U5450 (N_5450,N_4748,N_4717);
or U5451 (N_5451,N_4646,N_4519);
and U5452 (N_5452,N_4717,N_4905);
nand U5453 (N_5453,N_4523,N_4593);
or U5454 (N_5454,N_4527,N_4950);
or U5455 (N_5455,N_4802,N_4960);
and U5456 (N_5456,N_4925,N_4660);
xor U5457 (N_5457,N_4771,N_4609);
and U5458 (N_5458,N_4926,N_4832);
nor U5459 (N_5459,N_4753,N_4507);
and U5460 (N_5460,N_4716,N_4508);
or U5461 (N_5461,N_4749,N_4745);
nor U5462 (N_5462,N_4786,N_4822);
nor U5463 (N_5463,N_4715,N_4780);
or U5464 (N_5464,N_4911,N_4960);
or U5465 (N_5465,N_4626,N_4686);
xnor U5466 (N_5466,N_4990,N_4611);
or U5467 (N_5467,N_4675,N_4736);
or U5468 (N_5468,N_4757,N_4948);
or U5469 (N_5469,N_4546,N_4524);
nand U5470 (N_5470,N_4947,N_4720);
or U5471 (N_5471,N_4521,N_4913);
and U5472 (N_5472,N_4761,N_4540);
xor U5473 (N_5473,N_4797,N_4636);
and U5474 (N_5474,N_4822,N_4646);
nand U5475 (N_5475,N_4860,N_4807);
and U5476 (N_5476,N_4982,N_4692);
xor U5477 (N_5477,N_4836,N_4590);
nand U5478 (N_5478,N_4525,N_4659);
nor U5479 (N_5479,N_4508,N_4544);
nor U5480 (N_5480,N_4977,N_4945);
xor U5481 (N_5481,N_4569,N_4861);
nand U5482 (N_5482,N_4711,N_4784);
nand U5483 (N_5483,N_4705,N_4764);
or U5484 (N_5484,N_4627,N_4564);
or U5485 (N_5485,N_4889,N_4799);
and U5486 (N_5486,N_4729,N_4706);
nand U5487 (N_5487,N_4851,N_4612);
nand U5488 (N_5488,N_4769,N_4580);
nor U5489 (N_5489,N_4761,N_4651);
and U5490 (N_5490,N_4854,N_4612);
and U5491 (N_5491,N_4789,N_4696);
and U5492 (N_5492,N_4738,N_4534);
and U5493 (N_5493,N_4895,N_4542);
nor U5494 (N_5494,N_4517,N_4966);
nand U5495 (N_5495,N_4978,N_4919);
or U5496 (N_5496,N_4545,N_4758);
nor U5497 (N_5497,N_4866,N_4709);
nand U5498 (N_5498,N_4648,N_4504);
nand U5499 (N_5499,N_4806,N_4636);
nand U5500 (N_5500,N_5494,N_5300);
nand U5501 (N_5501,N_5089,N_5396);
or U5502 (N_5502,N_5073,N_5111);
and U5503 (N_5503,N_5035,N_5127);
and U5504 (N_5504,N_5098,N_5250);
nand U5505 (N_5505,N_5329,N_5397);
nor U5506 (N_5506,N_5371,N_5227);
nand U5507 (N_5507,N_5448,N_5225);
and U5508 (N_5508,N_5465,N_5357);
nand U5509 (N_5509,N_5125,N_5049);
xnor U5510 (N_5510,N_5251,N_5200);
and U5511 (N_5511,N_5462,N_5118);
or U5512 (N_5512,N_5279,N_5048);
nand U5513 (N_5513,N_5129,N_5176);
nor U5514 (N_5514,N_5420,N_5038);
nand U5515 (N_5515,N_5087,N_5156);
nor U5516 (N_5516,N_5275,N_5350);
nand U5517 (N_5517,N_5419,N_5495);
nand U5518 (N_5518,N_5015,N_5395);
xnor U5519 (N_5519,N_5179,N_5009);
or U5520 (N_5520,N_5075,N_5328);
xor U5521 (N_5521,N_5292,N_5005);
nand U5522 (N_5522,N_5139,N_5444);
and U5523 (N_5523,N_5276,N_5284);
xnor U5524 (N_5524,N_5099,N_5491);
or U5525 (N_5525,N_5457,N_5233);
and U5526 (N_5526,N_5271,N_5240);
and U5527 (N_5527,N_5499,N_5234);
nand U5528 (N_5528,N_5166,N_5126);
nor U5529 (N_5529,N_5394,N_5070);
nor U5530 (N_5530,N_5282,N_5363);
nand U5531 (N_5531,N_5223,N_5301);
or U5532 (N_5532,N_5025,N_5412);
or U5533 (N_5533,N_5431,N_5418);
nor U5534 (N_5534,N_5193,N_5290);
or U5535 (N_5535,N_5124,N_5201);
and U5536 (N_5536,N_5402,N_5304);
nand U5537 (N_5537,N_5196,N_5154);
and U5538 (N_5538,N_5265,N_5416);
and U5539 (N_5539,N_5135,N_5027);
xor U5540 (N_5540,N_5340,N_5051);
or U5541 (N_5541,N_5204,N_5105);
nor U5542 (N_5542,N_5298,N_5352);
nor U5543 (N_5543,N_5041,N_5345);
nand U5544 (N_5544,N_5059,N_5224);
nor U5545 (N_5545,N_5381,N_5342);
nand U5546 (N_5546,N_5390,N_5080);
or U5547 (N_5547,N_5237,N_5114);
and U5548 (N_5548,N_5456,N_5222);
and U5549 (N_5549,N_5113,N_5370);
or U5550 (N_5550,N_5461,N_5014);
nor U5551 (N_5551,N_5386,N_5071);
nor U5552 (N_5552,N_5407,N_5299);
xnor U5553 (N_5553,N_5187,N_5497);
or U5554 (N_5554,N_5410,N_5198);
nor U5555 (N_5555,N_5106,N_5205);
nand U5556 (N_5556,N_5472,N_5044);
nand U5557 (N_5557,N_5325,N_5092);
nor U5558 (N_5558,N_5459,N_5335);
nor U5559 (N_5559,N_5393,N_5324);
or U5560 (N_5560,N_5177,N_5373);
or U5561 (N_5561,N_5375,N_5440);
nand U5562 (N_5562,N_5278,N_5449);
nor U5563 (N_5563,N_5191,N_5389);
and U5564 (N_5564,N_5084,N_5319);
nand U5565 (N_5565,N_5110,N_5042);
xnor U5566 (N_5566,N_5426,N_5141);
nor U5567 (N_5567,N_5120,N_5088);
nand U5568 (N_5568,N_5483,N_5151);
and U5569 (N_5569,N_5019,N_5391);
nand U5570 (N_5570,N_5050,N_5182);
and U5571 (N_5571,N_5189,N_5377);
nand U5572 (N_5572,N_5045,N_5405);
nor U5573 (N_5573,N_5326,N_5441);
nor U5574 (N_5574,N_5257,N_5010);
nand U5575 (N_5575,N_5002,N_5433);
nor U5576 (N_5576,N_5327,N_5453);
nand U5577 (N_5577,N_5437,N_5309);
or U5578 (N_5578,N_5122,N_5012);
or U5579 (N_5579,N_5445,N_5195);
nand U5580 (N_5580,N_5085,N_5323);
or U5581 (N_5581,N_5142,N_5039);
nand U5582 (N_5582,N_5033,N_5277);
nand U5583 (N_5583,N_5003,N_5213);
nor U5584 (N_5584,N_5097,N_5210);
nor U5585 (N_5585,N_5493,N_5221);
or U5586 (N_5586,N_5314,N_5214);
nand U5587 (N_5587,N_5403,N_5374);
nor U5588 (N_5588,N_5115,N_5052);
and U5589 (N_5589,N_5147,N_5174);
nand U5590 (N_5590,N_5330,N_5435);
or U5591 (N_5591,N_5281,N_5194);
and U5592 (N_5592,N_5024,N_5358);
and U5593 (N_5593,N_5253,N_5215);
xnor U5594 (N_5594,N_5066,N_5447);
and U5595 (N_5595,N_5181,N_5392);
nor U5596 (N_5596,N_5285,N_5199);
nor U5597 (N_5597,N_5261,N_5414);
nor U5598 (N_5598,N_5256,N_5243);
and U5599 (N_5599,N_5354,N_5337);
xor U5600 (N_5600,N_5159,N_5294);
and U5601 (N_5601,N_5482,N_5490);
nand U5602 (N_5602,N_5272,N_5220);
and U5603 (N_5603,N_5007,N_5077);
and U5604 (N_5604,N_5247,N_5452);
nor U5605 (N_5605,N_5262,N_5400);
or U5606 (N_5606,N_5180,N_5242);
xor U5607 (N_5607,N_5362,N_5208);
nor U5608 (N_5608,N_5169,N_5442);
and U5609 (N_5609,N_5083,N_5158);
or U5610 (N_5610,N_5455,N_5434);
xor U5611 (N_5611,N_5026,N_5339);
or U5612 (N_5612,N_5382,N_5479);
nand U5613 (N_5613,N_5288,N_5104);
nor U5614 (N_5614,N_5460,N_5076);
nand U5615 (N_5615,N_5239,N_5331);
nand U5616 (N_5616,N_5361,N_5047);
and U5617 (N_5617,N_5086,N_5018);
nor U5618 (N_5618,N_5353,N_5178);
or U5619 (N_5619,N_5054,N_5093);
nand U5620 (N_5620,N_5226,N_5119);
or U5621 (N_5621,N_5101,N_5424);
nand U5622 (N_5622,N_5259,N_5476);
nand U5623 (N_5623,N_5032,N_5082);
nor U5624 (N_5624,N_5157,N_5100);
and U5625 (N_5625,N_5470,N_5450);
or U5626 (N_5626,N_5167,N_5152);
or U5627 (N_5627,N_5149,N_5322);
and U5628 (N_5628,N_5303,N_5245);
or U5629 (N_5629,N_5417,N_5367);
nor U5630 (N_5630,N_5332,N_5372);
xor U5631 (N_5631,N_5409,N_5020);
nor U5632 (N_5632,N_5171,N_5030);
nor U5633 (N_5633,N_5072,N_5146);
nand U5634 (N_5634,N_5004,N_5343);
nand U5635 (N_5635,N_5384,N_5108);
nor U5636 (N_5636,N_5474,N_5466);
nor U5637 (N_5637,N_5415,N_5219);
and U5638 (N_5638,N_5286,N_5197);
nand U5639 (N_5639,N_5287,N_5173);
nor U5640 (N_5640,N_5065,N_5378);
or U5641 (N_5641,N_5023,N_5074);
or U5642 (N_5642,N_5385,N_5321);
or U5643 (N_5643,N_5090,N_5091);
and U5644 (N_5644,N_5063,N_5346);
and U5645 (N_5645,N_5136,N_5383);
and U5646 (N_5646,N_5175,N_5218);
and U5647 (N_5647,N_5376,N_5280);
nand U5648 (N_5648,N_5464,N_5308);
and U5649 (N_5649,N_5170,N_5238);
xor U5650 (N_5650,N_5318,N_5305);
nand U5651 (N_5651,N_5430,N_5246);
nand U5652 (N_5652,N_5439,N_5011);
nor U5653 (N_5653,N_5478,N_5487);
or U5654 (N_5654,N_5366,N_5388);
or U5655 (N_5655,N_5469,N_5116);
nor U5656 (N_5656,N_5429,N_5477);
nand U5657 (N_5657,N_5061,N_5310);
nor U5658 (N_5658,N_5260,N_5001);
and U5659 (N_5659,N_5069,N_5132);
nor U5660 (N_5660,N_5150,N_5338);
nand U5661 (N_5661,N_5244,N_5291);
nand U5662 (N_5662,N_5209,N_5404);
nor U5663 (N_5663,N_5013,N_5046);
nor U5664 (N_5664,N_5312,N_5236);
and U5665 (N_5665,N_5496,N_5203);
nand U5666 (N_5666,N_5060,N_5094);
and U5667 (N_5667,N_5427,N_5359);
nor U5668 (N_5668,N_5317,N_5143);
xor U5669 (N_5669,N_5036,N_5188);
nand U5670 (N_5670,N_5422,N_5344);
and U5671 (N_5671,N_5006,N_5398);
nor U5672 (N_5672,N_5095,N_5163);
xnor U5673 (N_5673,N_5000,N_5207);
nand U5674 (N_5674,N_5216,N_5438);
and U5675 (N_5675,N_5485,N_5081);
nand U5676 (N_5676,N_5349,N_5168);
nor U5677 (N_5677,N_5421,N_5316);
and U5678 (N_5678,N_5133,N_5137);
and U5679 (N_5679,N_5096,N_5406);
and U5680 (N_5680,N_5123,N_5131);
nand U5681 (N_5681,N_5432,N_5162);
or U5682 (N_5682,N_5117,N_5172);
nand U5683 (N_5683,N_5369,N_5252);
nor U5684 (N_5684,N_5164,N_5356);
nor U5685 (N_5685,N_5365,N_5103);
nand U5686 (N_5686,N_5212,N_5190);
and U5687 (N_5687,N_5034,N_5368);
and U5688 (N_5688,N_5183,N_5128);
nor U5689 (N_5689,N_5267,N_5380);
xnor U5690 (N_5690,N_5056,N_5028);
or U5691 (N_5691,N_5296,N_5295);
xor U5692 (N_5692,N_5347,N_5401);
xnor U5693 (N_5693,N_5231,N_5241);
nand U5694 (N_5694,N_5232,N_5109);
xnor U5695 (N_5695,N_5017,N_5315);
and U5696 (N_5696,N_5008,N_5307);
nand U5697 (N_5697,N_5270,N_5079);
or U5698 (N_5698,N_5064,N_5254);
xnor U5699 (N_5699,N_5264,N_5269);
nor U5700 (N_5700,N_5186,N_5107);
nand U5701 (N_5701,N_5217,N_5387);
nor U5702 (N_5702,N_5228,N_5475);
nor U5703 (N_5703,N_5436,N_5202);
nand U5704 (N_5704,N_5153,N_5473);
and U5705 (N_5705,N_5229,N_5140);
and U5706 (N_5706,N_5443,N_5302);
nor U5707 (N_5707,N_5184,N_5454);
and U5708 (N_5708,N_5311,N_5306);
and U5709 (N_5709,N_5230,N_5058);
or U5710 (N_5710,N_5492,N_5399);
nor U5711 (N_5711,N_5165,N_5145);
nor U5712 (N_5712,N_5211,N_5078);
nor U5713 (N_5713,N_5185,N_5021);
and U5714 (N_5714,N_5258,N_5206);
nor U5715 (N_5715,N_5121,N_5268);
or U5716 (N_5716,N_5425,N_5022);
or U5717 (N_5717,N_5468,N_5334);
nor U5718 (N_5718,N_5263,N_5486);
nand U5719 (N_5719,N_5320,N_5289);
nand U5720 (N_5720,N_5266,N_5488);
nand U5721 (N_5721,N_5471,N_5255);
or U5722 (N_5722,N_5102,N_5248);
nand U5723 (N_5723,N_5355,N_5160);
and U5724 (N_5724,N_5379,N_5413);
nor U5725 (N_5725,N_5458,N_5283);
nor U5726 (N_5726,N_5293,N_5463);
nor U5727 (N_5727,N_5037,N_5040);
nor U5728 (N_5728,N_5446,N_5484);
nand U5729 (N_5729,N_5451,N_5031);
nand U5730 (N_5730,N_5341,N_5411);
and U5731 (N_5731,N_5364,N_5144);
or U5732 (N_5732,N_5274,N_5235);
or U5733 (N_5733,N_5130,N_5297);
and U5734 (N_5734,N_5062,N_5467);
and U5735 (N_5735,N_5161,N_5481);
nor U5736 (N_5736,N_5053,N_5192);
and U5737 (N_5737,N_5360,N_5351);
or U5738 (N_5738,N_5155,N_5067);
and U5739 (N_5739,N_5498,N_5423);
nand U5740 (N_5740,N_5336,N_5057);
xnor U5741 (N_5741,N_5273,N_5068);
nand U5742 (N_5742,N_5428,N_5148);
or U5743 (N_5743,N_5333,N_5055);
nand U5744 (N_5744,N_5480,N_5138);
nand U5745 (N_5745,N_5489,N_5134);
nand U5746 (N_5746,N_5348,N_5408);
nand U5747 (N_5747,N_5016,N_5313);
and U5748 (N_5748,N_5043,N_5249);
and U5749 (N_5749,N_5112,N_5029);
or U5750 (N_5750,N_5191,N_5085);
and U5751 (N_5751,N_5209,N_5405);
or U5752 (N_5752,N_5047,N_5271);
xor U5753 (N_5753,N_5239,N_5063);
or U5754 (N_5754,N_5091,N_5383);
or U5755 (N_5755,N_5431,N_5074);
nor U5756 (N_5756,N_5454,N_5254);
or U5757 (N_5757,N_5298,N_5336);
or U5758 (N_5758,N_5183,N_5489);
and U5759 (N_5759,N_5169,N_5302);
nand U5760 (N_5760,N_5266,N_5190);
nor U5761 (N_5761,N_5173,N_5283);
and U5762 (N_5762,N_5482,N_5013);
and U5763 (N_5763,N_5439,N_5197);
or U5764 (N_5764,N_5092,N_5020);
and U5765 (N_5765,N_5470,N_5321);
or U5766 (N_5766,N_5331,N_5129);
nor U5767 (N_5767,N_5196,N_5015);
or U5768 (N_5768,N_5009,N_5250);
nor U5769 (N_5769,N_5061,N_5035);
xor U5770 (N_5770,N_5439,N_5164);
xor U5771 (N_5771,N_5319,N_5088);
xnor U5772 (N_5772,N_5448,N_5056);
nand U5773 (N_5773,N_5297,N_5083);
and U5774 (N_5774,N_5346,N_5074);
nand U5775 (N_5775,N_5450,N_5495);
xnor U5776 (N_5776,N_5094,N_5259);
nor U5777 (N_5777,N_5219,N_5476);
nand U5778 (N_5778,N_5289,N_5414);
and U5779 (N_5779,N_5384,N_5430);
nor U5780 (N_5780,N_5141,N_5174);
nand U5781 (N_5781,N_5309,N_5264);
nor U5782 (N_5782,N_5405,N_5421);
or U5783 (N_5783,N_5241,N_5384);
nand U5784 (N_5784,N_5222,N_5497);
or U5785 (N_5785,N_5178,N_5124);
nand U5786 (N_5786,N_5109,N_5258);
xnor U5787 (N_5787,N_5243,N_5177);
nor U5788 (N_5788,N_5096,N_5364);
nor U5789 (N_5789,N_5325,N_5111);
and U5790 (N_5790,N_5480,N_5200);
xor U5791 (N_5791,N_5263,N_5007);
nand U5792 (N_5792,N_5195,N_5155);
or U5793 (N_5793,N_5454,N_5224);
or U5794 (N_5794,N_5297,N_5344);
nor U5795 (N_5795,N_5127,N_5147);
nand U5796 (N_5796,N_5088,N_5483);
or U5797 (N_5797,N_5119,N_5017);
nor U5798 (N_5798,N_5250,N_5126);
nand U5799 (N_5799,N_5117,N_5192);
nand U5800 (N_5800,N_5273,N_5427);
nor U5801 (N_5801,N_5144,N_5081);
and U5802 (N_5802,N_5157,N_5405);
xnor U5803 (N_5803,N_5318,N_5077);
and U5804 (N_5804,N_5416,N_5120);
or U5805 (N_5805,N_5060,N_5068);
nor U5806 (N_5806,N_5423,N_5246);
and U5807 (N_5807,N_5155,N_5132);
nand U5808 (N_5808,N_5076,N_5417);
nor U5809 (N_5809,N_5351,N_5434);
nor U5810 (N_5810,N_5375,N_5035);
nor U5811 (N_5811,N_5256,N_5239);
nand U5812 (N_5812,N_5229,N_5317);
or U5813 (N_5813,N_5129,N_5207);
or U5814 (N_5814,N_5053,N_5309);
or U5815 (N_5815,N_5056,N_5266);
nand U5816 (N_5816,N_5266,N_5086);
nand U5817 (N_5817,N_5042,N_5024);
nand U5818 (N_5818,N_5136,N_5177);
and U5819 (N_5819,N_5315,N_5166);
nor U5820 (N_5820,N_5422,N_5481);
nand U5821 (N_5821,N_5017,N_5293);
xnor U5822 (N_5822,N_5461,N_5085);
nor U5823 (N_5823,N_5435,N_5391);
or U5824 (N_5824,N_5422,N_5455);
and U5825 (N_5825,N_5173,N_5479);
nor U5826 (N_5826,N_5408,N_5398);
nor U5827 (N_5827,N_5302,N_5126);
or U5828 (N_5828,N_5079,N_5131);
nor U5829 (N_5829,N_5476,N_5068);
and U5830 (N_5830,N_5356,N_5348);
xor U5831 (N_5831,N_5398,N_5334);
and U5832 (N_5832,N_5043,N_5190);
nand U5833 (N_5833,N_5249,N_5051);
nor U5834 (N_5834,N_5236,N_5321);
nor U5835 (N_5835,N_5293,N_5220);
nor U5836 (N_5836,N_5005,N_5138);
or U5837 (N_5837,N_5114,N_5324);
and U5838 (N_5838,N_5383,N_5462);
nor U5839 (N_5839,N_5337,N_5024);
and U5840 (N_5840,N_5016,N_5426);
nor U5841 (N_5841,N_5149,N_5481);
nor U5842 (N_5842,N_5130,N_5057);
and U5843 (N_5843,N_5472,N_5128);
or U5844 (N_5844,N_5455,N_5281);
nor U5845 (N_5845,N_5158,N_5106);
and U5846 (N_5846,N_5236,N_5395);
xnor U5847 (N_5847,N_5219,N_5373);
nor U5848 (N_5848,N_5270,N_5471);
nor U5849 (N_5849,N_5176,N_5174);
nand U5850 (N_5850,N_5381,N_5191);
and U5851 (N_5851,N_5429,N_5260);
nor U5852 (N_5852,N_5381,N_5483);
nor U5853 (N_5853,N_5357,N_5059);
and U5854 (N_5854,N_5112,N_5470);
xor U5855 (N_5855,N_5280,N_5475);
or U5856 (N_5856,N_5466,N_5372);
nor U5857 (N_5857,N_5366,N_5423);
or U5858 (N_5858,N_5375,N_5081);
and U5859 (N_5859,N_5229,N_5032);
nor U5860 (N_5860,N_5108,N_5131);
xor U5861 (N_5861,N_5210,N_5199);
nor U5862 (N_5862,N_5068,N_5247);
or U5863 (N_5863,N_5266,N_5412);
nand U5864 (N_5864,N_5142,N_5029);
nand U5865 (N_5865,N_5006,N_5058);
and U5866 (N_5866,N_5130,N_5058);
and U5867 (N_5867,N_5106,N_5108);
nor U5868 (N_5868,N_5330,N_5250);
or U5869 (N_5869,N_5212,N_5263);
or U5870 (N_5870,N_5258,N_5448);
or U5871 (N_5871,N_5220,N_5339);
xnor U5872 (N_5872,N_5405,N_5267);
nor U5873 (N_5873,N_5402,N_5199);
nor U5874 (N_5874,N_5195,N_5036);
or U5875 (N_5875,N_5368,N_5443);
or U5876 (N_5876,N_5276,N_5175);
nor U5877 (N_5877,N_5306,N_5408);
xor U5878 (N_5878,N_5432,N_5342);
and U5879 (N_5879,N_5425,N_5301);
nand U5880 (N_5880,N_5350,N_5120);
nor U5881 (N_5881,N_5294,N_5428);
nor U5882 (N_5882,N_5172,N_5258);
nor U5883 (N_5883,N_5094,N_5240);
or U5884 (N_5884,N_5208,N_5256);
or U5885 (N_5885,N_5244,N_5050);
or U5886 (N_5886,N_5161,N_5170);
nor U5887 (N_5887,N_5373,N_5060);
xor U5888 (N_5888,N_5234,N_5186);
and U5889 (N_5889,N_5160,N_5310);
and U5890 (N_5890,N_5407,N_5318);
nand U5891 (N_5891,N_5491,N_5342);
and U5892 (N_5892,N_5083,N_5169);
and U5893 (N_5893,N_5062,N_5274);
nand U5894 (N_5894,N_5106,N_5328);
nor U5895 (N_5895,N_5057,N_5357);
or U5896 (N_5896,N_5120,N_5243);
xor U5897 (N_5897,N_5245,N_5456);
nor U5898 (N_5898,N_5433,N_5208);
nor U5899 (N_5899,N_5158,N_5010);
nand U5900 (N_5900,N_5153,N_5359);
nor U5901 (N_5901,N_5405,N_5413);
nand U5902 (N_5902,N_5006,N_5280);
nand U5903 (N_5903,N_5127,N_5157);
nor U5904 (N_5904,N_5138,N_5422);
or U5905 (N_5905,N_5318,N_5376);
and U5906 (N_5906,N_5124,N_5343);
or U5907 (N_5907,N_5023,N_5044);
xor U5908 (N_5908,N_5204,N_5091);
nand U5909 (N_5909,N_5165,N_5094);
xnor U5910 (N_5910,N_5134,N_5364);
or U5911 (N_5911,N_5334,N_5167);
nand U5912 (N_5912,N_5105,N_5323);
or U5913 (N_5913,N_5188,N_5003);
and U5914 (N_5914,N_5314,N_5433);
and U5915 (N_5915,N_5064,N_5473);
nand U5916 (N_5916,N_5011,N_5371);
or U5917 (N_5917,N_5413,N_5376);
nand U5918 (N_5918,N_5499,N_5160);
or U5919 (N_5919,N_5214,N_5305);
nand U5920 (N_5920,N_5190,N_5173);
xor U5921 (N_5921,N_5069,N_5264);
and U5922 (N_5922,N_5451,N_5225);
nor U5923 (N_5923,N_5476,N_5080);
and U5924 (N_5924,N_5475,N_5247);
nand U5925 (N_5925,N_5271,N_5408);
xnor U5926 (N_5926,N_5113,N_5366);
and U5927 (N_5927,N_5490,N_5252);
nand U5928 (N_5928,N_5105,N_5220);
nor U5929 (N_5929,N_5085,N_5429);
or U5930 (N_5930,N_5445,N_5134);
or U5931 (N_5931,N_5461,N_5120);
nand U5932 (N_5932,N_5216,N_5046);
or U5933 (N_5933,N_5454,N_5011);
or U5934 (N_5934,N_5282,N_5093);
or U5935 (N_5935,N_5086,N_5216);
xnor U5936 (N_5936,N_5243,N_5137);
or U5937 (N_5937,N_5275,N_5027);
and U5938 (N_5938,N_5137,N_5336);
and U5939 (N_5939,N_5049,N_5253);
and U5940 (N_5940,N_5412,N_5422);
xor U5941 (N_5941,N_5484,N_5121);
or U5942 (N_5942,N_5007,N_5288);
or U5943 (N_5943,N_5290,N_5160);
nand U5944 (N_5944,N_5297,N_5336);
and U5945 (N_5945,N_5471,N_5345);
nor U5946 (N_5946,N_5076,N_5316);
and U5947 (N_5947,N_5274,N_5482);
nor U5948 (N_5948,N_5325,N_5362);
or U5949 (N_5949,N_5123,N_5174);
or U5950 (N_5950,N_5454,N_5421);
and U5951 (N_5951,N_5367,N_5220);
nand U5952 (N_5952,N_5493,N_5429);
nor U5953 (N_5953,N_5456,N_5335);
nor U5954 (N_5954,N_5161,N_5085);
xnor U5955 (N_5955,N_5221,N_5498);
nand U5956 (N_5956,N_5151,N_5439);
nand U5957 (N_5957,N_5431,N_5292);
and U5958 (N_5958,N_5166,N_5254);
nand U5959 (N_5959,N_5375,N_5012);
nand U5960 (N_5960,N_5365,N_5472);
or U5961 (N_5961,N_5202,N_5121);
and U5962 (N_5962,N_5057,N_5356);
nor U5963 (N_5963,N_5384,N_5339);
nor U5964 (N_5964,N_5222,N_5340);
nor U5965 (N_5965,N_5395,N_5347);
or U5966 (N_5966,N_5435,N_5216);
nand U5967 (N_5967,N_5116,N_5268);
and U5968 (N_5968,N_5046,N_5107);
nor U5969 (N_5969,N_5098,N_5296);
nor U5970 (N_5970,N_5359,N_5481);
and U5971 (N_5971,N_5156,N_5349);
nor U5972 (N_5972,N_5380,N_5275);
or U5973 (N_5973,N_5113,N_5124);
and U5974 (N_5974,N_5354,N_5013);
and U5975 (N_5975,N_5062,N_5294);
nor U5976 (N_5976,N_5033,N_5238);
nand U5977 (N_5977,N_5321,N_5424);
nand U5978 (N_5978,N_5400,N_5246);
and U5979 (N_5979,N_5233,N_5299);
or U5980 (N_5980,N_5382,N_5286);
or U5981 (N_5981,N_5337,N_5082);
or U5982 (N_5982,N_5458,N_5358);
nand U5983 (N_5983,N_5126,N_5091);
or U5984 (N_5984,N_5443,N_5483);
or U5985 (N_5985,N_5253,N_5199);
or U5986 (N_5986,N_5295,N_5255);
and U5987 (N_5987,N_5318,N_5388);
and U5988 (N_5988,N_5248,N_5448);
and U5989 (N_5989,N_5094,N_5466);
nand U5990 (N_5990,N_5494,N_5215);
nand U5991 (N_5991,N_5316,N_5396);
nor U5992 (N_5992,N_5065,N_5483);
nor U5993 (N_5993,N_5084,N_5392);
nor U5994 (N_5994,N_5271,N_5255);
nor U5995 (N_5995,N_5178,N_5427);
or U5996 (N_5996,N_5409,N_5145);
nand U5997 (N_5997,N_5301,N_5225);
nor U5998 (N_5998,N_5396,N_5047);
and U5999 (N_5999,N_5210,N_5354);
nand U6000 (N_6000,N_5785,N_5698);
and U6001 (N_6001,N_5831,N_5817);
or U6002 (N_6002,N_5684,N_5699);
and U6003 (N_6003,N_5747,N_5982);
nand U6004 (N_6004,N_5595,N_5933);
nor U6005 (N_6005,N_5999,N_5763);
or U6006 (N_6006,N_5525,N_5709);
or U6007 (N_6007,N_5606,N_5591);
xor U6008 (N_6008,N_5618,N_5732);
xnor U6009 (N_6009,N_5562,N_5760);
nor U6010 (N_6010,N_5917,N_5737);
or U6011 (N_6011,N_5821,N_5717);
xnor U6012 (N_6012,N_5617,N_5846);
and U6013 (N_6013,N_5911,N_5955);
xnor U6014 (N_6014,N_5786,N_5539);
nand U6015 (N_6015,N_5956,N_5788);
or U6016 (N_6016,N_5688,N_5839);
and U6017 (N_6017,N_5513,N_5742);
nand U6018 (N_6018,N_5567,N_5870);
and U6019 (N_6019,N_5653,N_5694);
and U6020 (N_6020,N_5655,N_5540);
and U6021 (N_6021,N_5638,N_5945);
or U6022 (N_6022,N_5503,N_5892);
and U6023 (N_6023,N_5896,N_5860);
nand U6024 (N_6024,N_5529,N_5865);
and U6025 (N_6025,N_5922,N_5868);
nor U6026 (N_6026,N_5674,N_5599);
or U6027 (N_6027,N_5612,N_5613);
nand U6028 (N_6028,N_5780,N_5822);
xnor U6029 (N_6029,N_5985,N_5629);
nor U6030 (N_6030,N_5931,N_5908);
nand U6031 (N_6031,N_5748,N_5666);
nor U6032 (N_6032,N_5632,N_5576);
and U6033 (N_6033,N_5842,N_5987);
and U6034 (N_6034,N_5628,N_5872);
nor U6035 (N_6035,N_5967,N_5735);
nor U6036 (N_6036,N_5533,N_5824);
nand U6037 (N_6037,N_5965,N_5869);
xnor U6038 (N_6038,N_5871,N_5781);
nand U6039 (N_6039,N_5981,N_5507);
or U6040 (N_6040,N_5670,N_5657);
nand U6041 (N_6041,N_5947,N_5583);
and U6042 (N_6042,N_5608,N_5582);
xnor U6043 (N_6043,N_5844,N_5926);
nor U6044 (N_6044,N_5899,N_5849);
nand U6045 (N_6045,N_5816,N_5969);
xor U6046 (N_6046,N_5512,N_5675);
nand U6047 (N_6047,N_5719,N_5823);
or U6048 (N_6048,N_5704,N_5598);
nor U6049 (N_6049,N_5571,N_5972);
or U6050 (N_6050,N_5601,N_5886);
or U6051 (N_6051,N_5553,N_5827);
and U6052 (N_6052,N_5939,N_5700);
nor U6053 (N_6053,N_5993,N_5500);
nand U6054 (N_6054,N_5641,N_5723);
or U6055 (N_6055,N_5733,N_5703);
and U6056 (N_6056,N_5702,N_5797);
or U6057 (N_6057,N_5843,N_5961);
or U6058 (N_6058,N_5721,N_5537);
nor U6059 (N_6059,N_5555,N_5954);
or U6060 (N_6060,N_5552,N_5928);
or U6061 (N_6061,N_5957,N_5942);
nand U6062 (N_6062,N_5741,N_5861);
nor U6063 (N_6063,N_5751,N_5585);
or U6064 (N_6064,N_5623,N_5835);
xor U6065 (N_6065,N_5782,N_5720);
nand U6066 (N_6066,N_5610,N_5776);
nand U6067 (N_6067,N_5546,N_5715);
and U6068 (N_6068,N_5658,N_5864);
nor U6069 (N_6069,N_5665,N_5647);
nand U6070 (N_6070,N_5521,N_5668);
or U6071 (N_6071,N_5504,N_5907);
or U6072 (N_6072,N_5994,N_5897);
nand U6073 (N_6073,N_5958,N_5596);
nand U6074 (N_6074,N_5758,N_5547);
xor U6075 (N_6075,N_5990,N_5941);
xor U6076 (N_6076,N_5648,N_5976);
or U6077 (N_6077,N_5568,N_5590);
nor U6078 (N_6078,N_5573,N_5832);
nand U6079 (N_6079,N_5974,N_5853);
or U6080 (N_6080,N_5923,N_5882);
nor U6081 (N_6081,N_5646,N_5510);
xor U6082 (N_6082,N_5840,N_5676);
nor U6083 (N_6083,N_5627,N_5905);
nand U6084 (N_6084,N_5811,N_5631);
and U6085 (N_6085,N_5572,N_5960);
nor U6086 (N_6086,N_5910,N_5686);
nor U6087 (N_6087,N_5964,N_5501);
nand U6088 (N_6088,N_5511,N_5790);
and U6089 (N_6089,N_5691,N_5570);
nor U6090 (N_6090,N_5973,N_5649);
nand U6091 (N_6091,N_5837,N_5891);
nor U6092 (N_6092,N_5695,N_5847);
or U6093 (N_6093,N_5693,N_5640);
or U6094 (N_6094,N_5519,N_5789);
or U6095 (N_6095,N_5946,N_5671);
nor U6096 (N_6096,N_5597,N_5626);
nor U6097 (N_6097,N_5575,N_5743);
nand U6098 (N_6098,N_5867,N_5884);
nor U6099 (N_6099,N_5909,N_5902);
nand U6100 (N_6100,N_5997,N_5611);
nand U6101 (N_6101,N_5522,N_5669);
nand U6102 (N_6102,N_5600,N_5808);
nand U6103 (N_6103,N_5978,N_5834);
nand U6104 (N_6104,N_5784,N_5707);
nor U6105 (N_6105,N_5764,N_5722);
and U6106 (N_6106,N_5912,N_5901);
and U6107 (N_6107,N_5765,N_5635);
and U6108 (N_6108,N_5740,N_5662);
nor U6109 (N_6109,N_5651,N_5845);
and U6110 (N_6110,N_5953,N_5746);
nand U6111 (N_6111,N_5589,N_5544);
and U6112 (N_6112,N_5557,N_5794);
and U6113 (N_6113,N_5878,N_5564);
nand U6114 (N_6114,N_5754,N_5616);
nor U6115 (N_6115,N_5850,N_5535);
or U6116 (N_6116,N_5949,N_5929);
nor U6117 (N_6117,N_5932,N_5663);
or U6118 (N_6118,N_5614,N_5710);
nand U6119 (N_6119,N_5783,N_5724);
and U6120 (N_6120,N_5952,N_5545);
xnor U6121 (N_6121,N_5543,N_5636);
nand U6122 (N_6122,N_5855,N_5998);
or U6123 (N_6123,N_5558,N_5654);
or U6124 (N_6124,N_5859,N_5550);
nor U6125 (N_6125,N_5580,N_5975);
nand U6126 (N_6126,N_5678,N_5904);
nand U6127 (N_6127,N_5711,N_5752);
nand U6128 (N_6128,N_5734,N_5986);
or U6129 (N_6129,N_5778,N_5687);
and U6130 (N_6130,N_5992,N_5587);
nor U6131 (N_6131,N_5634,N_5894);
nor U6132 (N_6132,N_5716,N_5561);
and U6133 (N_6133,N_5906,N_5836);
xor U6134 (N_6134,N_5726,N_5615);
nand U6135 (N_6135,N_5875,N_5863);
or U6136 (N_6136,N_5744,N_5542);
or U6137 (N_6137,N_5528,N_5523);
xnor U6138 (N_6138,N_5714,N_5574);
nand U6139 (N_6139,N_5532,N_5996);
or U6140 (N_6140,N_5559,N_5963);
or U6141 (N_6141,N_5983,N_5852);
nor U6142 (N_6142,N_5536,N_5950);
or U6143 (N_6143,N_5738,N_5530);
xnor U6144 (N_6144,N_5795,N_5848);
nand U6145 (N_6145,N_5881,N_5889);
or U6146 (N_6146,N_5692,N_5779);
and U6147 (N_6147,N_5826,N_5727);
or U6148 (N_6148,N_5761,N_5560);
nand U6149 (N_6149,N_5913,N_5898);
nor U6150 (N_6150,N_5793,N_5526);
nand U6151 (N_6151,N_5877,N_5805);
nor U6152 (N_6152,N_5777,N_5527);
or U6153 (N_6153,N_5556,N_5566);
nand U6154 (N_6154,N_5622,N_5851);
or U6155 (N_6155,N_5745,N_5680);
nand U6156 (N_6156,N_5509,N_5773);
nand U6157 (N_6157,N_5885,N_5592);
and U6158 (N_6158,N_5645,N_5919);
or U6159 (N_6159,N_5768,N_5980);
and U6160 (N_6160,N_5605,N_5578);
and U6161 (N_6161,N_5639,N_5565);
nor U6162 (N_6162,N_5739,N_5959);
and U6163 (N_6163,N_5804,N_5991);
or U6164 (N_6164,N_5633,N_5594);
or U6165 (N_6165,N_5725,N_5841);
or U6166 (N_6166,N_5730,N_5798);
nand U6167 (N_6167,N_5799,N_5607);
nand U6168 (N_6168,N_5825,N_5979);
nand U6169 (N_6169,N_5637,N_5903);
nor U6170 (N_6170,N_5652,N_5938);
or U6171 (N_6171,N_5809,N_5642);
and U6172 (N_6172,N_5619,N_5951);
nand U6173 (N_6173,N_5829,N_5602);
and U6174 (N_6174,N_5820,N_5551);
or U6175 (N_6175,N_5879,N_5866);
and U6176 (N_6176,N_5888,N_5672);
and U6177 (N_6177,N_5854,N_5681);
xnor U6178 (N_6178,N_5689,N_5772);
nor U6179 (N_6179,N_5630,N_5792);
or U6180 (N_6180,N_5505,N_5940);
or U6181 (N_6181,N_5900,N_5696);
and U6182 (N_6182,N_5660,N_5819);
nand U6183 (N_6183,N_5531,N_5995);
or U6184 (N_6184,N_5769,N_5577);
and U6185 (N_6185,N_5818,N_5643);
xor U6186 (N_6186,N_5927,N_5971);
and U6187 (N_6187,N_5718,N_5857);
nand U6188 (N_6188,N_5858,N_5815);
and U6189 (N_6189,N_5581,N_5549);
nand U6190 (N_6190,N_5729,N_5810);
or U6191 (N_6191,N_5802,N_5563);
or U6192 (N_6192,N_5524,N_5988);
and U6193 (N_6193,N_5918,N_5862);
nor U6194 (N_6194,N_5874,N_5921);
nand U6195 (N_6195,N_5948,N_5893);
nor U6196 (N_6196,N_5708,N_5593);
nor U6197 (N_6197,N_5873,N_5621);
and U6198 (N_6198,N_5548,N_5506);
nand U6199 (N_6199,N_5673,N_5520);
nor U6200 (N_6200,N_5771,N_5759);
nand U6201 (N_6201,N_5838,N_5713);
xnor U6202 (N_6202,N_5977,N_5604);
nor U6203 (N_6203,N_5880,N_5516);
and U6204 (N_6204,N_5683,N_5968);
and U6205 (N_6205,N_5930,N_5728);
nand U6206 (N_6206,N_5753,N_5685);
xor U6207 (N_6207,N_5609,N_5706);
or U6208 (N_6208,N_5554,N_5937);
nor U6209 (N_6209,N_5661,N_5603);
nor U6210 (N_6210,N_5925,N_5762);
nand U6211 (N_6211,N_5755,N_5944);
nand U6212 (N_6212,N_5833,N_5518);
and U6213 (N_6213,N_5749,N_5812);
nor U6214 (N_6214,N_5962,N_5806);
xor U6215 (N_6215,N_5801,N_5656);
xor U6216 (N_6216,N_5796,N_5514);
nor U6217 (N_6217,N_5775,N_5701);
and U6218 (N_6218,N_5766,N_5924);
xor U6219 (N_6219,N_5787,N_5731);
or U6220 (N_6220,N_5807,N_5620);
nor U6221 (N_6221,N_5830,N_5586);
and U6222 (N_6222,N_5679,N_5757);
and U6223 (N_6223,N_5814,N_5736);
xor U6224 (N_6224,N_5502,N_5916);
or U6225 (N_6225,N_5774,N_5677);
xnor U6226 (N_6226,N_5659,N_5883);
or U6227 (N_6227,N_5828,N_5895);
or U6228 (N_6228,N_5579,N_5966);
or U6229 (N_6229,N_5690,N_5541);
and U6230 (N_6230,N_5705,N_5970);
nor U6231 (N_6231,N_5989,N_5920);
nor U6232 (N_6232,N_5943,N_5650);
nor U6233 (N_6233,N_5569,N_5813);
xnor U6234 (N_6234,N_5750,N_5682);
nor U6235 (N_6235,N_5664,N_5697);
or U6236 (N_6236,N_5876,N_5667);
or U6237 (N_6237,N_5803,N_5800);
and U6238 (N_6238,N_5890,N_5791);
nor U6239 (N_6239,N_5584,N_5935);
nand U6240 (N_6240,N_5914,N_5517);
nand U6241 (N_6241,N_5534,N_5624);
nor U6242 (N_6242,N_5538,N_5770);
and U6243 (N_6243,N_5588,N_5625);
xnor U6244 (N_6244,N_5856,N_5915);
and U6245 (N_6245,N_5515,N_5644);
xor U6246 (N_6246,N_5712,N_5936);
nor U6247 (N_6247,N_5984,N_5934);
and U6248 (N_6248,N_5756,N_5887);
nor U6249 (N_6249,N_5767,N_5508);
and U6250 (N_6250,N_5922,N_5791);
or U6251 (N_6251,N_5639,N_5677);
or U6252 (N_6252,N_5653,N_5672);
nand U6253 (N_6253,N_5768,N_5896);
nor U6254 (N_6254,N_5573,N_5992);
xor U6255 (N_6255,N_5985,N_5940);
nor U6256 (N_6256,N_5604,N_5972);
nor U6257 (N_6257,N_5747,N_5726);
or U6258 (N_6258,N_5884,N_5501);
and U6259 (N_6259,N_5839,N_5879);
or U6260 (N_6260,N_5575,N_5869);
and U6261 (N_6261,N_5530,N_5747);
or U6262 (N_6262,N_5867,N_5681);
or U6263 (N_6263,N_5631,N_5827);
nor U6264 (N_6264,N_5980,N_5859);
and U6265 (N_6265,N_5867,N_5642);
and U6266 (N_6266,N_5911,N_5684);
nand U6267 (N_6267,N_5980,N_5895);
nand U6268 (N_6268,N_5611,N_5985);
and U6269 (N_6269,N_5701,N_5624);
or U6270 (N_6270,N_5512,N_5626);
or U6271 (N_6271,N_5569,N_5894);
nor U6272 (N_6272,N_5646,N_5784);
or U6273 (N_6273,N_5996,N_5994);
and U6274 (N_6274,N_5575,N_5747);
nand U6275 (N_6275,N_5605,N_5612);
nor U6276 (N_6276,N_5695,N_5738);
nor U6277 (N_6277,N_5873,N_5822);
or U6278 (N_6278,N_5956,N_5784);
or U6279 (N_6279,N_5929,N_5937);
nand U6280 (N_6280,N_5596,N_5891);
nor U6281 (N_6281,N_5774,N_5872);
and U6282 (N_6282,N_5777,N_5956);
nor U6283 (N_6283,N_5680,N_5806);
and U6284 (N_6284,N_5732,N_5615);
or U6285 (N_6285,N_5531,N_5816);
nor U6286 (N_6286,N_5778,N_5766);
nor U6287 (N_6287,N_5822,N_5979);
nor U6288 (N_6288,N_5588,N_5788);
or U6289 (N_6289,N_5952,N_5714);
and U6290 (N_6290,N_5687,N_5608);
nand U6291 (N_6291,N_5758,N_5539);
nor U6292 (N_6292,N_5995,N_5790);
and U6293 (N_6293,N_5751,N_5956);
or U6294 (N_6294,N_5809,N_5983);
or U6295 (N_6295,N_5744,N_5630);
or U6296 (N_6296,N_5508,N_5936);
and U6297 (N_6297,N_5840,N_5968);
nor U6298 (N_6298,N_5932,N_5874);
xnor U6299 (N_6299,N_5677,N_5995);
or U6300 (N_6300,N_5646,N_5975);
or U6301 (N_6301,N_5623,N_5727);
and U6302 (N_6302,N_5513,N_5872);
or U6303 (N_6303,N_5501,N_5968);
and U6304 (N_6304,N_5932,N_5672);
or U6305 (N_6305,N_5851,N_5877);
xnor U6306 (N_6306,N_5873,N_5603);
and U6307 (N_6307,N_5650,N_5527);
nor U6308 (N_6308,N_5683,N_5900);
or U6309 (N_6309,N_5732,N_5612);
or U6310 (N_6310,N_5758,N_5967);
or U6311 (N_6311,N_5991,N_5524);
nor U6312 (N_6312,N_5539,N_5979);
nor U6313 (N_6313,N_5856,N_5818);
nand U6314 (N_6314,N_5574,N_5829);
xor U6315 (N_6315,N_5928,N_5706);
or U6316 (N_6316,N_5642,N_5783);
or U6317 (N_6317,N_5733,N_5843);
nor U6318 (N_6318,N_5559,N_5673);
and U6319 (N_6319,N_5716,N_5928);
nor U6320 (N_6320,N_5698,N_5632);
nor U6321 (N_6321,N_5993,N_5671);
nand U6322 (N_6322,N_5675,N_5751);
or U6323 (N_6323,N_5935,N_5790);
and U6324 (N_6324,N_5527,N_5910);
nand U6325 (N_6325,N_5521,N_5748);
and U6326 (N_6326,N_5915,N_5874);
and U6327 (N_6327,N_5831,N_5857);
and U6328 (N_6328,N_5820,N_5811);
nor U6329 (N_6329,N_5757,N_5717);
nor U6330 (N_6330,N_5580,N_5698);
or U6331 (N_6331,N_5932,N_5844);
nand U6332 (N_6332,N_5506,N_5894);
xor U6333 (N_6333,N_5808,N_5926);
or U6334 (N_6334,N_5767,N_5771);
nand U6335 (N_6335,N_5923,N_5917);
or U6336 (N_6336,N_5513,N_5548);
xnor U6337 (N_6337,N_5921,N_5699);
nand U6338 (N_6338,N_5581,N_5701);
or U6339 (N_6339,N_5875,N_5770);
nor U6340 (N_6340,N_5876,N_5788);
or U6341 (N_6341,N_5613,N_5669);
nand U6342 (N_6342,N_5963,N_5519);
nor U6343 (N_6343,N_5607,N_5690);
xnor U6344 (N_6344,N_5764,N_5901);
xnor U6345 (N_6345,N_5642,N_5854);
and U6346 (N_6346,N_5985,N_5615);
nand U6347 (N_6347,N_5942,N_5839);
or U6348 (N_6348,N_5910,N_5703);
nand U6349 (N_6349,N_5518,N_5895);
and U6350 (N_6350,N_5670,N_5514);
and U6351 (N_6351,N_5857,N_5520);
and U6352 (N_6352,N_5501,N_5855);
and U6353 (N_6353,N_5587,N_5876);
nand U6354 (N_6354,N_5550,N_5623);
or U6355 (N_6355,N_5734,N_5815);
nand U6356 (N_6356,N_5824,N_5569);
nor U6357 (N_6357,N_5585,N_5641);
nor U6358 (N_6358,N_5789,N_5502);
and U6359 (N_6359,N_5612,N_5520);
nand U6360 (N_6360,N_5636,N_5927);
nand U6361 (N_6361,N_5532,N_5960);
and U6362 (N_6362,N_5672,N_5783);
nor U6363 (N_6363,N_5878,N_5665);
and U6364 (N_6364,N_5975,N_5671);
and U6365 (N_6365,N_5633,N_5976);
or U6366 (N_6366,N_5874,N_5532);
and U6367 (N_6367,N_5960,N_5571);
nand U6368 (N_6368,N_5562,N_5529);
or U6369 (N_6369,N_5595,N_5778);
and U6370 (N_6370,N_5894,N_5675);
or U6371 (N_6371,N_5970,N_5926);
and U6372 (N_6372,N_5789,N_5714);
nand U6373 (N_6373,N_5901,N_5955);
xnor U6374 (N_6374,N_5809,N_5813);
nor U6375 (N_6375,N_5928,N_5549);
nor U6376 (N_6376,N_5561,N_5870);
nand U6377 (N_6377,N_5786,N_5719);
or U6378 (N_6378,N_5577,N_5664);
nand U6379 (N_6379,N_5753,N_5936);
and U6380 (N_6380,N_5602,N_5574);
or U6381 (N_6381,N_5556,N_5531);
or U6382 (N_6382,N_5637,N_5961);
and U6383 (N_6383,N_5884,N_5663);
and U6384 (N_6384,N_5932,N_5553);
nor U6385 (N_6385,N_5737,N_5829);
xor U6386 (N_6386,N_5809,N_5691);
nor U6387 (N_6387,N_5506,N_5663);
and U6388 (N_6388,N_5859,N_5600);
nand U6389 (N_6389,N_5761,N_5534);
xnor U6390 (N_6390,N_5881,N_5572);
or U6391 (N_6391,N_5774,N_5584);
or U6392 (N_6392,N_5744,N_5864);
nand U6393 (N_6393,N_5775,N_5850);
xor U6394 (N_6394,N_5550,N_5661);
or U6395 (N_6395,N_5881,N_5923);
nand U6396 (N_6396,N_5677,N_5950);
nor U6397 (N_6397,N_5759,N_5736);
or U6398 (N_6398,N_5903,N_5757);
and U6399 (N_6399,N_5995,N_5956);
or U6400 (N_6400,N_5528,N_5585);
nand U6401 (N_6401,N_5841,N_5610);
nand U6402 (N_6402,N_5740,N_5822);
and U6403 (N_6403,N_5943,N_5947);
or U6404 (N_6404,N_5949,N_5879);
nand U6405 (N_6405,N_5772,N_5747);
or U6406 (N_6406,N_5556,N_5652);
and U6407 (N_6407,N_5600,N_5736);
and U6408 (N_6408,N_5724,N_5568);
or U6409 (N_6409,N_5650,N_5592);
and U6410 (N_6410,N_5644,N_5590);
nand U6411 (N_6411,N_5651,N_5639);
or U6412 (N_6412,N_5891,N_5580);
and U6413 (N_6413,N_5591,N_5559);
xor U6414 (N_6414,N_5748,N_5792);
nand U6415 (N_6415,N_5564,N_5780);
nor U6416 (N_6416,N_5985,N_5594);
xnor U6417 (N_6417,N_5723,N_5886);
xnor U6418 (N_6418,N_5844,N_5633);
nand U6419 (N_6419,N_5874,N_5760);
nor U6420 (N_6420,N_5538,N_5729);
and U6421 (N_6421,N_5761,N_5624);
nor U6422 (N_6422,N_5566,N_5859);
and U6423 (N_6423,N_5674,N_5734);
and U6424 (N_6424,N_5584,N_5636);
nand U6425 (N_6425,N_5654,N_5639);
nor U6426 (N_6426,N_5716,N_5528);
or U6427 (N_6427,N_5799,N_5649);
and U6428 (N_6428,N_5719,N_5657);
and U6429 (N_6429,N_5639,N_5948);
nand U6430 (N_6430,N_5629,N_5815);
nor U6431 (N_6431,N_5801,N_5716);
nor U6432 (N_6432,N_5997,N_5646);
or U6433 (N_6433,N_5540,N_5604);
nor U6434 (N_6434,N_5807,N_5591);
nand U6435 (N_6435,N_5864,N_5566);
or U6436 (N_6436,N_5772,N_5537);
nor U6437 (N_6437,N_5570,N_5684);
nand U6438 (N_6438,N_5609,N_5846);
nand U6439 (N_6439,N_5845,N_5832);
and U6440 (N_6440,N_5779,N_5712);
and U6441 (N_6441,N_5670,N_5756);
nor U6442 (N_6442,N_5855,N_5844);
nand U6443 (N_6443,N_5667,N_5954);
nor U6444 (N_6444,N_5714,N_5794);
and U6445 (N_6445,N_5834,N_5554);
and U6446 (N_6446,N_5704,N_5542);
and U6447 (N_6447,N_5977,N_5761);
nand U6448 (N_6448,N_5874,N_5525);
or U6449 (N_6449,N_5504,N_5772);
or U6450 (N_6450,N_5806,N_5578);
xnor U6451 (N_6451,N_5921,N_5820);
or U6452 (N_6452,N_5640,N_5543);
nand U6453 (N_6453,N_5879,N_5831);
or U6454 (N_6454,N_5722,N_5894);
xor U6455 (N_6455,N_5608,N_5912);
or U6456 (N_6456,N_5993,N_5719);
and U6457 (N_6457,N_5948,N_5930);
or U6458 (N_6458,N_5839,N_5960);
or U6459 (N_6459,N_5552,N_5911);
and U6460 (N_6460,N_5732,N_5812);
or U6461 (N_6461,N_5714,N_5802);
nand U6462 (N_6462,N_5869,N_5753);
nand U6463 (N_6463,N_5919,N_5500);
nor U6464 (N_6464,N_5895,N_5929);
nand U6465 (N_6465,N_5906,N_5733);
nand U6466 (N_6466,N_5930,N_5920);
nor U6467 (N_6467,N_5662,N_5665);
nand U6468 (N_6468,N_5654,N_5981);
xnor U6469 (N_6469,N_5820,N_5996);
nand U6470 (N_6470,N_5921,N_5596);
and U6471 (N_6471,N_5626,N_5745);
or U6472 (N_6472,N_5639,N_5519);
and U6473 (N_6473,N_5659,N_5908);
and U6474 (N_6474,N_5937,N_5801);
nand U6475 (N_6475,N_5999,N_5625);
or U6476 (N_6476,N_5717,N_5926);
or U6477 (N_6477,N_5811,N_5920);
or U6478 (N_6478,N_5926,N_5858);
nor U6479 (N_6479,N_5744,N_5505);
nand U6480 (N_6480,N_5888,N_5927);
or U6481 (N_6481,N_5707,N_5599);
or U6482 (N_6482,N_5891,N_5586);
xnor U6483 (N_6483,N_5899,N_5992);
and U6484 (N_6484,N_5658,N_5923);
nor U6485 (N_6485,N_5957,N_5787);
nor U6486 (N_6486,N_5532,N_5985);
nor U6487 (N_6487,N_5582,N_5563);
xor U6488 (N_6488,N_5747,N_5612);
nor U6489 (N_6489,N_5866,N_5565);
nor U6490 (N_6490,N_5931,N_5965);
xnor U6491 (N_6491,N_5769,N_5522);
and U6492 (N_6492,N_5803,N_5617);
or U6493 (N_6493,N_5920,N_5772);
nor U6494 (N_6494,N_5524,N_5919);
or U6495 (N_6495,N_5964,N_5870);
nand U6496 (N_6496,N_5929,N_5650);
nand U6497 (N_6497,N_5531,N_5894);
nand U6498 (N_6498,N_5940,N_5952);
nor U6499 (N_6499,N_5918,N_5586);
or U6500 (N_6500,N_6494,N_6289);
nand U6501 (N_6501,N_6135,N_6389);
nor U6502 (N_6502,N_6234,N_6142);
nand U6503 (N_6503,N_6177,N_6496);
or U6504 (N_6504,N_6387,N_6174);
nor U6505 (N_6505,N_6036,N_6356);
and U6506 (N_6506,N_6286,N_6195);
or U6507 (N_6507,N_6445,N_6452);
nand U6508 (N_6508,N_6465,N_6398);
nor U6509 (N_6509,N_6091,N_6183);
nand U6510 (N_6510,N_6330,N_6053);
and U6511 (N_6511,N_6161,N_6369);
and U6512 (N_6512,N_6350,N_6487);
nor U6513 (N_6513,N_6360,N_6017);
nand U6514 (N_6514,N_6282,N_6170);
xor U6515 (N_6515,N_6086,N_6168);
nand U6516 (N_6516,N_6146,N_6213);
nand U6517 (N_6517,N_6429,N_6424);
nor U6518 (N_6518,N_6394,N_6007);
or U6519 (N_6519,N_6020,N_6442);
and U6520 (N_6520,N_6192,N_6284);
nor U6521 (N_6521,N_6175,N_6422);
nor U6522 (N_6522,N_6305,N_6241);
nand U6523 (N_6523,N_6497,N_6434);
nor U6524 (N_6524,N_6064,N_6019);
or U6525 (N_6525,N_6204,N_6140);
nor U6526 (N_6526,N_6029,N_6478);
nand U6527 (N_6527,N_6261,N_6331);
or U6528 (N_6528,N_6093,N_6155);
xnor U6529 (N_6529,N_6198,N_6426);
nand U6530 (N_6530,N_6358,N_6345);
or U6531 (N_6531,N_6315,N_6016);
or U6532 (N_6532,N_6062,N_6061);
and U6533 (N_6533,N_6105,N_6240);
nor U6534 (N_6534,N_6215,N_6132);
nand U6535 (N_6535,N_6436,N_6484);
and U6536 (N_6536,N_6216,N_6042);
and U6537 (N_6537,N_6208,N_6136);
nor U6538 (N_6538,N_6328,N_6413);
and U6539 (N_6539,N_6089,N_6226);
and U6540 (N_6540,N_6131,N_6334);
or U6541 (N_6541,N_6194,N_6110);
xnor U6542 (N_6542,N_6324,N_6073);
and U6543 (N_6543,N_6364,N_6302);
nand U6544 (N_6544,N_6291,N_6081);
or U6545 (N_6545,N_6092,N_6431);
and U6546 (N_6546,N_6269,N_6336);
nor U6547 (N_6547,N_6169,N_6023);
nand U6548 (N_6548,N_6124,N_6102);
or U6549 (N_6549,N_6243,N_6219);
or U6550 (N_6550,N_6475,N_6233);
and U6551 (N_6551,N_6108,N_6157);
or U6552 (N_6552,N_6236,N_6217);
nor U6553 (N_6553,N_6249,N_6248);
and U6554 (N_6554,N_6079,N_6392);
or U6555 (N_6555,N_6407,N_6099);
nor U6556 (N_6556,N_6279,N_6116);
or U6557 (N_6557,N_6164,N_6069);
nor U6558 (N_6558,N_6259,N_6461);
nor U6559 (N_6559,N_6239,N_6244);
and U6560 (N_6560,N_6276,N_6321);
or U6561 (N_6561,N_6154,N_6314);
xor U6562 (N_6562,N_6097,N_6372);
xnor U6563 (N_6563,N_6408,N_6067);
nand U6564 (N_6564,N_6375,N_6310);
or U6565 (N_6565,N_6415,N_6048);
nand U6566 (N_6566,N_6405,N_6171);
nor U6567 (N_6567,N_6278,N_6410);
and U6568 (N_6568,N_6256,N_6166);
and U6569 (N_6569,N_6211,N_6059);
or U6570 (N_6570,N_6128,N_6425);
nand U6571 (N_6571,N_6271,N_6160);
or U6572 (N_6572,N_6209,N_6404);
xnor U6573 (N_6573,N_6222,N_6148);
or U6574 (N_6574,N_6228,N_6270);
nor U6575 (N_6575,N_6125,N_6308);
nand U6576 (N_6576,N_6280,N_6285);
nor U6577 (N_6577,N_6218,N_6362);
xnor U6578 (N_6578,N_6423,N_6187);
nor U6579 (N_6579,N_6260,N_6316);
nand U6580 (N_6580,N_6051,N_6338);
nor U6581 (N_6581,N_6141,N_6273);
nor U6582 (N_6582,N_6022,N_6400);
nor U6583 (N_6583,N_6317,N_6201);
or U6584 (N_6584,N_6147,N_6298);
and U6585 (N_6585,N_6420,N_6185);
nand U6586 (N_6586,N_6004,N_6179);
or U6587 (N_6587,N_6403,N_6001);
nor U6588 (N_6588,N_6013,N_6223);
and U6589 (N_6589,N_6245,N_6045);
nor U6590 (N_6590,N_6072,N_6242);
or U6591 (N_6591,N_6439,N_6402);
nor U6592 (N_6592,N_6353,N_6459);
and U6593 (N_6593,N_6227,N_6491);
nand U6594 (N_6594,N_6390,N_6152);
nand U6595 (N_6595,N_6378,N_6320);
or U6596 (N_6596,N_6130,N_6176);
nor U6597 (N_6597,N_6368,N_6065);
or U6598 (N_6598,N_6082,N_6167);
nor U6599 (N_6599,N_6150,N_6457);
and U6600 (N_6600,N_6275,N_6351);
and U6601 (N_6601,N_6448,N_6447);
xor U6602 (N_6602,N_6458,N_6193);
nand U6603 (N_6603,N_6397,N_6078);
and U6604 (N_6604,N_6137,N_6266);
nand U6605 (N_6605,N_6467,N_6250);
nor U6606 (N_6606,N_6488,N_6262);
nand U6607 (N_6607,N_6230,N_6172);
and U6608 (N_6608,N_6033,N_6307);
nor U6609 (N_6609,N_6460,N_6277);
or U6610 (N_6610,N_6163,N_6455);
nor U6611 (N_6611,N_6388,N_6437);
nor U6612 (N_6612,N_6348,N_6258);
nand U6613 (N_6613,N_6470,N_6071);
or U6614 (N_6614,N_6114,N_6225);
nor U6615 (N_6615,N_6479,N_6237);
nor U6616 (N_6616,N_6432,N_6296);
nor U6617 (N_6617,N_6098,N_6210);
or U6618 (N_6618,N_6156,N_6083);
nand U6619 (N_6619,N_6224,N_6481);
or U6620 (N_6620,N_6034,N_6006);
and U6621 (N_6621,N_6035,N_6220);
xor U6622 (N_6622,N_6133,N_6354);
nand U6623 (N_6623,N_6367,N_6274);
nor U6624 (N_6624,N_6341,N_6121);
xnor U6625 (N_6625,N_6196,N_6363);
nor U6626 (N_6626,N_6463,N_6444);
and U6627 (N_6627,N_6009,N_6385);
nand U6628 (N_6628,N_6145,N_6323);
nor U6629 (N_6629,N_6018,N_6485);
and U6630 (N_6630,N_6039,N_6205);
nand U6631 (N_6631,N_6106,N_6382);
and U6632 (N_6632,N_6295,N_6028);
or U6633 (N_6633,N_6347,N_6199);
nor U6634 (N_6634,N_6293,N_6346);
or U6635 (N_6635,N_6438,N_6427);
or U6636 (N_6636,N_6104,N_6359);
nor U6637 (N_6637,N_6120,N_6085);
nor U6638 (N_6638,N_6464,N_6060);
nor U6639 (N_6639,N_6361,N_6200);
or U6640 (N_6640,N_6471,N_6326);
and U6641 (N_6641,N_6070,N_6096);
or U6642 (N_6642,N_6299,N_6221);
xnor U6643 (N_6643,N_6318,N_6232);
xor U6644 (N_6644,N_6474,N_6430);
or U6645 (N_6645,N_6376,N_6038);
nor U6646 (N_6646,N_6186,N_6134);
nand U6647 (N_6647,N_6342,N_6386);
nand U6648 (N_6648,N_6235,N_6265);
and U6649 (N_6649,N_6127,N_6068);
and U6650 (N_6650,N_6349,N_6483);
or U6651 (N_6651,N_6396,N_6477);
and U6652 (N_6652,N_6139,N_6181);
and U6653 (N_6653,N_6153,N_6165);
nor U6654 (N_6654,N_6428,N_6026);
and U6655 (N_6655,N_6066,N_6393);
nor U6656 (N_6656,N_6357,N_6272);
nand U6657 (N_6657,N_6063,N_6352);
nand U6658 (N_6658,N_6443,N_6419);
nor U6659 (N_6659,N_6313,N_6456);
or U6660 (N_6660,N_6008,N_6189);
nand U6661 (N_6661,N_6409,N_6468);
nor U6662 (N_6662,N_6057,N_6300);
nand U6663 (N_6663,N_6129,N_6080);
nor U6664 (N_6664,N_6406,N_6107);
and U6665 (N_6665,N_6040,N_6188);
xnor U6666 (N_6666,N_6319,N_6077);
nor U6667 (N_6667,N_6149,N_6476);
or U6668 (N_6668,N_6103,N_6311);
or U6669 (N_6669,N_6440,N_6325);
or U6670 (N_6670,N_6257,N_6414);
nor U6671 (N_6671,N_6399,N_6138);
nor U6672 (N_6672,N_6451,N_6301);
nor U6673 (N_6673,N_6123,N_6005);
nand U6674 (N_6674,N_6446,N_6012);
or U6675 (N_6675,N_6011,N_6044);
nor U6676 (N_6676,N_6290,N_6395);
or U6677 (N_6677,N_6037,N_6435);
and U6678 (N_6678,N_6370,N_6084);
or U6679 (N_6679,N_6094,N_6306);
nor U6680 (N_6680,N_6333,N_6251);
nor U6681 (N_6681,N_6117,N_6087);
or U6682 (N_6682,N_6109,N_6238);
nand U6683 (N_6683,N_6052,N_6203);
nand U6684 (N_6684,N_6229,N_6088);
nor U6685 (N_6685,N_6207,N_6214);
nand U6686 (N_6686,N_6264,N_6492);
and U6687 (N_6687,N_6100,N_6003);
and U6688 (N_6688,N_6373,N_6482);
and U6689 (N_6689,N_6281,N_6417);
nand U6690 (N_6690,N_6480,N_6441);
and U6691 (N_6691,N_6322,N_6113);
or U6692 (N_6692,N_6381,N_6355);
or U6693 (N_6693,N_6055,N_6499);
xnor U6694 (N_6694,N_6418,N_6252);
and U6695 (N_6695,N_6162,N_6056);
xnor U6696 (N_6696,N_6421,N_6283);
or U6697 (N_6697,N_6304,N_6118);
xnor U6698 (N_6698,N_6111,N_6294);
xor U6699 (N_6699,N_6000,N_6490);
nor U6700 (N_6700,N_6046,N_6473);
nand U6701 (N_6701,N_6493,N_6021);
nor U6702 (N_6702,N_6206,N_6365);
nand U6703 (N_6703,N_6015,N_6309);
or U6704 (N_6704,N_6495,N_6377);
nand U6705 (N_6705,N_6202,N_6246);
or U6706 (N_6706,N_6384,N_6090);
nand U6707 (N_6707,N_6247,N_6050);
nor U6708 (N_6708,N_6472,N_6058);
nand U6709 (N_6709,N_6151,N_6076);
or U6710 (N_6710,N_6380,N_6253);
and U6711 (N_6711,N_6374,N_6466);
or U6712 (N_6712,N_6335,N_6144);
nand U6713 (N_6713,N_6025,N_6344);
and U6714 (N_6714,N_6031,N_6498);
nor U6715 (N_6715,N_6416,N_6292);
and U6716 (N_6716,N_6332,N_6173);
nand U6717 (N_6717,N_6049,N_6371);
and U6718 (N_6718,N_6101,N_6054);
xor U6719 (N_6719,N_6433,N_6453);
nor U6720 (N_6720,N_6486,N_6343);
nand U6721 (N_6721,N_6297,N_6115);
or U6722 (N_6722,N_6391,N_6255);
nor U6723 (N_6723,N_6412,N_6047);
nand U6724 (N_6724,N_6191,N_6254);
xnor U6725 (N_6725,N_6288,N_6267);
nor U6726 (N_6726,N_6184,N_6027);
and U6727 (N_6727,N_6182,N_6450);
and U6728 (N_6728,N_6462,N_6329);
or U6729 (N_6729,N_6095,N_6024);
and U6730 (N_6730,N_6268,N_6411);
nand U6731 (N_6731,N_6340,N_6032);
or U6732 (N_6732,N_6180,N_6002);
xor U6733 (N_6733,N_6337,N_6143);
nor U6734 (N_6734,N_6231,N_6122);
nand U6735 (N_6735,N_6159,N_6449);
or U6736 (N_6736,N_6312,N_6075);
nand U6737 (N_6737,N_6158,N_6074);
xnor U6738 (N_6738,N_6263,N_6469);
xor U6739 (N_6739,N_6489,N_6112);
nor U6740 (N_6740,N_6327,N_6401);
or U6741 (N_6741,N_6366,N_6454);
nor U6742 (N_6742,N_6126,N_6303);
nor U6743 (N_6743,N_6383,N_6197);
xnor U6744 (N_6744,N_6190,N_6339);
or U6745 (N_6745,N_6014,N_6212);
nor U6746 (N_6746,N_6379,N_6287);
nand U6747 (N_6747,N_6178,N_6043);
and U6748 (N_6748,N_6030,N_6010);
and U6749 (N_6749,N_6041,N_6119);
and U6750 (N_6750,N_6005,N_6151);
nand U6751 (N_6751,N_6290,N_6335);
nor U6752 (N_6752,N_6140,N_6237);
or U6753 (N_6753,N_6390,N_6452);
and U6754 (N_6754,N_6389,N_6426);
and U6755 (N_6755,N_6125,N_6141);
or U6756 (N_6756,N_6499,N_6156);
nand U6757 (N_6757,N_6067,N_6364);
xor U6758 (N_6758,N_6437,N_6432);
nor U6759 (N_6759,N_6248,N_6254);
nor U6760 (N_6760,N_6400,N_6370);
or U6761 (N_6761,N_6460,N_6109);
nor U6762 (N_6762,N_6210,N_6477);
nor U6763 (N_6763,N_6388,N_6147);
xnor U6764 (N_6764,N_6150,N_6373);
or U6765 (N_6765,N_6244,N_6366);
nand U6766 (N_6766,N_6364,N_6170);
nor U6767 (N_6767,N_6310,N_6446);
and U6768 (N_6768,N_6457,N_6246);
nor U6769 (N_6769,N_6215,N_6317);
and U6770 (N_6770,N_6320,N_6498);
nand U6771 (N_6771,N_6185,N_6095);
and U6772 (N_6772,N_6227,N_6141);
and U6773 (N_6773,N_6070,N_6047);
nor U6774 (N_6774,N_6442,N_6174);
or U6775 (N_6775,N_6478,N_6209);
or U6776 (N_6776,N_6459,N_6182);
or U6777 (N_6777,N_6155,N_6103);
xnor U6778 (N_6778,N_6377,N_6384);
nor U6779 (N_6779,N_6296,N_6312);
nor U6780 (N_6780,N_6237,N_6067);
or U6781 (N_6781,N_6255,N_6493);
xor U6782 (N_6782,N_6261,N_6451);
or U6783 (N_6783,N_6107,N_6005);
or U6784 (N_6784,N_6212,N_6361);
or U6785 (N_6785,N_6443,N_6230);
nor U6786 (N_6786,N_6421,N_6439);
nand U6787 (N_6787,N_6042,N_6007);
or U6788 (N_6788,N_6498,N_6109);
and U6789 (N_6789,N_6468,N_6351);
and U6790 (N_6790,N_6371,N_6446);
nand U6791 (N_6791,N_6149,N_6394);
nand U6792 (N_6792,N_6429,N_6210);
or U6793 (N_6793,N_6133,N_6055);
xor U6794 (N_6794,N_6466,N_6245);
xnor U6795 (N_6795,N_6061,N_6473);
nand U6796 (N_6796,N_6416,N_6040);
and U6797 (N_6797,N_6309,N_6125);
or U6798 (N_6798,N_6333,N_6479);
nor U6799 (N_6799,N_6165,N_6424);
or U6800 (N_6800,N_6492,N_6100);
or U6801 (N_6801,N_6019,N_6088);
nand U6802 (N_6802,N_6086,N_6339);
or U6803 (N_6803,N_6039,N_6072);
or U6804 (N_6804,N_6218,N_6357);
and U6805 (N_6805,N_6272,N_6046);
nor U6806 (N_6806,N_6272,N_6211);
or U6807 (N_6807,N_6004,N_6210);
nor U6808 (N_6808,N_6455,N_6062);
nand U6809 (N_6809,N_6010,N_6437);
nand U6810 (N_6810,N_6348,N_6061);
nor U6811 (N_6811,N_6129,N_6156);
nor U6812 (N_6812,N_6004,N_6391);
or U6813 (N_6813,N_6083,N_6048);
nand U6814 (N_6814,N_6239,N_6073);
nand U6815 (N_6815,N_6429,N_6304);
xnor U6816 (N_6816,N_6340,N_6459);
nor U6817 (N_6817,N_6343,N_6385);
nand U6818 (N_6818,N_6048,N_6269);
nor U6819 (N_6819,N_6120,N_6406);
nand U6820 (N_6820,N_6314,N_6396);
and U6821 (N_6821,N_6105,N_6355);
or U6822 (N_6822,N_6489,N_6022);
nor U6823 (N_6823,N_6364,N_6291);
xnor U6824 (N_6824,N_6030,N_6346);
and U6825 (N_6825,N_6127,N_6027);
xnor U6826 (N_6826,N_6430,N_6076);
and U6827 (N_6827,N_6237,N_6124);
or U6828 (N_6828,N_6239,N_6309);
nand U6829 (N_6829,N_6024,N_6297);
xnor U6830 (N_6830,N_6056,N_6326);
nand U6831 (N_6831,N_6395,N_6057);
or U6832 (N_6832,N_6455,N_6227);
and U6833 (N_6833,N_6316,N_6204);
nand U6834 (N_6834,N_6330,N_6285);
nand U6835 (N_6835,N_6371,N_6265);
or U6836 (N_6836,N_6430,N_6196);
nand U6837 (N_6837,N_6485,N_6210);
or U6838 (N_6838,N_6194,N_6400);
nand U6839 (N_6839,N_6103,N_6285);
or U6840 (N_6840,N_6405,N_6183);
and U6841 (N_6841,N_6479,N_6008);
and U6842 (N_6842,N_6281,N_6457);
nor U6843 (N_6843,N_6476,N_6077);
nand U6844 (N_6844,N_6419,N_6136);
nand U6845 (N_6845,N_6361,N_6350);
or U6846 (N_6846,N_6499,N_6038);
nor U6847 (N_6847,N_6303,N_6496);
or U6848 (N_6848,N_6156,N_6257);
nand U6849 (N_6849,N_6363,N_6285);
nand U6850 (N_6850,N_6066,N_6039);
nand U6851 (N_6851,N_6002,N_6266);
nand U6852 (N_6852,N_6163,N_6402);
nand U6853 (N_6853,N_6214,N_6219);
and U6854 (N_6854,N_6027,N_6013);
nor U6855 (N_6855,N_6167,N_6079);
nor U6856 (N_6856,N_6112,N_6484);
nor U6857 (N_6857,N_6471,N_6120);
nand U6858 (N_6858,N_6401,N_6304);
or U6859 (N_6859,N_6090,N_6362);
nand U6860 (N_6860,N_6177,N_6474);
and U6861 (N_6861,N_6430,N_6371);
and U6862 (N_6862,N_6018,N_6355);
nor U6863 (N_6863,N_6407,N_6138);
or U6864 (N_6864,N_6244,N_6127);
or U6865 (N_6865,N_6339,N_6096);
or U6866 (N_6866,N_6281,N_6137);
or U6867 (N_6867,N_6028,N_6450);
and U6868 (N_6868,N_6016,N_6243);
and U6869 (N_6869,N_6341,N_6457);
nor U6870 (N_6870,N_6083,N_6257);
or U6871 (N_6871,N_6256,N_6018);
nand U6872 (N_6872,N_6375,N_6473);
and U6873 (N_6873,N_6283,N_6167);
xor U6874 (N_6874,N_6040,N_6250);
or U6875 (N_6875,N_6069,N_6103);
and U6876 (N_6876,N_6342,N_6192);
nand U6877 (N_6877,N_6308,N_6195);
xnor U6878 (N_6878,N_6017,N_6202);
nor U6879 (N_6879,N_6095,N_6099);
nor U6880 (N_6880,N_6086,N_6136);
and U6881 (N_6881,N_6311,N_6302);
nand U6882 (N_6882,N_6410,N_6274);
and U6883 (N_6883,N_6022,N_6141);
nand U6884 (N_6884,N_6117,N_6178);
nor U6885 (N_6885,N_6013,N_6330);
nor U6886 (N_6886,N_6463,N_6207);
nand U6887 (N_6887,N_6023,N_6340);
xnor U6888 (N_6888,N_6203,N_6390);
or U6889 (N_6889,N_6491,N_6380);
or U6890 (N_6890,N_6215,N_6346);
or U6891 (N_6891,N_6297,N_6396);
nand U6892 (N_6892,N_6332,N_6362);
nand U6893 (N_6893,N_6024,N_6404);
or U6894 (N_6894,N_6063,N_6398);
nand U6895 (N_6895,N_6283,N_6300);
and U6896 (N_6896,N_6204,N_6149);
xor U6897 (N_6897,N_6334,N_6044);
and U6898 (N_6898,N_6396,N_6097);
and U6899 (N_6899,N_6271,N_6482);
nor U6900 (N_6900,N_6364,N_6215);
nor U6901 (N_6901,N_6491,N_6003);
nand U6902 (N_6902,N_6442,N_6011);
nor U6903 (N_6903,N_6182,N_6481);
and U6904 (N_6904,N_6006,N_6431);
and U6905 (N_6905,N_6248,N_6288);
and U6906 (N_6906,N_6452,N_6393);
nor U6907 (N_6907,N_6395,N_6082);
or U6908 (N_6908,N_6431,N_6322);
nand U6909 (N_6909,N_6225,N_6468);
or U6910 (N_6910,N_6002,N_6056);
and U6911 (N_6911,N_6485,N_6234);
nor U6912 (N_6912,N_6307,N_6059);
nor U6913 (N_6913,N_6157,N_6216);
nand U6914 (N_6914,N_6428,N_6013);
and U6915 (N_6915,N_6411,N_6175);
nand U6916 (N_6916,N_6422,N_6344);
or U6917 (N_6917,N_6326,N_6481);
nand U6918 (N_6918,N_6095,N_6089);
or U6919 (N_6919,N_6491,N_6432);
nor U6920 (N_6920,N_6403,N_6018);
or U6921 (N_6921,N_6443,N_6001);
nand U6922 (N_6922,N_6181,N_6105);
and U6923 (N_6923,N_6471,N_6154);
xnor U6924 (N_6924,N_6489,N_6210);
xnor U6925 (N_6925,N_6365,N_6441);
or U6926 (N_6926,N_6078,N_6202);
nand U6927 (N_6927,N_6203,N_6374);
xor U6928 (N_6928,N_6408,N_6027);
nor U6929 (N_6929,N_6051,N_6073);
nand U6930 (N_6930,N_6188,N_6272);
and U6931 (N_6931,N_6446,N_6449);
nor U6932 (N_6932,N_6001,N_6355);
and U6933 (N_6933,N_6053,N_6353);
nor U6934 (N_6934,N_6046,N_6405);
nand U6935 (N_6935,N_6321,N_6017);
nor U6936 (N_6936,N_6345,N_6216);
nand U6937 (N_6937,N_6278,N_6418);
and U6938 (N_6938,N_6212,N_6203);
nand U6939 (N_6939,N_6345,N_6332);
nor U6940 (N_6940,N_6046,N_6203);
nor U6941 (N_6941,N_6400,N_6360);
nor U6942 (N_6942,N_6060,N_6455);
or U6943 (N_6943,N_6343,N_6247);
or U6944 (N_6944,N_6131,N_6162);
and U6945 (N_6945,N_6121,N_6279);
and U6946 (N_6946,N_6406,N_6464);
and U6947 (N_6947,N_6350,N_6277);
xnor U6948 (N_6948,N_6238,N_6452);
and U6949 (N_6949,N_6141,N_6380);
nand U6950 (N_6950,N_6118,N_6139);
nor U6951 (N_6951,N_6367,N_6447);
nand U6952 (N_6952,N_6218,N_6115);
or U6953 (N_6953,N_6199,N_6467);
nor U6954 (N_6954,N_6451,N_6032);
nor U6955 (N_6955,N_6338,N_6032);
nand U6956 (N_6956,N_6373,N_6243);
nand U6957 (N_6957,N_6116,N_6073);
and U6958 (N_6958,N_6005,N_6358);
or U6959 (N_6959,N_6301,N_6316);
and U6960 (N_6960,N_6146,N_6180);
nand U6961 (N_6961,N_6325,N_6109);
nor U6962 (N_6962,N_6079,N_6482);
xnor U6963 (N_6963,N_6190,N_6064);
and U6964 (N_6964,N_6107,N_6489);
or U6965 (N_6965,N_6360,N_6215);
nand U6966 (N_6966,N_6052,N_6286);
and U6967 (N_6967,N_6419,N_6014);
nand U6968 (N_6968,N_6404,N_6460);
nand U6969 (N_6969,N_6459,N_6228);
nor U6970 (N_6970,N_6188,N_6050);
nand U6971 (N_6971,N_6424,N_6059);
or U6972 (N_6972,N_6435,N_6092);
and U6973 (N_6973,N_6103,N_6328);
nor U6974 (N_6974,N_6411,N_6013);
nand U6975 (N_6975,N_6134,N_6315);
nand U6976 (N_6976,N_6017,N_6332);
nand U6977 (N_6977,N_6111,N_6053);
or U6978 (N_6978,N_6029,N_6471);
and U6979 (N_6979,N_6023,N_6376);
and U6980 (N_6980,N_6458,N_6450);
or U6981 (N_6981,N_6076,N_6295);
or U6982 (N_6982,N_6334,N_6280);
xor U6983 (N_6983,N_6340,N_6145);
nand U6984 (N_6984,N_6194,N_6050);
nor U6985 (N_6985,N_6068,N_6182);
or U6986 (N_6986,N_6378,N_6487);
xnor U6987 (N_6987,N_6179,N_6479);
nand U6988 (N_6988,N_6319,N_6072);
and U6989 (N_6989,N_6085,N_6099);
nand U6990 (N_6990,N_6302,N_6490);
nor U6991 (N_6991,N_6093,N_6204);
and U6992 (N_6992,N_6481,N_6264);
and U6993 (N_6993,N_6446,N_6478);
or U6994 (N_6994,N_6374,N_6123);
nor U6995 (N_6995,N_6015,N_6179);
nor U6996 (N_6996,N_6361,N_6221);
nor U6997 (N_6997,N_6042,N_6342);
nor U6998 (N_6998,N_6088,N_6193);
and U6999 (N_6999,N_6200,N_6073);
xor U7000 (N_7000,N_6748,N_6845);
or U7001 (N_7001,N_6516,N_6518);
nand U7002 (N_7002,N_6504,N_6618);
xnor U7003 (N_7003,N_6558,N_6958);
or U7004 (N_7004,N_6651,N_6529);
and U7005 (N_7005,N_6640,N_6714);
nor U7006 (N_7006,N_6637,N_6764);
nand U7007 (N_7007,N_6786,N_6696);
nor U7008 (N_7008,N_6898,N_6857);
xor U7009 (N_7009,N_6683,N_6660);
and U7010 (N_7010,N_6595,N_6545);
and U7011 (N_7011,N_6768,N_6820);
or U7012 (N_7012,N_6657,N_6578);
nand U7013 (N_7013,N_6589,N_6966);
nand U7014 (N_7014,N_6963,N_6724);
and U7015 (N_7015,N_6801,N_6766);
nor U7016 (N_7016,N_6612,N_6653);
nand U7017 (N_7017,N_6928,N_6987);
nand U7018 (N_7018,N_6508,N_6868);
and U7019 (N_7019,N_6909,N_6775);
and U7020 (N_7020,N_6541,N_6590);
xnor U7021 (N_7021,N_6770,N_6831);
nand U7022 (N_7022,N_6783,N_6995);
xnor U7023 (N_7023,N_6559,N_6893);
nor U7024 (N_7024,N_6846,N_6607);
nand U7025 (N_7025,N_6567,N_6955);
nor U7026 (N_7026,N_6742,N_6735);
or U7027 (N_7027,N_6732,N_6938);
nand U7028 (N_7028,N_6571,N_6933);
nand U7029 (N_7029,N_6645,N_6834);
and U7030 (N_7030,N_6745,N_6993);
and U7031 (N_7031,N_6982,N_6575);
xor U7032 (N_7032,N_6598,N_6581);
nand U7033 (N_7033,N_6599,N_6908);
and U7034 (N_7034,N_6899,N_6997);
nand U7035 (N_7035,N_6503,N_6673);
nand U7036 (N_7036,N_6750,N_6648);
nand U7037 (N_7037,N_6688,N_6897);
and U7038 (N_7038,N_6873,N_6716);
or U7039 (N_7039,N_6793,N_6782);
and U7040 (N_7040,N_6706,N_6551);
nor U7041 (N_7041,N_6836,N_6526);
nand U7042 (N_7042,N_6704,N_6668);
xor U7043 (N_7043,N_6540,N_6828);
nor U7044 (N_7044,N_6628,N_6697);
xor U7045 (N_7045,N_6659,N_6859);
and U7046 (N_7046,N_6729,N_6500);
or U7047 (N_7047,N_6794,N_6528);
and U7048 (N_7048,N_6725,N_6641);
or U7049 (N_7049,N_6813,N_6819);
or U7050 (N_7050,N_6656,N_6818);
and U7051 (N_7051,N_6988,N_6837);
and U7052 (N_7052,N_6989,N_6926);
and U7053 (N_7053,N_6821,N_6774);
nor U7054 (N_7054,N_6925,N_6755);
nor U7055 (N_7055,N_6597,N_6677);
nor U7056 (N_7056,N_6629,N_6727);
and U7057 (N_7057,N_6534,N_6773);
xnor U7058 (N_7058,N_6519,N_6515);
nor U7059 (N_7059,N_6736,N_6741);
nand U7060 (N_7060,N_6702,N_6544);
or U7061 (N_7061,N_6974,N_6728);
and U7062 (N_7062,N_6830,N_6743);
nand U7063 (N_7063,N_6666,N_6940);
nor U7064 (N_7064,N_6880,N_6754);
nor U7065 (N_7065,N_6761,N_6695);
or U7066 (N_7066,N_6879,N_6985);
and U7067 (N_7067,N_6979,N_6861);
or U7068 (N_7068,N_6901,N_6619);
or U7069 (N_7069,N_6603,N_6654);
nor U7070 (N_7070,N_6778,N_6611);
and U7071 (N_7071,N_6562,N_6717);
nand U7072 (N_7072,N_6751,N_6609);
or U7073 (N_7073,N_6864,N_6757);
nor U7074 (N_7074,N_6585,N_6892);
nand U7075 (N_7075,N_6701,N_6911);
nor U7076 (N_7076,N_6811,N_6682);
nor U7077 (N_7077,N_6721,N_6839);
nor U7078 (N_7078,N_6674,N_6984);
and U7079 (N_7079,N_6944,N_6825);
nand U7080 (N_7080,N_6552,N_6635);
nor U7081 (N_7081,N_6517,N_6872);
xor U7082 (N_7082,N_6905,N_6626);
nor U7083 (N_7083,N_6948,N_6690);
nand U7084 (N_7084,N_6891,N_6780);
nand U7085 (N_7085,N_6522,N_6885);
or U7086 (N_7086,N_6691,N_6887);
and U7087 (N_7087,N_6622,N_6588);
nor U7088 (N_7088,N_6882,N_6912);
and U7089 (N_7089,N_6527,N_6594);
nand U7090 (N_7090,N_6960,N_6554);
nor U7091 (N_7091,N_6835,N_6805);
nand U7092 (N_7092,N_6580,N_6903);
and U7093 (N_7093,N_6923,N_6951);
and U7094 (N_7094,N_6856,N_6680);
or U7095 (N_7095,N_6978,N_6665);
or U7096 (N_7096,N_6726,N_6624);
or U7097 (N_7097,N_6525,N_6556);
or U7098 (N_7098,N_6620,N_6920);
or U7099 (N_7099,N_6906,N_6514);
nand U7100 (N_7100,N_6917,N_6678);
nor U7101 (N_7101,N_6631,N_6924);
and U7102 (N_7102,N_6802,N_6639);
nand U7103 (N_7103,N_6907,N_6569);
nor U7104 (N_7104,N_6733,N_6711);
and U7105 (N_7105,N_6841,N_6535);
nand U7106 (N_7106,N_6664,N_6709);
or U7107 (N_7107,N_6740,N_6910);
and U7108 (N_7108,N_6600,N_6810);
nand U7109 (N_7109,N_6632,N_6814);
and U7110 (N_7110,N_6681,N_6705);
nand U7111 (N_7111,N_6798,N_6694);
nand U7112 (N_7112,N_6689,N_6918);
or U7113 (N_7113,N_6521,N_6916);
or U7114 (N_7114,N_6731,N_6855);
and U7115 (N_7115,N_6822,N_6809);
nor U7116 (N_7116,N_6779,N_6871);
nand U7117 (N_7117,N_6577,N_6593);
or U7118 (N_7118,N_6826,N_6663);
or U7119 (N_7119,N_6858,N_6760);
xnor U7120 (N_7120,N_6671,N_6539);
or U7121 (N_7121,N_6954,N_6915);
nand U7122 (N_7122,N_6712,N_6851);
and U7123 (N_7123,N_6902,N_6617);
or U7124 (N_7124,N_6867,N_6520);
or U7125 (N_7125,N_6881,N_6965);
nand U7126 (N_7126,N_6789,N_6538);
xnor U7127 (N_7127,N_6776,N_6981);
nor U7128 (N_7128,N_6548,N_6532);
nor U7129 (N_7129,N_6601,N_6537);
and U7130 (N_7130,N_6919,N_6992);
xor U7131 (N_7131,N_6847,N_6827);
nor U7132 (N_7132,N_6921,N_6772);
nor U7133 (N_7133,N_6968,N_6734);
and U7134 (N_7134,N_6904,N_6807);
nor U7135 (N_7135,N_6542,N_6623);
nand U7136 (N_7136,N_6959,N_6605);
nor U7137 (N_7137,N_6633,N_6679);
and U7138 (N_7138,N_6771,N_6693);
nand U7139 (N_7139,N_6713,N_6945);
nor U7140 (N_7140,N_6565,N_6964);
and U7141 (N_7141,N_6643,N_6913);
nand U7142 (N_7142,N_6844,N_6777);
nand U7143 (N_7143,N_6662,N_6583);
nor U7144 (N_7144,N_6934,N_6935);
nor U7145 (N_7145,N_6840,N_6853);
and U7146 (N_7146,N_6524,N_6610);
nor U7147 (N_7147,N_6523,N_6888);
or U7148 (N_7148,N_6672,N_6658);
or U7149 (N_7149,N_6896,N_6784);
or U7150 (N_7150,N_6790,N_6510);
xnor U7151 (N_7151,N_6596,N_6762);
xor U7152 (N_7152,N_6848,N_6922);
or U7153 (N_7153,N_6747,N_6843);
nor U7154 (N_7154,N_6568,N_6890);
nor U7155 (N_7155,N_6878,N_6803);
nand U7156 (N_7156,N_6833,N_6986);
or U7157 (N_7157,N_6591,N_6937);
and U7158 (N_7158,N_6883,N_6613);
and U7159 (N_7159,N_6686,N_6676);
and U7160 (N_7160,N_6999,N_6563);
xor U7161 (N_7161,N_6547,N_6719);
nor U7162 (N_7162,N_6698,N_6797);
nand U7163 (N_7163,N_6929,N_6953);
and U7164 (N_7164,N_6788,N_6630);
and U7165 (N_7165,N_6564,N_6574);
or U7166 (N_7166,N_6507,N_6675);
and U7167 (N_7167,N_6501,N_6650);
nand U7168 (N_7168,N_6866,N_6962);
nor U7169 (N_7169,N_6692,N_6557);
nor U7170 (N_7170,N_6980,N_6998);
xnor U7171 (N_7171,N_6983,N_6877);
nor U7172 (N_7172,N_6652,N_6949);
or U7173 (N_7173,N_6817,N_6533);
or U7174 (N_7174,N_6667,N_6849);
and U7175 (N_7175,N_6838,N_6975);
and U7176 (N_7176,N_6602,N_6710);
and U7177 (N_7177,N_6769,N_6570);
or U7178 (N_7178,N_6506,N_6730);
and U7179 (N_7179,N_6553,N_6792);
or U7180 (N_7180,N_6513,N_6546);
or U7181 (N_7181,N_6863,N_6616);
or U7182 (N_7182,N_6749,N_6531);
nor U7183 (N_7183,N_6530,N_6870);
and U7184 (N_7184,N_6576,N_6739);
xnor U7185 (N_7185,N_6957,N_6941);
nand U7186 (N_7186,N_6961,N_6894);
and U7187 (N_7187,N_6759,N_6869);
nor U7188 (N_7188,N_6823,N_6627);
nor U7189 (N_7189,N_6971,N_6854);
nand U7190 (N_7190,N_6943,N_6636);
and U7191 (N_7191,N_6621,N_6806);
xnor U7192 (N_7192,N_6874,N_6956);
nor U7193 (N_7193,N_6579,N_6646);
nor U7194 (N_7194,N_6781,N_6737);
nor U7195 (N_7195,N_6753,N_6808);
xor U7196 (N_7196,N_6994,N_6952);
and U7197 (N_7197,N_6895,N_6536);
or U7198 (N_7198,N_6625,N_6939);
nor U7199 (N_7199,N_6661,N_6991);
and U7200 (N_7200,N_6860,N_6990);
and U7201 (N_7201,N_6670,N_6914);
and U7202 (N_7202,N_6584,N_6876);
or U7203 (N_7203,N_6638,N_6608);
or U7204 (N_7204,N_6606,N_6832);
or U7205 (N_7205,N_6644,N_6829);
or U7206 (N_7206,N_6587,N_6634);
and U7207 (N_7207,N_6842,N_6604);
nand U7208 (N_7208,N_6573,N_6800);
or U7209 (N_7209,N_6720,N_6647);
xor U7210 (N_7210,N_6886,N_6505);
nor U7211 (N_7211,N_6723,N_6649);
xor U7212 (N_7212,N_6512,N_6763);
and U7213 (N_7213,N_6566,N_6572);
or U7214 (N_7214,N_6550,N_6722);
nor U7215 (N_7215,N_6752,N_6738);
and U7216 (N_7216,N_6718,N_6900);
and U7217 (N_7217,N_6549,N_6815);
xnor U7218 (N_7218,N_6996,N_6795);
nand U7219 (N_7219,N_6865,N_6850);
nand U7220 (N_7220,N_6758,N_6884);
nor U7221 (N_7221,N_6684,N_6715);
nand U7222 (N_7222,N_6687,N_6560);
nor U7223 (N_7223,N_6931,N_6669);
nor U7224 (N_7224,N_6511,N_6615);
nand U7225 (N_7225,N_6708,N_6561);
and U7226 (N_7226,N_6932,N_6927);
nor U7227 (N_7227,N_6586,N_6765);
and U7228 (N_7228,N_6799,N_6862);
xnor U7229 (N_7229,N_6582,N_6767);
nor U7230 (N_7230,N_6946,N_6947);
xor U7231 (N_7231,N_6930,N_6746);
nor U7232 (N_7232,N_6796,N_6972);
xnor U7233 (N_7233,N_6976,N_6977);
or U7234 (N_7234,N_6889,N_6950);
nand U7235 (N_7235,N_6543,N_6699);
and U7236 (N_7236,N_6936,N_6967);
xnor U7237 (N_7237,N_6852,N_6555);
nor U7238 (N_7238,N_6824,N_6816);
or U7239 (N_7239,N_6592,N_6700);
or U7240 (N_7240,N_6703,N_6509);
nand U7241 (N_7241,N_6969,N_6756);
or U7242 (N_7242,N_6787,N_6655);
xor U7243 (N_7243,N_6502,N_6875);
nand U7244 (N_7244,N_6785,N_6942);
nor U7245 (N_7245,N_6791,N_6970);
or U7246 (N_7246,N_6614,N_6642);
nand U7247 (N_7247,N_6804,N_6744);
nor U7248 (N_7248,N_6812,N_6707);
and U7249 (N_7249,N_6685,N_6973);
or U7250 (N_7250,N_6901,N_6714);
or U7251 (N_7251,N_6706,N_6548);
nor U7252 (N_7252,N_6980,N_6600);
xor U7253 (N_7253,N_6555,N_6573);
and U7254 (N_7254,N_6726,N_6540);
nand U7255 (N_7255,N_6566,N_6800);
nand U7256 (N_7256,N_6936,N_6648);
nand U7257 (N_7257,N_6768,N_6664);
or U7258 (N_7258,N_6667,N_6701);
or U7259 (N_7259,N_6532,N_6950);
nor U7260 (N_7260,N_6846,N_6546);
nand U7261 (N_7261,N_6578,N_6884);
nor U7262 (N_7262,N_6976,N_6988);
nor U7263 (N_7263,N_6908,N_6517);
nor U7264 (N_7264,N_6783,N_6926);
xnor U7265 (N_7265,N_6594,N_6796);
and U7266 (N_7266,N_6771,N_6627);
nor U7267 (N_7267,N_6969,N_6741);
nor U7268 (N_7268,N_6961,N_6633);
nand U7269 (N_7269,N_6633,N_6660);
and U7270 (N_7270,N_6636,N_6649);
or U7271 (N_7271,N_6741,N_6584);
or U7272 (N_7272,N_6803,N_6747);
and U7273 (N_7273,N_6669,N_6844);
nand U7274 (N_7274,N_6996,N_6572);
or U7275 (N_7275,N_6964,N_6817);
and U7276 (N_7276,N_6831,N_6995);
and U7277 (N_7277,N_6773,N_6506);
or U7278 (N_7278,N_6699,N_6773);
nand U7279 (N_7279,N_6651,N_6839);
and U7280 (N_7280,N_6701,N_6646);
xor U7281 (N_7281,N_6868,N_6956);
or U7282 (N_7282,N_6534,N_6986);
nand U7283 (N_7283,N_6580,N_6756);
or U7284 (N_7284,N_6784,N_6652);
nor U7285 (N_7285,N_6879,N_6798);
nand U7286 (N_7286,N_6620,N_6592);
and U7287 (N_7287,N_6722,N_6968);
and U7288 (N_7288,N_6563,N_6826);
or U7289 (N_7289,N_6872,N_6625);
and U7290 (N_7290,N_6822,N_6760);
and U7291 (N_7291,N_6901,N_6638);
xor U7292 (N_7292,N_6810,N_6844);
and U7293 (N_7293,N_6586,N_6632);
and U7294 (N_7294,N_6931,N_6920);
or U7295 (N_7295,N_6815,N_6994);
nor U7296 (N_7296,N_6929,N_6550);
and U7297 (N_7297,N_6843,N_6680);
or U7298 (N_7298,N_6878,N_6986);
nand U7299 (N_7299,N_6928,N_6830);
and U7300 (N_7300,N_6879,N_6728);
and U7301 (N_7301,N_6564,N_6606);
nor U7302 (N_7302,N_6508,N_6558);
or U7303 (N_7303,N_6956,N_6542);
or U7304 (N_7304,N_6996,N_6665);
or U7305 (N_7305,N_6700,N_6556);
and U7306 (N_7306,N_6842,N_6968);
or U7307 (N_7307,N_6517,N_6543);
xnor U7308 (N_7308,N_6556,N_6619);
or U7309 (N_7309,N_6549,N_6921);
nand U7310 (N_7310,N_6557,N_6940);
and U7311 (N_7311,N_6995,N_6928);
and U7312 (N_7312,N_6746,N_6618);
and U7313 (N_7313,N_6647,N_6548);
nand U7314 (N_7314,N_6636,N_6752);
and U7315 (N_7315,N_6842,N_6865);
or U7316 (N_7316,N_6812,N_6685);
nand U7317 (N_7317,N_6646,N_6501);
or U7318 (N_7318,N_6783,N_6962);
nor U7319 (N_7319,N_6815,N_6769);
nor U7320 (N_7320,N_6694,N_6625);
nor U7321 (N_7321,N_6873,N_6697);
nor U7322 (N_7322,N_6541,N_6565);
nand U7323 (N_7323,N_6597,N_6891);
nor U7324 (N_7324,N_6831,N_6981);
and U7325 (N_7325,N_6790,N_6957);
nor U7326 (N_7326,N_6893,N_6639);
nor U7327 (N_7327,N_6968,N_6880);
or U7328 (N_7328,N_6893,N_6552);
and U7329 (N_7329,N_6773,N_6693);
nand U7330 (N_7330,N_6594,N_6863);
nor U7331 (N_7331,N_6579,N_6753);
xor U7332 (N_7332,N_6812,N_6598);
and U7333 (N_7333,N_6565,N_6683);
nor U7334 (N_7334,N_6547,N_6693);
or U7335 (N_7335,N_6563,N_6873);
nor U7336 (N_7336,N_6826,N_6787);
nand U7337 (N_7337,N_6604,N_6925);
and U7338 (N_7338,N_6601,N_6776);
xor U7339 (N_7339,N_6644,N_6857);
nor U7340 (N_7340,N_6917,N_6832);
nand U7341 (N_7341,N_6682,N_6933);
or U7342 (N_7342,N_6860,N_6576);
nand U7343 (N_7343,N_6500,N_6606);
nand U7344 (N_7344,N_6900,N_6869);
xor U7345 (N_7345,N_6623,N_6740);
nor U7346 (N_7346,N_6531,N_6985);
xnor U7347 (N_7347,N_6788,N_6938);
or U7348 (N_7348,N_6502,N_6665);
or U7349 (N_7349,N_6501,N_6537);
nor U7350 (N_7350,N_6625,N_6596);
or U7351 (N_7351,N_6923,N_6537);
or U7352 (N_7352,N_6706,N_6536);
or U7353 (N_7353,N_6726,N_6707);
and U7354 (N_7354,N_6673,N_6754);
and U7355 (N_7355,N_6583,N_6825);
nor U7356 (N_7356,N_6738,N_6970);
xor U7357 (N_7357,N_6591,N_6715);
or U7358 (N_7358,N_6566,N_6957);
and U7359 (N_7359,N_6706,N_6500);
nand U7360 (N_7360,N_6968,N_6583);
or U7361 (N_7361,N_6685,N_6713);
or U7362 (N_7362,N_6990,N_6861);
or U7363 (N_7363,N_6739,N_6728);
and U7364 (N_7364,N_6548,N_6745);
nand U7365 (N_7365,N_6929,N_6642);
nor U7366 (N_7366,N_6937,N_6915);
or U7367 (N_7367,N_6648,N_6963);
or U7368 (N_7368,N_6897,N_6809);
xor U7369 (N_7369,N_6627,N_6866);
or U7370 (N_7370,N_6514,N_6798);
and U7371 (N_7371,N_6981,N_6900);
and U7372 (N_7372,N_6542,N_6568);
and U7373 (N_7373,N_6699,N_6907);
or U7374 (N_7374,N_6524,N_6853);
and U7375 (N_7375,N_6896,N_6731);
or U7376 (N_7376,N_6755,N_6766);
and U7377 (N_7377,N_6820,N_6812);
xor U7378 (N_7378,N_6681,N_6805);
and U7379 (N_7379,N_6995,N_6596);
nand U7380 (N_7380,N_6523,N_6907);
and U7381 (N_7381,N_6864,N_6852);
xor U7382 (N_7382,N_6813,N_6710);
nand U7383 (N_7383,N_6901,N_6899);
nand U7384 (N_7384,N_6765,N_6616);
and U7385 (N_7385,N_6848,N_6775);
or U7386 (N_7386,N_6607,N_6828);
nand U7387 (N_7387,N_6921,N_6500);
xnor U7388 (N_7388,N_6891,N_6884);
nor U7389 (N_7389,N_6810,N_6769);
or U7390 (N_7390,N_6791,N_6648);
and U7391 (N_7391,N_6671,N_6581);
and U7392 (N_7392,N_6855,N_6994);
and U7393 (N_7393,N_6922,N_6519);
and U7394 (N_7394,N_6832,N_6823);
nand U7395 (N_7395,N_6688,N_6775);
nand U7396 (N_7396,N_6689,N_6820);
xor U7397 (N_7397,N_6793,N_6976);
nand U7398 (N_7398,N_6655,N_6975);
and U7399 (N_7399,N_6611,N_6852);
nor U7400 (N_7400,N_6634,N_6807);
nor U7401 (N_7401,N_6993,N_6596);
nand U7402 (N_7402,N_6912,N_6616);
nand U7403 (N_7403,N_6871,N_6898);
xor U7404 (N_7404,N_6666,N_6742);
nand U7405 (N_7405,N_6790,N_6741);
and U7406 (N_7406,N_6796,N_6988);
xor U7407 (N_7407,N_6701,N_6612);
and U7408 (N_7408,N_6744,N_6940);
nand U7409 (N_7409,N_6796,N_6695);
nor U7410 (N_7410,N_6697,N_6916);
nor U7411 (N_7411,N_6504,N_6819);
or U7412 (N_7412,N_6657,N_6764);
nand U7413 (N_7413,N_6729,N_6740);
or U7414 (N_7414,N_6638,N_6758);
nand U7415 (N_7415,N_6743,N_6757);
nor U7416 (N_7416,N_6521,N_6973);
or U7417 (N_7417,N_6707,N_6798);
or U7418 (N_7418,N_6763,N_6533);
or U7419 (N_7419,N_6526,N_6888);
nor U7420 (N_7420,N_6634,N_6769);
or U7421 (N_7421,N_6710,N_6504);
and U7422 (N_7422,N_6736,N_6991);
nand U7423 (N_7423,N_6534,N_6731);
and U7424 (N_7424,N_6779,N_6700);
nor U7425 (N_7425,N_6581,N_6646);
and U7426 (N_7426,N_6795,N_6583);
and U7427 (N_7427,N_6628,N_6584);
or U7428 (N_7428,N_6836,N_6598);
nor U7429 (N_7429,N_6924,N_6933);
nand U7430 (N_7430,N_6934,N_6766);
or U7431 (N_7431,N_6712,N_6726);
and U7432 (N_7432,N_6809,N_6522);
nand U7433 (N_7433,N_6587,N_6972);
and U7434 (N_7434,N_6514,N_6664);
nand U7435 (N_7435,N_6650,N_6569);
nor U7436 (N_7436,N_6556,N_6867);
nor U7437 (N_7437,N_6661,N_6663);
nand U7438 (N_7438,N_6758,N_6702);
and U7439 (N_7439,N_6571,N_6521);
and U7440 (N_7440,N_6857,N_6839);
or U7441 (N_7441,N_6540,N_6705);
and U7442 (N_7442,N_6606,N_6712);
nand U7443 (N_7443,N_6909,N_6787);
xnor U7444 (N_7444,N_6570,N_6904);
or U7445 (N_7445,N_6703,N_6845);
and U7446 (N_7446,N_6695,N_6696);
nand U7447 (N_7447,N_6899,N_6645);
and U7448 (N_7448,N_6727,N_6788);
or U7449 (N_7449,N_6765,N_6678);
and U7450 (N_7450,N_6878,N_6576);
xnor U7451 (N_7451,N_6584,N_6956);
or U7452 (N_7452,N_6716,N_6857);
nand U7453 (N_7453,N_6524,N_6586);
and U7454 (N_7454,N_6505,N_6744);
or U7455 (N_7455,N_6586,N_6791);
and U7456 (N_7456,N_6527,N_6587);
and U7457 (N_7457,N_6763,N_6570);
xnor U7458 (N_7458,N_6813,N_6625);
and U7459 (N_7459,N_6691,N_6725);
or U7460 (N_7460,N_6796,N_6861);
xor U7461 (N_7461,N_6519,N_6878);
or U7462 (N_7462,N_6608,N_6637);
nand U7463 (N_7463,N_6856,N_6619);
and U7464 (N_7464,N_6557,N_6894);
nor U7465 (N_7465,N_6839,N_6962);
nand U7466 (N_7466,N_6926,N_6941);
or U7467 (N_7467,N_6678,N_6554);
nand U7468 (N_7468,N_6528,N_6936);
nand U7469 (N_7469,N_6667,N_6774);
and U7470 (N_7470,N_6981,N_6606);
nor U7471 (N_7471,N_6651,N_6623);
and U7472 (N_7472,N_6598,N_6881);
nand U7473 (N_7473,N_6946,N_6838);
or U7474 (N_7474,N_6908,N_6783);
and U7475 (N_7475,N_6845,N_6555);
or U7476 (N_7476,N_6527,N_6713);
nor U7477 (N_7477,N_6668,N_6597);
xnor U7478 (N_7478,N_6918,N_6676);
nor U7479 (N_7479,N_6986,N_6796);
and U7480 (N_7480,N_6923,N_6967);
xor U7481 (N_7481,N_6692,N_6879);
nor U7482 (N_7482,N_6701,N_6885);
nand U7483 (N_7483,N_6758,N_6828);
or U7484 (N_7484,N_6937,N_6699);
nor U7485 (N_7485,N_6704,N_6998);
nor U7486 (N_7486,N_6663,N_6709);
or U7487 (N_7487,N_6839,N_6611);
nand U7488 (N_7488,N_6871,N_6550);
nand U7489 (N_7489,N_6984,N_6941);
or U7490 (N_7490,N_6897,N_6590);
and U7491 (N_7491,N_6524,N_6879);
nand U7492 (N_7492,N_6607,N_6891);
and U7493 (N_7493,N_6628,N_6535);
and U7494 (N_7494,N_6500,N_6822);
or U7495 (N_7495,N_6643,N_6977);
xor U7496 (N_7496,N_6760,N_6743);
nand U7497 (N_7497,N_6670,N_6604);
and U7498 (N_7498,N_6817,N_6951);
and U7499 (N_7499,N_6999,N_6597);
and U7500 (N_7500,N_7247,N_7073);
and U7501 (N_7501,N_7477,N_7392);
and U7502 (N_7502,N_7099,N_7343);
and U7503 (N_7503,N_7316,N_7461);
xor U7504 (N_7504,N_7386,N_7165);
and U7505 (N_7505,N_7304,N_7267);
or U7506 (N_7506,N_7107,N_7375);
nand U7507 (N_7507,N_7434,N_7041);
nand U7508 (N_7508,N_7078,N_7359);
nand U7509 (N_7509,N_7429,N_7408);
nor U7510 (N_7510,N_7032,N_7416);
xor U7511 (N_7511,N_7398,N_7120);
or U7512 (N_7512,N_7478,N_7224);
nor U7513 (N_7513,N_7132,N_7308);
and U7514 (N_7514,N_7123,N_7001);
or U7515 (N_7515,N_7288,N_7468);
or U7516 (N_7516,N_7136,N_7455);
and U7517 (N_7517,N_7028,N_7020);
nand U7518 (N_7518,N_7071,N_7108);
and U7519 (N_7519,N_7184,N_7457);
and U7520 (N_7520,N_7122,N_7371);
xor U7521 (N_7521,N_7105,N_7109);
nor U7522 (N_7522,N_7326,N_7131);
nor U7523 (N_7523,N_7412,N_7365);
nor U7524 (N_7524,N_7005,N_7250);
nor U7525 (N_7525,N_7027,N_7066);
nand U7526 (N_7526,N_7315,N_7232);
or U7527 (N_7527,N_7060,N_7300);
and U7528 (N_7528,N_7160,N_7202);
and U7529 (N_7529,N_7355,N_7294);
nand U7530 (N_7530,N_7460,N_7007);
and U7531 (N_7531,N_7114,N_7469);
and U7532 (N_7532,N_7410,N_7113);
or U7533 (N_7533,N_7401,N_7072);
and U7534 (N_7534,N_7104,N_7443);
and U7535 (N_7535,N_7257,N_7427);
and U7536 (N_7536,N_7253,N_7038);
nor U7537 (N_7537,N_7498,N_7481);
nand U7538 (N_7538,N_7144,N_7342);
and U7539 (N_7539,N_7018,N_7210);
nand U7540 (N_7540,N_7459,N_7097);
and U7541 (N_7541,N_7065,N_7413);
nand U7542 (N_7542,N_7264,N_7360);
and U7543 (N_7543,N_7220,N_7391);
or U7544 (N_7544,N_7050,N_7118);
or U7545 (N_7545,N_7023,N_7083);
or U7546 (N_7546,N_7182,N_7130);
nand U7547 (N_7547,N_7381,N_7228);
nand U7548 (N_7548,N_7274,N_7008);
nor U7549 (N_7549,N_7011,N_7336);
nor U7550 (N_7550,N_7062,N_7035);
nand U7551 (N_7551,N_7317,N_7396);
or U7552 (N_7552,N_7252,N_7111);
nor U7553 (N_7553,N_7075,N_7465);
xor U7554 (N_7554,N_7306,N_7179);
and U7555 (N_7555,N_7070,N_7205);
and U7556 (N_7556,N_7081,N_7019);
xnor U7557 (N_7557,N_7263,N_7140);
and U7558 (N_7558,N_7289,N_7048);
or U7559 (N_7559,N_7320,N_7004);
nor U7560 (N_7560,N_7311,N_7246);
xnor U7561 (N_7561,N_7026,N_7482);
nor U7562 (N_7562,N_7353,N_7170);
or U7563 (N_7563,N_7142,N_7128);
or U7564 (N_7564,N_7159,N_7098);
nand U7565 (N_7565,N_7185,N_7363);
and U7566 (N_7566,N_7248,N_7080);
nand U7567 (N_7567,N_7162,N_7152);
and U7568 (N_7568,N_7373,N_7467);
or U7569 (N_7569,N_7287,N_7233);
nand U7570 (N_7570,N_7370,N_7197);
or U7571 (N_7571,N_7271,N_7053);
or U7572 (N_7572,N_7280,N_7454);
xnor U7573 (N_7573,N_7096,N_7422);
nand U7574 (N_7574,N_7446,N_7219);
nand U7575 (N_7575,N_7421,N_7329);
and U7576 (N_7576,N_7056,N_7237);
or U7577 (N_7577,N_7453,N_7243);
and U7578 (N_7578,N_7439,N_7217);
nand U7579 (N_7579,N_7172,N_7221);
nand U7580 (N_7580,N_7307,N_7334);
and U7581 (N_7581,N_7196,N_7497);
and U7582 (N_7582,N_7013,N_7442);
or U7583 (N_7583,N_7192,N_7082);
or U7584 (N_7584,N_7338,N_7054);
or U7585 (N_7585,N_7193,N_7333);
or U7586 (N_7586,N_7494,N_7174);
or U7587 (N_7587,N_7201,N_7324);
and U7588 (N_7588,N_7323,N_7110);
nand U7589 (N_7589,N_7225,N_7181);
nor U7590 (N_7590,N_7423,N_7068);
nor U7591 (N_7591,N_7278,N_7012);
or U7592 (N_7592,N_7491,N_7010);
and U7593 (N_7593,N_7437,N_7088);
or U7594 (N_7594,N_7094,N_7043);
xnor U7595 (N_7595,N_7244,N_7402);
nor U7596 (N_7596,N_7332,N_7474);
nor U7597 (N_7597,N_7156,N_7015);
or U7598 (N_7598,N_7450,N_7095);
nand U7599 (N_7599,N_7258,N_7266);
nand U7600 (N_7600,N_7039,N_7090);
and U7601 (N_7601,N_7417,N_7490);
nand U7602 (N_7602,N_7403,N_7178);
xor U7603 (N_7603,N_7480,N_7470);
and U7604 (N_7604,N_7021,N_7379);
xnor U7605 (N_7605,N_7061,N_7029);
nand U7606 (N_7606,N_7362,N_7321);
and U7607 (N_7607,N_7387,N_7199);
and U7608 (N_7608,N_7229,N_7414);
nand U7609 (N_7609,N_7301,N_7223);
or U7610 (N_7610,N_7030,N_7276);
xnor U7611 (N_7611,N_7431,N_7003);
or U7612 (N_7612,N_7125,N_7489);
nor U7613 (N_7613,N_7102,N_7286);
xnor U7614 (N_7614,N_7238,N_7269);
nor U7615 (N_7615,N_7433,N_7485);
nand U7616 (N_7616,N_7380,N_7337);
or U7617 (N_7617,N_7153,N_7372);
and U7618 (N_7618,N_7124,N_7231);
nand U7619 (N_7619,N_7218,N_7022);
or U7620 (N_7620,N_7495,N_7426);
or U7621 (N_7621,N_7283,N_7149);
and U7622 (N_7622,N_7399,N_7420);
and U7623 (N_7623,N_7309,N_7214);
nand U7624 (N_7624,N_7240,N_7087);
or U7625 (N_7625,N_7313,N_7499);
nand U7626 (N_7626,N_7348,N_7395);
or U7627 (N_7627,N_7055,N_7116);
or U7628 (N_7628,N_7374,N_7031);
or U7629 (N_7629,N_7037,N_7212);
and U7630 (N_7630,N_7345,N_7121);
nand U7631 (N_7631,N_7471,N_7208);
and U7632 (N_7632,N_7441,N_7077);
nor U7633 (N_7633,N_7188,N_7298);
nand U7634 (N_7634,N_7305,N_7206);
nand U7635 (N_7635,N_7361,N_7394);
or U7636 (N_7636,N_7261,N_7358);
nor U7637 (N_7637,N_7173,N_7473);
nor U7638 (N_7638,N_7262,N_7052);
or U7639 (N_7639,N_7302,N_7167);
or U7640 (N_7640,N_7466,N_7168);
nor U7641 (N_7641,N_7259,N_7195);
and U7642 (N_7642,N_7133,N_7346);
or U7643 (N_7643,N_7002,N_7135);
or U7644 (N_7644,N_7046,N_7207);
xnor U7645 (N_7645,N_7049,N_7452);
and U7646 (N_7646,N_7175,N_7384);
nand U7647 (N_7647,N_7166,N_7484);
nor U7648 (N_7648,N_7150,N_7293);
nor U7649 (N_7649,N_7155,N_7356);
xor U7650 (N_7650,N_7369,N_7444);
or U7651 (N_7651,N_7295,N_7024);
and U7652 (N_7652,N_7273,N_7322);
xnor U7653 (N_7653,N_7045,N_7047);
xor U7654 (N_7654,N_7376,N_7312);
xnor U7655 (N_7655,N_7245,N_7319);
nand U7656 (N_7656,N_7180,N_7138);
and U7657 (N_7657,N_7407,N_7009);
and U7658 (N_7658,N_7227,N_7169);
xnor U7659 (N_7659,N_7079,N_7239);
nor U7660 (N_7660,N_7101,N_7487);
and U7661 (N_7661,N_7328,N_7445);
nor U7662 (N_7662,N_7260,N_7255);
or U7663 (N_7663,N_7479,N_7222);
nand U7664 (N_7664,N_7119,N_7347);
nor U7665 (N_7665,N_7000,N_7236);
nand U7666 (N_7666,N_7103,N_7241);
and U7667 (N_7667,N_7213,N_7014);
and U7668 (N_7668,N_7314,N_7230);
nor U7669 (N_7669,N_7383,N_7025);
and U7670 (N_7670,N_7406,N_7404);
nor U7671 (N_7671,N_7226,N_7488);
or U7672 (N_7672,N_7275,N_7496);
nor U7673 (N_7673,N_7017,N_7279);
and U7674 (N_7674,N_7203,N_7158);
nor U7675 (N_7675,N_7393,N_7377);
nand U7676 (N_7676,N_7451,N_7390);
xnor U7677 (N_7677,N_7378,N_7006);
nand U7678 (N_7678,N_7281,N_7388);
xnor U7679 (N_7679,N_7074,N_7117);
nor U7680 (N_7680,N_7418,N_7341);
and U7681 (N_7681,N_7299,N_7069);
xnor U7682 (N_7682,N_7325,N_7187);
or U7683 (N_7683,N_7351,N_7335);
or U7684 (N_7684,N_7303,N_7190);
and U7685 (N_7685,N_7349,N_7063);
and U7686 (N_7686,N_7235,N_7164);
nor U7687 (N_7687,N_7285,N_7424);
and U7688 (N_7688,N_7146,N_7492);
nand U7689 (N_7689,N_7330,N_7141);
nor U7690 (N_7690,N_7076,N_7493);
nor U7691 (N_7691,N_7089,N_7216);
and U7692 (N_7692,N_7112,N_7157);
xnor U7693 (N_7693,N_7297,N_7486);
and U7694 (N_7694,N_7191,N_7448);
and U7695 (N_7695,N_7134,N_7389);
nor U7696 (N_7696,N_7292,N_7145);
nor U7697 (N_7697,N_7093,N_7367);
nand U7698 (N_7698,N_7483,N_7476);
and U7699 (N_7699,N_7344,N_7400);
xnor U7700 (N_7700,N_7215,N_7154);
and U7701 (N_7701,N_7475,N_7129);
or U7702 (N_7702,N_7463,N_7058);
or U7703 (N_7703,N_7409,N_7171);
and U7704 (N_7704,N_7251,N_7318);
nand U7705 (N_7705,N_7234,N_7051);
xor U7706 (N_7706,N_7368,N_7428);
nor U7707 (N_7707,N_7354,N_7447);
or U7708 (N_7708,N_7242,N_7091);
nand U7709 (N_7709,N_7127,N_7148);
xor U7710 (N_7710,N_7397,N_7456);
xnor U7711 (N_7711,N_7382,N_7067);
nand U7712 (N_7712,N_7357,N_7270);
nand U7713 (N_7713,N_7339,N_7265);
xnor U7714 (N_7714,N_7290,N_7411);
nor U7715 (N_7715,N_7189,N_7064);
nand U7716 (N_7716,N_7143,N_7183);
and U7717 (N_7717,N_7438,N_7115);
and U7718 (N_7718,N_7291,N_7163);
and U7719 (N_7719,N_7415,N_7435);
and U7720 (N_7720,N_7432,N_7186);
or U7721 (N_7721,N_7352,N_7209);
and U7722 (N_7722,N_7310,N_7044);
nor U7723 (N_7723,N_7364,N_7092);
xnor U7724 (N_7724,N_7327,N_7198);
or U7725 (N_7725,N_7425,N_7161);
nand U7726 (N_7726,N_7272,N_7204);
and U7727 (N_7727,N_7059,N_7385);
nand U7728 (N_7728,N_7268,N_7033);
nand U7729 (N_7729,N_7458,N_7177);
nand U7730 (N_7730,N_7350,N_7256);
or U7731 (N_7731,N_7211,N_7036);
and U7732 (N_7732,N_7151,N_7126);
nand U7733 (N_7733,N_7084,N_7086);
or U7734 (N_7734,N_7331,N_7137);
nand U7735 (N_7735,N_7200,N_7282);
or U7736 (N_7736,N_7464,N_7462);
and U7737 (N_7737,N_7284,N_7472);
nand U7738 (N_7738,N_7042,N_7436);
and U7739 (N_7739,N_7106,N_7340);
or U7740 (N_7740,N_7085,N_7194);
xor U7741 (N_7741,N_7366,N_7296);
xor U7742 (N_7742,N_7440,N_7139);
or U7743 (N_7743,N_7057,N_7254);
and U7744 (N_7744,N_7147,N_7016);
nand U7745 (N_7745,N_7249,N_7034);
or U7746 (N_7746,N_7449,N_7419);
and U7747 (N_7747,N_7277,N_7100);
or U7748 (N_7748,N_7040,N_7176);
and U7749 (N_7749,N_7405,N_7430);
or U7750 (N_7750,N_7196,N_7477);
or U7751 (N_7751,N_7147,N_7056);
or U7752 (N_7752,N_7184,N_7396);
nand U7753 (N_7753,N_7373,N_7254);
nand U7754 (N_7754,N_7484,N_7174);
xnor U7755 (N_7755,N_7446,N_7019);
nand U7756 (N_7756,N_7068,N_7039);
and U7757 (N_7757,N_7450,N_7280);
and U7758 (N_7758,N_7167,N_7362);
nand U7759 (N_7759,N_7408,N_7224);
nand U7760 (N_7760,N_7327,N_7498);
or U7761 (N_7761,N_7150,N_7257);
nand U7762 (N_7762,N_7107,N_7358);
nand U7763 (N_7763,N_7264,N_7326);
xnor U7764 (N_7764,N_7403,N_7275);
or U7765 (N_7765,N_7251,N_7454);
or U7766 (N_7766,N_7203,N_7084);
or U7767 (N_7767,N_7443,N_7209);
nor U7768 (N_7768,N_7438,N_7389);
nor U7769 (N_7769,N_7127,N_7173);
and U7770 (N_7770,N_7035,N_7370);
nor U7771 (N_7771,N_7078,N_7039);
nor U7772 (N_7772,N_7424,N_7024);
or U7773 (N_7773,N_7077,N_7150);
nor U7774 (N_7774,N_7149,N_7005);
xor U7775 (N_7775,N_7300,N_7489);
nand U7776 (N_7776,N_7335,N_7198);
and U7777 (N_7777,N_7421,N_7308);
nand U7778 (N_7778,N_7258,N_7341);
or U7779 (N_7779,N_7010,N_7100);
and U7780 (N_7780,N_7245,N_7042);
and U7781 (N_7781,N_7003,N_7260);
nand U7782 (N_7782,N_7374,N_7403);
or U7783 (N_7783,N_7356,N_7044);
nor U7784 (N_7784,N_7137,N_7379);
or U7785 (N_7785,N_7083,N_7046);
nand U7786 (N_7786,N_7279,N_7384);
and U7787 (N_7787,N_7336,N_7306);
and U7788 (N_7788,N_7094,N_7010);
nor U7789 (N_7789,N_7347,N_7333);
nand U7790 (N_7790,N_7094,N_7458);
xnor U7791 (N_7791,N_7046,N_7429);
xnor U7792 (N_7792,N_7212,N_7393);
xor U7793 (N_7793,N_7343,N_7336);
or U7794 (N_7794,N_7034,N_7286);
xnor U7795 (N_7795,N_7491,N_7469);
or U7796 (N_7796,N_7372,N_7410);
nand U7797 (N_7797,N_7006,N_7136);
and U7798 (N_7798,N_7482,N_7213);
xor U7799 (N_7799,N_7469,N_7235);
or U7800 (N_7800,N_7293,N_7458);
or U7801 (N_7801,N_7329,N_7158);
and U7802 (N_7802,N_7064,N_7083);
and U7803 (N_7803,N_7477,N_7110);
nand U7804 (N_7804,N_7144,N_7028);
or U7805 (N_7805,N_7128,N_7401);
nor U7806 (N_7806,N_7049,N_7279);
nand U7807 (N_7807,N_7044,N_7402);
nand U7808 (N_7808,N_7424,N_7481);
or U7809 (N_7809,N_7172,N_7243);
or U7810 (N_7810,N_7001,N_7471);
or U7811 (N_7811,N_7165,N_7309);
or U7812 (N_7812,N_7001,N_7156);
xnor U7813 (N_7813,N_7437,N_7060);
nor U7814 (N_7814,N_7299,N_7371);
nor U7815 (N_7815,N_7066,N_7242);
or U7816 (N_7816,N_7133,N_7109);
and U7817 (N_7817,N_7042,N_7109);
and U7818 (N_7818,N_7292,N_7399);
or U7819 (N_7819,N_7144,N_7244);
nor U7820 (N_7820,N_7373,N_7171);
nor U7821 (N_7821,N_7076,N_7146);
xor U7822 (N_7822,N_7270,N_7264);
nor U7823 (N_7823,N_7166,N_7094);
nand U7824 (N_7824,N_7223,N_7171);
or U7825 (N_7825,N_7025,N_7449);
nand U7826 (N_7826,N_7305,N_7400);
nor U7827 (N_7827,N_7387,N_7279);
and U7828 (N_7828,N_7000,N_7222);
and U7829 (N_7829,N_7182,N_7478);
and U7830 (N_7830,N_7492,N_7142);
nor U7831 (N_7831,N_7083,N_7004);
or U7832 (N_7832,N_7492,N_7153);
nand U7833 (N_7833,N_7051,N_7313);
and U7834 (N_7834,N_7339,N_7488);
xnor U7835 (N_7835,N_7346,N_7063);
or U7836 (N_7836,N_7085,N_7049);
or U7837 (N_7837,N_7011,N_7408);
nor U7838 (N_7838,N_7394,N_7053);
nand U7839 (N_7839,N_7116,N_7222);
and U7840 (N_7840,N_7018,N_7350);
nor U7841 (N_7841,N_7278,N_7410);
and U7842 (N_7842,N_7117,N_7220);
and U7843 (N_7843,N_7357,N_7343);
or U7844 (N_7844,N_7484,N_7495);
and U7845 (N_7845,N_7359,N_7323);
and U7846 (N_7846,N_7142,N_7427);
xor U7847 (N_7847,N_7341,N_7005);
or U7848 (N_7848,N_7258,N_7157);
or U7849 (N_7849,N_7380,N_7353);
or U7850 (N_7850,N_7281,N_7413);
xnor U7851 (N_7851,N_7277,N_7011);
or U7852 (N_7852,N_7024,N_7462);
and U7853 (N_7853,N_7199,N_7085);
or U7854 (N_7854,N_7419,N_7091);
xor U7855 (N_7855,N_7385,N_7402);
nor U7856 (N_7856,N_7024,N_7282);
nor U7857 (N_7857,N_7262,N_7233);
and U7858 (N_7858,N_7279,N_7133);
or U7859 (N_7859,N_7104,N_7173);
nor U7860 (N_7860,N_7404,N_7310);
and U7861 (N_7861,N_7184,N_7085);
nor U7862 (N_7862,N_7331,N_7471);
or U7863 (N_7863,N_7268,N_7231);
nor U7864 (N_7864,N_7472,N_7160);
nor U7865 (N_7865,N_7069,N_7109);
nand U7866 (N_7866,N_7269,N_7436);
and U7867 (N_7867,N_7232,N_7201);
and U7868 (N_7868,N_7198,N_7029);
nand U7869 (N_7869,N_7296,N_7234);
nand U7870 (N_7870,N_7421,N_7420);
nor U7871 (N_7871,N_7054,N_7494);
or U7872 (N_7872,N_7213,N_7258);
and U7873 (N_7873,N_7309,N_7173);
and U7874 (N_7874,N_7016,N_7449);
and U7875 (N_7875,N_7050,N_7487);
or U7876 (N_7876,N_7232,N_7355);
xor U7877 (N_7877,N_7193,N_7297);
xnor U7878 (N_7878,N_7166,N_7474);
and U7879 (N_7879,N_7409,N_7034);
and U7880 (N_7880,N_7396,N_7221);
xnor U7881 (N_7881,N_7222,N_7168);
nor U7882 (N_7882,N_7289,N_7308);
and U7883 (N_7883,N_7304,N_7339);
nor U7884 (N_7884,N_7083,N_7300);
and U7885 (N_7885,N_7252,N_7395);
or U7886 (N_7886,N_7445,N_7313);
xnor U7887 (N_7887,N_7020,N_7111);
or U7888 (N_7888,N_7223,N_7156);
or U7889 (N_7889,N_7384,N_7047);
nand U7890 (N_7890,N_7303,N_7318);
nor U7891 (N_7891,N_7433,N_7116);
or U7892 (N_7892,N_7079,N_7063);
or U7893 (N_7893,N_7276,N_7143);
or U7894 (N_7894,N_7202,N_7142);
or U7895 (N_7895,N_7266,N_7356);
and U7896 (N_7896,N_7254,N_7324);
or U7897 (N_7897,N_7262,N_7071);
and U7898 (N_7898,N_7002,N_7424);
nor U7899 (N_7899,N_7243,N_7313);
nor U7900 (N_7900,N_7226,N_7175);
or U7901 (N_7901,N_7310,N_7131);
nor U7902 (N_7902,N_7140,N_7059);
nor U7903 (N_7903,N_7035,N_7429);
nand U7904 (N_7904,N_7199,N_7420);
nand U7905 (N_7905,N_7273,N_7438);
xor U7906 (N_7906,N_7166,N_7338);
or U7907 (N_7907,N_7431,N_7491);
xor U7908 (N_7908,N_7404,N_7319);
or U7909 (N_7909,N_7382,N_7202);
nor U7910 (N_7910,N_7476,N_7461);
nand U7911 (N_7911,N_7100,N_7014);
nor U7912 (N_7912,N_7148,N_7400);
nor U7913 (N_7913,N_7173,N_7448);
and U7914 (N_7914,N_7192,N_7007);
and U7915 (N_7915,N_7187,N_7233);
nand U7916 (N_7916,N_7410,N_7108);
xor U7917 (N_7917,N_7060,N_7483);
nor U7918 (N_7918,N_7398,N_7130);
and U7919 (N_7919,N_7026,N_7499);
nand U7920 (N_7920,N_7406,N_7401);
or U7921 (N_7921,N_7006,N_7210);
or U7922 (N_7922,N_7194,N_7042);
nand U7923 (N_7923,N_7020,N_7462);
or U7924 (N_7924,N_7316,N_7315);
nand U7925 (N_7925,N_7289,N_7187);
nand U7926 (N_7926,N_7211,N_7268);
nor U7927 (N_7927,N_7465,N_7302);
or U7928 (N_7928,N_7045,N_7239);
nor U7929 (N_7929,N_7400,N_7339);
and U7930 (N_7930,N_7111,N_7460);
nand U7931 (N_7931,N_7023,N_7251);
nand U7932 (N_7932,N_7303,N_7217);
and U7933 (N_7933,N_7275,N_7281);
nor U7934 (N_7934,N_7431,N_7080);
and U7935 (N_7935,N_7272,N_7368);
nor U7936 (N_7936,N_7104,N_7143);
nor U7937 (N_7937,N_7414,N_7165);
nor U7938 (N_7938,N_7144,N_7043);
nor U7939 (N_7939,N_7491,N_7081);
and U7940 (N_7940,N_7368,N_7396);
or U7941 (N_7941,N_7326,N_7430);
nand U7942 (N_7942,N_7494,N_7066);
nand U7943 (N_7943,N_7341,N_7404);
or U7944 (N_7944,N_7494,N_7470);
nand U7945 (N_7945,N_7416,N_7435);
or U7946 (N_7946,N_7297,N_7070);
nor U7947 (N_7947,N_7145,N_7308);
nand U7948 (N_7948,N_7182,N_7022);
nand U7949 (N_7949,N_7152,N_7316);
and U7950 (N_7950,N_7209,N_7325);
and U7951 (N_7951,N_7462,N_7324);
nor U7952 (N_7952,N_7127,N_7195);
or U7953 (N_7953,N_7303,N_7442);
xnor U7954 (N_7954,N_7383,N_7298);
or U7955 (N_7955,N_7165,N_7196);
nand U7956 (N_7956,N_7304,N_7373);
nand U7957 (N_7957,N_7013,N_7460);
and U7958 (N_7958,N_7388,N_7032);
nand U7959 (N_7959,N_7247,N_7374);
nor U7960 (N_7960,N_7481,N_7340);
and U7961 (N_7961,N_7402,N_7230);
and U7962 (N_7962,N_7011,N_7216);
xor U7963 (N_7963,N_7387,N_7312);
xor U7964 (N_7964,N_7338,N_7061);
and U7965 (N_7965,N_7160,N_7132);
nor U7966 (N_7966,N_7280,N_7366);
or U7967 (N_7967,N_7243,N_7210);
nor U7968 (N_7968,N_7013,N_7132);
and U7969 (N_7969,N_7441,N_7070);
or U7970 (N_7970,N_7350,N_7430);
nor U7971 (N_7971,N_7297,N_7183);
xor U7972 (N_7972,N_7321,N_7047);
xor U7973 (N_7973,N_7360,N_7165);
and U7974 (N_7974,N_7044,N_7113);
and U7975 (N_7975,N_7081,N_7271);
and U7976 (N_7976,N_7441,N_7244);
nand U7977 (N_7977,N_7143,N_7439);
or U7978 (N_7978,N_7472,N_7372);
nand U7979 (N_7979,N_7388,N_7022);
xnor U7980 (N_7980,N_7352,N_7215);
or U7981 (N_7981,N_7199,N_7127);
nand U7982 (N_7982,N_7457,N_7296);
nand U7983 (N_7983,N_7325,N_7073);
and U7984 (N_7984,N_7231,N_7308);
or U7985 (N_7985,N_7015,N_7190);
or U7986 (N_7986,N_7486,N_7323);
or U7987 (N_7987,N_7339,N_7014);
nand U7988 (N_7988,N_7195,N_7489);
or U7989 (N_7989,N_7203,N_7209);
or U7990 (N_7990,N_7059,N_7323);
and U7991 (N_7991,N_7005,N_7384);
nor U7992 (N_7992,N_7018,N_7399);
nand U7993 (N_7993,N_7292,N_7096);
and U7994 (N_7994,N_7169,N_7153);
xnor U7995 (N_7995,N_7463,N_7264);
nor U7996 (N_7996,N_7303,N_7469);
nor U7997 (N_7997,N_7377,N_7105);
nor U7998 (N_7998,N_7393,N_7081);
and U7999 (N_7999,N_7381,N_7236);
nor U8000 (N_8000,N_7862,N_7867);
nor U8001 (N_8001,N_7677,N_7920);
and U8002 (N_8002,N_7560,N_7797);
or U8003 (N_8003,N_7755,N_7636);
nand U8004 (N_8004,N_7539,N_7641);
nand U8005 (N_8005,N_7620,N_7937);
or U8006 (N_8006,N_7799,N_7714);
xnor U8007 (N_8007,N_7932,N_7959);
or U8008 (N_8008,N_7515,N_7971);
or U8009 (N_8009,N_7773,N_7588);
or U8010 (N_8010,N_7671,N_7617);
and U8011 (N_8011,N_7860,N_7764);
nand U8012 (N_8012,N_7553,N_7682);
xnor U8013 (N_8013,N_7520,N_7784);
nor U8014 (N_8014,N_7643,N_7698);
and U8015 (N_8015,N_7625,N_7915);
or U8016 (N_8016,N_7640,N_7606);
nand U8017 (N_8017,N_7874,N_7756);
and U8018 (N_8018,N_7908,N_7930);
or U8019 (N_8019,N_7863,N_7957);
or U8020 (N_8020,N_7523,N_7612);
or U8021 (N_8021,N_7708,N_7857);
and U8022 (N_8022,N_7995,N_7647);
nor U8023 (N_8023,N_7711,N_7751);
or U8024 (N_8024,N_7883,N_7945);
nand U8025 (N_8025,N_7557,N_7804);
or U8026 (N_8026,N_7665,N_7554);
or U8027 (N_8027,N_7549,N_7652);
or U8028 (N_8028,N_7979,N_7722);
and U8029 (N_8029,N_7526,N_7964);
and U8030 (N_8030,N_7913,N_7693);
or U8031 (N_8031,N_7833,N_7914);
and U8032 (N_8032,N_7700,N_7710);
or U8033 (N_8033,N_7603,N_7583);
xnor U8034 (N_8034,N_7534,N_7848);
or U8035 (N_8035,N_7822,N_7907);
and U8036 (N_8036,N_7731,N_7760);
nor U8037 (N_8037,N_7992,N_7840);
xor U8038 (N_8038,N_7721,N_7977);
xnor U8039 (N_8039,N_7966,N_7938);
nand U8040 (N_8040,N_7655,N_7818);
nand U8041 (N_8041,N_7841,N_7859);
or U8042 (N_8042,N_7793,N_7781);
or U8043 (N_8043,N_7690,N_7517);
nor U8044 (N_8044,N_7741,N_7631);
xnor U8045 (N_8045,N_7765,N_7947);
nand U8046 (N_8046,N_7997,N_7511);
or U8047 (N_8047,N_7856,N_7988);
and U8048 (N_8048,N_7713,N_7661);
xor U8049 (N_8049,N_7675,N_7812);
nor U8050 (N_8050,N_7839,N_7504);
and U8051 (N_8051,N_7880,N_7745);
nand U8052 (N_8052,N_7884,N_7638);
nand U8053 (N_8053,N_7969,N_7974);
nand U8054 (N_8054,N_7628,N_7686);
nor U8055 (N_8055,N_7621,N_7771);
or U8056 (N_8056,N_7658,N_7536);
xnor U8057 (N_8057,N_7524,N_7936);
nand U8058 (N_8058,N_7794,N_7775);
nand U8059 (N_8059,N_7803,N_7712);
and U8060 (N_8060,N_7593,N_7779);
nand U8061 (N_8061,N_7963,N_7587);
nand U8062 (N_8062,N_7762,N_7666);
nor U8063 (N_8063,N_7852,N_7819);
xnor U8064 (N_8064,N_7739,N_7864);
and U8065 (N_8065,N_7723,N_7895);
xnor U8066 (N_8066,N_7735,N_7843);
nand U8067 (N_8067,N_7505,N_7702);
nor U8068 (N_8068,N_7570,N_7659);
and U8069 (N_8069,N_7627,N_7733);
or U8070 (N_8070,N_7935,N_7521);
or U8071 (N_8071,N_7574,N_7673);
and U8072 (N_8072,N_7835,N_7968);
and U8073 (N_8073,N_7847,N_7949);
xor U8074 (N_8074,N_7984,N_7951);
nand U8075 (N_8075,N_7830,N_7844);
nor U8076 (N_8076,N_7663,N_7887);
and U8077 (N_8077,N_7687,N_7900);
nor U8078 (N_8078,N_7726,N_7550);
or U8079 (N_8079,N_7967,N_7858);
nand U8080 (N_8080,N_7866,N_7757);
or U8081 (N_8081,N_7566,N_7540);
and U8082 (N_8082,N_7776,N_7525);
xnor U8083 (N_8083,N_7637,N_7991);
nor U8084 (N_8084,N_7846,N_7678);
and U8085 (N_8085,N_7898,N_7611);
or U8086 (N_8086,N_7728,N_7996);
and U8087 (N_8087,N_7565,N_7507);
or U8088 (N_8088,N_7545,N_7503);
nor U8089 (N_8089,N_7704,N_7777);
nand U8090 (N_8090,N_7747,N_7934);
nor U8091 (N_8091,N_7929,N_7868);
nand U8092 (N_8092,N_7601,N_7946);
and U8093 (N_8093,N_7685,N_7890);
or U8094 (N_8094,N_7886,N_7575);
and U8095 (N_8095,N_7662,N_7944);
xnor U8096 (N_8096,N_7814,N_7811);
xnor U8097 (N_8097,N_7633,N_7985);
and U8098 (N_8098,N_7925,N_7786);
nor U8099 (N_8099,N_7933,N_7650);
and U8100 (N_8100,N_7903,N_7928);
nor U8101 (N_8101,N_7740,N_7699);
nor U8102 (N_8102,N_7902,N_7892);
and U8103 (N_8103,N_7529,N_7805);
xnor U8104 (N_8104,N_7961,N_7796);
or U8105 (N_8105,N_7990,N_7834);
or U8106 (N_8106,N_7692,N_7849);
and U8107 (N_8107,N_7761,N_7622);
nor U8108 (N_8108,N_7894,N_7873);
nor U8109 (N_8109,N_7953,N_7876);
xor U8110 (N_8110,N_7749,N_7630);
nor U8111 (N_8111,N_7897,N_7854);
or U8112 (N_8112,N_7820,N_7558);
nor U8113 (N_8113,N_7589,N_7952);
nand U8114 (N_8114,N_7580,N_7501);
or U8115 (N_8115,N_7616,N_7768);
nand U8116 (N_8116,N_7769,N_7502);
nand U8117 (N_8117,N_7832,N_7734);
nand U8118 (N_8118,N_7748,N_7905);
nand U8119 (N_8119,N_7614,N_7842);
and U8120 (N_8120,N_7660,N_7871);
nor U8121 (N_8121,N_7626,N_7861);
xnor U8122 (N_8122,N_7865,N_7998);
or U8123 (N_8123,N_7738,N_7899);
nand U8124 (N_8124,N_7569,N_7592);
or U8125 (N_8125,N_7701,N_7911);
nand U8126 (N_8126,N_7705,N_7595);
nand U8127 (N_8127,N_7831,N_7889);
nand U8128 (N_8128,N_7736,N_7885);
and U8129 (N_8129,N_7730,N_7954);
or U8130 (N_8130,N_7674,N_7596);
nand U8131 (N_8131,N_7684,N_7855);
nand U8132 (N_8132,N_7763,N_7656);
xor U8133 (N_8133,N_7958,N_7717);
nor U8134 (N_8134,N_7602,N_7535);
nor U8135 (N_8135,N_7737,N_7715);
or U8136 (N_8136,N_7870,N_7827);
and U8137 (N_8137,N_7824,N_7916);
xor U8138 (N_8138,N_7821,N_7642);
nand U8139 (N_8139,N_7670,N_7576);
xor U8140 (N_8140,N_7563,N_7879);
or U8141 (N_8141,N_7987,N_7680);
nand U8142 (N_8142,N_7853,N_7906);
and U8143 (N_8143,N_7610,N_7623);
xnor U8144 (N_8144,N_7590,N_7567);
nor U8145 (N_8145,N_7767,N_7541);
nor U8146 (N_8146,N_7970,N_7645);
or U8147 (N_8147,N_7605,N_7980);
or U8148 (N_8148,N_7882,N_7586);
and U8149 (N_8149,N_7943,N_7573);
nand U8150 (N_8150,N_7815,N_7632);
and U8151 (N_8151,N_7615,N_7836);
nor U8152 (N_8152,N_7506,N_7696);
or U8153 (N_8153,N_7624,N_7828);
nand U8154 (N_8154,N_7917,N_7518);
or U8155 (N_8155,N_7538,N_7924);
nor U8156 (N_8156,N_7759,N_7667);
nand U8157 (N_8157,N_7795,N_7551);
or U8158 (N_8158,N_7960,N_7533);
xnor U8159 (N_8159,N_7579,N_7634);
and U8160 (N_8160,N_7718,N_7694);
nand U8161 (N_8161,N_7508,N_7800);
or U8162 (N_8162,N_7644,N_7926);
nand U8163 (N_8163,N_7801,N_7510);
nand U8164 (N_8164,N_7981,N_7845);
and U8165 (N_8165,N_7901,N_7808);
nand U8166 (N_8166,N_7532,N_7672);
nor U8167 (N_8167,N_7972,N_7976);
or U8168 (N_8168,N_7921,N_7697);
and U8169 (N_8169,N_7743,N_7619);
nor U8170 (N_8170,N_7584,N_7683);
nand U8171 (N_8171,N_7531,N_7649);
and U8172 (N_8172,N_7542,N_7999);
nor U8173 (N_8173,N_7581,N_7691);
and U8174 (N_8174,N_7530,N_7823);
nor U8175 (N_8175,N_7807,N_7568);
and U8176 (N_8176,N_7802,N_7891);
and U8177 (N_8177,N_7791,N_7706);
or U8178 (N_8178,N_7594,N_7837);
xnor U8179 (N_8179,N_7552,N_7516);
nand U8180 (N_8180,N_7695,N_7774);
or U8181 (N_8181,N_7578,N_7922);
nand U8182 (N_8182,N_7613,N_7732);
nand U8183 (N_8183,N_7798,N_7597);
and U8184 (N_8184,N_7888,N_7639);
and U8185 (N_8185,N_7754,N_7746);
or U8186 (N_8186,N_7881,N_7809);
or U8187 (N_8187,N_7772,N_7782);
and U8188 (N_8188,N_7850,N_7547);
xnor U8189 (N_8189,N_7725,N_7825);
nor U8190 (N_8190,N_7522,N_7766);
nand U8191 (N_8191,N_7657,N_7544);
nor U8192 (N_8192,N_7604,N_7651);
nand U8193 (N_8193,N_7720,N_7877);
or U8194 (N_8194,N_7681,N_7543);
nor U8195 (N_8195,N_7838,N_7729);
or U8196 (N_8196,N_7648,N_7927);
nand U8197 (N_8197,N_7956,N_7572);
and U8198 (N_8198,N_7744,N_7942);
nand U8199 (N_8199,N_7975,N_7679);
and U8200 (N_8200,N_7509,N_7635);
nor U8201 (N_8201,N_7896,N_7965);
or U8202 (N_8202,N_7910,N_7556);
nand U8203 (N_8203,N_7912,N_7653);
nand U8204 (N_8204,N_7591,N_7982);
nand U8205 (N_8205,N_7582,N_7500);
or U8206 (N_8206,N_7727,N_7585);
nand U8207 (N_8207,N_7941,N_7940);
nand U8208 (N_8208,N_7555,N_7709);
nand U8209 (N_8209,N_7537,N_7703);
and U8210 (N_8210,N_7608,N_7719);
or U8211 (N_8211,N_7931,N_7826);
nor U8212 (N_8212,N_7904,N_7688);
or U8213 (N_8213,N_7778,N_7973);
nand U8214 (N_8214,N_7919,N_7571);
nor U8215 (N_8215,N_7599,N_7724);
and U8216 (N_8216,N_7546,N_7810);
nand U8217 (N_8217,N_7789,N_7548);
or U8218 (N_8218,N_7654,N_7646);
nor U8219 (N_8219,N_7955,N_7813);
and U8220 (N_8220,N_7753,N_7707);
nor U8221 (N_8221,N_7788,N_7783);
nor U8222 (N_8222,N_7689,N_7787);
nand U8223 (N_8223,N_7559,N_7607);
xnor U8224 (N_8224,N_7785,N_7918);
or U8225 (N_8225,N_7770,N_7512);
or U8226 (N_8226,N_7829,N_7939);
and U8227 (N_8227,N_7676,N_7514);
nand U8228 (N_8228,N_7869,N_7792);
nor U8229 (N_8229,N_7609,N_7780);
nor U8230 (N_8230,N_7983,N_7562);
nor U8231 (N_8231,N_7519,N_7752);
or U8232 (N_8232,N_7669,N_7716);
or U8233 (N_8233,N_7664,N_7909);
nor U8234 (N_8234,N_7993,N_7893);
and U8235 (N_8235,N_7875,N_7528);
xor U8236 (N_8236,N_7923,N_7790);
and U8237 (N_8237,N_7950,N_7806);
nor U8238 (N_8238,N_7872,N_7600);
xnor U8239 (N_8239,N_7564,N_7668);
or U8240 (N_8240,N_7978,N_7948);
nand U8241 (N_8241,N_7561,N_7878);
nand U8242 (N_8242,N_7989,N_7816);
nor U8243 (N_8243,N_7618,N_7513);
nand U8244 (N_8244,N_7962,N_7527);
nor U8245 (N_8245,N_7758,N_7629);
nand U8246 (N_8246,N_7598,N_7750);
or U8247 (N_8247,N_7577,N_7817);
nand U8248 (N_8248,N_7986,N_7742);
nor U8249 (N_8249,N_7851,N_7994);
or U8250 (N_8250,N_7585,N_7779);
and U8251 (N_8251,N_7819,N_7553);
nor U8252 (N_8252,N_7701,N_7501);
nor U8253 (N_8253,N_7657,N_7815);
and U8254 (N_8254,N_7522,N_7521);
nand U8255 (N_8255,N_7790,N_7595);
nand U8256 (N_8256,N_7884,N_7935);
and U8257 (N_8257,N_7932,N_7771);
nand U8258 (N_8258,N_7720,N_7795);
nand U8259 (N_8259,N_7771,N_7626);
nor U8260 (N_8260,N_7533,N_7815);
nor U8261 (N_8261,N_7840,N_7617);
nand U8262 (N_8262,N_7931,N_7664);
nand U8263 (N_8263,N_7785,N_7616);
nand U8264 (N_8264,N_7684,N_7613);
nand U8265 (N_8265,N_7785,N_7950);
and U8266 (N_8266,N_7970,N_7505);
or U8267 (N_8267,N_7661,N_7566);
nor U8268 (N_8268,N_7892,N_7815);
nand U8269 (N_8269,N_7574,N_7946);
or U8270 (N_8270,N_7811,N_7783);
nor U8271 (N_8271,N_7936,N_7971);
nand U8272 (N_8272,N_7831,N_7803);
nand U8273 (N_8273,N_7962,N_7676);
nor U8274 (N_8274,N_7898,N_7685);
and U8275 (N_8275,N_7906,N_7528);
or U8276 (N_8276,N_7887,N_7563);
nand U8277 (N_8277,N_7840,N_7539);
xor U8278 (N_8278,N_7552,N_7568);
and U8279 (N_8279,N_7978,N_7907);
nor U8280 (N_8280,N_7852,N_7837);
nand U8281 (N_8281,N_7526,N_7520);
nor U8282 (N_8282,N_7724,N_7916);
nand U8283 (N_8283,N_7626,N_7977);
nor U8284 (N_8284,N_7967,N_7667);
and U8285 (N_8285,N_7754,N_7635);
or U8286 (N_8286,N_7656,N_7919);
or U8287 (N_8287,N_7514,N_7527);
or U8288 (N_8288,N_7871,N_7641);
nor U8289 (N_8289,N_7853,N_7998);
nor U8290 (N_8290,N_7914,N_7575);
xor U8291 (N_8291,N_7705,N_7856);
xor U8292 (N_8292,N_7831,N_7769);
xnor U8293 (N_8293,N_7571,N_7626);
and U8294 (N_8294,N_7689,N_7819);
nor U8295 (N_8295,N_7827,N_7709);
nand U8296 (N_8296,N_7963,N_7853);
nor U8297 (N_8297,N_7939,N_7813);
nand U8298 (N_8298,N_7648,N_7733);
nor U8299 (N_8299,N_7580,N_7665);
nor U8300 (N_8300,N_7671,N_7706);
and U8301 (N_8301,N_7558,N_7935);
or U8302 (N_8302,N_7561,N_7600);
nand U8303 (N_8303,N_7700,N_7767);
or U8304 (N_8304,N_7632,N_7770);
nand U8305 (N_8305,N_7731,N_7777);
and U8306 (N_8306,N_7675,N_7697);
or U8307 (N_8307,N_7848,N_7934);
nand U8308 (N_8308,N_7792,N_7639);
or U8309 (N_8309,N_7894,N_7877);
nor U8310 (N_8310,N_7947,N_7873);
or U8311 (N_8311,N_7962,N_7736);
nand U8312 (N_8312,N_7826,N_7699);
and U8313 (N_8313,N_7633,N_7872);
xnor U8314 (N_8314,N_7891,N_7834);
nor U8315 (N_8315,N_7713,N_7621);
nand U8316 (N_8316,N_7987,N_7968);
and U8317 (N_8317,N_7506,N_7790);
nor U8318 (N_8318,N_7552,N_7538);
or U8319 (N_8319,N_7816,N_7994);
nand U8320 (N_8320,N_7819,N_7853);
xnor U8321 (N_8321,N_7739,N_7606);
and U8322 (N_8322,N_7758,N_7747);
nor U8323 (N_8323,N_7598,N_7701);
xor U8324 (N_8324,N_7631,N_7929);
xnor U8325 (N_8325,N_7812,N_7658);
nand U8326 (N_8326,N_7794,N_7692);
nand U8327 (N_8327,N_7655,N_7946);
nor U8328 (N_8328,N_7761,N_7770);
nand U8329 (N_8329,N_7524,N_7805);
xor U8330 (N_8330,N_7673,N_7695);
or U8331 (N_8331,N_7757,N_7881);
or U8332 (N_8332,N_7821,N_7755);
nor U8333 (N_8333,N_7885,N_7991);
nand U8334 (N_8334,N_7958,N_7984);
nor U8335 (N_8335,N_7702,N_7958);
nor U8336 (N_8336,N_7764,N_7926);
or U8337 (N_8337,N_7745,N_7730);
nand U8338 (N_8338,N_7554,N_7607);
nand U8339 (N_8339,N_7948,N_7656);
nand U8340 (N_8340,N_7651,N_7637);
nand U8341 (N_8341,N_7654,N_7502);
and U8342 (N_8342,N_7690,N_7536);
or U8343 (N_8343,N_7564,N_7505);
or U8344 (N_8344,N_7568,N_7571);
xor U8345 (N_8345,N_7782,N_7509);
nor U8346 (N_8346,N_7519,N_7818);
nor U8347 (N_8347,N_7558,N_7980);
and U8348 (N_8348,N_7956,N_7942);
and U8349 (N_8349,N_7609,N_7562);
or U8350 (N_8350,N_7628,N_7723);
and U8351 (N_8351,N_7569,N_7922);
xor U8352 (N_8352,N_7682,N_7715);
or U8353 (N_8353,N_7681,N_7730);
or U8354 (N_8354,N_7809,N_7907);
nand U8355 (N_8355,N_7545,N_7932);
nand U8356 (N_8356,N_7615,N_7938);
or U8357 (N_8357,N_7551,N_7650);
or U8358 (N_8358,N_7638,N_7656);
xor U8359 (N_8359,N_7902,N_7914);
xnor U8360 (N_8360,N_7853,N_7878);
or U8361 (N_8361,N_7502,N_7717);
nor U8362 (N_8362,N_7902,N_7776);
or U8363 (N_8363,N_7969,N_7721);
nor U8364 (N_8364,N_7511,N_7994);
nor U8365 (N_8365,N_7657,N_7938);
xnor U8366 (N_8366,N_7551,N_7922);
and U8367 (N_8367,N_7932,N_7806);
nand U8368 (N_8368,N_7737,N_7668);
nor U8369 (N_8369,N_7584,N_7587);
and U8370 (N_8370,N_7585,N_7843);
nand U8371 (N_8371,N_7912,N_7816);
or U8372 (N_8372,N_7900,N_7617);
nor U8373 (N_8373,N_7846,N_7527);
nand U8374 (N_8374,N_7909,N_7713);
or U8375 (N_8375,N_7645,N_7561);
or U8376 (N_8376,N_7501,N_7793);
nor U8377 (N_8377,N_7531,N_7956);
and U8378 (N_8378,N_7906,N_7794);
and U8379 (N_8379,N_7977,N_7559);
nand U8380 (N_8380,N_7966,N_7898);
nand U8381 (N_8381,N_7782,N_7866);
nor U8382 (N_8382,N_7991,N_7934);
xor U8383 (N_8383,N_7514,N_7564);
and U8384 (N_8384,N_7692,N_7527);
and U8385 (N_8385,N_7614,N_7712);
nor U8386 (N_8386,N_7962,N_7963);
nor U8387 (N_8387,N_7959,N_7642);
and U8388 (N_8388,N_7988,N_7576);
or U8389 (N_8389,N_7804,N_7760);
nor U8390 (N_8390,N_7536,N_7816);
or U8391 (N_8391,N_7914,N_7602);
or U8392 (N_8392,N_7982,N_7677);
or U8393 (N_8393,N_7581,N_7846);
nor U8394 (N_8394,N_7796,N_7861);
nor U8395 (N_8395,N_7604,N_7543);
or U8396 (N_8396,N_7904,N_7676);
or U8397 (N_8397,N_7566,N_7515);
nor U8398 (N_8398,N_7553,N_7975);
or U8399 (N_8399,N_7817,N_7596);
xnor U8400 (N_8400,N_7783,N_7902);
and U8401 (N_8401,N_7858,N_7541);
nand U8402 (N_8402,N_7925,N_7701);
nand U8403 (N_8403,N_7768,N_7991);
and U8404 (N_8404,N_7559,N_7900);
nor U8405 (N_8405,N_7902,N_7602);
xnor U8406 (N_8406,N_7614,N_7872);
or U8407 (N_8407,N_7635,N_7675);
nand U8408 (N_8408,N_7536,N_7576);
and U8409 (N_8409,N_7732,N_7886);
xor U8410 (N_8410,N_7978,N_7561);
or U8411 (N_8411,N_7520,N_7779);
nand U8412 (N_8412,N_7723,N_7548);
nand U8413 (N_8413,N_7559,N_7889);
and U8414 (N_8414,N_7767,N_7589);
or U8415 (N_8415,N_7842,N_7941);
nand U8416 (N_8416,N_7776,N_7612);
nand U8417 (N_8417,N_7634,N_7638);
nand U8418 (N_8418,N_7561,N_7802);
nand U8419 (N_8419,N_7817,N_7946);
and U8420 (N_8420,N_7651,N_7648);
nand U8421 (N_8421,N_7946,N_7780);
and U8422 (N_8422,N_7883,N_7981);
xor U8423 (N_8423,N_7907,N_7581);
nor U8424 (N_8424,N_7956,N_7752);
nor U8425 (N_8425,N_7842,N_7603);
or U8426 (N_8426,N_7637,N_7919);
nor U8427 (N_8427,N_7594,N_7625);
nor U8428 (N_8428,N_7842,N_7921);
nand U8429 (N_8429,N_7609,N_7860);
or U8430 (N_8430,N_7719,N_7723);
or U8431 (N_8431,N_7514,N_7946);
or U8432 (N_8432,N_7608,N_7668);
and U8433 (N_8433,N_7997,N_7560);
nor U8434 (N_8434,N_7528,N_7558);
and U8435 (N_8435,N_7882,N_7663);
or U8436 (N_8436,N_7719,N_7661);
and U8437 (N_8437,N_7562,N_7980);
or U8438 (N_8438,N_7729,N_7599);
nand U8439 (N_8439,N_7527,N_7903);
nand U8440 (N_8440,N_7892,N_7739);
and U8441 (N_8441,N_7769,N_7504);
or U8442 (N_8442,N_7984,N_7690);
or U8443 (N_8443,N_7721,N_7768);
and U8444 (N_8444,N_7671,N_7592);
nor U8445 (N_8445,N_7947,N_7715);
nand U8446 (N_8446,N_7902,N_7860);
xor U8447 (N_8447,N_7692,N_7976);
and U8448 (N_8448,N_7841,N_7784);
or U8449 (N_8449,N_7627,N_7681);
xor U8450 (N_8450,N_7577,N_7987);
and U8451 (N_8451,N_7553,N_7774);
nand U8452 (N_8452,N_7650,N_7562);
nand U8453 (N_8453,N_7939,N_7661);
and U8454 (N_8454,N_7991,N_7716);
nand U8455 (N_8455,N_7682,N_7554);
nor U8456 (N_8456,N_7756,N_7579);
nor U8457 (N_8457,N_7952,N_7605);
nor U8458 (N_8458,N_7604,N_7964);
and U8459 (N_8459,N_7746,N_7925);
nor U8460 (N_8460,N_7937,N_7737);
nand U8461 (N_8461,N_7610,N_7546);
xor U8462 (N_8462,N_7837,N_7954);
or U8463 (N_8463,N_7702,N_7563);
nor U8464 (N_8464,N_7887,N_7707);
nand U8465 (N_8465,N_7738,N_7874);
nor U8466 (N_8466,N_7753,N_7537);
nand U8467 (N_8467,N_7921,N_7779);
and U8468 (N_8468,N_7731,N_7608);
xor U8469 (N_8469,N_7740,N_7847);
nand U8470 (N_8470,N_7790,N_7820);
xnor U8471 (N_8471,N_7635,N_7541);
and U8472 (N_8472,N_7813,N_7635);
nor U8473 (N_8473,N_7953,N_7500);
nand U8474 (N_8474,N_7902,N_7805);
or U8475 (N_8475,N_7621,N_7648);
nor U8476 (N_8476,N_7513,N_7946);
nand U8477 (N_8477,N_7757,N_7573);
and U8478 (N_8478,N_7792,N_7917);
nor U8479 (N_8479,N_7636,N_7566);
nand U8480 (N_8480,N_7773,N_7967);
and U8481 (N_8481,N_7995,N_7709);
and U8482 (N_8482,N_7506,N_7714);
or U8483 (N_8483,N_7624,N_7652);
and U8484 (N_8484,N_7754,N_7584);
nand U8485 (N_8485,N_7768,N_7814);
nand U8486 (N_8486,N_7701,N_7841);
nand U8487 (N_8487,N_7917,N_7741);
and U8488 (N_8488,N_7890,N_7703);
or U8489 (N_8489,N_7746,N_7820);
nor U8490 (N_8490,N_7770,N_7654);
xnor U8491 (N_8491,N_7996,N_7530);
or U8492 (N_8492,N_7648,N_7576);
xnor U8493 (N_8493,N_7881,N_7621);
and U8494 (N_8494,N_7798,N_7762);
or U8495 (N_8495,N_7782,N_7908);
nor U8496 (N_8496,N_7527,N_7863);
nand U8497 (N_8497,N_7982,N_7536);
and U8498 (N_8498,N_7858,N_7561);
and U8499 (N_8499,N_7543,N_7945);
nor U8500 (N_8500,N_8395,N_8102);
nand U8501 (N_8501,N_8356,N_8214);
nand U8502 (N_8502,N_8335,N_8343);
or U8503 (N_8503,N_8405,N_8412);
xnor U8504 (N_8504,N_8314,N_8017);
nor U8505 (N_8505,N_8059,N_8205);
or U8506 (N_8506,N_8424,N_8272);
nor U8507 (N_8507,N_8093,N_8260);
or U8508 (N_8508,N_8271,N_8270);
or U8509 (N_8509,N_8290,N_8193);
or U8510 (N_8510,N_8005,N_8147);
nor U8511 (N_8511,N_8004,N_8348);
and U8512 (N_8512,N_8153,N_8376);
and U8513 (N_8513,N_8083,N_8436);
nor U8514 (N_8514,N_8024,N_8247);
nand U8515 (N_8515,N_8457,N_8131);
nor U8516 (N_8516,N_8142,N_8306);
and U8517 (N_8517,N_8013,N_8374);
and U8518 (N_8518,N_8252,N_8105);
xnor U8519 (N_8519,N_8304,N_8345);
nor U8520 (N_8520,N_8162,N_8240);
nand U8521 (N_8521,N_8273,N_8163);
nor U8522 (N_8522,N_8367,N_8365);
or U8523 (N_8523,N_8313,N_8113);
nand U8524 (N_8524,N_8279,N_8074);
or U8525 (N_8525,N_8229,N_8026);
or U8526 (N_8526,N_8319,N_8032);
nand U8527 (N_8527,N_8009,N_8016);
and U8528 (N_8528,N_8164,N_8480);
nand U8529 (N_8529,N_8284,N_8328);
xnor U8530 (N_8530,N_8235,N_8409);
nand U8531 (N_8531,N_8010,N_8045);
and U8532 (N_8532,N_8497,N_8106);
xnor U8533 (N_8533,N_8188,N_8262);
and U8534 (N_8534,N_8408,N_8044);
nor U8535 (N_8535,N_8359,N_8478);
and U8536 (N_8536,N_8255,N_8261);
nand U8537 (N_8537,N_8419,N_8060);
nor U8538 (N_8538,N_8293,N_8054);
or U8539 (N_8539,N_8040,N_8406);
or U8540 (N_8540,N_8486,N_8307);
nand U8541 (N_8541,N_8310,N_8180);
and U8542 (N_8542,N_8015,N_8128);
nor U8543 (N_8543,N_8249,N_8047);
or U8544 (N_8544,N_8133,N_8366);
or U8545 (N_8545,N_8447,N_8484);
or U8546 (N_8546,N_8353,N_8487);
and U8547 (N_8547,N_8144,N_8337);
xor U8548 (N_8548,N_8455,N_8065);
and U8549 (N_8549,N_8096,N_8030);
or U8550 (N_8550,N_8159,N_8108);
nand U8551 (N_8551,N_8129,N_8226);
nor U8552 (N_8552,N_8172,N_8033);
xnor U8553 (N_8553,N_8372,N_8453);
and U8554 (N_8554,N_8426,N_8336);
and U8555 (N_8555,N_8377,N_8416);
nor U8556 (N_8556,N_8222,N_8362);
nor U8557 (N_8557,N_8422,N_8473);
nand U8558 (N_8558,N_8119,N_8115);
xnor U8559 (N_8559,N_8018,N_8434);
nand U8560 (N_8560,N_8090,N_8078);
xor U8561 (N_8561,N_8150,N_8461);
or U8562 (N_8562,N_8000,N_8458);
or U8563 (N_8563,N_8369,N_8389);
or U8564 (N_8564,N_8154,N_8138);
nor U8565 (N_8565,N_8498,N_8274);
and U8566 (N_8566,N_8267,N_8251);
and U8567 (N_8567,N_8479,N_8081);
nor U8568 (N_8568,N_8495,N_8287);
nor U8569 (N_8569,N_8371,N_8223);
or U8570 (N_8570,N_8349,N_8330);
nor U8571 (N_8571,N_8442,N_8325);
xor U8572 (N_8572,N_8415,N_8309);
or U8573 (N_8573,N_8396,N_8168);
nor U8574 (N_8574,N_8143,N_8097);
and U8575 (N_8575,N_8176,N_8241);
and U8576 (N_8576,N_8303,N_8340);
or U8577 (N_8577,N_8126,N_8470);
and U8578 (N_8578,N_8165,N_8069);
and U8579 (N_8579,N_8494,N_8450);
nand U8580 (N_8580,N_8316,N_8490);
nor U8581 (N_8581,N_8234,N_8114);
nand U8582 (N_8582,N_8347,N_8204);
and U8583 (N_8583,N_8427,N_8360);
or U8584 (N_8584,N_8301,N_8382);
nor U8585 (N_8585,N_8058,N_8116);
and U8586 (N_8586,N_8346,N_8051);
and U8587 (N_8587,N_8179,N_8275);
or U8588 (N_8588,N_8481,N_8437);
nor U8589 (N_8589,N_8338,N_8381);
or U8590 (N_8590,N_8370,N_8021);
xnor U8591 (N_8591,N_8292,N_8149);
nor U8592 (N_8592,N_8191,N_8035);
nor U8593 (N_8593,N_8469,N_8203);
nor U8594 (N_8594,N_8425,N_8094);
nand U8595 (N_8595,N_8111,N_8312);
or U8596 (N_8596,N_8390,N_8295);
and U8597 (N_8597,N_8167,N_8438);
xnor U8598 (N_8598,N_8326,N_8482);
or U8599 (N_8599,N_8254,N_8243);
nor U8600 (N_8600,N_8038,N_8091);
or U8601 (N_8601,N_8134,N_8029);
nand U8602 (N_8602,N_8070,N_8061);
and U8603 (N_8603,N_8189,N_8103);
or U8604 (N_8604,N_8207,N_8429);
xnor U8605 (N_8605,N_8196,N_8423);
and U8606 (N_8606,N_8146,N_8161);
or U8607 (N_8607,N_8407,N_8449);
nand U8608 (N_8608,N_8397,N_8151);
nor U8609 (N_8609,N_8075,N_8351);
nor U8610 (N_8610,N_8417,N_8403);
xor U8611 (N_8611,N_8012,N_8386);
nor U8612 (N_8612,N_8049,N_8098);
nand U8613 (N_8613,N_8368,N_8354);
nand U8614 (N_8614,N_8357,N_8084);
and U8615 (N_8615,N_8391,N_8462);
xnor U8616 (N_8616,N_8464,N_8192);
nand U8617 (N_8617,N_8334,N_8037);
nand U8618 (N_8618,N_8311,N_8472);
nand U8619 (N_8619,N_8410,N_8228);
xnor U8620 (N_8620,N_8291,N_8135);
and U8621 (N_8621,N_8099,N_8122);
and U8622 (N_8622,N_8210,N_8298);
xor U8623 (N_8623,N_8031,N_8242);
nor U8624 (N_8624,N_8110,N_8332);
and U8625 (N_8625,N_8392,N_8281);
nand U8626 (N_8626,N_8398,N_8130);
or U8627 (N_8627,N_8302,N_8411);
or U8628 (N_8628,N_8285,N_8460);
or U8629 (N_8629,N_8157,N_8198);
nand U8630 (N_8630,N_8175,N_8086);
nor U8631 (N_8631,N_8046,N_8118);
xor U8632 (N_8632,N_8089,N_8294);
nand U8633 (N_8633,N_8227,N_8466);
and U8634 (N_8634,N_8350,N_8171);
nand U8635 (N_8635,N_8231,N_8233);
or U8636 (N_8636,N_8394,N_8296);
or U8637 (N_8637,N_8197,N_8208);
or U8638 (N_8638,N_8217,N_8269);
and U8639 (N_8639,N_8001,N_8211);
nand U8640 (N_8640,N_8475,N_8341);
or U8641 (N_8641,N_8344,N_8324);
and U8642 (N_8642,N_8139,N_8331);
or U8643 (N_8643,N_8428,N_8363);
nor U8644 (N_8644,N_8430,N_8006);
nand U8645 (N_8645,N_8063,N_8441);
or U8646 (N_8646,N_8236,N_8297);
nand U8647 (N_8647,N_8280,N_8185);
and U8648 (N_8648,N_8431,N_8039);
or U8649 (N_8649,N_8025,N_8471);
and U8650 (N_8650,N_8265,N_8318);
nand U8651 (N_8651,N_8246,N_8257);
nand U8652 (N_8652,N_8219,N_8064);
and U8653 (N_8653,N_8433,N_8073);
nor U8654 (N_8654,N_8125,N_8259);
nand U8655 (N_8655,N_8399,N_8209);
or U8656 (N_8656,N_8380,N_8062);
nand U8657 (N_8657,N_8158,N_8352);
or U8658 (N_8658,N_8050,N_8104);
nand U8659 (N_8659,N_8170,N_8095);
nor U8660 (N_8660,N_8169,N_8420);
nor U8661 (N_8661,N_8156,N_8393);
nand U8662 (N_8662,N_8387,N_8072);
or U8663 (N_8663,N_8414,N_8003);
or U8664 (N_8664,N_8355,N_8463);
nor U8665 (N_8665,N_8439,N_8404);
xnor U8666 (N_8666,N_8446,N_8201);
nand U8667 (N_8667,N_8375,N_8076);
and U8668 (N_8668,N_8451,N_8087);
nand U8669 (N_8669,N_8238,N_8182);
nor U8670 (N_8670,N_8489,N_8286);
and U8671 (N_8671,N_8278,N_8027);
nand U8672 (N_8672,N_8100,N_8212);
xnor U8673 (N_8673,N_8183,N_8402);
and U8674 (N_8674,N_8456,N_8499);
nor U8675 (N_8675,N_8008,N_8358);
or U8676 (N_8676,N_8215,N_8256);
xnor U8677 (N_8677,N_8239,N_8007);
and U8678 (N_8678,N_8329,N_8401);
nor U8679 (N_8679,N_8277,N_8468);
nand U8680 (N_8680,N_8080,N_8283);
and U8681 (N_8681,N_8042,N_8444);
or U8682 (N_8682,N_8057,N_8079);
nand U8683 (N_8683,N_8485,N_8378);
nand U8684 (N_8684,N_8225,N_8383);
nand U8685 (N_8685,N_8220,N_8440);
xor U8686 (N_8686,N_8022,N_8052);
or U8687 (N_8687,N_8342,N_8048);
or U8688 (N_8688,N_8177,N_8121);
or U8689 (N_8689,N_8317,N_8492);
xnor U8690 (N_8690,N_8199,N_8476);
or U8691 (N_8691,N_8232,N_8379);
nand U8692 (N_8692,N_8361,N_8483);
nor U8693 (N_8693,N_8152,N_8184);
xor U8694 (N_8694,N_8132,N_8448);
and U8695 (N_8695,N_8245,N_8300);
xor U8696 (N_8696,N_8244,N_8493);
xor U8697 (N_8697,N_8195,N_8263);
nand U8698 (N_8698,N_8221,N_8202);
and U8699 (N_8699,N_8124,N_8034);
and U8700 (N_8700,N_8085,N_8088);
nor U8701 (N_8701,N_8068,N_8459);
nor U8702 (N_8702,N_8266,N_8173);
nand U8703 (N_8703,N_8299,N_8488);
or U8704 (N_8704,N_8077,N_8036);
or U8705 (N_8705,N_8019,N_8140);
and U8706 (N_8706,N_8200,N_8258);
or U8707 (N_8707,N_8230,N_8327);
and U8708 (N_8708,N_8043,N_8160);
nand U8709 (N_8709,N_8491,N_8385);
nand U8710 (N_8710,N_8289,N_8432);
or U8711 (N_8711,N_8454,N_8155);
or U8712 (N_8712,N_8218,N_8067);
nand U8713 (N_8713,N_8400,N_8092);
and U8714 (N_8714,N_8023,N_8137);
xor U8715 (N_8715,N_8276,N_8206);
xnor U8716 (N_8716,N_8216,N_8107);
xnor U8717 (N_8717,N_8053,N_8011);
or U8718 (N_8718,N_8477,N_8112);
or U8719 (N_8719,N_8213,N_8020);
nand U8720 (N_8720,N_8194,N_8333);
nor U8721 (N_8721,N_8384,N_8288);
nand U8722 (N_8722,N_8120,N_8339);
nand U8723 (N_8723,N_8181,N_8496);
nand U8724 (N_8724,N_8178,N_8320);
or U8725 (N_8725,N_8250,N_8145);
xor U8726 (N_8726,N_8109,N_8148);
or U8727 (N_8727,N_8123,N_8305);
and U8728 (N_8728,N_8101,N_8364);
and U8729 (N_8729,N_8071,N_8055);
and U8730 (N_8730,N_8467,N_8117);
and U8731 (N_8731,N_8465,N_8190);
nand U8732 (N_8732,N_8388,N_8474);
nor U8733 (N_8733,N_8248,N_8174);
and U8734 (N_8734,N_8056,N_8224);
or U8735 (N_8735,N_8435,N_8321);
or U8736 (N_8736,N_8014,N_8308);
or U8737 (N_8737,N_8253,N_8315);
xor U8738 (N_8738,N_8136,N_8186);
or U8739 (N_8739,N_8268,N_8141);
nor U8740 (N_8740,N_8166,N_8282);
or U8741 (N_8741,N_8127,N_8041);
and U8742 (N_8742,N_8452,N_8421);
nor U8743 (N_8743,N_8264,N_8323);
or U8744 (N_8744,N_8187,N_8002);
nand U8745 (N_8745,N_8413,N_8418);
or U8746 (N_8746,N_8028,N_8237);
nor U8747 (N_8747,N_8373,N_8082);
and U8748 (N_8748,N_8445,N_8322);
nand U8749 (N_8749,N_8066,N_8443);
nor U8750 (N_8750,N_8047,N_8005);
xnor U8751 (N_8751,N_8167,N_8344);
and U8752 (N_8752,N_8336,N_8246);
nand U8753 (N_8753,N_8210,N_8485);
nand U8754 (N_8754,N_8340,N_8173);
or U8755 (N_8755,N_8239,N_8445);
or U8756 (N_8756,N_8326,N_8230);
or U8757 (N_8757,N_8087,N_8164);
and U8758 (N_8758,N_8446,N_8372);
or U8759 (N_8759,N_8346,N_8259);
or U8760 (N_8760,N_8259,N_8273);
nor U8761 (N_8761,N_8036,N_8200);
nand U8762 (N_8762,N_8452,N_8174);
nand U8763 (N_8763,N_8024,N_8116);
and U8764 (N_8764,N_8450,N_8340);
nand U8765 (N_8765,N_8239,N_8132);
and U8766 (N_8766,N_8337,N_8038);
nor U8767 (N_8767,N_8417,N_8315);
or U8768 (N_8768,N_8030,N_8404);
or U8769 (N_8769,N_8483,N_8091);
or U8770 (N_8770,N_8052,N_8259);
nand U8771 (N_8771,N_8340,N_8133);
and U8772 (N_8772,N_8025,N_8493);
nor U8773 (N_8773,N_8434,N_8403);
or U8774 (N_8774,N_8317,N_8394);
nor U8775 (N_8775,N_8441,N_8108);
nand U8776 (N_8776,N_8376,N_8481);
or U8777 (N_8777,N_8453,N_8132);
nor U8778 (N_8778,N_8100,N_8167);
or U8779 (N_8779,N_8476,N_8036);
nand U8780 (N_8780,N_8031,N_8459);
nor U8781 (N_8781,N_8439,N_8302);
xor U8782 (N_8782,N_8128,N_8240);
or U8783 (N_8783,N_8034,N_8411);
nand U8784 (N_8784,N_8060,N_8481);
or U8785 (N_8785,N_8234,N_8418);
nor U8786 (N_8786,N_8425,N_8116);
nor U8787 (N_8787,N_8365,N_8304);
nand U8788 (N_8788,N_8418,N_8041);
or U8789 (N_8789,N_8172,N_8276);
nor U8790 (N_8790,N_8341,N_8418);
nor U8791 (N_8791,N_8287,N_8002);
and U8792 (N_8792,N_8272,N_8173);
or U8793 (N_8793,N_8205,N_8132);
nand U8794 (N_8794,N_8029,N_8326);
nand U8795 (N_8795,N_8105,N_8385);
nand U8796 (N_8796,N_8414,N_8201);
nand U8797 (N_8797,N_8354,N_8313);
nand U8798 (N_8798,N_8114,N_8274);
and U8799 (N_8799,N_8162,N_8410);
or U8800 (N_8800,N_8476,N_8401);
nor U8801 (N_8801,N_8467,N_8105);
nand U8802 (N_8802,N_8176,N_8395);
or U8803 (N_8803,N_8468,N_8460);
or U8804 (N_8804,N_8491,N_8338);
and U8805 (N_8805,N_8395,N_8149);
nor U8806 (N_8806,N_8382,N_8337);
nand U8807 (N_8807,N_8400,N_8282);
or U8808 (N_8808,N_8439,N_8012);
xnor U8809 (N_8809,N_8110,N_8151);
nor U8810 (N_8810,N_8159,N_8445);
and U8811 (N_8811,N_8483,N_8257);
nor U8812 (N_8812,N_8068,N_8062);
nand U8813 (N_8813,N_8381,N_8273);
or U8814 (N_8814,N_8418,N_8269);
nand U8815 (N_8815,N_8280,N_8192);
nand U8816 (N_8816,N_8422,N_8234);
nor U8817 (N_8817,N_8247,N_8460);
and U8818 (N_8818,N_8138,N_8272);
or U8819 (N_8819,N_8066,N_8042);
or U8820 (N_8820,N_8344,N_8012);
nand U8821 (N_8821,N_8462,N_8345);
xor U8822 (N_8822,N_8137,N_8477);
nor U8823 (N_8823,N_8311,N_8130);
nor U8824 (N_8824,N_8013,N_8468);
nor U8825 (N_8825,N_8341,N_8376);
and U8826 (N_8826,N_8247,N_8244);
nor U8827 (N_8827,N_8365,N_8017);
nand U8828 (N_8828,N_8123,N_8008);
and U8829 (N_8829,N_8465,N_8455);
and U8830 (N_8830,N_8099,N_8359);
xnor U8831 (N_8831,N_8136,N_8353);
nor U8832 (N_8832,N_8035,N_8479);
xnor U8833 (N_8833,N_8295,N_8168);
nand U8834 (N_8834,N_8033,N_8297);
nand U8835 (N_8835,N_8090,N_8001);
nor U8836 (N_8836,N_8405,N_8088);
or U8837 (N_8837,N_8142,N_8193);
nand U8838 (N_8838,N_8259,N_8196);
nor U8839 (N_8839,N_8028,N_8265);
or U8840 (N_8840,N_8211,N_8185);
nand U8841 (N_8841,N_8168,N_8178);
and U8842 (N_8842,N_8454,N_8013);
or U8843 (N_8843,N_8245,N_8234);
or U8844 (N_8844,N_8212,N_8029);
or U8845 (N_8845,N_8410,N_8059);
or U8846 (N_8846,N_8482,N_8306);
and U8847 (N_8847,N_8333,N_8308);
nand U8848 (N_8848,N_8432,N_8354);
nand U8849 (N_8849,N_8360,N_8340);
nand U8850 (N_8850,N_8055,N_8293);
nand U8851 (N_8851,N_8276,N_8344);
xnor U8852 (N_8852,N_8325,N_8136);
nand U8853 (N_8853,N_8363,N_8443);
or U8854 (N_8854,N_8008,N_8055);
nand U8855 (N_8855,N_8041,N_8113);
or U8856 (N_8856,N_8047,N_8304);
and U8857 (N_8857,N_8204,N_8142);
and U8858 (N_8858,N_8493,N_8077);
xor U8859 (N_8859,N_8006,N_8495);
and U8860 (N_8860,N_8305,N_8257);
nand U8861 (N_8861,N_8497,N_8002);
or U8862 (N_8862,N_8485,N_8288);
xor U8863 (N_8863,N_8147,N_8229);
nand U8864 (N_8864,N_8460,N_8191);
xnor U8865 (N_8865,N_8358,N_8432);
nor U8866 (N_8866,N_8437,N_8424);
nand U8867 (N_8867,N_8403,N_8397);
xor U8868 (N_8868,N_8006,N_8289);
nor U8869 (N_8869,N_8305,N_8186);
nand U8870 (N_8870,N_8075,N_8340);
or U8871 (N_8871,N_8237,N_8093);
nor U8872 (N_8872,N_8425,N_8424);
nor U8873 (N_8873,N_8125,N_8296);
and U8874 (N_8874,N_8469,N_8003);
nor U8875 (N_8875,N_8428,N_8406);
nand U8876 (N_8876,N_8145,N_8038);
nand U8877 (N_8877,N_8447,N_8251);
or U8878 (N_8878,N_8268,N_8160);
and U8879 (N_8879,N_8170,N_8441);
xnor U8880 (N_8880,N_8437,N_8359);
and U8881 (N_8881,N_8495,N_8256);
nand U8882 (N_8882,N_8447,N_8487);
and U8883 (N_8883,N_8329,N_8082);
nand U8884 (N_8884,N_8286,N_8354);
xnor U8885 (N_8885,N_8498,N_8338);
nor U8886 (N_8886,N_8416,N_8094);
nor U8887 (N_8887,N_8313,N_8106);
or U8888 (N_8888,N_8331,N_8301);
and U8889 (N_8889,N_8377,N_8311);
xor U8890 (N_8890,N_8184,N_8082);
nand U8891 (N_8891,N_8302,N_8391);
and U8892 (N_8892,N_8303,N_8087);
xor U8893 (N_8893,N_8172,N_8210);
nand U8894 (N_8894,N_8442,N_8090);
nand U8895 (N_8895,N_8100,N_8367);
nor U8896 (N_8896,N_8402,N_8110);
xor U8897 (N_8897,N_8020,N_8032);
and U8898 (N_8898,N_8229,N_8275);
nor U8899 (N_8899,N_8212,N_8276);
nor U8900 (N_8900,N_8434,N_8142);
nor U8901 (N_8901,N_8432,N_8304);
nand U8902 (N_8902,N_8071,N_8433);
nor U8903 (N_8903,N_8003,N_8396);
nor U8904 (N_8904,N_8167,N_8369);
nor U8905 (N_8905,N_8161,N_8263);
and U8906 (N_8906,N_8246,N_8134);
and U8907 (N_8907,N_8499,N_8205);
or U8908 (N_8908,N_8183,N_8315);
nor U8909 (N_8909,N_8171,N_8030);
nor U8910 (N_8910,N_8462,N_8078);
or U8911 (N_8911,N_8378,N_8291);
nand U8912 (N_8912,N_8461,N_8015);
nor U8913 (N_8913,N_8325,N_8247);
nand U8914 (N_8914,N_8099,N_8189);
nand U8915 (N_8915,N_8390,N_8062);
xor U8916 (N_8916,N_8293,N_8239);
or U8917 (N_8917,N_8244,N_8009);
and U8918 (N_8918,N_8375,N_8263);
nor U8919 (N_8919,N_8079,N_8301);
and U8920 (N_8920,N_8476,N_8198);
nor U8921 (N_8921,N_8253,N_8073);
nand U8922 (N_8922,N_8270,N_8379);
or U8923 (N_8923,N_8104,N_8278);
or U8924 (N_8924,N_8090,N_8209);
or U8925 (N_8925,N_8208,N_8384);
nor U8926 (N_8926,N_8214,N_8476);
nor U8927 (N_8927,N_8247,N_8485);
nand U8928 (N_8928,N_8474,N_8402);
nand U8929 (N_8929,N_8452,N_8347);
and U8930 (N_8930,N_8349,N_8058);
or U8931 (N_8931,N_8215,N_8414);
nand U8932 (N_8932,N_8030,N_8442);
xnor U8933 (N_8933,N_8173,N_8303);
nor U8934 (N_8934,N_8278,N_8346);
or U8935 (N_8935,N_8222,N_8143);
and U8936 (N_8936,N_8478,N_8311);
nor U8937 (N_8937,N_8353,N_8201);
or U8938 (N_8938,N_8088,N_8336);
xor U8939 (N_8939,N_8366,N_8109);
and U8940 (N_8940,N_8467,N_8154);
xnor U8941 (N_8941,N_8139,N_8269);
and U8942 (N_8942,N_8206,N_8117);
nand U8943 (N_8943,N_8436,N_8386);
or U8944 (N_8944,N_8024,N_8148);
nor U8945 (N_8945,N_8156,N_8248);
or U8946 (N_8946,N_8413,N_8324);
nor U8947 (N_8947,N_8287,N_8272);
nand U8948 (N_8948,N_8179,N_8418);
nand U8949 (N_8949,N_8393,N_8133);
and U8950 (N_8950,N_8269,N_8346);
nand U8951 (N_8951,N_8470,N_8274);
or U8952 (N_8952,N_8373,N_8037);
or U8953 (N_8953,N_8004,N_8151);
nor U8954 (N_8954,N_8288,N_8225);
nor U8955 (N_8955,N_8226,N_8463);
and U8956 (N_8956,N_8375,N_8485);
nand U8957 (N_8957,N_8086,N_8106);
or U8958 (N_8958,N_8340,N_8302);
or U8959 (N_8959,N_8272,N_8246);
nand U8960 (N_8960,N_8401,N_8048);
and U8961 (N_8961,N_8424,N_8372);
nor U8962 (N_8962,N_8471,N_8171);
or U8963 (N_8963,N_8375,N_8383);
or U8964 (N_8964,N_8374,N_8078);
and U8965 (N_8965,N_8300,N_8258);
or U8966 (N_8966,N_8282,N_8415);
or U8967 (N_8967,N_8477,N_8202);
and U8968 (N_8968,N_8023,N_8443);
xnor U8969 (N_8969,N_8021,N_8384);
nor U8970 (N_8970,N_8083,N_8053);
and U8971 (N_8971,N_8446,N_8219);
nor U8972 (N_8972,N_8336,N_8164);
and U8973 (N_8973,N_8023,N_8201);
nor U8974 (N_8974,N_8442,N_8121);
nor U8975 (N_8975,N_8023,N_8308);
or U8976 (N_8976,N_8113,N_8210);
nand U8977 (N_8977,N_8379,N_8114);
or U8978 (N_8978,N_8286,N_8016);
and U8979 (N_8979,N_8333,N_8132);
and U8980 (N_8980,N_8222,N_8181);
and U8981 (N_8981,N_8082,N_8490);
and U8982 (N_8982,N_8398,N_8364);
and U8983 (N_8983,N_8391,N_8479);
and U8984 (N_8984,N_8439,N_8045);
nor U8985 (N_8985,N_8184,N_8343);
nor U8986 (N_8986,N_8391,N_8130);
or U8987 (N_8987,N_8385,N_8401);
or U8988 (N_8988,N_8180,N_8103);
nand U8989 (N_8989,N_8067,N_8488);
xnor U8990 (N_8990,N_8380,N_8116);
nor U8991 (N_8991,N_8247,N_8369);
nand U8992 (N_8992,N_8294,N_8237);
or U8993 (N_8993,N_8142,N_8261);
or U8994 (N_8994,N_8308,N_8330);
and U8995 (N_8995,N_8348,N_8357);
nor U8996 (N_8996,N_8083,N_8338);
nand U8997 (N_8997,N_8106,N_8107);
nand U8998 (N_8998,N_8490,N_8215);
xor U8999 (N_8999,N_8236,N_8226);
or U9000 (N_9000,N_8957,N_8817);
nor U9001 (N_9001,N_8546,N_8852);
nand U9002 (N_9002,N_8800,N_8991);
or U9003 (N_9003,N_8646,N_8837);
nor U9004 (N_9004,N_8674,N_8879);
nand U9005 (N_9005,N_8983,N_8601);
nand U9006 (N_9006,N_8544,N_8966);
or U9007 (N_9007,N_8627,N_8736);
nor U9008 (N_9008,N_8662,N_8915);
nor U9009 (N_9009,N_8808,N_8774);
and U9010 (N_9010,N_8535,N_8805);
nor U9011 (N_9011,N_8625,N_8834);
and U9012 (N_9012,N_8593,N_8520);
xor U9013 (N_9013,N_8549,N_8637);
and U9014 (N_9014,N_8715,N_8610);
nand U9015 (N_9015,N_8998,N_8568);
nand U9016 (N_9016,N_8513,N_8695);
or U9017 (N_9017,N_8670,N_8575);
nand U9018 (N_9018,N_8502,N_8909);
nand U9019 (N_9019,N_8594,N_8894);
xor U9020 (N_9020,N_8986,N_8585);
nor U9021 (N_9021,N_8738,N_8865);
nor U9022 (N_9022,N_8723,N_8514);
or U9023 (N_9023,N_8776,N_8940);
nand U9024 (N_9024,N_8761,N_8950);
nor U9025 (N_9025,N_8503,N_8698);
nand U9026 (N_9026,N_8731,N_8821);
nand U9027 (N_9027,N_8807,N_8762);
nand U9028 (N_9028,N_8595,N_8725);
and U9029 (N_9029,N_8797,N_8939);
nor U9030 (N_9030,N_8883,N_8686);
or U9031 (N_9031,N_8641,N_8993);
xnor U9032 (N_9032,N_8908,N_8872);
nand U9033 (N_9033,N_8988,N_8848);
and U9034 (N_9034,N_8607,N_8948);
or U9035 (N_9035,N_8749,N_8841);
or U9036 (N_9036,N_8999,N_8878);
nor U9037 (N_9037,N_8525,N_8709);
xnor U9038 (N_9038,N_8666,N_8825);
nor U9039 (N_9039,N_8982,N_8540);
and U9040 (N_9040,N_8565,N_8985);
nand U9041 (N_9041,N_8693,N_8504);
or U9042 (N_9042,N_8953,N_8923);
nand U9043 (N_9043,N_8856,N_8614);
nand U9044 (N_9044,N_8927,N_8551);
and U9045 (N_9045,N_8510,N_8930);
nand U9046 (N_9046,N_8973,N_8645);
nand U9047 (N_9047,N_8789,N_8547);
nand U9048 (N_9048,N_8633,N_8810);
and U9049 (N_9049,N_8901,N_8959);
nand U9050 (N_9050,N_8592,N_8737);
nor U9051 (N_9051,N_8657,N_8941);
nand U9052 (N_9052,N_8877,N_8651);
nand U9053 (N_9053,N_8730,N_8820);
or U9054 (N_9054,N_8992,N_8963);
nor U9055 (N_9055,N_8919,N_8524);
and U9056 (N_9056,N_8669,N_8790);
and U9057 (N_9057,N_8951,N_8564);
or U9058 (N_9058,N_8580,N_8862);
nor U9059 (N_9059,N_8624,N_8728);
or U9060 (N_9060,N_8667,N_8965);
or U9061 (N_9061,N_8793,N_8716);
and U9062 (N_9062,N_8659,N_8557);
or U9063 (N_9063,N_8501,N_8591);
nand U9064 (N_9064,N_8896,N_8663);
nand U9065 (N_9065,N_8681,N_8753);
xor U9066 (N_9066,N_8765,N_8722);
nand U9067 (N_9067,N_8772,N_8828);
nor U9068 (N_9068,N_8553,N_8861);
nor U9069 (N_9069,N_8917,N_8881);
and U9070 (N_9070,N_8639,N_8745);
and U9071 (N_9071,N_8899,N_8928);
nor U9072 (N_9072,N_8717,N_8743);
or U9073 (N_9073,N_8644,N_8792);
and U9074 (N_9074,N_8739,N_8660);
xnor U9075 (N_9075,N_8542,N_8707);
and U9076 (N_9076,N_8888,N_8691);
xnor U9077 (N_9077,N_8532,N_8771);
nand U9078 (N_9078,N_8804,N_8802);
and U9079 (N_9079,N_8688,N_8947);
and U9080 (N_9080,N_8590,N_8523);
xnor U9081 (N_9081,N_8611,N_8935);
nor U9082 (N_9082,N_8665,N_8816);
nand U9083 (N_9083,N_8515,N_8826);
or U9084 (N_9084,N_8562,N_8705);
nor U9085 (N_9085,N_8823,N_8613);
nand U9086 (N_9086,N_8853,N_8572);
nor U9087 (N_9087,N_8934,N_8890);
nand U9088 (N_9088,N_8898,N_8618);
xnor U9089 (N_9089,N_8554,N_8638);
nand U9090 (N_9090,N_8766,N_8860);
and U9091 (N_9091,N_8757,N_8763);
nor U9092 (N_9092,N_8839,N_8573);
or U9093 (N_9093,N_8620,N_8996);
nand U9094 (N_9094,N_8897,N_8997);
nand U9095 (N_9095,N_8764,N_8740);
nor U9096 (N_9096,N_8664,N_8759);
and U9097 (N_9097,N_8543,N_8622);
nand U9098 (N_9098,N_8569,N_8720);
nand U9099 (N_9099,N_8902,N_8819);
nand U9100 (N_9100,N_8581,N_8527);
and U9101 (N_9101,N_8632,N_8972);
nand U9102 (N_9102,N_8714,N_8619);
xor U9103 (N_9103,N_8724,N_8995);
nor U9104 (N_9104,N_8752,N_8648);
xnor U9105 (N_9105,N_8608,N_8706);
nand U9106 (N_9106,N_8615,N_8956);
nor U9107 (N_9107,N_8529,N_8694);
nor U9108 (N_9108,N_8900,N_8975);
or U9109 (N_9109,N_8829,N_8799);
and U9110 (N_9110,N_8847,N_8617);
nor U9111 (N_9111,N_8584,N_8552);
and U9112 (N_9112,N_8711,N_8926);
nand U9113 (N_9113,N_8945,N_8741);
or U9114 (N_9114,N_8556,N_8954);
xor U9115 (N_9115,N_8747,N_8968);
and U9116 (N_9116,N_8893,N_8859);
nand U9117 (N_9117,N_8836,N_8567);
and U9118 (N_9118,N_8750,N_8978);
nand U9119 (N_9119,N_8606,N_8912);
xor U9120 (N_9120,N_8895,N_8708);
nor U9121 (N_9121,N_8885,N_8683);
or U9122 (N_9122,N_8964,N_8806);
nand U9123 (N_9123,N_8962,N_8563);
xnor U9124 (N_9124,N_8777,N_8721);
and U9125 (N_9125,N_8981,N_8931);
nand U9126 (N_9126,N_8631,N_8784);
nand U9127 (N_9127,N_8629,N_8668);
xor U9128 (N_9128,N_8851,N_8538);
or U9129 (N_9129,N_8558,N_8548);
nand U9130 (N_9130,N_8508,N_8586);
or U9131 (N_9131,N_8842,N_8849);
and U9132 (N_9132,N_8541,N_8636);
and U9133 (N_9133,N_8846,N_8531);
and U9134 (N_9134,N_8587,N_8609);
xor U9135 (N_9135,N_8642,N_8756);
or U9136 (N_9136,N_8976,N_8920);
nand U9137 (N_9137,N_8712,N_8652);
or U9138 (N_9138,N_8911,N_8518);
nor U9139 (N_9139,N_8655,N_8961);
nor U9140 (N_9140,N_8577,N_8943);
or U9141 (N_9141,N_8767,N_8867);
nand U9142 (N_9142,N_8889,N_8560);
nand U9143 (N_9143,N_8507,N_8775);
nand U9144 (N_9144,N_8628,N_8653);
nor U9145 (N_9145,N_8892,N_8522);
nor U9146 (N_9146,N_8571,N_8678);
or U9147 (N_9147,N_8868,N_8505);
xnor U9148 (N_9148,N_8697,N_8960);
nand U9149 (N_9149,N_8744,N_8718);
nand U9150 (N_9150,N_8843,N_8905);
nor U9151 (N_9151,N_8675,N_8994);
nand U9152 (N_9152,N_8719,N_8786);
nand U9153 (N_9153,N_8626,N_8822);
or U9154 (N_9154,N_8871,N_8984);
nand U9155 (N_9155,N_8914,N_8576);
and U9156 (N_9156,N_8788,N_8603);
nor U9157 (N_9157,N_8815,N_8809);
nand U9158 (N_9158,N_8755,N_8916);
or U9159 (N_9159,N_8734,N_8729);
nand U9160 (N_9160,N_8690,N_8979);
nor U9161 (N_9161,N_8891,N_8539);
nor U9162 (N_9162,N_8588,N_8811);
or U9163 (N_9163,N_8827,N_8870);
nand U9164 (N_9164,N_8528,N_8600);
xor U9165 (N_9165,N_8952,N_8785);
or U9166 (N_9166,N_8605,N_8699);
or U9167 (N_9167,N_8578,N_8929);
and U9168 (N_9168,N_8598,N_8589);
nor U9169 (N_9169,N_8903,N_8676);
xnor U9170 (N_9170,N_8924,N_8818);
or U9171 (N_9171,N_8936,N_8521);
or U9172 (N_9172,N_8574,N_8824);
and U9173 (N_9173,N_8801,N_8704);
nand U9174 (N_9174,N_8748,N_8794);
nand U9175 (N_9175,N_8884,N_8913);
nand U9176 (N_9176,N_8672,N_8673);
nor U9177 (N_9177,N_8536,N_8840);
or U9178 (N_9178,N_8742,N_8970);
nand U9179 (N_9179,N_8918,N_8977);
nor U9180 (N_9180,N_8887,N_8882);
and U9181 (N_9181,N_8779,N_8685);
and U9182 (N_9182,N_8783,N_8534);
or U9183 (N_9183,N_8746,N_8971);
or U9184 (N_9184,N_8796,N_8512);
nor U9185 (N_9185,N_8855,N_8798);
and U9186 (N_9186,N_8770,N_8864);
nand U9187 (N_9187,N_8782,N_8658);
nor U9188 (N_9188,N_8727,N_8754);
nor U9189 (N_9189,N_8687,N_8545);
xor U9190 (N_9190,N_8635,N_8679);
nand U9191 (N_9191,N_8987,N_8938);
or U9192 (N_9192,N_8932,N_8702);
nor U9193 (N_9193,N_8630,N_8526);
or U9194 (N_9194,N_8760,N_8967);
nor U9195 (N_9195,N_8949,N_8778);
nand U9196 (N_9196,N_8946,N_8634);
nor U9197 (N_9197,N_8516,N_8791);
nand U9198 (N_9198,N_8517,N_8886);
and U9199 (N_9199,N_8530,N_8661);
nand U9200 (N_9200,N_8990,N_8844);
nor U9201 (N_9201,N_8671,N_8597);
xor U9202 (N_9202,N_8944,N_8922);
nand U9203 (N_9203,N_8623,N_8726);
nor U9204 (N_9204,N_8696,N_8787);
nand U9205 (N_9205,N_8907,N_8735);
nor U9206 (N_9206,N_8733,N_8758);
nor U9207 (N_9207,N_8906,N_8863);
or U9208 (N_9208,N_8969,N_8781);
xnor U9209 (N_9209,N_8643,N_8559);
and U9210 (N_9210,N_8904,N_8680);
xor U9211 (N_9211,N_8511,N_8814);
nand U9212 (N_9212,N_8866,N_8845);
nand U9213 (N_9213,N_8768,N_8599);
or U9214 (N_9214,N_8974,N_8942);
nand U9215 (N_9215,N_8500,N_8832);
or U9216 (N_9216,N_8812,N_8555);
nor U9217 (N_9217,N_8869,N_8858);
or U9218 (N_9218,N_8857,N_8677);
nor U9219 (N_9219,N_8616,N_8835);
or U9220 (N_9220,N_8519,N_8921);
nor U9221 (N_9221,N_8732,N_8583);
and U9222 (N_9222,N_8854,N_8682);
nand U9223 (N_9223,N_8533,N_8640);
or U9224 (N_9224,N_8773,N_8769);
xnor U9225 (N_9225,N_8604,N_8647);
and U9226 (N_9226,N_8684,N_8780);
and U9227 (N_9227,N_8582,N_8692);
xnor U9228 (N_9228,N_8933,N_8831);
or U9229 (N_9229,N_8850,N_8537);
nand U9230 (N_9230,N_8700,N_8612);
and U9231 (N_9231,N_8910,N_8751);
nor U9232 (N_9232,N_8703,N_8654);
or U9233 (N_9233,N_8813,N_8989);
nand U9234 (N_9234,N_8876,N_8830);
nand U9235 (N_9235,N_8579,N_8561);
or U9236 (N_9236,N_8874,N_8701);
nand U9237 (N_9237,N_8566,N_8710);
and U9238 (N_9238,N_8838,N_8980);
and U9239 (N_9239,N_8880,N_8795);
nor U9240 (N_9240,N_8570,N_8550);
nand U9241 (N_9241,N_8602,N_8650);
nand U9242 (N_9242,N_8925,N_8689);
or U9243 (N_9243,N_8875,N_8873);
nor U9244 (N_9244,N_8713,N_8656);
and U9245 (N_9245,N_8955,N_8649);
xor U9246 (N_9246,N_8596,N_8621);
nand U9247 (N_9247,N_8509,N_8958);
and U9248 (N_9248,N_8937,N_8803);
nand U9249 (N_9249,N_8833,N_8506);
or U9250 (N_9250,N_8791,N_8765);
and U9251 (N_9251,N_8938,N_8983);
and U9252 (N_9252,N_8901,N_8710);
or U9253 (N_9253,N_8638,N_8781);
nand U9254 (N_9254,N_8688,N_8720);
or U9255 (N_9255,N_8628,N_8573);
or U9256 (N_9256,N_8878,N_8731);
nand U9257 (N_9257,N_8576,N_8508);
nor U9258 (N_9258,N_8615,N_8831);
and U9259 (N_9259,N_8828,N_8816);
nor U9260 (N_9260,N_8913,N_8980);
nor U9261 (N_9261,N_8645,N_8877);
nand U9262 (N_9262,N_8508,N_8668);
nor U9263 (N_9263,N_8950,N_8922);
and U9264 (N_9264,N_8597,N_8804);
xor U9265 (N_9265,N_8910,N_8846);
or U9266 (N_9266,N_8863,N_8714);
and U9267 (N_9267,N_8840,N_8770);
nor U9268 (N_9268,N_8789,N_8880);
nand U9269 (N_9269,N_8610,N_8874);
and U9270 (N_9270,N_8569,N_8638);
nand U9271 (N_9271,N_8958,N_8698);
nand U9272 (N_9272,N_8834,N_8872);
nor U9273 (N_9273,N_8533,N_8809);
nand U9274 (N_9274,N_8914,N_8683);
or U9275 (N_9275,N_8810,N_8790);
nand U9276 (N_9276,N_8704,N_8814);
nor U9277 (N_9277,N_8514,N_8753);
nand U9278 (N_9278,N_8628,N_8735);
nand U9279 (N_9279,N_8734,N_8666);
and U9280 (N_9280,N_8863,N_8982);
and U9281 (N_9281,N_8782,N_8834);
xor U9282 (N_9282,N_8768,N_8942);
xor U9283 (N_9283,N_8928,N_8504);
nand U9284 (N_9284,N_8900,N_8619);
nor U9285 (N_9285,N_8651,N_8741);
or U9286 (N_9286,N_8848,N_8998);
or U9287 (N_9287,N_8517,N_8725);
or U9288 (N_9288,N_8728,N_8510);
and U9289 (N_9289,N_8682,N_8750);
and U9290 (N_9290,N_8527,N_8720);
xor U9291 (N_9291,N_8529,N_8881);
and U9292 (N_9292,N_8635,N_8916);
or U9293 (N_9293,N_8842,N_8512);
and U9294 (N_9294,N_8697,N_8986);
or U9295 (N_9295,N_8953,N_8832);
or U9296 (N_9296,N_8569,N_8792);
nor U9297 (N_9297,N_8929,N_8909);
and U9298 (N_9298,N_8777,N_8956);
and U9299 (N_9299,N_8550,N_8661);
nand U9300 (N_9300,N_8928,N_8715);
nand U9301 (N_9301,N_8751,N_8575);
or U9302 (N_9302,N_8938,N_8618);
nand U9303 (N_9303,N_8922,N_8633);
xnor U9304 (N_9304,N_8924,N_8981);
nor U9305 (N_9305,N_8835,N_8830);
or U9306 (N_9306,N_8885,N_8555);
xnor U9307 (N_9307,N_8670,N_8655);
nor U9308 (N_9308,N_8823,N_8712);
or U9309 (N_9309,N_8503,N_8885);
and U9310 (N_9310,N_8572,N_8886);
and U9311 (N_9311,N_8833,N_8970);
xor U9312 (N_9312,N_8967,N_8945);
and U9313 (N_9313,N_8847,N_8643);
nand U9314 (N_9314,N_8783,N_8779);
nor U9315 (N_9315,N_8848,N_8920);
xnor U9316 (N_9316,N_8976,N_8921);
nor U9317 (N_9317,N_8838,N_8643);
or U9318 (N_9318,N_8974,N_8612);
or U9319 (N_9319,N_8567,N_8562);
xor U9320 (N_9320,N_8967,N_8516);
and U9321 (N_9321,N_8955,N_8657);
nand U9322 (N_9322,N_8935,N_8976);
xnor U9323 (N_9323,N_8752,N_8569);
nor U9324 (N_9324,N_8841,N_8912);
and U9325 (N_9325,N_8710,N_8567);
and U9326 (N_9326,N_8771,N_8717);
or U9327 (N_9327,N_8864,N_8863);
and U9328 (N_9328,N_8713,N_8912);
or U9329 (N_9329,N_8741,N_8660);
nor U9330 (N_9330,N_8780,N_8578);
nand U9331 (N_9331,N_8552,N_8867);
and U9332 (N_9332,N_8916,N_8672);
nand U9333 (N_9333,N_8827,N_8793);
and U9334 (N_9334,N_8814,N_8700);
nand U9335 (N_9335,N_8746,N_8547);
and U9336 (N_9336,N_8753,N_8583);
or U9337 (N_9337,N_8854,N_8813);
nor U9338 (N_9338,N_8624,N_8505);
and U9339 (N_9339,N_8553,N_8587);
and U9340 (N_9340,N_8800,N_8973);
nor U9341 (N_9341,N_8968,N_8910);
or U9342 (N_9342,N_8631,N_8646);
nand U9343 (N_9343,N_8542,N_8941);
nor U9344 (N_9344,N_8948,N_8831);
xor U9345 (N_9345,N_8760,N_8808);
nor U9346 (N_9346,N_8508,N_8547);
or U9347 (N_9347,N_8871,N_8967);
or U9348 (N_9348,N_8664,N_8749);
xor U9349 (N_9349,N_8823,N_8825);
and U9350 (N_9350,N_8865,N_8588);
and U9351 (N_9351,N_8917,N_8858);
xor U9352 (N_9352,N_8886,N_8660);
nor U9353 (N_9353,N_8833,N_8937);
nor U9354 (N_9354,N_8668,N_8798);
nand U9355 (N_9355,N_8773,N_8624);
or U9356 (N_9356,N_8811,N_8591);
nor U9357 (N_9357,N_8913,N_8531);
nor U9358 (N_9358,N_8735,N_8848);
nor U9359 (N_9359,N_8555,N_8700);
or U9360 (N_9360,N_8704,N_8536);
xor U9361 (N_9361,N_8839,N_8917);
nor U9362 (N_9362,N_8604,N_8750);
xnor U9363 (N_9363,N_8797,N_8941);
nand U9364 (N_9364,N_8520,N_8713);
or U9365 (N_9365,N_8674,N_8812);
or U9366 (N_9366,N_8516,N_8539);
and U9367 (N_9367,N_8756,N_8701);
or U9368 (N_9368,N_8707,N_8558);
or U9369 (N_9369,N_8659,N_8839);
xor U9370 (N_9370,N_8958,N_8510);
nor U9371 (N_9371,N_8835,N_8572);
xor U9372 (N_9372,N_8685,N_8895);
nand U9373 (N_9373,N_8613,N_8861);
nor U9374 (N_9374,N_8705,N_8608);
and U9375 (N_9375,N_8520,N_8684);
nand U9376 (N_9376,N_8715,N_8843);
xor U9377 (N_9377,N_8529,N_8963);
or U9378 (N_9378,N_8854,N_8889);
or U9379 (N_9379,N_8556,N_8946);
and U9380 (N_9380,N_8560,N_8847);
nand U9381 (N_9381,N_8861,N_8803);
xor U9382 (N_9382,N_8987,N_8917);
nor U9383 (N_9383,N_8650,N_8882);
or U9384 (N_9384,N_8703,N_8847);
nor U9385 (N_9385,N_8728,N_8616);
and U9386 (N_9386,N_8703,N_8652);
nor U9387 (N_9387,N_8616,N_8829);
and U9388 (N_9388,N_8769,N_8543);
or U9389 (N_9389,N_8751,N_8643);
nand U9390 (N_9390,N_8790,N_8851);
or U9391 (N_9391,N_8811,N_8662);
and U9392 (N_9392,N_8532,N_8742);
nand U9393 (N_9393,N_8567,N_8793);
or U9394 (N_9394,N_8673,N_8917);
xor U9395 (N_9395,N_8764,N_8992);
nand U9396 (N_9396,N_8901,N_8846);
nand U9397 (N_9397,N_8748,N_8793);
or U9398 (N_9398,N_8537,N_8578);
nand U9399 (N_9399,N_8650,N_8930);
or U9400 (N_9400,N_8641,N_8678);
nor U9401 (N_9401,N_8882,N_8960);
nor U9402 (N_9402,N_8995,N_8542);
and U9403 (N_9403,N_8972,N_8871);
nor U9404 (N_9404,N_8602,N_8717);
and U9405 (N_9405,N_8811,N_8919);
or U9406 (N_9406,N_8996,N_8539);
nor U9407 (N_9407,N_8527,N_8513);
or U9408 (N_9408,N_8983,N_8572);
nor U9409 (N_9409,N_8549,N_8746);
and U9410 (N_9410,N_8619,N_8890);
nor U9411 (N_9411,N_8550,N_8920);
xor U9412 (N_9412,N_8968,N_8679);
and U9413 (N_9413,N_8582,N_8885);
nand U9414 (N_9414,N_8755,N_8693);
or U9415 (N_9415,N_8911,N_8940);
nor U9416 (N_9416,N_8537,N_8628);
or U9417 (N_9417,N_8920,N_8707);
nand U9418 (N_9418,N_8636,N_8714);
and U9419 (N_9419,N_8679,N_8868);
nor U9420 (N_9420,N_8615,N_8852);
and U9421 (N_9421,N_8738,N_8661);
and U9422 (N_9422,N_8518,N_8736);
and U9423 (N_9423,N_8697,N_8648);
nand U9424 (N_9424,N_8811,N_8729);
nand U9425 (N_9425,N_8715,N_8982);
and U9426 (N_9426,N_8611,N_8635);
or U9427 (N_9427,N_8696,N_8948);
or U9428 (N_9428,N_8756,N_8728);
nand U9429 (N_9429,N_8622,N_8937);
and U9430 (N_9430,N_8824,N_8518);
nand U9431 (N_9431,N_8908,N_8723);
nor U9432 (N_9432,N_8518,N_8524);
nand U9433 (N_9433,N_8917,N_8829);
nand U9434 (N_9434,N_8941,N_8849);
nor U9435 (N_9435,N_8582,N_8892);
nor U9436 (N_9436,N_8682,N_8534);
nor U9437 (N_9437,N_8726,N_8779);
or U9438 (N_9438,N_8514,N_8654);
nor U9439 (N_9439,N_8751,N_8773);
and U9440 (N_9440,N_8761,N_8927);
and U9441 (N_9441,N_8537,N_8839);
nor U9442 (N_9442,N_8833,N_8632);
xnor U9443 (N_9443,N_8751,N_8800);
nor U9444 (N_9444,N_8724,N_8833);
xor U9445 (N_9445,N_8545,N_8676);
or U9446 (N_9446,N_8577,N_8986);
nand U9447 (N_9447,N_8818,N_8749);
or U9448 (N_9448,N_8811,N_8599);
and U9449 (N_9449,N_8901,N_8597);
nor U9450 (N_9450,N_8814,N_8524);
nor U9451 (N_9451,N_8918,N_8623);
nor U9452 (N_9452,N_8599,N_8547);
and U9453 (N_9453,N_8611,N_8552);
nor U9454 (N_9454,N_8566,N_8902);
nor U9455 (N_9455,N_8637,N_8542);
nand U9456 (N_9456,N_8704,N_8504);
and U9457 (N_9457,N_8727,N_8607);
nand U9458 (N_9458,N_8707,N_8907);
nand U9459 (N_9459,N_8907,N_8507);
or U9460 (N_9460,N_8538,N_8521);
and U9461 (N_9461,N_8639,N_8841);
and U9462 (N_9462,N_8641,N_8739);
and U9463 (N_9463,N_8538,N_8501);
nand U9464 (N_9464,N_8801,N_8691);
nor U9465 (N_9465,N_8927,N_8922);
and U9466 (N_9466,N_8643,N_8594);
or U9467 (N_9467,N_8717,N_8823);
nand U9468 (N_9468,N_8998,N_8689);
nor U9469 (N_9469,N_8896,N_8538);
nor U9470 (N_9470,N_8993,N_8515);
or U9471 (N_9471,N_8567,N_8708);
or U9472 (N_9472,N_8540,N_8527);
nor U9473 (N_9473,N_8519,N_8527);
nand U9474 (N_9474,N_8619,N_8852);
nor U9475 (N_9475,N_8655,N_8946);
nor U9476 (N_9476,N_8597,N_8653);
and U9477 (N_9477,N_8817,N_8562);
and U9478 (N_9478,N_8507,N_8872);
xor U9479 (N_9479,N_8636,N_8692);
or U9480 (N_9480,N_8976,N_8741);
and U9481 (N_9481,N_8685,N_8818);
nor U9482 (N_9482,N_8744,N_8616);
nand U9483 (N_9483,N_8784,N_8521);
nand U9484 (N_9484,N_8739,N_8563);
nor U9485 (N_9485,N_8952,N_8953);
and U9486 (N_9486,N_8808,N_8511);
nor U9487 (N_9487,N_8872,N_8816);
and U9488 (N_9488,N_8896,N_8550);
nor U9489 (N_9489,N_8989,N_8738);
and U9490 (N_9490,N_8864,N_8631);
nand U9491 (N_9491,N_8717,N_8903);
nand U9492 (N_9492,N_8898,N_8808);
xor U9493 (N_9493,N_8583,N_8907);
and U9494 (N_9494,N_8651,N_8919);
and U9495 (N_9495,N_8847,N_8629);
and U9496 (N_9496,N_8614,N_8604);
and U9497 (N_9497,N_8751,N_8739);
or U9498 (N_9498,N_8714,N_8991);
nor U9499 (N_9499,N_8608,N_8728);
and U9500 (N_9500,N_9102,N_9201);
nor U9501 (N_9501,N_9329,N_9082);
nor U9502 (N_9502,N_9096,N_9214);
nor U9503 (N_9503,N_9014,N_9033);
nor U9504 (N_9504,N_9177,N_9195);
or U9505 (N_9505,N_9018,N_9205);
nand U9506 (N_9506,N_9352,N_9489);
and U9507 (N_9507,N_9274,N_9200);
nand U9508 (N_9508,N_9485,N_9447);
nand U9509 (N_9509,N_9106,N_9460);
nand U9510 (N_9510,N_9377,N_9025);
nor U9511 (N_9511,N_9168,N_9066);
and U9512 (N_9512,N_9438,N_9349);
nand U9513 (N_9513,N_9246,N_9067);
nor U9514 (N_9514,N_9084,N_9367);
xor U9515 (N_9515,N_9334,N_9170);
nand U9516 (N_9516,N_9134,N_9482);
nand U9517 (N_9517,N_9258,N_9187);
and U9518 (N_9518,N_9426,N_9346);
nor U9519 (N_9519,N_9281,N_9494);
and U9520 (N_9520,N_9287,N_9468);
xnor U9521 (N_9521,N_9462,N_9213);
nand U9522 (N_9522,N_9094,N_9178);
nor U9523 (N_9523,N_9105,N_9010);
and U9524 (N_9524,N_9384,N_9415);
or U9525 (N_9525,N_9189,N_9356);
nand U9526 (N_9526,N_9408,N_9282);
or U9527 (N_9527,N_9028,N_9296);
and U9528 (N_9528,N_9219,N_9365);
nor U9529 (N_9529,N_9484,N_9027);
nand U9530 (N_9530,N_9459,N_9319);
xor U9531 (N_9531,N_9416,N_9076);
and U9532 (N_9532,N_9073,N_9292);
or U9533 (N_9533,N_9295,N_9256);
and U9534 (N_9534,N_9398,N_9095);
and U9535 (N_9535,N_9361,N_9330);
and U9536 (N_9536,N_9140,N_9357);
and U9537 (N_9537,N_9444,N_9031);
nand U9538 (N_9538,N_9314,N_9171);
or U9539 (N_9539,N_9491,N_9071);
and U9540 (N_9540,N_9045,N_9126);
nor U9541 (N_9541,N_9005,N_9032);
and U9542 (N_9542,N_9022,N_9407);
and U9543 (N_9543,N_9254,N_9222);
nor U9544 (N_9544,N_9078,N_9391);
nand U9545 (N_9545,N_9363,N_9336);
nand U9546 (N_9546,N_9308,N_9089);
nor U9547 (N_9547,N_9276,N_9477);
and U9548 (N_9548,N_9372,N_9364);
nor U9549 (N_9549,N_9184,N_9211);
nand U9550 (N_9550,N_9232,N_9449);
xor U9551 (N_9551,N_9175,N_9011);
nand U9552 (N_9552,N_9297,N_9463);
nand U9553 (N_9553,N_9075,N_9218);
nand U9554 (N_9554,N_9496,N_9320);
or U9555 (N_9555,N_9470,N_9107);
and U9556 (N_9556,N_9172,N_9412);
and U9557 (N_9557,N_9238,N_9202);
nor U9558 (N_9558,N_9400,N_9261);
and U9559 (N_9559,N_9008,N_9047);
nand U9560 (N_9560,N_9240,N_9247);
or U9561 (N_9561,N_9471,N_9006);
xnor U9562 (N_9562,N_9341,N_9225);
or U9563 (N_9563,N_9486,N_9139);
and U9564 (N_9564,N_9237,N_9059);
or U9565 (N_9565,N_9467,N_9118);
and U9566 (N_9566,N_9410,N_9393);
and U9567 (N_9567,N_9191,N_9166);
nor U9568 (N_9568,N_9186,N_9252);
nand U9569 (N_9569,N_9298,N_9358);
nor U9570 (N_9570,N_9279,N_9019);
nor U9571 (N_9571,N_9098,N_9419);
nand U9572 (N_9572,N_9239,N_9079);
nand U9573 (N_9573,N_9249,N_9072);
or U9574 (N_9574,N_9268,N_9023);
nor U9575 (N_9575,N_9145,N_9390);
or U9576 (N_9576,N_9348,N_9355);
or U9577 (N_9577,N_9004,N_9149);
or U9578 (N_9578,N_9192,N_9487);
or U9579 (N_9579,N_9473,N_9453);
and U9580 (N_9580,N_9403,N_9037);
and U9581 (N_9581,N_9425,N_9262);
nand U9582 (N_9582,N_9051,N_9490);
or U9583 (N_9583,N_9446,N_9136);
nand U9584 (N_9584,N_9307,N_9378);
and U9585 (N_9585,N_9411,N_9338);
nor U9586 (N_9586,N_9212,N_9266);
nor U9587 (N_9587,N_9120,N_9207);
or U9588 (N_9588,N_9369,N_9452);
nand U9589 (N_9589,N_9235,N_9324);
or U9590 (N_9590,N_9381,N_9479);
nor U9591 (N_9591,N_9049,N_9360);
nand U9592 (N_9592,N_9480,N_9414);
nand U9593 (N_9593,N_9432,N_9242);
nor U9594 (N_9594,N_9316,N_9302);
and U9595 (N_9595,N_9038,N_9183);
and U9596 (N_9596,N_9339,N_9443);
and U9597 (N_9597,N_9228,N_9472);
and U9598 (N_9598,N_9215,N_9041);
nor U9599 (N_9599,N_9318,N_9128);
or U9600 (N_9600,N_9269,N_9176);
and U9601 (N_9601,N_9163,N_9280);
nor U9602 (N_9602,N_9223,N_9430);
and U9603 (N_9603,N_9345,N_9376);
nor U9604 (N_9604,N_9000,N_9193);
or U9605 (N_9605,N_9224,N_9284);
and U9606 (N_9606,N_9208,N_9030);
or U9607 (N_9607,N_9115,N_9283);
or U9608 (N_9608,N_9185,N_9405);
or U9609 (N_9609,N_9423,N_9399);
nand U9610 (N_9610,N_9179,N_9257);
and U9611 (N_9611,N_9464,N_9481);
or U9612 (N_9612,N_9090,N_9270);
or U9613 (N_9613,N_9271,N_9289);
and U9614 (N_9614,N_9001,N_9233);
and U9615 (N_9615,N_9035,N_9497);
nand U9616 (N_9616,N_9164,N_9131);
xor U9617 (N_9617,N_9099,N_9043);
nor U9618 (N_9618,N_9231,N_9182);
nand U9619 (N_9619,N_9150,N_9431);
nand U9620 (N_9620,N_9161,N_9190);
nor U9621 (N_9621,N_9456,N_9125);
and U9622 (N_9622,N_9110,N_9124);
nor U9623 (N_9623,N_9229,N_9148);
nand U9624 (N_9624,N_9162,N_9077);
nor U9625 (N_9625,N_9340,N_9159);
nand U9626 (N_9626,N_9379,N_9042);
nand U9627 (N_9627,N_9152,N_9108);
or U9628 (N_9628,N_9109,N_9112);
and U9629 (N_9629,N_9389,N_9442);
xnor U9630 (N_9630,N_9044,N_9100);
or U9631 (N_9631,N_9333,N_9243);
nor U9632 (N_9632,N_9209,N_9331);
or U9633 (N_9633,N_9306,N_9475);
nor U9634 (N_9634,N_9437,N_9458);
xnor U9635 (N_9635,N_9450,N_9169);
xnor U9636 (N_9636,N_9344,N_9068);
and U9637 (N_9637,N_9127,N_9465);
and U9638 (N_9638,N_9111,N_9310);
nor U9639 (N_9639,N_9013,N_9315);
xor U9640 (N_9640,N_9382,N_9245);
nor U9641 (N_9641,N_9409,N_9080);
and U9642 (N_9642,N_9373,N_9495);
nand U9643 (N_9643,N_9074,N_9064);
or U9644 (N_9644,N_9267,N_9278);
or U9645 (N_9645,N_9137,N_9180);
nand U9646 (N_9646,N_9198,N_9288);
and U9647 (N_9647,N_9337,N_9040);
nand U9648 (N_9648,N_9474,N_9368);
or U9649 (N_9649,N_9113,N_9466);
nor U9650 (N_9650,N_9101,N_9359);
or U9651 (N_9651,N_9396,N_9386);
nand U9652 (N_9652,N_9050,N_9142);
or U9653 (N_9653,N_9081,N_9234);
and U9654 (N_9654,N_9092,N_9220);
nand U9655 (N_9655,N_9053,N_9476);
and U9656 (N_9656,N_9328,N_9158);
and U9657 (N_9657,N_9498,N_9342);
nand U9658 (N_9658,N_9350,N_9291);
nand U9659 (N_9659,N_9293,N_9427);
and U9660 (N_9660,N_9285,N_9087);
and U9661 (N_9661,N_9146,N_9129);
nand U9662 (N_9662,N_9353,N_9277);
or U9663 (N_9663,N_9194,N_9060);
nand U9664 (N_9664,N_9133,N_9457);
nor U9665 (N_9665,N_9230,N_9394);
nand U9666 (N_9666,N_9418,N_9086);
or U9667 (N_9667,N_9065,N_9039);
nand U9668 (N_9668,N_9174,N_9070);
xor U9669 (N_9669,N_9313,N_9097);
nand U9670 (N_9670,N_9299,N_9196);
and U9671 (N_9671,N_9251,N_9123);
nand U9672 (N_9672,N_9250,N_9448);
and U9673 (N_9673,N_9454,N_9451);
and U9674 (N_9674,N_9499,N_9088);
or U9675 (N_9675,N_9343,N_9304);
nor U9676 (N_9676,N_9488,N_9317);
xor U9677 (N_9677,N_9007,N_9144);
nor U9678 (N_9678,N_9156,N_9428);
nand U9679 (N_9679,N_9199,N_9221);
nor U9680 (N_9680,N_9439,N_9305);
and U9681 (N_9681,N_9483,N_9009);
nand U9682 (N_9682,N_9052,N_9138);
xor U9683 (N_9683,N_9012,N_9354);
and U9684 (N_9684,N_9311,N_9054);
and U9685 (N_9685,N_9021,N_9058);
and U9686 (N_9686,N_9434,N_9024);
nor U9687 (N_9687,N_9347,N_9327);
and U9688 (N_9688,N_9263,N_9273);
and U9689 (N_9689,N_9083,N_9121);
or U9690 (N_9690,N_9433,N_9217);
or U9691 (N_9691,N_9181,N_9445);
xor U9692 (N_9692,N_9401,N_9119);
or U9693 (N_9693,N_9167,N_9265);
nand U9694 (N_9694,N_9244,N_9026);
and U9695 (N_9695,N_9420,N_9093);
and U9696 (N_9696,N_9264,N_9335);
or U9697 (N_9697,N_9141,N_9303);
nor U9698 (N_9698,N_9272,N_9160);
and U9699 (N_9699,N_9241,N_9421);
or U9700 (N_9700,N_9029,N_9154);
xor U9701 (N_9701,N_9061,N_9062);
nor U9702 (N_9702,N_9204,N_9056);
nor U9703 (N_9703,N_9383,N_9114);
or U9704 (N_9704,N_9020,N_9469);
nor U9705 (N_9705,N_9157,N_9290);
nand U9706 (N_9706,N_9063,N_9255);
nand U9707 (N_9707,N_9455,N_9371);
or U9708 (N_9708,N_9332,N_9402);
xnor U9709 (N_9709,N_9103,N_9322);
xor U9710 (N_9710,N_9435,N_9493);
xor U9711 (N_9711,N_9300,N_9362);
nand U9712 (N_9712,N_9206,N_9151);
and U9713 (N_9713,N_9392,N_9321);
and U9714 (N_9714,N_9003,N_9260);
and U9715 (N_9715,N_9397,N_9380);
nand U9716 (N_9716,N_9351,N_9301);
xnor U9717 (N_9717,N_9326,N_9441);
nor U9718 (N_9718,N_9227,N_9461);
and U9719 (N_9719,N_9057,N_9203);
xnor U9720 (N_9720,N_9036,N_9424);
nor U9721 (N_9721,N_9429,N_9370);
nor U9722 (N_9722,N_9034,N_9153);
or U9723 (N_9723,N_9155,N_9286);
and U9724 (N_9724,N_9165,N_9002);
nand U9725 (N_9725,N_9236,N_9122);
nand U9726 (N_9726,N_9132,N_9135);
and U9727 (N_9727,N_9406,N_9404);
nand U9728 (N_9728,N_9259,N_9374);
xnor U9729 (N_9729,N_9325,N_9248);
nor U9730 (N_9730,N_9069,N_9323);
xor U9731 (N_9731,N_9375,N_9226);
and U9732 (N_9732,N_9388,N_9117);
nand U9733 (N_9733,N_9417,N_9436);
and U9734 (N_9734,N_9143,N_9216);
nand U9735 (N_9735,N_9440,N_9275);
nand U9736 (N_9736,N_9210,N_9309);
or U9737 (N_9737,N_9085,N_9173);
or U9738 (N_9738,N_9046,N_9015);
and U9739 (N_9739,N_9130,N_9422);
nor U9740 (N_9740,N_9091,N_9253);
nor U9741 (N_9741,N_9366,N_9294);
xnor U9742 (N_9742,N_9312,N_9116);
nor U9743 (N_9743,N_9016,N_9188);
or U9744 (N_9744,N_9017,N_9413);
nand U9745 (N_9745,N_9197,N_9492);
nand U9746 (N_9746,N_9478,N_9387);
nand U9747 (N_9747,N_9385,N_9147);
and U9748 (N_9748,N_9104,N_9055);
and U9749 (N_9749,N_9048,N_9395);
nor U9750 (N_9750,N_9394,N_9101);
and U9751 (N_9751,N_9100,N_9011);
nand U9752 (N_9752,N_9177,N_9363);
nand U9753 (N_9753,N_9468,N_9393);
or U9754 (N_9754,N_9140,N_9472);
nand U9755 (N_9755,N_9173,N_9401);
or U9756 (N_9756,N_9175,N_9378);
and U9757 (N_9757,N_9207,N_9398);
and U9758 (N_9758,N_9041,N_9060);
nor U9759 (N_9759,N_9104,N_9200);
xnor U9760 (N_9760,N_9339,N_9234);
and U9761 (N_9761,N_9203,N_9410);
xor U9762 (N_9762,N_9473,N_9202);
and U9763 (N_9763,N_9469,N_9042);
and U9764 (N_9764,N_9092,N_9205);
or U9765 (N_9765,N_9090,N_9336);
and U9766 (N_9766,N_9468,N_9255);
nor U9767 (N_9767,N_9003,N_9026);
nor U9768 (N_9768,N_9372,N_9265);
nand U9769 (N_9769,N_9215,N_9473);
and U9770 (N_9770,N_9115,N_9463);
or U9771 (N_9771,N_9091,N_9345);
or U9772 (N_9772,N_9261,N_9059);
xnor U9773 (N_9773,N_9086,N_9248);
and U9774 (N_9774,N_9158,N_9015);
or U9775 (N_9775,N_9158,N_9267);
and U9776 (N_9776,N_9185,N_9217);
nor U9777 (N_9777,N_9079,N_9203);
or U9778 (N_9778,N_9463,N_9177);
nand U9779 (N_9779,N_9442,N_9350);
and U9780 (N_9780,N_9101,N_9377);
and U9781 (N_9781,N_9275,N_9364);
nand U9782 (N_9782,N_9425,N_9422);
or U9783 (N_9783,N_9315,N_9015);
and U9784 (N_9784,N_9082,N_9301);
xnor U9785 (N_9785,N_9234,N_9376);
and U9786 (N_9786,N_9008,N_9094);
nand U9787 (N_9787,N_9120,N_9442);
xnor U9788 (N_9788,N_9051,N_9202);
nor U9789 (N_9789,N_9184,N_9002);
or U9790 (N_9790,N_9394,N_9133);
nand U9791 (N_9791,N_9046,N_9344);
nand U9792 (N_9792,N_9240,N_9075);
nand U9793 (N_9793,N_9187,N_9068);
or U9794 (N_9794,N_9154,N_9397);
nor U9795 (N_9795,N_9038,N_9388);
or U9796 (N_9796,N_9347,N_9110);
and U9797 (N_9797,N_9328,N_9267);
nand U9798 (N_9798,N_9431,N_9112);
or U9799 (N_9799,N_9208,N_9369);
nand U9800 (N_9800,N_9162,N_9161);
or U9801 (N_9801,N_9202,N_9241);
or U9802 (N_9802,N_9205,N_9428);
nor U9803 (N_9803,N_9324,N_9396);
nand U9804 (N_9804,N_9250,N_9311);
nor U9805 (N_9805,N_9008,N_9254);
nor U9806 (N_9806,N_9111,N_9198);
or U9807 (N_9807,N_9375,N_9307);
xor U9808 (N_9808,N_9324,N_9473);
and U9809 (N_9809,N_9238,N_9289);
or U9810 (N_9810,N_9045,N_9333);
and U9811 (N_9811,N_9479,N_9079);
and U9812 (N_9812,N_9399,N_9416);
nor U9813 (N_9813,N_9103,N_9405);
and U9814 (N_9814,N_9497,N_9399);
or U9815 (N_9815,N_9199,N_9228);
nand U9816 (N_9816,N_9464,N_9442);
or U9817 (N_9817,N_9282,N_9021);
nor U9818 (N_9818,N_9275,N_9435);
xor U9819 (N_9819,N_9044,N_9094);
nand U9820 (N_9820,N_9275,N_9084);
nor U9821 (N_9821,N_9200,N_9392);
xor U9822 (N_9822,N_9478,N_9127);
nand U9823 (N_9823,N_9389,N_9455);
nand U9824 (N_9824,N_9118,N_9446);
nor U9825 (N_9825,N_9098,N_9036);
nor U9826 (N_9826,N_9345,N_9412);
or U9827 (N_9827,N_9387,N_9453);
or U9828 (N_9828,N_9334,N_9406);
xnor U9829 (N_9829,N_9401,N_9360);
nor U9830 (N_9830,N_9492,N_9097);
or U9831 (N_9831,N_9368,N_9250);
and U9832 (N_9832,N_9242,N_9422);
and U9833 (N_9833,N_9288,N_9385);
nand U9834 (N_9834,N_9066,N_9133);
or U9835 (N_9835,N_9466,N_9220);
and U9836 (N_9836,N_9028,N_9053);
or U9837 (N_9837,N_9094,N_9060);
nor U9838 (N_9838,N_9400,N_9009);
and U9839 (N_9839,N_9240,N_9074);
and U9840 (N_9840,N_9175,N_9395);
or U9841 (N_9841,N_9317,N_9282);
xnor U9842 (N_9842,N_9206,N_9308);
nor U9843 (N_9843,N_9265,N_9332);
nand U9844 (N_9844,N_9489,N_9315);
xor U9845 (N_9845,N_9421,N_9054);
or U9846 (N_9846,N_9406,N_9416);
or U9847 (N_9847,N_9053,N_9188);
nor U9848 (N_9848,N_9332,N_9279);
or U9849 (N_9849,N_9127,N_9345);
nor U9850 (N_9850,N_9055,N_9380);
xor U9851 (N_9851,N_9299,N_9213);
or U9852 (N_9852,N_9397,N_9007);
and U9853 (N_9853,N_9005,N_9186);
nor U9854 (N_9854,N_9242,N_9048);
nor U9855 (N_9855,N_9104,N_9125);
or U9856 (N_9856,N_9492,N_9481);
nor U9857 (N_9857,N_9124,N_9287);
nand U9858 (N_9858,N_9096,N_9437);
and U9859 (N_9859,N_9041,N_9366);
nor U9860 (N_9860,N_9469,N_9152);
nand U9861 (N_9861,N_9061,N_9192);
or U9862 (N_9862,N_9065,N_9254);
nand U9863 (N_9863,N_9011,N_9494);
nor U9864 (N_9864,N_9302,N_9297);
and U9865 (N_9865,N_9021,N_9390);
or U9866 (N_9866,N_9411,N_9099);
nand U9867 (N_9867,N_9007,N_9420);
nand U9868 (N_9868,N_9481,N_9388);
and U9869 (N_9869,N_9190,N_9421);
nand U9870 (N_9870,N_9144,N_9355);
or U9871 (N_9871,N_9461,N_9210);
nand U9872 (N_9872,N_9223,N_9167);
or U9873 (N_9873,N_9252,N_9124);
and U9874 (N_9874,N_9443,N_9364);
or U9875 (N_9875,N_9220,N_9212);
and U9876 (N_9876,N_9132,N_9442);
and U9877 (N_9877,N_9233,N_9248);
xnor U9878 (N_9878,N_9487,N_9340);
nor U9879 (N_9879,N_9285,N_9192);
or U9880 (N_9880,N_9287,N_9102);
or U9881 (N_9881,N_9305,N_9496);
and U9882 (N_9882,N_9445,N_9379);
or U9883 (N_9883,N_9364,N_9403);
nor U9884 (N_9884,N_9384,N_9330);
and U9885 (N_9885,N_9298,N_9094);
or U9886 (N_9886,N_9191,N_9432);
or U9887 (N_9887,N_9396,N_9000);
or U9888 (N_9888,N_9438,N_9045);
nand U9889 (N_9889,N_9375,N_9099);
nand U9890 (N_9890,N_9423,N_9155);
xor U9891 (N_9891,N_9400,N_9340);
or U9892 (N_9892,N_9109,N_9013);
nand U9893 (N_9893,N_9258,N_9284);
nor U9894 (N_9894,N_9123,N_9170);
nor U9895 (N_9895,N_9338,N_9379);
or U9896 (N_9896,N_9121,N_9476);
xor U9897 (N_9897,N_9360,N_9166);
and U9898 (N_9898,N_9211,N_9439);
nand U9899 (N_9899,N_9424,N_9491);
or U9900 (N_9900,N_9361,N_9112);
or U9901 (N_9901,N_9372,N_9439);
or U9902 (N_9902,N_9067,N_9185);
and U9903 (N_9903,N_9291,N_9302);
nor U9904 (N_9904,N_9040,N_9463);
or U9905 (N_9905,N_9349,N_9310);
xor U9906 (N_9906,N_9477,N_9168);
and U9907 (N_9907,N_9129,N_9199);
nand U9908 (N_9908,N_9460,N_9378);
or U9909 (N_9909,N_9065,N_9020);
nor U9910 (N_9910,N_9173,N_9450);
and U9911 (N_9911,N_9116,N_9305);
nand U9912 (N_9912,N_9221,N_9154);
xnor U9913 (N_9913,N_9334,N_9434);
and U9914 (N_9914,N_9243,N_9229);
nor U9915 (N_9915,N_9366,N_9317);
nand U9916 (N_9916,N_9400,N_9199);
nand U9917 (N_9917,N_9233,N_9134);
nand U9918 (N_9918,N_9268,N_9017);
nand U9919 (N_9919,N_9156,N_9367);
and U9920 (N_9920,N_9253,N_9485);
nand U9921 (N_9921,N_9469,N_9316);
and U9922 (N_9922,N_9028,N_9099);
nor U9923 (N_9923,N_9072,N_9024);
nor U9924 (N_9924,N_9133,N_9225);
nor U9925 (N_9925,N_9267,N_9045);
nand U9926 (N_9926,N_9131,N_9069);
or U9927 (N_9927,N_9184,N_9244);
and U9928 (N_9928,N_9340,N_9369);
or U9929 (N_9929,N_9113,N_9242);
or U9930 (N_9930,N_9479,N_9208);
and U9931 (N_9931,N_9251,N_9099);
nand U9932 (N_9932,N_9027,N_9366);
nor U9933 (N_9933,N_9016,N_9060);
nand U9934 (N_9934,N_9123,N_9136);
and U9935 (N_9935,N_9090,N_9296);
or U9936 (N_9936,N_9138,N_9005);
nand U9937 (N_9937,N_9057,N_9161);
or U9938 (N_9938,N_9139,N_9222);
and U9939 (N_9939,N_9042,N_9087);
or U9940 (N_9940,N_9466,N_9104);
nand U9941 (N_9941,N_9242,N_9015);
nand U9942 (N_9942,N_9225,N_9156);
nor U9943 (N_9943,N_9196,N_9101);
nand U9944 (N_9944,N_9348,N_9170);
nor U9945 (N_9945,N_9280,N_9491);
xor U9946 (N_9946,N_9376,N_9148);
and U9947 (N_9947,N_9473,N_9221);
or U9948 (N_9948,N_9322,N_9237);
nand U9949 (N_9949,N_9049,N_9313);
xor U9950 (N_9950,N_9007,N_9423);
and U9951 (N_9951,N_9433,N_9098);
and U9952 (N_9952,N_9268,N_9447);
or U9953 (N_9953,N_9492,N_9228);
and U9954 (N_9954,N_9318,N_9127);
nor U9955 (N_9955,N_9079,N_9488);
nor U9956 (N_9956,N_9449,N_9070);
nor U9957 (N_9957,N_9044,N_9154);
or U9958 (N_9958,N_9270,N_9412);
or U9959 (N_9959,N_9118,N_9126);
or U9960 (N_9960,N_9238,N_9343);
nand U9961 (N_9961,N_9478,N_9175);
xor U9962 (N_9962,N_9324,N_9117);
and U9963 (N_9963,N_9436,N_9457);
and U9964 (N_9964,N_9088,N_9226);
or U9965 (N_9965,N_9336,N_9489);
nand U9966 (N_9966,N_9013,N_9061);
nor U9967 (N_9967,N_9110,N_9218);
or U9968 (N_9968,N_9424,N_9263);
xor U9969 (N_9969,N_9065,N_9053);
nor U9970 (N_9970,N_9332,N_9251);
and U9971 (N_9971,N_9444,N_9495);
and U9972 (N_9972,N_9360,N_9358);
nor U9973 (N_9973,N_9257,N_9190);
and U9974 (N_9974,N_9301,N_9373);
nor U9975 (N_9975,N_9023,N_9361);
xnor U9976 (N_9976,N_9120,N_9444);
or U9977 (N_9977,N_9137,N_9169);
and U9978 (N_9978,N_9332,N_9460);
and U9979 (N_9979,N_9295,N_9416);
nor U9980 (N_9980,N_9401,N_9298);
or U9981 (N_9981,N_9427,N_9403);
and U9982 (N_9982,N_9071,N_9042);
xnor U9983 (N_9983,N_9459,N_9221);
nor U9984 (N_9984,N_9477,N_9466);
and U9985 (N_9985,N_9413,N_9177);
and U9986 (N_9986,N_9037,N_9343);
or U9987 (N_9987,N_9146,N_9138);
or U9988 (N_9988,N_9406,N_9103);
nand U9989 (N_9989,N_9218,N_9464);
and U9990 (N_9990,N_9021,N_9162);
or U9991 (N_9991,N_9060,N_9223);
nand U9992 (N_9992,N_9074,N_9364);
or U9993 (N_9993,N_9280,N_9046);
nand U9994 (N_9994,N_9448,N_9339);
or U9995 (N_9995,N_9201,N_9042);
or U9996 (N_9996,N_9190,N_9268);
nand U9997 (N_9997,N_9460,N_9019);
nand U9998 (N_9998,N_9107,N_9401);
or U9999 (N_9999,N_9473,N_9105);
nand UO_0 (O_0,N_9939,N_9765);
and UO_1 (O_1,N_9592,N_9615);
nand UO_2 (O_2,N_9676,N_9910);
xnor UO_3 (O_3,N_9990,N_9512);
nor UO_4 (O_4,N_9651,N_9761);
and UO_5 (O_5,N_9543,N_9997);
and UO_6 (O_6,N_9613,N_9909);
and UO_7 (O_7,N_9976,N_9649);
nor UO_8 (O_8,N_9867,N_9769);
nor UO_9 (O_9,N_9748,N_9754);
xor UO_10 (O_10,N_9724,N_9784);
and UO_11 (O_11,N_9688,N_9915);
and UO_12 (O_12,N_9590,N_9908);
or UO_13 (O_13,N_9515,N_9745);
xor UO_14 (O_14,N_9710,N_9820);
or UO_15 (O_15,N_9921,N_9542);
or UO_16 (O_16,N_9893,N_9587);
nand UO_17 (O_17,N_9575,N_9794);
nand UO_18 (O_18,N_9624,N_9768);
nand UO_19 (O_19,N_9617,N_9559);
or UO_20 (O_20,N_9975,N_9798);
xnor UO_21 (O_21,N_9716,N_9595);
nor UO_22 (O_22,N_9995,N_9660);
nor UO_23 (O_23,N_9989,N_9726);
xor UO_24 (O_24,N_9556,N_9695);
nor UO_25 (O_25,N_9630,N_9770);
or UO_26 (O_26,N_9987,N_9608);
nor UO_27 (O_27,N_9672,N_9747);
nand UO_28 (O_28,N_9718,N_9520);
nand UO_29 (O_29,N_9534,N_9802);
or UO_30 (O_30,N_9550,N_9925);
or UO_31 (O_31,N_9952,N_9558);
nand UO_32 (O_32,N_9571,N_9873);
or UO_33 (O_33,N_9993,N_9998);
nor UO_34 (O_34,N_9898,N_9551);
and UO_35 (O_35,N_9848,N_9854);
nand UO_36 (O_36,N_9846,N_9874);
nand UO_37 (O_37,N_9766,N_9823);
or UO_38 (O_38,N_9830,N_9657);
or UO_39 (O_39,N_9585,N_9962);
nor UO_40 (O_40,N_9896,N_9771);
and UO_41 (O_41,N_9954,N_9831);
nor UO_42 (O_42,N_9859,N_9659);
nand UO_43 (O_43,N_9546,N_9806);
or UO_44 (O_44,N_9828,N_9713);
nor UO_45 (O_45,N_9918,N_9774);
nand UO_46 (O_46,N_9632,N_9978);
nand UO_47 (O_47,N_9776,N_9679);
or UO_48 (O_48,N_9833,N_9689);
nand UO_49 (O_49,N_9963,N_9904);
nor UO_50 (O_50,N_9922,N_9788);
nand UO_51 (O_51,N_9715,N_9879);
and UO_52 (O_52,N_9865,N_9742);
nand UO_53 (O_53,N_9808,N_9662);
and UO_54 (O_54,N_9641,N_9647);
and UO_55 (O_55,N_9717,N_9753);
or UO_56 (O_56,N_9725,N_9580);
xnor UO_57 (O_57,N_9616,N_9604);
and UO_58 (O_58,N_9965,N_9905);
and UO_59 (O_59,N_9889,N_9562);
or UO_60 (O_60,N_9834,N_9863);
nor UO_61 (O_61,N_9596,N_9755);
and UO_62 (O_62,N_9654,N_9957);
and UO_63 (O_63,N_9611,N_9787);
nand UO_64 (O_64,N_9886,N_9914);
nor UO_65 (O_65,N_9735,N_9936);
or UO_66 (O_66,N_9884,N_9927);
xnor UO_67 (O_67,N_9933,N_9700);
nor UO_68 (O_68,N_9693,N_9540);
and UO_69 (O_69,N_9871,N_9665);
and UO_70 (O_70,N_9593,N_9500);
or UO_71 (O_71,N_9658,N_9955);
and UO_72 (O_72,N_9907,N_9972);
and UO_73 (O_73,N_9699,N_9775);
nand UO_74 (O_74,N_9967,N_9866);
or UO_75 (O_75,N_9762,N_9720);
or UO_76 (O_76,N_9574,N_9644);
nand UO_77 (O_77,N_9796,N_9738);
nor UO_78 (O_78,N_9875,N_9988);
nor UO_79 (O_79,N_9639,N_9569);
and UO_80 (O_80,N_9882,N_9721);
nand UO_81 (O_81,N_9712,N_9844);
nor UO_82 (O_82,N_9505,N_9818);
nor UO_83 (O_83,N_9671,N_9812);
nand UO_84 (O_84,N_9779,N_9638);
or UO_85 (O_85,N_9504,N_9750);
nor UO_86 (O_86,N_9937,N_9953);
xor UO_87 (O_87,N_9736,N_9810);
xnor UO_88 (O_88,N_9573,N_9842);
or UO_89 (O_89,N_9881,N_9814);
xor UO_90 (O_90,N_9714,N_9877);
nand UO_91 (O_91,N_9917,N_9803);
and UO_92 (O_92,N_9829,N_9723);
or UO_93 (O_93,N_9981,N_9843);
nor UO_94 (O_94,N_9730,N_9897);
nor UO_95 (O_95,N_9951,N_9675);
and UO_96 (O_96,N_9883,N_9570);
and UO_97 (O_97,N_9661,N_9502);
or UO_98 (O_98,N_9885,N_9870);
or UO_99 (O_99,N_9986,N_9618);
nor UO_100 (O_100,N_9652,N_9579);
nand UO_101 (O_101,N_9743,N_9532);
nand UO_102 (O_102,N_9789,N_9912);
or UO_103 (O_103,N_9599,N_9940);
and UO_104 (O_104,N_9824,N_9746);
and UO_105 (O_105,N_9992,N_9956);
nand UO_106 (O_106,N_9816,N_9529);
or UO_107 (O_107,N_9602,N_9553);
nand UO_108 (O_108,N_9821,N_9627);
nand UO_109 (O_109,N_9522,N_9985);
and UO_110 (O_110,N_9944,N_9872);
or UO_111 (O_111,N_9648,N_9880);
and UO_112 (O_112,N_9841,N_9878);
or UO_113 (O_113,N_9681,N_9759);
and UO_114 (O_114,N_9612,N_9966);
and UO_115 (O_115,N_9778,N_9623);
nand UO_116 (O_116,N_9800,N_9733);
nor UO_117 (O_117,N_9786,N_9669);
and UO_118 (O_118,N_9568,N_9892);
nand UO_119 (O_119,N_9541,N_9506);
xnor UO_120 (O_120,N_9516,N_9847);
and UO_121 (O_121,N_9763,N_9603);
or UO_122 (O_122,N_9835,N_9974);
nor UO_123 (O_123,N_9977,N_9605);
or UO_124 (O_124,N_9792,N_9582);
nor UO_125 (O_125,N_9911,N_9837);
and UO_126 (O_126,N_9622,N_9801);
and UO_127 (O_127,N_9737,N_9561);
xor UO_128 (O_128,N_9584,N_9567);
nor UO_129 (O_129,N_9697,N_9822);
nor UO_130 (O_130,N_9752,N_9729);
or UO_131 (O_131,N_9996,N_9677);
nor UO_132 (O_132,N_9509,N_9513);
nor UO_133 (O_133,N_9811,N_9862);
xnor UO_134 (O_134,N_9864,N_9591);
xnor UO_135 (O_135,N_9781,N_9524);
nor UO_136 (O_136,N_9619,N_9838);
and UO_137 (O_137,N_9626,N_9948);
and UO_138 (O_138,N_9704,N_9935);
nor UO_139 (O_139,N_9678,N_9899);
nand UO_140 (O_140,N_9851,N_9970);
nand UO_141 (O_141,N_9514,N_9674);
and UO_142 (O_142,N_9682,N_9598);
and UO_143 (O_143,N_9741,N_9663);
and UO_144 (O_144,N_9533,N_9791);
and UO_145 (O_145,N_9817,N_9857);
and UO_146 (O_146,N_9519,N_9760);
nand UO_147 (O_147,N_9827,N_9924);
nor UO_148 (O_148,N_9727,N_9926);
and UO_149 (O_149,N_9629,N_9780);
and UO_150 (O_150,N_9653,N_9511);
nor UO_151 (O_151,N_9959,N_9890);
nor UO_152 (O_152,N_9508,N_9691);
nor UO_153 (O_153,N_9999,N_9849);
xnor UO_154 (O_154,N_9578,N_9526);
nand UO_155 (O_155,N_9566,N_9538);
or UO_156 (O_156,N_9709,N_9795);
or UO_157 (O_157,N_9528,N_9941);
or UO_158 (O_158,N_9903,N_9902);
and UO_159 (O_159,N_9635,N_9523);
xnor UO_160 (O_160,N_9544,N_9757);
nand UO_161 (O_161,N_9839,N_9895);
xnor UO_162 (O_162,N_9606,N_9968);
nand UO_163 (O_163,N_9906,N_9620);
nand UO_164 (O_164,N_9913,N_9625);
nor UO_165 (O_165,N_9518,N_9637);
nand UO_166 (O_166,N_9852,N_9557);
nor UO_167 (O_167,N_9785,N_9900);
and UO_168 (O_168,N_9517,N_9836);
nand UO_169 (O_169,N_9692,N_9655);
and UO_170 (O_170,N_9832,N_9583);
nand UO_171 (O_171,N_9799,N_9797);
and UO_172 (O_172,N_9938,N_9530);
nand UO_173 (O_173,N_9636,N_9813);
nand UO_174 (O_174,N_9577,N_9614);
or UO_175 (O_175,N_9706,N_9764);
nand UO_176 (O_176,N_9740,N_9767);
nor UO_177 (O_177,N_9525,N_9973);
and UO_178 (O_178,N_9868,N_9855);
nor UO_179 (O_179,N_9645,N_9640);
and UO_180 (O_180,N_9804,N_9609);
nor UO_181 (O_181,N_9531,N_9698);
and UO_182 (O_182,N_9929,N_9731);
nor UO_183 (O_183,N_9634,N_9790);
nand UO_184 (O_184,N_9961,N_9673);
and UO_185 (O_185,N_9930,N_9739);
nor UO_186 (O_186,N_9979,N_9923);
nand UO_187 (O_187,N_9610,N_9749);
and UO_188 (O_188,N_9949,N_9744);
xor UO_189 (O_189,N_9950,N_9670);
nand UO_190 (O_190,N_9958,N_9946);
or UO_191 (O_191,N_9964,N_9631);
nand UO_192 (O_192,N_9643,N_9667);
nor UO_193 (O_193,N_9728,N_9861);
and UO_194 (O_194,N_9586,N_9825);
or UO_195 (O_195,N_9850,N_9711);
xor UO_196 (O_196,N_9758,N_9805);
nand UO_197 (O_197,N_9971,N_9680);
or UO_198 (O_198,N_9945,N_9607);
and UO_199 (O_199,N_9826,N_9919);
or UO_200 (O_200,N_9537,N_9600);
nand UO_201 (O_201,N_9685,N_9708);
or UO_202 (O_202,N_9980,N_9983);
nand UO_203 (O_203,N_9621,N_9510);
and UO_204 (O_204,N_9777,N_9809);
nor UO_205 (O_205,N_9793,N_9666);
nor UO_206 (O_206,N_9894,N_9901);
or UO_207 (O_207,N_9701,N_9782);
nand UO_208 (O_208,N_9860,N_9840);
nand UO_209 (O_209,N_9783,N_9932);
nand UO_210 (O_210,N_9994,N_9560);
nand UO_211 (O_211,N_9597,N_9686);
nor UO_212 (O_212,N_9819,N_9734);
nor UO_213 (O_213,N_9547,N_9934);
nor UO_214 (O_214,N_9960,N_9694);
xor UO_215 (O_215,N_9845,N_9539);
xnor UO_216 (O_216,N_9548,N_9703);
and UO_217 (O_217,N_9521,N_9722);
nand UO_218 (O_218,N_9555,N_9507);
nand UO_219 (O_219,N_9888,N_9991);
and UO_220 (O_220,N_9656,N_9719);
and UO_221 (O_221,N_9581,N_9690);
nor UO_222 (O_222,N_9984,N_9869);
or UO_223 (O_223,N_9527,N_9942);
nand UO_224 (O_224,N_9588,N_9552);
and UO_225 (O_225,N_9549,N_9687);
and UO_226 (O_226,N_9650,N_9982);
nand UO_227 (O_227,N_9943,N_9684);
nand UO_228 (O_228,N_9576,N_9732);
nor UO_229 (O_229,N_9642,N_9535);
nor UO_230 (O_230,N_9887,N_9920);
nand UO_231 (O_231,N_9858,N_9969);
and UO_232 (O_232,N_9589,N_9702);
nand UO_233 (O_233,N_9947,N_9628);
and UO_234 (O_234,N_9565,N_9696);
nand UO_235 (O_235,N_9773,N_9668);
nand UO_236 (O_236,N_9928,N_9683);
nand UO_237 (O_237,N_9633,N_9772);
nand UO_238 (O_238,N_9756,N_9807);
and UO_239 (O_239,N_9891,N_9601);
or UO_240 (O_240,N_9563,N_9536);
or UO_241 (O_241,N_9707,N_9705);
and UO_242 (O_242,N_9916,N_9931);
xor UO_243 (O_243,N_9856,N_9853);
nor UO_244 (O_244,N_9876,N_9545);
nor UO_245 (O_245,N_9572,N_9664);
nand UO_246 (O_246,N_9594,N_9815);
nand UO_247 (O_247,N_9554,N_9564);
nor UO_248 (O_248,N_9501,N_9751);
xor UO_249 (O_249,N_9646,N_9503);
and UO_250 (O_250,N_9935,N_9666);
and UO_251 (O_251,N_9607,N_9732);
and UO_252 (O_252,N_9508,N_9886);
or UO_253 (O_253,N_9929,N_9566);
or UO_254 (O_254,N_9875,N_9569);
or UO_255 (O_255,N_9807,N_9872);
or UO_256 (O_256,N_9963,N_9655);
or UO_257 (O_257,N_9573,N_9681);
or UO_258 (O_258,N_9992,N_9832);
and UO_259 (O_259,N_9827,N_9757);
nor UO_260 (O_260,N_9723,N_9624);
nor UO_261 (O_261,N_9964,N_9585);
nor UO_262 (O_262,N_9548,N_9872);
or UO_263 (O_263,N_9973,N_9728);
or UO_264 (O_264,N_9940,N_9901);
or UO_265 (O_265,N_9981,N_9564);
nor UO_266 (O_266,N_9875,N_9876);
xor UO_267 (O_267,N_9708,N_9619);
and UO_268 (O_268,N_9776,N_9658);
or UO_269 (O_269,N_9746,N_9992);
xnor UO_270 (O_270,N_9811,N_9679);
nand UO_271 (O_271,N_9803,N_9938);
or UO_272 (O_272,N_9658,N_9952);
and UO_273 (O_273,N_9865,N_9988);
nor UO_274 (O_274,N_9501,N_9597);
or UO_275 (O_275,N_9775,N_9788);
or UO_276 (O_276,N_9601,N_9808);
nand UO_277 (O_277,N_9922,N_9617);
nor UO_278 (O_278,N_9583,N_9997);
nor UO_279 (O_279,N_9689,N_9918);
and UO_280 (O_280,N_9613,N_9534);
nand UO_281 (O_281,N_9884,N_9945);
nor UO_282 (O_282,N_9984,N_9977);
xor UO_283 (O_283,N_9571,N_9943);
and UO_284 (O_284,N_9512,N_9893);
or UO_285 (O_285,N_9900,N_9973);
nor UO_286 (O_286,N_9635,N_9841);
nand UO_287 (O_287,N_9516,N_9508);
nor UO_288 (O_288,N_9557,N_9771);
and UO_289 (O_289,N_9661,N_9962);
nand UO_290 (O_290,N_9871,N_9893);
nand UO_291 (O_291,N_9835,N_9709);
xor UO_292 (O_292,N_9700,N_9975);
nand UO_293 (O_293,N_9904,N_9768);
or UO_294 (O_294,N_9703,N_9638);
or UO_295 (O_295,N_9873,N_9768);
or UO_296 (O_296,N_9618,N_9787);
nand UO_297 (O_297,N_9683,N_9642);
and UO_298 (O_298,N_9983,N_9695);
xor UO_299 (O_299,N_9830,N_9920);
nand UO_300 (O_300,N_9882,N_9992);
and UO_301 (O_301,N_9552,N_9649);
and UO_302 (O_302,N_9980,N_9678);
nor UO_303 (O_303,N_9728,N_9558);
nor UO_304 (O_304,N_9828,N_9683);
nand UO_305 (O_305,N_9920,N_9818);
nand UO_306 (O_306,N_9592,N_9727);
nand UO_307 (O_307,N_9608,N_9696);
xnor UO_308 (O_308,N_9835,N_9641);
or UO_309 (O_309,N_9999,N_9969);
nand UO_310 (O_310,N_9504,N_9719);
and UO_311 (O_311,N_9545,N_9988);
xor UO_312 (O_312,N_9673,N_9715);
and UO_313 (O_313,N_9605,N_9663);
and UO_314 (O_314,N_9550,N_9618);
nor UO_315 (O_315,N_9886,N_9999);
nand UO_316 (O_316,N_9538,N_9617);
and UO_317 (O_317,N_9556,N_9781);
and UO_318 (O_318,N_9851,N_9537);
nand UO_319 (O_319,N_9639,N_9576);
or UO_320 (O_320,N_9929,N_9552);
nand UO_321 (O_321,N_9682,N_9521);
or UO_322 (O_322,N_9843,N_9971);
or UO_323 (O_323,N_9782,N_9814);
nor UO_324 (O_324,N_9672,N_9804);
and UO_325 (O_325,N_9685,N_9619);
xor UO_326 (O_326,N_9644,N_9610);
or UO_327 (O_327,N_9963,N_9891);
xnor UO_328 (O_328,N_9829,N_9923);
and UO_329 (O_329,N_9821,N_9794);
or UO_330 (O_330,N_9916,N_9940);
xnor UO_331 (O_331,N_9582,N_9725);
and UO_332 (O_332,N_9596,N_9844);
or UO_333 (O_333,N_9784,N_9982);
nand UO_334 (O_334,N_9510,N_9500);
or UO_335 (O_335,N_9711,N_9939);
nand UO_336 (O_336,N_9795,N_9816);
and UO_337 (O_337,N_9877,N_9698);
nand UO_338 (O_338,N_9726,N_9694);
or UO_339 (O_339,N_9935,N_9882);
nand UO_340 (O_340,N_9689,N_9928);
xnor UO_341 (O_341,N_9953,N_9805);
nand UO_342 (O_342,N_9623,N_9994);
nand UO_343 (O_343,N_9607,N_9541);
and UO_344 (O_344,N_9513,N_9647);
nor UO_345 (O_345,N_9519,N_9945);
or UO_346 (O_346,N_9590,N_9587);
and UO_347 (O_347,N_9754,N_9951);
and UO_348 (O_348,N_9780,N_9715);
nor UO_349 (O_349,N_9764,N_9647);
and UO_350 (O_350,N_9784,N_9810);
nand UO_351 (O_351,N_9770,N_9884);
and UO_352 (O_352,N_9786,N_9746);
nand UO_353 (O_353,N_9768,N_9572);
and UO_354 (O_354,N_9691,N_9593);
and UO_355 (O_355,N_9783,N_9909);
or UO_356 (O_356,N_9839,N_9960);
or UO_357 (O_357,N_9847,N_9676);
or UO_358 (O_358,N_9637,N_9717);
and UO_359 (O_359,N_9594,N_9994);
xnor UO_360 (O_360,N_9559,N_9902);
xor UO_361 (O_361,N_9522,N_9598);
or UO_362 (O_362,N_9528,N_9976);
or UO_363 (O_363,N_9551,N_9554);
nand UO_364 (O_364,N_9867,N_9831);
nor UO_365 (O_365,N_9635,N_9675);
or UO_366 (O_366,N_9839,N_9816);
and UO_367 (O_367,N_9993,N_9500);
or UO_368 (O_368,N_9662,N_9824);
and UO_369 (O_369,N_9650,N_9611);
nor UO_370 (O_370,N_9770,N_9694);
nor UO_371 (O_371,N_9511,N_9794);
or UO_372 (O_372,N_9803,N_9825);
and UO_373 (O_373,N_9614,N_9674);
nand UO_374 (O_374,N_9530,N_9820);
nand UO_375 (O_375,N_9922,N_9664);
and UO_376 (O_376,N_9803,N_9652);
or UO_377 (O_377,N_9791,N_9503);
nor UO_378 (O_378,N_9932,N_9996);
and UO_379 (O_379,N_9729,N_9634);
or UO_380 (O_380,N_9663,N_9686);
or UO_381 (O_381,N_9738,N_9507);
and UO_382 (O_382,N_9516,N_9506);
and UO_383 (O_383,N_9978,N_9546);
nand UO_384 (O_384,N_9682,N_9743);
or UO_385 (O_385,N_9582,N_9880);
nand UO_386 (O_386,N_9719,N_9871);
nor UO_387 (O_387,N_9553,N_9533);
nand UO_388 (O_388,N_9885,N_9859);
nor UO_389 (O_389,N_9683,N_9655);
nor UO_390 (O_390,N_9547,N_9858);
nand UO_391 (O_391,N_9703,N_9827);
or UO_392 (O_392,N_9581,N_9751);
nor UO_393 (O_393,N_9658,N_9974);
or UO_394 (O_394,N_9624,N_9774);
or UO_395 (O_395,N_9953,N_9985);
and UO_396 (O_396,N_9700,N_9608);
and UO_397 (O_397,N_9510,N_9673);
and UO_398 (O_398,N_9676,N_9514);
nor UO_399 (O_399,N_9859,N_9670);
or UO_400 (O_400,N_9888,N_9747);
nor UO_401 (O_401,N_9692,N_9750);
xnor UO_402 (O_402,N_9871,N_9570);
nor UO_403 (O_403,N_9691,N_9662);
nand UO_404 (O_404,N_9768,N_9555);
nor UO_405 (O_405,N_9610,N_9894);
or UO_406 (O_406,N_9635,N_9543);
xnor UO_407 (O_407,N_9792,N_9674);
and UO_408 (O_408,N_9791,N_9775);
and UO_409 (O_409,N_9511,N_9731);
or UO_410 (O_410,N_9904,N_9657);
and UO_411 (O_411,N_9599,N_9617);
and UO_412 (O_412,N_9858,N_9857);
and UO_413 (O_413,N_9631,N_9773);
nand UO_414 (O_414,N_9632,N_9504);
nor UO_415 (O_415,N_9562,N_9644);
nor UO_416 (O_416,N_9608,N_9633);
or UO_417 (O_417,N_9642,N_9737);
or UO_418 (O_418,N_9647,N_9630);
or UO_419 (O_419,N_9524,N_9643);
nand UO_420 (O_420,N_9770,N_9939);
or UO_421 (O_421,N_9593,N_9912);
nor UO_422 (O_422,N_9509,N_9933);
xor UO_423 (O_423,N_9658,N_9917);
nand UO_424 (O_424,N_9959,N_9811);
nand UO_425 (O_425,N_9983,N_9994);
and UO_426 (O_426,N_9715,N_9506);
and UO_427 (O_427,N_9523,N_9509);
nor UO_428 (O_428,N_9543,N_9506);
and UO_429 (O_429,N_9570,N_9733);
and UO_430 (O_430,N_9712,N_9654);
or UO_431 (O_431,N_9777,N_9571);
or UO_432 (O_432,N_9945,N_9758);
or UO_433 (O_433,N_9918,N_9643);
and UO_434 (O_434,N_9542,N_9958);
nand UO_435 (O_435,N_9819,N_9987);
nor UO_436 (O_436,N_9555,N_9500);
nand UO_437 (O_437,N_9902,N_9925);
and UO_438 (O_438,N_9587,N_9574);
nor UO_439 (O_439,N_9828,N_9741);
xnor UO_440 (O_440,N_9870,N_9625);
and UO_441 (O_441,N_9986,N_9599);
and UO_442 (O_442,N_9864,N_9672);
nand UO_443 (O_443,N_9547,N_9667);
nor UO_444 (O_444,N_9627,N_9630);
or UO_445 (O_445,N_9580,N_9726);
xnor UO_446 (O_446,N_9603,N_9540);
nand UO_447 (O_447,N_9770,N_9627);
nor UO_448 (O_448,N_9963,N_9908);
nand UO_449 (O_449,N_9729,N_9639);
nor UO_450 (O_450,N_9659,N_9903);
and UO_451 (O_451,N_9929,N_9911);
nand UO_452 (O_452,N_9681,N_9623);
xor UO_453 (O_453,N_9706,N_9506);
and UO_454 (O_454,N_9710,N_9559);
and UO_455 (O_455,N_9989,N_9884);
or UO_456 (O_456,N_9640,N_9715);
xnor UO_457 (O_457,N_9877,N_9772);
nor UO_458 (O_458,N_9697,N_9920);
and UO_459 (O_459,N_9717,N_9617);
or UO_460 (O_460,N_9537,N_9690);
xnor UO_461 (O_461,N_9952,N_9716);
and UO_462 (O_462,N_9536,N_9835);
nor UO_463 (O_463,N_9944,N_9519);
or UO_464 (O_464,N_9780,N_9579);
or UO_465 (O_465,N_9861,N_9980);
xnor UO_466 (O_466,N_9915,N_9820);
and UO_467 (O_467,N_9761,N_9733);
nand UO_468 (O_468,N_9547,N_9602);
nand UO_469 (O_469,N_9612,N_9936);
nor UO_470 (O_470,N_9991,N_9885);
and UO_471 (O_471,N_9691,N_9630);
nor UO_472 (O_472,N_9953,N_9956);
nor UO_473 (O_473,N_9968,N_9771);
nor UO_474 (O_474,N_9574,N_9930);
nor UO_475 (O_475,N_9924,N_9669);
nor UO_476 (O_476,N_9651,N_9538);
xor UO_477 (O_477,N_9821,N_9612);
and UO_478 (O_478,N_9879,N_9809);
nand UO_479 (O_479,N_9904,N_9686);
nor UO_480 (O_480,N_9991,N_9702);
and UO_481 (O_481,N_9675,N_9859);
xor UO_482 (O_482,N_9557,N_9816);
or UO_483 (O_483,N_9974,N_9894);
and UO_484 (O_484,N_9986,N_9899);
or UO_485 (O_485,N_9583,N_9783);
nor UO_486 (O_486,N_9623,N_9615);
or UO_487 (O_487,N_9827,N_9603);
or UO_488 (O_488,N_9820,N_9953);
and UO_489 (O_489,N_9912,N_9665);
xor UO_490 (O_490,N_9712,N_9514);
nand UO_491 (O_491,N_9517,N_9732);
and UO_492 (O_492,N_9772,N_9541);
nand UO_493 (O_493,N_9779,N_9629);
and UO_494 (O_494,N_9790,N_9809);
and UO_495 (O_495,N_9911,N_9723);
nor UO_496 (O_496,N_9768,N_9781);
nor UO_497 (O_497,N_9570,N_9930);
nor UO_498 (O_498,N_9587,N_9876);
nand UO_499 (O_499,N_9523,N_9622);
nor UO_500 (O_500,N_9779,N_9758);
or UO_501 (O_501,N_9518,N_9940);
or UO_502 (O_502,N_9747,N_9909);
nor UO_503 (O_503,N_9580,N_9691);
and UO_504 (O_504,N_9712,N_9863);
nand UO_505 (O_505,N_9575,N_9880);
nand UO_506 (O_506,N_9582,N_9920);
nand UO_507 (O_507,N_9825,N_9828);
or UO_508 (O_508,N_9827,N_9717);
and UO_509 (O_509,N_9695,N_9840);
nand UO_510 (O_510,N_9993,N_9661);
or UO_511 (O_511,N_9644,N_9998);
and UO_512 (O_512,N_9697,N_9602);
nand UO_513 (O_513,N_9741,N_9730);
or UO_514 (O_514,N_9858,N_9863);
and UO_515 (O_515,N_9978,N_9838);
xor UO_516 (O_516,N_9767,N_9792);
xor UO_517 (O_517,N_9621,N_9727);
xnor UO_518 (O_518,N_9975,N_9569);
nand UO_519 (O_519,N_9679,N_9503);
and UO_520 (O_520,N_9509,N_9864);
nand UO_521 (O_521,N_9651,N_9855);
xnor UO_522 (O_522,N_9946,N_9898);
and UO_523 (O_523,N_9870,N_9536);
xnor UO_524 (O_524,N_9589,N_9898);
nor UO_525 (O_525,N_9987,N_9733);
nor UO_526 (O_526,N_9665,N_9853);
nand UO_527 (O_527,N_9595,N_9664);
nand UO_528 (O_528,N_9700,N_9815);
and UO_529 (O_529,N_9569,N_9623);
nor UO_530 (O_530,N_9694,N_9559);
nand UO_531 (O_531,N_9876,N_9509);
nor UO_532 (O_532,N_9747,N_9858);
and UO_533 (O_533,N_9838,N_9580);
nand UO_534 (O_534,N_9809,N_9768);
and UO_535 (O_535,N_9595,N_9890);
nand UO_536 (O_536,N_9951,N_9501);
nor UO_537 (O_537,N_9760,N_9666);
or UO_538 (O_538,N_9911,N_9545);
or UO_539 (O_539,N_9518,N_9576);
and UO_540 (O_540,N_9942,N_9532);
and UO_541 (O_541,N_9665,N_9586);
nor UO_542 (O_542,N_9541,N_9633);
or UO_543 (O_543,N_9535,N_9828);
or UO_544 (O_544,N_9750,N_9712);
or UO_545 (O_545,N_9536,N_9565);
nand UO_546 (O_546,N_9549,N_9883);
nand UO_547 (O_547,N_9673,N_9545);
and UO_548 (O_548,N_9720,N_9605);
and UO_549 (O_549,N_9617,N_9603);
nor UO_550 (O_550,N_9694,N_9741);
nand UO_551 (O_551,N_9726,N_9759);
nor UO_552 (O_552,N_9709,N_9759);
nor UO_553 (O_553,N_9848,N_9832);
and UO_554 (O_554,N_9764,N_9776);
or UO_555 (O_555,N_9847,N_9954);
nand UO_556 (O_556,N_9867,N_9636);
nor UO_557 (O_557,N_9842,N_9663);
xnor UO_558 (O_558,N_9814,N_9530);
xnor UO_559 (O_559,N_9807,N_9781);
or UO_560 (O_560,N_9831,N_9958);
nand UO_561 (O_561,N_9631,N_9833);
nor UO_562 (O_562,N_9919,N_9715);
and UO_563 (O_563,N_9873,N_9877);
nor UO_564 (O_564,N_9805,N_9550);
xor UO_565 (O_565,N_9719,N_9766);
and UO_566 (O_566,N_9798,N_9690);
xor UO_567 (O_567,N_9816,N_9619);
nor UO_568 (O_568,N_9771,N_9589);
nand UO_569 (O_569,N_9933,N_9869);
and UO_570 (O_570,N_9622,N_9570);
and UO_571 (O_571,N_9920,N_9895);
xnor UO_572 (O_572,N_9620,N_9655);
or UO_573 (O_573,N_9709,N_9700);
nor UO_574 (O_574,N_9850,N_9593);
or UO_575 (O_575,N_9568,N_9902);
nand UO_576 (O_576,N_9557,N_9616);
and UO_577 (O_577,N_9962,N_9855);
nor UO_578 (O_578,N_9901,N_9903);
and UO_579 (O_579,N_9926,N_9734);
xnor UO_580 (O_580,N_9965,N_9861);
nor UO_581 (O_581,N_9518,N_9505);
nor UO_582 (O_582,N_9992,N_9522);
nand UO_583 (O_583,N_9959,N_9734);
nand UO_584 (O_584,N_9513,N_9831);
or UO_585 (O_585,N_9519,N_9721);
nand UO_586 (O_586,N_9785,N_9866);
and UO_587 (O_587,N_9733,N_9992);
or UO_588 (O_588,N_9910,N_9793);
nor UO_589 (O_589,N_9773,N_9759);
nand UO_590 (O_590,N_9750,N_9847);
or UO_591 (O_591,N_9691,N_9640);
nand UO_592 (O_592,N_9503,N_9713);
nor UO_593 (O_593,N_9706,N_9587);
xnor UO_594 (O_594,N_9581,N_9551);
nand UO_595 (O_595,N_9936,N_9619);
xor UO_596 (O_596,N_9614,N_9855);
nor UO_597 (O_597,N_9940,N_9853);
or UO_598 (O_598,N_9680,N_9675);
xnor UO_599 (O_599,N_9535,N_9770);
or UO_600 (O_600,N_9632,N_9690);
and UO_601 (O_601,N_9733,N_9546);
nor UO_602 (O_602,N_9615,N_9827);
or UO_603 (O_603,N_9900,N_9764);
nand UO_604 (O_604,N_9502,N_9633);
or UO_605 (O_605,N_9995,N_9605);
and UO_606 (O_606,N_9528,N_9718);
or UO_607 (O_607,N_9726,N_9627);
or UO_608 (O_608,N_9717,N_9636);
nor UO_609 (O_609,N_9554,N_9530);
nor UO_610 (O_610,N_9948,N_9517);
xnor UO_611 (O_611,N_9838,N_9592);
nor UO_612 (O_612,N_9566,N_9577);
or UO_613 (O_613,N_9683,N_9882);
nor UO_614 (O_614,N_9568,N_9924);
and UO_615 (O_615,N_9886,N_9970);
and UO_616 (O_616,N_9895,N_9696);
xnor UO_617 (O_617,N_9914,N_9500);
nand UO_618 (O_618,N_9892,N_9830);
and UO_619 (O_619,N_9807,N_9682);
nor UO_620 (O_620,N_9911,N_9868);
and UO_621 (O_621,N_9818,N_9598);
and UO_622 (O_622,N_9873,N_9813);
nor UO_623 (O_623,N_9858,N_9727);
nand UO_624 (O_624,N_9820,N_9595);
nand UO_625 (O_625,N_9538,N_9976);
nand UO_626 (O_626,N_9733,N_9684);
and UO_627 (O_627,N_9976,N_9733);
nor UO_628 (O_628,N_9817,N_9810);
and UO_629 (O_629,N_9586,N_9961);
or UO_630 (O_630,N_9833,N_9690);
or UO_631 (O_631,N_9694,N_9840);
or UO_632 (O_632,N_9730,N_9783);
nor UO_633 (O_633,N_9860,N_9815);
nor UO_634 (O_634,N_9997,N_9914);
nand UO_635 (O_635,N_9500,N_9930);
and UO_636 (O_636,N_9608,N_9814);
and UO_637 (O_637,N_9525,N_9689);
xnor UO_638 (O_638,N_9542,N_9649);
and UO_639 (O_639,N_9813,N_9998);
and UO_640 (O_640,N_9823,N_9893);
nor UO_641 (O_641,N_9538,N_9756);
nor UO_642 (O_642,N_9830,N_9532);
nor UO_643 (O_643,N_9844,N_9941);
or UO_644 (O_644,N_9800,N_9929);
and UO_645 (O_645,N_9926,N_9649);
and UO_646 (O_646,N_9993,N_9829);
or UO_647 (O_647,N_9808,N_9528);
nor UO_648 (O_648,N_9512,N_9667);
nor UO_649 (O_649,N_9801,N_9850);
and UO_650 (O_650,N_9969,N_9963);
nand UO_651 (O_651,N_9538,N_9985);
nor UO_652 (O_652,N_9576,N_9550);
and UO_653 (O_653,N_9662,N_9757);
nand UO_654 (O_654,N_9597,N_9968);
nand UO_655 (O_655,N_9786,N_9784);
nor UO_656 (O_656,N_9556,N_9521);
xor UO_657 (O_657,N_9643,N_9798);
nand UO_658 (O_658,N_9983,N_9882);
nor UO_659 (O_659,N_9991,N_9584);
or UO_660 (O_660,N_9532,N_9990);
and UO_661 (O_661,N_9714,N_9999);
nand UO_662 (O_662,N_9791,N_9909);
xor UO_663 (O_663,N_9820,N_9923);
or UO_664 (O_664,N_9678,N_9646);
nor UO_665 (O_665,N_9718,N_9944);
or UO_666 (O_666,N_9970,N_9668);
or UO_667 (O_667,N_9945,N_9968);
nor UO_668 (O_668,N_9513,N_9657);
nor UO_669 (O_669,N_9783,N_9985);
xor UO_670 (O_670,N_9794,N_9504);
or UO_671 (O_671,N_9545,N_9938);
nor UO_672 (O_672,N_9851,N_9740);
nor UO_673 (O_673,N_9949,N_9650);
or UO_674 (O_674,N_9585,N_9909);
nand UO_675 (O_675,N_9504,N_9723);
xor UO_676 (O_676,N_9782,N_9806);
or UO_677 (O_677,N_9542,N_9987);
nand UO_678 (O_678,N_9854,N_9903);
xor UO_679 (O_679,N_9636,N_9629);
or UO_680 (O_680,N_9895,N_9851);
or UO_681 (O_681,N_9978,N_9513);
nor UO_682 (O_682,N_9843,N_9544);
and UO_683 (O_683,N_9891,N_9616);
nor UO_684 (O_684,N_9775,N_9539);
xor UO_685 (O_685,N_9864,N_9553);
nand UO_686 (O_686,N_9729,N_9632);
or UO_687 (O_687,N_9835,N_9983);
or UO_688 (O_688,N_9658,N_9622);
nand UO_689 (O_689,N_9759,N_9853);
nand UO_690 (O_690,N_9537,N_9705);
or UO_691 (O_691,N_9549,N_9931);
or UO_692 (O_692,N_9837,N_9729);
and UO_693 (O_693,N_9599,N_9884);
nand UO_694 (O_694,N_9552,N_9544);
xnor UO_695 (O_695,N_9716,N_9732);
and UO_696 (O_696,N_9525,N_9849);
or UO_697 (O_697,N_9586,N_9535);
nor UO_698 (O_698,N_9629,N_9877);
xnor UO_699 (O_699,N_9757,N_9946);
nand UO_700 (O_700,N_9635,N_9940);
nand UO_701 (O_701,N_9645,N_9677);
xnor UO_702 (O_702,N_9524,N_9597);
nand UO_703 (O_703,N_9639,N_9724);
nor UO_704 (O_704,N_9518,N_9908);
and UO_705 (O_705,N_9590,N_9515);
nand UO_706 (O_706,N_9909,N_9891);
or UO_707 (O_707,N_9849,N_9965);
nor UO_708 (O_708,N_9792,N_9645);
and UO_709 (O_709,N_9628,N_9908);
nor UO_710 (O_710,N_9511,N_9728);
and UO_711 (O_711,N_9509,N_9718);
or UO_712 (O_712,N_9841,N_9982);
or UO_713 (O_713,N_9747,N_9710);
or UO_714 (O_714,N_9770,N_9945);
xor UO_715 (O_715,N_9815,N_9583);
xor UO_716 (O_716,N_9944,N_9839);
nor UO_717 (O_717,N_9737,N_9505);
xor UO_718 (O_718,N_9769,N_9958);
nor UO_719 (O_719,N_9538,N_9890);
nand UO_720 (O_720,N_9960,N_9517);
and UO_721 (O_721,N_9694,N_9670);
nand UO_722 (O_722,N_9596,N_9687);
and UO_723 (O_723,N_9697,N_9812);
nor UO_724 (O_724,N_9765,N_9872);
or UO_725 (O_725,N_9572,N_9702);
nand UO_726 (O_726,N_9680,N_9545);
or UO_727 (O_727,N_9747,N_9925);
nand UO_728 (O_728,N_9656,N_9710);
nand UO_729 (O_729,N_9501,N_9572);
xnor UO_730 (O_730,N_9606,N_9934);
xor UO_731 (O_731,N_9541,N_9560);
and UO_732 (O_732,N_9505,N_9638);
and UO_733 (O_733,N_9548,N_9751);
nand UO_734 (O_734,N_9757,N_9665);
and UO_735 (O_735,N_9630,N_9806);
xor UO_736 (O_736,N_9576,N_9594);
xor UO_737 (O_737,N_9867,N_9574);
xnor UO_738 (O_738,N_9539,N_9790);
and UO_739 (O_739,N_9945,N_9694);
nand UO_740 (O_740,N_9765,N_9885);
or UO_741 (O_741,N_9594,N_9622);
xor UO_742 (O_742,N_9993,N_9530);
nand UO_743 (O_743,N_9611,N_9744);
nor UO_744 (O_744,N_9599,N_9892);
nand UO_745 (O_745,N_9722,N_9552);
or UO_746 (O_746,N_9920,N_9593);
or UO_747 (O_747,N_9526,N_9606);
or UO_748 (O_748,N_9586,N_9872);
or UO_749 (O_749,N_9806,N_9765);
and UO_750 (O_750,N_9799,N_9629);
xor UO_751 (O_751,N_9759,N_9863);
or UO_752 (O_752,N_9555,N_9833);
and UO_753 (O_753,N_9793,N_9587);
or UO_754 (O_754,N_9866,N_9836);
and UO_755 (O_755,N_9941,N_9753);
nor UO_756 (O_756,N_9638,N_9961);
or UO_757 (O_757,N_9754,N_9812);
xor UO_758 (O_758,N_9712,N_9885);
and UO_759 (O_759,N_9627,N_9857);
nand UO_760 (O_760,N_9654,N_9814);
xor UO_761 (O_761,N_9987,N_9890);
or UO_762 (O_762,N_9601,N_9885);
and UO_763 (O_763,N_9732,N_9896);
nand UO_764 (O_764,N_9989,N_9990);
and UO_765 (O_765,N_9565,N_9852);
nand UO_766 (O_766,N_9741,N_9923);
nor UO_767 (O_767,N_9735,N_9901);
xor UO_768 (O_768,N_9920,N_9741);
xnor UO_769 (O_769,N_9838,N_9776);
and UO_770 (O_770,N_9760,N_9586);
or UO_771 (O_771,N_9542,N_9780);
nor UO_772 (O_772,N_9999,N_9564);
and UO_773 (O_773,N_9823,N_9905);
and UO_774 (O_774,N_9869,N_9809);
and UO_775 (O_775,N_9833,N_9977);
or UO_776 (O_776,N_9764,N_9566);
or UO_777 (O_777,N_9937,N_9554);
and UO_778 (O_778,N_9818,N_9988);
nor UO_779 (O_779,N_9722,N_9996);
and UO_780 (O_780,N_9610,N_9666);
xnor UO_781 (O_781,N_9519,N_9867);
or UO_782 (O_782,N_9874,N_9951);
nor UO_783 (O_783,N_9815,N_9942);
and UO_784 (O_784,N_9728,N_9718);
or UO_785 (O_785,N_9769,N_9823);
and UO_786 (O_786,N_9665,N_9518);
nand UO_787 (O_787,N_9898,N_9668);
xor UO_788 (O_788,N_9771,N_9671);
xnor UO_789 (O_789,N_9631,N_9930);
xor UO_790 (O_790,N_9824,N_9603);
or UO_791 (O_791,N_9959,N_9640);
nor UO_792 (O_792,N_9827,N_9598);
and UO_793 (O_793,N_9943,N_9660);
or UO_794 (O_794,N_9745,N_9778);
nand UO_795 (O_795,N_9633,N_9524);
and UO_796 (O_796,N_9971,N_9654);
nor UO_797 (O_797,N_9766,N_9642);
xor UO_798 (O_798,N_9591,N_9986);
nor UO_799 (O_799,N_9539,N_9731);
nand UO_800 (O_800,N_9646,N_9554);
nor UO_801 (O_801,N_9657,N_9891);
and UO_802 (O_802,N_9949,N_9766);
nand UO_803 (O_803,N_9709,N_9935);
nor UO_804 (O_804,N_9796,N_9860);
and UO_805 (O_805,N_9723,N_9872);
nor UO_806 (O_806,N_9628,N_9790);
xor UO_807 (O_807,N_9809,N_9887);
nand UO_808 (O_808,N_9848,N_9827);
or UO_809 (O_809,N_9956,N_9559);
nand UO_810 (O_810,N_9706,N_9994);
and UO_811 (O_811,N_9897,N_9656);
or UO_812 (O_812,N_9611,N_9564);
or UO_813 (O_813,N_9768,N_9639);
or UO_814 (O_814,N_9736,N_9852);
or UO_815 (O_815,N_9742,N_9838);
nand UO_816 (O_816,N_9714,N_9786);
and UO_817 (O_817,N_9851,N_9852);
nor UO_818 (O_818,N_9625,N_9689);
or UO_819 (O_819,N_9629,N_9601);
nand UO_820 (O_820,N_9763,N_9777);
or UO_821 (O_821,N_9616,N_9825);
and UO_822 (O_822,N_9739,N_9563);
nor UO_823 (O_823,N_9850,N_9699);
nand UO_824 (O_824,N_9520,N_9659);
nor UO_825 (O_825,N_9692,N_9715);
or UO_826 (O_826,N_9756,N_9912);
nor UO_827 (O_827,N_9739,N_9541);
and UO_828 (O_828,N_9515,N_9903);
or UO_829 (O_829,N_9748,N_9535);
and UO_830 (O_830,N_9533,N_9988);
or UO_831 (O_831,N_9986,N_9702);
or UO_832 (O_832,N_9690,N_9735);
xnor UO_833 (O_833,N_9848,N_9907);
nand UO_834 (O_834,N_9830,N_9720);
nand UO_835 (O_835,N_9649,N_9503);
or UO_836 (O_836,N_9539,N_9972);
and UO_837 (O_837,N_9912,N_9773);
nor UO_838 (O_838,N_9730,N_9848);
nor UO_839 (O_839,N_9731,N_9823);
nand UO_840 (O_840,N_9757,N_9858);
xnor UO_841 (O_841,N_9824,N_9535);
nor UO_842 (O_842,N_9813,N_9732);
and UO_843 (O_843,N_9627,N_9564);
nand UO_844 (O_844,N_9715,N_9894);
or UO_845 (O_845,N_9539,N_9807);
nor UO_846 (O_846,N_9717,N_9595);
xnor UO_847 (O_847,N_9940,N_9784);
or UO_848 (O_848,N_9796,N_9789);
nor UO_849 (O_849,N_9887,N_9821);
nor UO_850 (O_850,N_9898,N_9753);
or UO_851 (O_851,N_9634,N_9724);
or UO_852 (O_852,N_9631,N_9648);
nand UO_853 (O_853,N_9988,N_9652);
xor UO_854 (O_854,N_9951,N_9563);
nand UO_855 (O_855,N_9813,N_9761);
nor UO_856 (O_856,N_9602,N_9755);
nor UO_857 (O_857,N_9726,N_9767);
and UO_858 (O_858,N_9940,N_9566);
nor UO_859 (O_859,N_9924,N_9533);
or UO_860 (O_860,N_9632,N_9839);
nand UO_861 (O_861,N_9891,N_9716);
or UO_862 (O_862,N_9791,N_9959);
xnor UO_863 (O_863,N_9703,N_9893);
nand UO_864 (O_864,N_9643,N_9565);
nand UO_865 (O_865,N_9763,N_9563);
nor UO_866 (O_866,N_9627,N_9636);
nand UO_867 (O_867,N_9746,N_9842);
nor UO_868 (O_868,N_9757,N_9500);
and UO_869 (O_869,N_9937,N_9875);
xor UO_870 (O_870,N_9820,N_9709);
nor UO_871 (O_871,N_9559,N_9998);
and UO_872 (O_872,N_9973,N_9720);
or UO_873 (O_873,N_9787,N_9525);
or UO_874 (O_874,N_9588,N_9879);
nand UO_875 (O_875,N_9740,N_9952);
nand UO_876 (O_876,N_9502,N_9874);
and UO_877 (O_877,N_9618,N_9624);
xor UO_878 (O_878,N_9851,N_9741);
nor UO_879 (O_879,N_9769,N_9657);
and UO_880 (O_880,N_9645,N_9876);
or UO_881 (O_881,N_9676,N_9667);
nor UO_882 (O_882,N_9838,N_9681);
nand UO_883 (O_883,N_9891,N_9761);
or UO_884 (O_884,N_9724,N_9803);
nor UO_885 (O_885,N_9910,N_9508);
or UO_886 (O_886,N_9556,N_9826);
xnor UO_887 (O_887,N_9817,N_9885);
or UO_888 (O_888,N_9762,N_9690);
nand UO_889 (O_889,N_9702,N_9834);
and UO_890 (O_890,N_9589,N_9763);
and UO_891 (O_891,N_9701,N_9853);
or UO_892 (O_892,N_9941,N_9733);
nor UO_893 (O_893,N_9841,N_9591);
and UO_894 (O_894,N_9839,N_9636);
and UO_895 (O_895,N_9763,N_9915);
xnor UO_896 (O_896,N_9659,N_9537);
or UO_897 (O_897,N_9505,N_9573);
and UO_898 (O_898,N_9769,N_9837);
nor UO_899 (O_899,N_9647,N_9650);
nand UO_900 (O_900,N_9972,N_9546);
nand UO_901 (O_901,N_9871,N_9649);
and UO_902 (O_902,N_9552,N_9684);
and UO_903 (O_903,N_9646,N_9717);
or UO_904 (O_904,N_9902,N_9964);
nand UO_905 (O_905,N_9730,N_9692);
and UO_906 (O_906,N_9604,N_9971);
and UO_907 (O_907,N_9643,N_9910);
nor UO_908 (O_908,N_9644,N_9758);
xor UO_909 (O_909,N_9853,N_9901);
xnor UO_910 (O_910,N_9655,N_9585);
nor UO_911 (O_911,N_9738,N_9915);
or UO_912 (O_912,N_9882,N_9937);
or UO_913 (O_913,N_9758,N_9835);
or UO_914 (O_914,N_9502,N_9891);
nand UO_915 (O_915,N_9895,N_9554);
or UO_916 (O_916,N_9709,N_9567);
nand UO_917 (O_917,N_9971,N_9586);
and UO_918 (O_918,N_9778,N_9503);
or UO_919 (O_919,N_9885,N_9722);
nor UO_920 (O_920,N_9575,N_9505);
xnor UO_921 (O_921,N_9930,N_9513);
or UO_922 (O_922,N_9811,N_9830);
nor UO_923 (O_923,N_9973,N_9520);
and UO_924 (O_924,N_9881,N_9869);
nand UO_925 (O_925,N_9562,N_9923);
nand UO_926 (O_926,N_9770,N_9528);
and UO_927 (O_927,N_9766,N_9742);
nor UO_928 (O_928,N_9910,N_9865);
nand UO_929 (O_929,N_9986,N_9979);
or UO_930 (O_930,N_9818,N_9660);
nor UO_931 (O_931,N_9928,N_9917);
xor UO_932 (O_932,N_9522,N_9955);
nand UO_933 (O_933,N_9611,N_9873);
xnor UO_934 (O_934,N_9879,N_9839);
and UO_935 (O_935,N_9567,N_9693);
xor UO_936 (O_936,N_9834,N_9594);
nand UO_937 (O_937,N_9553,N_9710);
nor UO_938 (O_938,N_9575,N_9720);
nor UO_939 (O_939,N_9537,N_9785);
nand UO_940 (O_940,N_9976,N_9591);
nor UO_941 (O_941,N_9587,N_9681);
or UO_942 (O_942,N_9669,N_9836);
nand UO_943 (O_943,N_9864,N_9583);
and UO_944 (O_944,N_9678,N_9880);
nand UO_945 (O_945,N_9876,N_9985);
or UO_946 (O_946,N_9721,N_9834);
and UO_947 (O_947,N_9775,N_9565);
nor UO_948 (O_948,N_9968,N_9870);
nor UO_949 (O_949,N_9589,N_9686);
or UO_950 (O_950,N_9511,N_9646);
and UO_951 (O_951,N_9976,N_9706);
or UO_952 (O_952,N_9789,N_9648);
nor UO_953 (O_953,N_9563,N_9695);
and UO_954 (O_954,N_9766,N_9539);
and UO_955 (O_955,N_9945,N_9720);
nor UO_956 (O_956,N_9747,N_9627);
nand UO_957 (O_957,N_9631,N_9812);
xnor UO_958 (O_958,N_9688,N_9833);
nor UO_959 (O_959,N_9937,N_9773);
or UO_960 (O_960,N_9970,N_9723);
nor UO_961 (O_961,N_9820,N_9571);
or UO_962 (O_962,N_9728,N_9976);
nand UO_963 (O_963,N_9654,N_9646);
nand UO_964 (O_964,N_9831,N_9773);
or UO_965 (O_965,N_9500,N_9815);
or UO_966 (O_966,N_9674,N_9859);
and UO_967 (O_967,N_9503,N_9826);
nand UO_968 (O_968,N_9825,N_9667);
nor UO_969 (O_969,N_9810,N_9797);
and UO_970 (O_970,N_9671,N_9667);
or UO_971 (O_971,N_9962,N_9784);
xnor UO_972 (O_972,N_9926,N_9678);
nor UO_973 (O_973,N_9722,N_9985);
and UO_974 (O_974,N_9608,N_9980);
nor UO_975 (O_975,N_9664,N_9592);
or UO_976 (O_976,N_9887,N_9896);
nand UO_977 (O_977,N_9540,N_9635);
nand UO_978 (O_978,N_9594,N_9842);
or UO_979 (O_979,N_9832,N_9714);
nor UO_980 (O_980,N_9923,N_9700);
and UO_981 (O_981,N_9512,N_9678);
nor UO_982 (O_982,N_9655,N_9872);
or UO_983 (O_983,N_9704,N_9615);
nor UO_984 (O_984,N_9787,N_9994);
xnor UO_985 (O_985,N_9617,N_9926);
or UO_986 (O_986,N_9532,N_9591);
and UO_987 (O_987,N_9507,N_9824);
nor UO_988 (O_988,N_9856,N_9536);
and UO_989 (O_989,N_9632,N_9989);
nand UO_990 (O_990,N_9700,N_9513);
nor UO_991 (O_991,N_9646,N_9556);
nor UO_992 (O_992,N_9702,N_9684);
nand UO_993 (O_993,N_9553,N_9700);
and UO_994 (O_994,N_9758,N_9816);
or UO_995 (O_995,N_9612,N_9961);
xor UO_996 (O_996,N_9888,N_9941);
and UO_997 (O_997,N_9974,N_9713);
or UO_998 (O_998,N_9712,N_9871);
and UO_999 (O_999,N_9726,N_9733);
xnor UO_1000 (O_1000,N_9508,N_9521);
nand UO_1001 (O_1001,N_9704,N_9719);
or UO_1002 (O_1002,N_9529,N_9772);
or UO_1003 (O_1003,N_9945,N_9815);
xor UO_1004 (O_1004,N_9586,N_9568);
or UO_1005 (O_1005,N_9500,N_9609);
nand UO_1006 (O_1006,N_9874,N_9604);
or UO_1007 (O_1007,N_9627,N_9524);
and UO_1008 (O_1008,N_9676,N_9976);
nor UO_1009 (O_1009,N_9621,N_9822);
nor UO_1010 (O_1010,N_9850,N_9703);
and UO_1011 (O_1011,N_9692,N_9837);
nand UO_1012 (O_1012,N_9591,N_9582);
xor UO_1013 (O_1013,N_9889,N_9692);
and UO_1014 (O_1014,N_9548,N_9670);
and UO_1015 (O_1015,N_9885,N_9851);
or UO_1016 (O_1016,N_9864,N_9699);
and UO_1017 (O_1017,N_9615,N_9753);
nand UO_1018 (O_1018,N_9627,N_9844);
and UO_1019 (O_1019,N_9672,N_9685);
nor UO_1020 (O_1020,N_9619,N_9879);
nand UO_1021 (O_1021,N_9628,N_9997);
or UO_1022 (O_1022,N_9561,N_9783);
or UO_1023 (O_1023,N_9628,N_9979);
and UO_1024 (O_1024,N_9584,N_9744);
and UO_1025 (O_1025,N_9895,N_9921);
and UO_1026 (O_1026,N_9849,N_9649);
and UO_1027 (O_1027,N_9624,N_9730);
nand UO_1028 (O_1028,N_9814,N_9698);
nor UO_1029 (O_1029,N_9854,N_9767);
xnor UO_1030 (O_1030,N_9501,N_9973);
and UO_1031 (O_1031,N_9680,N_9563);
or UO_1032 (O_1032,N_9946,N_9592);
nor UO_1033 (O_1033,N_9777,N_9841);
nor UO_1034 (O_1034,N_9766,N_9733);
or UO_1035 (O_1035,N_9734,N_9719);
nand UO_1036 (O_1036,N_9964,N_9517);
nand UO_1037 (O_1037,N_9697,N_9744);
and UO_1038 (O_1038,N_9700,N_9778);
or UO_1039 (O_1039,N_9662,N_9649);
or UO_1040 (O_1040,N_9881,N_9724);
or UO_1041 (O_1041,N_9619,N_9680);
and UO_1042 (O_1042,N_9552,N_9940);
nor UO_1043 (O_1043,N_9919,N_9933);
and UO_1044 (O_1044,N_9612,N_9804);
or UO_1045 (O_1045,N_9949,N_9855);
xnor UO_1046 (O_1046,N_9852,N_9820);
nor UO_1047 (O_1047,N_9599,N_9664);
or UO_1048 (O_1048,N_9856,N_9593);
xor UO_1049 (O_1049,N_9562,N_9904);
and UO_1050 (O_1050,N_9829,N_9803);
or UO_1051 (O_1051,N_9826,N_9976);
xor UO_1052 (O_1052,N_9711,N_9617);
nand UO_1053 (O_1053,N_9731,N_9808);
nand UO_1054 (O_1054,N_9701,N_9603);
nor UO_1055 (O_1055,N_9777,N_9554);
xnor UO_1056 (O_1056,N_9927,N_9560);
xnor UO_1057 (O_1057,N_9895,N_9711);
and UO_1058 (O_1058,N_9691,N_9989);
and UO_1059 (O_1059,N_9534,N_9609);
or UO_1060 (O_1060,N_9794,N_9748);
or UO_1061 (O_1061,N_9663,N_9908);
or UO_1062 (O_1062,N_9577,N_9642);
nor UO_1063 (O_1063,N_9571,N_9762);
or UO_1064 (O_1064,N_9563,N_9995);
or UO_1065 (O_1065,N_9790,N_9682);
nand UO_1066 (O_1066,N_9837,N_9812);
or UO_1067 (O_1067,N_9505,N_9643);
and UO_1068 (O_1068,N_9533,N_9964);
xor UO_1069 (O_1069,N_9875,N_9779);
and UO_1070 (O_1070,N_9858,N_9997);
xor UO_1071 (O_1071,N_9650,N_9903);
nand UO_1072 (O_1072,N_9777,N_9853);
nand UO_1073 (O_1073,N_9769,N_9733);
and UO_1074 (O_1074,N_9796,N_9703);
nand UO_1075 (O_1075,N_9669,N_9538);
nor UO_1076 (O_1076,N_9563,N_9875);
or UO_1077 (O_1077,N_9639,N_9730);
and UO_1078 (O_1078,N_9563,N_9694);
nor UO_1079 (O_1079,N_9669,N_9817);
xor UO_1080 (O_1080,N_9745,N_9699);
nand UO_1081 (O_1081,N_9906,N_9976);
nand UO_1082 (O_1082,N_9537,N_9694);
xnor UO_1083 (O_1083,N_9946,N_9649);
and UO_1084 (O_1084,N_9603,N_9526);
or UO_1085 (O_1085,N_9695,N_9761);
nand UO_1086 (O_1086,N_9717,N_9976);
nor UO_1087 (O_1087,N_9816,N_9913);
nand UO_1088 (O_1088,N_9745,N_9717);
nor UO_1089 (O_1089,N_9979,N_9662);
nor UO_1090 (O_1090,N_9832,N_9833);
xnor UO_1091 (O_1091,N_9761,N_9693);
nor UO_1092 (O_1092,N_9882,N_9848);
or UO_1093 (O_1093,N_9616,N_9862);
xnor UO_1094 (O_1094,N_9609,N_9956);
nor UO_1095 (O_1095,N_9911,N_9609);
nand UO_1096 (O_1096,N_9532,N_9964);
nand UO_1097 (O_1097,N_9546,N_9657);
or UO_1098 (O_1098,N_9950,N_9641);
nand UO_1099 (O_1099,N_9541,N_9980);
and UO_1100 (O_1100,N_9814,N_9892);
and UO_1101 (O_1101,N_9799,N_9662);
nor UO_1102 (O_1102,N_9595,N_9808);
xor UO_1103 (O_1103,N_9786,N_9767);
and UO_1104 (O_1104,N_9946,N_9795);
or UO_1105 (O_1105,N_9937,N_9990);
and UO_1106 (O_1106,N_9505,N_9983);
or UO_1107 (O_1107,N_9531,N_9909);
xor UO_1108 (O_1108,N_9953,N_9852);
nand UO_1109 (O_1109,N_9902,N_9542);
nor UO_1110 (O_1110,N_9770,N_9859);
nand UO_1111 (O_1111,N_9741,N_9696);
nor UO_1112 (O_1112,N_9912,N_9527);
nand UO_1113 (O_1113,N_9614,N_9586);
or UO_1114 (O_1114,N_9526,N_9775);
and UO_1115 (O_1115,N_9734,N_9556);
nand UO_1116 (O_1116,N_9967,N_9837);
and UO_1117 (O_1117,N_9893,N_9995);
nand UO_1118 (O_1118,N_9689,N_9605);
nor UO_1119 (O_1119,N_9616,N_9780);
nor UO_1120 (O_1120,N_9620,N_9709);
nor UO_1121 (O_1121,N_9528,N_9674);
and UO_1122 (O_1122,N_9547,N_9530);
and UO_1123 (O_1123,N_9912,N_9867);
and UO_1124 (O_1124,N_9840,N_9530);
nand UO_1125 (O_1125,N_9820,N_9951);
or UO_1126 (O_1126,N_9672,N_9618);
or UO_1127 (O_1127,N_9772,N_9603);
nand UO_1128 (O_1128,N_9699,N_9727);
or UO_1129 (O_1129,N_9821,N_9986);
and UO_1130 (O_1130,N_9578,N_9629);
or UO_1131 (O_1131,N_9507,N_9872);
or UO_1132 (O_1132,N_9871,N_9556);
and UO_1133 (O_1133,N_9730,N_9954);
and UO_1134 (O_1134,N_9902,N_9920);
nor UO_1135 (O_1135,N_9976,N_9827);
xnor UO_1136 (O_1136,N_9742,N_9619);
or UO_1137 (O_1137,N_9896,N_9777);
nand UO_1138 (O_1138,N_9993,N_9887);
nand UO_1139 (O_1139,N_9767,N_9879);
xor UO_1140 (O_1140,N_9546,N_9809);
xor UO_1141 (O_1141,N_9637,N_9779);
nand UO_1142 (O_1142,N_9626,N_9576);
nand UO_1143 (O_1143,N_9671,N_9701);
or UO_1144 (O_1144,N_9972,N_9688);
or UO_1145 (O_1145,N_9735,N_9616);
nor UO_1146 (O_1146,N_9640,N_9534);
nor UO_1147 (O_1147,N_9887,N_9839);
xnor UO_1148 (O_1148,N_9914,N_9874);
nand UO_1149 (O_1149,N_9913,N_9550);
and UO_1150 (O_1150,N_9561,N_9755);
or UO_1151 (O_1151,N_9971,N_9567);
nand UO_1152 (O_1152,N_9868,N_9604);
and UO_1153 (O_1153,N_9636,N_9980);
and UO_1154 (O_1154,N_9737,N_9889);
nor UO_1155 (O_1155,N_9564,N_9660);
nor UO_1156 (O_1156,N_9928,N_9885);
and UO_1157 (O_1157,N_9697,N_9726);
nand UO_1158 (O_1158,N_9851,N_9988);
or UO_1159 (O_1159,N_9935,N_9929);
nand UO_1160 (O_1160,N_9938,N_9751);
and UO_1161 (O_1161,N_9870,N_9716);
or UO_1162 (O_1162,N_9904,N_9518);
nand UO_1163 (O_1163,N_9994,N_9974);
nor UO_1164 (O_1164,N_9833,N_9539);
or UO_1165 (O_1165,N_9875,N_9744);
and UO_1166 (O_1166,N_9643,N_9652);
xor UO_1167 (O_1167,N_9975,N_9956);
or UO_1168 (O_1168,N_9791,N_9716);
nor UO_1169 (O_1169,N_9790,N_9806);
nand UO_1170 (O_1170,N_9638,N_9792);
or UO_1171 (O_1171,N_9663,N_9729);
or UO_1172 (O_1172,N_9803,N_9544);
and UO_1173 (O_1173,N_9728,N_9504);
and UO_1174 (O_1174,N_9676,N_9547);
or UO_1175 (O_1175,N_9900,N_9649);
and UO_1176 (O_1176,N_9629,N_9915);
and UO_1177 (O_1177,N_9974,N_9718);
or UO_1178 (O_1178,N_9724,N_9992);
nor UO_1179 (O_1179,N_9525,N_9856);
or UO_1180 (O_1180,N_9860,N_9725);
nor UO_1181 (O_1181,N_9949,N_9950);
or UO_1182 (O_1182,N_9504,N_9991);
nand UO_1183 (O_1183,N_9646,N_9742);
nand UO_1184 (O_1184,N_9947,N_9606);
and UO_1185 (O_1185,N_9854,N_9870);
and UO_1186 (O_1186,N_9559,N_9958);
or UO_1187 (O_1187,N_9801,N_9797);
nand UO_1188 (O_1188,N_9605,N_9550);
nand UO_1189 (O_1189,N_9877,N_9712);
nand UO_1190 (O_1190,N_9920,N_9731);
and UO_1191 (O_1191,N_9699,N_9650);
or UO_1192 (O_1192,N_9664,N_9667);
nand UO_1193 (O_1193,N_9861,N_9798);
nor UO_1194 (O_1194,N_9577,N_9513);
nand UO_1195 (O_1195,N_9640,N_9747);
nor UO_1196 (O_1196,N_9973,N_9792);
nor UO_1197 (O_1197,N_9750,N_9909);
nand UO_1198 (O_1198,N_9629,N_9501);
nand UO_1199 (O_1199,N_9764,N_9611);
or UO_1200 (O_1200,N_9569,N_9544);
and UO_1201 (O_1201,N_9742,N_9570);
nor UO_1202 (O_1202,N_9527,N_9517);
nand UO_1203 (O_1203,N_9633,N_9865);
or UO_1204 (O_1204,N_9792,N_9862);
nand UO_1205 (O_1205,N_9775,N_9806);
or UO_1206 (O_1206,N_9719,N_9727);
and UO_1207 (O_1207,N_9567,N_9588);
and UO_1208 (O_1208,N_9736,N_9849);
and UO_1209 (O_1209,N_9585,N_9658);
nand UO_1210 (O_1210,N_9900,N_9614);
nor UO_1211 (O_1211,N_9701,N_9904);
and UO_1212 (O_1212,N_9602,N_9622);
nand UO_1213 (O_1213,N_9725,N_9949);
xnor UO_1214 (O_1214,N_9807,N_9502);
nor UO_1215 (O_1215,N_9998,N_9672);
nand UO_1216 (O_1216,N_9805,N_9941);
nor UO_1217 (O_1217,N_9592,N_9553);
and UO_1218 (O_1218,N_9970,N_9763);
nand UO_1219 (O_1219,N_9758,N_9995);
xor UO_1220 (O_1220,N_9840,N_9772);
nand UO_1221 (O_1221,N_9840,N_9935);
or UO_1222 (O_1222,N_9678,N_9734);
nor UO_1223 (O_1223,N_9546,N_9717);
or UO_1224 (O_1224,N_9861,N_9757);
or UO_1225 (O_1225,N_9683,N_9542);
nor UO_1226 (O_1226,N_9527,N_9975);
nand UO_1227 (O_1227,N_9590,N_9738);
nor UO_1228 (O_1228,N_9987,N_9797);
and UO_1229 (O_1229,N_9894,N_9759);
nand UO_1230 (O_1230,N_9520,N_9701);
and UO_1231 (O_1231,N_9946,N_9623);
or UO_1232 (O_1232,N_9668,N_9956);
and UO_1233 (O_1233,N_9661,N_9514);
and UO_1234 (O_1234,N_9771,N_9885);
nor UO_1235 (O_1235,N_9926,N_9871);
and UO_1236 (O_1236,N_9786,N_9756);
nand UO_1237 (O_1237,N_9588,N_9939);
or UO_1238 (O_1238,N_9593,N_9819);
or UO_1239 (O_1239,N_9671,N_9720);
and UO_1240 (O_1240,N_9898,N_9686);
nor UO_1241 (O_1241,N_9889,N_9872);
or UO_1242 (O_1242,N_9771,N_9854);
or UO_1243 (O_1243,N_9608,N_9709);
nor UO_1244 (O_1244,N_9731,N_9944);
xor UO_1245 (O_1245,N_9917,N_9932);
or UO_1246 (O_1246,N_9650,N_9616);
nor UO_1247 (O_1247,N_9885,N_9788);
and UO_1248 (O_1248,N_9732,N_9780);
nor UO_1249 (O_1249,N_9889,N_9576);
nand UO_1250 (O_1250,N_9659,N_9901);
or UO_1251 (O_1251,N_9912,N_9850);
nor UO_1252 (O_1252,N_9991,N_9934);
or UO_1253 (O_1253,N_9577,N_9711);
and UO_1254 (O_1254,N_9998,N_9946);
nand UO_1255 (O_1255,N_9957,N_9799);
and UO_1256 (O_1256,N_9953,N_9710);
nand UO_1257 (O_1257,N_9513,N_9684);
and UO_1258 (O_1258,N_9939,N_9921);
nor UO_1259 (O_1259,N_9698,N_9936);
xnor UO_1260 (O_1260,N_9594,N_9758);
nor UO_1261 (O_1261,N_9656,N_9755);
and UO_1262 (O_1262,N_9939,N_9534);
xor UO_1263 (O_1263,N_9875,N_9647);
nor UO_1264 (O_1264,N_9640,N_9769);
and UO_1265 (O_1265,N_9503,N_9866);
and UO_1266 (O_1266,N_9628,N_9994);
and UO_1267 (O_1267,N_9618,N_9849);
nand UO_1268 (O_1268,N_9689,N_9778);
xnor UO_1269 (O_1269,N_9590,N_9781);
nor UO_1270 (O_1270,N_9668,N_9863);
nor UO_1271 (O_1271,N_9868,N_9738);
xnor UO_1272 (O_1272,N_9903,N_9961);
xnor UO_1273 (O_1273,N_9529,N_9783);
nand UO_1274 (O_1274,N_9867,N_9528);
and UO_1275 (O_1275,N_9628,N_9781);
nor UO_1276 (O_1276,N_9876,N_9735);
or UO_1277 (O_1277,N_9912,N_9508);
nand UO_1278 (O_1278,N_9762,N_9515);
and UO_1279 (O_1279,N_9915,N_9964);
nand UO_1280 (O_1280,N_9909,N_9803);
nand UO_1281 (O_1281,N_9546,N_9527);
and UO_1282 (O_1282,N_9588,N_9942);
or UO_1283 (O_1283,N_9897,N_9590);
nand UO_1284 (O_1284,N_9903,N_9549);
or UO_1285 (O_1285,N_9828,N_9587);
nor UO_1286 (O_1286,N_9533,N_9972);
xnor UO_1287 (O_1287,N_9859,N_9572);
nor UO_1288 (O_1288,N_9850,N_9816);
or UO_1289 (O_1289,N_9983,N_9580);
and UO_1290 (O_1290,N_9773,N_9521);
and UO_1291 (O_1291,N_9630,N_9990);
or UO_1292 (O_1292,N_9845,N_9961);
xor UO_1293 (O_1293,N_9571,N_9564);
and UO_1294 (O_1294,N_9794,N_9642);
xnor UO_1295 (O_1295,N_9507,N_9625);
xor UO_1296 (O_1296,N_9972,N_9997);
and UO_1297 (O_1297,N_9950,N_9846);
nor UO_1298 (O_1298,N_9867,N_9880);
or UO_1299 (O_1299,N_9736,N_9537);
nand UO_1300 (O_1300,N_9813,N_9887);
nor UO_1301 (O_1301,N_9979,N_9874);
nor UO_1302 (O_1302,N_9825,N_9750);
nand UO_1303 (O_1303,N_9994,N_9896);
and UO_1304 (O_1304,N_9581,N_9834);
nand UO_1305 (O_1305,N_9974,N_9964);
and UO_1306 (O_1306,N_9716,N_9983);
nor UO_1307 (O_1307,N_9600,N_9567);
nand UO_1308 (O_1308,N_9995,N_9542);
or UO_1309 (O_1309,N_9842,N_9907);
or UO_1310 (O_1310,N_9859,N_9701);
nand UO_1311 (O_1311,N_9994,N_9773);
and UO_1312 (O_1312,N_9804,N_9769);
xnor UO_1313 (O_1313,N_9702,N_9767);
nand UO_1314 (O_1314,N_9762,N_9565);
and UO_1315 (O_1315,N_9653,N_9816);
nand UO_1316 (O_1316,N_9654,N_9870);
and UO_1317 (O_1317,N_9787,N_9830);
nand UO_1318 (O_1318,N_9750,N_9764);
or UO_1319 (O_1319,N_9713,N_9970);
xnor UO_1320 (O_1320,N_9914,N_9593);
xor UO_1321 (O_1321,N_9713,N_9946);
nor UO_1322 (O_1322,N_9958,N_9636);
nand UO_1323 (O_1323,N_9574,N_9708);
and UO_1324 (O_1324,N_9852,N_9873);
and UO_1325 (O_1325,N_9570,N_9638);
xnor UO_1326 (O_1326,N_9548,N_9892);
nor UO_1327 (O_1327,N_9963,N_9753);
or UO_1328 (O_1328,N_9708,N_9965);
nor UO_1329 (O_1329,N_9645,N_9550);
or UO_1330 (O_1330,N_9856,N_9924);
nor UO_1331 (O_1331,N_9811,N_9553);
xor UO_1332 (O_1332,N_9512,N_9547);
and UO_1333 (O_1333,N_9806,N_9866);
nor UO_1334 (O_1334,N_9513,N_9950);
nand UO_1335 (O_1335,N_9534,N_9744);
and UO_1336 (O_1336,N_9579,N_9903);
nor UO_1337 (O_1337,N_9778,N_9753);
nand UO_1338 (O_1338,N_9504,N_9855);
xnor UO_1339 (O_1339,N_9994,N_9613);
and UO_1340 (O_1340,N_9621,N_9543);
or UO_1341 (O_1341,N_9590,N_9667);
xnor UO_1342 (O_1342,N_9808,N_9537);
or UO_1343 (O_1343,N_9692,N_9916);
or UO_1344 (O_1344,N_9953,N_9612);
nor UO_1345 (O_1345,N_9707,N_9821);
or UO_1346 (O_1346,N_9796,N_9818);
nand UO_1347 (O_1347,N_9645,N_9542);
or UO_1348 (O_1348,N_9936,N_9686);
nand UO_1349 (O_1349,N_9874,N_9771);
or UO_1350 (O_1350,N_9862,N_9947);
and UO_1351 (O_1351,N_9913,N_9930);
nor UO_1352 (O_1352,N_9684,N_9859);
and UO_1353 (O_1353,N_9918,N_9589);
nand UO_1354 (O_1354,N_9924,N_9512);
nand UO_1355 (O_1355,N_9639,N_9960);
nand UO_1356 (O_1356,N_9804,N_9764);
nand UO_1357 (O_1357,N_9978,N_9884);
nor UO_1358 (O_1358,N_9816,N_9977);
nand UO_1359 (O_1359,N_9884,N_9752);
nor UO_1360 (O_1360,N_9532,N_9872);
and UO_1361 (O_1361,N_9683,N_9747);
nor UO_1362 (O_1362,N_9539,N_9769);
nand UO_1363 (O_1363,N_9814,N_9666);
and UO_1364 (O_1364,N_9931,N_9835);
and UO_1365 (O_1365,N_9565,N_9885);
or UO_1366 (O_1366,N_9988,N_9500);
or UO_1367 (O_1367,N_9761,N_9923);
or UO_1368 (O_1368,N_9794,N_9665);
and UO_1369 (O_1369,N_9613,N_9756);
nand UO_1370 (O_1370,N_9807,N_9952);
xnor UO_1371 (O_1371,N_9567,N_9993);
or UO_1372 (O_1372,N_9997,N_9910);
nor UO_1373 (O_1373,N_9654,N_9892);
nand UO_1374 (O_1374,N_9723,N_9714);
nor UO_1375 (O_1375,N_9833,N_9882);
nand UO_1376 (O_1376,N_9510,N_9883);
or UO_1377 (O_1377,N_9871,N_9806);
and UO_1378 (O_1378,N_9658,N_9760);
nor UO_1379 (O_1379,N_9855,N_9684);
xor UO_1380 (O_1380,N_9643,N_9593);
and UO_1381 (O_1381,N_9712,N_9947);
nand UO_1382 (O_1382,N_9632,N_9907);
or UO_1383 (O_1383,N_9663,N_9883);
nor UO_1384 (O_1384,N_9633,N_9844);
nor UO_1385 (O_1385,N_9680,N_9637);
xor UO_1386 (O_1386,N_9570,N_9701);
nand UO_1387 (O_1387,N_9808,N_9997);
and UO_1388 (O_1388,N_9970,N_9563);
xor UO_1389 (O_1389,N_9517,N_9928);
or UO_1390 (O_1390,N_9772,N_9909);
or UO_1391 (O_1391,N_9762,N_9735);
and UO_1392 (O_1392,N_9681,N_9916);
nand UO_1393 (O_1393,N_9859,N_9831);
or UO_1394 (O_1394,N_9586,N_9913);
and UO_1395 (O_1395,N_9597,N_9898);
xnor UO_1396 (O_1396,N_9570,N_9971);
nor UO_1397 (O_1397,N_9602,N_9784);
or UO_1398 (O_1398,N_9594,N_9871);
or UO_1399 (O_1399,N_9542,N_9888);
nor UO_1400 (O_1400,N_9928,N_9688);
or UO_1401 (O_1401,N_9530,N_9599);
or UO_1402 (O_1402,N_9799,N_9512);
and UO_1403 (O_1403,N_9606,N_9608);
or UO_1404 (O_1404,N_9546,N_9697);
or UO_1405 (O_1405,N_9669,N_9866);
and UO_1406 (O_1406,N_9916,N_9913);
nand UO_1407 (O_1407,N_9693,N_9541);
or UO_1408 (O_1408,N_9779,N_9711);
xor UO_1409 (O_1409,N_9870,N_9725);
nand UO_1410 (O_1410,N_9803,N_9565);
nand UO_1411 (O_1411,N_9556,N_9512);
nand UO_1412 (O_1412,N_9703,N_9825);
nand UO_1413 (O_1413,N_9666,N_9546);
nor UO_1414 (O_1414,N_9661,N_9757);
nor UO_1415 (O_1415,N_9791,N_9598);
nor UO_1416 (O_1416,N_9873,N_9821);
xor UO_1417 (O_1417,N_9551,N_9943);
xnor UO_1418 (O_1418,N_9869,N_9516);
or UO_1419 (O_1419,N_9648,N_9863);
nand UO_1420 (O_1420,N_9722,N_9759);
or UO_1421 (O_1421,N_9883,N_9572);
nor UO_1422 (O_1422,N_9909,N_9604);
nand UO_1423 (O_1423,N_9641,N_9625);
or UO_1424 (O_1424,N_9552,N_9662);
nand UO_1425 (O_1425,N_9708,N_9926);
xnor UO_1426 (O_1426,N_9950,N_9882);
nand UO_1427 (O_1427,N_9656,N_9569);
nor UO_1428 (O_1428,N_9932,N_9803);
nor UO_1429 (O_1429,N_9767,N_9853);
nor UO_1430 (O_1430,N_9603,N_9965);
and UO_1431 (O_1431,N_9984,N_9619);
nor UO_1432 (O_1432,N_9579,N_9762);
and UO_1433 (O_1433,N_9771,N_9877);
xnor UO_1434 (O_1434,N_9655,N_9633);
and UO_1435 (O_1435,N_9587,N_9652);
nor UO_1436 (O_1436,N_9965,N_9753);
nand UO_1437 (O_1437,N_9824,N_9500);
nor UO_1438 (O_1438,N_9627,N_9827);
or UO_1439 (O_1439,N_9959,N_9744);
nand UO_1440 (O_1440,N_9849,N_9724);
xor UO_1441 (O_1441,N_9835,N_9611);
nor UO_1442 (O_1442,N_9726,N_9707);
nand UO_1443 (O_1443,N_9531,N_9923);
nor UO_1444 (O_1444,N_9611,N_9754);
nor UO_1445 (O_1445,N_9851,N_9612);
nor UO_1446 (O_1446,N_9966,N_9720);
nor UO_1447 (O_1447,N_9502,N_9750);
and UO_1448 (O_1448,N_9641,N_9936);
nor UO_1449 (O_1449,N_9790,N_9601);
and UO_1450 (O_1450,N_9650,N_9641);
nor UO_1451 (O_1451,N_9692,N_9594);
and UO_1452 (O_1452,N_9791,N_9787);
and UO_1453 (O_1453,N_9823,N_9715);
and UO_1454 (O_1454,N_9553,N_9568);
xnor UO_1455 (O_1455,N_9912,N_9951);
nand UO_1456 (O_1456,N_9724,N_9833);
nor UO_1457 (O_1457,N_9546,N_9967);
or UO_1458 (O_1458,N_9932,N_9554);
and UO_1459 (O_1459,N_9996,N_9598);
nor UO_1460 (O_1460,N_9917,N_9594);
and UO_1461 (O_1461,N_9892,N_9596);
nor UO_1462 (O_1462,N_9886,N_9786);
and UO_1463 (O_1463,N_9715,N_9701);
nor UO_1464 (O_1464,N_9810,N_9991);
nor UO_1465 (O_1465,N_9690,N_9754);
xor UO_1466 (O_1466,N_9876,N_9585);
or UO_1467 (O_1467,N_9588,N_9650);
and UO_1468 (O_1468,N_9908,N_9559);
nor UO_1469 (O_1469,N_9617,N_9671);
or UO_1470 (O_1470,N_9788,N_9641);
nor UO_1471 (O_1471,N_9537,N_9611);
or UO_1472 (O_1472,N_9618,N_9789);
nand UO_1473 (O_1473,N_9508,N_9780);
nand UO_1474 (O_1474,N_9844,N_9963);
nand UO_1475 (O_1475,N_9636,N_9624);
and UO_1476 (O_1476,N_9516,N_9552);
xnor UO_1477 (O_1477,N_9795,N_9845);
nand UO_1478 (O_1478,N_9789,N_9811);
or UO_1479 (O_1479,N_9843,N_9644);
or UO_1480 (O_1480,N_9550,N_9846);
or UO_1481 (O_1481,N_9691,N_9709);
nor UO_1482 (O_1482,N_9567,N_9654);
or UO_1483 (O_1483,N_9846,N_9833);
nor UO_1484 (O_1484,N_9583,N_9841);
xnor UO_1485 (O_1485,N_9960,N_9764);
nor UO_1486 (O_1486,N_9909,N_9748);
and UO_1487 (O_1487,N_9856,N_9738);
or UO_1488 (O_1488,N_9656,N_9666);
xnor UO_1489 (O_1489,N_9692,N_9787);
xor UO_1490 (O_1490,N_9633,N_9755);
nand UO_1491 (O_1491,N_9575,N_9815);
and UO_1492 (O_1492,N_9875,N_9996);
and UO_1493 (O_1493,N_9550,N_9725);
nor UO_1494 (O_1494,N_9549,N_9922);
and UO_1495 (O_1495,N_9838,N_9747);
and UO_1496 (O_1496,N_9513,N_9673);
nor UO_1497 (O_1497,N_9646,N_9899);
and UO_1498 (O_1498,N_9642,N_9809);
xor UO_1499 (O_1499,N_9625,N_9879);
endmodule